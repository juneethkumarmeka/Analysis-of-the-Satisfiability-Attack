module basic_2500_25000_3000_5_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
or U0 (N_0,In_2450,In_1742);
xnor U1 (N_1,In_1802,In_729);
nand U2 (N_2,In_362,In_714);
nor U3 (N_3,In_757,In_1275);
nand U4 (N_4,In_1976,In_1206);
nand U5 (N_5,In_1954,In_2264);
and U6 (N_6,In_1747,In_213);
nor U7 (N_7,In_816,In_2249);
xor U8 (N_8,In_1544,In_2011);
or U9 (N_9,In_605,In_257);
nor U10 (N_10,In_26,In_741);
or U11 (N_11,In_949,In_830);
nor U12 (N_12,In_541,In_566);
xor U13 (N_13,In_922,In_601);
nor U14 (N_14,In_774,In_1228);
xnor U15 (N_15,In_1308,In_759);
or U16 (N_16,In_1093,In_2217);
nand U17 (N_17,In_825,In_1799);
xnor U18 (N_18,In_2034,In_1555);
and U19 (N_19,In_1639,In_1651);
or U20 (N_20,In_576,In_892);
or U21 (N_21,In_701,In_1643);
nand U22 (N_22,In_323,In_241);
xnor U23 (N_23,In_1508,In_77);
and U24 (N_24,In_68,In_1444);
and U25 (N_25,In_887,In_1850);
nor U26 (N_26,In_519,In_327);
or U27 (N_27,In_48,In_2036);
and U28 (N_28,In_1609,In_2277);
and U29 (N_29,In_1195,In_1505);
xor U30 (N_30,In_2216,In_113);
xor U31 (N_31,In_509,In_764);
nand U32 (N_32,In_683,In_1718);
and U33 (N_33,In_1266,In_2395);
and U34 (N_34,In_2051,In_1709);
xnor U35 (N_35,In_1224,In_703);
and U36 (N_36,In_1983,In_2195);
nor U37 (N_37,In_1038,In_1011);
xor U38 (N_38,In_93,In_2441);
and U39 (N_39,In_2311,In_1201);
and U40 (N_40,In_2353,In_133);
nand U41 (N_41,In_2,In_1851);
or U42 (N_42,In_1236,In_85);
and U43 (N_43,In_1149,In_915);
nor U44 (N_44,In_795,In_466);
or U45 (N_45,In_1340,In_857);
xor U46 (N_46,In_98,In_219);
and U47 (N_47,In_1970,In_1288);
xnor U48 (N_48,In_211,In_754);
nor U49 (N_49,In_1830,In_1488);
xor U50 (N_50,In_2272,In_1596);
nand U51 (N_51,In_1120,In_348);
nand U52 (N_52,In_1673,In_2172);
or U53 (N_53,In_990,In_24);
or U54 (N_54,In_183,In_693);
nand U55 (N_55,In_293,In_1410);
or U56 (N_56,In_1924,In_1200);
nor U57 (N_57,In_875,In_2374);
nor U58 (N_58,In_2002,In_261);
nor U59 (N_59,In_579,In_1398);
nor U60 (N_60,In_1197,In_244);
or U61 (N_61,In_1390,In_57);
xor U62 (N_62,In_462,In_641);
and U63 (N_63,In_1600,In_2173);
and U64 (N_64,In_1392,In_2359);
nor U65 (N_65,In_518,In_1357);
and U66 (N_66,In_2267,In_1650);
and U67 (N_67,In_963,In_361);
or U68 (N_68,In_567,In_1780);
nand U69 (N_69,In_992,In_2273);
nand U70 (N_70,In_1040,In_1907);
or U71 (N_71,In_1857,In_880);
xnor U72 (N_72,In_1946,In_419);
nand U73 (N_73,In_288,In_2468);
and U74 (N_74,In_191,In_1761);
or U75 (N_75,In_2384,In_1529);
xor U76 (N_76,In_1371,In_2138);
or U77 (N_77,In_1890,In_625);
or U78 (N_78,In_1530,In_1346);
and U79 (N_79,In_2143,In_850);
nor U80 (N_80,In_1872,In_53);
nor U81 (N_81,In_1077,In_1937);
and U82 (N_82,In_2372,In_1406);
and U83 (N_83,In_2206,In_2198);
nand U84 (N_84,In_2293,In_888);
nor U85 (N_85,In_1382,In_835);
nor U86 (N_86,In_1617,In_676);
xnor U87 (N_87,In_1723,In_1743);
and U88 (N_88,In_433,In_2428);
or U89 (N_89,In_457,In_269);
and U90 (N_90,In_1625,In_2163);
nand U91 (N_91,In_1214,In_784);
or U92 (N_92,In_1817,In_2191);
or U93 (N_93,In_454,In_105);
nand U94 (N_94,In_2244,In_1549);
and U95 (N_95,In_1685,In_467);
nor U96 (N_96,In_2412,In_1668);
and U97 (N_97,In_1623,In_1364);
or U98 (N_98,In_1178,In_1283);
or U99 (N_99,In_1183,In_386);
nand U100 (N_100,In_1334,In_1328);
nor U101 (N_101,In_1130,In_1194);
nor U102 (N_102,In_1669,In_1079);
xor U103 (N_103,In_1196,In_1518);
xnor U104 (N_104,In_2453,In_672);
nor U105 (N_105,In_1582,In_588);
nand U106 (N_106,In_793,In_110);
or U107 (N_107,In_2480,In_684);
nor U108 (N_108,In_2376,In_91);
nor U109 (N_109,In_1359,In_1587);
or U110 (N_110,In_393,In_1523);
nand U111 (N_111,In_1642,In_1863);
nand U112 (N_112,In_1285,In_1873);
or U113 (N_113,In_2079,In_2477);
xor U114 (N_114,In_2368,In_414);
xor U115 (N_115,In_218,In_1867);
nand U116 (N_116,In_2303,In_2445);
and U117 (N_117,In_472,In_115);
xnor U118 (N_118,In_882,In_2120);
nor U119 (N_119,In_2177,In_2419);
nor U120 (N_120,In_432,In_125);
and U121 (N_121,In_2227,In_846);
nor U122 (N_122,In_112,In_1648);
nand U123 (N_123,In_1373,In_2078);
nand U124 (N_124,In_786,In_1785);
xor U125 (N_125,In_14,In_2127);
xor U126 (N_126,In_2461,In_2095);
nor U127 (N_127,In_1565,In_2123);
nor U128 (N_128,In_893,In_1317);
xor U129 (N_129,In_1900,In_1706);
nor U130 (N_130,In_2052,In_485);
xor U131 (N_131,In_2346,In_2306);
and U132 (N_132,In_2247,In_429);
or U133 (N_133,In_148,In_2114);
nand U134 (N_134,In_1935,In_561);
or U135 (N_135,In_1811,In_549);
nand U136 (N_136,In_2314,In_2398);
nand U137 (N_137,In_1217,In_145);
nor U138 (N_138,In_629,In_777);
nor U139 (N_139,In_985,In_814);
nor U140 (N_140,In_1633,In_33);
nor U141 (N_141,In_1855,In_411);
xnor U142 (N_142,In_2471,In_546);
nor U143 (N_143,In_1076,In_89);
nor U144 (N_144,In_1920,In_2358);
nor U145 (N_145,In_1003,In_228);
or U146 (N_146,In_917,In_1386);
or U147 (N_147,In_1672,In_488);
nor U148 (N_148,In_39,In_1240);
nand U149 (N_149,In_205,In_1984);
xor U150 (N_150,In_1828,In_688);
xnor U151 (N_151,In_1688,In_494);
and U152 (N_152,In_1979,In_1934);
and U153 (N_153,In_1923,In_40);
or U154 (N_154,In_16,In_1166);
and U155 (N_155,In_751,In_1919);
nor U156 (N_156,In_307,In_868);
and U157 (N_157,In_504,In_2084);
or U158 (N_158,In_2416,In_2141);
and U159 (N_159,In_858,In_1221);
nand U160 (N_160,In_1703,In_1414);
and U161 (N_161,In_2248,In_706);
nor U162 (N_162,In_736,In_2067);
or U163 (N_163,In_1475,In_1354);
or U164 (N_164,In_2119,In_685);
nor U165 (N_165,In_1454,In_872);
nor U166 (N_166,In_1512,In_1043);
xnor U167 (N_167,In_2048,In_2188);
nor U168 (N_168,In_1132,In_1891);
nand U169 (N_169,In_175,In_55);
or U170 (N_170,In_1961,In_132);
and U171 (N_171,In_1020,In_2109);
or U172 (N_172,In_2165,In_1594);
and U173 (N_173,In_193,In_2491);
nor U174 (N_174,In_1428,In_802);
nand U175 (N_175,In_2271,In_707);
nor U176 (N_176,In_45,In_2229);
or U177 (N_177,In_1948,In_63);
and U178 (N_178,In_568,In_438);
nand U179 (N_179,In_734,In_1628);
xnor U180 (N_180,In_294,In_920);
xor U181 (N_181,In_1306,In_324);
or U182 (N_182,In_538,In_347);
or U183 (N_183,In_2377,In_1062);
and U184 (N_184,In_11,In_1626);
nor U185 (N_185,In_130,In_1074);
and U186 (N_186,In_885,In_769);
and U187 (N_187,In_420,In_197);
nand U188 (N_188,In_1179,In_2403);
xnor U189 (N_189,In_662,In_38);
or U190 (N_190,In_746,In_726);
nand U191 (N_191,In_2014,In_713);
xnor U192 (N_192,In_96,In_21);
or U193 (N_193,In_2105,In_1035);
xnor U194 (N_194,In_2202,In_1490);
xor U195 (N_195,In_1744,In_1363);
or U196 (N_196,In_280,In_529);
and U197 (N_197,In_630,In_989);
nand U198 (N_198,In_957,In_1528);
nand U199 (N_199,In_1345,In_1289);
nor U200 (N_200,In_937,In_1615);
nor U201 (N_201,In_1165,In_574);
xor U202 (N_202,In_1586,In_221);
or U203 (N_203,In_1234,In_1491);
or U204 (N_204,In_792,In_1479);
or U205 (N_205,In_2145,In_520);
and U206 (N_206,In_1998,In_645);
or U207 (N_207,In_942,In_680);
nand U208 (N_208,In_2117,In_972);
xnor U209 (N_209,In_25,In_1932);
nor U210 (N_210,In_773,In_2423);
and U211 (N_211,In_1404,In_285);
nand U212 (N_212,In_543,In_100);
nor U213 (N_213,In_719,In_2390);
xnor U214 (N_214,In_1046,In_1696);
nand U215 (N_215,In_1975,In_603);
or U216 (N_216,In_861,In_266);
xor U217 (N_217,In_1333,In_1239);
or U218 (N_218,In_1438,In_2409);
nand U219 (N_219,In_891,In_691);
or U220 (N_220,In_712,In_1805);
xnor U221 (N_221,In_2486,In_1313);
and U222 (N_222,In_260,In_2396);
or U223 (N_223,In_497,In_1350);
xnor U224 (N_224,In_1945,In_10);
and U225 (N_225,In_1142,In_818);
and U226 (N_226,In_2467,In_1848);
or U227 (N_227,In_1699,In_1492);
nor U228 (N_228,In_345,In_901);
and U229 (N_229,In_550,In_560);
nor U230 (N_230,In_441,In_335);
and U231 (N_231,In_514,In_916);
nand U232 (N_232,In_1847,In_1692);
or U233 (N_233,In_2268,In_1520);
nor U234 (N_234,In_1409,In_614);
xnor U235 (N_235,In_918,In_2347);
nor U236 (N_236,In_945,In_290);
nand U237 (N_237,In_2493,In_154);
nor U238 (N_238,In_2252,In_1816);
xor U239 (N_239,In_2386,In_246);
xor U240 (N_240,In_116,In_1792);
nor U241 (N_241,In_1424,In_1790);
xnor U242 (N_242,In_1487,In_1383);
and U243 (N_243,In_364,In_1127);
nand U244 (N_244,In_2193,In_2410);
nor U245 (N_245,In_2285,In_1379);
or U246 (N_246,In_461,In_785);
xnor U247 (N_247,In_1049,In_1112);
nor U248 (N_248,In_1052,In_140);
xor U249 (N_249,In_1061,In_416);
and U250 (N_250,In_167,In_1230);
nand U251 (N_251,In_1418,In_1547);
and U252 (N_252,In_1461,In_6);
nand U253 (N_253,In_286,In_1331);
nor U254 (N_254,In_2381,In_1389);
nor U255 (N_255,In_681,In_1366);
and U256 (N_256,In_632,In_863);
xnor U257 (N_257,In_2054,In_2464);
or U258 (N_258,In_1676,In_813);
nor U259 (N_259,In_1930,In_1813);
and U260 (N_260,In_2475,In_1644);
nand U261 (N_261,In_117,In_770);
and U262 (N_262,In_1941,In_1420);
nand U263 (N_263,In_589,In_1353);
xnor U264 (N_264,In_995,In_2380);
nand U265 (N_265,In_476,In_2402);
nor U266 (N_266,In_2253,In_1577);
or U267 (N_267,In_512,In_1874);
and U268 (N_268,In_801,In_1798);
and U269 (N_269,In_2434,In_849);
and U270 (N_270,In_2135,In_1808);
and U271 (N_271,In_1395,In_1169);
nor U272 (N_272,In_1322,In_725);
and U273 (N_273,In_1750,In_1771);
and U274 (N_274,In_106,In_400);
or U275 (N_275,In_1121,In_297);
and U276 (N_276,In_1116,In_1304);
nand U277 (N_277,In_1645,In_2379);
nand U278 (N_278,In_1636,In_2016);
and U279 (N_279,In_1796,In_1015);
or U280 (N_280,In_296,In_1909);
and U281 (N_281,In_1307,In_1327);
nor U282 (N_282,In_1219,In_161);
and U283 (N_283,In_1952,In_1903);
or U284 (N_284,In_960,In_1784);
or U285 (N_285,In_2334,In_231);
xnor U286 (N_286,In_227,In_1341);
or U287 (N_287,In_388,In_1012);
and U288 (N_288,In_368,In_745);
nor U289 (N_289,In_1926,In_1002);
xor U290 (N_290,In_377,In_1287);
nor U291 (N_291,In_1233,In_2137);
nor U292 (N_292,In_1232,In_483);
xnor U293 (N_293,In_1377,In_337);
and U294 (N_294,In_1971,In_2487);
or U295 (N_295,In_146,In_2481);
xnor U296 (N_296,In_958,In_690);
nand U297 (N_297,In_2019,In_1325);
and U298 (N_298,In_908,In_203);
and U299 (N_299,In_253,In_1474);
xnor U300 (N_300,In_1362,In_1978);
nand U301 (N_301,In_2199,In_1385);
nor U302 (N_302,In_1915,In_1447);
and U303 (N_303,In_1731,In_934);
xnor U304 (N_304,In_1078,In_1211);
xor U305 (N_305,In_607,In_940);
or U306 (N_306,In_1963,In_1494);
or U307 (N_307,In_310,In_619);
nor U308 (N_308,In_84,In_2088);
and U309 (N_309,In_1955,In_2363);
and U310 (N_310,In_1527,In_2460);
xnor U311 (N_311,In_1768,In_178);
or U312 (N_312,In_2013,In_446);
nand U313 (N_313,In_2157,In_422);
xnor U314 (N_314,In_1734,In_982);
nand U315 (N_315,In_2077,In_954);
xnor U316 (N_316,In_1973,In_1203);
or U317 (N_317,In_637,In_845);
xnor U318 (N_318,In_914,In_111);
nor U319 (N_319,In_356,In_141);
and U320 (N_320,In_836,In_1571);
nand U321 (N_321,In_363,In_1167);
and U322 (N_322,In_182,In_698);
xnor U323 (N_323,In_679,In_2415);
xor U324 (N_324,In_1683,In_156);
and U325 (N_325,In_598,In_1212);
nand U326 (N_326,In_372,In_1028);
nand U327 (N_327,In_824,In_1870);
nor U328 (N_328,In_181,In_762);
nor U329 (N_329,In_1007,In_1421);
and U330 (N_330,In_2276,In_128);
and U331 (N_331,In_1913,In_41);
nand U332 (N_332,In_613,In_2443);
or U333 (N_333,In_1517,In_1425);
xor U334 (N_334,In_2295,In_235);
nor U335 (N_335,In_2394,In_750);
xor U336 (N_336,In_1122,In_275);
nand U337 (N_337,In_1966,In_1177);
xnor U338 (N_338,In_43,In_354);
nand U339 (N_339,In_2254,In_1831);
nor U340 (N_340,In_249,In_1301);
or U341 (N_341,In_2329,In_710);
nand U342 (N_342,In_2178,In_2160);
and U343 (N_343,In_1807,In_1837);
xor U344 (N_344,In_522,In_1752);
nand U345 (N_345,In_239,In_2087);
and U346 (N_346,In_90,In_1423);
nor U347 (N_347,In_951,In_2166);
nor U348 (N_348,In_447,In_1767);
and U349 (N_349,In_2495,In_2404);
or U350 (N_350,In_176,In_12);
and U351 (N_351,In_1982,In_212);
nor U352 (N_352,In_610,In_597);
and U353 (N_353,In_932,In_1439);
xnor U354 (N_354,In_187,In_1158);
xor U355 (N_355,In_991,In_256);
or U356 (N_356,In_1916,In_2232);
xor U357 (N_357,In_1845,In_217);
xnor U358 (N_358,In_2071,In_1455);
and U359 (N_359,In_596,In_646);
nand U360 (N_360,In_1336,In_1069);
or U361 (N_361,In_240,In_1562);
xnor U362 (N_362,In_1724,In_964);
xnor U363 (N_363,In_2008,In_548);
xor U364 (N_364,In_1290,In_1931);
or U365 (N_365,In_2065,In_775);
nor U366 (N_366,In_1272,In_1801);
and U367 (N_367,In_1575,In_1921);
or U368 (N_368,In_1170,In_314);
xnor U369 (N_369,In_649,In_81);
or U370 (N_370,In_318,In_552);
or U371 (N_371,In_427,In_1381);
xor U372 (N_372,In_974,In_1564);
nor U373 (N_373,In_544,In_97);
nor U374 (N_374,In_484,In_2148);
or U375 (N_375,In_1021,In_209);
nand U376 (N_376,In_1933,In_1044);
xor U377 (N_377,In_190,In_2279);
and U378 (N_378,In_2239,In_2357);
or U379 (N_379,In_1297,In_58);
nand U380 (N_380,In_907,In_540);
nor U381 (N_381,In_1879,In_413);
and U382 (N_382,In_841,In_352);
nor U383 (N_383,In_1893,In_925);
nand U384 (N_384,In_826,In_1720);
xnor U385 (N_385,In_1260,In_1251);
or U386 (N_386,In_2497,In_559);
nand U387 (N_387,In_2341,In_696);
nor U388 (N_388,In_1431,In_1400);
nor U389 (N_389,In_1841,In_1281);
and U390 (N_390,In_709,In_2282);
nor U391 (N_391,In_1852,In_2305);
nor U392 (N_392,In_1795,In_501);
nor U393 (N_393,In_933,In_2061);
nand U394 (N_394,In_1186,In_2124);
nor U395 (N_395,In_22,In_2496);
or U396 (N_396,In_502,In_1789);
or U397 (N_397,In_636,In_1188);
or U398 (N_398,In_2458,In_1519);
xnor U399 (N_399,In_1499,In_2122);
xnor U400 (N_400,In_19,In_439);
and U401 (N_401,In_643,In_262);
and U402 (N_402,In_34,In_1988);
or U403 (N_403,In_2144,In_2125);
xor U404 (N_404,In_1717,In_2287);
and U405 (N_405,In_2197,In_967);
nor U406 (N_406,In_810,In_1180);
or U407 (N_407,In_234,In_358);
nand U408 (N_408,In_1993,In_15);
nor U409 (N_409,In_749,In_1888);
nor U410 (N_410,In_947,In_2243);
xor U411 (N_411,In_1257,In_2236);
or U412 (N_412,In_1119,In_2366);
or U413 (N_413,In_1638,In_1883);
nand U414 (N_414,In_2047,In_465);
and U415 (N_415,In_367,In_69);
or U416 (N_416,In_900,In_1991);
and U417 (N_417,In_946,In_399);
nand U418 (N_418,In_2397,In_723);
xor U419 (N_419,In_1840,In_1738);
xnor U420 (N_420,In_1820,In_1225);
nor U421 (N_421,In_1791,In_778);
nand U422 (N_422,In_886,In_64);
nand U423 (N_423,In_304,In_2203);
nor U424 (N_424,In_2399,In_245);
and U425 (N_425,In_50,In_51);
and U426 (N_426,In_2133,In_1509);
and U427 (N_427,In_1522,In_1176);
nor U428 (N_428,In_927,In_1774);
and U429 (N_429,In_2213,In_1205);
xor U430 (N_430,In_49,In_1797);
and U431 (N_431,In_1819,In_254);
and U432 (N_432,In_1548,In_404);
xnor U433 (N_433,In_1110,In_1370);
nor U434 (N_434,In_1656,In_1640);
nor U435 (N_435,In_620,In_1678);
nor U436 (N_436,In_1846,In_1);
nor U437 (N_437,In_1449,In_1779);
or U438 (N_438,In_1315,In_491);
xor U439 (N_439,In_1143,In_1770);
and U440 (N_440,In_1442,In_2275);
and U441 (N_441,In_1914,In_2288);
and U442 (N_442,In_401,In_226);
nor U443 (N_443,In_2308,In_1254);
nand U444 (N_444,In_788,In_1472);
and U445 (N_445,In_87,In_2092);
or U446 (N_446,In_73,In_101);
and U447 (N_447,In_1099,In_1606);
and U448 (N_448,In_1017,In_2332);
and U449 (N_449,In_2089,In_1605);
nor U450 (N_450,In_2161,In_2129);
or U451 (N_451,In_44,In_525);
or U452 (N_452,In_2192,In_135);
nor U453 (N_453,In_744,In_1375);
nand U454 (N_454,In_27,In_66);
or U455 (N_455,In_2324,In_1632);
or U456 (N_456,In_2041,In_1545);
xor U457 (N_457,In_1405,In_1960);
xnor U458 (N_458,In_626,In_811);
nor U459 (N_459,In_1125,In_1515);
nor U460 (N_460,In_374,In_1726);
xor U461 (N_461,In_761,In_445);
nor U462 (N_462,In_1433,In_1860);
xnor U463 (N_463,In_1759,In_1056);
or U464 (N_464,In_2167,In_1469);
xnor U465 (N_465,In_2302,In_1026);
xor U466 (N_466,In_2436,In_371);
and U467 (N_467,In_1560,In_1838);
xnor U468 (N_468,In_196,In_516);
xnor U469 (N_469,In_1235,In_107);
nor U470 (N_470,In_944,In_896);
nor U471 (N_471,In_155,In_1653);
xnor U472 (N_472,In_578,In_1990);
or U473 (N_473,In_606,In_171);
xor U474 (N_474,In_1607,In_1507);
xor U475 (N_475,In_1446,In_1621);
or U476 (N_476,In_1708,In_539);
nand U477 (N_477,In_1342,In_2291);
nor U478 (N_478,In_1160,In_1013);
and U479 (N_479,In_201,In_1552);
or U480 (N_480,In_558,In_798);
or U481 (N_481,In_1980,In_265);
nor U482 (N_482,In_1063,In_585);
or U483 (N_483,In_2246,In_1922);
xor U484 (N_484,In_2000,In_1065);
nand U485 (N_485,In_640,In_527);
or U486 (N_486,In_71,In_547);
xor U487 (N_487,In_418,In_966);
nand U488 (N_488,In_263,In_1713);
and U489 (N_489,In_536,In_2345);
xor U490 (N_490,In_1686,In_2435);
and U491 (N_491,In_122,In_134);
nor U492 (N_492,In_2074,In_1725);
or U493 (N_493,In_317,In_1256);
or U494 (N_494,In_981,In_1153);
nor U495 (N_495,In_2184,In_631);
xnor U496 (N_496,In_1016,In_2083);
nor U497 (N_497,In_36,In_392);
and U498 (N_498,In_847,In_76);
nand U499 (N_499,In_2024,In_837);
nand U500 (N_500,In_748,In_2297);
xnor U501 (N_501,In_657,In_1352);
and U502 (N_502,In_20,In_2489);
or U503 (N_503,In_531,In_1557);
and U504 (N_504,In_2111,In_387);
or U505 (N_505,In_1070,In_1493);
and U506 (N_506,In_2100,In_852);
xor U507 (N_507,In_1175,In_1977);
xor U508 (N_508,In_1458,In_31);
nor U509 (N_509,In_573,In_650);
xor U510 (N_510,In_862,In_1159);
nand U511 (N_511,In_2220,In_486);
xor U512 (N_512,In_385,In_2454);
nand U513 (N_513,In_2010,In_2408);
or U514 (N_514,In_840,In_1111);
and U515 (N_515,In_2375,In_2281);
xnor U516 (N_516,In_2072,In_1733);
or U517 (N_517,In_1361,In_1674);
nand U518 (N_518,In_586,In_274);
or U519 (N_519,In_984,In_1427);
nor U520 (N_520,In_870,In_2286);
and U521 (N_521,In_664,In_1876);
nand U522 (N_522,In_2201,In_0);
nor U523 (N_523,In_131,In_102);
and U524 (N_524,In_2060,In_833);
nor U525 (N_525,In_2164,In_517);
or U526 (N_526,In_479,In_1721);
nand U527 (N_527,In_2361,In_1113);
nand U528 (N_528,In_1652,In_2262);
or U529 (N_529,In_587,In_551);
and U530 (N_530,In_123,In_407);
and U531 (N_531,In_634,In_879);
nand U532 (N_532,In_2230,In_1343);
or U533 (N_533,In_435,In_332);
nor U534 (N_534,In_943,In_1800);
or U535 (N_535,In_1154,In_1858);
and U536 (N_536,In_1868,In_1314);
and U537 (N_537,In_2270,In_424);
and U538 (N_538,In_628,In_1220);
or U539 (N_539,In_236,In_738);
nor U540 (N_540,In_2371,In_2225);
xnor U541 (N_541,In_2266,In_2320);
nand U542 (N_542,In_1332,In_1402);
and U543 (N_543,In_1525,In_215);
nor U544 (N_544,In_1193,In_1263);
xnor U545 (N_545,In_464,In_1880);
nand U546 (N_546,In_584,In_1292);
nand U547 (N_547,In_881,In_794);
and U548 (N_548,In_1746,In_2106);
and U549 (N_549,In_88,In_2170);
xor U550 (N_550,In_200,In_1722);
xor U551 (N_551,In_8,In_866);
and U552 (N_552,In_1511,In_765);
nand U553 (N_553,In_1698,In_987);
xor U554 (N_554,In_287,In_2007);
xor U555 (N_555,In_214,In_1054);
nand U556 (N_556,In_306,In_1546);
nor U557 (N_557,In_2231,In_17);
nor U558 (N_558,In_1660,In_415);
xnor U559 (N_559,In_1441,In_2037);
nand U560 (N_560,In_1451,In_295);
nor U561 (N_561,In_1215,In_2049);
nand U562 (N_562,In_815,In_1115);
xor U563 (N_563,In_1965,In_61);
and U564 (N_564,In_160,In_475);
xnor U565 (N_565,In_2090,In_1483);
nor U566 (N_566,In_1702,In_860);
nand U567 (N_567,In_997,In_1574);
nor U568 (N_568,In_1700,In_1209);
and U569 (N_569,In_819,In_232);
nand U570 (N_570,In_37,In_577);
or U571 (N_571,In_2301,In_1255);
and U572 (N_572,In_1773,In_149);
nor U573 (N_573,In_158,In_1267);
and U574 (N_574,In_2278,In_812);
or U575 (N_575,In_1906,In_790);
and U576 (N_576,In_1925,In_2330);
nor U577 (N_577,In_2070,In_1008);
or U578 (N_578,In_654,In_2499);
nor U579 (N_579,In_611,In_1391);
nor U580 (N_580,In_2098,In_2068);
nand U581 (N_581,In_2257,In_452);
nor U582 (N_582,In_2029,In_2001);
or U583 (N_583,In_1413,In_1897);
or U584 (N_584,In_1495,In_78);
or U585 (N_585,In_594,In_909);
xor U586 (N_586,In_903,In_394);
xnor U587 (N_587,In_2128,In_699);
xor U588 (N_588,In_1677,In_2452);
xnor U589 (N_589,In_682,In_5);
nand U590 (N_590,In_2189,In_1202);
nor U591 (N_591,In_988,In_2112);
or U592 (N_592,In_18,In_460);
nor U593 (N_593,In_1681,In_1904);
and U594 (N_594,In_557,In_204);
or U595 (N_595,In_2073,In_1419);
xor U596 (N_596,In_2490,In_1465);
nand U597 (N_597,In_397,In_272);
and U598 (N_598,In_883,In_1460);
nor U599 (N_599,In_1611,In_308);
nand U600 (N_600,In_1995,In_2028);
xor U601 (N_601,In_2099,In_1140);
xnor U602 (N_602,In_1622,In_2082);
or U603 (N_603,In_855,In_1558);
nand U604 (N_604,In_692,In_1503);
nand U605 (N_605,In_1736,In_339);
nor U606 (N_606,In_13,In_2044);
or U607 (N_607,In_1189,In_1550);
nor U608 (N_608,In_456,In_137);
xnor U609 (N_609,In_2298,In_177);
nor U610 (N_610,In_2113,In_869);
or U611 (N_611,In_329,In_1023);
nor U612 (N_612,In_1348,In_1060);
xnor U613 (N_613,In_1156,In_1612);
nand U614 (N_614,In_1905,In_2317);
nor U615 (N_615,In_521,In_583);
and U616 (N_616,In_1136,In_59);
xnor U617 (N_617,In_2440,In_2261);
and U618 (N_618,In_1833,In_581);
xor U619 (N_619,In_2056,In_2414);
or U620 (N_620,In_2043,In_526);
nand U621 (N_621,In_838,In_2233);
and U622 (N_622,In_671,In_1630);
nand U623 (N_623,In_609,In_384);
nor U624 (N_624,In_931,In_398);
xnor U625 (N_625,In_2406,In_499);
nor U626 (N_626,In_189,In_854);
and U627 (N_627,In_1655,In_1765);
nand U628 (N_628,In_350,In_1000);
or U629 (N_629,In_804,In_1786);
or U630 (N_630,In_638,In_1397);
xor U631 (N_631,In_542,In_1707);
nand U632 (N_632,In_1032,In_1432);
nor U633 (N_633,In_1243,In_360);
or U634 (N_634,In_2096,In_35);
xnor U635 (N_635,In_1351,In_768);
xnor U636 (N_636,In_1729,In_42);
nand U637 (N_637,In_1714,In_1942);
or U638 (N_638,In_440,In_2430);
nand U639 (N_639,In_2492,In_2149);
and U640 (N_640,In_174,In_1252);
or U641 (N_641,In_562,In_1080);
or U642 (N_642,In_1665,In_2299);
nor U643 (N_643,In_2063,In_1064);
xnor U644 (N_644,In_2064,In_2449);
nand U645 (N_645,In_771,In_975);
nand U646 (N_646,In_2026,In_2108);
nor U647 (N_647,In_1981,In_259);
nand U648 (N_648,In_720,In_1335);
or U649 (N_649,In_575,In_663);
nand U650 (N_650,In_1462,In_496);
xnor U651 (N_651,In_1782,In_2457);
or U652 (N_652,In_165,In_1992);
and U653 (N_653,In_1881,In_2405);
and U654 (N_654,In_1697,In_1477);
xor U655 (N_655,In_142,In_1075);
and U656 (N_656,In_2355,In_1101);
nand U657 (N_657,In_781,In_1486);
xnor U658 (N_658,In_2018,In_647);
or U659 (N_659,In_642,In_1889);
xor U660 (N_660,In_570,In_342);
and U661 (N_661,In_599,In_1603);
nand U662 (N_662,In_1705,In_1827);
xnor U663 (N_663,In_2140,In_279);
or U664 (N_664,In_1962,In_2290);
nand U665 (N_665,In_1242,In_1886);
nor U666 (N_666,In_1027,In_92);
xnor U667 (N_667,In_1053,In_406);
nand U668 (N_668,In_528,In_1741);
and U669 (N_669,In_1055,In_1355);
nand U670 (N_670,In_1730,In_1208);
or U671 (N_671,In_1299,In_1001);
nor U672 (N_672,In_1399,In_180);
xnor U673 (N_673,In_844,In_1098);
nor U674 (N_674,In_1986,In_1809);
xor U675 (N_675,In_1854,In_1666);
nand U676 (N_676,In_299,In_1794);
nand U677 (N_677,In_2182,In_2316);
nor U678 (N_678,In_1309,In_2318);
and U679 (N_679,In_1776,In_1745);
or U680 (N_680,In_1936,In_492);
and U681 (N_681,In_1300,In_506);
xor U682 (N_682,In_2319,In_264);
or U683 (N_683,In_463,In_302);
nor U684 (N_684,In_1658,In_978);
xor U685 (N_685,In_2351,In_2085);
or U686 (N_686,In_1237,In_569);
nor U687 (N_687,In_1513,In_979);
or U688 (N_688,In_1259,In_722);
nor U689 (N_689,In_2035,In_1539);
or U690 (N_690,In_1155,In_1265);
nor U691 (N_691,In_878,In_1661);
or U692 (N_692,In_732,In_1105);
and U693 (N_693,In_1619,In_248);
nand U694 (N_694,In_147,In_1277);
nand U695 (N_695,In_1629,In_67);
nor U696 (N_696,In_2142,In_402);
nor U697 (N_697,In_172,In_1748);
nor U698 (N_698,In_1740,In_2205);
and U699 (N_699,In_2331,In_2327);
xnor U700 (N_700,In_482,In_1663);
nand U701 (N_701,In_1985,In_1394);
nor U702 (N_702,In_513,In_2210);
nor U703 (N_703,In_2367,In_242);
or U704 (N_704,In_2446,In_1103);
xnor U705 (N_705,In_939,In_998);
xor U706 (N_706,In_1559,In_952);
nand U707 (N_707,In_1504,In_1553);
nand U708 (N_708,In_1092,In_1368);
and U709 (N_709,In_1590,In_1566);
and U710 (N_710,In_508,In_1403);
xor U711 (N_711,In_772,In_1261);
nand U712 (N_712,In_2228,In_1911);
or U713 (N_713,In_1089,In_1387);
or U714 (N_714,In_62,In_1216);
or U715 (N_715,In_129,In_1133);
nor U716 (N_716,In_2283,In_623);
xor U717 (N_717,In_791,In_592);
nor U718 (N_718,In_52,In_1510);
nand U719 (N_719,In_756,In_853);
nor U720 (N_720,In_1452,In_1249);
and U721 (N_721,In_29,In_2168);
or U722 (N_722,In_498,In_595);
and U723 (N_723,In_1181,In_1100);
xor U724 (N_724,In_1554,In_1601);
nand U725 (N_725,In_1269,In_1887);
xnor U726 (N_726,In_2240,In_436);
or U727 (N_727,In_291,In_206);
nor U728 (N_728,In_633,In_627);
xnor U729 (N_729,In_2433,In_806);
or U730 (N_730,In_468,In_2315);
and U731 (N_731,In_715,In_1464);
or U732 (N_732,In_994,In_103);
nand U733 (N_733,In_571,In_28);
nand U734 (N_734,In_251,In_2159);
xor U735 (N_735,In_1614,In_1949);
or U736 (N_736,In_328,In_1781);
nor U737 (N_737,In_2066,In_1572);
nor U738 (N_738,In_1329,In_223);
nor U739 (N_739,In_1457,In_1576);
or U740 (N_740,In_969,In_152);
nand U741 (N_741,In_1592,In_379);
nor U742 (N_742,In_2343,In_2350);
nand U743 (N_743,In_1047,In_1408);
nand U744 (N_744,In_1597,In_1124);
or U745 (N_745,In_1088,In_1164);
and U746 (N_746,In_1320,In_1019);
nor U747 (N_747,In_839,In_2218);
nand U748 (N_748,In_877,In_1271);
xnor U749 (N_749,In_2420,In_686);
xnor U750 (N_750,In_807,In_1241);
or U751 (N_751,In_1938,In_1727);
xnor U752 (N_752,In_1861,In_1689);
or U753 (N_753,In_2494,In_104);
nor U754 (N_754,In_1139,In_1839);
nand U755 (N_755,In_505,In_648);
nor U756 (N_756,In_2321,In_2265);
or U757 (N_757,In_1453,In_2190);
or U758 (N_758,In_495,In_383);
nand U759 (N_759,In_2259,In_1940);
and U760 (N_760,In_1033,In_1258);
nand U761 (N_761,In_1997,In_1066);
or U762 (N_762,In_1969,In_340);
nor U763 (N_763,In_1579,In_1687);
xnor U764 (N_764,In_2158,In_2333);
xor U765 (N_765,In_2059,In_1072);
or U766 (N_766,In_2115,In_1303);
nor U767 (N_767,In_2365,In_2344);
xor U768 (N_768,In_1174,In_2176);
or U769 (N_769,In_2004,In_1567);
xor U770 (N_770,In_1144,In_2296);
or U771 (N_771,In_1025,In_1593);
or U772 (N_772,In_1859,In_7);
or U773 (N_773,In_1635,In_1624);
xor U774 (N_774,In_507,In_1018);
or U775 (N_775,In_1456,In_250);
and U776 (N_776,In_1095,In_1608);
nor U777 (N_777,In_2050,In_1532);
xor U778 (N_778,In_2221,In_1134);
nand U779 (N_779,In_298,In_1245);
nor U780 (N_780,In_1864,In_624);
xnor U781 (N_781,In_1824,In_338);
or U782 (N_782,In_895,In_678);
nand U783 (N_783,In_1030,In_2241);
or U784 (N_784,In_1102,In_1369);
nor U785 (N_785,In_941,In_556);
nand U786 (N_786,In_1561,In_2223);
nand U787 (N_787,In_1022,In_913);
xnor U788 (N_788,In_2300,In_1616);
xor U789 (N_789,In_735,In_890);
xor U790 (N_790,In_238,In_1885);
xnor U791 (N_791,In_2472,In_351);
or U792 (N_792,In_935,In_1246);
nor U793 (N_793,In_1291,In_1803);
or U794 (N_794,In_2094,In_1146);
or U795 (N_795,In_1264,In_1953);
xnor U796 (N_796,In_2101,In_1106);
or U797 (N_797,In_2455,In_904);
xor U798 (N_798,In_2187,In_1145);
nor U799 (N_799,In_316,In_2183);
nor U800 (N_800,In_448,In_277);
and U801 (N_801,In_898,In_1536);
and U802 (N_802,In_1484,In_1360);
xnor U803 (N_803,In_79,In_382);
nand U804 (N_804,In_822,In_1280);
nand U805 (N_805,In_1701,In_1766);
nor U806 (N_806,In_1832,In_1711);
nand U807 (N_807,In_1126,In_805);
nand U808 (N_808,In_1478,In_1467);
nand U809 (N_809,In_2479,In_2269);
xor U810 (N_810,In_1866,In_186);
and U811 (N_811,In_1434,In_1436);
and U812 (N_812,In_2107,In_412);
or U813 (N_813,In_2057,In_1910);
or U814 (N_814,In_2425,In_2258);
nand U815 (N_815,In_1463,In_602);
and U816 (N_816,In_2383,In_473);
and U817 (N_817,In_2046,In_188);
or U818 (N_818,In_1210,In_1118);
nand U819 (N_819,In_2407,In_1367);
nand U820 (N_820,In_355,In_1048);
nor U821 (N_821,In_2153,In_851);
nand U822 (N_822,In_1637,In_1244);
or U823 (N_823,In_2304,In_1094);
nand U824 (N_824,In_1849,In_313);
and U825 (N_825,In_1422,In_1540);
or U826 (N_826,In_2292,In_2103);
nand U827 (N_827,In_535,In_2069);
and U828 (N_828,In_616,In_593);
nand U829 (N_829,In_1305,In_1892);
or U830 (N_830,In_843,In_899);
nor U831 (N_831,In_2476,In_2130);
xor U832 (N_832,In_1598,In_1059);
nor U833 (N_833,In_391,In_2250);
or U834 (N_834,In_1757,In_948);
nand U835 (N_835,In_333,In_2200);
xor U836 (N_836,In_1199,In_2309);
nand U837 (N_837,In_126,In_243);
xor U838 (N_838,In_2017,In_1222);
nand U839 (N_839,In_1295,In_1514);
nand U840 (N_840,In_500,In_1396);
nand U841 (N_841,In_1631,In_1950);
nor U842 (N_842,In_2055,In_1667);
nand U843 (N_843,In_1337,In_553);
xor U844 (N_844,In_82,In_2474);
and U845 (N_845,In_192,In_1818);
nor U846 (N_846,In_1378,In_2025);
xnor U847 (N_847,In_2020,In_687);
xor U848 (N_848,In_4,In_1671);
nor U849 (N_849,In_1204,In_827);
xnor U850 (N_850,In_2023,In_1108);
or U851 (N_851,In_320,In_2062);
xnor U852 (N_852,In_1213,In_1131);
nand U853 (N_853,In_554,In_1569);
nor U854 (N_854,In_2473,In_1675);
or U855 (N_855,In_2485,In_1836);
and U856 (N_856,In_1737,In_622);
or U857 (N_857,In_480,In_831);
nor U858 (N_858,In_2369,In_1627);
xor U859 (N_859,In_2370,In_1450);
xor U860 (N_860,In_1589,In_936);
nor U861 (N_861,In_255,In_1783);
and U862 (N_862,In_1247,In_859);
nand U863 (N_863,In_1031,In_470);
and U864 (N_864,In_390,In_1182);
nand U865 (N_865,In_271,In_163);
and U866 (N_866,In_704,In_2389);
and U867 (N_867,In_1412,In_1282);
or U868 (N_868,In_580,In_2427);
or U869 (N_869,In_740,In_1989);
or U870 (N_870,In_1647,In_237);
xor U871 (N_871,In_1939,In_1943);
nand U872 (N_872,In_996,In_343);
and U873 (N_873,In_2180,In_1273);
and U874 (N_874,In_797,In_767);
xnor U875 (N_875,In_151,In_871);
or U876 (N_876,In_747,In_537);
nand U877 (N_877,In_670,In_1429);
xnor U878 (N_878,In_1326,In_1968);
nand U879 (N_879,In_1613,In_2208);
or U880 (N_880,In_1497,In_1058);
nand U881 (N_881,In_1591,In_1097);
or U882 (N_882,In_565,In_1944);
xor U883 (N_883,In_760,In_1763);
nor U884 (N_884,In_2326,In_1401);
xor U885 (N_885,In_1664,In_1679);
and U886 (N_886,In_1957,In_1481);
and U887 (N_887,In_1086,In_897);
and U888 (N_888,In_2132,In_2097);
nand U889 (N_889,In_72,In_222);
nand U890 (N_890,In_2356,In_65);
and U891 (N_891,In_1037,In_658);
xor U892 (N_892,In_1253,In_832);
xor U893 (N_893,In_1999,In_1821);
nand U894 (N_894,In_2393,In_1151);
or U895 (N_895,In_1231,In_341);
xnor U896 (N_896,In_873,In_2139);
nand U897 (N_897,In_2147,In_1083);
or U898 (N_898,In_208,In_2134);
nor U899 (N_899,In_2352,In_673);
nand U900 (N_900,In_1764,In_2245);
nor U901 (N_901,In_1042,In_258);
xnor U902 (N_902,In_2151,In_799);
and U903 (N_903,In_1476,In_2451);
or U904 (N_904,In_1620,In_1471);
xnor U905 (N_905,In_405,In_2042);
xnor U906 (N_906,In_373,In_1695);
xor U907 (N_907,In_2186,In_162);
or U908 (N_908,In_1416,In_910);
xnor U909 (N_909,In_442,In_1715);
or U910 (N_910,In_1787,In_1440);
xor U911 (N_911,In_2448,In_1073);
xnor U912 (N_912,In_2310,In_1091);
nor U913 (N_913,In_1485,In_1610);
and U914 (N_914,In_2006,In_2162);
xnor U915 (N_915,In_2126,In_1223);
or U916 (N_916,In_2469,In_1349);
and U917 (N_917,In_656,In_1339);
xnor U918 (N_918,In_1344,In_1769);
nor U919 (N_919,In_555,In_166);
and U920 (N_920,In_1312,In_301);
or U921 (N_921,In_344,In_1762);
and U922 (N_922,In_635,In_1284);
and U923 (N_923,In_428,In_1583);
xor U924 (N_924,In_207,In_2021);
nand U925 (N_925,In_2385,In_2378);
or U926 (N_926,In_119,In_1229);
or U927 (N_927,In_1959,In_330);
nand U928 (N_928,In_2444,In_1321);
nor U929 (N_929,In_282,In_283);
nand U930 (N_930,In_782,In_953);
xor U931 (N_931,In_1810,In_2429);
nor U932 (N_932,In_1347,In_1716);
nand U933 (N_933,In_1162,In_1896);
nand U934 (N_934,In_2349,In_346);
nand U935 (N_935,In_926,In_2364);
and U936 (N_936,In_80,In_961);
or U937 (N_937,In_702,In_157);
nand U938 (N_938,In_1662,In_1535);
or U939 (N_939,In_986,In_487);
and U940 (N_940,In_2260,In_1128);
and U941 (N_941,In_1319,In_1372);
or U942 (N_942,In_1356,In_864);
nor U943 (N_943,In_766,In_2214);
nor U944 (N_944,In_1238,In_1691);
nand U945 (N_945,In_1445,In_2238);
nor U946 (N_946,In_474,In_74);
nor U947 (N_947,In_1137,In_1568);
nor U948 (N_948,In_2015,In_1168);
or U949 (N_949,In_481,In_224);
nand U950 (N_950,In_2032,In_321);
xor U951 (N_951,In_2226,In_2354);
nand U952 (N_952,In_906,In_1657);
nor U953 (N_953,In_114,In_737);
nand U954 (N_954,In_2338,In_600);
and U955 (N_955,In_2426,In_289);
nor U956 (N_956,In_471,In_2263);
nor U957 (N_957,In_2154,In_1684);
and U958 (N_958,In_515,In_2146);
and U959 (N_959,In_1835,In_489);
nor U960 (N_960,In_1690,In_1500);
or U961 (N_961,In_524,In_315);
nand U962 (N_962,In_139,In_660);
nor U963 (N_963,In_743,In_1526);
xor U964 (N_964,In_380,In_1994);
nand U965 (N_965,In_708,In_1172);
or U966 (N_966,In_705,In_426);
or U967 (N_967,In_2294,In_225);
and U968 (N_968,In_1584,In_281);
and U969 (N_969,In_353,In_2342);
xor U970 (N_970,In_1036,In_396);
and U971 (N_971,In_453,In_1085);
nand U972 (N_972,In_381,In_533);
nand U973 (N_973,In_1045,In_1646);
xnor U974 (N_974,In_669,In_1010);
nand U975 (N_975,In_1218,In_2104);
or U976 (N_976,In_1634,In_1602);
nand U977 (N_977,In_136,In_677);
and U978 (N_978,In_2387,In_1756);
xor U979 (N_979,In_2483,In_1129);
nand U980 (N_980,In_1749,In_604);
nor U981 (N_981,In_728,In_23);
or U982 (N_982,In_919,In_2086);
or U983 (N_983,In_911,In_437);
or U984 (N_984,In_1928,In_999);
xor U985 (N_985,In_787,In_977);
and U986 (N_986,In_2388,In_1071);
nor U987 (N_987,In_118,In_75);
xor U988 (N_988,In_2194,In_144);
nor U989 (N_989,In_1894,In_1533);
nand U990 (N_990,In_2196,In_2040);
or U991 (N_991,In_449,In_2152);
nor U992 (N_992,In_865,In_618);
and U993 (N_993,In_305,In_727);
or U994 (N_994,In_1987,In_1298);
nor U995 (N_995,In_530,In_395);
and U996 (N_996,In_653,In_828);
xnor U997 (N_997,In_733,In_410);
nor U998 (N_998,In_867,In_1082);
xnor U999 (N_999,In_1437,In_1693);
and U1000 (N_1000,In_856,In_458);
xor U1001 (N_1001,In_1161,In_2442);
or U1002 (N_1002,In_956,In_2417);
and U1003 (N_1003,In_2337,In_970);
xnor U1004 (N_1004,In_1468,In_170);
nand U1005 (N_1005,In_1812,In_1466);
nor U1006 (N_1006,In_1141,In_1753);
nor U1007 (N_1007,In_1563,In_1057);
nor U1008 (N_1008,In_523,In_2093);
nand U1009 (N_1009,In_1190,In_668);
nand U1010 (N_1010,In_1311,In_1822);
nor U1011 (N_1011,In_1912,In_1618);
and U1012 (N_1012,In_1899,In_276);
nor U1013 (N_1013,In_2325,In_511);
and U1014 (N_1014,In_1279,In_2209);
and U1015 (N_1015,In_2027,In_1365);
or U1016 (N_1016,In_1068,In_2411);
nand U1017 (N_1017,In_2289,In_336);
nand U1018 (N_1018,In_1735,In_86);
nor U1019 (N_1019,In_1135,In_2009);
or U1020 (N_1020,In_1895,In_312);
nand U1021 (N_1021,In_796,In_2204);
nor U1022 (N_1022,In_1293,In_2058);
and U1023 (N_1023,In_876,In_247);
nand U1024 (N_1024,In_2207,In_950);
nand U1025 (N_1025,In_2174,In_1869);
xnor U1026 (N_1026,In_1996,In_1388);
and U1027 (N_1027,In_2478,In_2033);
or U1028 (N_1028,In_1834,In_2212);
nand U1029 (N_1029,In_2465,In_1084);
nand U1030 (N_1030,In_2116,In_1393);
or U1031 (N_1031,In_1908,In_2039);
or U1032 (N_1032,In_311,In_612);
xor U1033 (N_1033,In_444,In_1480);
xor U1034 (N_1034,In_1148,In_973);
nand U1035 (N_1035,In_1929,In_2284);
nor U1036 (N_1036,In_2110,In_1844);
nand U1037 (N_1037,In_108,In_1947);
or U1038 (N_1038,In_403,In_109);
nand U1039 (N_1039,In_724,In_2022);
or U1040 (N_1040,In_1825,In_1793);
xor U1041 (N_1041,In_971,In_1185);
or U1042 (N_1042,In_1595,In_2312);
xor U1043 (N_1043,In_1826,In_572);
xor U1044 (N_1044,In_425,In_591);
nor U1045 (N_1045,In_639,In_675);
nor U1046 (N_1046,In_1278,In_1710);
nand U1047 (N_1047,In_273,In_2075);
and U1048 (N_1048,In_1659,In_2155);
xor U1049 (N_1049,In_783,In_1649);
and U1050 (N_1050,In_216,In_621);
xnor U1051 (N_1051,In_615,In_1435);
xor U1052 (N_1052,In_2431,In_1814);
nor U1053 (N_1053,In_803,In_730);
and U1054 (N_1054,In_1173,In_1578);
xnor U1055 (N_1055,In_834,In_1358);
and U1056 (N_1056,In_2421,In_1728);
nor U1057 (N_1057,In_924,In_1184);
xor U1058 (N_1058,In_1823,In_1538);
and U1059 (N_1059,In_2076,In_1654);
nor U1060 (N_1060,In_928,In_2185);
xnor U1061 (N_1061,In_1829,In_1751);
and U1062 (N_1062,In_1192,In_1157);
and U1063 (N_1063,In_1041,In_370);
or U1064 (N_1064,In_477,In_780);
xnor U1065 (N_1065,In_2255,In_252);
nand U1066 (N_1066,In_1296,In_303);
or U1067 (N_1067,In_1330,In_124);
nand U1068 (N_1068,In_168,In_1537);
nor U1069 (N_1069,In_1407,In_2348);
nand U1070 (N_1070,In_2012,In_1516);
nor U1071 (N_1071,In_121,In_1878);
xor U1072 (N_1072,In_776,In_1524);
nand U1073 (N_1073,In_1760,In_1534);
xnor U1074 (N_1074,In_1029,In_842);
xor U1075 (N_1075,In_493,In_590);
nand U1076 (N_1076,In_1163,In_752);
nor U1077 (N_1077,In_1843,In_1302);
and U1078 (N_1078,In_450,In_1778);
nor U1079 (N_1079,In_1191,In_1882);
nand U1080 (N_1080,In_1050,In_1732);
xor U1081 (N_1081,In_2392,In_1918);
and U1082 (N_1082,In_582,In_976);
xor U1083 (N_1083,In_326,In_779);
or U1084 (N_1084,In_376,In_1286);
and U1085 (N_1085,In_534,In_1506);
and U1086 (N_1086,In_2005,In_1324);
and U1087 (N_1087,In_1815,In_46);
or U1088 (N_1088,In_2215,In_1542);
nand U1089 (N_1089,In_2336,In_2482);
xor U1090 (N_1090,In_1448,In_2424);
xor U1091 (N_1091,In_532,In_921);
xor U1092 (N_1092,In_1489,In_1067);
and U1093 (N_1093,In_2235,In_1117);
nand U1094 (N_1094,In_2466,In_1316);
nand U1095 (N_1095,In_1884,In_2382);
or U1096 (N_1096,In_2031,In_1270);
or U1097 (N_1097,In_2175,In_742);
or U1098 (N_1098,In_959,In_233);
xnor U1099 (N_1099,In_1551,In_667);
nand U1100 (N_1100,In_1758,In_9);
and U1101 (N_1101,In_1004,In_889);
nand U1102 (N_1102,In_1411,In_758);
nand U1103 (N_1103,In_2456,In_1498);
or U1104 (N_1104,In_763,In_1788);
xnor U1105 (N_1105,In_198,In_1443);
nor U1106 (N_1106,In_94,In_423);
or U1107 (N_1107,In_2081,In_292);
xor U1108 (N_1108,In_503,In_2459);
and U1109 (N_1109,In_455,In_2156);
or U1110 (N_1110,In_309,In_95);
nor U1111 (N_1111,In_1323,In_809);
nand U1112 (N_1112,In_564,In_1248);
nor U1113 (N_1113,In_2322,In_366);
nand U1114 (N_1114,In_1123,In_202);
or U1115 (N_1115,In_2169,In_718);
nand U1116 (N_1116,In_2498,In_1338);
nor U1117 (N_1117,In_644,In_2335);
nand U1118 (N_1118,In_54,In_2470);
or U1119 (N_1119,In_1806,In_659);
xnor U1120 (N_1120,In_2150,In_30);
nor U1121 (N_1121,In_1772,In_1415);
nor U1122 (N_1122,In_1262,In_1641);
xor U1123 (N_1123,In_2313,In_1581);
and U1124 (N_1124,In_545,In_2030);
nand U1125 (N_1125,In_56,In_120);
xor U1126 (N_1126,In_70,In_2400);
nor U1127 (N_1127,In_1107,In_331);
xnor U1128 (N_1128,In_1034,In_375);
or U1129 (N_1129,In_1754,In_325);
or U1130 (N_1130,In_1531,In_1877);
and U1131 (N_1131,In_2484,In_284);
nand U1132 (N_1132,In_2256,In_1014);
xor U1133 (N_1133,In_938,In_185);
nand U1134 (N_1134,In_800,In_608);
or U1135 (N_1135,In_2118,In_1482);
and U1136 (N_1136,In_2222,In_1898);
or U1137 (N_1137,In_159,In_2422);
nor U1138 (N_1138,In_617,In_2438);
xor U1139 (N_1139,In_2373,In_1096);
xnor U1140 (N_1140,In_655,In_1380);
nand U1141 (N_1141,In_1039,In_365);
nor U1142 (N_1142,In_2391,In_1604);
nand U1143 (N_1143,In_1150,In_184);
nor U1144 (N_1144,In_1682,In_697);
nand U1145 (N_1145,In_194,In_902);
nand U1146 (N_1146,In_153,In_1580);
nand U1147 (N_1147,In_651,In_1376);
xor U1148 (N_1148,In_2053,In_817);
nand U1149 (N_1149,In_359,In_1024);
and U1150 (N_1150,In_2418,In_408);
nor U1151 (N_1151,In_1009,In_150);
nand U1152 (N_1152,In_1171,In_195);
xor U1153 (N_1153,In_721,In_434);
or U1154 (N_1154,In_731,In_1958);
nand U1155 (N_1155,In_2171,In_2274);
xor U1156 (N_1156,In_478,In_60);
nand U1157 (N_1157,In_674,In_1570);
nand U1158 (N_1158,In_2432,In_1501);
and U1159 (N_1159,In_789,In_1502);
nor U1160 (N_1160,In_1543,In_357);
xor U1161 (N_1161,In_980,In_1081);
and U1162 (N_1162,In_848,In_717);
nand U1163 (N_1163,In_965,In_923);
xnor U1164 (N_1164,In_1901,In_2234);
nor U1165 (N_1165,In_829,In_143);
and U1166 (N_1166,In_164,In_2439);
nand U1167 (N_1167,In_1680,In_173);
xor U1168 (N_1168,In_1417,In_2462);
xnor U1169 (N_1169,In_99,In_930);
or U1170 (N_1170,In_820,In_1104);
nor U1171 (N_1171,In_369,In_711);
nor U1172 (N_1172,In_1964,In_739);
or U1173 (N_1173,In_1109,In_1974);
or U1174 (N_1174,In_2102,In_1871);
and U1175 (N_1175,In_32,In_2280);
nand U1176 (N_1176,In_1268,In_1704);
or U1177 (N_1177,In_1187,In_1374);
nor U1178 (N_1178,In_169,In_2080);
nor U1179 (N_1179,In_1152,In_1147);
and U1180 (N_1180,In_1719,In_127);
nand U1181 (N_1181,In_929,In_2437);
or U1182 (N_1182,In_2038,In_1902);
nand U1183 (N_1183,In_2003,In_962);
nor U1184 (N_1184,In_665,In_334);
xor U1185 (N_1185,In_1090,In_716);
or U1186 (N_1186,In_2488,In_319);
and U1187 (N_1187,In_1712,In_1967);
and U1188 (N_1188,In_1804,In_1842);
xor U1189 (N_1189,In_179,In_1585);
and U1190 (N_1190,In_1294,In_2339);
nand U1191 (N_1191,In_1917,In_993);
xor U1192 (N_1192,In_1430,In_469);
or U1193 (N_1193,In_808,In_1384);
and U1194 (N_1194,In_47,In_2091);
nor U1195 (N_1195,In_1226,In_955);
and U1196 (N_1196,In_270,In_2307);
nor U1197 (N_1197,In_1853,In_300);
nor U1198 (N_1198,In_210,In_3);
nor U1199 (N_1199,In_874,In_1138);
and U1200 (N_1200,In_138,In_2323);
xor U1201 (N_1201,In_694,In_490);
nand U1202 (N_1202,In_1198,In_700);
and U1203 (N_1203,In_199,In_1777);
nand U1204 (N_1204,In_83,In_409);
or U1205 (N_1205,In_278,In_1459);
nor U1206 (N_1206,In_1541,In_2413);
and U1207 (N_1207,In_884,In_1521);
xor U1208 (N_1208,In_2251,In_1599);
nand U1209 (N_1209,In_1775,In_1856);
or U1210 (N_1210,In_1473,In_821);
and U1211 (N_1211,In_905,In_2045);
or U1212 (N_1212,In_1114,In_378);
nand U1213 (N_1213,In_2447,In_1496);
and U1214 (N_1214,In_1862,In_1310);
nor U1215 (N_1215,In_2136,In_459);
or U1216 (N_1216,In_417,In_1694);
nand U1217 (N_1217,In_2237,In_451);
xnor U1218 (N_1218,In_1972,In_421);
nor U1219 (N_1219,In_1588,In_1739);
nor U1220 (N_1220,In_2179,In_563);
nand U1221 (N_1221,In_652,In_1927);
nand U1222 (N_1222,In_2242,In_968);
or U1223 (N_1223,In_1227,In_1250);
nand U1224 (N_1224,In_2121,In_2131);
and U1225 (N_1225,In_267,In_2401);
xnor U1226 (N_1226,In_2340,In_1005);
or U1227 (N_1227,In_268,In_689);
and U1228 (N_1228,In_1951,In_2181);
xor U1229 (N_1229,In_220,In_1276);
and U1230 (N_1230,In_389,In_349);
or U1231 (N_1231,In_2463,In_661);
or U1232 (N_1232,In_1573,In_2360);
nand U1233 (N_1233,In_1274,In_2362);
nand U1234 (N_1234,In_823,In_894);
or U1235 (N_1235,In_443,In_1426);
or U1236 (N_1236,In_2328,In_755);
nor U1237 (N_1237,In_510,In_1470);
nand U1238 (N_1238,In_1556,In_1956);
nor U1239 (N_1239,In_666,In_2224);
nand U1240 (N_1240,In_230,In_1006);
and U1241 (N_1241,In_431,In_1318);
nor U1242 (N_1242,In_2219,In_2211);
nand U1243 (N_1243,In_1670,In_695);
nor U1244 (N_1244,In_229,In_430);
and U1245 (N_1245,In_1051,In_1875);
nand U1246 (N_1246,In_753,In_1087);
nand U1247 (N_1247,In_1755,In_1865);
and U1248 (N_1248,In_983,In_322);
or U1249 (N_1249,In_1207,In_912);
nor U1250 (N_1250,In_1412,In_684);
or U1251 (N_1251,In_1113,In_2375);
nor U1252 (N_1252,In_611,In_518);
nor U1253 (N_1253,In_1657,In_1669);
xnor U1254 (N_1254,In_1652,In_351);
or U1255 (N_1255,In_1121,In_1224);
nor U1256 (N_1256,In_8,In_1572);
xor U1257 (N_1257,In_290,In_415);
or U1258 (N_1258,In_2034,In_1737);
nor U1259 (N_1259,In_200,In_876);
and U1260 (N_1260,In_754,In_335);
xor U1261 (N_1261,In_619,In_1636);
or U1262 (N_1262,In_1273,In_297);
xor U1263 (N_1263,In_637,In_510);
nor U1264 (N_1264,In_2210,In_2036);
xor U1265 (N_1265,In_2195,In_947);
nand U1266 (N_1266,In_923,In_2255);
nand U1267 (N_1267,In_826,In_2338);
nand U1268 (N_1268,In_1383,In_1467);
and U1269 (N_1269,In_1158,In_2316);
nand U1270 (N_1270,In_2050,In_1530);
and U1271 (N_1271,In_1224,In_1798);
xor U1272 (N_1272,In_890,In_1424);
nor U1273 (N_1273,In_2486,In_266);
and U1274 (N_1274,In_2284,In_911);
nor U1275 (N_1275,In_1934,In_1765);
nor U1276 (N_1276,In_921,In_1401);
or U1277 (N_1277,In_1433,In_1185);
xnor U1278 (N_1278,In_934,In_1612);
xor U1279 (N_1279,In_880,In_1054);
xor U1280 (N_1280,In_190,In_1672);
xor U1281 (N_1281,In_1138,In_1071);
nor U1282 (N_1282,In_133,In_696);
nand U1283 (N_1283,In_1301,In_465);
nor U1284 (N_1284,In_1735,In_160);
and U1285 (N_1285,In_560,In_360);
xor U1286 (N_1286,In_1519,In_497);
and U1287 (N_1287,In_660,In_584);
or U1288 (N_1288,In_1312,In_836);
nand U1289 (N_1289,In_1893,In_1072);
xor U1290 (N_1290,In_560,In_1829);
xnor U1291 (N_1291,In_1618,In_1554);
nand U1292 (N_1292,In_557,In_2143);
or U1293 (N_1293,In_1420,In_1383);
nor U1294 (N_1294,In_589,In_25);
or U1295 (N_1295,In_1252,In_236);
nand U1296 (N_1296,In_2259,In_2322);
nand U1297 (N_1297,In_534,In_872);
xnor U1298 (N_1298,In_512,In_646);
or U1299 (N_1299,In_1577,In_1233);
or U1300 (N_1300,In_1180,In_1341);
or U1301 (N_1301,In_1800,In_1841);
xnor U1302 (N_1302,In_2479,In_713);
nor U1303 (N_1303,In_1278,In_913);
nand U1304 (N_1304,In_1597,In_543);
nand U1305 (N_1305,In_2017,In_1863);
nand U1306 (N_1306,In_1598,In_57);
and U1307 (N_1307,In_2119,In_979);
nand U1308 (N_1308,In_414,In_1617);
or U1309 (N_1309,In_181,In_162);
xnor U1310 (N_1310,In_2377,In_768);
nand U1311 (N_1311,In_915,In_1351);
and U1312 (N_1312,In_131,In_386);
nor U1313 (N_1313,In_2067,In_1279);
xnor U1314 (N_1314,In_1715,In_690);
or U1315 (N_1315,In_2261,In_289);
xor U1316 (N_1316,In_1682,In_1923);
xnor U1317 (N_1317,In_410,In_1009);
nor U1318 (N_1318,In_390,In_1715);
xnor U1319 (N_1319,In_1583,In_1937);
or U1320 (N_1320,In_1569,In_2292);
or U1321 (N_1321,In_1449,In_1396);
or U1322 (N_1322,In_2061,In_1241);
and U1323 (N_1323,In_1945,In_282);
nor U1324 (N_1324,In_1037,In_782);
nand U1325 (N_1325,In_2117,In_1350);
nor U1326 (N_1326,In_409,In_2012);
or U1327 (N_1327,In_850,In_1755);
or U1328 (N_1328,In_2095,In_314);
and U1329 (N_1329,In_2298,In_620);
or U1330 (N_1330,In_2403,In_1996);
nor U1331 (N_1331,In_1329,In_163);
xor U1332 (N_1332,In_1930,In_1908);
nor U1333 (N_1333,In_566,In_2038);
nand U1334 (N_1334,In_142,In_1291);
or U1335 (N_1335,In_1120,In_8);
and U1336 (N_1336,In_959,In_400);
or U1337 (N_1337,In_1467,In_1785);
nand U1338 (N_1338,In_1123,In_921);
or U1339 (N_1339,In_308,In_1974);
nand U1340 (N_1340,In_1104,In_1114);
and U1341 (N_1341,In_781,In_799);
nand U1342 (N_1342,In_2023,In_587);
nand U1343 (N_1343,In_2292,In_1282);
or U1344 (N_1344,In_2094,In_2271);
xor U1345 (N_1345,In_108,In_1220);
and U1346 (N_1346,In_111,In_2123);
and U1347 (N_1347,In_2395,In_1264);
or U1348 (N_1348,In_1015,In_988);
nand U1349 (N_1349,In_1083,In_433);
nand U1350 (N_1350,In_2101,In_2411);
or U1351 (N_1351,In_2174,In_2044);
xnor U1352 (N_1352,In_416,In_1258);
or U1353 (N_1353,In_1488,In_432);
nand U1354 (N_1354,In_1262,In_755);
xor U1355 (N_1355,In_2390,In_2090);
nor U1356 (N_1356,In_1302,In_1977);
nand U1357 (N_1357,In_704,In_1412);
xnor U1358 (N_1358,In_569,In_178);
nor U1359 (N_1359,In_1481,In_901);
nand U1360 (N_1360,In_1358,In_391);
or U1361 (N_1361,In_1178,In_1373);
or U1362 (N_1362,In_505,In_2114);
xor U1363 (N_1363,In_1476,In_997);
and U1364 (N_1364,In_1364,In_2003);
and U1365 (N_1365,In_2090,In_2071);
and U1366 (N_1366,In_879,In_851);
xnor U1367 (N_1367,In_2382,In_17);
xnor U1368 (N_1368,In_1438,In_1145);
nand U1369 (N_1369,In_1176,In_813);
nor U1370 (N_1370,In_424,In_965);
nor U1371 (N_1371,In_973,In_1835);
nand U1372 (N_1372,In_2071,In_2067);
nand U1373 (N_1373,In_1068,In_1303);
xnor U1374 (N_1374,In_632,In_33);
or U1375 (N_1375,In_768,In_1606);
or U1376 (N_1376,In_2125,In_669);
or U1377 (N_1377,In_904,In_687);
xor U1378 (N_1378,In_617,In_1191);
or U1379 (N_1379,In_2453,In_368);
xnor U1380 (N_1380,In_1232,In_2251);
nor U1381 (N_1381,In_1118,In_1944);
xnor U1382 (N_1382,In_1018,In_262);
xor U1383 (N_1383,In_675,In_2148);
nor U1384 (N_1384,In_1681,In_1075);
xnor U1385 (N_1385,In_117,In_1985);
or U1386 (N_1386,In_1690,In_1945);
xor U1387 (N_1387,In_35,In_1459);
nor U1388 (N_1388,In_2012,In_1424);
xnor U1389 (N_1389,In_889,In_2389);
or U1390 (N_1390,In_1731,In_554);
xor U1391 (N_1391,In_153,In_881);
nand U1392 (N_1392,In_1755,In_2492);
nand U1393 (N_1393,In_2110,In_247);
and U1394 (N_1394,In_11,In_1536);
nor U1395 (N_1395,In_2038,In_1538);
nand U1396 (N_1396,In_421,In_398);
or U1397 (N_1397,In_1830,In_1174);
and U1398 (N_1398,In_402,In_1202);
and U1399 (N_1399,In_1352,In_2223);
xnor U1400 (N_1400,In_1255,In_1518);
xnor U1401 (N_1401,In_309,In_960);
or U1402 (N_1402,In_2279,In_2024);
nor U1403 (N_1403,In_1807,In_7);
nand U1404 (N_1404,In_763,In_1855);
xor U1405 (N_1405,In_862,In_2360);
nor U1406 (N_1406,In_1712,In_950);
and U1407 (N_1407,In_1006,In_1578);
nor U1408 (N_1408,In_1389,In_2117);
and U1409 (N_1409,In_2351,In_2283);
nand U1410 (N_1410,In_1402,In_50);
nand U1411 (N_1411,In_1005,In_1695);
nor U1412 (N_1412,In_2339,In_26);
nand U1413 (N_1413,In_2456,In_895);
nor U1414 (N_1414,In_1360,In_1216);
and U1415 (N_1415,In_802,In_1052);
nor U1416 (N_1416,In_137,In_370);
or U1417 (N_1417,In_949,In_842);
nand U1418 (N_1418,In_1486,In_2277);
xor U1419 (N_1419,In_1283,In_1508);
xnor U1420 (N_1420,In_295,In_2384);
nand U1421 (N_1421,In_2011,In_1354);
nand U1422 (N_1422,In_967,In_601);
and U1423 (N_1423,In_1677,In_197);
nand U1424 (N_1424,In_1462,In_802);
nand U1425 (N_1425,In_364,In_2013);
xnor U1426 (N_1426,In_601,In_2088);
or U1427 (N_1427,In_829,In_1451);
nand U1428 (N_1428,In_645,In_1346);
and U1429 (N_1429,In_528,In_484);
nor U1430 (N_1430,In_2153,In_433);
or U1431 (N_1431,In_1587,In_2295);
nor U1432 (N_1432,In_965,In_1641);
and U1433 (N_1433,In_1526,In_89);
nor U1434 (N_1434,In_199,In_754);
or U1435 (N_1435,In_2210,In_1425);
nand U1436 (N_1436,In_2209,In_940);
nor U1437 (N_1437,In_683,In_847);
or U1438 (N_1438,In_2210,In_2489);
nand U1439 (N_1439,In_269,In_109);
or U1440 (N_1440,In_2491,In_813);
nor U1441 (N_1441,In_2043,In_1545);
or U1442 (N_1442,In_348,In_1328);
nor U1443 (N_1443,In_891,In_1915);
nor U1444 (N_1444,In_1249,In_2405);
nor U1445 (N_1445,In_1625,In_1384);
xor U1446 (N_1446,In_164,In_1054);
nor U1447 (N_1447,In_1342,In_1790);
and U1448 (N_1448,In_212,In_2150);
nor U1449 (N_1449,In_1989,In_456);
nor U1450 (N_1450,In_741,In_32);
or U1451 (N_1451,In_1464,In_650);
and U1452 (N_1452,In_2419,In_720);
nor U1453 (N_1453,In_2308,In_2075);
nand U1454 (N_1454,In_1231,In_1750);
or U1455 (N_1455,In_2491,In_699);
nor U1456 (N_1456,In_2161,In_2181);
or U1457 (N_1457,In_1286,In_1919);
xor U1458 (N_1458,In_610,In_2279);
xor U1459 (N_1459,In_2332,In_62);
and U1460 (N_1460,In_2424,In_544);
xnor U1461 (N_1461,In_342,In_2117);
xor U1462 (N_1462,In_1968,In_2437);
nor U1463 (N_1463,In_1848,In_619);
and U1464 (N_1464,In_383,In_78);
nor U1465 (N_1465,In_109,In_1651);
or U1466 (N_1466,In_1204,In_1836);
or U1467 (N_1467,In_2434,In_2035);
and U1468 (N_1468,In_2420,In_1568);
nor U1469 (N_1469,In_1318,In_2154);
and U1470 (N_1470,In_2280,In_1405);
xor U1471 (N_1471,In_1736,In_544);
nand U1472 (N_1472,In_1669,In_166);
and U1473 (N_1473,In_2413,In_967);
nand U1474 (N_1474,In_399,In_395);
nand U1475 (N_1475,In_917,In_628);
or U1476 (N_1476,In_220,In_1184);
nand U1477 (N_1477,In_1448,In_839);
and U1478 (N_1478,In_229,In_1027);
xor U1479 (N_1479,In_1149,In_2401);
nor U1480 (N_1480,In_2243,In_469);
and U1481 (N_1481,In_1902,In_1079);
and U1482 (N_1482,In_478,In_388);
and U1483 (N_1483,In_1790,In_2201);
or U1484 (N_1484,In_1248,In_927);
or U1485 (N_1485,In_359,In_1107);
and U1486 (N_1486,In_1768,In_1059);
and U1487 (N_1487,In_524,In_850);
nand U1488 (N_1488,In_1881,In_2434);
and U1489 (N_1489,In_1504,In_2412);
and U1490 (N_1490,In_2025,In_2273);
nor U1491 (N_1491,In_240,In_2441);
nand U1492 (N_1492,In_1925,In_1270);
nor U1493 (N_1493,In_1287,In_271);
nor U1494 (N_1494,In_1673,In_1335);
nand U1495 (N_1495,In_623,In_948);
nand U1496 (N_1496,In_2036,In_920);
xnor U1497 (N_1497,In_658,In_1919);
nand U1498 (N_1498,In_377,In_2099);
or U1499 (N_1499,In_863,In_1642);
and U1500 (N_1500,In_1250,In_1693);
or U1501 (N_1501,In_115,In_1063);
and U1502 (N_1502,In_2281,In_1117);
or U1503 (N_1503,In_231,In_1980);
or U1504 (N_1504,In_856,In_1839);
xor U1505 (N_1505,In_433,In_1102);
or U1506 (N_1506,In_315,In_1704);
nor U1507 (N_1507,In_1562,In_1978);
or U1508 (N_1508,In_1803,In_1087);
xor U1509 (N_1509,In_1046,In_1142);
nand U1510 (N_1510,In_463,In_2011);
or U1511 (N_1511,In_1074,In_237);
or U1512 (N_1512,In_1931,In_203);
or U1513 (N_1513,In_2317,In_833);
xor U1514 (N_1514,In_384,In_1558);
nor U1515 (N_1515,In_1038,In_185);
nor U1516 (N_1516,In_1319,In_2376);
xnor U1517 (N_1517,In_2431,In_2089);
nor U1518 (N_1518,In_1197,In_2315);
or U1519 (N_1519,In_1279,In_214);
or U1520 (N_1520,In_1205,In_1367);
or U1521 (N_1521,In_2139,In_1538);
nor U1522 (N_1522,In_437,In_2496);
nor U1523 (N_1523,In_1529,In_1095);
xor U1524 (N_1524,In_1218,In_103);
or U1525 (N_1525,In_17,In_1553);
xor U1526 (N_1526,In_1912,In_413);
nand U1527 (N_1527,In_134,In_2103);
xor U1528 (N_1528,In_791,In_1188);
and U1529 (N_1529,In_893,In_900);
xor U1530 (N_1530,In_492,In_60);
nor U1531 (N_1531,In_1482,In_842);
or U1532 (N_1532,In_1339,In_102);
nor U1533 (N_1533,In_1308,In_1991);
nor U1534 (N_1534,In_2460,In_1641);
nand U1535 (N_1535,In_1184,In_693);
xnor U1536 (N_1536,In_1138,In_1541);
or U1537 (N_1537,In_805,In_928);
and U1538 (N_1538,In_2290,In_160);
and U1539 (N_1539,In_1302,In_2451);
xnor U1540 (N_1540,In_829,In_2197);
nand U1541 (N_1541,In_1407,In_1941);
nand U1542 (N_1542,In_589,In_908);
xor U1543 (N_1543,In_53,In_1094);
xor U1544 (N_1544,In_188,In_1855);
or U1545 (N_1545,In_1251,In_320);
xor U1546 (N_1546,In_1429,In_1832);
xor U1547 (N_1547,In_1496,In_1124);
nor U1548 (N_1548,In_2022,In_1827);
nor U1549 (N_1549,In_694,In_2318);
and U1550 (N_1550,In_1537,In_2415);
xor U1551 (N_1551,In_2016,In_893);
and U1552 (N_1552,In_167,In_1730);
nor U1553 (N_1553,In_2304,In_15);
nand U1554 (N_1554,In_2383,In_2409);
and U1555 (N_1555,In_764,In_2281);
xnor U1556 (N_1556,In_2010,In_1216);
nor U1557 (N_1557,In_2349,In_2195);
nand U1558 (N_1558,In_1357,In_875);
or U1559 (N_1559,In_1968,In_380);
xor U1560 (N_1560,In_486,In_2378);
or U1561 (N_1561,In_1934,In_535);
nor U1562 (N_1562,In_1021,In_1528);
nand U1563 (N_1563,In_113,In_363);
nand U1564 (N_1564,In_2242,In_653);
and U1565 (N_1565,In_402,In_2186);
nand U1566 (N_1566,In_2445,In_1158);
nor U1567 (N_1567,In_739,In_2439);
or U1568 (N_1568,In_440,In_1196);
nand U1569 (N_1569,In_1388,In_958);
xor U1570 (N_1570,In_551,In_2433);
and U1571 (N_1571,In_2202,In_984);
xor U1572 (N_1572,In_1209,In_2106);
xor U1573 (N_1573,In_288,In_878);
nor U1574 (N_1574,In_32,In_387);
nand U1575 (N_1575,In_1671,In_592);
and U1576 (N_1576,In_208,In_591);
or U1577 (N_1577,In_347,In_2028);
xor U1578 (N_1578,In_1584,In_1061);
and U1579 (N_1579,In_424,In_813);
and U1580 (N_1580,In_1258,In_2224);
xor U1581 (N_1581,In_1782,In_1955);
xor U1582 (N_1582,In_1743,In_1273);
nor U1583 (N_1583,In_410,In_1799);
and U1584 (N_1584,In_2158,In_1815);
nor U1585 (N_1585,In_646,In_35);
xor U1586 (N_1586,In_1717,In_117);
xnor U1587 (N_1587,In_570,In_697);
or U1588 (N_1588,In_1309,In_339);
and U1589 (N_1589,In_665,In_1729);
and U1590 (N_1590,In_1253,In_670);
xor U1591 (N_1591,In_1456,In_418);
or U1592 (N_1592,In_46,In_2360);
and U1593 (N_1593,In_2403,In_1201);
or U1594 (N_1594,In_1678,In_988);
xor U1595 (N_1595,In_2126,In_248);
and U1596 (N_1596,In_213,In_34);
xnor U1597 (N_1597,In_1814,In_1880);
and U1598 (N_1598,In_529,In_875);
and U1599 (N_1599,In_1937,In_1091);
nand U1600 (N_1600,In_1292,In_1399);
nand U1601 (N_1601,In_18,In_929);
xnor U1602 (N_1602,In_1089,In_1463);
nor U1603 (N_1603,In_2099,In_963);
xnor U1604 (N_1604,In_1622,In_1705);
nor U1605 (N_1605,In_31,In_1998);
nor U1606 (N_1606,In_157,In_47);
nor U1607 (N_1607,In_740,In_19);
nand U1608 (N_1608,In_1175,In_817);
nand U1609 (N_1609,In_403,In_1577);
nand U1610 (N_1610,In_1687,In_1077);
and U1611 (N_1611,In_1461,In_1126);
or U1612 (N_1612,In_1393,In_170);
or U1613 (N_1613,In_209,In_1475);
xor U1614 (N_1614,In_886,In_2122);
and U1615 (N_1615,In_1055,In_377);
nor U1616 (N_1616,In_616,In_1299);
and U1617 (N_1617,In_1899,In_1227);
nand U1618 (N_1618,In_1689,In_1924);
nand U1619 (N_1619,In_955,In_1325);
or U1620 (N_1620,In_1784,In_1399);
nand U1621 (N_1621,In_1828,In_1545);
and U1622 (N_1622,In_836,In_1267);
xnor U1623 (N_1623,In_2434,In_343);
and U1624 (N_1624,In_1205,In_2200);
or U1625 (N_1625,In_1705,In_1945);
or U1626 (N_1626,In_33,In_1792);
or U1627 (N_1627,In_1230,In_1881);
nand U1628 (N_1628,In_424,In_921);
and U1629 (N_1629,In_722,In_2055);
or U1630 (N_1630,In_337,In_689);
xor U1631 (N_1631,In_1578,In_1082);
nand U1632 (N_1632,In_862,In_2302);
and U1633 (N_1633,In_2084,In_2295);
nand U1634 (N_1634,In_1687,In_326);
and U1635 (N_1635,In_2454,In_1974);
xnor U1636 (N_1636,In_684,In_665);
nand U1637 (N_1637,In_246,In_1437);
nand U1638 (N_1638,In_2068,In_548);
or U1639 (N_1639,In_2272,In_446);
nand U1640 (N_1640,In_963,In_946);
and U1641 (N_1641,In_1729,In_1829);
and U1642 (N_1642,In_1206,In_1120);
nor U1643 (N_1643,In_372,In_2282);
nand U1644 (N_1644,In_1107,In_111);
and U1645 (N_1645,In_2454,In_942);
and U1646 (N_1646,In_195,In_1855);
nand U1647 (N_1647,In_1567,In_2472);
or U1648 (N_1648,In_1793,In_281);
or U1649 (N_1649,In_956,In_1463);
nor U1650 (N_1650,In_1274,In_1468);
nand U1651 (N_1651,In_35,In_587);
nand U1652 (N_1652,In_1965,In_589);
nand U1653 (N_1653,In_1441,In_1207);
and U1654 (N_1654,In_368,In_413);
nor U1655 (N_1655,In_1931,In_211);
or U1656 (N_1656,In_1721,In_2244);
nand U1657 (N_1657,In_1164,In_1392);
nor U1658 (N_1658,In_399,In_1709);
nand U1659 (N_1659,In_1826,In_1495);
nand U1660 (N_1660,In_2227,In_2073);
xor U1661 (N_1661,In_1548,In_1688);
or U1662 (N_1662,In_1304,In_535);
or U1663 (N_1663,In_2430,In_1);
or U1664 (N_1664,In_2297,In_1697);
and U1665 (N_1665,In_813,In_1799);
nor U1666 (N_1666,In_1305,In_2193);
or U1667 (N_1667,In_1945,In_2078);
nor U1668 (N_1668,In_1777,In_2276);
or U1669 (N_1669,In_2194,In_1156);
nor U1670 (N_1670,In_461,In_1787);
and U1671 (N_1671,In_189,In_1787);
or U1672 (N_1672,In_683,In_1225);
xnor U1673 (N_1673,In_868,In_966);
and U1674 (N_1674,In_1255,In_1766);
and U1675 (N_1675,In_1828,In_2487);
nand U1676 (N_1676,In_2309,In_1597);
nand U1677 (N_1677,In_996,In_1105);
and U1678 (N_1678,In_1250,In_2198);
or U1679 (N_1679,In_1613,In_474);
or U1680 (N_1680,In_581,In_2206);
nor U1681 (N_1681,In_460,In_1365);
and U1682 (N_1682,In_1797,In_1564);
nand U1683 (N_1683,In_500,In_156);
xor U1684 (N_1684,In_1314,In_1159);
nor U1685 (N_1685,In_2242,In_720);
nor U1686 (N_1686,In_430,In_1730);
xor U1687 (N_1687,In_1601,In_137);
xnor U1688 (N_1688,In_1066,In_2389);
nor U1689 (N_1689,In_843,In_456);
nand U1690 (N_1690,In_2071,In_897);
and U1691 (N_1691,In_1858,In_1126);
xnor U1692 (N_1692,In_2068,In_1492);
xor U1693 (N_1693,In_706,In_2236);
xor U1694 (N_1694,In_2212,In_2389);
or U1695 (N_1695,In_332,In_2241);
nand U1696 (N_1696,In_2002,In_2435);
nand U1697 (N_1697,In_1104,In_2002);
or U1698 (N_1698,In_722,In_343);
nor U1699 (N_1699,In_353,In_1716);
nor U1700 (N_1700,In_850,In_1522);
xor U1701 (N_1701,In_1290,In_669);
and U1702 (N_1702,In_1311,In_2177);
xor U1703 (N_1703,In_773,In_688);
nand U1704 (N_1704,In_1086,In_1801);
and U1705 (N_1705,In_2379,In_211);
xnor U1706 (N_1706,In_1957,In_2100);
and U1707 (N_1707,In_1610,In_235);
nand U1708 (N_1708,In_1180,In_248);
nor U1709 (N_1709,In_1701,In_1938);
and U1710 (N_1710,In_647,In_357);
nor U1711 (N_1711,In_1804,In_1117);
nand U1712 (N_1712,In_24,In_1929);
or U1713 (N_1713,In_1378,In_648);
nand U1714 (N_1714,In_2216,In_1938);
nand U1715 (N_1715,In_2350,In_1110);
or U1716 (N_1716,In_360,In_254);
nor U1717 (N_1717,In_1397,In_1526);
nor U1718 (N_1718,In_790,In_718);
nor U1719 (N_1719,In_1185,In_798);
or U1720 (N_1720,In_2034,In_640);
nand U1721 (N_1721,In_1645,In_208);
xnor U1722 (N_1722,In_1937,In_8);
or U1723 (N_1723,In_881,In_2397);
xor U1724 (N_1724,In_109,In_532);
or U1725 (N_1725,In_2457,In_2332);
nor U1726 (N_1726,In_1706,In_307);
or U1727 (N_1727,In_1751,In_686);
nor U1728 (N_1728,In_2121,In_190);
xnor U1729 (N_1729,In_581,In_2350);
nor U1730 (N_1730,In_681,In_2102);
xor U1731 (N_1731,In_972,In_1578);
nor U1732 (N_1732,In_1317,In_1010);
nand U1733 (N_1733,In_1827,In_2331);
and U1734 (N_1734,In_1664,In_907);
and U1735 (N_1735,In_732,In_1642);
nor U1736 (N_1736,In_359,In_2252);
nand U1737 (N_1737,In_305,In_1510);
or U1738 (N_1738,In_1662,In_657);
or U1739 (N_1739,In_2451,In_1158);
xor U1740 (N_1740,In_2430,In_616);
and U1741 (N_1741,In_631,In_521);
nor U1742 (N_1742,In_1992,In_2143);
nor U1743 (N_1743,In_1625,In_525);
nor U1744 (N_1744,In_1035,In_2077);
and U1745 (N_1745,In_2189,In_242);
nand U1746 (N_1746,In_171,In_100);
xor U1747 (N_1747,In_683,In_2423);
xor U1748 (N_1748,In_605,In_2478);
or U1749 (N_1749,In_1259,In_1321);
nand U1750 (N_1750,In_590,In_2214);
nand U1751 (N_1751,In_1218,In_2225);
xnor U1752 (N_1752,In_2051,In_133);
and U1753 (N_1753,In_471,In_1295);
xor U1754 (N_1754,In_1547,In_584);
nand U1755 (N_1755,In_1217,In_324);
xor U1756 (N_1756,In_1235,In_204);
nand U1757 (N_1757,In_1572,In_1667);
nor U1758 (N_1758,In_1345,In_1116);
xor U1759 (N_1759,In_2367,In_1130);
and U1760 (N_1760,In_2496,In_31);
nand U1761 (N_1761,In_1817,In_983);
or U1762 (N_1762,In_1529,In_1531);
xnor U1763 (N_1763,In_630,In_1435);
or U1764 (N_1764,In_452,In_2167);
xnor U1765 (N_1765,In_1354,In_1058);
and U1766 (N_1766,In_487,In_1589);
xor U1767 (N_1767,In_1659,In_1658);
nor U1768 (N_1768,In_679,In_140);
xnor U1769 (N_1769,In_969,In_1474);
or U1770 (N_1770,In_472,In_1839);
nor U1771 (N_1771,In_692,In_1978);
nand U1772 (N_1772,In_1956,In_1337);
xor U1773 (N_1773,In_2083,In_326);
or U1774 (N_1774,In_1319,In_123);
xor U1775 (N_1775,In_1565,In_2237);
nand U1776 (N_1776,In_1929,In_321);
and U1777 (N_1777,In_1417,In_1957);
and U1778 (N_1778,In_1475,In_1693);
nand U1779 (N_1779,In_1183,In_1088);
nand U1780 (N_1780,In_882,In_1339);
nor U1781 (N_1781,In_1632,In_1092);
xnor U1782 (N_1782,In_173,In_1537);
or U1783 (N_1783,In_748,In_674);
nor U1784 (N_1784,In_227,In_734);
or U1785 (N_1785,In_417,In_1337);
nand U1786 (N_1786,In_362,In_806);
and U1787 (N_1787,In_1514,In_1576);
and U1788 (N_1788,In_1635,In_1000);
and U1789 (N_1789,In_761,In_591);
nor U1790 (N_1790,In_35,In_1794);
nand U1791 (N_1791,In_1565,In_1527);
and U1792 (N_1792,In_1426,In_401);
and U1793 (N_1793,In_1435,In_1459);
xnor U1794 (N_1794,In_75,In_2296);
or U1795 (N_1795,In_457,In_2144);
and U1796 (N_1796,In_901,In_1817);
xor U1797 (N_1797,In_225,In_1794);
xnor U1798 (N_1798,In_1810,In_684);
nand U1799 (N_1799,In_1722,In_2208);
and U1800 (N_1800,In_2220,In_2257);
or U1801 (N_1801,In_2103,In_1384);
and U1802 (N_1802,In_1416,In_626);
and U1803 (N_1803,In_2448,In_106);
nor U1804 (N_1804,In_571,In_507);
nand U1805 (N_1805,In_1523,In_1725);
or U1806 (N_1806,In_636,In_1367);
or U1807 (N_1807,In_836,In_922);
nor U1808 (N_1808,In_278,In_970);
nor U1809 (N_1809,In_2251,In_2116);
nand U1810 (N_1810,In_1122,In_2421);
xnor U1811 (N_1811,In_1697,In_805);
nor U1812 (N_1812,In_2226,In_1359);
or U1813 (N_1813,In_785,In_783);
xnor U1814 (N_1814,In_1738,In_1336);
or U1815 (N_1815,In_1148,In_476);
and U1816 (N_1816,In_1345,In_150);
nand U1817 (N_1817,In_324,In_136);
and U1818 (N_1818,In_439,In_2114);
or U1819 (N_1819,In_1810,In_357);
nand U1820 (N_1820,In_1924,In_390);
or U1821 (N_1821,In_2478,In_1350);
nand U1822 (N_1822,In_13,In_944);
xnor U1823 (N_1823,In_1341,In_60);
or U1824 (N_1824,In_195,In_98);
xor U1825 (N_1825,In_930,In_1098);
nor U1826 (N_1826,In_1825,In_1190);
xor U1827 (N_1827,In_1341,In_628);
and U1828 (N_1828,In_2404,In_1774);
xnor U1829 (N_1829,In_1108,In_2354);
or U1830 (N_1830,In_1372,In_769);
xnor U1831 (N_1831,In_32,In_1665);
nor U1832 (N_1832,In_1300,In_821);
xnor U1833 (N_1833,In_211,In_1175);
xor U1834 (N_1834,In_445,In_492);
xor U1835 (N_1835,In_1044,In_1454);
and U1836 (N_1836,In_1727,In_134);
nand U1837 (N_1837,In_1649,In_1138);
nand U1838 (N_1838,In_532,In_407);
xor U1839 (N_1839,In_242,In_1004);
or U1840 (N_1840,In_1998,In_419);
nand U1841 (N_1841,In_455,In_1798);
xnor U1842 (N_1842,In_917,In_1068);
nor U1843 (N_1843,In_2079,In_1761);
nand U1844 (N_1844,In_1293,In_1014);
and U1845 (N_1845,In_2010,In_106);
and U1846 (N_1846,In_1466,In_76);
or U1847 (N_1847,In_976,In_1445);
xor U1848 (N_1848,In_420,In_281);
nand U1849 (N_1849,In_1329,In_1508);
or U1850 (N_1850,In_1471,In_2399);
nor U1851 (N_1851,In_1464,In_1167);
and U1852 (N_1852,In_2222,In_972);
nor U1853 (N_1853,In_1870,In_892);
nand U1854 (N_1854,In_2133,In_665);
and U1855 (N_1855,In_1695,In_211);
or U1856 (N_1856,In_770,In_1625);
or U1857 (N_1857,In_1185,In_443);
or U1858 (N_1858,In_787,In_2236);
nand U1859 (N_1859,In_1192,In_761);
xor U1860 (N_1860,In_1043,In_2289);
xnor U1861 (N_1861,In_2199,In_1025);
nand U1862 (N_1862,In_315,In_2002);
or U1863 (N_1863,In_305,In_1354);
nand U1864 (N_1864,In_271,In_70);
or U1865 (N_1865,In_2303,In_772);
and U1866 (N_1866,In_1614,In_1850);
or U1867 (N_1867,In_1102,In_66);
nor U1868 (N_1868,In_2236,In_1002);
and U1869 (N_1869,In_1770,In_143);
xor U1870 (N_1870,In_1144,In_166);
nand U1871 (N_1871,In_212,In_1540);
xor U1872 (N_1872,In_743,In_767);
or U1873 (N_1873,In_1845,In_1170);
nand U1874 (N_1874,In_834,In_850);
or U1875 (N_1875,In_2305,In_1105);
xor U1876 (N_1876,In_589,In_2224);
nand U1877 (N_1877,In_1128,In_854);
or U1878 (N_1878,In_2171,In_837);
nand U1879 (N_1879,In_1169,In_1860);
nor U1880 (N_1880,In_1192,In_864);
or U1881 (N_1881,In_1819,In_2233);
or U1882 (N_1882,In_1354,In_1777);
xnor U1883 (N_1883,In_1626,In_1228);
and U1884 (N_1884,In_911,In_262);
nand U1885 (N_1885,In_1188,In_2424);
xor U1886 (N_1886,In_1550,In_1718);
nor U1887 (N_1887,In_934,In_659);
or U1888 (N_1888,In_412,In_761);
or U1889 (N_1889,In_1454,In_1672);
or U1890 (N_1890,In_1476,In_469);
xnor U1891 (N_1891,In_13,In_716);
nor U1892 (N_1892,In_2082,In_1742);
or U1893 (N_1893,In_1591,In_2096);
or U1894 (N_1894,In_577,In_1908);
nor U1895 (N_1895,In_306,In_202);
or U1896 (N_1896,In_1723,In_2272);
nand U1897 (N_1897,In_975,In_491);
xnor U1898 (N_1898,In_741,In_632);
nor U1899 (N_1899,In_1091,In_2169);
or U1900 (N_1900,In_703,In_1467);
nand U1901 (N_1901,In_171,In_309);
xor U1902 (N_1902,In_2326,In_2357);
nor U1903 (N_1903,In_677,In_1024);
and U1904 (N_1904,In_2108,In_2042);
nand U1905 (N_1905,In_2151,In_2211);
and U1906 (N_1906,In_272,In_993);
and U1907 (N_1907,In_189,In_1211);
nor U1908 (N_1908,In_1162,In_946);
xor U1909 (N_1909,In_1548,In_497);
nand U1910 (N_1910,In_1301,In_1498);
xor U1911 (N_1911,In_31,In_1508);
or U1912 (N_1912,In_1119,In_1664);
xnor U1913 (N_1913,In_136,In_351);
or U1914 (N_1914,In_2016,In_344);
nand U1915 (N_1915,In_1326,In_1916);
xor U1916 (N_1916,In_31,In_1849);
and U1917 (N_1917,In_1021,In_1637);
nor U1918 (N_1918,In_18,In_150);
nor U1919 (N_1919,In_985,In_1936);
and U1920 (N_1920,In_69,In_1769);
nor U1921 (N_1921,In_2099,In_439);
xor U1922 (N_1922,In_2115,In_1036);
or U1923 (N_1923,In_494,In_815);
or U1924 (N_1924,In_2226,In_87);
nor U1925 (N_1925,In_1773,In_1479);
xor U1926 (N_1926,In_42,In_508);
and U1927 (N_1927,In_588,In_1688);
nor U1928 (N_1928,In_1772,In_2377);
or U1929 (N_1929,In_1822,In_2128);
or U1930 (N_1930,In_852,In_1034);
xnor U1931 (N_1931,In_611,In_2426);
or U1932 (N_1932,In_802,In_479);
and U1933 (N_1933,In_377,In_996);
nand U1934 (N_1934,In_1430,In_1209);
xor U1935 (N_1935,In_2249,In_502);
and U1936 (N_1936,In_2062,In_501);
nor U1937 (N_1937,In_1175,In_795);
nand U1938 (N_1938,In_2476,In_30);
and U1939 (N_1939,In_2301,In_2194);
nor U1940 (N_1940,In_1397,In_524);
or U1941 (N_1941,In_697,In_1594);
or U1942 (N_1942,In_443,In_222);
nand U1943 (N_1943,In_1580,In_1512);
nor U1944 (N_1944,In_764,In_982);
or U1945 (N_1945,In_1092,In_1050);
and U1946 (N_1946,In_485,In_418);
and U1947 (N_1947,In_1654,In_1093);
nand U1948 (N_1948,In_1944,In_1438);
nor U1949 (N_1949,In_1856,In_65);
nand U1950 (N_1950,In_14,In_752);
and U1951 (N_1951,In_585,In_1314);
or U1952 (N_1952,In_356,In_997);
and U1953 (N_1953,In_2073,In_1595);
nand U1954 (N_1954,In_636,In_2407);
xnor U1955 (N_1955,In_4,In_227);
nor U1956 (N_1956,In_972,In_1696);
or U1957 (N_1957,In_1773,In_487);
or U1958 (N_1958,In_1315,In_1167);
xnor U1959 (N_1959,In_2125,In_595);
and U1960 (N_1960,In_637,In_2457);
nand U1961 (N_1961,In_366,In_467);
xor U1962 (N_1962,In_1066,In_442);
nand U1963 (N_1963,In_867,In_2020);
nor U1964 (N_1964,In_2203,In_1441);
xor U1965 (N_1965,In_1247,In_681);
and U1966 (N_1966,In_1905,In_535);
nand U1967 (N_1967,In_961,In_1688);
or U1968 (N_1968,In_1500,In_1547);
nand U1969 (N_1969,In_1188,In_829);
and U1970 (N_1970,In_2067,In_1448);
xor U1971 (N_1971,In_1395,In_2145);
or U1972 (N_1972,In_1468,In_1373);
and U1973 (N_1973,In_484,In_468);
nand U1974 (N_1974,In_2346,In_2298);
and U1975 (N_1975,In_1643,In_1115);
or U1976 (N_1976,In_2490,In_29);
nor U1977 (N_1977,In_1762,In_2397);
nand U1978 (N_1978,In_1373,In_800);
xor U1979 (N_1979,In_273,In_233);
and U1980 (N_1980,In_673,In_2263);
or U1981 (N_1981,In_2248,In_504);
nand U1982 (N_1982,In_1807,In_137);
nor U1983 (N_1983,In_887,In_687);
and U1984 (N_1984,In_117,In_1072);
or U1985 (N_1985,In_1536,In_669);
nand U1986 (N_1986,In_2357,In_660);
xnor U1987 (N_1987,In_1718,In_2024);
nor U1988 (N_1988,In_2226,In_180);
xor U1989 (N_1989,In_1255,In_1576);
or U1990 (N_1990,In_1597,In_717);
or U1991 (N_1991,In_921,In_2149);
xnor U1992 (N_1992,In_166,In_2009);
nand U1993 (N_1993,In_1342,In_529);
xnor U1994 (N_1994,In_883,In_1341);
nor U1995 (N_1995,In_960,In_1968);
and U1996 (N_1996,In_2325,In_349);
xnor U1997 (N_1997,In_323,In_1270);
xor U1998 (N_1998,In_1450,In_1892);
and U1999 (N_1999,In_1601,In_281);
xnor U2000 (N_2000,In_2146,In_261);
xor U2001 (N_2001,In_2423,In_794);
and U2002 (N_2002,In_632,In_2483);
xnor U2003 (N_2003,In_2348,In_1539);
nand U2004 (N_2004,In_1399,In_2207);
or U2005 (N_2005,In_1795,In_727);
nor U2006 (N_2006,In_1308,In_2248);
nand U2007 (N_2007,In_2255,In_1425);
nor U2008 (N_2008,In_1435,In_277);
nor U2009 (N_2009,In_587,In_1499);
and U2010 (N_2010,In_659,In_51);
or U2011 (N_2011,In_1847,In_601);
xnor U2012 (N_2012,In_2274,In_893);
nand U2013 (N_2013,In_1005,In_674);
and U2014 (N_2014,In_1202,In_1449);
and U2015 (N_2015,In_2386,In_1491);
and U2016 (N_2016,In_2022,In_1871);
and U2017 (N_2017,In_1896,In_934);
and U2018 (N_2018,In_1863,In_726);
xor U2019 (N_2019,In_1691,In_1951);
xnor U2020 (N_2020,In_1815,In_705);
and U2021 (N_2021,In_10,In_1079);
and U2022 (N_2022,In_2482,In_1765);
nor U2023 (N_2023,In_2187,In_110);
and U2024 (N_2024,In_185,In_991);
or U2025 (N_2025,In_1422,In_973);
or U2026 (N_2026,In_1804,In_1559);
nand U2027 (N_2027,In_2081,In_507);
xnor U2028 (N_2028,In_525,In_1850);
and U2029 (N_2029,In_2393,In_1127);
or U2030 (N_2030,In_427,In_1056);
and U2031 (N_2031,In_1709,In_737);
nor U2032 (N_2032,In_2157,In_368);
or U2033 (N_2033,In_130,In_87);
or U2034 (N_2034,In_1518,In_541);
nor U2035 (N_2035,In_456,In_1863);
xnor U2036 (N_2036,In_2372,In_1803);
or U2037 (N_2037,In_1387,In_1725);
or U2038 (N_2038,In_2246,In_428);
nand U2039 (N_2039,In_2233,In_1319);
and U2040 (N_2040,In_713,In_605);
nand U2041 (N_2041,In_2483,In_2356);
and U2042 (N_2042,In_1485,In_1029);
nand U2043 (N_2043,In_2047,In_2488);
xnor U2044 (N_2044,In_552,In_2248);
and U2045 (N_2045,In_1934,In_986);
xor U2046 (N_2046,In_502,In_1766);
or U2047 (N_2047,In_873,In_1920);
nor U2048 (N_2048,In_423,In_1778);
and U2049 (N_2049,In_2144,In_2313);
nand U2050 (N_2050,In_248,In_1875);
and U2051 (N_2051,In_338,In_1632);
nand U2052 (N_2052,In_1413,In_913);
nand U2053 (N_2053,In_1354,In_585);
nand U2054 (N_2054,In_1153,In_1168);
or U2055 (N_2055,In_1779,In_1686);
or U2056 (N_2056,In_2294,In_1062);
nand U2057 (N_2057,In_1338,In_1370);
or U2058 (N_2058,In_441,In_418);
or U2059 (N_2059,In_1302,In_509);
xnor U2060 (N_2060,In_1938,In_1356);
or U2061 (N_2061,In_112,In_1104);
nand U2062 (N_2062,In_1421,In_489);
or U2063 (N_2063,In_753,In_1585);
or U2064 (N_2064,In_2106,In_926);
or U2065 (N_2065,In_1809,In_1277);
nand U2066 (N_2066,In_300,In_2059);
xnor U2067 (N_2067,In_1116,In_2257);
nand U2068 (N_2068,In_1857,In_1700);
or U2069 (N_2069,In_877,In_401);
and U2070 (N_2070,In_1408,In_381);
and U2071 (N_2071,In_784,In_981);
xor U2072 (N_2072,In_2339,In_623);
nor U2073 (N_2073,In_1272,In_311);
nor U2074 (N_2074,In_1198,In_881);
and U2075 (N_2075,In_1305,In_843);
nand U2076 (N_2076,In_2141,In_263);
xnor U2077 (N_2077,In_935,In_171);
and U2078 (N_2078,In_1917,In_886);
nand U2079 (N_2079,In_7,In_1900);
nor U2080 (N_2080,In_506,In_1542);
or U2081 (N_2081,In_2463,In_2205);
nand U2082 (N_2082,In_1228,In_1463);
and U2083 (N_2083,In_10,In_1335);
nor U2084 (N_2084,In_2233,In_378);
nor U2085 (N_2085,In_2157,In_2277);
or U2086 (N_2086,In_761,In_1733);
and U2087 (N_2087,In_2488,In_869);
and U2088 (N_2088,In_1553,In_294);
or U2089 (N_2089,In_2004,In_1374);
and U2090 (N_2090,In_2027,In_1381);
or U2091 (N_2091,In_1124,In_2250);
xnor U2092 (N_2092,In_1513,In_757);
nand U2093 (N_2093,In_1970,In_1378);
nand U2094 (N_2094,In_1179,In_1953);
xnor U2095 (N_2095,In_1280,In_362);
and U2096 (N_2096,In_1206,In_1916);
and U2097 (N_2097,In_904,In_1246);
xnor U2098 (N_2098,In_2288,In_1186);
nand U2099 (N_2099,In_2379,In_1563);
nor U2100 (N_2100,In_1388,In_813);
nand U2101 (N_2101,In_1307,In_1428);
or U2102 (N_2102,In_2390,In_459);
nor U2103 (N_2103,In_1984,In_11);
and U2104 (N_2104,In_727,In_1156);
nor U2105 (N_2105,In_84,In_2252);
nor U2106 (N_2106,In_1866,In_2260);
xnor U2107 (N_2107,In_1118,In_2288);
or U2108 (N_2108,In_1928,In_206);
or U2109 (N_2109,In_1937,In_2374);
nor U2110 (N_2110,In_1767,In_898);
or U2111 (N_2111,In_1608,In_2041);
or U2112 (N_2112,In_2080,In_2322);
nand U2113 (N_2113,In_464,In_1476);
or U2114 (N_2114,In_2271,In_1161);
nor U2115 (N_2115,In_1027,In_1531);
or U2116 (N_2116,In_2052,In_1555);
xnor U2117 (N_2117,In_1520,In_883);
nor U2118 (N_2118,In_568,In_1227);
or U2119 (N_2119,In_1818,In_924);
nor U2120 (N_2120,In_1423,In_290);
or U2121 (N_2121,In_376,In_1699);
or U2122 (N_2122,In_84,In_188);
or U2123 (N_2123,In_968,In_1232);
or U2124 (N_2124,In_1587,In_1038);
nor U2125 (N_2125,In_1360,In_928);
and U2126 (N_2126,In_2075,In_58);
nor U2127 (N_2127,In_319,In_135);
xor U2128 (N_2128,In_362,In_911);
nand U2129 (N_2129,In_1103,In_2374);
nand U2130 (N_2130,In_1937,In_1238);
xnor U2131 (N_2131,In_1201,In_477);
and U2132 (N_2132,In_387,In_2133);
xor U2133 (N_2133,In_642,In_1783);
and U2134 (N_2134,In_1291,In_1019);
nor U2135 (N_2135,In_424,In_460);
and U2136 (N_2136,In_664,In_2300);
nand U2137 (N_2137,In_462,In_172);
and U2138 (N_2138,In_1411,In_1283);
nor U2139 (N_2139,In_300,In_77);
nor U2140 (N_2140,In_1407,In_1402);
nor U2141 (N_2141,In_1684,In_918);
nor U2142 (N_2142,In_222,In_835);
nor U2143 (N_2143,In_1790,In_901);
nor U2144 (N_2144,In_1711,In_1848);
nor U2145 (N_2145,In_989,In_229);
xor U2146 (N_2146,In_1942,In_1084);
nand U2147 (N_2147,In_204,In_633);
nand U2148 (N_2148,In_2226,In_1973);
nand U2149 (N_2149,In_1082,In_619);
nand U2150 (N_2150,In_220,In_2037);
nor U2151 (N_2151,In_1151,In_1619);
nor U2152 (N_2152,In_2275,In_1848);
xor U2153 (N_2153,In_316,In_2381);
or U2154 (N_2154,In_1096,In_1684);
nand U2155 (N_2155,In_961,In_2335);
or U2156 (N_2156,In_997,In_432);
nand U2157 (N_2157,In_2216,In_1624);
xnor U2158 (N_2158,In_1291,In_2011);
and U2159 (N_2159,In_2290,In_1097);
xor U2160 (N_2160,In_1982,In_1552);
nor U2161 (N_2161,In_253,In_2456);
xor U2162 (N_2162,In_1480,In_1991);
and U2163 (N_2163,In_482,In_542);
and U2164 (N_2164,In_1000,In_2015);
xnor U2165 (N_2165,In_424,In_2468);
nor U2166 (N_2166,In_45,In_1050);
or U2167 (N_2167,In_187,In_837);
nand U2168 (N_2168,In_868,In_1406);
nor U2169 (N_2169,In_89,In_1236);
nor U2170 (N_2170,In_681,In_1885);
or U2171 (N_2171,In_2029,In_2006);
and U2172 (N_2172,In_532,In_1726);
or U2173 (N_2173,In_2012,In_2199);
nor U2174 (N_2174,In_1971,In_1145);
xnor U2175 (N_2175,In_2402,In_2389);
nor U2176 (N_2176,In_207,In_1978);
and U2177 (N_2177,In_604,In_2429);
nor U2178 (N_2178,In_823,In_981);
nor U2179 (N_2179,In_981,In_679);
or U2180 (N_2180,In_1430,In_1758);
or U2181 (N_2181,In_1033,In_115);
and U2182 (N_2182,In_1129,In_994);
and U2183 (N_2183,In_1959,In_741);
or U2184 (N_2184,In_1715,In_1735);
and U2185 (N_2185,In_1151,In_1812);
nand U2186 (N_2186,In_742,In_999);
nor U2187 (N_2187,In_619,In_1994);
and U2188 (N_2188,In_1442,In_1997);
nand U2189 (N_2189,In_560,In_2443);
nand U2190 (N_2190,In_2284,In_862);
or U2191 (N_2191,In_875,In_215);
nand U2192 (N_2192,In_1717,In_2450);
nand U2193 (N_2193,In_1075,In_2094);
xor U2194 (N_2194,In_303,In_1047);
nor U2195 (N_2195,In_224,In_1878);
nor U2196 (N_2196,In_1362,In_919);
or U2197 (N_2197,In_974,In_1889);
or U2198 (N_2198,In_1433,In_1148);
or U2199 (N_2199,In_1562,In_614);
nor U2200 (N_2200,In_283,In_2086);
and U2201 (N_2201,In_402,In_1621);
or U2202 (N_2202,In_2020,In_1401);
or U2203 (N_2203,In_1845,In_501);
nor U2204 (N_2204,In_2039,In_2153);
or U2205 (N_2205,In_809,In_1878);
nand U2206 (N_2206,In_976,In_920);
nand U2207 (N_2207,In_450,In_2388);
or U2208 (N_2208,In_1779,In_1311);
and U2209 (N_2209,In_52,In_225);
or U2210 (N_2210,In_2347,In_2252);
nor U2211 (N_2211,In_334,In_967);
nor U2212 (N_2212,In_143,In_289);
and U2213 (N_2213,In_2111,In_1433);
nand U2214 (N_2214,In_1924,In_424);
xnor U2215 (N_2215,In_91,In_543);
nor U2216 (N_2216,In_1137,In_1009);
nor U2217 (N_2217,In_858,In_1277);
or U2218 (N_2218,In_1762,In_1821);
and U2219 (N_2219,In_477,In_236);
xor U2220 (N_2220,In_1290,In_686);
xor U2221 (N_2221,In_1955,In_794);
nor U2222 (N_2222,In_1990,In_1982);
or U2223 (N_2223,In_244,In_1550);
nand U2224 (N_2224,In_1895,In_60);
nand U2225 (N_2225,In_652,In_129);
or U2226 (N_2226,In_539,In_843);
nor U2227 (N_2227,In_1368,In_2033);
or U2228 (N_2228,In_705,In_832);
or U2229 (N_2229,In_1221,In_1804);
nor U2230 (N_2230,In_1712,In_381);
nand U2231 (N_2231,In_1730,In_2039);
or U2232 (N_2232,In_1962,In_2318);
nand U2233 (N_2233,In_718,In_280);
and U2234 (N_2234,In_1328,In_120);
or U2235 (N_2235,In_285,In_2399);
and U2236 (N_2236,In_1557,In_1864);
nor U2237 (N_2237,In_2372,In_2137);
and U2238 (N_2238,In_801,In_2477);
or U2239 (N_2239,In_784,In_995);
and U2240 (N_2240,In_1854,In_54);
xor U2241 (N_2241,In_1853,In_2172);
nor U2242 (N_2242,In_2063,In_1939);
nor U2243 (N_2243,In_1730,In_46);
xor U2244 (N_2244,In_704,In_661);
nor U2245 (N_2245,In_333,In_259);
nand U2246 (N_2246,In_178,In_1224);
xor U2247 (N_2247,In_1780,In_1599);
and U2248 (N_2248,In_371,In_866);
and U2249 (N_2249,In_2306,In_1052);
or U2250 (N_2250,In_431,In_1637);
or U2251 (N_2251,In_917,In_2485);
xnor U2252 (N_2252,In_1203,In_1455);
and U2253 (N_2253,In_107,In_433);
or U2254 (N_2254,In_498,In_320);
xor U2255 (N_2255,In_442,In_887);
and U2256 (N_2256,In_2271,In_1210);
or U2257 (N_2257,In_503,In_729);
or U2258 (N_2258,In_344,In_1030);
nor U2259 (N_2259,In_1190,In_473);
nand U2260 (N_2260,In_290,In_1467);
xnor U2261 (N_2261,In_1289,In_1864);
and U2262 (N_2262,In_1126,In_2021);
xor U2263 (N_2263,In_434,In_1390);
and U2264 (N_2264,In_1629,In_1895);
and U2265 (N_2265,In_114,In_724);
xor U2266 (N_2266,In_2041,In_1223);
nand U2267 (N_2267,In_1841,In_1334);
and U2268 (N_2268,In_1509,In_1697);
nor U2269 (N_2269,In_1331,In_1498);
and U2270 (N_2270,In_1783,In_47);
and U2271 (N_2271,In_2324,In_27);
xnor U2272 (N_2272,In_518,In_254);
or U2273 (N_2273,In_2397,In_2086);
nand U2274 (N_2274,In_646,In_1027);
or U2275 (N_2275,In_2234,In_2330);
and U2276 (N_2276,In_741,In_1825);
nand U2277 (N_2277,In_627,In_1192);
and U2278 (N_2278,In_1642,In_1764);
xor U2279 (N_2279,In_51,In_702);
nor U2280 (N_2280,In_1456,In_455);
and U2281 (N_2281,In_2319,In_539);
xor U2282 (N_2282,In_2450,In_2115);
or U2283 (N_2283,In_624,In_692);
nand U2284 (N_2284,In_818,In_370);
nand U2285 (N_2285,In_1505,In_1512);
xnor U2286 (N_2286,In_1046,In_1119);
nand U2287 (N_2287,In_1816,In_982);
xnor U2288 (N_2288,In_825,In_425);
or U2289 (N_2289,In_209,In_1354);
xnor U2290 (N_2290,In_2289,In_1376);
or U2291 (N_2291,In_899,In_195);
xnor U2292 (N_2292,In_780,In_2289);
xor U2293 (N_2293,In_1740,In_1246);
nand U2294 (N_2294,In_1561,In_2334);
and U2295 (N_2295,In_2269,In_1551);
nor U2296 (N_2296,In_2188,In_2158);
or U2297 (N_2297,In_2305,In_2441);
nor U2298 (N_2298,In_591,In_2446);
nand U2299 (N_2299,In_58,In_2053);
nand U2300 (N_2300,In_2344,In_406);
or U2301 (N_2301,In_1734,In_2091);
nand U2302 (N_2302,In_787,In_1069);
and U2303 (N_2303,In_1291,In_132);
or U2304 (N_2304,In_206,In_678);
or U2305 (N_2305,In_1764,In_2480);
xnor U2306 (N_2306,In_2008,In_423);
xor U2307 (N_2307,In_187,In_968);
or U2308 (N_2308,In_718,In_320);
nor U2309 (N_2309,In_1288,In_789);
nor U2310 (N_2310,In_220,In_822);
and U2311 (N_2311,In_1999,In_2447);
nand U2312 (N_2312,In_1351,In_1017);
nand U2313 (N_2313,In_1247,In_1630);
and U2314 (N_2314,In_1514,In_213);
or U2315 (N_2315,In_2352,In_508);
nor U2316 (N_2316,In_184,In_532);
and U2317 (N_2317,In_1659,In_2273);
and U2318 (N_2318,In_1307,In_2204);
xnor U2319 (N_2319,In_1190,In_1599);
and U2320 (N_2320,In_2422,In_971);
or U2321 (N_2321,In_810,In_1182);
and U2322 (N_2322,In_651,In_421);
or U2323 (N_2323,In_2497,In_667);
and U2324 (N_2324,In_1360,In_2471);
xnor U2325 (N_2325,In_837,In_1544);
nand U2326 (N_2326,In_1959,In_1475);
and U2327 (N_2327,In_1536,In_847);
nor U2328 (N_2328,In_1396,In_1093);
or U2329 (N_2329,In_47,In_2426);
nand U2330 (N_2330,In_2299,In_1439);
nand U2331 (N_2331,In_2383,In_1369);
nand U2332 (N_2332,In_1002,In_771);
nand U2333 (N_2333,In_1824,In_68);
nand U2334 (N_2334,In_1969,In_2157);
or U2335 (N_2335,In_1504,In_108);
or U2336 (N_2336,In_2125,In_56);
or U2337 (N_2337,In_953,In_1799);
nand U2338 (N_2338,In_2107,In_1291);
xnor U2339 (N_2339,In_2095,In_1016);
xnor U2340 (N_2340,In_1223,In_270);
nand U2341 (N_2341,In_1619,In_178);
and U2342 (N_2342,In_1366,In_986);
nor U2343 (N_2343,In_233,In_2387);
and U2344 (N_2344,In_291,In_824);
or U2345 (N_2345,In_128,In_1253);
or U2346 (N_2346,In_962,In_2195);
and U2347 (N_2347,In_100,In_495);
nor U2348 (N_2348,In_1676,In_1427);
nand U2349 (N_2349,In_2269,In_938);
nor U2350 (N_2350,In_125,In_707);
nor U2351 (N_2351,In_786,In_411);
xor U2352 (N_2352,In_106,In_1424);
and U2353 (N_2353,In_283,In_2257);
or U2354 (N_2354,In_961,In_1175);
nand U2355 (N_2355,In_1242,In_2028);
xnor U2356 (N_2356,In_894,In_850);
nor U2357 (N_2357,In_1971,In_463);
and U2358 (N_2358,In_1802,In_1509);
xor U2359 (N_2359,In_1935,In_434);
or U2360 (N_2360,In_2264,In_441);
nor U2361 (N_2361,In_2013,In_2291);
and U2362 (N_2362,In_1658,In_1930);
and U2363 (N_2363,In_470,In_1243);
nor U2364 (N_2364,In_2249,In_2376);
xor U2365 (N_2365,In_1864,In_1717);
or U2366 (N_2366,In_1525,In_1711);
xor U2367 (N_2367,In_786,In_659);
or U2368 (N_2368,In_324,In_740);
nor U2369 (N_2369,In_2122,In_604);
nand U2370 (N_2370,In_1029,In_1876);
nor U2371 (N_2371,In_2165,In_372);
nor U2372 (N_2372,In_2372,In_1456);
or U2373 (N_2373,In_1194,In_2013);
nor U2374 (N_2374,In_2490,In_2133);
nor U2375 (N_2375,In_1733,In_823);
nand U2376 (N_2376,In_1777,In_1794);
nand U2377 (N_2377,In_2157,In_956);
nand U2378 (N_2378,In_1812,In_1134);
and U2379 (N_2379,In_676,In_520);
or U2380 (N_2380,In_1503,In_996);
nor U2381 (N_2381,In_173,In_291);
and U2382 (N_2382,In_372,In_283);
xor U2383 (N_2383,In_1484,In_1082);
and U2384 (N_2384,In_2222,In_788);
and U2385 (N_2385,In_232,In_74);
and U2386 (N_2386,In_2408,In_1367);
nand U2387 (N_2387,In_1817,In_213);
nand U2388 (N_2388,In_1817,In_265);
nand U2389 (N_2389,In_707,In_950);
nand U2390 (N_2390,In_2428,In_1322);
or U2391 (N_2391,In_961,In_591);
nand U2392 (N_2392,In_1019,In_139);
nor U2393 (N_2393,In_315,In_2038);
nand U2394 (N_2394,In_2227,In_1693);
and U2395 (N_2395,In_1005,In_1358);
or U2396 (N_2396,In_0,In_2302);
xor U2397 (N_2397,In_1751,In_2373);
nand U2398 (N_2398,In_1260,In_2487);
and U2399 (N_2399,In_1889,In_2214);
nor U2400 (N_2400,In_1302,In_577);
nor U2401 (N_2401,In_491,In_819);
and U2402 (N_2402,In_2011,In_1594);
nand U2403 (N_2403,In_1080,In_1674);
nor U2404 (N_2404,In_501,In_1321);
nand U2405 (N_2405,In_148,In_171);
nand U2406 (N_2406,In_988,In_45);
nor U2407 (N_2407,In_575,In_2445);
and U2408 (N_2408,In_798,In_2257);
xor U2409 (N_2409,In_124,In_1480);
nor U2410 (N_2410,In_269,In_1614);
nand U2411 (N_2411,In_2303,In_752);
or U2412 (N_2412,In_2447,In_599);
or U2413 (N_2413,In_262,In_1990);
and U2414 (N_2414,In_80,In_362);
nand U2415 (N_2415,In_750,In_1771);
nand U2416 (N_2416,In_420,In_1518);
nor U2417 (N_2417,In_3,In_2174);
nor U2418 (N_2418,In_650,In_602);
nand U2419 (N_2419,In_1264,In_1779);
or U2420 (N_2420,In_2274,In_1739);
xnor U2421 (N_2421,In_189,In_138);
or U2422 (N_2422,In_46,In_1483);
or U2423 (N_2423,In_1720,In_643);
nor U2424 (N_2424,In_806,In_2311);
or U2425 (N_2425,In_2441,In_310);
and U2426 (N_2426,In_1001,In_1318);
and U2427 (N_2427,In_1802,In_1881);
nand U2428 (N_2428,In_2442,In_1625);
and U2429 (N_2429,In_1868,In_1107);
nor U2430 (N_2430,In_231,In_125);
nor U2431 (N_2431,In_1693,In_2176);
nand U2432 (N_2432,In_1322,In_2481);
nand U2433 (N_2433,In_1563,In_2055);
xor U2434 (N_2434,In_1485,In_449);
nor U2435 (N_2435,In_2484,In_2160);
nand U2436 (N_2436,In_1365,In_786);
or U2437 (N_2437,In_608,In_1962);
xor U2438 (N_2438,In_310,In_13);
or U2439 (N_2439,In_1506,In_11);
nor U2440 (N_2440,In_1809,In_121);
nand U2441 (N_2441,In_2296,In_2381);
nor U2442 (N_2442,In_2030,In_1675);
or U2443 (N_2443,In_1651,In_1916);
nand U2444 (N_2444,In_972,In_331);
nand U2445 (N_2445,In_256,In_1289);
and U2446 (N_2446,In_1851,In_1208);
nor U2447 (N_2447,In_1175,In_985);
or U2448 (N_2448,In_310,In_266);
and U2449 (N_2449,In_1551,In_1931);
nand U2450 (N_2450,In_1726,In_2361);
nor U2451 (N_2451,In_2466,In_1679);
xnor U2452 (N_2452,In_189,In_1434);
and U2453 (N_2453,In_1424,In_1730);
xor U2454 (N_2454,In_1458,In_1247);
or U2455 (N_2455,In_856,In_1273);
xor U2456 (N_2456,In_108,In_690);
xnor U2457 (N_2457,In_1462,In_898);
or U2458 (N_2458,In_2212,In_863);
xnor U2459 (N_2459,In_1549,In_1352);
or U2460 (N_2460,In_138,In_2204);
or U2461 (N_2461,In_1575,In_203);
xnor U2462 (N_2462,In_1940,In_860);
xor U2463 (N_2463,In_1375,In_1397);
and U2464 (N_2464,In_1384,In_121);
nand U2465 (N_2465,In_2278,In_858);
nor U2466 (N_2466,In_2383,In_416);
xor U2467 (N_2467,In_1904,In_610);
nor U2468 (N_2468,In_1652,In_1861);
or U2469 (N_2469,In_9,In_1982);
nor U2470 (N_2470,In_893,In_1763);
xor U2471 (N_2471,In_2199,In_1123);
xor U2472 (N_2472,In_1029,In_1940);
and U2473 (N_2473,In_2231,In_2187);
or U2474 (N_2474,In_1218,In_1479);
or U2475 (N_2475,In_652,In_1317);
xnor U2476 (N_2476,In_1981,In_636);
and U2477 (N_2477,In_2318,In_361);
xnor U2478 (N_2478,In_1781,In_506);
and U2479 (N_2479,In_918,In_862);
or U2480 (N_2480,In_1322,In_1393);
xnor U2481 (N_2481,In_1303,In_857);
xnor U2482 (N_2482,In_2148,In_1298);
and U2483 (N_2483,In_1821,In_1172);
and U2484 (N_2484,In_1101,In_2369);
nor U2485 (N_2485,In_732,In_771);
or U2486 (N_2486,In_2059,In_1419);
or U2487 (N_2487,In_446,In_2392);
nor U2488 (N_2488,In_453,In_88);
nor U2489 (N_2489,In_998,In_1995);
and U2490 (N_2490,In_1265,In_1348);
xor U2491 (N_2491,In_2492,In_444);
or U2492 (N_2492,In_1670,In_252);
xor U2493 (N_2493,In_128,In_927);
nand U2494 (N_2494,In_1590,In_2452);
and U2495 (N_2495,In_1474,In_738);
nand U2496 (N_2496,In_1002,In_928);
and U2497 (N_2497,In_1054,In_1297);
nor U2498 (N_2498,In_1545,In_1607);
and U2499 (N_2499,In_1686,In_1495);
xnor U2500 (N_2500,In_1351,In_2188);
nor U2501 (N_2501,In_1143,In_390);
nor U2502 (N_2502,In_124,In_189);
xor U2503 (N_2503,In_65,In_1463);
or U2504 (N_2504,In_1853,In_556);
xor U2505 (N_2505,In_1922,In_275);
nor U2506 (N_2506,In_1069,In_1351);
xor U2507 (N_2507,In_2387,In_185);
nor U2508 (N_2508,In_1268,In_2415);
or U2509 (N_2509,In_224,In_1591);
nand U2510 (N_2510,In_596,In_1034);
xnor U2511 (N_2511,In_2366,In_845);
nor U2512 (N_2512,In_1459,In_922);
and U2513 (N_2513,In_1709,In_2403);
nor U2514 (N_2514,In_910,In_343);
and U2515 (N_2515,In_2305,In_187);
nor U2516 (N_2516,In_759,In_801);
and U2517 (N_2517,In_859,In_449);
xor U2518 (N_2518,In_2185,In_1982);
xnor U2519 (N_2519,In_2420,In_2352);
xor U2520 (N_2520,In_327,In_175);
and U2521 (N_2521,In_336,In_454);
nor U2522 (N_2522,In_1731,In_1289);
xnor U2523 (N_2523,In_71,In_1672);
nor U2524 (N_2524,In_1778,In_1285);
nand U2525 (N_2525,In_1703,In_49);
or U2526 (N_2526,In_119,In_1442);
nor U2527 (N_2527,In_1633,In_1748);
and U2528 (N_2528,In_1413,In_366);
and U2529 (N_2529,In_400,In_2128);
nor U2530 (N_2530,In_1474,In_1589);
nand U2531 (N_2531,In_1930,In_1387);
nor U2532 (N_2532,In_135,In_1626);
nand U2533 (N_2533,In_678,In_1324);
nand U2534 (N_2534,In_1751,In_825);
nand U2535 (N_2535,In_1767,In_1172);
nor U2536 (N_2536,In_1893,In_2275);
nor U2537 (N_2537,In_736,In_2114);
or U2538 (N_2538,In_101,In_443);
xor U2539 (N_2539,In_1775,In_477);
or U2540 (N_2540,In_1287,In_2183);
nor U2541 (N_2541,In_1866,In_2146);
and U2542 (N_2542,In_2156,In_2445);
nor U2543 (N_2543,In_1636,In_333);
or U2544 (N_2544,In_1268,In_2302);
nor U2545 (N_2545,In_854,In_2060);
xnor U2546 (N_2546,In_1022,In_154);
nand U2547 (N_2547,In_1820,In_2222);
nor U2548 (N_2548,In_729,In_63);
or U2549 (N_2549,In_34,In_279);
xnor U2550 (N_2550,In_770,In_976);
nor U2551 (N_2551,In_1045,In_31);
or U2552 (N_2552,In_1227,In_137);
or U2553 (N_2553,In_2128,In_1754);
nor U2554 (N_2554,In_918,In_1131);
and U2555 (N_2555,In_2386,In_2092);
nor U2556 (N_2556,In_907,In_1200);
or U2557 (N_2557,In_1500,In_231);
nor U2558 (N_2558,In_1647,In_1351);
nor U2559 (N_2559,In_1027,In_678);
xnor U2560 (N_2560,In_327,In_138);
or U2561 (N_2561,In_2207,In_348);
or U2562 (N_2562,In_1967,In_2084);
or U2563 (N_2563,In_1538,In_1193);
nor U2564 (N_2564,In_1189,In_1236);
and U2565 (N_2565,In_1895,In_194);
nor U2566 (N_2566,In_1842,In_471);
or U2567 (N_2567,In_2411,In_373);
nor U2568 (N_2568,In_2276,In_529);
nand U2569 (N_2569,In_2059,In_1360);
and U2570 (N_2570,In_2066,In_2274);
and U2571 (N_2571,In_652,In_713);
and U2572 (N_2572,In_1468,In_294);
nand U2573 (N_2573,In_2455,In_1943);
nor U2574 (N_2574,In_1226,In_1579);
nand U2575 (N_2575,In_386,In_1211);
nand U2576 (N_2576,In_1666,In_1945);
or U2577 (N_2577,In_1816,In_2310);
nor U2578 (N_2578,In_2366,In_2014);
and U2579 (N_2579,In_1594,In_1718);
xor U2580 (N_2580,In_2420,In_895);
nand U2581 (N_2581,In_2294,In_681);
and U2582 (N_2582,In_1806,In_431);
and U2583 (N_2583,In_1879,In_2419);
nor U2584 (N_2584,In_1781,In_1860);
nand U2585 (N_2585,In_571,In_2479);
nand U2586 (N_2586,In_293,In_2290);
or U2587 (N_2587,In_340,In_2395);
or U2588 (N_2588,In_971,In_1415);
and U2589 (N_2589,In_1208,In_568);
or U2590 (N_2590,In_970,In_1646);
or U2591 (N_2591,In_1514,In_1546);
or U2592 (N_2592,In_909,In_2264);
and U2593 (N_2593,In_1115,In_1225);
xor U2594 (N_2594,In_717,In_104);
xor U2595 (N_2595,In_503,In_2049);
or U2596 (N_2596,In_1418,In_2284);
or U2597 (N_2597,In_2234,In_2321);
nand U2598 (N_2598,In_2218,In_270);
or U2599 (N_2599,In_995,In_406);
nor U2600 (N_2600,In_776,In_187);
or U2601 (N_2601,In_642,In_2351);
nor U2602 (N_2602,In_1718,In_2435);
or U2603 (N_2603,In_1902,In_1807);
nand U2604 (N_2604,In_1410,In_19);
xor U2605 (N_2605,In_1670,In_381);
nor U2606 (N_2606,In_35,In_1489);
xnor U2607 (N_2607,In_2467,In_2283);
nand U2608 (N_2608,In_1482,In_288);
nand U2609 (N_2609,In_1965,In_227);
nor U2610 (N_2610,In_1277,In_297);
and U2611 (N_2611,In_1949,In_1803);
nor U2612 (N_2612,In_51,In_2306);
nor U2613 (N_2613,In_1613,In_2000);
xnor U2614 (N_2614,In_755,In_2388);
xnor U2615 (N_2615,In_804,In_984);
and U2616 (N_2616,In_1116,In_2413);
xor U2617 (N_2617,In_1039,In_2049);
nor U2618 (N_2618,In_2274,In_719);
nand U2619 (N_2619,In_545,In_155);
and U2620 (N_2620,In_1434,In_1800);
or U2621 (N_2621,In_910,In_1070);
and U2622 (N_2622,In_993,In_98);
nor U2623 (N_2623,In_2466,In_1828);
or U2624 (N_2624,In_1117,In_1648);
nor U2625 (N_2625,In_818,In_2356);
xnor U2626 (N_2626,In_1797,In_297);
nand U2627 (N_2627,In_1485,In_1692);
xnor U2628 (N_2628,In_798,In_2222);
nand U2629 (N_2629,In_1623,In_831);
xor U2630 (N_2630,In_450,In_558);
xnor U2631 (N_2631,In_1884,In_1098);
nand U2632 (N_2632,In_1526,In_526);
nand U2633 (N_2633,In_1265,In_1036);
nand U2634 (N_2634,In_598,In_572);
nor U2635 (N_2635,In_571,In_2182);
xor U2636 (N_2636,In_1933,In_1075);
nand U2637 (N_2637,In_504,In_2273);
nor U2638 (N_2638,In_1530,In_1486);
or U2639 (N_2639,In_1401,In_18);
or U2640 (N_2640,In_331,In_1680);
or U2641 (N_2641,In_1430,In_1333);
xor U2642 (N_2642,In_16,In_1224);
xnor U2643 (N_2643,In_223,In_1945);
xor U2644 (N_2644,In_135,In_91);
nand U2645 (N_2645,In_1586,In_1072);
nand U2646 (N_2646,In_2210,In_117);
nand U2647 (N_2647,In_589,In_275);
and U2648 (N_2648,In_1231,In_2020);
or U2649 (N_2649,In_1815,In_489);
nor U2650 (N_2650,In_1541,In_2361);
nor U2651 (N_2651,In_2461,In_1189);
and U2652 (N_2652,In_1873,In_474);
xor U2653 (N_2653,In_518,In_2002);
and U2654 (N_2654,In_361,In_238);
nor U2655 (N_2655,In_2495,In_1980);
and U2656 (N_2656,In_1693,In_2333);
xor U2657 (N_2657,In_73,In_1698);
nand U2658 (N_2658,In_1971,In_2356);
or U2659 (N_2659,In_2188,In_2273);
and U2660 (N_2660,In_135,In_2119);
nand U2661 (N_2661,In_970,In_1784);
nor U2662 (N_2662,In_618,In_885);
or U2663 (N_2663,In_224,In_2451);
nor U2664 (N_2664,In_1712,In_963);
and U2665 (N_2665,In_1452,In_2085);
xnor U2666 (N_2666,In_20,In_1100);
xnor U2667 (N_2667,In_1977,In_904);
and U2668 (N_2668,In_302,In_212);
or U2669 (N_2669,In_74,In_694);
and U2670 (N_2670,In_226,In_2203);
nor U2671 (N_2671,In_2244,In_2453);
and U2672 (N_2672,In_1487,In_2358);
or U2673 (N_2673,In_1775,In_422);
xor U2674 (N_2674,In_2064,In_1745);
or U2675 (N_2675,In_1578,In_1074);
nand U2676 (N_2676,In_1152,In_2000);
and U2677 (N_2677,In_1702,In_1376);
xor U2678 (N_2678,In_1065,In_1074);
or U2679 (N_2679,In_952,In_1651);
or U2680 (N_2680,In_2373,In_1596);
and U2681 (N_2681,In_557,In_1911);
and U2682 (N_2682,In_468,In_578);
or U2683 (N_2683,In_1570,In_697);
and U2684 (N_2684,In_473,In_697);
nor U2685 (N_2685,In_697,In_2135);
and U2686 (N_2686,In_1324,In_2022);
nand U2687 (N_2687,In_2059,In_2341);
and U2688 (N_2688,In_1806,In_1537);
or U2689 (N_2689,In_1670,In_1278);
nand U2690 (N_2690,In_1673,In_491);
and U2691 (N_2691,In_190,In_979);
nand U2692 (N_2692,In_2348,In_1000);
nor U2693 (N_2693,In_2483,In_357);
and U2694 (N_2694,In_1518,In_479);
nand U2695 (N_2695,In_717,In_2283);
nand U2696 (N_2696,In_2133,In_1562);
nand U2697 (N_2697,In_1811,In_776);
xor U2698 (N_2698,In_168,In_13);
and U2699 (N_2699,In_2285,In_2132);
xnor U2700 (N_2700,In_1397,In_2320);
or U2701 (N_2701,In_2252,In_1144);
nand U2702 (N_2702,In_65,In_265);
xnor U2703 (N_2703,In_2097,In_1836);
nand U2704 (N_2704,In_633,In_1864);
nor U2705 (N_2705,In_1242,In_1543);
or U2706 (N_2706,In_2301,In_793);
nor U2707 (N_2707,In_2196,In_89);
xor U2708 (N_2708,In_578,In_1181);
or U2709 (N_2709,In_762,In_1660);
or U2710 (N_2710,In_2153,In_2152);
and U2711 (N_2711,In_225,In_1642);
xnor U2712 (N_2712,In_2491,In_788);
nand U2713 (N_2713,In_2287,In_2034);
nand U2714 (N_2714,In_576,In_136);
or U2715 (N_2715,In_1123,In_692);
and U2716 (N_2716,In_392,In_1006);
xor U2717 (N_2717,In_1490,In_1987);
nand U2718 (N_2718,In_1720,In_53);
xnor U2719 (N_2719,In_1148,In_1187);
and U2720 (N_2720,In_1035,In_1943);
nor U2721 (N_2721,In_1700,In_1589);
nand U2722 (N_2722,In_94,In_1786);
nor U2723 (N_2723,In_1278,In_1969);
xnor U2724 (N_2724,In_362,In_1522);
nor U2725 (N_2725,In_1593,In_886);
nand U2726 (N_2726,In_1063,In_402);
or U2727 (N_2727,In_137,In_144);
nand U2728 (N_2728,In_875,In_527);
and U2729 (N_2729,In_1822,In_2474);
nor U2730 (N_2730,In_306,In_705);
nand U2731 (N_2731,In_96,In_1217);
or U2732 (N_2732,In_50,In_2349);
nor U2733 (N_2733,In_2468,In_381);
xor U2734 (N_2734,In_2457,In_312);
nor U2735 (N_2735,In_830,In_1490);
nor U2736 (N_2736,In_1127,In_150);
nor U2737 (N_2737,In_2460,In_1883);
xnor U2738 (N_2738,In_846,In_1582);
nor U2739 (N_2739,In_306,In_752);
nand U2740 (N_2740,In_1780,In_2282);
nor U2741 (N_2741,In_1814,In_2417);
nor U2742 (N_2742,In_799,In_2259);
nor U2743 (N_2743,In_2020,In_2264);
and U2744 (N_2744,In_1786,In_1009);
and U2745 (N_2745,In_1097,In_1460);
xor U2746 (N_2746,In_6,In_1179);
or U2747 (N_2747,In_188,In_1202);
and U2748 (N_2748,In_242,In_32);
nand U2749 (N_2749,In_2026,In_1313);
nand U2750 (N_2750,In_2324,In_270);
nor U2751 (N_2751,In_663,In_1882);
or U2752 (N_2752,In_715,In_1792);
or U2753 (N_2753,In_806,In_1318);
and U2754 (N_2754,In_2088,In_1722);
nor U2755 (N_2755,In_1607,In_2273);
xor U2756 (N_2756,In_2178,In_1196);
and U2757 (N_2757,In_2413,In_954);
and U2758 (N_2758,In_1123,In_239);
nor U2759 (N_2759,In_1362,In_311);
or U2760 (N_2760,In_571,In_1525);
nor U2761 (N_2761,In_1436,In_1827);
or U2762 (N_2762,In_204,In_1953);
nand U2763 (N_2763,In_2442,In_1590);
or U2764 (N_2764,In_1162,In_541);
or U2765 (N_2765,In_947,In_1679);
nor U2766 (N_2766,In_344,In_836);
and U2767 (N_2767,In_1000,In_1204);
nor U2768 (N_2768,In_1908,In_1728);
xor U2769 (N_2769,In_2059,In_836);
and U2770 (N_2770,In_1912,In_1985);
or U2771 (N_2771,In_1332,In_2184);
nor U2772 (N_2772,In_172,In_2372);
xor U2773 (N_2773,In_949,In_1266);
xor U2774 (N_2774,In_731,In_1453);
and U2775 (N_2775,In_477,In_0);
or U2776 (N_2776,In_1792,In_100);
nand U2777 (N_2777,In_397,In_2242);
nand U2778 (N_2778,In_2420,In_651);
or U2779 (N_2779,In_1510,In_1557);
and U2780 (N_2780,In_2115,In_856);
nand U2781 (N_2781,In_25,In_249);
and U2782 (N_2782,In_1942,In_1950);
nor U2783 (N_2783,In_426,In_1936);
xnor U2784 (N_2784,In_1954,In_2035);
xnor U2785 (N_2785,In_913,In_438);
or U2786 (N_2786,In_178,In_1032);
xor U2787 (N_2787,In_761,In_1912);
or U2788 (N_2788,In_1634,In_210);
nor U2789 (N_2789,In_535,In_1549);
nand U2790 (N_2790,In_1782,In_737);
and U2791 (N_2791,In_2368,In_1850);
nand U2792 (N_2792,In_1972,In_139);
or U2793 (N_2793,In_13,In_880);
and U2794 (N_2794,In_359,In_1747);
or U2795 (N_2795,In_2001,In_402);
xnor U2796 (N_2796,In_2386,In_86);
or U2797 (N_2797,In_740,In_1601);
nand U2798 (N_2798,In_2425,In_2045);
nor U2799 (N_2799,In_1528,In_2045);
xor U2800 (N_2800,In_2453,In_305);
nand U2801 (N_2801,In_1869,In_1340);
xor U2802 (N_2802,In_1617,In_1625);
nor U2803 (N_2803,In_1156,In_1249);
and U2804 (N_2804,In_1038,In_1380);
nor U2805 (N_2805,In_425,In_1002);
or U2806 (N_2806,In_172,In_917);
xnor U2807 (N_2807,In_16,In_1690);
xor U2808 (N_2808,In_1384,In_1498);
and U2809 (N_2809,In_1038,In_431);
nand U2810 (N_2810,In_158,In_63);
nand U2811 (N_2811,In_378,In_879);
nor U2812 (N_2812,In_113,In_978);
nand U2813 (N_2813,In_1521,In_1452);
xor U2814 (N_2814,In_419,In_108);
nand U2815 (N_2815,In_2090,In_1317);
nor U2816 (N_2816,In_619,In_64);
and U2817 (N_2817,In_1912,In_2048);
nand U2818 (N_2818,In_2244,In_1913);
xor U2819 (N_2819,In_2372,In_153);
nand U2820 (N_2820,In_2110,In_1319);
xnor U2821 (N_2821,In_784,In_541);
or U2822 (N_2822,In_1307,In_1691);
nor U2823 (N_2823,In_2321,In_904);
or U2824 (N_2824,In_582,In_1500);
or U2825 (N_2825,In_553,In_505);
and U2826 (N_2826,In_1407,In_587);
or U2827 (N_2827,In_741,In_2116);
and U2828 (N_2828,In_2195,In_1665);
or U2829 (N_2829,In_1402,In_1582);
and U2830 (N_2830,In_2057,In_648);
nand U2831 (N_2831,In_262,In_642);
nor U2832 (N_2832,In_673,In_143);
and U2833 (N_2833,In_335,In_814);
or U2834 (N_2834,In_1609,In_1232);
xor U2835 (N_2835,In_755,In_913);
nor U2836 (N_2836,In_1626,In_1897);
nor U2837 (N_2837,In_2222,In_2258);
nor U2838 (N_2838,In_1404,In_2120);
and U2839 (N_2839,In_1892,In_2042);
or U2840 (N_2840,In_2242,In_1068);
xor U2841 (N_2841,In_2197,In_488);
nor U2842 (N_2842,In_1006,In_18);
or U2843 (N_2843,In_48,In_350);
nand U2844 (N_2844,In_1247,In_1405);
nor U2845 (N_2845,In_1888,In_1542);
or U2846 (N_2846,In_2109,In_907);
xnor U2847 (N_2847,In_351,In_2432);
and U2848 (N_2848,In_2167,In_1831);
xnor U2849 (N_2849,In_920,In_26);
xnor U2850 (N_2850,In_774,In_2019);
and U2851 (N_2851,In_1416,In_1987);
and U2852 (N_2852,In_2063,In_370);
or U2853 (N_2853,In_1252,In_1292);
or U2854 (N_2854,In_485,In_171);
nand U2855 (N_2855,In_2422,In_578);
and U2856 (N_2856,In_111,In_2144);
xnor U2857 (N_2857,In_339,In_1160);
xor U2858 (N_2858,In_1688,In_967);
or U2859 (N_2859,In_2078,In_1786);
nand U2860 (N_2860,In_790,In_385);
xnor U2861 (N_2861,In_1052,In_1500);
nand U2862 (N_2862,In_68,In_608);
xor U2863 (N_2863,In_625,In_424);
or U2864 (N_2864,In_1909,In_1657);
and U2865 (N_2865,In_415,In_1266);
and U2866 (N_2866,In_1230,In_1097);
and U2867 (N_2867,In_1339,In_1436);
and U2868 (N_2868,In_2060,In_1390);
nand U2869 (N_2869,In_1586,In_2493);
xnor U2870 (N_2870,In_251,In_140);
xnor U2871 (N_2871,In_2293,In_1850);
or U2872 (N_2872,In_1671,In_1275);
nor U2873 (N_2873,In_1223,In_2267);
nand U2874 (N_2874,In_863,In_1789);
nor U2875 (N_2875,In_1106,In_1968);
or U2876 (N_2876,In_625,In_566);
and U2877 (N_2877,In_1389,In_243);
and U2878 (N_2878,In_1825,In_1313);
nand U2879 (N_2879,In_408,In_801);
nand U2880 (N_2880,In_862,In_1311);
nor U2881 (N_2881,In_517,In_1908);
xnor U2882 (N_2882,In_86,In_585);
or U2883 (N_2883,In_1931,In_2189);
and U2884 (N_2884,In_160,In_1113);
nor U2885 (N_2885,In_604,In_1593);
nor U2886 (N_2886,In_102,In_1370);
and U2887 (N_2887,In_761,In_973);
nand U2888 (N_2888,In_370,In_2171);
nor U2889 (N_2889,In_1923,In_339);
and U2890 (N_2890,In_2296,In_842);
and U2891 (N_2891,In_1755,In_1852);
and U2892 (N_2892,In_897,In_1083);
or U2893 (N_2893,In_2043,In_46);
or U2894 (N_2894,In_180,In_148);
nand U2895 (N_2895,In_0,In_2350);
nor U2896 (N_2896,In_1965,In_1684);
nand U2897 (N_2897,In_1988,In_1222);
nor U2898 (N_2898,In_416,In_2124);
and U2899 (N_2899,In_1858,In_1878);
and U2900 (N_2900,In_1134,In_1058);
nand U2901 (N_2901,In_1464,In_2330);
and U2902 (N_2902,In_388,In_1413);
xor U2903 (N_2903,In_48,In_1208);
and U2904 (N_2904,In_999,In_1731);
nor U2905 (N_2905,In_576,In_2214);
or U2906 (N_2906,In_1692,In_1591);
and U2907 (N_2907,In_739,In_1371);
nand U2908 (N_2908,In_1617,In_652);
nor U2909 (N_2909,In_1781,In_1367);
nor U2910 (N_2910,In_2219,In_943);
or U2911 (N_2911,In_951,In_2379);
and U2912 (N_2912,In_1367,In_56);
xor U2913 (N_2913,In_962,In_1483);
nand U2914 (N_2914,In_1080,In_176);
or U2915 (N_2915,In_726,In_1047);
xor U2916 (N_2916,In_551,In_1368);
and U2917 (N_2917,In_261,In_116);
xnor U2918 (N_2918,In_1031,In_443);
or U2919 (N_2919,In_2428,In_4);
and U2920 (N_2920,In_884,In_283);
xnor U2921 (N_2921,In_1603,In_1855);
xnor U2922 (N_2922,In_2484,In_1507);
nand U2923 (N_2923,In_1842,In_1461);
or U2924 (N_2924,In_505,In_193);
nand U2925 (N_2925,In_892,In_2210);
and U2926 (N_2926,In_828,In_1008);
nor U2927 (N_2927,In_2215,In_695);
or U2928 (N_2928,In_1932,In_2035);
and U2929 (N_2929,In_1628,In_662);
nor U2930 (N_2930,In_966,In_1666);
nand U2931 (N_2931,In_2200,In_488);
or U2932 (N_2932,In_1034,In_1006);
or U2933 (N_2933,In_1836,In_2488);
xnor U2934 (N_2934,In_1813,In_2297);
nand U2935 (N_2935,In_1583,In_1129);
nor U2936 (N_2936,In_964,In_1444);
nor U2937 (N_2937,In_1471,In_2454);
or U2938 (N_2938,In_2397,In_2145);
xor U2939 (N_2939,In_1306,In_1075);
nand U2940 (N_2940,In_1427,In_902);
and U2941 (N_2941,In_1611,In_1529);
or U2942 (N_2942,In_1745,In_2441);
and U2943 (N_2943,In_1488,In_470);
or U2944 (N_2944,In_367,In_1259);
xor U2945 (N_2945,In_1681,In_638);
or U2946 (N_2946,In_945,In_1360);
and U2947 (N_2947,In_1993,In_119);
xor U2948 (N_2948,In_2000,In_161);
or U2949 (N_2949,In_2135,In_437);
nand U2950 (N_2950,In_1187,In_1970);
nand U2951 (N_2951,In_352,In_255);
nor U2952 (N_2952,In_1099,In_327);
or U2953 (N_2953,In_1282,In_2199);
and U2954 (N_2954,In_959,In_1371);
xor U2955 (N_2955,In_1179,In_2296);
or U2956 (N_2956,In_327,In_1378);
nand U2957 (N_2957,In_942,In_1188);
nand U2958 (N_2958,In_2171,In_1872);
nor U2959 (N_2959,In_92,In_1616);
and U2960 (N_2960,In_2380,In_1566);
or U2961 (N_2961,In_1133,In_1169);
and U2962 (N_2962,In_1148,In_744);
nand U2963 (N_2963,In_1130,In_1026);
nand U2964 (N_2964,In_598,In_1165);
xor U2965 (N_2965,In_695,In_2431);
or U2966 (N_2966,In_2254,In_931);
xnor U2967 (N_2967,In_2483,In_708);
or U2968 (N_2968,In_1290,In_315);
nor U2969 (N_2969,In_985,In_1133);
xor U2970 (N_2970,In_843,In_1679);
nand U2971 (N_2971,In_861,In_839);
nor U2972 (N_2972,In_1890,In_1848);
nand U2973 (N_2973,In_1072,In_650);
nand U2974 (N_2974,In_791,In_1011);
and U2975 (N_2975,In_2072,In_1698);
and U2976 (N_2976,In_91,In_337);
or U2977 (N_2977,In_1008,In_1844);
xor U2978 (N_2978,In_77,In_862);
nor U2979 (N_2979,In_2434,In_2399);
or U2980 (N_2980,In_1694,In_2291);
or U2981 (N_2981,In_1034,In_1450);
nor U2982 (N_2982,In_1860,In_2321);
nor U2983 (N_2983,In_2091,In_179);
nor U2984 (N_2984,In_240,In_1700);
xor U2985 (N_2985,In_1401,In_1898);
and U2986 (N_2986,In_1986,In_716);
xor U2987 (N_2987,In_2359,In_65);
nor U2988 (N_2988,In_503,In_1178);
nor U2989 (N_2989,In_575,In_1660);
nor U2990 (N_2990,In_1115,In_512);
xnor U2991 (N_2991,In_1635,In_2482);
xnor U2992 (N_2992,In_2374,In_1661);
xnor U2993 (N_2993,In_920,In_274);
or U2994 (N_2994,In_774,In_2258);
or U2995 (N_2995,In_844,In_119);
xnor U2996 (N_2996,In_1241,In_1354);
or U2997 (N_2997,In_1393,In_418);
and U2998 (N_2998,In_2071,In_2323);
nor U2999 (N_2999,In_248,In_735);
or U3000 (N_3000,In_121,In_348);
or U3001 (N_3001,In_2394,In_1222);
or U3002 (N_3002,In_1683,In_1531);
and U3003 (N_3003,In_2320,In_1904);
xnor U3004 (N_3004,In_2092,In_2086);
nand U3005 (N_3005,In_883,In_954);
nor U3006 (N_3006,In_1757,In_2294);
xnor U3007 (N_3007,In_1910,In_2114);
nand U3008 (N_3008,In_2464,In_620);
and U3009 (N_3009,In_1016,In_511);
xnor U3010 (N_3010,In_2430,In_1506);
nor U3011 (N_3011,In_747,In_154);
and U3012 (N_3012,In_2148,In_1503);
nor U3013 (N_3013,In_1801,In_2390);
and U3014 (N_3014,In_1823,In_873);
nand U3015 (N_3015,In_2406,In_1702);
and U3016 (N_3016,In_942,In_1537);
nand U3017 (N_3017,In_618,In_1859);
or U3018 (N_3018,In_2150,In_869);
and U3019 (N_3019,In_1014,In_2262);
nor U3020 (N_3020,In_1231,In_1056);
nor U3021 (N_3021,In_780,In_1127);
nand U3022 (N_3022,In_1232,In_213);
or U3023 (N_3023,In_2247,In_1079);
xnor U3024 (N_3024,In_2313,In_1766);
xor U3025 (N_3025,In_1286,In_1536);
and U3026 (N_3026,In_954,In_1002);
nor U3027 (N_3027,In_1004,In_2251);
xor U3028 (N_3028,In_154,In_442);
or U3029 (N_3029,In_1115,In_487);
nand U3030 (N_3030,In_758,In_151);
nand U3031 (N_3031,In_468,In_1651);
nand U3032 (N_3032,In_1319,In_32);
xor U3033 (N_3033,In_1392,In_1991);
nand U3034 (N_3034,In_1244,In_1164);
nor U3035 (N_3035,In_603,In_1919);
and U3036 (N_3036,In_1599,In_737);
and U3037 (N_3037,In_1736,In_917);
or U3038 (N_3038,In_1868,In_639);
and U3039 (N_3039,In_1899,In_773);
nor U3040 (N_3040,In_492,In_1588);
and U3041 (N_3041,In_904,In_2076);
and U3042 (N_3042,In_1740,In_1039);
nor U3043 (N_3043,In_1220,In_0);
nand U3044 (N_3044,In_2436,In_846);
nor U3045 (N_3045,In_336,In_2175);
and U3046 (N_3046,In_2181,In_1864);
or U3047 (N_3047,In_116,In_937);
or U3048 (N_3048,In_457,In_1618);
and U3049 (N_3049,In_1314,In_2277);
nor U3050 (N_3050,In_2394,In_503);
xnor U3051 (N_3051,In_875,In_342);
and U3052 (N_3052,In_1725,In_2097);
xor U3053 (N_3053,In_94,In_321);
and U3054 (N_3054,In_2109,In_866);
xnor U3055 (N_3055,In_165,In_1691);
nand U3056 (N_3056,In_1823,In_223);
nor U3057 (N_3057,In_1399,In_1216);
or U3058 (N_3058,In_1198,In_1335);
nor U3059 (N_3059,In_1872,In_1796);
nand U3060 (N_3060,In_589,In_1602);
nor U3061 (N_3061,In_788,In_2359);
nor U3062 (N_3062,In_496,In_1691);
or U3063 (N_3063,In_710,In_1626);
or U3064 (N_3064,In_761,In_2253);
or U3065 (N_3065,In_1991,In_1432);
xnor U3066 (N_3066,In_1492,In_148);
or U3067 (N_3067,In_2171,In_2470);
nor U3068 (N_3068,In_1127,In_2053);
nor U3069 (N_3069,In_1046,In_2387);
nand U3070 (N_3070,In_123,In_1938);
xnor U3071 (N_3071,In_1782,In_2434);
and U3072 (N_3072,In_585,In_870);
nand U3073 (N_3073,In_662,In_1691);
or U3074 (N_3074,In_1734,In_534);
nor U3075 (N_3075,In_1895,In_599);
nor U3076 (N_3076,In_866,In_1790);
or U3077 (N_3077,In_1720,In_471);
nand U3078 (N_3078,In_1519,In_290);
nand U3079 (N_3079,In_1094,In_1684);
and U3080 (N_3080,In_2323,In_2291);
xor U3081 (N_3081,In_1748,In_386);
or U3082 (N_3082,In_2014,In_158);
nand U3083 (N_3083,In_2371,In_1800);
xor U3084 (N_3084,In_694,In_1907);
nand U3085 (N_3085,In_2201,In_1708);
and U3086 (N_3086,In_406,In_1600);
and U3087 (N_3087,In_1197,In_2213);
nor U3088 (N_3088,In_758,In_273);
nand U3089 (N_3089,In_108,In_204);
nand U3090 (N_3090,In_556,In_2153);
nor U3091 (N_3091,In_1731,In_1495);
and U3092 (N_3092,In_313,In_1287);
xor U3093 (N_3093,In_1787,In_221);
nand U3094 (N_3094,In_1584,In_2193);
nand U3095 (N_3095,In_1122,In_945);
nor U3096 (N_3096,In_2202,In_519);
and U3097 (N_3097,In_2237,In_2072);
xnor U3098 (N_3098,In_2374,In_2157);
or U3099 (N_3099,In_516,In_464);
xnor U3100 (N_3100,In_1544,In_1298);
or U3101 (N_3101,In_494,In_1510);
xnor U3102 (N_3102,In_2470,In_975);
or U3103 (N_3103,In_952,In_501);
or U3104 (N_3104,In_1789,In_759);
xnor U3105 (N_3105,In_385,In_1630);
nor U3106 (N_3106,In_66,In_1843);
xor U3107 (N_3107,In_1836,In_278);
and U3108 (N_3108,In_2150,In_1345);
or U3109 (N_3109,In_833,In_1633);
or U3110 (N_3110,In_1310,In_1216);
and U3111 (N_3111,In_604,In_2499);
and U3112 (N_3112,In_800,In_816);
nand U3113 (N_3113,In_211,In_1636);
or U3114 (N_3114,In_723,In_1398);
nor U3115 (N_3115,In_2431,In_617);
xor U3116 (N_3116,In_529,In_48);
xor U3117 (N_3117,In_1926,In_1805);
nor U3118 (N_3118,In_1656,In_1155);
nand U3119 (N_3119,In_926,In_2477);
nor U3120 (N_3120,In_151,In_39);
nor U3121 (N_3121,In_903,In_321);
and U3122 (N_3122,In_1619,In_1212);
nor U3123 (N_3123,In_1669,In_403);
nor U3124 (N_3124,In_2106,In_174);
and U3125 (N_3125,In_1530,In_2387);
xnor U3126 (N_3126,In_1343,In_2278);
nor U3127 (N_3127,In_2131,In_1977);
and U3128 (N_3128,In_1366,In_923);
and U3129 (N_3129,In_434,In_160);
nand U3130 (N_3130,In_1368,In_1621);
xnor U3131 (N_3131,In_1507,In_1178);
and U3132 (N_3132,In_518,In_433);
or U3133 (N_3133,In_1488,In_852);
xor U3134 (N_3134,In_1346,In_2453);
nor U3135 (N_3135,In_1491,In_1465);
nand U3136 (N_3136,In_2306,In_1482);
or U3137 (N_3137,In_1530,In_1225);
xor U3138 (N_3138,In_452,In_1192);
nand U3139 (N_3139,In_2348,In_254);
and U3140 (N_3140,In_1483,In_1346);
xor U3141 (N_3141,In_1795,In_2359);
xor U3142 (N_3142,In_1235,In_1297);
or U3143 (N_3143,In_682,In_968);
nor U3144 (N_3144,In_1211,In_297);
and U3145 (N_3145,In_1364,In_1693);
and U3146 (N_3146,In_600,In_96);
and U3147 (N_3147,In_432,In_1088);
nor U3148 (N_3148,In_737,In_1231);
nor U3149 (N_3149,In_384,In_930);
nor U3150 (N_3150,In_945,In_564);
nand U3151 (N_3151,In_1197,In_1124);
and U3152 (N_3152,In_2048,In_231);
or U3153 (N_3153,In_1137,In_1962);
nor U3154 (N_3154,In_664,In_493);
nor U3155 (N_3155,In_927,In_1072);
xnor U3156 (N_3156,In_2346,In_576);
xor U3157 (N_3157,In_964,In_2364);
or U3158 (N_3158,In_992,In_1297);
or U3159 (N_3159,In_1638,In_1958);
or U3160 (N_3160,In_395,In_1333);
nand U3161 (N_3161,In_2085,In_339);
or U3162 (N_3162,In_2342,In_1286);
or U3163 (N_3163,In_294,In_12);
nor U3164 (N_3164,In_14,In_628);
xnor U3165 (N_3165,In_2101,In_1240);
or U3166 (N_3166,In_2177,In_1456);
nand U3167 (N_3167,In_812,In_125);
or U3168 (N_3168,In_1380,In_913);
nor U3169 (N_3169,In_338,In_1016);
nor U3170 (N_3170,In_2192,In_642);
xnor U3171 (N_3171,In_2475,In_646);
nor U3172 (N_3172,In_2450,In_512);
or U3173 (N_3173,In_1260,In_1880);
and U3174 (N_3174,In_2370,In_1850);
nand U3175 (N_3175,In_1879,In_87);
and U3176 (N_3176,In_1056,In_2202);
and U3177 (N_3177,In_323,In_88);
xor U3178 (N_3178,In_1055,In_2406);
and U3179 (N_3179,In_1659,In_670);
or U3180 (N_3180,In_1470,In_1482);
or U3181 (N_3181,In_2488,In_226);
nand U3182 (N_3182,In_1023,In_1367);
or U3183 (N_3183,In_652,In_343);
nand U3184 (N_3184,In_516,In_1707);
and U3185 (N_3185,In_1596,In_1623);
and U3186 (N_3186,In_2264,In_1524);
nand U3187 (N_3187,In_997,In_2112);
and U3188 (N_3188,In_554,In_1092);
nor U3189 (N_3189,In_951,In_2329);
and U3190 (N_3190,In_2207,In_1096);
or U3191 (N_3191,In_450,In_920);
xnor U3192 (N_3192,In_848,In_150);
nand U3193 (N_3193,In_1220,In_553);
nand U3194 (N_3194,In_1974,In_630);
or U3195 (N_3195,In_2049,In_1979);
nand U3196 (N_3196,In_1764,In_2498);
and U3197 (N_3197,In_1449,In_1319);
or U3198 (N_3198,In_2349,In_73);
or U3199 (N_3199,In_2160,In_232);
and U3200 (N_3200,In_2045,In_1319);
nor U3201 (N_3201,In_794,In_1943);
xor U3202 (N_3202,In_464,In_2218);
or U3203 (N_3203,In_499,In_2193);
nor U3204 (N_3204,In_152,In_372);
and U3205 (N_3205,In_12,In_1930);
nor U3206 (N_3206,In_788,In_706);
and U3207 (N_3207,In_1397,In_2374);
nor U3208 (N_3208,In_1580,In_1828);
nand U3209 (N_3209,In_972,In_1837);
or U3210 (N_3210,In_1792,In_244);
or U3211 (N_3211,In_613,In_60);
nand U3212 (N_3212,In_905,In_836);
nand U3213 (N_3213,In_1724,In_298);
or U3214 (N_3214,In_1782,In_758);
xnor U3215 (N_3215,In_1786,In_2358);
nand U3216 (N_3216,In_800,In_1883);
nor U3217 (N_3217,In_218,In_2223);
and U3218 (N_3218,In_1037,In_366);
or U3219 (N_3219,In_2058,In_1170);
xnor U3220 (N_3220,In_1929,In_1735);
nor U3221 (N_3221,In_1233,In_436);
and U3222 (N_3222,In_1481,In_2428);
nand U3223 (N_3223,In_1303,In_340);
and U3224 (N_3224,In_737,In_1144);
nand U3225 (N_3225,In_1115,In_1701);
or U3226 (N_3226,In_2084,In_1618);
xor U3227 (N_3227,In_1883,In_914);
nand U3228 (N_3228,In_276,In_1548);
nor U3229 (N_3229,In_157,In_113);
xnor U3230 (N_3230,In_1269,In_2169);
or U3231 (N_3231,In_1559,In_1485);
and U3232 (N_3232,In_435,In_445);
xnor U3233 (N_3233,In_858,In_1800);
or U3234 (N_3234,In_954,In_649);
xor U3235 (N_3235,In_57,In_2478);
xnor U3236 (N_3236,In_1233,In_1327);
or U3237 (N_3237,In_1930,In_965);
nor U3238 (N_3238,In_252,In_2420);
nor U3239 (N_3239,In_2176,In_2154);
nor U3240 (N_3240,In_2457,In_464);
xnor U3241 (N_3241,In_1758,In_1992);
or U3242 (N_3242,In_1115,In_216);
or U3243 (N_3243,In_500,In_538);
nor U3244 (N_3244,In_991,In_1618);
nor U3245 (N_3245,In_886,In_1690);
and U3246 (N_3246,In_681,In_1376);
or U3247 (N_3247,In_1789,In_60);
or U3248 (N_3248,In_1982,In_969);
xnor U3249 (N_3249,In_2121,In_516);
xnor U3250 (N_3250,In_1304,In_907);
or U3251 (N_3251,In_1215,In_730);
nor U3252 (N_3252,In_1955,In_1564);
nand U3253 (N_3253,In_843,In_2320);
nand U3254 (N_3254,In_683,In_1343);
nand U3255 (N_3255,In_2256,In_2294);
nor U3256 (N_3256,In_1728,In_647);
xnor U3257 (N_3257,In_1917,In_88);
nand U3258 (N_3258,In_1320,In_2314);
nand U3259 (N_3259,In_1695,In_1308);
xnor U3260 (N_3260,In_2439,In_1448);
nor U3261 (N_3261,In_1572,In_672);
nor U3262 (N_3262,In_2465,In_199);
and U3263 (N_3263,In_1387,In_1101);
or U3264 (N_3264,In_2394,In_359);
nand U3265 (N_3265,In_1649,In_483);
nand U3266 (N_3266,In_396,In_358);
and U3267 (N_3267,In_123,In_604);
xnor U3268 (N_3268,In_1716,In_2238);
and U3269 (N_3269,In_16,In_117);
or U3270 (N_3270,In_1197,In_925);
or U3271 (N_3271,In_959,In_1018);
or U3272 (N_3272,In_738,In_539);
nand U3273 (N_3273,In_980,In_1671);
nand U3274 (N_3274,In_1153,In_495);
nand U3275 (N_3275,In_1492,In_1266);
xor U3276 (N_3276,In_782,In_879);
and U3277 (N_3277,In_1686,In_631);
nand U3278 (N_3278,In_1329,In_1767);
nand U3279 (N_3279,In_1209,In_2240);
nor U3280 (N_3280,In_1335,In_1215);
xor U3281 (N_3281,In_131,In_928);
nand U3282 (N_3282,In_1600,In_1226);
and U3283 (N_3283,In_809,In_789);
xor U3284 (N_3284,In_741,In_656);
and U3285 (N_3285,In_2198,In_359);
or U3286 (N_3286,In_1143,In_1125);
and U3287 (N_3287,In_214,In_1090);
and U3288 (N_3288,In_2243,In_42);
or U3289 (N_3289,In_1399,In_1929);
or U3290 (N_3290,In_1501,In_1901);
xor U3291 (N_3291,In_1573,In_1112);
nor U3292 (N_3292,In_76,In_83);
nand U3293 (N_3293,In_1346,In_2007);
nand U3294 (N_3294,In_873,In_324);
nand U3295 (N_3295,In_1495,In_1984);
xor U3296 (N_3296,In_1375,In_2080);
or U3297 (N_3297,In_2281,In_2418);
or U3298 (N_3298,In_1191,In_958);
xor U3299 (N_3299,In_545,In_806);
nand U3300 (N_3300,In_293,In_483);
xnor U3301 (N_3301,In_2044,In_2363);
xor U3302 (N_3302,In_2494,In_1027);
or U3303 (N_3303,In_1976,In_1119);
nand U3304 (N_3304,In_1577,In_719);
nor U3305 (N_3305,In_518,In_1929);
nand U3306 (N_3306,In_1964,In_395);
xor U3307 (N_3307,In_407,In_681);
xor U3308 (N_3308,In_420,In_310);
nand U3309 (N_3309,In_1462,In_1050);
and U3310 (N_3310,In_260,In_2246);
and U3311 (N_3311,In_1034,In_1915);
nand U3312 (N_3312,In_1458,In_285);
nand U3313 (N_3313,In_2031,In_162);
and U3314 (N_3314,In_717,In_64);
and U3315 (N_3315,In_582,In_645);
and U3316 (N_3316,In_239,In_165);
xor U3317 (N_3317,In_372,In_1778);
nor U3318 (N_3318,In_1794,In_2373);
nand U3319 (N_3319,In_1139,In_1928);
and U3320 (N_3320,In_1720,In_855);
and U3321 (N_3321,In_453,In_2110);
nor U3322 (N_3322,In_2185,In_2123);
xor U3323 (N_3323,In_1465,In_1082);
nand U3324 (N_3324,In_2438,In_2475);
nand U3325 (N_3325,In_2436,In_1077);
nor U3326 (N_3326,In_1823,In_1587);
xnor U3327 (N_3327,In_2122,In_2082);
and U3328 (N_3328,In_959,In_2153);
nand U3329 (N_3329,In_1062,In_2114);
nand U3330 (N_3330,In_126,In_39);
xnor U3331 (N_3331,In_1321,In_478);
xnor U3332 (N_3332,In_382,In_1587);
nor U3333 (N_3333,In_363,In_790);
and U3334 (N_3334,In_2451,In_289);
nor U3335 (N_3335,In_2425,In_1106);
or U3336 (N_3336,In_2406,In_1045);
nor U3337 (N_3337,In_1548,In_1552);
nand U3338 (N_3338,In_2396,In_2373);
and U3339 (N_3339,In_593,In_1577);
xnor U3340 (N_3340,In_1537,In_1692);
nor U3341 (N_3341,In_1642,In_354);
or U3342 (N_3342,In_1890,In_1737);
and U3343 (N_3343,In_1915,In_2048);
nand U3344 (N_3344,In_1630,In_985);
and U3345 (N_3345,In_1857,In_828);
xnor U3346 (N_3346,In_2406,In_1700);
nand U3347 (N_3347,In_1435,In_771);
nor U3348 (N_3348,In_183,In_1834);
xor U3349 (N_3349,In_134,In_951);
and U3350 (N_3350,In_471,In_584);
or U3351 (N_3351,In_596,In_2204);
nor U3352 (N_3352,In_1972,In_1302);
xnor U3353 (N_3353,In_2495,In_2086);
nand U3354 (N_3354,In_1299,In_585);
xnor U3355 (N_3355,In_2051,In_1546);
nor U3356 (N_3356,In_1378,In_4);
nor U3357 (N_3357,In_1765,In_1723);
nand U3358 (N_3358,In_1806,In_900);
nand U3359 (N_3359,In_1707,In_1924);
nor U3360 (N_3360,In_1277,In_1205);
or U3361 (N_3361,In_1442,In_1102);
or U3362 (N_3362,In_552,In_1093);
xnor U3363 (N_3363,In_1959,In_1977);
xor U3364 (N_3364,In_684,In_1272);
or U3365 (N_3365,In_756,In_1196);
and U3366 (N_3366,In_366,In_1674);
xor U3367 (N_3367,In_2271,In_519);
or U3368 (N_3368,In_240,In_2079);
xnor U3369 (N_3369,In_481,In_702);
or U3370 (N_3370,In_1024,In_1150);
or U3371 (N_3371,In_1220,In_1041);
nor U3372 (N_3372,In_59,In_1667);
nor U3373 (N_3373,In_166,In_9);
xnor U3374 (N_3374,In_1199,In_1714);
xnor U3375 (N_3375,In_2208,In_475);
or U3376 (N_3376,In_2174,In_950);
xnor U3377 (N_3377,In_1082,In_1437);
nor U3378 (N_3378,In_377,In_1026);
nand U3379 (N_3379,In_1436,In_2308);
or U3380 (N_3380,In_350,In_2091);
xor U3381 (N_3381,In_1106,In_717);
nor U3382 (N_3382,In_418,In_1361);
xor U3383 (N_3383,In_435,In_578);
or U3384 (N_3384,In_1125,In_1750);
and U3385 (N_3385,In_1249,In_2160);
and U3386 (N_3386,In_1058,In_813);
nand U3387 (N_3387,In_1686,In_2477);
xnor U3388 (N_3388,In_344,In_2043);
and U3389 (N_3389,In_716,In_284);
nor U3390 (N_3390,In_1305,In_1905);
and U3391 (N_3391,In_231,In_1358);
and U3392 (N_3392,In_358,In_2486);
or U3393 (N_3393,In_437,In_733);
xor U3394 (N_3394,In_1231,In_1726);
or U3395 (N_3395,In_260,In_816);
xnor U3396 (N_3396,In_675,In_2277);
and U3397 (N_3397,In_1872,In_152);
xnor U3398 (N_3398,In_1754,In_1149);
nand U3399 (N_3399,In_260,In_1668);
nand U3400 (N_3400,In_2473,In_2219);
or U3401 (N_3401,In_170,In_1996);
nor U3402 (N_3402,In_1938,In_733);
nor U3403 (N_3403,In_255,In_694);
nand U3404 (N_3404,In_83,In_1185);
and U3405 (N_3405,In_1016,In_835);
xnor U3406 (N_3406,In_2435,In_1325);
nand U3407 (N_3407,In_2080,In_103);
xnor U3408 (N_3408,In_59,In_2237);
nor U3409 (N_3409,In_2404,In_786);
nor U3410 (N_3410,In_1357,In_33);
nand U3411 (N_3411,In_610,In_260);
and U3412 (N_3412,In_2091,In_310);
nand U3413 (N_3413,In_1298,In_1314);
or U3414 (N_3414,In_1896,In_1069);
and U3415 (N_3415,In_2355,In_403);
or U3416 (N_3416,In_571,In_1554);
xnor U3417 (N_3417,In_1788,In_2309);
nor U3418 (N_3418,In_1169,In_1578);
and U3419 (N_3419,In_2030,In_1599);
nor U3420 (N_3420,In_44,In_1005);
nand U3421 (N_3421,In_700,In_288);
xnor U3422 (N_3422,In_825,In_1703);
and U3423 (N_3423,In_84,In_1268);
or U3424 (N_3424,In_2491,In_2059);
xnor U3425 (N_3425,In_860,In_1375);
and U3426 (N_3426,In_127,In_409);
xor U3427 (N_3427,In_2279,In_2318);
nand U3428 (N_3428,In_108,In_416);
or U3429 (N_3429,In_2002,In_2024);
xnor U3430 (N_3430,In_2122,In_1584);
or U3431 (N_3431,In_2112,In_1993);
or U3432 (N_3432,In_1522,In_875);
nor U3433 (N_3433,In_716,In_1384);
and U3434 (N_3434,In_526,In_1463);
nor U3435 (N_3435,In_1903,In_2223);
and U3436 (N_3436,In_1069,In_1892);
xnor U3437 (N_3437,In_2467,In_305);
nand U3438 (N_3438,In_1611,In_2154);
nor U3439 (N_3439,In_2407,In_1331);
xnor U3440 (N_3440,In_1870,In_839);
and U3441 (N_3441,In_486,In_1012);
xor U3442 (N_3442,In_2396,In_2301);
nand U3443 (N_3443,In_1975,In_2312);
or U3444 (N_3444,In_1310,In_1343);
nor U3445 (N_3445,In_619,In_464);
nand U3446 (N_3446,In_2422,In_1119);
nor U3447 (N_3447,In_1426,In_2314);
nand U3448 (N_3448,In_138,In_1063);
nor U3449 (N_3449,In_1804,In_1372);
or U3450 (N_3450,In_1198,In_1730);
and U3451 (N_3451,In_1749,In_2362);
nand U3452 (N_3452,In_335,In_2360);
nand U3453 (N_3453,In_2320,In_257);
nor U3454 (N_3454,In_1486,In_613);
nor U3455 (N_3455,In_2205,In_2327);
nor U3456 (N_3456,In_1312,In_1937);
nor U3457 (N_3457,In_385,In_596);
or U3458 (N_3458,In_2122,In_2493);
xnor U3459 (N_3459,In_590,In_2163);
xnor U3460 (N_3460,In_1640,In_357);
nand U3461 (N_3461,In_1396,In_131);
nor U3462 (N_3462,In_594,In_1590);
or U3463 (N_3463,In_1724,In_866);
and U3464 (N_3464,In_994,In_1882);
and U3465 (N_3465,In_68,In_506);
nor U3466 (N_3466,In_716,In_956);
or U3467 (N_3467,In_1290,In_2337);
and U3468 (N_3468,In_2298,In_1923);
nor U3469 (N_3469,In_2345,In_2070);
nor U3470 (N_3470,In_2277,In_476);
or U3471 (N_3471,In_2404,In_621);
nand U3472 (N_3472,In_400,In_1254);
nor U3473 (N_3473,In_2408,In_1519);
or U3474 (N_3474,In_774,In_972);
and U3475 (N_3475,In_1071,In_1346);
nand U3476 (N_3476,In_775,In_55);
and U3477 (N_3477,In_2079,In_2302);
nor U3478 (N_3478,In_1544,In_1616);
xor U3479 (N_3479,In_942,In_269);
xnor U3480 (N_3480,In_1320,In_318);
nand U3481 (N_3481,In_1888,In_694);
and U3482 (N_3482,In_944,In_503);
or U3483 (N_3483,In_221,In_17);
nand U3484 (N_3484,In_1550,In_2128);
and U3485 (N_3485,In_1165,In_1196);
or U3486 (N_3486,In_157,In_2320);
or U3487 (N_3487,In_1037,In_102);
and U3488 (N_3488,In_2247,In_810);
nand U3489 (N_3489,In_2179,In_324);
xnor U3490 (N_3490,In_375,In_1285);
xnor U3491 (N_3491,In_770,In_1007);
nor U3492 (N_3492,In_547,In_2417);
and U3493 (N_3493,In_1927,In_2010);
nor U3494 (N_3494,In_2179,In_1981);
nand U3495 (N_3495,In_49,In_617);
xnor U3496 (N_3496,In_1364,In_124);
nand U3497 (N_3497,In_1495,In_2237);
xor U3498 (N_3498,In_281,In_2094);
xor U3499 (N_3499,In_1340,In_274);
or U3500 (N_3500,In_1768,In_2075);
nor U3501 (N_3501,In_507,In_167);
or U3502 (N_3502,In_618,In_1154);
nand U3503 (N_3503,In_1247,In_1183);
and U3504 (N_3504,In_512,In_2465);
and U3505 (N_3505,In_2317,In_555);
nand U3506 (N_3506,In_1994,In_468);
and U3507 (N_3507,In_1600,In_1355);
or U3508 (N_3508,In_1769,In_398);
nand U3509 (N_3509,In_1195,In_88);
nand U3510 (N_3510,In_666,In_1088);
nor U3511 (N_3511,In_1020,In_1878);
xnor U3512 (N_3512,In_2104,In_936);
xor U3513 (N_3513,In_1861,In_1991);
or U3514 (N_3514,In_509,In_1524);
xor U3515 (N_3515,In_733,In_2055);
nor U3516 (N_3516,In_517,In_1958);
nor U3517 (N_3517,In_1202,In_2220);
or U3518 (N_3518,In_747,In_2105);
xor U3519 (N_3519,In_2013,In_2220);
nand U3520 (N_3520,In_925,In_2246);
nand U3521 (N_3521,In_19,In_1087);
or U3522 (N_3522,In_2375,In_1544);
nand U3523 (N_3523,In_1888,In_1859);
and U3524 (N_3524,In_258,In_2295);
nor U3525 (N_3525,In_405,In_581);
nand U3526 (N_3526,In_937,In_155);
and U3527 (N_3527,In_778,In_1451);
nand U3528 (N_3528,In_924,In_2216);
or U3529 (N_3529,In_1828,In_761);
and U3530 (N_3530,In_2191,In_372);
xnor U3531 (N_3531,In_1242,In_2178);
or U3532 (N_3532,In_1937,In_440);
and U3533 (N_3533,In_634,In_250);
nor U3534 (N_3534,In_1524,In_2089);
or U3535 (N_3535,In_1377,In_1463);
nor U3536 (N_3536,In_2358,In_1140);
and U3537 (N_3537,In_998,In_120);
xor U3538 (N_3538,In_1397,In_81);
nor U3539 (N_3539,In_1690,In_1057);
or U3540 (N_3540,In_545,In_1481);
xor U3541 (N_3541,In_1061,In_2367);
and U3542 (N_3542,In_997,In_590);
nor U3543 (N_3543,In_121,In_945);
xor U3544 (N_3544,In_13,In_417);
or U3545 (N_3545,In_1908,In_1369);
nor U3546 (N_3546,In_901,In_217);
xor U3547 (N_3547,In_22,In_321);
nand U3548 (N_3548,In_1348,In_1552);
nor U3549 (N_3549,In_2257,In_2425);
and U3550 (N_3550,In_1018,In_1092);
and U3551 (N_3551,In_491,In_1824);
or U3552 (N_3552,In_47,In_64);
nor U3553 (N_3553,In_834,In_2416);
nand U3554 (N_3554,In_437,In_709);
xor U3555 (N_3555,In_713,In_37);
nor U3556 (N_3556,In_1179,In_2354);
and U3557 (N_3557,In_1682,In_1328);
or U3558 (N_3558,In_1154,In_384);
nor U3559 (N_3559,In_1907,In_2057);
nor U3560 (N_3560,In_1086,In_500);
or U3561 (N_3561,In_1435,In_1768);
and U3562 (N_3562,In_1907,In_1825);
xor U3563 (N_3563,In_1883,In_281);
nor U3564 (N_3564,In_869,In_1205);
and U3565 (N_3565,In_664,In_1054);
nor U3566 (N_3566,In_2418,In_2433);
and U3567 (N_3567,In_1615,In_1256);
xnor U3568 (N_3568,In_113,In_1855);
xnor U3569 (N_3569,In_269,In_253);
or U3570 (N_3570,In_855,In_712);
nand U3571 (N_3571,In_2174,In_483);
or U3572 (N_3572,In_2495,In_2342);
nand U3573 (N_3573,In_1646,In_372);
nor U3574 (N_3574,In_450,In_57);
nor U3575 (N_3575,In_1642,In_1049);
nand U3576 (N_3576,In_2291,In_827);
and U3577 (N_3577,In_1294,In_1587);
nand U3578 (N_3578,In_2165,In_830);
and U3579 (N_3579,In_816,In_1322);
and U3580 (N_3580,In_2294,In_1421);
nor U3581 (N_3581,In_2429,In_1878);
and U3582 (N_3582,In_1684,In_2404);
and U3583 (N_3583,In_1218,In_790);
nor U3584 (N_3584,In_1412,In_2195);
or U3585 (N_3585,In_1413,In_2484);
nor U3586 (N_3586,In_1984,In_1893);
xnor U3587 (N_3587,In_1412,In_2212);
nor U3588 (N_3588,In_2294,In_1186);
and U3589 (N_3589,In_2376,In_2461);
nand U3590 (N_3590,In_1409,In_2039);
and U3591 (N_3591,In_1166,In_1652);
nand U3592 (N_3592,In_1293,In_2377);
nor U3593 (N_3593,In_934,In_247);
and U3594 (N_3594,In_1012,In_708);
nor U3595 (N_3595,In_2474,In_1999);
nand U3596 (N_3596,In_1555,In_1622);
nand U3597 (N_3597,In_577,In_2318);
nand U3598 (N_3598,In_1197,In_789);
or U3599 (N_3599,In_1557,In_655);
nor U3600 (N_3600,In_2076,In_1118);
and U3601 (N_3601,In_1385,In_2359);
xor U3602 (N_3602,In_701,In_145);
xor U3603 (N_3603,In_674,In_2329);
xor U3604 (N_3604,In_1523,In_2400);
or U3605 (N_3605,In_2475,In_2480);
nor U3606 (N_3606,In_32,In_864);
and U3607 (N_3607,In_1798,In_898);
nor U3608 (N_3608,In_1428,In_707);
nor U3609 (N_3609,In_2136,In_1298);
xor U3610 (N_3610,In_26,In_600);
nor U3611 (N_3611,In_810,In_2179);
nor U3612 (N_3612,In_2402,In_376);
and U3613 (N_3613,In_2271,In_1992);
nor U3614 (N_3614,In_545,In_2247);
and U3615 (N_3615,In_40,In_1526);
and U3616 (N_3616,In_2200,In_1320);
and U3617 (N_3617,In_211,In_616);
or U3618 (N_3618,In_1271,In_1768);
or U3619 (N_3619,In_1300,In_2221);
or U3620 (N_3620,In_1702,In_1416);
or U3621 (N_3621,In_744,In_20);
nor U3622 (N_3622,In_2013,In_1942);
and U3623 (N_3623,In_601,In_1727);
nor U3624 (N_3624,In_320,In_2415);
xnor U3625 (N_3625,In_79,In_1367);
xor U3626 (N_3626,In_1139,In_1828);
xnor U3627 (N_3627,In_1623,In_1433);
nor U3628 (N_3628,In_2053,In_2495);
nor U3629 (N_3629,In_2032,In_1515);
xor U3630 (N_3630,In_9,In_1709);
or U3631 (N_3631,In_891,In_866);
or U3632 (N_3632,In_498,In_627);
and U3633 (N_3633,In_953,In_1898);
or U3634 (N_3634,In_548,In_250);
nand U3635 (N_3635,In_1975,In_1001);
or U3636 (N_3636,In_709,In_2166);
and U3637 (N_3637,In_1089,In_1568);
and U3638 (N_3638,In_303,In_297);
xor U3639 (N_3639,In_1083,In_1924);
nand U3640 (N_3640,In_2399,In_2447);
and U3641 (N_3641,In_361,In_1850);
and U3642 (N_3642,In_2227,In_1266);
nor U3643 (N_3643,In_468,In_1537);
and U3644 (N_3644,In_165,In_1522);
nor U3645 (N_3645,In_1980,In_1480);
nor U3646 (N_3646,In_1291,In_147);
and U3647 (N_3647,In_1953,In_1370);
and U3648 (N_3648,In_135,In_1982);
nand U3649 (N_3649,In_272,In_149);
or U3650 (N_3650,In_1845,In_260);
or U3651 (N_3651,In_871,In_1192);
nand U3652 (N_3652,In_2284,In_1028);
nor U3653 (N_3653,In_263,In_2273);
or U3654 (N_3654,In_2101,In_2029);
or U3655 (N_3655,In_199,In_715);
nand U3656 (N_3656,In_2495,In_2324);
xor U3657 (N_3657,In_1697,In_2404);
nand U3658 (N_3658,In_1309,In_182);
or U3659 (N_3659,In_386,In_309);
nand U3660 (N_3660,In_113,In_856);
nand U3661 (N_3661,In_2296,In_307);
nor U3662 (N_3662,In_1258,In_681);
or U3663 (N_3663,In_1833,In_1976);
nor U3664 (N_3664,In_1373,In_2357);
or U3665 (N_3665,In_1083,In_2404);
and U3666 (N_3666,In_2171,In_1744);
and U3667 (N_3667,In_417,In_1577);
xor U3668 (N_3668,In_2205,In_647);
and U3669 (N_3669,In_2324,In_2176);
nand U3670 (N_3670,In_1158,In_568);
nand U3671 (N_3671,In_971,In_2267);
nand U3672 (N_3672,In_114,In_954);
or U3673 (N_3673,In_1227,In_176);
and U3674 (N_3674,In_1128,In_1896);
or U3675 (N_3675,In_1017,In_1111);
nand U3676 (N_3676,In_93,In_1194);
nand U3677 (N_3677,In_1307,In_903);
or U3678 (N_3678,In_1886,In_2227);
nand U3679 (N_3679,In_2329,In_528);
nor U3680 (N_3680,In_434,In_317);
and U3681 (N_3681,In_1358,In_441);
or U3682 (N_3682,In_2086,In_2266);
or U3683 (N_3683,In_2055,In_483);
nand U3684 (N_3684,In_1214,In_1639);
or U3685 (N_3685,In_2404,In_2131);
nand U3686 (N_3686,In_1099,In_2459);
nor U3687 (N_3687,In_2467,In_1897);
and U3688 (N_3688,In_2485,In_213);
xor U3689 (N_3689,In_233,In_56);
xor U3690 (N_3690,In_1792,In_70);
xnor U3691 (N_3691,In_1051,In_56);
and U3692 (N_3692,In_984,In_1166);
nand U3693 (N_3693,In_2499,In_1254);
and U3694 (N_3694,In_2344,In_191);
nand U3695 (N_3695,In_1432,In_2103);
and U3696 (N_3696,In_310,In_1038);
nor U3697 (N_3697,In_1003,In_1638);
or U3698 (N_3698,In_2243,In_1390);
nand U3699 (N_3699,In_1069,In_2472);
nand U3700 (N_3700,In_2383,In_1084);
nor U3701 (N_3701,In_1490,In_1765);
xnor U3702 (N_3702,In_743,In_575);
and U3703 (N_3703,In_263,In_1130);
nor U3704 (N_3704,In_1062,In_2362);
nor U3705 (N_3705,In_493,In_1225);
and U3706 (N_3706,In_1107,In_862);
nor U3707 (N_3707,In_492,In_935);
or U3708 (N_3708,In_988,In_2028);
nand U3709 (N_3709,In_1102,In_982);
nand U3710 (N_3710,In_1206,In_251);
nor U3711 (N_3711,In_1007,In_1585);
or U3712 (N_3712,In_1067,In_899);
nand U3713 (N_3713,In_51,In_1745);
nor U3714 (N_3714,In_1183,In_333);
and U3715 (N_3715,In_1985,In_2153);
or U3716 (N_3716,In_1812,In_1144);
nor U3717 (N_3717,In_1368,In_1061);
nor U3718 (N_3718,In_1947,In_309);
xor U3719 (N_3719,In_1892,In_2347);
xor U3720 (N_3720,In_324,In_821);
xor U3721 (N_3721,In_2492,In_1937);
nand U3722 (N_3722,In_351,In_621);
xnor U3723 (N_3723,In_908,In_37);
and U3724 (N_3724,In_2107,In_1681);
nor U3725 (N_3725,In_879,In_305);
or U3726 (N_3726,In_1578,In_892);
nor U3727 (N_3727,In_840,In_2338);
nor U3728 (N_3728,In_2289,In_2266);
nor U3729 (N_3729,In_1346,In_2053);
xnor U3730 (N_3730,In_1916,In_170);
and U3731 (N_3731,In_356,In_1692);
and U3732 (N_3732,In_1717,In_1460);
nand U3733 (N_3733,In_1575,In_1712);
nand U3734 (N_3734,In_765,In_2302);
and U3735 (N_3735,In_915,In_764);
and U3736 (N_3736,In_1739,In_2070);
nand U3737 (N_3737,In_2160,In_765);
and U3738 (N_3738,In_47,In_977);
nor U3739 (N_3739,In_1507,In_1993);
nand U3740 (N_3740,In_629,In_2350);
nand U3741 (N_3741,In_80,In_39);
or U3742 (N_3742,In_1721,In_634);
and U3743 (N_3743,In_2267,In_656);
or U3744 (N_3744,In_1144,In_410);
nor U3745 (N_3745,In_349,In_654);
or U3746 (N_3746,In_1317,In_1624);
nand U3747 (N_3747,In_2018,In_237);
and U3748 (N_3748,In_707,In_163);
or U3749 (N_3749,In_1659,In_2081);
nor U3750 (N_3750,In_261,In_346);
nand U3751 (N_3751,In_26,In_16);
xnor U3752 (N_3752,In_2074,In_1570);
and U3753 (N_3753,In_2074,In_945);
or U3754 (N_3754,In_69,In_1134);
and U3755 (N_3755,In_1678,In_1691);
and U3756 (N_3756,In_679,In_620);
xnor U3757 (N_3757,In_208,In_253);
nor U3758 (N_3758,In_1828,In_1349);
nor U3759 (N_3759,In_399,In_443);
xor U3760 (N_3760,In_1164,In_1429);
or U3761 (N_3761,In_644,In_2163);
xor U3762 (N_3762,In_661,In_1503);
or U3763 (N_3763,In_836,In_1711);
xor U3764 (N_3764,In_2430,In_262);
or U3765 (N_3765,In_1095,In_1993);
nor U3766 (N_3766,In_1569,In_1757);
xor U3767 (N_3767,In_1742,In_259);
xor U3768 (N_3768,In_509,In_1103);
and U3769 (N_3769,In_2481,In_233);
nor U3770 (N_3770,In_876,In_572);
and U3771 (N_3771,In_2188,In_969);
or U3772 (N_3772,In_445,In_1949);
nand U3773 (N_3773,In_313,In_820);
nand U3774 (N_3774,In_2254,In_2334);
or U3775 (N_3775,In_1149,In_2255);
or U3776 (N_3776,In_7,In_2119);
xnor U3777 (N_3777,In_736,In_491);
nand U3778 (N_3778,In_48,In_467);
xnor U3779 (N_3779,In_1639,In_246);
nor U3780 (N_3780,In_1525,In_1875);
nor U3781 (N_3781,In_2329,In_113);
xor U3782 (N_3782,In_2451,In_1710);
xnor U3783 (N_3783,In_1877,In_306);
xor U3784 (N_3784,In_2240,In_60);
xor U3785 (N_3785,In_1823,In_214);
nor U3786 (N_3786,In_1364,In_1388);
or U3787 (N_3787,In_1109,In_321);
nand U3788 (N_3788,In_1155,In_881);
xnor U3789 (N_3789,In_1416,In_29);
nor U3790 (N_3790,In_1987,In_20);
nor U3791 (N_3791,In_1202,In_1230);
or U3792 (N_3792,In_106,In_1019);
nor U3793 (N_3793,In_3,In_51);
and U3794 (N_3794,In_1600,In_177);
nor U3795 (N_3795,In_1480,In_971);
or U3796 (N_3796,In_1020,In_379);
xnor U3797 (N_3797,In_1050,In_2365);
xor U3798 (N_3798,In_212,In_1496);
xor U3799 (N_3799,In_2144,In_1192);
nand U3800 (N_3800,In_1392,In_1255);
xor U3801 (N_3801,In_2462,In_656);
xor U3802 (N_3802,In_490,In_2201);
or U3803 (N_3803,In_2086,In_913);
xnor U3804 (N_3804,In_748,In_1822);
xnor U3805 (N_3805,In_1863,In_2066);
or U3806 (N_3806,In_1470,In_1984);
nor U3807 (N_3807,In_1176,In_2211);
nand U3808 (N_3808,In_106,In_648);
xor U3809 (N_3809,In_944,In_830);
and U3810 (N_3810,In_1000,In_882);
nand U3811 (N_3811,In_224,In_697);
xor U3812 (N_3812,In_1819,In_1267);
nor U3813 (N_3813,In_1918,In_637);
and U3814 (N_3814,In_85,In_650);
nand U3815 (N_3815,In_2233,In_1988);
xnor U3816 (N_3816,In_976,In_1136);
nand U3817 (N_3817,In_2158,In_1577);
and U3818 (N_3818,In_1051,In_24);
xnor U3819 (N_3819,In_105,In_1472);
nor U3820 (N_3820,In_1594,In_1704);
nor U3821 (N_3821,In_2298,In_2473);
nand U3822 (N_3822,In_185,In_1622);
or U3823 (N_3823,In_277,In_691);
or U3824 (N_3824,In_457,In_1617);
nand U3825 (N_3825,In_2133,In_235);
nand U3826 (N_3826,In_2105,In_1739);
or U3827 (N_3827,In_906,In_1866);
or U3828 (N_3828,In_1958,In_1634);
or U3829 (N_3829,In_601,In_2123);
xor U3830 (N_3830,In_2391,In_1379);
or U3831 (N_3831,In_1742,In_1510);
or U3832 (N_3832,In_1191,In_1214);
nand U3833 (N_3833,In_828,In_352);
or U3834 (N_3834,In_566,In_1324);
nand U3835 (N_3835,In_394,In_626);
nor U3836 (N_3836,In_1393,In_157);
nand U3837 (N_3837,In_2441,In_625);
nand U3838 (N_3838,In_1942,In_1955);
xor U3839 (N_3839,In_1399,In_1538);
or U3840 (N_3840,In_945,In_1539);
nor U3841 (N_3841,In_1625,In_1941);
nand U3842 (N_3842,In_1143,In_2480);
nor U3843 (N_3843,In_2110,In_10);
nand U3844 (N_3844,In_1893,In_2413);
nor U3845 (N_3845,In_1380,In_233);
nor U3846 (N_3846,In_1726,In_1119);
nor U3847 (N_3847,In_1820,In_2159);
and U3848 (N_3848,In_1828,In_1511);
and U3849 (N_3849,In_1657,In_754);
and U3850 (N_3850,In_378,In_454);
or U3851 (N_3851,In_506,In_2215);
xor U3852 (N_3852,In_2040,In_1191);
nor U3853 (N_3853,In_1488,In_996);
xor U3854 (N_3854,In_1744,In_1511);
nor U3855 (N_3855,In_2061,In_2375);
nand U3856 (N_3856,In_2385,In_387);
and U3857 (N_3857,In_278,In_63);
nor U3858 (N_3858,In_336,In_2216);
and U3859 (N_3859,In_2146,In_1739);
nand U3860 (N_3860,In_1457,In_112);
nor U3861 (N_3861,In_258,In_2307);
nand U3862 (N_3862,In_617,In_146);
or U3863 (N_3863,In_2193,In_1336);
xor U3864 (N_3864,In_1589,In_366);
and U3865 (N_3865,In_1225,In_761);
nand U3866 (N_3866,In_888,In_545);
nor U3867 (N_3867,In_902,In_121);
xor U3868 (N_3868,In_1784,In_1150);
or U3869 (N_3869,In_776,In_625);
or U3870 (N_3870,In_1298,In_943);
nand U3871 (N_3871,In_2238,In_1918);
xor U3872 (N_3872,In_1630,In_172);
xor U3873 (N_3873,In_2088,In_2236);
or U3874 (N_3874,In_1694,In_682);
xnor U3875 (N_3875,In_1245,In_1563);
nor U3876 (N_3876,In_1038,In_2434);
or U3877 (N_3877,In_1615,In_1321);
or U3878 (N_3878,In_1147,In_2260);
xor U3879 (N_3879,In_1150,In_2357);
nor U3880 (N_3880,In_98,In_2491);
nand U3881 (N_3881,In_582,In_2307);
nand U3882 (N_3882,In_1835,In_1548);
or U3883 (N_3883,In_1465,In_381);
xor U3884 (N_3884,In_876,In_1631);
or U3885 (N_3885,In_1657,In_960);
nand U3886 (N_3886,In_2472,In_2004);
and U3887 (N_3887,In_1938,In_1493);
nor U3888 (N_3888,In_556,In_2118);
nor U3889 (N_3889,In_2088,In_1637);
or U3890 (N_3890,In_1950,In_1821);
nand U3891 (N_3891,In_323,In_1399);
xor U3892 (N_3892,In_1775,In_1400);
xor U3893 (N_3893,In_1327,In_2438);
xnor U3894 (N_3894,In_442,In_1459);
and U3895 (N_3895,In_1955,In_1330);
nor U3896 (N_3896,In_2320,In_2244);
nor U3897 (N_3897,In_1898,In_88);
nand U3898 (N_3898,In_1127,In_1199);
or U3899 (N_3899,In_2456,In_808);
nand U3900 (N_3900,In_197,In_999);
or U3901 (N_3901,In_2309,In_517);
and U3902 (N_3902,In_479,In_1350);
nor U3903 (N_3903,In_134,In_2284);
or U3904 (N_3904,In_1589,In_957);
or U3905 (N_3905,In_39,In_778);
and U3906 (N_3906,In_1104,In_287);
nand U3907 (N_3907,In_92,In_611);
or U3908 (N_3908,In_988,In_963);
nor U3909 (N_3909,In_1365,In_1983);
nor U3910 (N_3910,In_1197,In_463);
xnor U3911 (N_3911,In_1271,In_1755);
xnor U3912 (N_3912,In_1334,In_388);
nand U3913 (N_3913,In_2136,In_1160);
nor U3914 (N_3914,In_826,In_1909);
or U3915 (N_3915,In_669,In_683);
xor U3916 (N_3916,In_925,In_616);
nand U3917 (N_3917,In_2256,In_45);
and U3918 (N_3918,In_1337,In_1682);
xor U3919 (N_3919,In_8,In_1755);
nand U3920 (N_3920,In_1534,In_996);
or U3921 (N_3921,In_1278,In_952);
nor U3922 (N_3922,In_1255,In_2197);
nor U3923 (N_3923,In_795,In_1629);
nand U3924 (N_3924,In_172,In_295);
xor U3925 (N_3925,In_1145,In_702);
nor U3926 (N_3926,In_1028,In_2268);
nor U3927 (N_3927,In_951,In_1603);
xnor U3928 (N_3928,In_1928,In_574);
and U3929 (N_3929,In_1882,In_1484);
nand U3930 (N_3930,In_1606,In_530);
nand U3931 (N_3931,In_1096,In_359);
and U3932 (N_3932,In_57,In_1527);
nand U3933 (N_3933,In_2104,In_242);
and U3934 (N_3934,In_1757,In_905);
nor U3935 (N_3935,In_387,In_504);
xnor U3936 (N_3936,In_1371,In_1512);
or U3937 (N_3937,In_1983,In_247);
and U3938 (N_3938,In_1975,In_100);
nor U3939 (N_3939,In_798,In_917);
xnor U3940 (N_3940,In_321,In_2377);
nand U3941 (N_3941,In_628,In_1659);
nor U3942 (N_3942,In_1465,In_2344);
nand U3943 (N_3943,In_534,In_99);
and U3944 (N_3944,In_1348,In_1620);
and U3945 (N_3945,In_869,In_2455);
or U3946 (N_3946,In_1057,In_1126);
or U3947 (N_3947,In_91,In_842);
nand U3948 (N_3948,In_1195,In_1988);
nand U3949 (N_3949,In_1209,In_1771);
nor U3950 (N_3950,In_2295,In_1887);
or U3951 (N_3951,In_129,In_977);
xnor U3952 (N_3952,In_1357,In_2165);
or U3953 (N_3953,In_308,In_2410);
and U3954 (N_3954,In_486,In_2292);
nand U3955 (N_3955,In_252,In_2348);
nand U3956 (N_3956,In_1467,In_2175);
and U3957 (N_3957,In_2426,In_2101);
nand U3958 (N_3958,In_2380,In_882);
nand U3959 (N_3959,In_988,In_2075);
nand U3960 (N_3960,In_349,In_1896);
and U3961 (N_3961,In_1533,In_2292);
nor U3962 (N_3962,In_1791,In_938);
and U3963 (N_3963,In_1474,In_1251);
xor U3964 (N_3964,In_1737,In_2165);
or U3965 (N_3965,In_1030,In_407);
xor U3966 (N_3966,In_1574,In_1524);
and U3967 (N_3967,In_1093,In_2148);
and U3968 (N_3968,In_1186,In_686);
or U3969 (N_3969,In_1680,In_2188);
nand U3970 (N_3970,In_382,In_1434);
nand U3971 (N_3971,In_1712,In_756);
nor U3972 (N_3972,In_1376,In_1270);
and U3973 (N_3973,In_192,In_2159);
nor U3974 (N_3974,In_489,In_2333);
and U3975 (N_3975,In_1239,In_534);
xnor U3976 (N_3976,In_5,In_401);
and U3977 (N_3977,In_2011,In_1458);
nor U3978 (N_3978,In_747,In_1902);
or U3979 (N_3979,In_1255,In_766);
nor U3980 (N_3980,In_2119,In_228);
or U3981 (N_3981,In_2020,In_1900);
nand U3982 (N_3982,In_774,In_848);
and U3983 (N_3983,In_1416,In_325);
nor U3984 (N_3984,In_714,In_1885);
xor U3985 (N_3985,In_1985,In_1554);
and U3986 (N_3986,In_1680,In_2199);
nor U3987 (N_3987,In_936,In_336);
xor U3988 (N_3988,In_1638,In_1250);
and U3989 (N_3989,In_1337,In_443);
xnor U3990 (N_3990,In_265,In_1253);
xor U3991 (N_3991,In_1383,In_797);
nor U3992 (N_3992,In_2366,In_818);
or U3993 (N_3993,In_1984,In_1628);
nand U3994 (N_3994,In_1286,In_2020);
xor U3995 (N_3995,In_962,In_304);
nand U3996 (N_3996,In_477,In_923);
nand U3997 (N_3997,In_2033,In_1623);
nand U3998 (N_3998,In_403,In_198);
or U3999 (N_3999,In_212,In_507);
and U4000 (N_4000,In_2013,In_2487);
nor U4001 (N_4001,In_2324,In_1735);
nor U4002 (N_4002,In_553,In_847);
and U4003 (N_4003,In_116,In_468);
nand U4004 (N_4004,In_371,In_1863);
and U4005 (N_4005,In_2414,In_2271);
and U4006 (N_4006,In_664,In_2386);
or U4007 (N_4007,In_1412,In_2312);
xor U4008 (N_4008,In_729,In_616);
nor U4009 (N_4009,In_616,In_855);
and U4010 (N_4010,In_1623,In_560);
nor U4011 (N_4011,In_628,In_2483);
nand U4012 (N_4012,In_2249,In_1101);
and U4013 (N_4013,In_1729,In_1860);
nor U4014 (N_4014,In_1269,In_35);
nand U4015 (N_4015,In_1087,In_47);
xor U4016 (N_4016,In_1869,In_1321);
nand U4017 (N_4017,In_661,In_848);
xor U4018 (N_4018,In_1687,In_878);
and U4019 (N_4019,In_1801,In_398);
or U4020 (N_4020,In_1885,In_2202);
xor U4021 (N_4021,In_2431,In_15);
nor U4022 (N_4022,In_1351,In_1474);
nand U4023 (N_4023,In_1799,In_2435);
nand U4024 (N_4024,In_2195,In_1639);
xnor U4025 (N_4025,In_213,In_1719);
xor U4026 (N_4026,In_99,In_139);
or U4027 (N_4027,In_739,In_345);
xnor U4028 (N_4028,In_2473,In_1172);
nor U4029 (N_4029,In_2152,In_1807);
and U4030 (N_4030,In_944,In_2447);
nand U4031 (N_4031,In_2113,In_116);
nand U4032 (N_4032,In_1304,In_468);
xnor U4033 (N_4033,In_1358,In_2312);
nor U4034 (N_4034,In_309,In_1688);
or U4035 (N_4035,In_1143,In_498);
xor U4036 (N_4036,In_889,In_2056);
nand U4037 (N_4037,In_1665,In_1784);
nor U4038 (N_4038,In_597,In_2054);
and U4039 (N_4039,In_1014,In_1463);
nor U4040 (N_4040,In_405,In_2417);
nor U4041 (N_4041,In_489,In_1748);
and U4042 (N_4042,In_1820,In_2066);
nand U4043 (N_4043,In_150,In_2285);
xor U4044 (N_4044,In_1937,In_1386);
and U4045 (N_4045,In_2400,In_322);
or U4046 (N_4046,In_684,In_1714);
nor U4047 (N_4047,In_2020,In_1185);
nand U4048 (N_4048,In_457,In_429);
xnor U4049 (N_4049,In_1215,In_1500);
and U4050 (N_4050,In_774,In_637);
or U4051 (N_4051,In_181,In_1780);
or U4052 (N_4052,In_453,In_1917);
nand U4053 (N_4053,In_354,In_497);
or U4054 (N_4054,In_1101,In_2080);
xnor U4055 (N_4055,In_1589,In_446);
or U4056 (N_4056,In_633,In_1321);
and U4057 (N_4057,In_186,In_698);
nor U4058 (N_4058,In_1772,In_2170);
nand U4059 (N_4059,In_2471,In_2108);
or U4060 (N_4060,In_1737,In_2390);
nor U4061 (N_4061,In_703,In_1735);
xnor U4062 (N_4062,In_2031,In_1452);
nor U4063 (N_4063,In_1804,In_335);
xnor U4064 (N_4064,In_1678,In_1940);
nor U4065 (N_4065,In_633,In_679);
nor U4066 (N_4066,In_2276,In_1675);
nand U4067 (N_4067,In_1625,In_572);
or U4068 (N_4068,In_2072,In_829);
xor U4069 (N_4069,In_183,In_1640);
nand U4070 (N_4070,In_629,In_2444);
xnor U4071 (N_4071,In_1326,In_1878);
xnor U4072 (N_4072,In_613,In_871);
and U4073 (N_4073,In_1822,In_99);
and U4074 (N_4074,In_678,In_765);
nor U4075 (N_4075,In_1230,In_2224);
nand U4076 (N_4076,In_1168,In_704);
nor U4077 (N_4077,In_454,In_1094);
nand U4078 (N_4078,In_1485,In_359);
and U4079 (N_4079,In_1161,In_2264);
or U4080 (N_4080,In_1411,In_2476);
xor U4081 (N_4081,In_2488,In_2372);
or U4082 (N_4082,In_1275,In_1273);
nand U4083 (N_4083,In_1344,In_1560);
nor U4084 (N_4084,In_1432,In_1372);
nand U4085 (N_4085,In_804,In_936);
nand U4086 (N_4086,In_2459,In_1719);
nor U4087 (N_4087,In_752,In_1498);
nor U4088 (N_4088,In_1639,In_854);
and U4089 (N_4089,In_1319,In_348);
nor U4090 (N_4090,In_1434,In_1587);
or U4091 (N_4091,In_835,In_324);
xor U4092 (N_4092,In_1229,In_1728);
nor U4093 (N_4093,In_615,In_597);
nor U4094 (N_4094,In_1442,In_2137);
nand U4095 (N_4095,In_274,In_411);
xnor U4096 (N_4096,In_2408,In_610);
and U4097 (N_4097,In_755,In_811);
nor U4098 (N_4098,In_304,In_1664);
nor U4099 (N_4099,In_1127,In_2338);
or U4100 (N_4100,In_1570,In_1915);
nor U4101 (N_4101,In_1006,In_869);
nor U4102 (N_4102,In_896,In_2311);
nor U4103 (N_4103,In_1545,In_586);
xor U4104 (N_4104,In_22,In_1619);
and U4105 (N_4105,In_1501,In_2199);
nor U4106 (N_4106,In_17,In_874);
nor U4107 (N_4107,In_841,In_1117);
xnor U4108 (N_4108,In_1140,In_73);
and U4109 (N_4109,In_1811,In_93);
xnor U4110 (N_4110,In_1511,In_770);
or U4111 (N_4111,In_380,In_300);
or U4112 (N_4112,In_54,In_388);
nor U4113 (N_4113,In_346,In_386);
or U4114 (N_4114,In_1311,In_702);
xnor U4115 (N_4115,In_1788,In_1204);
or U4116 (N_4116,In_1628,In_198);
xnor U4117 (N_4117,In_1706,In_2249);
nand U4118 (N_4118,In_891,In_1238);
nor U4119 (N_4119,In_1035,In_2323);
nand U4120 (N_4120,In_1346,In_1306);
nor U4121 (N_4121,In_289,In_2469);
xor U4122 (N_4122,In_2405,In_15);
xnor U4123 (N_4123,In_196,In_1051);
nor U4124 (N_4124,In_1969,In_1505);
or U4125 (N_4125,In_388,In_1058);
and U4126 (N_4126,In_1017,In_1543);
and U4127 (N_4127,In_713,In_777);
and U4128 (N_4128,In_1311,In_447);
and U4129 (N_4129,In_933,In_1945);
or U4130 (N_4130,In_1836,In_535);
and U4131 (N_4131,In_855,In_347);
nor U4132 (N_4132,In_1955,In_275);
and U4133 (N_4133,In_2407,In_1732);
or U4134 (N_4134,In_914,In_1455);
or U4135 (N_4135,In_945,In_1954);
nor U4136 (N_4136,In_2289,In_554);
xor U4137 (N_4137,In_348,In_2205);
nor U4138 (N_4138,In_1920,In_1038);
nor U4139 (N_4139,In_2214,In_463);
and U4140 (N_4140,In_737,In_1908);
or U4141 (N_4141,In_783,In_1163);
and U4142 (N_4142,In_1781,In_861);
xor U4143 (N_4143,In_1387,In_1498);
and U4144 (N_4144,In_2375,In_1419);
and U4145 (N_4145,In_2476,In_195);
or U4146 (N_4146,In_564,In_2484);
and U4147 (N_4147,In_769,In_1700);
xnor U4148 (N_4148,In_1230,In_1120);
xor U4149 (N_4149,In_1521,In_1511);
nor U4150 (N_4150,In_94,In_1948);
nor U4151 (N_4151,In_986,In_333);
nor U4152 (N_4152,In_2317,In_23);
nand U4153 (N_4153,In_1667,In_1668);
nand U4154 (N_4154,In_1504,In_2136);
and U4155 (N_4155,In_2209,In_837);
nand U4156 (N_4156,In_1183,In_2150);
and U4157 (N_4157,In_576,In_2156);
xor U4158 (N_4158,In_1039,In_2164);
nand U4159 (N_4159,In_1709,In_1834);
nor U4160 (N_4160,In_792,In_1701);
or U4161 (N_4161,In_750,In_947);
xor U4162 (N_4162,In_1011,In_2378);
xnor U4163 (N_4163,In_1132,In_1013);
or U4164 (N_4164,In_1011,In_570);
and U4165 (N_4165,In_2104,In_2220);
nor U4166 (N_4166,In_1088,In_1723);
nor U4167 (N_4167,In_832,In_2232);
nand U4168 (N_4168,In_934,In_83);
nor U4169 (N_4169,In_2072,In_929);
nor U4170 (N_4170,In_1032,In_1642);
xor U4171 (N_4171,In_2263,In_1989);
and U4172 (N_4172,In_1042,In_318);
xnor U4173 (N_4173,In_710,In_130);
or U4174 (N_4174,In_2333,In_1795);
nor U4175 (N_4175,In_724,In_1421);
xnor U4176 (N_4176,In_2467,In_376);
and U4177 (N_4177,In_1440,In_1445);
or U4178 (N_4178,In_397,In_1138);
xnor U4179 (N_4179,In_1723,In_48);
or U4180 (N_4180,In_2375,In_1800);
nor U4181 (N_4181,In_2046,In_1518);
xnor U4182 (N_4182,In_78,In_74);
xnor U4183 (N_4183,In_1148,In_1252);
xnor U4184 (N_4184,In_1480,In_1734);
nor U4185 (N_4185,In_2048,In_800);
nor U4186 (N_4186,In_1992,In_1563);
and U4187 (N_4187,In_1829,In_1771);
nand U4188 (N_4188,In_183,In_1233);
nand U4189 (N_4189,In_582,In_1966);
nor U4190 (N_4190,In_906,In_306);
nor U4191 (N_4191,In_26,In_503);
and U4192 (N_4192,In_1386,In_1495);
nor U4193 (N_4193,In_981,In_660);
nand U4194 (N_4194,In_917,In_1932);
or U4195 (N_4195,In_486,In_1052);
nand U4196 (N_4196,In_300,In_1775);
xor U4197 (N_4197,In_2341,In_2307);
xor U4198 (N_4198,In_152,In_2125);
xor U4199 (N_4199,In_1594,In_271);
or U4200 (N_4200,In_157,In_577);
nand U4201 (N_4201,In_2065,In_198);
nand U4202 (N_4202,In_909,In_414);
nand U4203 (N_4203,In_12,In_2067);
nand U4204 (N_4204,In_480,In_2346);
xnor U4205 (N_4205,In_1101,In_1685);
nor U4206 (N_4206,In_1968,In_505);
nand U4207 (N_4207,In_2312,In_1110);
nand U4208 (N_4208,In_1839,In_713);
nor U4209 (N_4209,In_1752,In_1239);
xnor U4210 (N_4210,In_2380,In_1559);
and U4211 (N_4211,In_1419,In_1542);
or U4212 (N_4212,In_1419,In_1657);
and U4213 (N_4213,In_1112,In_108);
and U4214 (N_4214,In_1014,In_816);
and U4215 (N_4215,In_1923,In_2479);
or U4216 (N_4216,In_2078,In_154);
xor U4217 (N_4217,In_122,In_2129);
xnor U4218 (N_4218,In_1590,In_280);
or U4219 (N_4219,In_471,In_661);
nand U4220 (N_4220,In_31,In_1891);
nand U4221 (N_4221,In_1071,In_649);
nand U4222 (N_4222,In_1582,In_1308);
xor U4223 (N_4223,In_2107,In_832);
or U4224 (N_4224,In_2292,In_2038);
nand U4225 (N_4225,In_1111,In_1173);
or U4226 (N_4226,In_2454,In_1725);
xnor U4227 (N_4227,In_1596,In_928);
xnor U4228 (N_4228,In_1828,In_55);
or U4229 (N_4229,In_451,In_414);
xnor U4230 (N_4230,In_901,In_983);
or U4231 (N_4231,In_1076,In_1959);
nor U4232 (N_4232,In_103,In_346);
nor U4233 (N_4233,In_1995,In_368);
or U4234 (N_4234,In_1491,In_125);
xor U4235 (N_4235,In_2407,In_870);
or U4236 (N_4236,In_2125,In_2448);
nand U4237 (N_4237,In_922,In_1636);
nor U4238 (N_4238,In_1095,In_535);
and U4239 (N_4239,In_2237,In_1324);
xor U4240 (N_4240,In_1757,In_963);
xnor U4241 (N_4241,In_78,In_2486);
and U4242 (N_4242,In_257,In_1731);
nand U4243 (N_4243,In_1820,In_2047);
xor U4244 (N_4244,In_2131,In_1619);
xor U4245 (N_4245,In_1982,In_324);
and U4246 (N_4246,In_410,In_66);
nand U4247 (N_4247,In_370,In_2240);
and U4248 (N_4248,In_1860,In_847);
nor U4249 (N_4249,In_1710,In_830);
and U4250 (N_4250,In_2002,In_2247);
and U4251 (N_4251,In_1477,In_543);
xnor U4252 (N_4252,In_1196,In_819);
nor U4253 (N_4253,In_737,In_1630);
and U4254 (N_4254,In_1153,In_1061);
and U4255 (N_4255,In_1950,In_1704);
and U4256 (N_4256,In_1805,In_1061);
and U4257 (N_4257,In_1328,In_341);
nand U4258 (N_4258,In_1241,In_1513);
nor U4259 (N_4259,In_1236,In_500);
nand U4260 (N_4260,In_1719,In_2118);
or U4261 (N_4261,In_688,In_834);
and U4262 (N_4262,In_499,In_2071);
nor U4263 (N_4263,In_2098,In_774);
nor U4264 (N_4264,In_862,In_817);
nor U4265 (N_4265,In_2123,In_1574);
nor U4266 (N_4266,In_541,In_864);
or U4267 (N_4267,In_375,In_613);
xor U4268 (N_4268,In_149,In_1826);
or U4269 (N_4269,In_515,In_1551);
xnor U4270 (N_4270,In_1361,In_1329);
or U4271 (N_4271,In_657,In_651);
xnor U4272 (N_4272,In_1598,In_1769);
nand U4273 (N_4273,In_1155,In_1292);
nand U4274 (N_4274,In_858,In_116);
or U4275 (N_4275,In_405,In_2368);
nand U4276 (N_4276,In_200,In_1318);
or U4277 (N_4277,In_1978,In_178);
nand U4278 (N_4278,In_2205,In_1741);
and U4279 (N_4279,In_823,In_218);
nor U4280 (N_4280,In_275,In_2484);
nand U4281 (N_4281,In_883,In_1089);
or U4282 (N_4282,In_1119,In_1168);
nor U4283 (N_4283,In_1000,In_1675);
xor U4284 (N_4284,In_2073,In_624);
or U4285 (N_4285,In_821,In_1144);
nor U4286 (N_4286,In_354,In_2231);
and U4287 (N_4287,In_650,In_1459);
and U4288 (N_4288,In_637,In_1103);
xnor U4289 (N_4289,In_2295,In_1279);
nor U4290 (N_4290,In_1331,In_155);
nor U4291 (N_4291,In_1105,In_582);
xnor U4292 (N_4292,In_2110,In_965);
nand U4293 (N_4293,In_171,In_1875);
or U4294 (N_4294,In_2208,In_548);
and U4295 (N_4295,In_1773,In_1716);
and U4296 (N_4296,In_1577,In_2013);
or U4297 (N_4297,In_582,In_2321);
nor U4298 (N_4298,In_419,In_337);
nor U4299 (N_4299,In_1620,In_366);
or U4300 (N_4300,In_2322,In_1416);
and U4301 (N_4301,In_914,In_760);
or U4302 (N_4302,In_1417,In_2417);
nand U4303 (N_4303,In_445,In_195);
or U4304 (N_4304,In_1374,In_1060);
nand U4305 (N_4305,In_112,In_76);
or U4306 (N_4306,In_2075,In_363);
xor U4307 (N_4307,In_2268,In_203);
and U4308 (N_4308,In_573,In_2153);
or U4309 (N_4309,In_1324,In_1712);
nand U4310 (N_4310,In_1838,In_1029);
nand U4311 (N_4311,In_1533,In_1732);
xnor U4312 (N_4312,In_2395,In_1479);
nor U4313 (N_4313,In_2305,In_230);
nor U4314 (N_4314,In_2158,In_534);
nor U4315 (N_4315,In_464,In_693);
nor U4316 (N_4316,In_362,In_244);
xnor U4317 (N_4317,In_1068,In_2010);
xnor U4318 (N_4318,In_2241,In_1765);
xor U4319 (N_4319,In_1181,In_1189);
and U4320 (N_4320,In_338,In_2149);
and U4321 (N_4321,In_2184,In_932);
nor U4322 (N_4322,In_1418,In_732);
nor U4323 (N_4323,In_705,In_798);
xor U4324 (N_4324,In_1047,In_1027);
and U4325 (N_4325,In_2434,In_1212);
xnor U4326 (N_4326,In_1056,In_2365);
nor U4327 (N_4327,In_1482,In_1336);
nand U4328 (N_4328,In_1275,In_1987);
and U4329 (N_4329,In_2050,In_790);
or U4330 (N_4330,In_614,In_407);
nand U4331 (N_4331,In_1097,In_2164);
and U4332 (N_4332,In_1129,In_1305);
xor U4333 (N_4333,In_645,In_1398);
nand U4334 (N_4334,In_1545,In_1734);
or U4335 (N_4335,In_989,In_2157);
and U4336 (N_4336,In_1216,In_2462);
or U4337 (N_4337,In_1590,In_1571);
and U4338 (N_4338,In_2041,In_814);
or U4339 (N_4339,In_140,In_1694);
nor U4340 (N_4340,In_554,In_2261);
nor U4341 (N_4341,In_73,In_939);
or U4342 (N_4342,In_747,In_1081);
xnor U4343 (N_4343,In_2047,In_1180);
or U4344 (N_4344,In_1091,In_112);
and U4345 (N_4345,In_1216,In_1590);
nor U4346 (N_4346,In_815,In_1187);
nor U4347 (N_4347,In_1930,In_1373);
nand U4348 (N_4348,In_1559,In_1440);
or U4349 (N_4349,In_237,In_2271);
xor U4350 (N_4350,In_707,In_1577);
and U4351 (N_4351,In_1845,In_258);
and U4352 (N_4352,In_1689,In_601);
nor U4353 (N_4353,In_1951,In_114);
xnor U4354 (N_4354,In_1439,In_1242);
nand U4355 (N_4355,In_2361,In_595);
or U4356 (N_4356,In_1668,In_312);
nor U4357 (N_4357,In_1875,In_888);
or U4358 (N_4358,In_1317,In_2454);
nor U4359 (N_4359,In_376,In_1674);
nand U4360 (N_4360,In_1305,In_1684);
xnor U4361 (N_4361,In_2185,In_2346);
nand U4362 (N_4362,In_282,In_705);
or U4363 (N_4363,In_1439,In_1873);
and U4364 (N_4364,In_2319,In_838);
nor U4365 (N_4365,In_346,In_1247);
and U4366 (N_4366,In_1904,In_1540);
nand U4367 (N_4367,In_1789,In_2463);
or U4368 (N_4368,In_1494,In_1594);
xor U4369 (N_4369,In_1067,In_1517);
xnor U4370 (N_4370,In_1385,In_1326);
nor U4371 (N_4371,In_2443,In_266);
nor U4372 (N_4372,In_1170,In_493);
nand U4373 (N_4373,In_1027,In_1414);
nor U4374 (N_4374,In_600,In_519);
and U4375 (N_4375,In_741,In_2484);
nor U4376 (N_4376,In_440,In_551);
nand U4377 (N_4377,In_2107,In_1307);
nor U4378 (N_4378,In_733,In_544);
nand U4379 (N_4379,In_1968,In_1564);
xor U4380 (N_4380,In_1931,In_914);
xor U4381 (N_4381,In_122,In_728);
xnor U4382 (N_4382,In_658,In_1409);
nand U4383 (N_4383,In_416,In_51);
or U4384 (N_4384,In_1944,In_1472);
nand U4385 (N_4385,In_1435,In_568);
or U4386 (N_4386,In_130,In_1162);
nor U4387 (N_4387,In_1045,In_836);
or U4388 (N_4388,In_2386,In_922);
and U4389 (N_4389,In_1663,In_322);
xor U4390 (N_4390,In_1882,In_184);
xor U4391 (N_4391,In_520,In_2020);
nand U4392 (N_4392,In_747,In_1340);
or U4393 (N_4393,In_1184,In_2183);
or U4394 (N_4394,In_477,In_1581);
and U4395 (N_4395,In_607,In_369);
xor U4396 (N_4396,In_374,In_2296);
xor U4397 (N_4397,In_2186,In_745);
or U4398 (N_4398,In_2404,In_278);
and U4399 (N_4399,In_721,In_626);
nand U4400 (N_4400,In_34,In_1997);
nand U4401 (N_4401,In_1819,In_1031);
or U4402 (N_4402,In_164,In_1260);
nor U4403 (N_4403,In_853,In_1412);
nand U4404 (N_4404,In_1898,In_482);
nand U4405 (N_4405,In_2371,In_1459);
and U4406 (N_4406,In_226,In_301);
or U4407 (N_4407,In_1850,In_1164);
nor U4408 (N_4408,In_115,In_1999);
xnor U4409 (N_4409,In_644,In_2106);
or U4410 (N_4410,In_147,In_80);
nor U4411 (N_4411,In_2493,In_1618);
nand U4412 (N_4412,In_516,In_248);
xor U4413 (N_4413,In_2456,In_1238);
xnor U4414 (N_4414,In_390,In_861);
or U4415 (N_4415,In_2361,In_1679);
xnor U4416 (N_4416,In_7,In_210);
nor U4417 (N_4417,In_2271,In_17);
nor U4418 (N_4418,In_2435,In_873);
xor U4419 (N_4419,In_191,In_1490);
nand U4420 (N_4420,In_786,In_460);
or U4421 (N_4421,In_374,In_1071);
and U4422 (N_4422,In_2212,In_1231);
or U4423 (N_4423,In_1189,In_1226);
nand U4424 (N_4424,In_1251,In_1794);
nor U4425 (N_4425,In_1750,In_48);
nand U4426 (N_4426,In_633,In_2059);
and U4427 (N_4427,In_408,In_2238);
and U4428 (N_4428,In_1171,In_1076);
nor U4429 (N_4429,In_425,In_2102);
xor U4430 (N_4430,In_777,In_1026);
or U4431 (N_4431,In_2423,In_981);
nand U4432 (N_4432,In_693,In_2059);
nand U4433 (N_4433,In_2316,In_306);
nand U4434 (N_4434,In_858,In_10);
and U4435 (N_4435,In_2424,In_1700);
xnor U4436 (N_4436,In_2085,In_1177);
nor U4437 (N_4437,In_449,In_890);
xnor U4438 (N_4438,In_673,In_657);
or U4439 (N_4439,In_171,In_1186);
nor U4440 (N_4440,In_1163,In_1594);
xor U4441 (N_4441,In_2312,In_22);
xnor U4442 (N_4442,In_1344,In_965);
xnor U4443 (N_4443,In_2426,In_1252);
nor U4444 (N_4444,In_573,In_1643);
xnor U4445 (N_4445,In_1083,In_452);
nor U4446 (N_4446,In_858,In_1481);
xor U4447 (N_4447,In_1568,In_2257);
xor U4448 (N_4448,In_2259,In_1430);
and U4449 (N_4449,In_1414,In_575);
and U4450 (N_4450,In_2042,In_371);
or U4451 (N_4451,In_1885,In_1582);
or U4452 (N_4452,In_1932,In_1190);
and U4453 (N_4453,In_1212,In_1872);
nor U4454 (N_4454,In_192,In_486);
and U4455 (N_4455,In_1415,In_2449);
nand U4456 (N_4456,In_2152,In_1417);
nand U4457 (N_4457,In_2499,In_97);
nor U4458 (N_4458,In_1804,In_477);
and U4459 (N_4459,In_470,In_282);
xor U4460 (N_4460,In_1260,In_733);
and U4461 (N_4461,In_1955,In_2059);
xor U4462 (N_4462,In_1681,In_490);
xnor U4463 (N_4463,In_1344,In_1256);
nand U4464 (N_4464,In_101,In_2404);
xnor U4465 (N_4465,In_2008,In_2378);
or U4466 (N_4466,In_2087,In_577);
and U4467 (N_4467,In_1641,In_303);
or U4468 (N_4468,In_2084,In_2076);
nor U4469 (N_4469,In_1341,In_1772);
or U4470 (N_4470,In_1396,In_2133);
xnor U4471 (N_4471,In_1402,In_1327);
nor U4472 (N_4472,In_2043,In_352);
xnor U4473 (N_4473,In_435,In_1487);
nand U4474 (N_4474,In_615,In_362);
and U4475 (N_4475,In_1004,In_2129);
xor U4476 (N_4476,In_1481,In_974);
and U4477 (N_4477,In_684,In_1881);
and U4478 (N_4478,In_69,In_1286);
nor U4479 (N_4479,In_1333,In_1819);
xor U4480 (N_4480,In_1436,In_1303);
nor U4481 (N_4481,In_2002,In_2119);
nor U4482 (N_4482,In_130,In_2402);
xnor U4483 (N_4483,In_2054,In_449);
nor U4484 (N_4484,In_1613,In_2049);
xnor U4485 (N_4485,In_1647,In_1901);
or U4486 (N_4486,In_189,In_1364);
nand U4487 (N_4487,In_1752,In_1036);
xnor U4488 (N_4488,In_2206,In_1008);
nor U4489 (N_4489,In_1218,In_1203);
or U4490 (N_4490,In_2062,In_2256);
or U4491 (N_4491,In_1875,In_1579);
and U4492 (N_4492,In_800,In_756);
xor U4493 (N_4493,In_2250,In_433);
and U4494 (N_4494,In_852,In_477);
nand U4495 (N_4495,In_807,In_2124);
and U4496 (N_4496,In_346,In_1751);
nand U4497 (N_4497,In_1625,In_1920);
nand U4498 (N_4498,In_579,In_2244);
or U4499 (N_4499,In_875,In_2231);
and U4500 (N_4500,In_502,In_153);
and U4501 (N_4501,In_1289,In_1551);
or U4502 (N_4502,In_1948,In_1835);
nand U4503 (N_4503,In_1936,In_245);
nand U4504 (N_4504,In_793,In_637);
nor U4505 (N_4505,In_1542,In_147);
or U4506 (N_4506,In_1784,In_1953);
xnor U4507 (N_4507,In_637,In_639);
and U4508 (N_4508,In_2304,In_964);
or U4509 (N_4509,In_49,In_1289);
and U4510 (N_4510,In_1509,In_1338);
or U4511 (N_4511,In_1526,In_2287);
and U4512 (N_4512,In_212,In_1678);
nor U4513 (N_4513,In_1451,In_1217);
nand U4514 (N_4514,In_2488,In_2402);
or U4515 (N_4515,In_1321,In_2433);
nand U4516 (N_4516,In_538,In_1028);
xor U4517 (N_4517,In_2253,In_1313);
or U4518 (N_4518,In_232,In_680);
nor U4519 (N_4519,In_2465,In_797);
xnor U4520 (N_4520,In_1071,In_879);
nand U4521 (N_4521,In_936,In_17);
nand U4522 (N_4522,In_1817,In_1230);
and U4523 (N_4523,In_968,In_828);
xor U4524 (N_4524,In_84,In_651);
nand U4525 (N_4525,In_0,In_1779);
nand U4526 (N_4526,In_588,In_165);
and U4527 (N_4527,In_142,In_1190);
nand U4528 (N_4528,In_665,In_1266);
or U4529 (N_4529,In_490,In_2154);
nor U4530 (N_4530,In_1607,In_2240);
and U4531 (N_4531,In_367,In_1885);
xor U4532 (N_4532,In_808,In_2044);
or U4533 (N_4533,In_1085,In_1225);
nand U4534 (N_4534,In_2457,In_1636);
nor U4535 (N_4535,In_205,In_890);
nand U4536 (N_4536,In_2314,In_1010);
nand U4537 (N_4537,In_1352,In_1815);
xor U4538 (N_4538,In_391,In_2287);
nand U4539 (N_4539,In_1587,In_1792);
nor U4540 (N_4540,In_827,In_663);
nor U4541 (N_4541,In_86,In_1952);
or U4542 (N_4542,In_2365,In_65);
and U4543 (N_4543,In_1530,In_2419);
nor U4544 (N_4544,In_32,In_2065);
xor U4545 (N_4545,In_2214,In_2102);
nand U4546 (N_4546,In_106,In_696);
and U4547 (N_4547,In_212,In_1048);
or U4548 (N_4548,In_2491,In_1506);
nand U4549 (N_4549,In_885,In_1818);
or U4550 (N_4550,In_1470,In_1180);
or U4551 (N_4551,In_924,In_2155);
xor U4552 (N_4552,In_1395,In_2374);
or U4553 (N_4553,In_1481,In_654);
or U4554 (N_4554,In_550,In_1485);
or U4555 (N_4555,In_813,In_386);
or U4556 (N_4556,In_344,In_1045);
xnor U4557 (N_4557,In_809,In_1762);
and U4558 (N_4558,In_2344,In_1022);
nor U4559 (N_4559,In_2177,In_1983);
and U4560 (N_4560,In_1822,In_1709);
nand U4561 (N_4561,In_362,In_1435);
nand U4562 (N_4562,In_2091,In_1635);
xnor U4563 (N_4563,In_1480,In_1255);
nor U4564 (N_4564,In_1967,In_1659);
nand U4565 (N_4565,In_1821,In_1566);
xor U4566 (N_4566,In_369,In_1196);
nor U4567 (N_4567,In_2230,In_1498);
nand U4568 (N_4568,In_1550,In_787);
nor U4569 (N_4569,In_683,In_2075);
nor U4570 (N_4570,In_328,In_1170);
and U4571 (N_4571,In_1730,In_2483);
or U4572 (N_4572,In_86,In_649);
or U4573 (N_4573,In_1213,In_386);
nand U4574 (N_4574,In_678,In_1858);
nor U4575 (N_4575,In_1786,In_163);
nand U4576 (N_4576,In_606,In_922);
or U4577 (N_4577,In_2086,In_2289);
and U4578 (N_4578,In_2360,In_2208);
nand U4579 (N_4579,In_987,In_405);
nand U4580 (N_4580,In_872,In_2387);
or U4581 (N_4581,In_606,In_763);
xor U4582 (N_4582,In_808,In_1816);
and U4583 (N_4583,In_1357,In_423);
or U4584 (N_4584,In_1688,In_2284);
nand U4585 (N_4585,In_1522,In_914);
or U4586 (N_4586,In_1736,In_940);
or U4587 (N_4587,In_1967,In_279);
or U4588 (N_4588,In_219,In_2362);
nor U4589 (N_4589,In_2098,In_2332);
nor U4590 (N_4590,In_2083,In_2033);
nand U4591 (N_4591,In_1312,In_1386);
and U4592 (N_4592,In_330,In_2004);
and U4593 (N_4593,In_612,In_358);
nand U4594 (N_4594,In_623,In_301);
and U4595 (N_4595,In_126,In_512);
xnor U4596 (N_4596,In_1872,In_2196);
and U4597 (N_4597,In_2396,In_1409);
and U4598 (N_4598,In_1444,In_1354);
nand U4599 (N_4599,In_1749,In_2006);
nand U4600 (N_4600,In_530,In_1020);
xor U4601 (N_4601,In_1440,In_1460);
xnor U4602 (N_4602,In_2351,In_1197);
nand U4603 (N_4603,In_259,In_114);
and U4604 (N_4604,In_2492,In_397);
xor U4605 (N_4605,In_2318,In_1858);
or U4606 (N_4606,In_1345,In_2020);
xor U4607 (N_4607,In_228,In_1172);
or U4608 (N_4608,In_403,In_445);
or U4609 (N_4609,In_1586,In_1362);
xnor U4610 (N_4610,In_2117,In_1078);
and U4611 (N_4611,In_1770,In_337);
nand U4612 (N_4612,In_722,In_643);
or U4613 (N_4613,In_646,In_275);
and U4614 (N_4614,In_1665,In_1583);
nor U4615 (N_4615,In_1902,In_1822);
nand U4616 (N_4616,In_1362,In_1663);
or U4617 (N_4617,In_495,In_186);
and U4618 (N_4618,In_840,In_2127);
and U4619 (N_4619,In_2027,In_353);
nor U4620 (N_4620,In_1005,In_236);
nand U4621 (N_4621,In_606,In_521);
or U4622 (N_4622,In_983,In_414);
xnor U4623 (N_4623,In_1531,In_1776);
and U4624 (N_4624,In_364,In_193);
or U4625 (N_4625,In_2477,In_700);
or U4626 (N_4626,In_212,In_2130);
xor U4627 (N_4627,In_2134,In_2354);
nor U4628 (N_4628,In_1108,In_1822);
and U4629 (N_4629,In_1283,In_1585);
xnor U4630 (N_4630,In_1187,In_1420);
or U4631 (N_4631,In_2179,In_924);
and U4632 (N_4632,In_2348,In_391);
or U4633 (N_4633,In_2045,In_1911);
and U4634 (N_4634,In_1767,In_2446);
and U4635 (N_4635,In_1454,In_2316);
xnor U4636 (N_4636,In_2476,In_2052);
and U4637 (N_4637,In_789,In_1796);
or U4638 (N_4638,In_460,In_1138);
nand U4639 (N_4639,In_672,In_343);
and U4640 (N_4640,In_1715,In_156);
nor U4641 (N_4641,In_407,In_1579);
or U4642 (N_4642,In_524,In_1919);
and U4643 (N_4643,In_1806,In_77);
nand U4644 (N_4644,In_1211,In_921);
or U4645 (N_4645,In_1662,In_1392);
nand U4646 (N_4646,In_519,In_1376);
or U4647 (N_4647,In_1735,In_1289);
or U4648 (N_4648,In_1230,In_622);
nand U4649 (N_4649,In_20,In_1811);
nor U4650 (N_4650,In_731,In_1951);
nand U4651 (N_4651,In_397,In_2385);
xor U4652 (N_4652,In_774,In_1626);
and U4653 (N_4653,In_340,In_53);
nand U4654 (N_4654,In_436,In_1769);
nand U4655 (N_4655,In_1148,In_1925);
or U4656 (N_4656,In_502,In_1350);
nand U4657 (N_4657,In_635,In_1117);
xnor U4658 (N_4658,In_337,In_783);
nor U4659 (N_4659,In_1611,In_75);
nor U4660 (N_4660,In_1902,In_1280);
nand U4661 (N_4661,In_705,In_823);
or U4662 (N_4662,In_1820,In_904);
nor U4663 (N_4663,In_1542,In_1090);
nand U4664 (N_4664,In_2046,In_1050);
nor U4665 (N_4665,In_2432,In_1877);
xnor U4666 (N_4666,In_2478,In_1445);
xor U4667 (N_4667,In_544,In_1878);
nand U4668 (N_4668,In_1344,In_1020);
xnor U4669 (N_4669,In_1396,In_2234);
and U4670 (N_4670,In_917,In_2145);
or U4671 (N_4671,In_528,In_1729);
xor U4672 (N_4672,In_1977,In_1713);
and U4673 (N_4673,In_2057,In_1325);
xnor U4674 (N_4674,In_532,In_1275);
nor U4675 (N_4675,In_2010,In_733);
nand U4676 (N_4676,In_2454,In_1710);
and U4677 (N_4677,In_1391,In_1462);
and U4678 (N_4678,In_2410,In_1711);
xor U4679 (N_4679,In_1860,In_1603);
xnor U4680 (N_4680,In_1807,In_2424);
and U4681 (N_4681,In_1373,In_1889);
nand U4682 (N_4682,In_2453,In_531);
nand U4683 (N_4683,In_2257,In_1826);
or U4684 (N_4684,In_2270,In_625);
nor U4685 (N_4685,In_7,In_1432);
nand U4686 (N_4686,In_1076,In_100);
xnor U4687 (N_4687,In_369,In_1292);
or U4688 (N_4688,In_856,In_169);
nor U4689 (N_4689,In_679,In_2051);
nor U4690 (N_4690,In_1565,In_1508);
nand U4691 (N_4691,In_2144,In_2392);
nor U4692 (N_4692,In_2017,In_1375);
and U4693 (N_4693,In_831,In_1645);
nand U4694 (N_4694,In_1465,In_1593);
nor U4695 (N_4695,In_1382,In_2488);
nor U4696 (N_4696,In_933,In_1526);
nor U4697 (N_4697,In_817,In_750);
nand U4698 (N_4698,In_86,In_2496);
xor U4699 (N_4699,In_1361,In_1053);
nor U4700 (N_4700,In_2294,In_1443);
nand U4701 (N_4701,In_2311,In_476);
nand U4702 (N_4702,In_2238,In_2344);
and U4703 (N_4703,In_1293,In_1074);
or U4704 (N_4704,In_472,In_403);
nor U4705 (N_4705,In_183,In_1035);
nand U4706 (N_4706,In_2055,In_1569);
nor U4707 (N_4707,In_377,In_2301);
nand U4708 (N_4708,In_1561,In_1214);
xor U4709 (N_4709,In_1919,In_2177);
nor U4710 (N_4710,In_1659,In_2038);
nor U4711 (N_4711,In_602,In_982);
xor U4712 (N_4712,In_1663,In_1475);
xnor U4713 (N_4713,In_2097,In_1027);
or U4714 (N_4714,In_486,In_2173);
xor U4715 (N_4715,In_2415,In_251);
or U4716 (N_4716,In_317,In_1081);
or U4717 (N_4717,In_896,In_273);
xnor U4718 (N_4718,In_2137,In_1248);
xnor U4719 (N_4719,In_1642,In_303);
xor U4720 (N_4720,In_140,In_197);
or U4721 (N_4721,In_2353,In_575);
xor U4722 (N_4722,In_1482,In_2026);
nand U4723 (N_4723,In_2446,In_814);
and U4724 (N_4724,In_364,In_2111);
xor U4725 (N_4725,In_1310,In_1858);
xnor U4726 (N_4726,In_575,In_586);
nor U4727 (N_4727,In_2103,In_1355);
and U4728 (N_4728,In_81,In_146);
nand U4729 (N_4729,In_2000,In_1303);
xor U4730 (N_4730,In_1992,In_1054);
xor U4731 (N_4731,In_241,In_1860);
and U4732 (N_4732,In_2467,In_565);
xor U4733 (N_4733,In_1384,In_801);
and U4734 (N_4734,In_646,In_1683);
xor U4735 (N_4735,In_879,In_1468);
nand U4736 (N_4736,In_639,In_1916);
and U4737 (N_4737,In_399,In_1339);
and U4738 (N_4738,In_305,In_1894);
or U4739 (N_4739,In_1644,In_1515);
nor U4740 (N_4740,In_2191,In_1555);
or U4741 (N_4741,In_1047,In_2215);
xor U4742 (N_4742,In_1694,In_1075);
nand U4743 (N_4743,In_1683,In_79);
xor U4744 (N_4744,In_431,In_1673);
nand U4745 (N_4745,In_1985,In_1876);
nor U4746 (N_4746,In_134,In_2112);
nand U4747 (N_4747,In_208,In_474);
or U4748 (N_4748,In_597,In_272);
nor U4749 (N_4749,In_1000,In_628);
or U4750 (N_4750,In_737,In_475);
nand U4751 (N_4751,In_968,In_356);
nor U4752 (N_4752,In_649,In_12);
nor U4753 (N_4753,In_1898,In_2489);
nor U4754 (N_4754,In_2287,In_736);
nand U4755 (N_4755,In_1388,In_137);
nor U4756 (N_4756,In_758,In_610);
and U4757 (N_4757,In_1283,In_1260);
nand U4758 (N_4758,In_1266,In_1735);
or U4759 (N_4759,In_1100,In_1388);
nor U4760 (N_4760,In_44,In_1737);
and U4761 (N_4761,In_169,In_2114);
or U4762 (N_4762,In_764,In_2009);
or U4763 (N_4763,In_1692,In_2352);
nor U4764 (N_4764,In_534,In_178);
nor U4765 (N_4765,In_1564,In_822);
nor U4766 (N_4766,In_577,In_320);
and U4767 (N_4767,In_1057,In_2313);
xnor U4768 (N_4768,In_2424,In_1984);
nand U4769 (N_4769,In_99,In_1052);
and U4770 (N_4770,In_898,In_142);
and U4771 (N_4771,In_1702,In_465);
xnor U4772 (N_4772,In_667,In_2159);
and U4773 (N_4773,In_2452,In_1098);
nor U4774 (N_4774,In_1490,In_333);
and U4775 (N_4775,In_2437,In_529);
and U4776 (N_4776,In_2272,In_2020);
or U4777 (N_4777,In_1662,In_2011);
nor U4778 (N_4778,In_487,In_1664);
nand U4779 (N_4779,In_341,In_788);
xor U4780 (N_4780,In_1882,In_1010);
nor U4781 (N_4781,In_2387,In_2163);
xor U4782 (N_4782,In_2486,In_1852);
xnor U4783 (N_4783,In_669,In_2189);
and U4784 (N_4784,In_2470,In_1837);
or U4785 (N_4785,In_456,In_1504);
or U4786 (N_4786,In_820,In_641);
and U4787 (N_4787,In_1067,In_280);
or U4788 (N_4788,In_2151,In_2163);
or U4789 (N_4789,In_539,In_1616);
or U4790 (N_4790,In_915,In_1732);
xor U4791 (N_4791,In_452,In_77);
and U4792 (N_4792,In_2396,In_753);
nor U4793 (N_4793,In_1705,In_1452);
or U4794 (N_4794,In_457,In_217);
xnor U4795 (N_4795,In_1990,In_2006);
nor U4796 (N_4796,In_641,In_2444);
nor U4797 (N_4797,In_620,In_1267);
xnor U4798 (N_4798,In_2178,In_1954);
xor U4799 (N_4799,In_1487,In_1089);
xor U4800 (N_4800,In_2154,In_881);
xnor U4801 (N_4801,In_1078,In_791);
and U4802 (N_4802,In_2098,In_2157);
nor U4803 (N_4803,In_1765,In_1229);
and U4804 (N_4804,In_483,In_2160);
and U4805 (N_4805,In_729,In_191);
xnor U4806 (N_4806,In_1850,In_737);
nand U4807 (N_4807,In_35,In_2380);
nor U4808 (N_4808,In_478,In_1888);
nand U4809 (N_4809,In_1674,In_764);
nand U4810 (N_4810,In_1883,In_1700);
or U4811 (N_4811,In_584,In_286);
and U4812 (N_4812,In_2164,In_2179);
nor U4813 (N_4813,In_1885,In_2244);
or U4814 (N_4814,In_1414,In_2205);
nor U4815 (N_4815,In_143,In_1760);
and U4816 (N_4816,In_1905,In_2165);
nand U4817 (N_4817,In_2126,In_1727);
nand U4818 (N_4818,In_203,In_1186);
nand U4819 (N_4819,In_580,In_1232);
xnor U4820 (N_4820,In_1465,In_14);
and U4821 (N_4821,In_151,In_1001);
or U4822 (N_4822,In_759,In_730);
xnor U4823 (N_4823,In_383,In_2472);
nand U4824 (N_4824,In_2165,In_445);
and U4825 (N_4825,In_1704,In_1312);
nor U4826 (N_4826,In_2210,In_1549);
xor U4827 (N_4827,In_1277,In_2239);
and U4828 (N_4828,In_1618,In_2033);
or U4829 (N_4829,In_1857,In_335);
xnor U4830 (N_4830,In_1306,In_1855);
xnor U4831 (N_4831,In_2043,In_1586);
xnor U4832 (N_4832,In_2320,In_993);
or U4833 (N_4833,In_2455,In_339);
and U4834 (N_4834,In_213,In_1624);
nand U4835 (N_4835,In_514,In_1224);
nor U4836 (N_4836,In_318,In_797);
or U4837 (N_4837,In_1614,In_2459);
nor U4838 (N_4838,In_2215,In_1154);
nor U4839 (N_4839,In_24,In_1147);
nor U4840 (N_4840,In_2128,In_1290);
nand U4841 (N_4841,In_1915,In_2315);
nor U4842 (N_4842,In_1631,In_266);
nor U4843 (N_4843,In_864,In_544);
and U4844 (N_4844,In_254,In_65);
nor U4845 (N_4845,In_2205,In_825);
or U4846 (N_4846,In_1031,In_698);
xnor U4847 (N_4847,In_450,In_58);
or U4848 (N_4848,In_2431,In_488);
xor U4849 (N_4849,In_1431,In_433);
and U4850 (N_4850,In_73,In_1856);
or U4851 (N_4851,In_691,In_2338);
nor U4852 (N_4852,In_1354,In_1877);
xor U4853 (N_4853,In_1947,In_2454);
xor U4854 (N_4854,In_1719,In_2109);
and U4855 (N_4855,In_2396,In_597);
and U4856 (N_4856,In_961,In_1596);
and U4857 (N_4857,In_468,In_667);
xnor U4858 (N_4858,In_1754,In_2146);
and U4859 (N_4859,In_1138,In_297);
or U4860 (N_4860,In_941,In_428);
or U4861 (N_4861,In_860,In_1392);
and U4862 (N_4862,In_2225,In_1637);
nor U4863 (N_4863,In_1737,In_1610);
xnor U4864 (N_4864,In_947,In_1604);
nand U4865 (N_4865,In_936,In_2380);
nand U4866 (N_4866,In_1342,In_2211);
and U4867 (N_4867,In_672,In_144);
nor U4868 (N_4868,In_729,In_1638);
xnor U4869 (N_4869,In_1094,In_2496);
or U4870 (N_4870,In_965,In_450);
xor U4871 (N_4871,In_1955,In_1476);
nand U4872 (N_4872,In_568,In_2456);
or U4873 (N_4873,In_1172,In_391);
nand U4874 (N_4874,In_1548,In_122);
and U4875 (N_4875,In_1666,In_317);
and U4876 (N_4876,In_115,In_421);
and U4877 (N_4877,In_107,In_2485);
xnor U4878 (N_4878,In_1814,In_868);
or U4879 (N_4879,In_635,In_2204);
nor U4880 (N_4880,In_233,In_396);
nand U4881 (N_4881,In_1540,In_1551);
nor U4882 (N_4882,In_67,In_1055);
nand U4883 (N_4883,In_1177,In_890);
nor U4884 (N_4884,In_272,In_2316);
xnor U4885 (N_4885,In_921,In_2395);
or U4886 (N_4886,In_1764,In_730);
xor U4887 (N_4887,In_1686,In_100);
nand U4888 (N_4888,In_1823,In_1352);
nand U4889 (N_4889,In_895,In_2161);
or U4890 (N_4890,In_511,In_1613);
xor U4891 (N_4891,In_882,In_1178);
nor U4892 (N_4892,In_1250,In_1935);
nand U4893 (N_4893,In_2075,In_1912);
or U4894 (N_4894,In_20,In_387);
nor U4895 (N_4895,In_1456,In_638);
nand U4896 (N_4896,In_1454,In_2252);
nand U4897 (N_4897,In_2190,In_109);
nand U4898 (N_4898,In_1832,In_1348);
and U4899 (N_4899,In_166,In_367);
and U4900 (N_4900,In_1905,In_1800);
xor U4901 (N_4901,In_1166,In_225);
nor U4902 (N_4902,In_410,In_435);
and U4903 (N_4903,In_60,In_2006);
or U4904 (N_4904,In_464,In_1519);
nand U4905 (N_4905,In_1686,In_678);
and U4906 (N_4906,In_1746,In_1588);
and U4907 (N_4907,In_1663,In_2001);
or U4908 (N_4908,In_1368,In_602);
nand U4909 (N_4909,In_1791,In_2242);
and U4910 (N_4910,In_726,In_305);
nor U4911 (N_4911,In_329,In_2354);
nor U4912 (N_4912,In_241,In_200);
xor U4913 (N_4913,In_278,In_1495);
xnor U4914 (N_4914,In_980,In_2411);
nor U4915 (N_4915,In_1367,In_1056);
and U4916 (N_4916,In_1299,In_822);
nor U4917 (N_4917,In_973,In_971);
xor U4918 (N_4918,In_1239,In_124);
or U4919 (N_4919,In_1946,In_849);
and U4920 (N_4920,In_1537,In_1265);
nand U4921 (N_4921,In_422,In_108);
xor U4922 (N_4922,In_262,In_2137);
xnor U4923 (N_4923,In_2278,In_1368);
nor U4924 (N_4924,In_30,In_253);
nand U4925 (N_4925,In_266,In_1606);
xor U4926 (N_4926,In_1856,In_1945);
xor U4927 (N_4927,In_2001,In_879);
or U4928 (N_4928,In_2475,In_1459);
xnor U4929 (N_4929,In_2498,In_360);
and U4930 (N_4930,In_337,In_810);
nand U4931 (N_4931,In_1347,In_645);
nand U4932 (N_4932,In_379,In_1801);
nand U4933 (N_4933,In_2034,In_1789);
nor U4934 (N_4934,In_712,In_2222);
xnor U4935 (N_4935,In_1642,In_468);
or U4936 (N_4936,In_2415,In_222);
xor U4937 (N_4937,In_1025,In_1906);
nand U4938 (N_4938,In_674,In_489);
or U4939 (N_4939,In_1911,In_413);
nor U4940 (N_4940,In_110,In_293);
nor U4941 (N_4941,In_313,In_1308);
nor U4942 (N_4942,In_1421,In_1636);
nor U4943 (N_4943,In_1477,In_1895);
xnor U4944 (N_4944,In_2268,In_842);
nand U4945 (N_4945,In_949,In_1771);
nor U4946 (N_4946,In_1009,In_1533);
or U4947 (N_4947,In_1467,In_132);
or U4948 (N_4948,In_1776,In_827);
xnor U4949 (N_4949,In_978,In_1990);
nor U4950 (N_4950,In_784,In_1568);
and U4951 (N_4951,In_101,In_1082);
and U4952 (N_4952,In_1076,In_1684);
or U4953 (N_4953,In_2248,In_1354);
or U4954 (N_4954,In_920,In_395);
and U4955 (N_4955,In_1817,In_1410);
xnor U4956 (N_4956,In_896,In_279);
or U4957 (N_4957,In_1922,In_2488);
or U4958 (N_4958,In_485,In_2267);
nand U4959 (N_4959,In_917,In_848);
xor U4960 (N_4960,In_1805,In_1683);
xnor U4961 (N_4961,In_2126,In_2452);
nor U4962 (N_4962,In_706,In_314);
or U4963 (N_4963,In_2211,In_982);
nor U4964 (N_4964,In_1566,In_2112);
xnor U4965 (N_4965,In_2091,In_705);
and U4966 (N_4966,In_2458,In_610);
nand U4967 (N_4967,In_728,In_187);
xnor U4968 (N_4968,In_1804,In_1157);
and U4969 (N_4969,In_1787,In_349);
xor U4970 (N_4970,In_1122,In_2405);
xnor U4971 (N_4971,In_397,In_1837);
nor U4972 (N_4972,In_996,In_1656);
or U4973 (N_4973,In_838,In_1839);
xor U4974 (N_4974,In_74,In_2188);
or U4975 (N_4975,In_808,In_1222);
nand U4976 (N_4976,In_801,In_996);
nor U4977 (N_4977,In_701,In_714);
nand U4978 (N_4978,In_2368,In_1259);
nor U4979 (N_4979,In_2250,In_1146);
or U4980 (N_4980,In_2079,In_1062);
nand U4981 (N_4981,In_2482,In_747);
nand U4982 (N_4982,In_957,In_712);
nor U4983 (N_4983,In_1431,In_143);
xor U4984 (N_4984,In_2298,In_1971);
nand U4985 (N_4985,In_2412,In_523);
nand U4986 (N_4986,In_1827,In_1029);
xor U4987 (N_4987,In_1963,In_1479);
and U4988 (N_4988,In_724,In_704);
nor U4989 (N_4989,In_54,In_1240);
or U4990 (N_4990,In_1189,In_1858);
nand U4991 (N_4991,In_322,In_1271);
nor U4992 (N_4992,In_1027,In_953);
nand U4993 (N_4993,In_2,In_898);
or U4994 (N_4994,In_825,In_114);
nor U4995 (N_4995,In_2002,In_1138);
xnor U4996 (N_4996,In_326,In_1676);
nand U4997 (N_4997,In_168,In_396);
and U4998 (N_4998,In_2144,In_744);
nand U4999 (N_4999,In_1542,In_226);
nand U5000 (N_5000,N_1644,N_3869);
or U5001 (N_5001,N_887,N_444);
nor U5002 (N_5002,N_174,N_3921);
or U5003 (N_5003,N_1491,N_1762);
xor U5004 (N_5004,N_2332,N_2964);
and U5005 (N_5005,N_74,N_1541);
and U5006 (N_5006,N_283,N_752);
and U5007 (N_5007,N_833,N_1376);
nand U5008 (N_5008,N_1709,N_620);
nand U5009 (N_5009,N_908,N_2911);
or U5010 (N_5010,N_1521,N_4047);
or U5011 (N_5011,N_4207,N_923);
nor U5012 (N_5012,N_1140,N_4567);
or U5013 (N_5013,N_4635,N_4757);
nand U5014 (N_5014,N_2074,N_3237);
or U5015 (N_5015,N_195,N_4241);
xnor U5016 (N_5016,N_4524,N_1134);
and U5017 (N_5017,N_323,N_3002);
and U5018 (N_5018,N_2054,N_4147);
xnor U5019 (N_5019,N_3733,N_458);
nand U5020 (N_5020,N_3997,N_301);
nand U5021 (N_5021,N_2661,N_2608);
or U5022 (N_5022,N_4281,N_555);
or U5023 (N_5023,N_188,N_2961);
nand U5024 (N_5024,N_1595,N_2772);
nor U5025 (N_5025,N_3969,N_4965);
nand U5026 (N_5026,N_29,N_1857);
nor U5027 (N_5027,N_4776,N_3666);
xor U5028 (N_5028,N_3612,N_2918);
or U5029 (N_5029,N_2299,N_4943);
xnor U5030 (N_5030,N_1648,N_2938);
and U5031 (N_5031,N_1518,N_3147);
xor U5032 (N_5032,N_3582,N_3179);
and U5033 (N_5033,N_3896,N_4068);
or U5034 (N_5034,N_4800,N_4665);
and U5035 (N_5035,N_1933,N_280);
xor U5036 (N_5036,N_3392,N_66);
and U5037 (N_5037,N_1751,N_1574);
xor U5038 (N_5038,N_1139,N_3359);
or U5039 (N_5039,N_281,N_2977);
xnor U5040 (N_5040,N_1112,N_1668);
xor U5041 (N_5041,N_4124,N_2687);
xor U5042 (N_5042,N_1611,N_4354);
xnor U5043 (N_5043,N_4317,N_3708);
or U5044 (N_5044,N_4177,N_2878);
and U5045 (N_5045,N_1961,N_1510);
and U5046 (N_5046,N_1717,N_825);
nor U5047 (N_5047,N_890,N_3668);
xnor U5048 (N_5048,N_4821,N_884);
xnor U5049 (N_5049,N_519,N_1216);
or U5050 (N_5050,N_2417,N_2239);
nand U5051 (N_5051,N_2044,N_1602);
or U5052 (N_5052,N_581,N_3916);
xnor U5053 (N_5053,N_1699,N_1393);
xnor U5054 (N_5054,N_661,N_2951);
or U5055 (N_5055,N_3994,N_4153);
nor U5056 (N_5056,N_1652,N_851);
nor U5057 (N_5057,N_872,N_2512);
and U5058 (N_5058,N_2526,N_1424);
and U5059 (N_5059,N_2462,N_2719);
nand U5060 (N_5060,N_3979,N_1353);
or U5061 (N_5061,N_2221,N_2415);
and U5062 (N_5062,N_1358,N_3320);
nor U5063 (N_5063,N_1629,N_2115);
or U5064 (N_5064,N_350,N_2756);
or U5065 (N_5065,N_3105,N_1210);
and U5066 (N_5066,N_3630,N_952);
and U5067 (N_5067,N_1303,N_2544);
nor U5068 (N_5068,N_3739,N_4631);
and U5069 (N_5069,N_2550,N_1223);
xor U5070 (N_5070,N_62,N_2319);
xor U5071 (N_5071,N_4441,N_2706);
nor U5072 (N_5072,N_4710,N_127);
nor U5073 (N_5073,N_3923,N_1990);
nor U5074 (N_5074,N_4802,N_4179);
nor U5075 (N_5075,N_2580,N_4095);
xor U5076 (N_5076,N_2017,N_891);
nand U5077 (N_5077,N_1721,N_502);
nand U5078 (N_5078,N_1664,N_2540);
or U5079 (N_5079,N_3177,N_4211);
nand U5080 (N_5080,N_2869,N_1076);
nand U5081 (N_5081,N_3611,N_4127);
nor U5082 (N_5082,N_1401,N_2351);
nand U5083 (N_5083,N_1890,N_968);
nor U5084 (N_5084,N_3955,N_4442);
and U5085 (N_5085,N_1119,N_4597);
nor U5086 (N_5086,N_107,N_4148);
and U5087 (N_5087,N_3149,N_1658);
or U5088 (N_5088,N_1632,N_1921);
xnor U5089 (N_5089,N_3245,N_284);
xnor U5090 (N_5090,N_3389,N_1844);
xnor U5091 (N_5091,N_3401,N_2454);
xor U5092 (N_5092,N_1916,N_4426);
and U5093 (N_5093,N_332,N_114);
nand U5094 (N_5094,N_935,N_2638);
and U5095 (N_5095,N_3057,N_1350);
and U5096 (N_5096,N_623,N_1368);
xor U5097 (N_5097,N_456,N_1555);
and U5098 (N_5098,N_4964,N_4120);
or U5099 (N_5099,N_1593,N_2065);
nand U5100 (N_5100,N_4592,N_4036);
xor U5101 (N_5101,N_3367,N_582);
and U5102 (N_5102,N_1863,N_2585);
nor U5103 (N_5103,N_1600,N_4909);
and U5104 (N_5104,N_4937,N_3629);
nor U5105 (N_5105,N_3614,N_4480);
xnor U5106 (N_5106,N_1724,N_4850);
or U5107 (N_5107,N_4297,N_2433);
nand U5108 (N_5108,N_2457,N_2675);
nor U5109 (N_5109,N_2244,N_123);
xnor U5110 (N_5110,N_2262,N_3269);
or U5111 (N_5111,N_4612,N_3220);
nor U5112 (N_5112,N_3112,N_4764);
and U5113 (N_5113,N_4078,N_2695);
and U5114 (N_5114,N_4141,N_3837);
nand U5115 (N_5115,N_3381,N_2212);
nor U5116 (N_5116,N_3360,N_530);
nor U5117 (N_5117,N_4942,N_1737);
xnor U5118 (N_5118,N_4131,N_2743);
nand U5119 (N_5119,N_1716,N_98);
nand U5120 (N_5120,N_3510,N_3476);
or U5121 (N_5121,N_4791,N_1498);
nor U5122 (N_5122,N_4958,N_233);
or U5123 (N_5123,N_1581,N_2431);
nand U5124 (N_5124,N_941,N_2223);
or U5125 (N_5125,N_2396,N_737);
nor U5126 (N_5126,N_4194,N_4687);
nor U5127 (N_5127,N_1936,N_983);
nand U5128 (N_5128,N_2592,N_4707);
or U5129 (N_5129,N_4443,N_3142);
or U5130 (N_5130,N_2984,N_4672);
and U5131 (N_5131,N_4115,N_848);
nor U5132 (N_5132,N_554,N_3995);
xnor U5133 (N_5133,N_2099,N_2724);
and U5134 (N_5134,N_4572,N_1516);
nand U5135 (N_5135,N_3346,N_1601);
xnor U5136 (N_5136,N_550,N_2407);
or U5137 (N_5137,N_2149,N_683);
or U5138 (N_5138,N_1887,N_2901);
and U5139 (N_5139,N_4960,N_2643);
nor U5140 (N_5140,N_770,N_3227);
or U5141 (N_5141,N_3079,N_1000);
nand U5142 (N_5142,N_2755,N_408);
or U5143 (N_5143,N_4178,N_1261);
and U5144 (N_5144,N_788,N_4807);
nor U5145 (N_5145,N_1725,N_4984);
nand U5146 (N_5146,N_3628,N_3230);
nand U5147 (N_5147,N_3756,N_2032);
and U5148 (N_5148,N_4013,N_1435);
nor U5149 (N_5149,N_1964,N_466);
nand U5150 (N_5150,N_3566,N_1983);
nor U5151 (N_5151,N_1421,N_2078);
xor U5152 (N_5152,N_3802,N_1116);
nor U5153 (N_5153,N_599,N_398);
or U5154 (N_5154,N_3115,N_808);
and U5155 (N_5155,N_565,N_3194);
nor U5156 (N_5156,N_3729,N_538);
or U5157 (N_5157,N_447,N_4638);
nor U5158 (N_5158,N_4461,N_616);
or U5159 (N_5159,N_1084,N_347);
nor U5160 (N_5160,N_1826,N_871);
nand U5161 (N_5161,N_2047,N_901);
xnor U5162 (N_5162,N_3011,N_3328);
and U5163 (N_5163,N_1092,N_4067);
xnor U5164 (N_5164,N_2980,N_3319);
nor U5165 (N_5165,N_1337,N_3085);
nor U5166 (N_5166,N_4470,N_433);
nand U5167 (N_5167,N_4840,N_4420);
nand U5168 (N_5168,N_1094,N_3981);
nor U5169 (N_5169,N_1646,N_4924);
nand U5170 (N_5170,N_4111,N_2944);
nor U5171 (N_5171,N_4272,N_694);
xnor U5172 (N_5172,N_1722,N_4903);
xnor U5173 (N_5173,N_2628,N_1891);
or U5174 (N_5174,N_747,N_2776);
nand U5175 (N_5175,N_1038,N_2558);
and U5176 (N_5176,N_978,N_4323);
xnor U5177 (N_5177,N_1158,N_4431);
nor U5178 (N_5178,N_3196,N_4228);
nor U5179 (N_5179,N_4140,N_3260);
nor U5180 (N_5180,N_2525,N_4787);
nor U5181 (N_5181,N_2303,N_4182);
or U5182 (N_5182,N_3838,N_3405);
or U5183 (N_5183,N_2258,N_2910);
nor U5184 (N_5184,N_416,N_4428);
and U5185 (N_5185,N_200,N_3373);
nor U5186 (N_5186,N_4049,N_757);
or U5187 (N_5187,N_1986,N_4401);
nor U5188 (N_5188,N_4042,N_86);
and U5189 (N_5189,N_4685,N_1788);
xnor U5190 (N_5190,N_101,N_972);
or U5191 (N_5191,N_2718,N_3407);
and U5192 (N_5192,N_239,N_4172);
and U5193 (N_5193,N_4970,N_3096);
or U5194 (N_5194,N_80,N_3604);
and U5195 (N_5195,N_4726,N_847);
or U5196 (N_5196,N_4129,N_2921);
and U5197 (N_5197,N_4669,N_2682);
xnor U5198 (N_5198,N_4076,N_4879);
xor U5199 (N_5199,N_3781,N_758);
xnor U5200 (N_5200,N_1163,N_1911);
or U5201 (N_5201,N_393,N_1448);
and U5202 (N_5202,N_1395,N_4526);
nor U5203 (N_5203,N_4366,N_63);
or U5204 (N_5204,N_453,N_489);
or U5205 (N_5205,N_4195,N_2022);
or U5206 (N_5206,N_4571,N_994);
nand U5207 (N_5207,N_1364,N_1228);
and U5208 (N_5208,N_4629,N_1299);
xor U5209 (N_5209,N_4652,N_3014);
xnor U5210 (N_5210,N_3832,N_2084);
or U5211 (N_5211,N_627,N_2676);
nor U5212 (N_5212,N_1948,N_4870);
and U5213 (N_5213,N_3337,N_4615);
xor U5214 (N_5214,N_1615,N_763);
nor U5215 (N_5215,N_3653,N_3546);
xnor U5216 (N_5216,N_3287,N_4214);
xor U5217 (N_5217,N_3038,N_3141);
or U5218 (N_5218,N_1314,N_2920);
nand U5219 (N_5219,N_729,N_1344);
or U5220 (N_5220,N_2722,N_491);
xnor U5221 (N_5221,N_4093,N_3847);
nand U5222 (N_5222,N_3491,N_3762);
xor U5223 (N_5223,N_4543,N_4642);
nand U5224 (N_5224,N_3641,N_108);
and U5225 (N_5225,N_2527,N_2036);
and U5226 (N_5226,N_4537,N_787);
nor U5227 (N_5227,N_2751,N_2232);
xor U5228 (N_5228,N_3732,N_51);
and U5229 (N_5229,N_2173,N_1509);
and U5230 (N_5230,N_897,N_1482);
or U5231 (N_5231,N_4,N_4413);
nand U5232 (N_5232,N_256,N_1870);
and U5233 (N_5233,N_1682,N_2157);
nor U5234 (N_5234,N_2038,N_2874);
nor U5235 (N_5235,N_3228,N_3270);
nor U5236 (N_5236,N_849,N_3284);
nand U5237 (N_5237,N_2632,N_3345);
nor U5238 (N_5238,N_4768,N_120);
or U5239 (N_5239,N_1693,N_1930);
or U5240 (N_5240,N_4482,N_2147);
and U5241 (N_5241,N_109,N_4722);
nand U5242 (N_5242,N_1757,N_1627);
xnor U5243 (N_5243,N_471,N_3996);
and U5244 (N_5244,N_3503,N_861);
nand U5245 (N_5245,N_641,N_883);
nand U5246 (N_5246,N_1355,N_1322);
and U5247 (N_5247,N_2161,N_512);
xor U5248 (N_5248,N_1548,N_3253);
xnor U5249 (N_5249,N_2761,N_2859);
and U5250 (N_5250,N_4923,N_922);
and U5251 (N_5251,N_3616,N_2474);
and U5252 (N_5252,N_2081,N_2946);
or U5253 (N_5253,N_2420,N_3517);
or U5254 (N_5254,N_2636,N_2919);
xor U5255 (N_5255,N_4041,N_544);
nand U5256 (N_5256,N_2736,N_4070);
nor U5257 (N_5257,N_4103,N_1504);
and U5258 (N_5258,N_2563,N_2680);
xnor U5259 (N_5259,N_3882,N_2155);
and U5260 (N_5260,N_663,N_638);
xor U5261 (N_5261,N_1069,N_569);
nand U5262 (N_5262,N_682,N_4250);
and U5263 (N_5263,N_3782,N_1767);
nor U5264 (N_5264,N_4318,N_1590);
nand U5265 (N_5265,N_1256,N_1404);
xnor U5266 (N_5266,N_4562,N_1596);
and U5267 (N_5267,N_56,N_2520);
nor U5268 (N_5268,N_1825,N_3192);
xor U5269 (N_5269,N_1955,N_3158);
and U5270 (N_5270,N_331,N_2904);
nand U5271 (N_5271,N_3601,N_3099);
and U5272 (N_5272,N_1289,N_1793);
or U5273 (N_5273,N_1397,N_2335);
nand U5274 (N_5274,N_3827,N_3674);
nor U5275 (N_5275,N_804,N_2483);
nor U5276 (N_5276,N_1283,N_1422);
and U5277 (N_5277,N_946,N_4555);
xor U5278 (N_5278,N_4065,N_4229);
nand U5279 (N_5279,N_754,N_859);
or U5280 (N_5280,N_4775,N_2488);
and U5281 (N_5281,N_4026,N_4398);
nand U5282 (N_5282,N_828,N_4027);
or U5283 (N_5283,N_2350,N_2179);
or U5284 (N_5284,N_4458,N_2088);
xnor U5285 (N_5285,N_4678,N_4599);
xor U5286 (N_5286,N_4873,N_4434);
nand U5287 (N_5287,N_103,N_2400);
nor U5288 (N_5288,N_2289,N_1202);
and U5289 (N_5289,N_1102,N_3458);
or U5290 (N_5290,N_3252,N_412);
xnor U5291 (N_5291,N_617,N_4163);
nor U5292 (N_5292,N_3723,N_1711);
and U5293 (N_5293,N_2589,N_4002);
nor U5294 (N_5294,N_3800,N_699);
or U5295 (N_5295,N_401,N_3484);
nor U5296 (N_5296,N_3754,N_4106);
xnor U5297 (N_5297,N_3265,N_4288);
nand U5298 (N_5298,N_3817,N_2456);
or U5299 (N_5299,N_571,N_4948);
xor U5300 (N_5300,N_2178,N_141);
nor U5301 (N_5301,N_3243,N_2771);
nand U5302 (N_5302,N_3530,N_2711);
nor U5303 (N_5303,N_2056,N_2143);
nor U5304 (N_5304,N_1053,N_2669);
or U5305 (N_5305,N_4711,N_3526);
and U5306 (N_5306,N_1583,N_1044);
and U5307 (N_5307,N_3578,N_335);
nand U5308 (N_5308,N_2333,N_1399);
nand U5309 (N_5309,N_1829,N_3675);
xor U5310 (N_5310,N_693,N_1167);
and U5311 (N_5311,N_2037,N_2658);
and U5312 (N_5312,N_3884,N_1425);
nand U5313 (N_5313,N_710,N_2269);
nor U5314 (N_5314,N_4114,N_3704);
xor U5315 (N_5315,N_25,N_1275);
xor U5316 (N_5316,N_1057,N_765);
nor U5317 (N_5317,N_1334,N_372);
nand U5318 (N_5318,N_4246,N_1315);
and U5319 (N_5319,N_1070,N_834);
xor U5320 (N_5320,N_1673,N_2180);
xor U5321 (N_5321,N_1237,N_3101);
xnor U5322 (N_5322,N_3790,N_3306);
xor U5323 (N_5323,N_50,N_4940);
xor U5324 (N_5324,N_723,N_1843);
and U5325 (N_5325,N_4059,N_1129);
xnor U5326 (N_5326,N_1416,N_4337);
or U5327 (N_5327,N_2888,N_839);
and U5328 (N_5328,N_1628,N_3998);
and U5329 (N_5329,N_3543,N_3071);
and U5330 (N_5330,N_591,N_4892);
or U5331 (N_5331,N_465,N_2359);
and U5332 (N_5332,N_2356,N_3792);
or U5333 (N_5333,N_1471,N_3555);
nand U5334 (N_5334,N_4077,N_4038);
or U5335 (N_5335,N_12,N_662);
and U5336 (N_5336,N_2610,N_3326);
and U5337 (N_5337,N_23,N_3308);
nor U5338 (N_5338,N_4959,N_2519);
and U5339 (N_5339,N_1492,N_1527);
and U5340 (N_5340,N_1390,N_3868);
and U5341 (N_5341,N_2045,N_905);
and U5342 (N_5342,N_4302,N_572);
nand U5343 (N_5343,N_4412,N_4770);
xnor U5344 (N_5344,N_4116,N_4183);
and U5345 (N_5345,N_159,N_3897);
or U5346 (N_5346,N_2413,N_1433);
nand U5347 (N_5347,N_2322,N_2987);
nand U5348 (N_5348,N_131,N_3039);
xnor U5349 (N_5349,N_337,N_1319);
and U5350 (N_5350,N_3056,N_1382);
and U5351 (N_5351,N_4432,N_4508);
nor U5352 (N_5352,N_4450,N_448);
nand U5353 (N_5353,N_3086,N_3008);
and U5354 (N_5354,N_61,N_4706);
or U5355 (N_5355,N_4738,N_1500);
nand U5356 (N_5356,N_2886,N_2272);
nand U5357 (N_5357,N_3174,N_944);
xor U5358 (N_5358,N_810,N_966);
nand U5359 (N_5359,N_4545,N_4831);
nand U5360 (N_5360,N_1502,N_1079);
or U5361 (N_5361,N_4590,N_1061);
nor U5362 (N_5362,N_1630,N_4091);
nor U5363 (N_5363,N_318,N_1852);
nor U5364 (N_5364,N_2264,N_3931);
nor U5365 (N_5365,N_4627,N_235);
or U5366 (N_5366,N_1209,N_786);
xnor U5367 (N_5367,N_2249,N_2963);
or U5368 (N_5368,N_3957,N_1943);
nor U5369 (N_5369,N_3028,N_2891);
or U5370 (N_5370,N_2915,N_1408);
and U5371 (N_5371,N_958,N_313);
or U5372 (N_5372,N_230,N_509);
or U5373 (N_5373,N_4805,N_1525);
nor U5374 (N_5374,N_4836,N_4573);
or U5375 (N_5375,N_1173,N_2954);
nand U5376 (N_5376,N_516,N_4872);
or U5377 (N_5377,N_3460,N_4989);
nand U5378 (N_5378,N_494,N_77);
and U5379 (N_5379,N_410,N_3844);
xor U5380 (N_5380,N_2300,N_3579);
nor U5381 (N_5381,N_2428,N_1293);
nor U5382 (N_5382,N_3662,N_138);
nor U5383 (N_5383,N_88,N_4644);
and U5384 (N_5384,N_422,N_4210);
nand U5385 (N_5385,N_3833,N_4634);
xnor U5386 (N_5386,N_2040,N_3089);
and U5387 (N_5387,N_1241,N_3342);
or U5388 (N_5388,N_1288,N_3788);
or U5389 (N_5389,N_2740,N_304);
nand U5390 (N_5390,N_943,N_3077);
xor U5391 (N_5391,N_3163,N_4176);
xnor U5392 (N_5392,N_3670,N_4294);
or U5393 (N_5393,N_4563,N_1892);
xnor U5394 (N_5394,N_367,N_2288);
nand U5395 (N_5395,N_608,N_1147);
xnor U5396 (N_5396,N_1812,N_1791);
and U5397 (N_5397,N_1406,N_1015);
and U5398 (N_5398,N_237,N_495);
or U5399 (N_5399,N_4857,N_6);
nor U5400 (N_5400,N_4453,N_3676);
nand U5401 (N_5401,N_170,N_689);
or U5402 (N_5402,N_4957,N_2245);
nor U5403 (N_5403,N_3726,N_1675);
nand U5404 (N_5404,N_3766,N_4395);
or U5405 (N_5405,N_999,N_2256);
nor U5406 (N_5406,N_3903,N_4976);
and U5407 (N_5407,N_3883,N_329);
and U5408 (N_5408,N_17,N_3499);
xnor U5409 (N_5409,N_250,N_3962);
and U5410 (N_5410,N_567,N_48);
nand U5411 (N_5411,N_4589,N_2116);
nor U5412 (N_5412,N_1691,N_1940);
or U5413 (N_5413,N_4494,N_2323);
or U5414 (N_5414,N_2897,N_4978);
nand U5415 (N_5415,N_576,N_3712);
nand U5416 (N_5416,N_360,N_1765);
nor U5417 (N_5417,N_135,N_1871);
and U5418 (N_5418,N_3012,N_1437);
or U5419 (N_5419,N_388,N_3631);
and U5420 (N_5420,N_4454,N_1861);
nand U5421 (N_5421,N_3752,N_4295);
or U5422 (N_5422,N_180,N_252);
nand U5423 (N_5423,N_612,N_1731);
nand U5424 (N_5424,N_52,N_1515);
or U5425 (N_5425,N_3574,N_1589);
and U5426 (N_5426,N_3561,N_2279);
and U5427 (N_5427,N_1313,N_4818);
nand U5428 (N_5428,N_2294,N_1227);
nor U5429 (N_5429,N_1738,N_1698);
nand U5430 (N_5430,N_3169,N_4033);
nor U5431 (N_5431,N_3030,N_1660);
nor U5432 (N_5432,N_603,N_2554);
nand U5433 (N_5433,N_2739,N_4209);
nor U5434 (N_5434,N_4783,N_124);
nor U5435 (N_5435,N_115,N_1306);
xor U5436 (N_5436,N_4702,N_24);
or U5437 (N_5437,N_4915,N_2060);
nor U5438 (N_5438,N_1872,N_2206);
or U5439 (N_5439,N_1957,N_4919);
nor U5440 (N_5440,N_3070,N_724);
and U5441 (N_5441,N_1584,N_3727);
and U5442 (N_5442,N_1922,N_3454);
nor U5443 (N_5443,N_832,N_3785);
nor U5444 (N_5444,N_579,N_2847);
and U5445 (N_5445,N_163,N_1618);
and U5446 (N_5446,N_4893,N_3182);
xor U5447 (N_5447,N_3572,N_54);
or U5448 (N_5448,N_3534,N_2260);
xor U5449 (N_5449,N_525,N_2418);
nand U5450 (N_5450,N_4826,N_2731);
xor U5451 (N_5451,N_1184,N_2553);
nand U5452 (N_5452,N_3294,N_3563);
or U5453 (N_5453,N_4012,N_3855);
nand U5454 (N_5454,N_3451,N_2893);
and U5455 (N_5455,N_4032,N_764);
and U5456 (N_5456,N_698,N_2637);
nand U5457 (N_5457,N_2020,N_4137);
xor U5458 (N_5458,N_1349,N_2672);
nor U5459 (N_5459,N_288,N_1992);
or U5460 (N_5460,N_182,N_4489);
or U5461 (N_5461,N_4866,N_1131);
nor U5462 (N_5462,N_4372,N_4773);
nand U5463 (N_5463,N_278,N_1530);
nor U5464 (N_5464,N_625,N_113);
nand U5465 (N_5465,N_2744,N_4752);
and U5466 (N_5466,N_2076,N_1066);
xor U5467 (N_5467,N_813,N_4739);
nor U5468 (N_5468,N_366,N_3836);
nand U5469 (N_5469,N_153,N_2985);
and U5470 (N_5470,N_4686,N_4784);
or U5471 (N_5471,N_656,N_3398);
nor U5472 (N_5472,N_3799,N_1217);
nand U5473 (N_5473,N_3016,N_3324);
nor U5474 (N_5474,N_3544,N_2242);
nor U5475 (N_5475,N_1456,N_319);
nand U5476 (N_5476,N_2586,N_3303);
and U5477 (N_5477,N_3041,N_2966);
or U5478 (N_5478,N_2114,N_31);
and U5479 (N_5479,N_2538,N_2923);
nor U5480 (N_5480,N_3371,N_4650);
nor U5481 (N_5481,N_4336,N_1187);
and U5482 (N_5482,N_4522,N_1233);
xor U5483 (N_5483,N_122,N_3632);
nor U5484 (N_5484,N_4104,N_1444);
and U5485 (N_5485,N_2535,N_3468);
or U5486 (N_5486,N_481,N_2998);
and U5487 (N_5487,N_1847,N_4368);
and U5488 (N_5488,N_1330,N_3531);
nand U5489 (N_5489,N_2500,N_3549);
xor U5490 (N_5490,N_1674,N_4024);
xor U5491 (N_5491,N_3536,N_472);
nand U5492 (N_5492,N_3767,N_427);
and U5493 (N_5493,N_3552,N_3840);
and U5494 (N_5494,N_4161,N_455);
nor U5495 (N_5495,N_3821,N_735);
nand U5496 (N_5496,N_1272,N_2183);
and U5497 (N_5497,N_2318,N_2925);
or U5498 (N_5498,N_2517,N_2854);
xnor U5499 (N_5499,N_2600,N_3852);
nor U5500 (N_5500,N_4728,N_1128);
xor U5501 (N_5501,N_2930,N_2363);
nor U5502 (N_5502,N_3031,N_4171);
or U5503 (N_5503,N_60,N_2066);
nand U5504 (N_5504,N_1914,N_3048);
and U5505 (N_5505,N_3864,N_1333);
or U5506 (N_5506,N_4794,N_1320);
nor U5507 (N_5507,N_2702,N_2077);
nor U5508 (N_5508,N_2492,N_387);
nand U5509 (N_5509,N_2493,N_3044);
xor U5510 (N_5510,N_2422,N_4198);
xnor U5511 (N_5511,N_2873,N_2927);
and U5512 (N_5512,N_3256,N_3627);
nand U5513 (N_5513,N_1478,N_669);
nor U5514 (N_5514,N_2425,N_2956);
nor U5515 (N_5515,N_2969,N_3849);
and U5516 (N_5516,N_1969,N_3238);
nand U5517 (N_5517,N_1305,N_2111);
nand U5518 (N_5518,N_97,N_1833);
and U5519 (N_5519,N_4259,N_2807);
or U5520 (N_5520,N_4158,N_1533);
and U5521 (N_5521,N_2399,N_3281);
nor U5522 (N_5522,N_775,N_1952);
nand U5523 (N_5523,N_4814,N_4689);
nor U5524 (N_5524,N_4564,N_78);
nor U5525 (N_5525,N_2973,N_1490);
and U5526 (N_5526,N_2354,N_1879);
nand U5527 (N_5527,N_2806,N_4896);
nand U5528 (N_5528,N_2626,N_478);
or U5529 (N_5529,N_2764,N_231);
and U5530 (N_5530,N_1035,N_916);
nand U5531 (N_5531,N_4889,N_3184);
xnor U5532 (N_5532,N_3592,N_2835);
xnor U5533 (N_5533,N_2565,N_3143);
nand U5534 (N_5534,N_110,N_1481);
nor U5535 (N_5535,N_328,N_240);
or U5536 (N_5536,N_973,N_1263);
xnor U5537 (N_5537,N_1090,N_4394);
nand U5538 (N_5538,N_792,N_3535);
and U5539 (N_5539,N_3477,N_1214);
xnor U5540 (N_5540,N_79,N_2466);
and U5541 (N_5541,N_2340,N_1204);
nor U5542 (N_5542,N_4125,N_479);
and U5543 (N_5543,N_1985,N_4823);
nand U5544 (N_5544,N_333,N_2331);
nor U5545 (N_5545,N_1146,N_5);
or U5546 (N_5546,N_3266,N_1034);
nand U5547 (N_5547,N_556,N_867);
and U5548 (N_5548,N_862,N_1150);
nor U5549 (N_5549,N_1866,N_671);
nand U5550 (N_5550,N_2041,N_192);
nor U5551 (N_5551,N_4046,N_869);
nand U5552 (N_5552,N_2827,N_3651);
nand U5553 (N_5553,N_435,N_4619);
nand U5554 (N_5554,N_2617,N_982);
nor U5555 (N_5555,N_484,N_2344);
nor U5556 (N_5556,N_2660,N_4484);
nand U5557 (N_5557,N_3106,N_3195);
nor U5558 (N_5558,N_1098,N_3267);
or U5559 (N_5559,N_1794,N_4513);
or U5560 (N_5560,N_3737,N_2372);
nand U5561 (N_5561,N_1127,N_962);
xnor U5562 (N_5562,N_2129,N_541);
nor U5563 (N_5563,N_2169,N_2614);
nand U5564 (N_5564,N_4227,N_1949);
and U5565 (N_5565,N_3125,N_4254);
xnor U5566 (N_5566,N_3626,N_4375);
xnor U5567 (N_5567,N_1447,N_1040);
or U5568 (N_5568,N_1556,N_3709);
and U5569 (N_5569,N_371,N_2487);
nand U5570 (N_5570,N_322,N_815);
nand U5571 (N_5571,N_1373,N_508);
and U5572 (N_5572,N_1752,N_71);
or U5573 (N_5573,N_3483,N_452);
nand U5574 (N_5574,N_2276,N_104);
or U5575 (N_5575,N_3374,N_3);
nand U5576 (N_5576,N_3482,N_4843);
xnor U5577 (N_5577,N_778,N_4704);
nor U5578 (N_5578,N_695,N_4056);
nand U5579 (N_5579,N_2884,N_1982);
xor U5580 (N_5580,N_628,N_1697);
nor U5581 (N_5581,N_1571,N_4865);
nand U5582 (N_5582,N_4858,N_2068);
or U5583 (N_5583,N_722,N_3839);
nand U5584 (N_5584,N_2278,N_1497);
nor U5585 (N_5585,N_2324,N_73);
nand U5586 (N_5586,N_133,N_1666);
xor U5587 (N_5587,N_2320,N_4031);
or U5588 (N_5588,N_1739,N_1782);
xnor U5589 (N_5589,N_4875,N_186);
nand U5590 (N_5590,N_4512,N_1645);
xor U5591 (N_5591,N_1008,N_4192);
nor U5592 (N_5592,N_4312,N_1389);
nand U5593 (N_5593,N_4954,N_2330);
xor U5594 (N_5594,N_2864,N_4260);
nor U5595 (N_5595,N_684,N_4400);
or U5596 (N_5596,N_2788,N_315);
xor U5597 (N_5597,N_2478,N_2189);
or U5598 (N_5598,N_3380,N_3478);
nand U5599 (N_5599,N_2922,N_193);
nand U5600 (N_5600,N_805,N_4092);
or U5601 (N_5601,N_776,N_2063);
xor U5602 (N_5602,N_3545,N_4636);
or U5603 (N_5603,N_4891,N_95);
or U5604 (N_5604,N_2735,N_1551);
or U5605 (N_5605,N_4086,N_2463);
nand U5606 (N_5606,N_1032,N_3431);
nand U5607 (N_5607,N_4403,N_907);
or U5608 (N_5608,N_932,N_1348);
and U5609 (N_5609,N_68,N_16);
xnor U5610 (N_5610,N_4066,N_1249);
and U5611 (N_5611,N_4112,N_4661);
nand U5612 (N_5612,N_2866,N_4014);
xor U5613 (N_5613,N_4011,N_209);
and U5614 (N_5614,N_2642,N_4521);
xnor U5615 (N_5615,N_3502,N_659);
or U5616 (N_5616,N_3654,N_1191);
xor U5617 (N_5617,N_2397,N_342);
nand U5618 (N_5618,N_2468,N_1199);
and U5619 (N_5619,N_1719,N_515);
nand U5620 (N_5620,N_4607,N_717);
nand U5621 (N_5621,N_3402,N_3362);
xnor U5622 (N_5622,N_1513,N_4737);
nor U5623 (N_5623,N_1436,N_562);
xor U5624 (N_5624,N_1662,N_3516);
nand U5625 (N_5625,N_4469,N_777);
or U5626 (N_5626,N_128,N_1784);
nand U5627 (N_5627,N_1748,N_1365);
or U5628 (N_5628,N_254,N_1544);
or U5629 (N_5629,N_850,N_3826);
and U5630 (N_5630,N_3498,N_3049);
or U5631 (N_5631,N_2750,N_1643);
xnor U5632 (N_5632,N_716,N_3129);
nor U5633 (N_5633,N_314,N_877);
or U5634 (N_5634,N_4315,N_977);
or U5635 (N_5635,N_3313,N_457);
or U5636 (N_5636,N_2308,N_2624);
xnor U5637 (N_5637,N_1222,N_3134);
nand U5638 (N_5638,N_3879,N_560);
xor U5639 (N_5639,N_3642,N_1997);
xor U5640 (N_5640,N_2948,N_201);
nand U5641 (N_5641,N_441,N_4170);
or U5642 (N_5642,N_2846,N_3088);
or U5643 (N_5643,N_632,N_2392);
and U5644 (N_5644,N_4824,N_2725);
nand U5645 (N_5645,N_227,N_1770);
xor U5646 (N_5646,N_176,N_4912);
and U5647 (N_5647,N_1667,N_2381);
and U5648 (N_5648,N_2549,N_4174);
xor U5649 (N_5649,N_3532,N_2694);
and U5650 (N_5650,N_1559,N_4985);
nand U5651 (N_5651,N_4988,N_3892);
nand U5652 (N_5652,N_3848,N_1732);
and U5653 (N_5653,N_4595,N_3160);
or U5654 (N_5654,N_537,N_2405);
or U5655 (N_5655,N_2914,N_299);
nor U5656 (N_5656,N_997,N_497);
xor U5657 (N_5657,N_2082,N_3091);
nor U5658 (N_5658,N_4223,N_2230);
and U5659 (N_5659,N_3927,N_117);
and U5660 (N_5660,N_3055,N_2625);
xnor U5661 (N_5661,N_1300,N_563);
nand U5662 (N_5662,N_2419,N_2887);
xnor U5663 (N_5663,N_359,N_4558);
and U5664 (N_5664,N_2296,N_4997);
nand U5665 (N_5665,N_4119,N_498);
nand U5666 (N_5666,N_679,N_262);
xor U5667 (N_5667,N_2170,N_1203);
nand U5668 (N_5668,N_2635,N_4914);
or U5669 (N_5669,N_2653,N_3467);
nor U5670 (N_5670,N_2416,N_3857);
and U5671 (N_5671,N_1818,N_4109);
or U5672 (N_5672,N_2831,N_1718);
nor U5673 (N_5673,N_2699,N_1514);
xor U5674 (N_5674,N_2411,N_4621);
nand U5675 (N_5675,N_4765,N_4212);
xor U5676 (N_5676,N_2684,N_1246);
nand U5677 (N_5677,N_1004,N_4222);
nand U5678 (N_5678,N_3914,N_3470);
and U5679 (N_5679,N_734,N_3671);
and U5680 (N_5680,N_312,N_4234);
or U5681 (N_5681,N_402,N_3297);
or U5682 (N_5682,N_2747,N_2528);
xnor U5683 (N_5683,N_4733,N_1048);
nand U5684 (N_5684,N_1624,N_635);
nor U5685 (N_5685,N_4684,N_3051);
xor U5686 (N_5686,N_3784,N_2234);
nand U5687 (N_5687,N_4200,N_2823);
xor U5688 (N_5688,N_1457,N_1115);
and U5689 (N_5689,N_1764,N_1610);
xor U5690 (N_5690,N_3067,N_3617);
nor U5691 (N_5691,N_1535,N_1710);
or U5692 (N_5692,N_3464,N_3907);
nand U5693 (N_5693,N_2314,N_4520);
and U5694 (N_5694,N_1942,N_4496);
nand U5695 (N_5695,N_2227,N_704);
and U5696 (N_5696,N_4392,N_2679);
nor U5697 (N_5697,N_3279,N_1519);
and U5698 (N_5698,N_1713,N_2681);
and U5699 (N_5699,N_2412,N_2039);
nor U5700 (N_5700,N_1438,N_1772);
nand U5701 (N_5701,N_3584,N_4527);
xor U5702 (N_5702,N_4708,N_4574);
and U5703 (N_5703,N_2561,N_536);
xor U5704 (N_5704,N_2190,N_4864);
xor U5705 (N_5705,N_1270,N_3548);
and U5706 (N_5706,N_843,N_2138);
and U5707 (N_5707,N_3634,N_3309);
and U5708 (N_5708,N_956,N_2510);
or U5709 (N_5709,N_1407,N_2275);
nand U5710 (N_5710,N_2757,N_4569);
nand U5711 (N_5711,N_1137,N_896);
and U5712 (N_5712,N_4362,N_2004);
or U5713 (N_5713,N_846,N_1790);
or U5714 (N_5714,N_2470,N_2877);
and U5715 (N_5715,N_2898,N_630);
xor U5716 (N_5716,N_1111,N_2214);
xor U5717 (N_5717,N_4551,N_4927);
and U5718 (N_5718,N_2810,N_1686);
and U5719 (N_5719,N_741,N_1157);
xor U5720 (N_5720,N_4301,N_2267);
xnor U5721 (N_5721,N_4916,N_3673);
nor U5722 (N_5722,N_2467,N_2513);
and U5723 (N_5723,N_2187,N_4249);
and U5724 (N_5724,N_685,N_2453);
and U5725 (N_5725,N_3379,N_305);
or U5726 (N_5726,N_4913,N_3154);
nor U5727 (N_5727,N_425,N_3151);
and U5728 (N_5728,N_4734,N_4763);
nand U5729 (N_5729,N_3707,N_3062);
and U5730 (N_5730,N_981,N_306);
nor U5731 (N_5731,N_2174,N_1946);
nor U5732 (N_5732,N_796,N_2640);
nand U5733 (N_5733,N_1856,N_345);
xor U5734 (N_5734,N_4803,N_271);
xor U5735 (N_5735,N_276,N_4242);
or U5736 (N_5736,N_1367,N_1064);
nand U5737 (N_5737,N_2295,N_2633);
nand U5738 (N_5738,N_1680,N_824);
nand U5739 (N_5739,N_1284,N_203);
nand U5740 (N_5740,N_4507,N_3240);
nand U5741 (N_5741,N_424,N_822);
nor U5742 (N_5742,N_4348,N_3080);
nor U5743 (N_5743,N_1845,N_1340);
and U5744 (N_5744,N_1894,N_3694);
nand U5745 (N_5745,N_3081,N_4440);
and U5746 (N_5746,N_3542,N_211);
xnor U5747 (N_5747,N_803,N_507);
or U5748 (N_5748,N_1378,N_2634);
or U5749 (N_5749,N_4911,N_816);
nand U5750 (N_5750,N_2763,N_3424);
nor U5751 (N_5751,N_4529,N_1685);
nor U5752 (N_5752,N_4735,N_3411);
or U5753 (N_5753,N_1778,N_2668);
nor U5754 (N_5754,N_626,N_3037);
or U5755 (N_5755,N_185,N_2790);
nor U5756 (N_5756,N_2102,N_4550);
nor U5757 (N_5757,N_4671,N_2429);
nor U5758 (N_5758,N_2657,N_1380);
xnor U5759 (N_5759,N_94,N_4966);
nand U5760 (N_5760,N_462,N_1734);
and U5761 (N_5761,N_1043,N_1443);
nor U5762 (N_5762,N_2620,N_3958);
or U5763 (N_5763,N_4094,N_3200);
nor U5764 (N_5764,N_4992,N_751);
or U5765 (N_5765,N_341,N_3167);
and U5766 (N_5766,N_4639,N_3146);
or U5767 (N_5767,N_3459,N_3199);
nor U5768 (N_5768,N_4326,N_3609);
xor U5769 (N_5769,N_1049,N_2793);
nor U5770 (N_5770,N_3396,N_4518);
and U5771 (N_5771,N_2250,N_4338);
xor U5772 (N_5772,N_3557,N_370);
or U5773 (N_5773,N_2814,N_84);
and U5774 (N_5774,N_1162,N_2186);
nand U5775 (N_5775,N_217,N_149);
or U5776 (N_5776,N_2616,N_4949);
and U5777 (N_5777,N_3835,N_866);
nor U5778 (N_5778,N_1205,N_3400);
nand U5779 (N_5779,N_3985,N_3203);
and U5780 (N_5780,N_2247,N_1200);
nand U5781 (N_5781,N_1415,N_1650);
or U5782 (N_5782,N_1065,N_1987);
and U5783 (N_5783,N_2421,N_2875);
nor U5784 (N_5784,N_720,N_3202);
nor U5785 (N_5785,N_3808,N_2388);
nand U5786 (N_5786,N_4559,N_789);
and U5787 (N_5787,N_4651,N_3523);
nand U5788 (N_5788,N_951,N_1439);
xor U5789 (N_5789,N_3554,N_3357);
nor U5790 (N_5790,N_2683,N_2843);
or U5791 (N_5791,N_4793,N_1234);
xnor U5792 (N_5792,N_4601,N_4416);
nand U5793 (N_5793,N_277,N_1265);
or U5794 (N_5794,N_1493,N_4986);
xor U5795 (N_5795,N_1430,N_3299);
xnor U5796 (N_5796,N_785,N_3103);
nor U5797 (N_5797,N_4050,N_1798);
nand U5798 (N_5798,N_3035,N_2907);
nor U5799 (N_5799,N_1537,N_4376);
nand U5800 (N_5800,N_368,N_2341);
xor U5801 (N_5801,N_4233,N_232);
xnor U5802 (N_5802,N_4667,N_1001);
and U5803 (N_5803,N_730,N_1977);
or U5804 (N_5804,N_1072,N_950);
nor U5805 (N_5805,N_2917,N_2703);
nor U5806 (N_5806,N_1708,N_2815);
nor U5807 (N_5807,N_4682,N_2498);
xor U5808 (N_5808,N_4152,N_384);
and U5809 (N_5809,N_784,N_3599);
or U5810 (N_5810,N_2618,N_1375);
nand U5811 (N_5811,N_4645,N_2369);
or U5812 (N_5812,N_3001,N_0);
nor U5813 (N_5813,N_4079,N_3047);
nand U5814 (N_5814,N_568,N_904);
and U5815 (N_5815,N_1105,N_611);
nor U5816 (N_5816,N_3949,N_3722);
xnor U5817 (N_5817,N_400,N_2880);
nand U5818 (N_5818,N_1050,N_2562);
or U5819 (N_5819,N_3640,N_3986);
or U5820 (N_5820,N_1155,N_4849);
nor U5821 (N_5821,N_1181,N_1999);
or U5822 (N_5822,N_4418,N_3300);
nor U5823 (N_5823,N_2109,N_1298);
nor U5824 (N_5824,N_1036,N_1483);
xnor U5825 (N_5825,N_4806,N_1432);
nand U5826 (N_5826,N_594,N_2137);
or U5827 (N_5827,N_965,N_2560);
nor U5828 (N_5828,N_4727,N_2536);
xnor U5829 (N_5829,N_2305,N_1741);
and U5830 (N_5830,N_4721,N_4901);
xnor U5831 (N_5831,N_4754,N_3972);
or U5832 (N_5832,N_1165,N_4731);
xnor U5833 (N_5833,N_4990,N_112);
nor U5834 (N_5834,N_1931,N_2828);
nand U5835 (N_5835,N_4598,N_640);
or U5836 (N_5836,N_3394,N_428);
xor U5837 (N_5837,N_2541,N_4253);
nor U5838 (N_5838,N_175,N_4538);
nor U5839 (N_5839,N_2151,N_501);
nand U5840 (N_5840,N_1141,N_986);
nor U5841 (N_5841,N_2594,N_4264);
xnor U5842 (N_5842,N_3778,N_2177);
nor U5843 (N_5843,N_4245,N_2357);
nor U5844 (N_5844,N_4291,N_3597);
xnor U5845 (N_5845,N_1851,N_3633);
and U5846 (N_5846,N_1178,N_1858);
and U5847 (N_5847,N_4080,N_4055);
and U5848 (N_5848,N_921,N_2362);
nand U5849 (N_5849,N_762,N_1736);
and U5850 (N_5850,N_3658,N_4438);
xor U5851 (N_5851,N_4492,N_1291);
xor U5852 (N_5852,N_3113,N_1391);
nor U5853 (N_5853,N_1835,N_1927);
or U5854 (N_5854,N_3944,N_2717);
nand U5855 (N_5855,N_4844,N_2009);
nand U5856 (N_5856,N_4660,N_4097);
or U5857 (N_5857,N_4658,N_4579);
nor U5858 (N_5858,N_2906,N_199);
nor U5859 (N_5859,N_3692,N_374);
xnor U5860 (N_5860,N_4261,N_1783);
nor U5861 (N_5861,N_4855,N_4540);
nand U5862 (N_5862,N_1840,N_881);
or U5863 (N_5863,N_3824,N_3865);
xnor U5864 (N_5864,N_995,N_2046);
and U5865 (N_5865,N_4303,N_3255);
and U5866 (N_5866,N_2876,N_2055);
xor U5867 (N_5867,N_3842,N_1995);
nand U5868 (N_5868,N_2304,N_1805);
nor U5869 (N_5869,N_2371,N_1808);
xnor U5870 (N_5870,N_3819,N_1984);
nor U5871 (N_5871,N_2808,N_3263);
and U5872 (N_5872,N_2774,N_1392);
nor U5873 (N_5873,N_4421,N_4025);
and U5874 (N_5874,N_1009,N_2446);
or U5875 (N_5875,N_1442,N_4231);
xor U5876 (N_5876,N_1396,N_156);
xor U5877 (N_5877,N_2645,N_4075);
xor U5878 (N_5878,N_2460,N_2593);
and U5879 (N_5879,N_1896,N_4121);
xnor U5880 (N_5880,N_296,N_655);
or U5881 (N_5881,N_96,N_3570);
and U5882 (N_5882,N_2233,N_2002);
nor U5883 (N_5883,N_1280,N_3881);
and U5884 (N_5884,N_876,N_275);
and U5885 (N_5885,N_878,N_1882);
nand U5886 (N_5886,N_3429,N_4262);
or U5887 (N_5887,N_1062,N_2733);
or U5888 (N_5888,N_4385,N_3350);
nor U5889 (N_5889,N_3567,N_4130);
or U5890 (N_5890,N_2570,N_75);
and U5891 (N_5891,N_1838,N_2542);
or U5892 (N_5892,N_4387,N_918);
nand U5893 (N_5893,N_2720,N_1042);
xnor U5894 (N_5894,N_2779,N_3109);
or U5895 (N_5895,N_3677,N_1179);
nor U5896 (N_5896,N_1193,N_1113);
and U5897 (N_5897,N_1122,N_2979);
or U5898 (N_5898,N_2613,N_4532);
and U5899 (N_5899,N_4409,N_1900);
and U5900 (N_5900,N_2336,N_214);
or U5901 (N_5901,N_3514,N_3032);
nor U5902 (N_5902,N_316,N_395);
nand U5903 (N_5903,N_2805,N_585);
nor U5904 (N_5904,N_2274,N_3624);
xor U5905 (N_5905,N_4769,N_1558);
nand U5906 (N_5906,N_4475,N_4560);
and U5907 (N_5907,N_915,N_1797);
nand U5908 (N_5908,N_1370,N_766);
nand U5909 (N_5909,N_3880,N_2903);
nor U5910 (N_5910,N_3978,N_4625);
nor U5911 (N_5911,N_251,N_3244);
or U5912 (N_5912,N_32,N_3638);
or U5913 (N_5913,N_3042,N_4333);
xnor U5914 (N_5914,N_527,N_2662);
or U5915 (N_5915,N_2800,N_4828);
and U5916 (N_5916,N_731,N_1363);
nor U5917 (N_5917,N_672,N_3487);
or U5918 (N_5918,N_551,N_2133);
nor U5919 (N_5919,N_4827,N_3325);
nor U5920 (N_5920,N_4289,N_373);
xnor U5921 (N_5921,N_3335,N_1097);
xnor U5922 (N_5922,N_1347,N_454);
nor U5923 (N_5923,N_1117,N_290);
nand U5924 (N_5924,N_3234,N_1873);
nor U5925 (N_5925,N_2311,N_4554);
or U5926 (N_5926,N_1878,N_818);
xor U5927 (N_5927,N_303,N_1677);
or U5928 (N_5928,N_821,N_2858);
and U5929 (N_5929,N_3550,N_4777);
nor U5930 (N_5930,N_3672,N_2164);
nor U5931 (N_5931,N_1604,N_2551);
and U5932 (N_5932,N_1665,N_2994);
nand U5933 (N_5933,N_4054,N_889);
and U5934 (N_5934,N_3083,N_3247);
and U5935 (N_5935,N_3017,N_523);
or U5936 (N_5936,N_2059,N_4947);
and U5937 (N_5937,N_2014,N_1932);
xor U5938 (N_5938,N_1135,N_2479);
nor U5939 (N_5939,N_1281,N_2402);
or U5940 (N_5940,N_3229,N_1694);
and U5941 (N_5941,N_1007,N_3870);
and U5942 (N_5942,N_2167,N_4018);
and U5943 (N_5943,N_3383,N_1366);
or U5944 (N_5944,N_566,N_2939);
nor U5945 (N_5945,N_2967,N_1080);
and U5946 (N_5946,N_2582,N_3904);
nand U5947 (N_5947,N_3760,N_3003);
or U5948 (N_5948,N_1449,N_673);
or U5949 (N_5949,N_677,N_588);
xor U5950 (N_5950,N_4691,N_4202);
xnor U5951 (N_5951,N_4724,N_3311);
or U5952 (N_5952,N_2781,N_1153);
xor U5953 (N_5953,N_1753,N_3022);
nor U5954 (N_5954,N_1232,N_470);
nor U5955 (N_5955,N_3909,N_3757);
nand U5956 (N_5956,N_4009,N_1877);
xor U5957 (N_5957,N_155,N_3681);
and U5958 (N_5958,N_4330,N_3846);
or U5959 (N_5959,N_2890,N_4363);
or U5960 (N_5960,N_2339,N_172);
nor U5961 (N_5961,N_4962,N_909);
and U5962 (N_5962,N_2619,N_1869);
and U5963 (N_5963,N_20,N_1190);
nor U5964 (N_5964,N_3805,N_1011);
nor U5965 (N_5965,N_4929,N_3144);
nand U5966 (N_5966,N_1464,N_4602);
or U5967 (N_5967,N_4345,N_475);
nor U5968 (N_5968,N_4643,N_4834);
nor U5969 (N_5969,N_4467,N_1745);
or U5970 (N_5970,N_1166,N_469);
xor U5971 (N_5971,N_1622,N_1705);
xor U5972 (N_5972,N_2850,N_2152);
nor U5973 (N_5973,N_1534,N_4961);
xnor U5974 (N_5974,N_4090,N_945);
xnor U5975 (N_5975,N_624,N_1587);
and U5976 (N_5976,N_405,N_1565);
or U5977 (N_5977,N_3643,N_228);
and U5978 (N_5978,N_3170,N_3361);
or U5979 (N_5979,N_330,N_989);
and U5980 (N_5980,N_3059,N_4613);
and U5981 (N_5981,N_1312,N_3775);
nor U5982 (N_5982,N_4820,N_1195);
xnor U5983 (N_5983,N_4584,N_1428);
and U5984 (N_5984,N_4608,N_3509);
xor U5985 (N_5985,N_324,N_417);
nor U5986 (N_5986,N_4675,N_1459);
or U5987 (N_5987,N_795,N_1728);
nand U5988 (N_5988,N_1304,N_1411);
nor U5989 (N_5989,N_4196,N_2328);
or U5990 (N_5990,N_1174,N_1229);
or U5991 (N_5991,N_1470,N_3043);
and U5992 (N_5992,N_2548,N_2567);
nor U5993 (N_5993,N_343,N_1935);
and U5994 (N_5994,N_1779,N_320);
xnor U5995 (N_5995,N_2005,N_2708);
nand U5996 (N_5996,N_2726,N_4286);
and U5997 (N_5997,N_947,N_4199);
xor U5998 (N_5998,N_2494,N_474);
or U5999 (N_5999,N_2727,N_1950);
xor U6000 (N_6000,N_3655,N_1172);
or U6001 (N_6001,N_2530,N_2432);
or U6002 (N_6002,N_1440,N_3488);
nand U6003 (N_6003,N_2424,N_2785);
and U6004 (N_6004,N_4083,N_1938);
nand U6005 (N_6005,N_3173,N_1170);
or U6006 (N_6006,N_4666,N_376);
and U6007 (N_6007,N_1801,N_2598);
xor U6008 (N_6008,N_4269,N_4968);
nor U6009 (N_6009,N_4256,N_2057);
nor U6010 (N_6010,N_1455,N_3976);
or U6011 (N_6011,N_584,N_4833);
or U6012 (N_6012,N_4030,N_853);
nand U6013 (N_6013,N_1538,N_2832);
xnor U6014 (N_6014,N_3235,N_243);
or U6015 (N_6015,N_2885,N_2692);
or U6016 (N_6016,N_3330,N_3780);
and U6017 (N_6017,N_3222,N_344);
nand U6018 (N_6018,N_2307,N_2958);
nand U6019 (N_6019,N_292,N_4931);
and U6020 (N_6020,N_1126,N_468);
or U6021 (N_6021,N_4206,N_4447);
nor U6022 (N_6022,N_4576,N_3878);
nand U6023 (N_6023,N_4938,N_2773);
nor U6024 (N_6024,N_28,N_334);
and U6025 (N_6025,N_3551,N_3183);
or U6026 (N_6026,N_1671,N_961);
xnor U6027 (N_6027,N_4128,N_842);
and U6028 (N_6028,N_3327,N_1463);
nand U6029 (N_6029,N_1786,N_1635);
and U6030 (N_6030,N_1219,N_753);
and U6031 (N_6031,N_4881,N_2955);
or U6032 (N_6032,N_4604,N_3254);
and U6033 (N_6033,N_4606,N_2867);
nand U6034 (N_6034,N_3285,N_55);
xor U6035 (N_6035,N_2203,N_2612);
or U6036 (N_6036,N_3524,N_2952);
or U6037 (N_6037,N_119,N_4071);
or U6038 (N_6038,N_2863,N_1889);
nor U6039 (N_6039,N_3452,N_4466);
xnor U6040 (N_6040,N_3812,N_1499);
nor U6041 (N_6041,N_1104,N_294);
and U6042 (N_6042,N_2933,N_4051);
and U6043 (N_6043,N_3385,N_1083);
or U6044 (N_6044,N_1575,N_1188);
and U6045 (N_6045,N_4630,N_2124);
nor U6046 (N_6046,N_4812,N_4393);
and U6047 (N_6047,N_3420,N_2112);
nand U6048 (N_6048,N_3745,N_476);
and U6049 (N_6049,N_4015,N_4994);
xnor U6050 (N_6050,N_1917,N_2345);
nand U6051 (N_6051,N_139,N_3006);
or U6052 (N_6052,N_3210,N_3278);
and U6053 (N_6053,N_1372,N_3935);
nor U6054 (N_6054,N_2997,N_1789);
xnor U6055 (N_6055,N_3471,N_4549);
or U6056 (N_6056,N_2097,N_1248);
or U6057 (N_6057,N_162,N_794);
nand U6058 (N_6058,N_1522,N_4531);
or U6059 (N_6059,N_732,N_1875);
xnor U6060 (N_6060,N_3462,N_3122);
and U6061 (N_6061,N_3418,N_3902);
or U6062 (N_6062,N_3421,N_3967);
and U6063 (N_6063,N_100,N_3859);
and U6064 (N_6064,N_4582,N_3947);
nand U6065 (N_6065,N_3660,N_3970);
xor U6066 (N_6066,N_1920,N_3872);
xnor U6067 (N_6067,N_4043,N_1259);
nand U6068 (N_6068,N_2957,N_147);
and U6069 (N_6069,N_960,N_4908);
or U6070 (N_6070,N_1754,N_3093);
or U6071 (N_6071,N_4880,N_4151);
or U6072 (N_6072,N_1026,N_3368);
xnor U6073 (N_6073,N_3576,N_3720);
nor U6074 (N_6074,N_4971,N_4504);
and U6075 (N_6075,N_4377,N_2949);
or U6076 (N_6076,N_3399,N_464);
and U6077 (N_6077,N_2427,N_1966);
or U6078 (N_6078,N_4117,N_893);
nor U6079 (N_6079,N_3241,N_2691);
or U6080 (N_6080,N_4197,N_522);
or U6081 (N_6081,N_37,N_4327);
xor U6082 (N_6082,N_917,N_3020);
nand U6083 (N_6083,N_356,N_4503);
or U6084 (N_6084,N_2837,N_2280);
and U6085 (N_6085,N_2516,N_4244);
nand U6086 (N_6086,N_3971,N_3132);
xnor U6087 (N_6087,N_2355,N_2524);
and U6088 (N_6088,N_1915,N_1051);
and U6089 (N_6089,N_2366,N_406);
nand U6090 (N_6090,N_4930,N_2485);
and U6091 (N_6091,N_3803,N_1441);
xnor U6092 (N_6092,N_3656,N_759);
nor U6093 (N_6093,N_4611,N_1218);
xor U6094 (N_6094,N_420,N_703);
and U6095 (N_6095,N_1089,N_1316);
or U6096 (N_6096,N_4479,N_806);
xnor U6097 (N_6097,N_4700,N_1780);
nand U6098 (N_6098,N_3268,N_2053);
and U6099 (N_6099,N_3384,N_2091);
nand U6100 (N_6100,N_1374,N_1423);
xnor U6101 (N_6101,N_4785,N_1620);
or U6102 (N_6102,N_2584,N_3433);
xor U6103 (N_6103,N_645,N_2856);
and U6104 (N_6104,N_2812,N_2709);
xor U6105 (N_6105,N_65,N_727);
or U6106 (N_6106,N_696,N_3343);
nor U6107 (N_6107,N_3314,N_3329);
nand U6108 (N_6108,N_3525,N_3890);
and U6109 (N_6109,N_4314,N_4279);
or U6110 (N_6110,N_2268,N_942);
nor U6111 (N_6111,N_142,N_3435);
nand U6112 (N_6112,N_4519,N_4465);
or U6113 (N_6113,N_3097,N_1176);
xnor U6114 (N_6114,N_2648,N_4628);
xnor U6115 (N_6115,N_3193,N_205);
or U6116 (N_6116,N_3964,N_3393);
or U6117 (N_6117,N_3286,N_4852);
xor U6118 (N_6118,N_4185,N_2601);
and U6119 (N_6119,N_2166,N_2899);
nor U6120 (N_6120,N_3930,N_3975);
nand U6121 (N_6121,N_4305,N_1760);
nand U6122 (N_6122,N_1169,N_1769);
xor U6123 (N_6123,N_1746,N_4448);
nand U6124 (N_6124,N_1905,N_1);
nor U6125 (N_6125,N_3809,N_2865);
or U6126 (N_6126,N_3547,N_2678);
or U6127 (N_6127,N_1118,N_4168);
xnor U6128 (N_6128,N_3000,N_300);
nand U6129 (N_6129,N_854,N_4975);
and U6130 (N_6130,N_4498,N_3899);
or U6131 (N_6131,N_1427,N_2261);
or U6132 (N_6132,N_4358,N_459);
nand U6133 (N_6133,N_1771,N_3273);
xnor U6134 (N_6134,N_619,N_2881);
xor U6135 (N_6135,N_4339,N_4203);
or U6136 (N_6136,N_245,N_4328);
xnor U6137 (N_6137,N_1088,N_76);
xor U6138 (N_6138,N_807,N_4240);
xnor U6139 (N_6139,N_4404,N_2663);
and U6140 (N_6140,N_3069,N_2);
or U6141 (N_6141,N_129,N_4313);
and U6142 (N_6142,N_2313,N_21);
nand U6143 (N_6143,N_390,N_3591);
xnor U6144 (N_6144,N_4255,N_3159);
or U6145 (N_6145,N_3442,N_3717);
or U6146 (N_6146,N_4974,N_4624);
nor U6147 (N_6147,N_309,N_2627);
and U6148 (N_6148,N_800,N_3889);
nor U6149 (N_6149,N_409,N_559);
or U6150 (N_6150,N_4268,N_539);
and U6151 (N_6151,N_1037,N_3178);
or U6152 (N_6152,N_873,N_4786);
nor U6153 (N_6153,N_4353,N_89);
nand U6154 (N_6154,N_4743,N_2010);
nand U6155 (N_6155,N_1554,N_1108);
nor U6156 (N_6156,N_3137,N_2545);
and U6157 (N_6157,N_1567,N_3912);
and U6158 (N_6158,N_3119,N_3225);
nand U6159 (N_6159,N_3893,N_1381);
or U6160 (N_6160,N_2882,N_4087);
and U6161 (N_6161,N_3863,N_2021);
xor U6162 (N_6162,N_744,N_4714);
xnor U6163 (N_6163,N_3165,N_4502);
nand U6164 (N_6164,N_307,N_3779);
nand U6165 (N_6165,N_3201,N_545);
or U6166 (N_6166,N_1785,N_480);
xnor U6167 (N_6167,N_2801,N_2758);
xnor U6168 (N_6168,N_1434,N_987);
xor U6169 (N_6169,N_3213,N_2760);
and U6170 (N_6170,N_4237,N_2630);
and U6171 (N_6171,N_2855,N_4670);
nand U6172 (N_6172,N_3305,N_39);
and U6173 (N_6173,N_3226,N_2395);
xnor U6174 (N_6174,N_1849,N_974);
and U6175 (N_6175,N_4745,N_2080);
xnor U6176 (N_6176,N_386,N_1346);
xnor U6177 (N_6177,N_1182,N_4074);
nor U6178 (N_6178,N_3507,N_1161);
and U6179 (N_6179,N_1225,N_173);
xor U6180 (N_6180,N_3352,N_979);
and U6181 (N_6181,N_4488,N_4877);
nand U6182 (N_6182,N_3118,N_2802);
nand U6183 (N_6183,N_2629,N_3558);
nand U6184 (N_6184,N_4000,N_1531);
xor U6185 (N_6185,N_4213,N_1212);
or U6186 (N_6186,N_2537,N_2451);
nor U6187 (N_6187,N_3751,N_3341);
nor U6188 (N_6188,N_3344,N_4019);
and U6189 (N_6189,N_1235,N_2481);
or U6190 (N_6190,N_3636,N_1394);
or U6191 (N_6191,N_4306,N_2030);
or U6192 (N_6192,N_3372,N_2896);
xnor U6193 (N_6193,N_2581,N_4058);
nand U6194 (N_6194,N_3351,N_2217);
or U6195 (N_6195,N_4276,N_1403);
or U6196 (N_6196,N_3033,N_2822);
xnor U6197 (N_6197,N_3942,N_473);
nor U6198 (N_6198,N_167,N_3353);
nand U6199 (N_6199,N_3155,N_3058);
xnor U6200 (N_6200,N_2386,N_70);
nor U6201 (N_6201,N_514,N_4751);
and U6202 (N_6202,N_2142,N_1608);
and U6203 (N_6203,N_802,N_2905);
nor U6204 (N_6204,N_3804,N_4941);
nand U6205 (N_6205,N_3339,N_1761);
or U6206 (N_6206,N_1339,N_4139);
or U6207 (N_6207,N_3830,N_4135);
nand U6208 (N_6208,N_3427,N_2941);
and U6209 (N_6209,N_1454,N_4887);
xor U6210 (N_6210,N_2639,N_1484);
xnor U6211 (N_6211,N_4126,N_4232);
and U6212 (N_6212,N_811,N_2968);
and U6213 (N_6213,N_4557,N_1091);
nand U6214 (N_6214,N_2851,N_1816);
and U6215 (N_6215,N_4514,N_4444);
or U6216 (N_6216,N_574,N_1707);
nor U6217 (N_6217,N_40,N_647);
nand U6218 (N_6218,N_1020,N_1903);
xnor U6219 (N_6219,N_4842,N_1876);
nor U6220 (N_6220,N_3439,N_3659);
and U6221 (N_6221,N_1657,N_618);
nor U6222 (N_6222,N_4906,N_3426);
nand U6223 (N_6223,N_3443,N_2759);
nor U6224 (N_6224,N_4263,N_609);
nand U6225 (N_6225,N_3375,N_1189);
xor U6226 (N_6226,N_34,N_3098);
or U6227 (N_6227,N_4593,N_2654);
nand U6228 (N_6228,N_3845,N_1251);
xor U6229 (N_6229,N_3615,N_3843);
nand U6230 (N_6230,N_2292,N_3382);
nand U6231 (N_6231,N_702,N_4542);
or U6232 (N_6232,N_631,N_1465);
nand U6233 (N_6233,N_2291,N_587);
xnor U6234 (N_6234,N_4034,N_1154);
and U6235 (N_6235,N_4799,N_4340);
xnor U6236 (N_6236,N_2950,N_2576);
nor U6237 (N_6237,N_2532,N_1591);
and U6238 (N_6238,N_3215,N_1317);
and U6239 (N_6239,N_3166,N_1487);
nand U6240 (N_6240,N_2615,N_2965);
and U6241 (N_6241,N_4096,N_3714);
xor U6242 (N_6242,N_831,N_2458);
nand U6243 (N_6243,N_2373,N_1093);
nor U6244 (N_6244,N_2988,N_4021);
or U6245 (N_6245,N_2165,N_59);
or U6246 (N_6246,N_451,N_4944);
nand U6247 (N_6247,N_1880,N_1243);
nand U6248 (N_6248,N_3511,N_1078);
nor U6249 (N_6249,N_2786,N_1909);
nand U6250 (N_6250,N_2659,N_1024);
and U6251 (N_6251,N_577,N_1221);
or U6252 (N_6252,N_3716,N_488);
xor U6253 (N_6253,N_643,N_4154);
nor U6254 (N_6254,N_3569,N_198);
nor U6255 (N_6255,N_483,N_3124);
nor U6256 (N_6256,N_2723,N_1965);
and U6257 (N_6257,N_179,N_1972);
xor U6258 (N_6258,N_1405,N_1956);
xor U6259 (N_6259,N_4371,N_1461);
or U6260 (N_6260,N_670,N_3710);
nor U6261 (N_6261,N_3015,N_1580);
and U6262 (N_6262,N_622,N_1526);
nor U6263 (N_6263,N_3437,N_4101);
xnor U6264 (N_6264,N_150,N_2310);
and U6265 (N_6265,N_1945,N_1639);
xor U6266 (N_6266,N_3687,N_90);
nor U6267 (N_6267,N_197,N_3974);
and U6268 (N_6268,N_1264,N_7);
nand U6269 (N_6269,N_4397,N_3456);
and U6270 (N_6270,N_3490,N_1795);
or U6271 (N_6271,N_4759,N_3212);
nand U6272 (N_6272,N_1832,N_2798);
nand U6273 (N_6273,N_1045,N_3755);
or U6274 (N_6274,N_4082,N_817);
nor U6275 (N_6275,N_1827,N_711);
xor U6276 (N_6276,N_2281,N_3625);
and U6277 (N_6277,N_879,N_3715);
nand U6278 (N_6278,N_1107,N_1640);
or U6279 (N_6279,N_1369,N_3123);
nand U6280 (N_6280,N_1022,N_2001);
and U6281 (N_6281,N_3620,N_1557);
and U6282 (N_6282,N_1703,N_4698);
and U6283 (N_6283,N_4695,N_521);
nor U6284 (N_6284,N_4252,N_132);
nor U6285 (N_6285,N_3054,N_996);
nor U6286 (N_6286,N_3251,N_1775);
or U6287 (N_6287,N_2337,N_580);
and U6288 (N_6288,N_593,N_4585);
nand U6289 (N_6289,N_2049,N_238);
xnor U6290 (N_6290,N_14,N_3275);
and U6291 (N_6291,N_4568,N_1168);
xnor U6292 (N_6292,N_3217,N_3913);
nor U6293 (N_6293,N_4979,N_3894);
and U6294 (N_6294,N_2370,N_2193);
and U6295 (N_6295,N_1362,N_3472);
and U6296 (N_6296,N_4219,N_4167);
nor U6297 (N_6297,N_532,N_4720);
nor U6298 (N_6298,N_3198,N_4771);
or U6299 (N_6299,N_4516,N_3156);
nand U6300 (N_6300,N_769,N_2666);
or U6301 (N_6301,N_1302,N_3152);
or U6302 (N_6302,N_2821,N_3453);
nor U6303 (N_6303,N_3934,N_3274);
nor U6304 (N_6304,N_3395,N_4274);
nor U6305 (N_6305,N_2443,N_2438);
and U6306 (N_6306,N_1959,N_4406);
xnor U6307 (N_6307,N_934,N_189);
nand U6308 (N_6308,N_2849,N_2768);
and U6309 (N_6309,N_902,N_3121);
and U6310 (N_6310,N_4779,N_4188);
and U6311 (N_6311,N_1862,N_4894);
or U6312 (N_6312,N_3117,N_4829);
nor U6313 (N_6313,N_3602,N_1297);
and U6314 (N_6314,N_642,N_3494);
or U6315 (N_6315,N_2509,N_41);
nand U6316 (N_6316,N_2900,N_2783);
and U6317 (N_6317,N_4851,N_701);
xnor U6318 (N_6318,N_4981,N_2225);
nand U6319 (N_6319,N_2385,N_3232);
nand U6320 (N_6320,N_1082,N_4694);
nand U6321 (N_6321,N_136,N_1385);
nor U6322 (N_6322,N_4904,N_2871);
xnor U6323 (N_6323,N_2622,N_1201);
nand U6324 (N_6324,N_2732,N_4618);
xor U6325 (N_6325,N_273,N_3943);
nand U6326 (N_6326,N_1796,N_45);
and U6327 (N_6327,N_2434,N_3929);
nand U6328 (N_6328,N_11,N_1342);
or U6329 (N_6329,N_3764,N_3680);
xor U6330 (N_6330,N_2231,N_4723);
nor U6331 (N_6331,N_1254,N_2459);
and U6332 (N_6332,N_4265,N_658);
nand U6333 (N_6333,N_1310,N_3911);
nand U6334 (N_6334,N_4057,N_2609);
xor U6335 (N_6335,N_1968,N_1768);
and U6336 (N_6336,N_4594,N_2290);
nand U6337 (N_6337,N_3528,N_2266);
xor U6338 (N_6338,N_2597,N_2495);
xnor U6339 (N_6339,N_1612,N_3293);
or U6340 (N_6340,N_92,N_3679);
or U6341 (N_6341,N_210,N_583);
xor U6342 (N_6342,N_2972,N_351);
xnor U6343 (N_6343,N_4424,N_4899);
or U6344 (N_6344,N_3290,N_874);
xnor U6345 (N_6345,N_2442,N_2853);
nor U6346 (N_6346,N_1925,N_4552);
nand U6347 (N_6347,N_411,N_144);
nor U6348 (N_6348,N_116,N_1160);
nor U6349 (N_6349,N_2839,N_2931);
nor U6350 (N_6350,N_326,N_1301);
or U6351 (N_6351,N_4577,N_1585);
and U6352 (N_6352,N_604,N_3735);
nor U6353 (N_6353,N_990,N_2090);
xnor U6354 (N_6354,N_780,N_2590);
xnor U6355 (N_6355,N_4145,N_4108);
nor U6356 (N_6356,N_1542,N_3197);
xnor U6357 (N_6357,N_4882,N_605);
nand U6358 (N_6358,N_2534,N_4546);
and U6359 (N_6359,N_4048,N_3951);
xor U6360 (N_6360,N_2148,N_2156);
nor U6361 (N_6361,N_3264,N_4350);
nor U6362 (N_6362,N_1021,N_2346);
and U6363 (N_6363,N_3605,N_3231);
nand U6364 (N_6364,N_111,N_285);
and U6365 (N_6365,N_4487,N_652);
xor U6366 (N_6366,N_705,N_2029);
or U6367 (N_6367,N_4267,N_3414);
nor U6368 (N_6368,N_1597,N_13);
nor U6369 (N_6369,N_3610,N_3753);
xor U6370 (N_6370,N_3771,N_4186);
nand U6371 (N_6371,N_3082,N_2293);
nor U6372 (N_6372,N_4692,N_1295);
or U6373 (N_6373,N_852,N_2441);
xor U6374 (N_6374,N_2176,N_664);
or U6375 (N_6375,N_4464,N_287);
xnor U6376 (N_6376,N_2309,N_3665);
nor U6377 (N_6377,N_1837,N_3954);
or U6378 (N_6378,N_4838,N_2440);
or U6379 (N_6379,N_4505,N_403);
or U6380 (N_6380,N_2348,N_4283);
nor U6381 (N_6381,N_181,N_2926);
nand U6382 (N_6382,N_246,N_3242);
or U6383 (N_6383,N_2986,N_3527);
and U6384 (N_6384,N_4819,N_2697);
and U6385 (N_6385,N_4510,N_4335);
xnor U6386 (N_6386,N_4801,N_4884);
xnor U6387 (N_6387,N_1888,N_208);
and U6388 (N_6388,N_1029,N_4023);
and U6389 (N_6389,N_3513,N_4956);
nor U6390 (N_6390,N_2748,N_430);
and U6391 (N_6391,N_4429,N_1563);
nand U6392 (N_6392,N_3983,N_4243);
and U6393 (N_6393,N_4709,N_1562);
nand U6394 (N_6394,N_3461,N_4760);
xnor U6395 (N_6395,N_1913,N_4839);
nand U6396 (N_6396,N_4367,N_524);
nand U6397 (N_6397,N_1343,N_4523);
xor U6398 (N_6398,N_1729,N_939);
and U6399 (N_6399,N_461,N_3408);
or U6400 (N_6400,N_827,N_4907);
xnor U6401 (N_6401,N_955,N_561);
or U6402 (N_6402,N_3417,N_3973);
xnor U6403 (N_6403,N_2048,N_2316);
and U6404 (N_6404,N_1164,N_4217);
xor U6405 (N_6405,N_3559,N_742);
or U6406 (N_6406,N_2192,N_3952);
nand U6407 (N_6407,N_3588,N_798);
nor U6408 (N_6408,N_2216,N_1018);
xnor U6409 (N_6409,N_586,N_3189);
nand U6410 (N_6410,N_1588,N_3652);
xor U6411 (N_6411,N_797,N_3905);
nand U6412 (N_6412,N_1177,N_1676);
xor U6413 (N_6413,N_4614,N_2497);
xnor U6414 (N_6414,N_570,N_3564);
or U6415 (N_6415,N_1325,N_1807);
or U6416 (N_6416,N_3825,N_644);
xnor U6417 (N_6417,N_187,N_2650);
xor U6418 (N_6418,N_1252,N_8);
xnor U6419 (N_6419,N_540,N_2334);
nand U6420 (N_6420,N_3828,N_549);
xor U6421 (N_6421,N_2252,N_2820);
nand U6422 (N_6422,N_1152,N_844);
nand U6423 (N_6423,N_3661,N_4439);
nor U6424 (N_6424,N_3315,N_164);
nor U6425 (N_6425,N_674,N_2883);
or U6426 (N_6426,N_1475,N_2766);
xor U6427 (N_6427,N_1669,N_1929);
and U6428 (N_6428,N_4973,N_348);
or U6429 (N_6429,N_415,N_2991);
or U6430 (N_6430,N_2484,N_613);
or U6431 (N_6431,N_4717,N_244);
xor U6432 (N_6432,N_3877,N_1953);
nor U6433 (N_6433,N_728,N_1352);
xnor U6434 (N_6434,N_2263,N_1831);
or U6435 (N_6435,N_3724,N_3465);
xnor U6436 (N_6436,N_352,N_1864);
and U6437 (N_6437,N_2664,N_1701);
xor U6438 (N_6438,N_4457,N_4378);
xnor U6439 (N_6439,N_1255,N_1414);
nor U6440 (N_6440,N_2071,N_1656);
nand U6441 (N_6441,N_2701,N_2838);
xor U6442 (N_6442,N_3110,N_3485);
nor U6443 (N_6443,N_4616,N_1874);
nand U6444 (N_6444,N_985,N_636);
and U6445 (N_6445,N_346,N_4460);
and U6446 (N_6446,N_47,N_1960);
nor U6447 (N_6447,N_1285,N_4405);
and U6448 (N_6448,N_3053,N_4918);
nor U6449 (N_6449,N_35,N_3953);
and U6450 (N_6450,N_2974,N_2083);
nand U6451 (N_6451,N_648,N_1654);
nor U6452 (N_6452,N_1569,N_2942);
or U6453 (N_6453,N_4905,N_4647);
xor U6454 (N_6454,N_3820,N_1063);
xnor U6455 (N_6455,N_3938,N_3980);
or U6456 (N_6456,N_3338,N_2848);
nand U6457 (N_6457,N_2811,N_3711);
and U6458 (N_6458,N_3386,N_2945);
nand U6459 (N_6459,N_709,N_4459);
or U6460 (N_6460,N_1918,N_654);
xor U6461 (N_6461,N_592,N_2051);
xor U6462 (N_6462,N_3321,N_3246);
and U6463 (N_6463,N_4663,N_1578);
xnor U6464 (N_6464,N_3860,N_3162);
or U6465 (N_6465,N_161,N_3596);
xnor U6466 (N_6466,N_4308,N_1899);
nor U6467 (N_6467,N_1759,N_4040);
or U6468 (N_6468,N_1242,N_2317);
xnor U6469 (N_6469,N_1619,N_3856);
or U6470 (N_6470,N_3102,N_3519);
and U6471 (N_6471,N_4581,N_3706);
and U6472 (N_6472,N_3721,N_125);
xnor U6473 (N_6473,N_1971,N_1410);
and U6474 (N_6474,N_4972,N_4928);
xnor U6475 (N_6475,N_3770,N_3131);
nand U6476 (N_6476,N_4384,N_106);
and U6477 (N_6477,N_4790,N_268);
or U6478 (N_6478,N_4778,N_2000);
nor U6479 (N_6479,N_253,N_357);
and U6480 (N_6480,N_4100,N_1466);
or U6481 (N_6481,N_575,N_743);
or U6482 (N_6482,N_894,N_3333);
xnor U6483 (N_6483,N_3148,N_600);
or U6484 (N_6484,N_4134,N_446);
or U6485 (N_6485,N_4236,N_1327);
and U6486 (N_6486,N_130,N_2670);
and U6487 (N_6487,N_4180,N_3423);
nor U6488 (N_6488,N_3693,N_1910);
xnor U6489 (N_6489,N_2981,N_2064);
or U6490 (N_6490,N_3072,N_868);
and U6491 (N_6491,N_289,N_936);
xnor U6492 (N_6492,N_3066,N_2436);
nand U6493 (N_6493,N_3575,N_3446);
xnor U6494 (N_6494,N_3851,N_2257);
nand U6495 (N_6495,N_2254,N_2729);
or U6496 (N_6496,N_2248,N_1617);
and U6497 (N_6497,N_678,N_650);
nor U6498 (N_6498,N_2591,N_4878);
xnor U6499 (N_6499,N_274,N_4566);
nand U6500 (N_6500,N_1420,N_911);
xor U6501 (N_6501,N_38,N_3205);
nor U6502 (N_6502,N_2690,N_3901);
nor U6503 (N_6503,N_4932,N_4676);
and U6504 (N_6504,N_222,N_4204);
or U6505 (N_6505,N_774,N_4732);
nor U6506 (N_6506,N_2665,N_2978);
nor U6507 (N_6507,N_2572,N_3926);
nor U6508 (N_6508,N_99,N_2222);
or U6509 (N_6509,N_2445,N_1014);
nor U6510 (N_6510,N_3219,N_1706);
and U6511 (N_6511,N_148,N_1806);
xnor U6512 (N_6512,N_597,N_1991);
nand U6513 (N_6513,N_3791,N_2673);
nor U6514 (N_6514,N_2283,N_595);
or U6515 (N_6515,N_814,N_2845);
nand U6516 (N_6516,N_2749,N_4810);
nor U6517 (N_6517,N_2025,N_2126);
and U6518 (N_6518,N_1413,N_2557);
and U6519 (N_6519,N_1642,N_397);
and U6520 (N_6520,N_42,N_266);
nand U6521 (N_6521,N_3594,N_3518);
nand U6522 (N_6522,N_1336,N_528);
and U6523 (N_6523,N_4382,N_3932);
or U6524 (N_6524,N_4900,N_1244);
nor U6525 (N_6525,N_1962,N_3858);
and U6526 (N_6526,N_4478,N_2195);
or U6527 (N_6527,N_4285,N_2298);
nand U6528 (N_6528,N_3428,N_2651);
and U6529 (N_6529,N_526,N_2499);
nor U6530 (N_6530,N_10,N_3013);
nor U6531 (N_6531,N_3811,N_2238);
and U6532 (N_6532,N_4730,N_2202);
or U6533 (N_6533,N_190,N_830);
or U6534 (N_6534,N_505,N_2533);
or U6535 (N_6535,N_1121,N_3135);
and U6536 (N_6536,N_1125,N_426);
or U6537 (N_6537,N_418,N_589);
and U6538 (N_6538,N_264,N_4287);
xnor U6539 (N_6539,N_3139,N_3992);
or U6540 (N_6540,N_2809,N_143);
and U6541 (N_6541,N_4664,N_4797);
nand U6542 (N_6542,N_4346,N_1452);
nor U6543 (N_6543,N_4102,N_4792);
or U6544 (N_6544,N_1472,N_4788);
xnor U6545 (N_6545,N_3910,N_3331);
and U6546 (N_6546,N_4848,N_3795);
nand U6547 (N_6547,N_4225,N_4072);
nor U6548 (N_6548,N_4637,N_1476);
and U6549 (N_6549,N_4795,N_4561);
and U6550 (N_6550,N_4525,N_1081);
xor U6551 (N_6551,N_2448,N_1332);
and U6552 (N_6552,N_836,N_3489);
nor U6553 (N_6553,N_926,N_213);
nand U6554 (N_6554,N_3999,N_3369);
and U6555 (N_6555,N_2093,N_790);
or U6556 (N_6556,N_1670,N_3695);
and U6557 (N_6557,N_2042,N_3356);
nand U6558 (N_6558,N_4422,N_4247);
or U6559 (N_6559,N_548,N_377);
and U6560 (N_6560,N_4220,N_518);
nand U6561 (N_6561,N_302,N_4251);
nor U6562 (N_6562,N_3185,N_1815);
or U6563 (N_6563,N_2475,N_2817);
and U6564 (N_6564,N_1477,N_3114);
xnor U6565 (N_6565,N_4085,N_4370);
nand U6566 (N_6566,N_394,N_1151);
xnor U6567 (N_6567,N_3168,N_2408);
and U6568 (N_6568,N_3444,N_2437);
nor U6569 (N_6569,N_4407,N_4996);
or U6570 (N_6570,N_4044,N_4874);
xor U6571 (N_6571,N_4809,N_1981);
nor U6572 (N_6572,N_4910,N_2361);
xor U6573 (N_6573,N_2224,N_2104);
nor U6574 (N_6574,N_4853,N_1883);
or U6575 (N_6575,N_3568,N_1501);
xor U6576 (N_6576,N_4713,N_2204);
or U6577 (N_6577,N_183,N_2208);
xor U6578 (N_6578,N_311,N_1338);
xnor U6579 (N_6579,N_920,N_206);
nand U6580 (N_6580,N_2127,N_2990);
nor U6581 (N_6581,N_4863,N_3920);
nor U6582 (N_6582,N_1980,N_4587);
xor U6583 (N_6583,N_3334,N_621);
nor U6584 (N_6584,N_2426,N_1842);
or U6585 (N_6585,N_2862,N_3291);
nand U6586 (N_6586,N_925,N_4758);
and U6587 (N_6587,N_3153,N_4544);
nand U6588 (N_6588,N_3649,N_267);
nor U6589 (N_6589,N_1653,N_3412);
nand U6590 (N_6590,N_2035,N_3988);
and U6591 (N_6591,N_4084,N_140);
or U6592 (N_6592,N_3046,N_4169);
or U6593 (N_6593,N_4284,N_838);
xor U6594 (N_6594,N_3318,N_2132);
nand U6595 (N_6595,N_1192,N_3806);
nand U6596 (N_6596,N_4683,N_4860);
nor U6597 (N_6597,N_2704,N_382);
nor U6598 (N_6598,N_1749,N_1473);
and U6599 (N_6599,N_1085,N_2105);
nand U6600 (N_6600,N_739,N_726);
nor U6601 (N_6601,N_1354,N_2430);
or U6602 (N_6602,N_1068,N_241);
nor U6603 (N_6603,N_369,N_2098);
or U6604 (N_6604,N_499,N_1975);
xnor U6605 (N_6605,N_2611,N_4998);
xor U6606 (N_6606,N_3078,N_1149);
and U6607 (N_6607,N_3540,N_4895);
nand U6608 (N_6608,N_3060,N_4113);
xor U6609 (N_6609,N_3104,N_4374);
xor U6610 (N_6610,N_4934,N_4410);
or U6611 (N_6611,N_4774,N_1726);
nor U6612 (N_6612,N_1308,N_2461);
nand U6613 (N_6613,N_404,N_4357);
nor U6614 (N_6614,N_665,N_4832);
and U6615 (N_6615,N_91,N_2435);
and U6616 (N_6616,N_3747,N_3818);
xnor U6617 (N_6617,N_615,N_4662);
and U6618 (N_6618,N_4925,N_4716);
or U6619 (N_6619,N_971,N_1431);
and U6620 (N_6620,N_4445,N_1508);
nand U6621 (N_6621,N_1379,N_3875);
or U6622 (N_6622,N_4813,N_1054);
nand U6623 (N_6623,N_3211,N_3815);
or U6624 (N_6624,N_4299,N_234);
xnor U6625 (N_6625,N_3936,N_4536);
or U6626 (N_6626,N_4747,N_3298);
nand U6627 (N_6627,N_137,N_3292);
or U6628 (N_6628,N_3761,N_242);
and U6629 (N_6629,N_1171,N_81);
nor U6630 (N_6630,N_2546,N_1400);
and U6631 (N_6631,N_3797,N_1958);
xor U6632 (N_6632,N_3455,N_2730);
or U6633 (N_6633,N_3765,N_1468);
nand U6634 (N_6634,N_4037,N_2715);
and U6635 (N_6635,N_4187,N_2501);
nand U6636 (N_6636,N_1649,N_4991);
xnor U6637 (N_6637,N_4282,N_3434);
nor U6638 (N_6638,N_2312,N_1025);
nor U6639 (N_6639,N_2125,N_614);
or U6640 (N_6640,N_2403,N_1377);
xnor U6641 (N_6641,N_4110,N_3607);
nand U6642 (N_6642,N_383,N_1356);
and U6643 (N_6643,N_485,N_4693);
and U6644 (N_6644,N_1800,N_4028);
nand U6645 (N_6645,N_2196,N_4088);
and U6646 (N_6646,N_938,N_1926);
nor U6647 (N_6647,N_4868,N_4696);
xor U6648 (N_6648,N_3138,N_1142);
nand U6649 (N_6649,N_4257,N_3618);
or U6650 (N_6650,N_1351,N_4712);
nand U6651 (N_6651,N_1550,N_1867);
or U6652 (N_6652,N_216,N_1055);
nor U6653 (N_6653,N_4946,N_2667);
xor U6654 (N_6654,N_1636,N_856);
or U6655 (N_6655,N_906,N_3111);
nand U6656 (N_6656,N_496,N_3387);
or U6657 (N_6657,N_4845,N_2777);
nand U6658 (N_6658,N_707,N_1279);
or U6659 (N_6659,N_2338,N_4740);
and U6660 (N_6660,N_4105,N_3685);
nand U6661 (N_6661,N_1854,N_146);
nor U6662 (N_6662,N_4610,N_2599);
and U6663 (N_6663,N_2762,N_1103);
nand U6664 (N_6664,N_3019,N_2573);
or U6665 (N_6665,N_3713,N_1750);
and U6666 (N_6666,N_3562,N_2031);
nor U6667 (N_6667,N_2503,N_969);
nor U6668 (N_6668,N_2841,N_3571);
xor U6669 (N_6669,N_1902,N_4310);
nor U6670 (N_6670,N_2569,N_4600);
nand U6671 (N_6671,N_4679,N_1714);
or U6672 (N_6672,N_697,N_1973);
or U6673 (N_6673,N_2976,N_3187);
or U6674 (N_6674,N_49,N_3786);
or U6675 (N_6675,N_3758,N_3438);
nor U6676 (N_6676,N_3409,N_4474);
nand U6677 (N_6677,N_885,N_3036);
and U6678 (N_6678,N_2960,N_134);
nand U6679 (N_6679,N_2253,N_4854);
or U6680 (N_6680,N_450,N_3249);
nand U6681 (N_6681,N_3191,N_1206);
and U6682 (N_6682,N_1690,N_2181);
and U6683 (N_6683,N_1774,N_215);
xnor U6684 (N_6684,N_1307,N_421);
nor U6685 (N_6685,N_2518,N_3127);
or U6686 (N_6686,N_2789,N_295);
nand U6687 (N_6687,N_3796,N_4122);
nor U6688 (N_6688,N_4239,N_1641);
xnor U6689 (N_6689,N_3403,N_3390);
nor U6690 (N_6690,N_358,N_4939);
nor U6691 (N_6691,N_1185,N_2121);
nor U6692 (N_6692,N_4003,N_4380);
and U6693 (N_6693,N_651,N_1810);
nand U6694 (N_6694,N_3529,N_3521);
and U6695 (N_6695,N_3271,N_3419);
xnor U6696 (N_6696,N_740,N_3959);
or U6697 (N_6697,N_257,N_169);
nor U6698 (N_6698,N_2389,N_1607);
nand U6699 (N_6699,N_3908,N_1412);
nand U6700 (N_6700,N_308,N_2621);
nor U6701 (N_6701,N_4718,N_4456);
nand U6702 (N_6702,N_3814,N_691);
or U6703 (N_6703,N_3772,N_4053);
nor U6704 (N_6704,N_4069,N_1033);
xor U6705 (N_6705,N_2529,N_1777);
xor U6706 (N_6706,N_4383,N_3508);
and U6707 (N_6707,N_1978,N_993);
and U6708 (N_6708,N_4623,N_3176);
and U6709 (N_6709,N_3600,N_736);
nor U6710 (N_6710,N_2027,N_4609);
or U6711 (N_6711,N_2119,N_2236);
or U6712 (N_6712,N_2842,N_2473);
and U6713 (N_6713,N_279,N_2652);
and U6714 (N_6714,N_1625,N_2282);
nor U6715 (N_6715,N_1361,N_639);
and U6716 (N_6716,N_2943,N_2834);
nand U6717 (N_6717,N_3608,N_2780);
nor U6718 (N_6718,N_1445,N_4553);
nor U6719 (N_6719,N_2058,N_1529);
nor U6720 (N_6720,N_82,N_1616);
or U6721 (N_6721,N_3065,N_1884);
nand U6722 (N_6722,N_4680,N_1683);
nor U6723 (N_6723,N_310,N_4688);
or U6724 (N_6724,N_3406,N_596);
nand U6725 (N_6725,N_4064,N_1071);
xnor U6726 (N_6726,N_2205,N_3463);
or U6727 (N_6727,N_1294,N_2139);
or U6728 (N_6728,N_2394,N_1951);
or U6729 (N_6729,N_927,N_2013);
xnor U6730 (N_6730,N_44,N_414);
or U6731 (N_6731,N_4155,N_749);
nand U6732 (N_6732,N_2696,N_1819);
nor U6733 (N_6733,N_1853,N_1898);
xnor U6734 (N_6734,N_381,N_364);
and U6735 (N_6735,N_1143,N_2531);
nor U6736 (N_6736,N_799,N_2587);
or U6737 (N_6737,N_1830,N_1799);
nor U6738 (N_6738,N_2211,N_2277);
nor U6739 (N_6739,N_924,N_3736);
nand U6740 (N_6740,N_4605,N_72);
and U6741 (N_6741,N_4226,N_4238);
or U6742 (N_6742,N_2404,N_3007);
or U6743 (N_6743,N_4321,N_1687);
nor U6744 (N_6744,N_3664,N_1568);
and U6745 (N_6745,N_4746,N_1970);
and U6746 (N_6746,N_700,N_261);
nor U6747 (N_6747,N_2819,N_3900);
xnor U6748 (N_6748,N_4189,N_1371);
xnor U6749 (N_6749,N_2329,N_1110);
nand U6750 (N_6750,N_841,N_3924);
nor U6751 (N_6751,N_4649,N_336);
or U6752 (N_6752,N_738,N_4193);
and U6753 (N_6753,N_423,N_3956);
and U6754 (N_6754,N_2574,N_2450);
or U6755 (N_6755,N_2096,N_2103);
nor U6756 (N_6756,N_1988,N_2647);
and U6757 (N_6757,N_4162,N_2379);
xor U6758 (N_6758,N_2813,N_2836);
nand U6759 (N_6759,N_3646,N_220);
nand U6760 (N_6760,N_2128,N_4677);
nand U6761 (N_6761,N_2962,N_733);
or U6762 (N_6762,N_3984,N_3841);
nand U6763 (N_6763,N_3776,N_4452);
nor U6764 (N_6764,N_2583,N_4191);
xor U6765 (N_6765,N_2932,N_686);
or U6766 (N_6766,N_3340,N_4580);
and U6767 (N_6767,N_2163,N_991);
nor U6768 (N_6768,N_1885,N_829);
nor U6769 (N_6769,N_2118,N_2753);
and U6770 (N_6770,N_2131,N_2671);
nand U6771 (N_6771,N_3370,N_4655);
and U6772 (N_6772,N_1402,N_865);
nor U6773 (N_6773,N_1047,N_4622);
nor U6774 (N_6774,N_4293,N_1692);
and U6775 (N_6775,N_1073,N_4275);
and U6776 (N_6776,N_4138,N_2508);
nand U6777 (N_6777,N_3296,N_3701);
and U6778 (N_6778,N_1740,N_2539);
xnor U6779 (N_6779,N_4674,N_3416);
xnor U6780 (N_6780,N_4399,N_3209);
nor U6781 (N_6781,N_2769,N_2511);
xor U6782 (N_6782,N_439,N_4493);
or U6783 (N_6783,N_3731,N_1267);
nand U6784 (N_6784,N_4324,N_1939);
xnor U6785 (N_6785,N_4390,N_4455);
and U6786 (N_6786,N_4166,N_3702);
nor U6787 (N_6787,N_1834,N_4136);
xor U6788 (N_6788,N_4098,N_1100);
nand U6789 (N_6789,N_3573,N_2377);
nand U6790 (N_6790,N_4472,N_1114);
or U6791 (N_6791,N_2860,N_2321);
nor U6792 (N_6792,N_1954,N_4062);
and U6793 (N_6793,N_1266,N_4007);
nand U6794 (N_6794,N_3635,N_2390);
or U6795 (N_6795,N_1747,N_1865);
nand U6796 (N_6796,N_4369,N_46);
nor U6797 (N_6797,N_223,N_4364);
and U6798 (N_6798,N_1904,N_3214);
xnor U6799 (N_6799,N_3307,N_928);
nand U6800 (N_6800,N_1647,N_3023);
or U6801 (N_6801,N_67,N_429);
or U6802 (N_6802,N_2490,N_165);
nand U6803 (N_6803,N_3064,N_145);
nand U6804 (N_6804,N_486,N_4922);
xnor U6805 (N_6805,N_954,N_1006);
and U6806 (N_6806,N_1689,N_598);
xnor U6807 (N_6807,N_2393,N_2378);
and U6808 (N_6808,N_1238,N_2188);
xor U6809 (N_6809,N_3364,N_4277);
nor U6810 (N_6810,N_2989,N_2816);
nor U6811 (N_6811,N_692,N_2934);
xor U6812 (N_6812,N_3175,N_2024);
nor U6813 (N_6813,N_4334,N_1326);
and U6814 (N_6814,N_782,N_1897);
xnor U6815 (N_6815,N_1287,N_4804);
and U6816 (N_6816,N_2089,N_3301);
or U6817 (N_6817,N_4081,N_2387);
and U6818 (N_6818,N_1733,N_4876);
and U6819 (N_6819,N_4715,N_3140);
nor U6820 (N_6820,N_3440,N_3553);
nand U6821 (N_6821,N_2383,N_4653);
and U6822 (N_6822,N_2913,N_204);
nor U6823 (N_6823,N_4969,N_3798);
nor U6824 (N_6824,N_4360,N_2079);
xor U6825 (N_6825,N_1429,N_1239);
and U6826 (N_6826,N_3886,N_2588);
nand U6827 (N_6827,N_4356,N_4808);
or U6828 (N_6828,N_3738,N_1186);
xnor U6829 (N_6829,N_1730,N_2255);
and U6830 (N_6830,N_948,N_2507);
and U6831 (N_6831,N_1419,N_171);
nor U6832 (N_6832,N_1528,N_504);
and U6833 (N_6833,N_715,N_9);
and U6834 (N_6834,N_791,N_3040);
nand U6835 (N_6835,N_1688,N_4146);
nor U6836 (N_6836,N_3376,N_3145);
xor U6837 (N_6837,N_657,N_3497);
nor U6838 (N_6838,N_1341,N_2062);
or U6839 (N_6839,N_967,N_226);
or U6840 (N_6840,N_3948,N_4311);
or U6841 (N_6841,N_3657,N_325);
or U6842 (N_6842,N_3323,N_4355);
and U6843 (N_6843,N_2929,N_3749);
or U6844 (N_6844,N_1318,N_2741);
or U6845 (N_6845,N_2375,N_2578);
or U6846 (N_6846,N_984,N_353);
nor U6847 (N_6847,N_1309,N_2286);
or U6848 (N_6848,N_1451,N_864);
nor U6849 (N_6849,N_2326,N_910);
xor U6850 (N_6850,N_746,N_1994);
nand U6851 (N_6851,N_3794,N_2674);
nand U6852 (N_6852,N_4133,N_2171);
or U6853 (N_6853,N_4690,N_247);
or U6854 (N_6854,N_3450,N_4830);
or U6855 (N_6855,N_2607,N_248);
or U6856 (N_6856,N_4586,N_931);
nand U6857 (N_6857,N_3026,N_338);
or U6858 (N_6858,N_1776,N_2219);
and U6859 (N_6859,N_4008,N_2146);
nor U6860 (N_6860,N_1623,N_1505);
nand U6861 (N_6861,N_1817,N_1684);
or U6862 (N_6862,N_4159,N_2852);
and U6863 (N_6863,N_725,N_2754);
nor U6864 (N_6864,N_4388,N_4936);
and U6865 (N_6865,N_4352,N_4201);
nor U6866 (N_6866,N_3895,N_442);
nand U6867 (N_6867,N_4184,N_3696);
and U6868 (N_6868,N_1886,N_477);
nor U6869 (N_6869,N_3968,N_668);
nor U6870 (N_6870,N_431,N_396);
xnor U6871 (N_6871,N_1028,N_207);
nand U6872 (N_6872,N_2342,N_2649);
nand U6873 (N_6873,N_2368,N_4499);
nand U6874 (N_6874,N_4320,N_1323);
and U6875 (N_6875,N_2085,N_2069);
xor U6876 (N_6876,N_3565,N_4230);
or U6877 (N_6877,N_4132,N_2285);
nand U6878 (N_6878,N_467,N_4500);
or U6879 (N_6879,N_3933,N_3595);
or U6880 (N_6880,N_2721,N_438);
nor U6881 (N_6881,N_4298,N_249);
nor U6882 (N_6882,N_1727,N_2409);
and U6883 (N_6883,N_1075,N_880);
xor U6884 (N_6884,N_2686,N_2075);
or U6885 (N_6885,N_534,N_2472);
nor U6886 (N_6886,N_2471,N_157);
and U6887 (N_6887,N_1663,N_4107);
xor U6888 (N_6888,N_2123,N_2229);
xor U6889 (N_6889,N_4725,N_1268);
nand U6890 (N_6890,N_529,N_1802);
or U6891 (N_6891,N_4386,N_4648);
xor U6892 (N_6892,N_69,N_2018);
and U6893 (N_6893,N_557,N_3705);
nor U6894 (N_6894,N_4144,N_4533);
and U6895 (N_6895,N_4837,N_4657);
or U6896 (N_6896,N_212,N_1335);
xnor U6897 (N_6897,N_1859,N_4248);
nand U6898 (N_6898,N_937,N_1912);
or U6899 (N_6899,N_2410,N_282);
and U6900 (N_6900,N_3768,N_1947);
nor U6901 (N_6901,N_3171,N_1523);
xor U6902 (N_6902,N_543,N_291);
nor U6903 (N_6903,N_219,N_399);
xor U6904 (N_6904,N_3493,N_2241);
or U6905 (N_6905,N_3580,N_4856);
xor U6906 (N_6906,N_3317,N_4871);
nor U6907 (N_6907,N_2824,N_4528);
nor U6908 (N_6908,N_3667,N_3250);
or U6909 (N_6909,N_2902,N_3853);
or U6910 (N_6910,N_2547,N_4547);
nor U6911 (N_6911,N_437,N_449);
and U6912 (N_6912,N_2689,N_4273);
and U6913 (N_6913,N_1974,N_4045);
or U6914 (N_6914,N_1230,N_3095);
or U6915 (N_6915,N_126,N_3276);
nand U6916 (N_6916,N_637,N_1712);
xnor U6917 (N_6917,N_3639,N_2220);
and U6918 (N_6918,N_3725,N_3585);
xnor U6919 (N_6919,N_121,N_1924);
or U6920 (N_6920,N_3221,N_3774);
and U6921 (N_6921,N_1387,N_4530);
nor U6922 (N_6922,N_1681,N_4659);
nand U6923 (N_6923,N_2784,N_1633);
and U6924 (N_6924,N_4099,N_4342);
xor U6925 (N_6925,N_2092,N_33);
or U6926 (N_6926,N_2374,N_4920);
xor U6927 (N_6927,N_1820,N_3404);
nand U6928 (N_6928,N_520,N_2714);
nand U6929 (N_6929,N_1803,N_1276);
nor U6930 (N_6930,N_1787,N_1144);
or U6931 (N_6931,N_3366,N_1934);
nor U6932 (N_6932,N_755,N_4835);
nor U6933 (N_6933,N_4373,N_2240);
xor U6934 (N_6934,N_4449,N_4483);
xnor U6935 (N_6935,N_3586,N_4570);
nor U6936 (N_6936,N_1566,N_3703);
nor U6937 (N_6937,N_1183,N_3891);
and U6938 (N_6938,N_4296,N_2352);
or U6939 (N_6939,N_1494,N_4235);
xor U6940 (N_6940,N_3316,N_4902);
nand U6941 (N_6941,N_3698,N_2380);
nand U6942 (N_6942,N_718,N_2343);
nor U6943 (N_6943,N_2928,N_3094);
and U6944 (N_6944,N_3436,N_327);
nor U6945 (N_6945,N_772,N_419);
and U6946 (N_6946,N_3918,N_4029);
xor U6947 (N_6947,N_2384,N_2028);
and U6948 (N_6948,N_57,N_1220);
nor U6949 (N_6949,N_3623,N_4006);
nor U6950 (N_6950,N_2012,N_2868);
nor U6951 (N_6951,N_2215,N_3190);
xnor U6952 (N_6952,N_3005,N_4022);
and U6953 (N_6953,N_2521,N_3637);
xnor U6954 (N_6954,N_3697,N_1893);
xor U6955 (N_6955,N_4476,N_3834);
or U6956 (N_6956,N_1213,N_3336);
or U6957 (N_6957,N_2916,N_1561);
nor U6958 (N_6958,N_4142,N_3977);
nand U6959 (N_6959,N_500,N_4951);
nand U6960 (N_6960,N_2423,N_1572);
nor U6961 (N_6961,N_3993,N_1937);
nand U6962 (N_6962,N_2175,N_3823);
and U6963 (N_6963,N_443,N_1809);
or U6964 (N_6964,N_4744,N_1474);
nor U6965 (N_6965,N_2141,N_3074);
nand U6966 (N_6966,N_4052,N_2870);
nor U6967 (N_6967,N_601,N_2444);
and U6968 (N_6968,N_1480,N_634);
nand U6969 (N_6969,N_2251,N_1023);
xor U6970 (N_6970,N_2153,N_826);
xnor U6971 (N_6971,N_2050,N_1467);
or U6972 (N_6972,N_2107,N_2579);
and U6973 (N_6973,N_1621,N_2198);
or U6974 (N_6974,N_2504,N_1659);
and U6975 (N_6975,N_4535,N_4796);
xor U6976 (N_6976,N_4697,N_2975);
or U6977 (N_6977,N_2476,N_3018);
nor U6978 (N_6978,N_4926,N_4341);
nor U6979 (N_6979,N_3684,N_3925);
nor U6980 (N_6980,N_2136,N_3295);
nor U6981 (N_6981,N_1993,N_3010);
or U6982 (N_6982,N_4539,N_2015);
or U6983 (N_6983,N_1507,N_781);
or U6984 (N_6984,N_3987,N_1120);
and U6985 (N_6985,N_2770,N_3783);
xor U6986 (N_6986,N_3289,N_375);
nor U6987 (N_6987,N_2496,N_3937);
nor U6988 (N_6988,N_2199,N_1489);
xor U6989 (N_6989,N_1019,N_202);
nor U6990 (N_6990,N_1577,N_4898);
nor U6991 (N_6991,N_4175,N_3619);
and U6992 (N_6992,N_3034,N_900);
or U6993 (N_6993,N_988,N_1967);
xnor U6994 (N_6994,N_1606,N_3691);
or U6995 (N_6995,N_4118,N_380);
and U6996 (N_6996,N_666,N_2857);
xnor U6997 (N_6997,N_1207,N_3539);
nand U6998 (N_6998,N_3866,N_2117);
and U6999 (N_6999,N_1360,N_2455);
nand U7000 (N_7000,N_1979,N_1919);
or U7001 (N_7001,N_3475,N_914);
nor U7002 (N_7002,N_3590,N_3447);
xnor U7003 (N_7003,N_3480,N_4945);
and U7004 (N_7004,N_4150,N_4982);
xor U7005 (N_7005,N_1357,N_4035);
or U7006 (N_7006,N_980,N_511);
nand U7007 (N_7007,N_1792,N_4789);
or U7008 (N_7008,N_713,N_4216);
or U7009 (N_7009,N_3259,N_3589);
xor U7010 (N_7010,N_4749,N_1231);
xor U7011 (N_7011,N_4772,N_4017);
and U7012 (N_7012,N_3746,N_4798);
or U7013 (N_7013,N_1060,N_976);
nor U7014 (N_7014,N_779,N_3495);
nor U7015 (N_7015,N_1546,N_1138);
xor U7016 (N_7016,N_3683,N_4123);
and U7017 (N_7017,N_3915,N_1495);
xor U7018 (N_7018,N_2575,N_3719);
nand U7019 (N_7019,N_2641,N_2113);
nand U7020 (N_7020,N_1462,N_1460);
nand U7021 (N_7021,N_1198,N_919);
and U7022 (N_7022,N_1637,N_2228);
xor U7023 (N_7023,N_3128,N_1758);
nand U7024 (N_7024,N_4862,N_4089);
and U7025 (N_7025,N_3473,N_3810);
nand U7026 (N_7026,N_3262,N_1702);
xnor U7027 (N_7027,N_4736,N_2505);
or U7028 (N_7028,N_558,N_1996);
nand U7029 (N_7029,N_1720,N_1030);
and U7030 (N_7030,N_4290,N_3107);
nand U7031 (N_7031,N_4501,N_2999);
xor U7032 (N_7032,N_3862,N_3678);
nand U7033 (N_7033,N_1564,N_3950);
nand U7034 (N_7034,N_2543,N_321);
or U7035 (N_7035,N_3410,N_3172);
nor U7036 (N_7036,N_4149,N_463);
nor U7037 (N_7037,N_349,N_3917);
xor U7038 (N_7038,N_2564,N_2364);
nor U7039 (N_7039,N_1553,N_2894);
nand U7040 (N_7040,N_4556,N_259);
or U7041 (N_7041,N_3061,N_4668);
and U7042 (N_7042,N_4063,N_1511);
xor U7043 (N_7043,N_2026,N_2016);
nand U7044 (N_7044,N_492,N_286);
or U7045 (N_7045,N_2003,N_3378);
nor U7046 (N_7046,N_4319,N_1086);
and U7047 (N_7047,N_460,N_3283);
or U7048 (N_7048,N_3541,N_2778);
nor U7049 (N_7049,N_1180,N_3239);
or U7050 (N_7050,N_3730,N_708);
nor U7051 (N_7051,N_85,N_3577);
nor U7052 (N_7052,N_1539,N_4396);
nor U7053 (N_7053,N_4490,N_168);
and U7054 (N_7054,N_4767,N_4073);
or U7055 (N_7055,N_4933,N_2606);
xnor U7056 (N_7056,N_2218,N_2265);
and U7057 (N_7057,N_2365,N_855);
or U7058 (N_7058,N_1828,N_1016);
xnor U7059 (N_7059,N_482,N_3939);
nand U7060 (N_7060,N_2184,N_2447);
and U7061 (N_7061,N_4541,N_2134);
or U7062 (N_7062,N_681,N_1130);
or U7063 (N_7063,N_2100,N_4304);
nand U7064 (N_7064,N_1823,N_4869);
nand U7065 (N_7065,N_1634,N_2008);
and U7066 (N_7066,N_270,N_3365);
nor U7067 (N_7067,N_1592,N_4766);
nand U7068 (N_7068,N_3888,N_1586);
and U7069 (N_7069,N_3816,N_4258);
or U7070 (N_7070,N_178,N_2207);
and U7071 (N_7071,N_4506,N_1271);
or U7072 (N_7072,N_2391,N_4215);
xnor U7073 (N_7073,N_1486,N_2825);
xnor U7074 (N_7074,N_2712,N_1742);
xnor U7075 (N_7075,N_236,N_4010);
or U7076 (N_7076,N_3024,N_3873);
or U7077 (N_7077,N_1106,N_2398);
or U7078 (N_7078,N_4999,N_2297);
or U7079 (N_7079,N_1417,N_1570);
and U7080 (N_7080,N_2237,N_4473);
xor U7081 (N_7081,N_1386,N_3854);
nor U7082 (N_7082,N_1773,N_687);
and U7083 (N_7083,N_1331,N_4681);
xnor U7084 (N_7084,N_646,N_3009);
nor U7085 (N_7085,N_354,N_3556);
nor U7086 (N_7086,N_4753,N_2971);
or U7087 (N_7087,N_1290,N_4952);
and U7088 (N_7088,N_2070,N_4782);
xnor U7089 (N_7089,N_4729,N_2007);
and U7090 (N_7090,N_4471,N_1576);
and U7091 (N_7091,N_1398,N_949);
and U7092 (N_7092,N_564,N_3560);
or U7093 (N_7093,N_809,N_2765);
and U7094 (N_7094,N_2284,N_3945);
nor U7095 (N_7095,N_4427,N_4888);
xnor U7096 (N_7096,N_2970,N_3004);
nor U7097 (N_7097,N_1626,N_30);
xnor U7098 (N_7098,N_2829,N_2201);
nand U7099 (N_7099,N_963,N_3861);
xor U7100 (N_7100,N_1506,N_1010);
nand U7101 (N_7101,N_2191,N_3347);
nor U7102 (N_7102,N_712,N_3164);
nand U7103 (N_7103,N_1868,N_3644);
nand U7104 (N_7104,N_3277,N_783);
and U7105 (N_7105,N_1901,N_823);
nor U7106 (N_7106,N_1409,N_2287);
nand U7107 (N_7107,N_1197,N_1613);
xnor U7108 (N_7108,N_2700,N_2552);
xnor U7109 (N_7109,N_3989,N_2246);
or U7110 (N_7110,N_750,N_793);
nor U7111 (N_7111,N_4883,N_2301);
nand U7112 (N_7112,N_959,N_3136);
nand U7113 (N_7113,N_2830,N_4811);
nand U7114 (N_7114,N_2325,N_2515);
and U7115 (N_7115,N_3492,N_1418);
xor U7116 (N_7116,N_1928,N_1781);
or U7117 (N_7117,N_3092,N_2106);
or U7118 (N_7118,N_2159,N_4633);
and U7119 (N_7119,N_940,N_801);
and U7120 (N_7120,N_64,N_3598);
xnor U7121 (N_7121,N_3469,N_903);
nor U7122 (N_7122,N_2644,N_1638);
nand U7123 (N_7123,N_3441,N_3581);
and U7124 (N_7124,N_2145,N_36);
and U7125 (N_7125,N_653,N_4867);
and U7126 (N_7126,N_166,N_391);
xor U7127 (N_7127,N_4987,N_2086);
nand U7128 (N_7128,N_263,N_4433);
xor U7129 (N_7129,N_4391,N_3302);
nor U7130 (N_7130,N_2259,N_845);
or U7131 (N_7131,N_3622,N_3100);
nor U7132 (N_7132,N_819,N_2482);
or U7133 (N_7133,N_4415,N_2150);
nor U7134 (N_7134,N_3397,N_858);
or U7135 (N_7135,N_2502,N_970);
xnor U7136 (N_7136,N_3288,N_4435);
nor U7137 (N_7137,N_4816,N_1850);
and U7138 (N_7138,N_2168,N_667);
nand U7139 (N_7139,N_2872,N_2908);
and U7140 (N_7140,N_1855,N_1735);
or U7141 (N_7141,N_490,N_4160);
nand U7142 (N_7142,N_4548,N_2566);
nor U7143 (N_7143,N_2154,N_2677);
nor U7144 (N_7144,N_1087,N_2693);
or U7145 (N_7145,N_3505,N_4361);
and U7146 (N_7146,N_1536,N_4656);
nor U7147 (N_7147,N_3686,N_2947);
xor U7148 (N_7148,N_1058,N_3647);
nor U7149 (N_7149,N_3108,N_2737);
xor U7150 (N_7150,N_2469,N_2568);
or U7151 (N_7151,N_1704,N_3310);
and U7152 (N_7152,N_1923,N_3537);
nand U7153 (N_7153,N_2270,N_1067);
and U7154 (N_7154,N_4742,N_933);
xor U7155 (N_7155,N_1672,N_265);
and U7156 (N_7156,N_3621,N_1041);
nor U7157 (N_7157,N_4534,N_43);
or U7158 (N_7158,N_2936,N_3075);
nor U7159 (N_7159,N_160,N_4640);
or U7160 (N_7160,N_1661,N_4495);
nor U7161 (N_7161,N_1743,N_3898);
and U7162 (N_7162,N_3457,N_4143);
xnor U7163 (N_7163,N_899,N_3425);
xor U7164 (N_7164,N_4020,N_4316);
nor U7165 (N_7165,N_4389,N_4300);
xor U7166 (N_7166,N_1906,N_3186);
nor U7167 (N_7167,N_3312,N_1257);
nand U7168 (N_7168,N_3928,N_4343);
nor U7169 (N_7169,N_1074,N_1031);
nor U7170 (N_7170,N_4654,N_2135);
xnor U7171 (N_7171,N_4463,N_2937);
xor U7172 (N_7172,N_767,N_2043);
xor U7173 (N_7173,N_542,N_3748);
nor U7174 (N_7174,N_434,N_2603);
nor U7175 (N_7175,N_4016,N_1039);
nand U7176 (N_7176,N_2595,N_690);
nor U7177 (N_7177,N_2094,N_3027);
or U7178 (N_7178,N_820,N_1594);
and U7179 (N_7179,N_2302,N_255);
nand U7180 (N_7180,N_2315,N_4861);
and U7181 (N_7181,N_1560,N_355);
nor U7182 (N_7182,N_3777,N_1077);
or U7183 (N_7183,N_531,N_3188);
and U7184 (N_7184,N_4221,N_3084);
nand U7185 (N_7185,N_535,N_835);
nand U7186 (N_7186,N_3223,N_2464);
xnor U7187 (N_7187,N_2486,N_1545);
nor U7188 (N_7188,N_2799,N_4436);
and U7189 (N_7189,N_3741,N_3363);
xnor U7190 (N_7190,N_1547,N_3887);
or U7191 (N_7191,N_93,N_4309);
nor U7192 (N_7192,N_3500,N_649);
and U7193 (N_7193,N_1240,N_3740);
or U7194 (N_7194,N_2087,N_1196);
or U7195 (N_7195,N_3533,N_4156);
and U7196 (N_7196,N_3688,N_225);
and U7197 (N_7197,N_2095,N_998);
or U7198 (N_7198,N_1056,N_930);
and U7199 (N_7199,N_4402,N_2019);
xor U7200 (N_7200,N_1292,N_3025);
and U7201 (N_7201,N_1532,N_339);
xnor U7202 (N_7202,N_3087,N_4967);
nor U7203 (N_7203,N_1766,N_184);
or U7204 (N_7204,N_224,N_4481);
nand U7205 (N_7205,N_2158,N_4165);
nor U7206 (N_7206,N_4859,N_975);
nand U7207 (N_7207,N_1998,N_3700);
nor U7208 (N_7208,N_3133,N_2023);
nor U7209 (N_7209,N_2401,N_2376);
or U7210 (N_7210,N_1598,N_837);
and U7211 (N_7211,N_2646,N_1109);
nand U7212 (N_7212,N_4344,N_4596);
xnor U7213 (N_7213,N_3150,N_875);
nand U7214 (N_7214,N_3506,N_2833);
xor U7215 (N_7215,N_1822,N_4699);
nand U7216 (N_7216,N_4705,N_3224);
xor U7217 (N_7217,N_1695,N_4451);
nor U7218 (N_7218,N_2555,N_2738);
and U7219 (N_7219,N_1426,N_4004);
nand U7220 (N_7220,N_4632,N_3940);
nor U7221 (N_7221,N_1132,N_3743);
xor U7222 (N_7222,N_3966,N_1095);
nand U7223 (N_7223,N_2522,N_4292);
or U7224 (N_7224,N_298,N_3742);
and U7225 (N_7225,N_4437,N_4885);
nand U7226 (N_7226,N_2122,N_3272);
xor U7227 (N_7227,N_4423,N_3871);
xor U7228 (N_7228,N_553,N_2072);
nor U7229 (N_7229,N_4486,N_4761);
or U7230 (N_7230,N_2571,N_432);
xor U7231 (N_7231,N_3501,N_3699);
or U7232 (N_7232,N_578,N_3415);
nand U7233 (N_7233,N_4280,N_517);
nor U7234 (N_7234,N_2818,N_1458);
nor U7235 (N_7235,N_3793,N_4381);
or U7236 (N_7236,N_3648,N_1124);
xor U7237 (N_7237,N_913,N_1821);
nand U7238 (N_7238,N_340,N_3669);
or U7239 (N_7239,N_1696,N_882);
and U7240 (N_7240,N_2796,N_1245);
xor U7241 (N_7241,N_2782,N_363);
xnor U7242 (N_7242,N_3645,N_3750);
or U7243 (N_7243,N_3479,N_2477);
or U7244 (N_7244,N_546,N_2144);
xor U7245 (N_7245,N_4886,N_3258);
or U7246 (N_7246,N_3734,N_4061);
nor U7247 (N_7247,N_1976,N_4270);
xnor U7248 (N_7248,N_761,N_1450);
nand U7249 (N_7249,N_2449,N_4349);
and U7250 (N_7250,N_272,N_3813);
or U7251 (N_7251,N_675,N_4039);
and U7252 (N_7252,N_4617,N_2353);
nor U7253 (N_7253,N_4565,N_857);
xnor U7254 (N_7254,N_4485,N_3045);
and U7255 (N_7255,N_2367,N_493);
xnor U7256 (N_7256,N_3388,N_3718);
or U7257 (N_7257,N_1278,N_2452);
or U7258 (N_7258,N_1579,N_196);
and U7259 (N_7259,N_1388,N_2912);
nand U7260 (N_7260,N_3874,N_118);
xor U7261 (N_7261,N_964,N_2514);
or U7262 (N_7262,N_773,N_1813);
nor U7263 (N_7263,N_4578,N_389);
or U7264 (N_7264,N_2360,N_2489);
nand U7265 (N_7265,N_154,N_1226);
nand U7266 (N_7266,N_218,N_4953);
nand U7267 (N_7267,N_1269,N_2775);
xor U7268 (N_7268,N_1027,N_102);
nand U7269 (N_7269,N_151,N_3822);
or U7270 (N_7270,N_3126,N_3906);
or U7271 (N_7271,N_2382,N_1860);
or U7272 (N_7272,N_3763,N_4815);
and U7273 (N_7273,N_4641,N_1123);
xor U7274 (N_7274,N_3207,N_2685);
nor U7275 (N_7275,N_503,N_4603);
or U7276 (N_7276,N_317,N_3538);
xnor U7277 (N_7277,N_1941,N_3603);
and U7278 (N_7278,N_4060,N_2795);
and U7279 (N_7279,N_3204,N_1159);
or U7280 (N_7280,N_2140,N_4408);
and U7281 (N_7281,N_260,N_3282);
and U7282 (N_7282,N_2993,N_680);
xnor U7283 (N_7283,N_3515,N_2698);
or U7284 (N_7284,N_929,N_221);
or U7285 (N_7285,N_895,N_3960);
xor U7286 (N_7286,N_2491,N_3689);
nand U7287 (N_7287,N_3496,N_4379);
and U7288 (N_7288,N_4755,N_269);
and U7289 (N_7289,N_1224,N_4575);
xor U7290 (N_7290,N_3358,N_4762);
and U7291 (N_7291,N_2235,N_3090);
nor U7292 (N_7292,N_4646,N_19);
or U7293 (N_7293,N_1175,N_385);
nor U7294 (N_7294,N_1503,N_870);
nand U7295 (N_7295,N_2506,N_362);
or U7296 (N_7296,N_1756,N_4322);
nand U7297 (N_7297,N_2656,N_1059);
nor U7298 (N_7298,N_1446,N_2953);
and U7299 (N_7299,N_4417,N_4841);
xor U7300 (N_7300,N_4351,N_3650);
and U7301 (N_7301,N_2577,N_3801);
and U7302 (N_7302,N_1543,N_2767);
nand U7303 (N_7303,N_2596,N_1744);
or U7304 (N_7304,N_1488,N_2710);
nand U7305 (N_7305,N_2791,N_2861);
xnor U7306 (N_7306,N_552,N_4983);
and U7307 (N_7307,N_2006,N_2605);
or U7308 (N_7308,N_2480,N_4703);
or U7309 (N_7309,N_440,N_3850);
nor U7310 (N_7310,N_4224,N_3466);
or U7311 (N_7311,N_4497,N_3789);
and U7312 (N_7312,N_3432,N_1345);
or U7313 (N_7313,N_3304,N_1824);
nand U7314 (N_7314,N_1763,N_606);
or U7315 (N_7315,N_2787,N_1012);
or U7316 (N_7316,N_4331,N_1384);
xor U7317 (N_7317,N_2924,N_1247);
xnor U7318 (N_7318,N_3587,N_2120);
nor U7319 (N_7319,N_4517,N_3504);
and U7320 (N_7320,N_3181,N_1359);
xnor U7321 (N_7321,N_3354,N_4995);
or U7322 (N_7322,N_3073,N_4817);
nand U7323 (N_7323,N_27,N_3161);
nor U7324 (N_7324,N_892,N_2983);
nor U7325 (N_7325,N_2895,N_607);
nand U7326 (N_7326,N_3885,N_2110);
or U7327 (N_7327,N_4509,N_2347);
or U7328 (N_7328,N_1582,N_258);
and U7329 (N_7329,N_2792,N_3831);
nand U7330 (N_7330,N_2982,N_3963);
xor U7331 (N_7331,N_2631,N_1286);
xor U7332 (N_7332,N_158,N_1603);
and U7333 (N_7333,N_660,N_2358);
xnor U7334 (N_7334,N_407,N_2745);
or U7335 (N_7335,N_15,N_2889);
or U7336 (N_7336,N_152,N_1846);
nor U7337 (N_7337,N_3116,N_1549);
or U7338 (N_7338,N_1678,N_2194);
and U7339 (N_7339,N_1814,N_898);
nor U7340 (N_7340,N_1839,N_2271);
or U7341 (N_7341,N_2200,N_2073);
and U7342 (N_7342,N_4583,N_2797);
nor U7343 (N_7343,N_1848,N_3991);
xor U7344 (N_7344,N_2101,N_293);
nor U7345 (N_7345,N_2182,N_3990);
nand U7346 (N_7346,N_361,N_3322);
or U7347 (N_7347,N_4164,N_1651);
xor U7348 (N_7348,N_3021,N_436);
or U7349 (N_7349,N_1496,N_1609);
or U7350 (N_7350,N_4173,N_4266);
and U7351 (N_7351,N_4511,N_229);
nand U7352 (N_7352,N_3261,N_2067);
nor U7353 (N_7353,N_2623,N_992);
and U7354 (N_7354,N_4846,N_2959);
or U7355 (N_7355,N_2213,N_4780);
and U7356 (N_7356,N_860,N_4847);
xnor U7357 (N_7357,N_533,N_1145);
xor U7358 (N_7358,N_760,N_3208);
xor U7359 (N_7359,N_4748,N_2844);
and U7360 (N_7360,N_1046,N_2209);
nor U7361 (N_7361,N_3728,N_1895);
and U7362 (N_7362,N_4332,N_4963);
nand U7363 (N_7363,N_2935,N_4307);
nand U7364 (N_7364,N_745,N_3216);
and U7365 (N_7365,N_1907,N_2243);
or U7366 (N_7366,N_2746,N_4977);
nand U7367 (N_7367,N_4477,N_2052);
or U7368 (N_7368,N_1540,N_3965);
and U7369 (N_7369,N_4365,N_1715);
or U7370 (N_7370,N_3520,N_2327);
xor U7371 (N_7371,N_2688,N_3807);
and U7372 (N_7372,N_1944,N_413);
nand U7373 (N_7373,N_2655,N_2160);
or U7374 (N_7374,N_2716,N_953);
nor U7375 (N_7375,N_3919,N_4993);
or U7376 (N_7376,N_365,N_4411);
xnor U7377 (N_7377,N_513,N_87);
xor U7378 (N_7378,N_2162,N_1236);
and U7379 (N_7379,N_1485,N_4325);
or U7380 (N_7380,N_1512,N_4980);
nor U7381 (N_7381,N_1963,N_768);
nor U7382 (N_7382,N_3280,N_1328);
or U7383 (N_7383,N_1383,N_1002);
xnor U7384 (N_7384,N_1282,N_2523);
nand U7385 (N_7385,N_1099,N_1003);
or U7386 (N_7386,N_4271,N_1723);
and U7387 (N_7387,N_1614,N_3076);
xnor U7388 (N_7388,N_1552,N_610);
or U7389 (N_7389,N_1599,N_1096);
nand U7390 (N_7390,N_1679,N_3430);
xor U7391 (N_7391,N_1262,N_1989);
nor U7392 (N_7392,N_3355,N_3474);
nor U7393 (N_7393,N_1311,N_378);
xnor U7394 (N_7394,N_3348,N_445);
and U7395 (N_7395,N_3445,N_2996);
or U7396 (N_7396,N_4515,N_1836);
nor U7397 (N_7397,N_2804,N_191);
xor U7398 (N_7398,N_1329,N_4917);
and U7399 (N_7399,N_1101,N_2940);
xnor U7400 (N_7400,N_3759,N_3063);
nand U7401 (N_7401,N_4955,N_3486);
xnor U7402 (N_7402,N_4781,N_3218);
xnor U7403 (N_7403,N_4359,N_3029);
or U7404 (N_7404,N_2742,N_83);
or U7405 (N_7405,N_756,N_1520);
nand U7406 (N_7406,N_2108,N_4921);
xor U7407 (N_7407,N_3941,N_3583);
nor U7408 (N_7408,N_4419,N_2992);
xnor U7409 (N_7409,N_4190,N_2840);
and U7410 (N_7410,N_510,N_4825);
xor U7411 (N_7411,N_4278,N_748);
xor U7412 (N_7412,N_3522,N_1258);
and U7413 (N_7413,N_2803,N_4329);
and U7414 (N_7414,N_2034,N_379);
xor U7415 (N_7415,N_4208,N_3481);
and U7416 (N_7416,N_1841,N_3512);
nand U7417 (N_7417,N_3867,N_3391);
or U7418 (N_7418,N_3422,N_688);
and U7419 (N_7419,N_4756,N_1453);
nand U7420 (N_7420,N_3682,N_2713);
xnor U7421 (N_7421,N_2349,N_2130);
nor U7422 (N_7422,N_2061,N_3052);
nor U7423 (N_7423,N_2185,N_3257);
nor U7424 (N_7424,N_4414,N_4890);
xnor U7425 (N_7425,N_1524,N_4446);
xnor U7426 (N_7426,N_2707,N_1215);
or U7427 (N_7427,N_22,N_863);
and U7428 (N_7428,N_1469,N_706);
and U7429 (N_7429,N_1133,N_4491);
nand U7430 (N_7430,N_3157,N_2226);
nand U7431 (N_7431,N_3332,N_2752);
nand U7432 (N_7432,N_1700,N_1005);
xor U7433 (N_7433,N_771,N_4741);
and U7434 (N_7434,N_4205,N_2011);
xnor U7435 (N_7435,N_4347,N_1755);
or U7436 (N_7436,N_633,N_2306);
and U7437 (N_7437,N_888,N_1605);
and U7438 (N_7438,N_3773,N_1655);
xor U7439 (N_7439,N_1250,N_3593);
and U7440 (N_7440,N_4588,N_4001);
and U7441 (N_7441,N_3377,N_3829);
and U7442 (N_7442,N_812,N_3744);
and U7443 (N_7443,N_1273,N_3206);
or U7444 (N_7444,N_3663,N_4591);
and U7445 (N_7445,N_1274,N_4701);
and U7446 (N_7446,N_2995,N_2604);
xnor U7447 (N_7447,N_1811,N_4181);
or U7448 (N_7448,N_1573,N_912);
nand U7449 (N_7449,N_2826,N_3236);
or U7450 (N_7450,N_714,N_3787);
nor U7451 (N_7451,N_3449,N_2172);
nor U7452 (N_7452,N_2602,N_105);
and U7453 (N_7453,N_4430,N_1253);
xor U7454 (N_7454,N_58,N_573);
nand U7455 (N_7455,N_4425,N_4950);
or U7456 (N_7456,N_177,N_3233);
or U7457 (N_7457,N_1517,N_3413);
nand U7458 (N_7458,N_2033,N_53);
or U7459 (N_7459,N_1324,N_4157);
nand U7460 (N_7460,N_840,N_4005);
nand U7461 (N_7461,N_2406,N_2559);
nand U7462 (N_7462,N_1148,N_3606);
and U7463 (N_7463,N_1881,N_487);
xnor U7464 (N_7464,N_4935,N_297);
and U7465 (N_7465,N_3876,N_4673);
xor U7466 (N_7466,N_4750,N_4626);
nor U7467 (N_7467,N_2439,N_1013);
nand U7468 (N_7468,N_2892,N_3448);
nand U7469 (N_7469,N_721,N_1479);
and U7470 (N_7470,N_2465,N_3068);
and U7471 (N_7471,N_3982,N_602);
or U7472 (N_7472,N_392,N_2879);
and U7473 (N_7473,N_4822,N_194);
and U7474 (N_7474,N_886,N_2909);
xnor U7475 (N_7475,N_1321,N_590);
xor U7476 (N_7476,N_1260,N_4719);
xor U7477 (N_7477,N_629,N_1208);
and U7478 (N_7478,N_1156,N_4620);
nor U7479 (N_7479,N_3961,N_1194);
and U7480 (N_7480,N_1296,N_676);
or U7481 (N_7481,N_1052,N_3946);
nand U7482 (N_7482,N_3690,N_2414);
nand U7483 (N_7483,N_3613,N_719);
nor U7484 (N_7484,N_1804,N_1631);
nor U7485 (N_7485,N_957,N_2273);
or U7486 (N_7486,N_2210,N_3922);
nor U7487 (N_7487,N_1136,N_3180);
nand U7488 (N_7488,N_3248,N_4468);
or U7489 (N_7489,N_4218,N_3130);
xnor U7490 (N_7490,N_1277,N_1017);
nand U7491 (N_7491,N_2728,N_3120);
nand U7492 (N_7492,N_3769,N_2556);
or U7493 (N_7493,N_18,N_4897);
xor U7494 (N_7494,N_26,N_1211);
nand U7495 (N_7495,N_2197,N_506);
xnor U7496 (N_7496,N_2734,N_547);
and U7497 (N_7497,N_1908,N_2705);
nor U7498 (N_7498,N_2794,N_4462);
nor U7499 (N_7499,N_3349,N_3050);
nor U7500 (N_7500,N_2291,N_1008);
and U7501 (N_7501,N_1138,N_4699);
nand U7502 (N_7502,N_2600,N_3434);
nand U7503 (N_7503,N_4987,N_2525);
xnor U7504 (N_7504,N_3124,N_495);
nor U7505 (N_7505,N_3124,N_2551);
nor U7506 (N_7506,N_717,N_2825);
xnor U7507 (N_7507,N_1805,N_351);
xor U7508 (N_7508,N_4475,N_3974);
and U7509 (N_7509,N_3226,N_4161);
nor U7510 (N_7510,N_2254,N_4302);
nor U7511 (N_7511,N_1170,N_3005);
nand U7512 (N_7512,N_2122,N_4277);
xor U7513 (N_7513,N_4949,N_2896);
or U7514 (N_7514,N_80,N_2150);
nand U7515 (N_7515,N_202,N_879);
and U7516 (N_7516,N_1263,N_4793);
xnor U7517 (N_7517,N_2610,N_3952);
nand U7518 (N_7518,N_1931,N_2676);
xor U7519 (N_7519,N_3588,N_3720);
or U7520 (N_7520,N_1320,N_503);
nor U7521 (N_7521,N_3580,N_1197);
nand U7522 (N_7522,N_821,N_788);
and U7523 (N_7523,N_573,N_2086);
xnor U7524 (N_7524,N_4778,N_3018);
and U7525 (N_7525,N_4008,N_941);
or U7526 (N_7526,N_1884,N_3872);
xnor U7527 (N_7527,N_4425,N_4265);
nand U7528 (N_7528,N_1492,N_2797);
xnor U7529 (N_7529,N_4040,N_1803);
or U7530 (N_7530,N_4783,N_333);
or U7531 (N_7531,N_1303,N_4595);
nand U7532 (N_7532,N_2426,N_308);
nor U7533 (N_7533,N_4553,N_3607);
xor U7534 (N_7534,N_1047,N_820);
nand U7535 (N_7535,N_510,N_4262);
and U7536 (N_7536,N_3501,N_3992);
and U7537 (N_7537,N_1547,N_4665);
or U7538 (N_7538,N_780,N_1293);
nor U7539 (N_7539,N_3134,N_4996);
xor U7540 (N_7540,N_2905,N_783);
or U7541 (N_7541,N_798,N_3569);
or U7542 (N_7542,N_2278,N_77);
or U7543 (N_7543,N_2880,N_4344);
nor U7544 (N_7544,N_2511,N_951);
and U7545 (N_7545,N_471,N_3496);
or U7546 (N_7546,N_1066,N_367);
nand U7547 (N_7547,N_4593,N_1714);
or U7548 (N_7548,N_2701,N_561);
nor U7549 (N_7549,N_1563,N_1389);
or U7550 (N_7550,N_1113,N_1385);
nor U7551 (N_7551,N_539,N_4566);
nand U7552 (N_7552,N_2251,N_3680);
or U7553 (N_7553,N_3797,N_1244);
nand U7554 (N_7554,N_2114,N_4956);
xor U7555 (N_7555,N_4403,N_61);
or U7556 (N_7556,N_4820,N_1426);
or U7557 (N_7557,N_1478,N_4445);
nor U7558 (N_7558,N_2058,N_2310);
and U7559 (N_7559,N_171,N_2830);
or U7560 (N_7560,N_4966,N_522);
nor U7561 (N_7561,N_2545,N_1611);
or U7562 (N_7562,N_539,N_2957);
and U7563 (N_7563,N_2798,N_222);
nor U7564 (N_7564,N_316,N_2222);
nand U7565 (N_7565,N_265,N_4862);
xnor U7566 (N_7566,N_225,N_4087);
and U7567 (N_7567,N_3947,N_4649);
xnor U7568 (N_7568,N_49,N_377);
nand U7569 (N_7569,N_238,N_1462);
nand U7570 (N_7570,N_4592,N_4116);
or U7571 (N_7571,N_409,N_1674);
nor U7572 (N_7572,N_1838,N_3225);
nor U7573 (N_7573,N_2483,N_1445);
or U7574 (N_7574,N_4610,N_449);
and U7575 (N_7575,N_4739,N_2728);
and U7576 (N_7576,N_3502,N_1419);
nand U7577 (N_7577,N_3028,N_4873);
or U7578 (N_7578,N_240,N_1567);
nor U7579 (N_7579,N_3440,N_3617);
nor U7580 (N_7580,N_4078,N_3338);
or U7581 (N_7581,N_4529,N_3430);
xor U7582 (N_7582,N_614,N_2011);
xnor U7583 (N_7583,N_1567,N_4543);
nor U7584 (N_7584,N_1633,N_4736);
nor U7585 (N_7585,N_1864,N_1763);
nand U7586 (N_7586,N_4659,N_1531);
xor U7587 (N_7587,N_1114,N_3737);
nand U7588 (N_7588,N_4273,N_4135);
nor U7589 (N_7589,N_4330,N_3932);
and U7590 (N_7590,N_2345,N_2132);
and U7591 (N_7591,N_541,N_3958);
nand U7592 (N_7592,N_3087,N_527);
nor U7593 (N_7593,N_3323,N_2177);
or U7594 (N_7594,N_2582,N_3517);
nand U7595 (N_7595,N_4913,N_678);
and U7596 (N_7596,N_4518,N_1651);
and U7597 (N_7597,N_2393,N_1572);
or U7598 (N_7598,N_4503,N_3895);
nand U7599 (N_7599,N_99,N_3023);
nor U7600 (N_7600,N_2114,N_641);
and U7601 (N_7601,N_4102,N_3072);
xor U7602 (N_7602,N_2453,N_4267);
or U7603 (N_7603,N_4262,N_3846);
xnor U7604 (N_7604,N_2141,N_3030);
xnor U7605 (N_7605,N_4318,N_1514);
and U7606 (N_7606,N_4446,N_1534);
nand U7607 (N_7607,N_230,N_2258);
nand U7608 (N_7608,N_259,N_3890);
and U7609 (N_7609,N_3575,N_2425);
or U7610 (N_7610,N_395,N_4002);
and U7611 (N_7611,N_3780,N_3857);
xnor U7612 (N_7612,N_3747,N_2617);
or U7613 (N_7613,N_2891,N_2319);
nor U7614 (N_7614,N_3702,N_1142);
nand U7615 (N_7615,N_4543,N_4278);
nor U7616 (N_7616,N_589,N_3185);
or U7617 (N_7617,N_4846,N_1900);
nor U7618 (N_7618,N_1578,N_4645);
xnor U7619 (N_7619,N_1507,N_4933);
nand U7620 (N_7620,N_1400,N_1203);
xnor U7621 (N_7621,N_978,N_2463);
xnor U7622 (N_7622,N_1139,N_3563);
nor U7623 (N_7623,N_1170,N_4882);
nand U7624 (N_7624,N_375,N_4677);
nand U7625 (N_7625,N_4778,N_1975);
xnor U7626 (N_7626,N_3065,N_1986);
nand U7627 (N_7627,N_1552,N_1179);
nor U7628 (N_7628,N_548,N_3362);
and U7629 (N_7629,N_4540,N_198);
and U7630 (N_7630,N_2172,N_3900);
xor U7631 (N_7631,N_3273,N_4671);
xnor U7632 (N_7632,N_3050,N_4779);
xor U7633 (N_7633,N_1410,N_4350);
xnor U7634 (N_7634,N_3158,N_4273);
or U7635 (N_7635,N_1341,N_143);
nand U7636 (N_7636,N_2002,N_3171);
and U7637 (N_7637,N_4920,N_996);
and U7638 (N_7638,N_2093,N_3689);
and U7639 (N_7639,N_2407,N_3073);
xor U7640 (N_7640,N_1568,N_3796);
xnor U7641 (N_7641,N_4106,N_567);
or U7642 (N_7642,N_391,N_2709);
or U7643 (N_7643,N_4652,N_1529);
or U7644 (N_7644,N_59,N_1982);
or U7645 (N_7645,N_3225,N_3902);
and U7646 (N_7646,N_3366,N_4121);
or U7647 (N_7647,N_4175,N_680);
or U7648 (N_7648,N_1730,N_4372);
and U7649 (N_7649,N_3231,N_1662);
xnor U7650 (N_7650,N_4136,N_145);
nand U7651 (N_7651,N_4534,N_2166);
xnor U7652 (N_7652,N_3353,N_3756);
nand U7653 (N_7653,N_4511,N_1281);
nor U7654 (N_7654,N_3812,N_2426);
nand U7655 (N_7655,N_3829,N_4258);
xnor U7656 (N_7656,N_1786,N_2705);
xor U7657 (N_7657,N_2471,N_210);
nand U7658 (N_7658,N_3413,N_4681);
and U7659 (N_7659,N_2387,N_3650);
nor U7660 (N_7660,N_1357,N_165);
nand U7661 (N_7661,N_3629,N_1082);
nor U7662 (N_7662,N_3857,N_2757);
nand U7663 (N_7663,N_4962,N_3173);
nor U7664 (N_7664,N_224,N_2718);
or U7665 (N_7665,N_4827,N_3780);
nand U7666 (N_7666,N_3383,N_452);
nand U7667 (N_7667,N_4083,N_4476);
nor U7668 (N_7668,N_4561,N_4803);
and U7669 (N_7669,N_4763,N_3271);
and U7670 (N_7670,N_1141,N_3186);
and U7671 (N_7671,N_1916,N_3173);
xnor U7672 (N_7672,N_3790,N_4020);
nor U7673 (N_7673,N_4063,N_3139);
and U7674 (N_7674,N_160,N_110);
nand U7675 (N_7675,N_4575,N_3321);
nor U7676 (N_7676,N_1075,N_754);
xor U7677 (N_7677,N_4101,N_3903);
xnor U7678 (N_7678,N_520,N_308);
and U7679 (N_7679,N_1471,N_3864);
and U7680 (N_7680,N_2967,N_177);
nand U7681 (N_7681,N_4294,N_928);
nor U7682 (N_7682,N_1877,N_689);
or U7683 (N_7683,N_2468,N_3882);
xor U7684 (N_7684,N_1813,N_348);
nor U7685 (N_7685,N_3159,N_400);
nand U7686 (N_7686,N_122,N_718);
nor U7687 (N_7687,N_3030,N_3385);
or U7688 (N_7688,N_1905,N_642);
nand U7689 (N_7689,N_576,N_107);
or U7690 (N_7690,N_4268,N_1971);
nor U7691 (N_7691,N_3011,N_3697);
nand U7692 (N_7692,N_360,N_1972);
nand U7693 (N_7693,N_2827,N_3532);
nand U7694 (N_7694,N_1219,N_1805);
nand U7695 (N_7695,N_25,N_3545);
nor U7696 (N_7696,N_2823,N_2835);
and U7697 (N_7697,N_352,N_3479);
xnor U7698 (N_7698,N_363,N_1474);
or U7699 (N_7699,N_802,N_4736);
nand U7700 (N_7700,N_2233,N_3229);
or U7701 (N_7701,N_317,N_3574);
nand U7702 (N_7702,N_216,N_1931);
nand U7703 (N_7703,N_1432,N_4244);
nand U7704 (N_7704,N_2896,N_3387);
xnor U7705 (N_7705,N_2174,N_4497);
xnor U7706 (N_7706,N_2788,N_3687);
xnor U7707 (N_7707,N_3417,N_4106);
nor U7708 (N_7708,N_2332,N_3538);
and U7709 (N_7709,N_468,N_1175);
nor U7710 (N_7710,N_3388,N_1462);
nor U7711 (N_7711,N_2004,N_1656);
or U7712 (N_7712,N_1127,N_854);
nand U7713 (N_7713,N_2467,N_1699);
or U7714 (N_7714,N_1081,N_2323);
xnor U7715 (N_7715,N_2486,N_627);
nand U7716 (N_7716,N_588,N_4676);
nand U7717 (N_7717,N_3697,N_3739);
nand U7718 (N_7718,N_699,N_4173);
nand U7719 (N_7719,N_288,N_426);
nand U7720 (N_7720,N_964,N_2378);
nand U7721 (N_7721,N_3735,N_2484);
xnor U7722 (N_7722,N_3027,N_4682);
xnor U7723 (N_7723,N_2493,N_3581);
xor U7724 (N_7724,N_1490,N_1253);
or U7725 (N_7725,N_3410,N_484);
or U7726 (N_7726,N_2031,N_3640);
nor U7727 (N_7727,N_2365,N_4118);
and U7728 (N_7728,N_2561,N_3168);
nor U7729 (N_7729,N_4697,N_3668);
xor U7730 (N_7730,N_1060,N_4247);
or U7731 (N_7731,N_1288,N_347);
xor U7732 (N_7732,N_2393,N_2903);
xnor U7733 (N_7733,N_4107,N_1354);
nor U7734 (N_7734,N_511,N_2097);
nand U7735 (N_7735,N_725,N_3423);
or U7736 (N_7736,N_1973,N_898);
and U7737 (N_7737,N_4421,N_474);
and U7738 (N_7738,N_3950,N_1591);
nand U7739 (N_7739,N_32,N_3413);
xnor U7740 (N_7740,N_4348,N_33);
nor U7741 (N_7741,N_4714,N_3785);
xnor U7742 (N_7742,N_2950,N_1034);
xor U7743 (N_7743,N_4809,N_3742);
xor U7744 (N_7744,N_477,N_4900);
nor U7745 (N_7745,N_3815,N_3246);
nand U7746 (N_7746,N_1180,N_3267);
and U7747 (N_7747,N_1340,N_4408);
xnor U7748 (N_7748,N_875,N_412);
nor U7749 (N_7749,N_4064,N_2358);
nand U7750 (N_7750,N_2094,N_1267);
xnor U7751 (N_7751,N_4329,N_3330);
or U7752 (N_7752,N_701,N_1178);
xor U7753 (N_7753,N_2146,N_3500);
or U7754 (N_7754,N_4877,N_4445);
xnor U7755 (N_7755,N_3118,N_1611);
or U7756 (N_7756,N_1429,N_3263);
nand U7757 (N_7757,N_145,N_2413);
and U7758 (N_7758,N_343,N_3834);
or U7759 (N_7759,N_3965,N_1139);
or U7760 (N_7760,N_3342,N_724);
nor U7761 (N_7761,N_4095,N_1104);
nor U7762 (N_7762,N_4731,N_4493);
or U7763 (N_7763,N_286,N_500);
xor U7764 (N_7764,N_832,N_1482);
or U7765 (N_7765,N_4508,N_3949);
nand U7766 (N_7766,N_1524,N_1357);
nand U7767 (N_7767,N_1776,N_1150);
xnor U7768 (N_7768,N_1548,N_1884);
and U7769 (N_7769,N_369,N_4580);
nor U7770 (N_7770,N_3949,N_253);
nor U7771 (N_7771,N_1410,N_1512);
or U7772 (N_7772,N_3852,N_1729);
xnor U7773 (N_7773,N_2544,N_4599);
nand U7774 (N_7774,N_4792,N_1400);
or U7775 (N_7775,N_2210,N_1439);
nor U7776 (N_7776,N_2066,N_665);
or U7777 (N_7777,N_4700,N_507);
and U7778 (N_7778,N_3233,N_1968);
xor U7779 (N_7779,N_4923,N_173);
nor U7780 (N_7780,N_4439,N_3125);
xor U7781 (N_7781,N_1277,N_1552);
or U7782 (N_7782,N_3514,N_3178);
nor U7783 (N_7783,N_671,N_2279);
xor U7784 (N_7784,N_4786,N_1165);
and U7785 (N_7785,N_4868,N_2069);
nand U7786 (N_7786,N_721,N_3964);
and U7787 (N_7787,N_3724,N_155);
or U7788 (N_7788,N_4936,N_1481);
xnor U7789 (N_7789,N_2056,N_780);
and U7790 (N_7790,N_3720,N_2093);
and U7791 (N_7791,N_947,N_4408);
or U7792 (N_7792,N_1178,N_4272);
xnor U7793 (N_7793,N_3277,N_780);
nor U7794 (N_7794,N_2216,N_4908);
xnor U7795 (N_7795,N_3688,N_4517);
nand U7796 (N_7796,N_3060,N_3992);
nor U7797 (N_7797,N_4440,N_3823);
or U7798 (N_7798,N_172,N_3335);
or U7799 (N_7799,N_2900,N_4888);
nand U7800 (N_7800,N_1516,N_3535);
xnor U7801 (N_7801,N_610,N_1778);
nand U7802 (N_7802,N_1533,N_577);
and U7803 (N_7803,N_2253,N_2481);
nand U7804 (N_7804,N_2126,N_3788);
xnor U7805 (N_7805,N_527,N_4848);
or U7806 (N_7806,N_4028,N_3853);
and U7807 (N_7807,N_373,N_3282);
and U7808 (N_7808,N_4926,N_1844);
nor U7809 (N_7809,N_95,N_868);
and U7810 (N_7810,N_1559,N_4229);
nor U7811 (N_7811,N_1817,N_3872);
xor U7812 (N_7812,N_3964,N_4959);
or U7813 (N_7813,N_910,N_4978);
and U7814 (N_7814,N_4554,N_4755);
or U7815 (N_7815,N_4641,N_2462);
or U7816 (N_7816,N_2313,N_1611);
xor U7817 (N_7817,N_2986,N_3323);
or U7818 (N_7818,N_2891,N_1333);
nor U7819 (N_7819,N_2532,N_2198);
nor U7820 (N_7820,N_3192,N_3473);
or U7821 (N_7821,N_4072,N_2276);
or U7822 (N_7822,N_2815,N_1369);
nand U7823 (N_7823,N_4497,N_725);
and U7824 (N_7824,N_4538,N_2537);
and U7825 (N_7825,N_3112,N_1279);
or U7826 (N_7826,N_2990,N_1304);
and U7827 (N_7827,N_3614,N_2481);
or U7828 (N_7828,N_2618,N_4308);
nand U7829 (N_7829,N_1992,N_1799);
and U7830 (N_7830,N_168,N_3413);
xnor U7831 (N_7831,N_3733,N_4833);
nor U7832 (N_7832,N_3246,N_3713);
and U7833 (N_7833,N_3067,N_3929);
and U7834 (N_7834,N_898,N_2384);
nor U7835 (N_7835,N_1753,N_3034);
xor U7836 (N_7836,N_228,N_3723);
nor U7837 (N_7837,N_2054,N_2452);
xor U7838 (N_7838,N_86,N_1909);
and U7839 (N_7839,N_1005,N_421);
nor U7840 (N_7840,N_2803,N_2075);
nand U7841 (N_7841,N_555,N_4073);
xor U7842 (N_7842,N_574,N_4340);
or U7843 (N_7843,N_2693,N_1991);
and U7844 (N_7844,N_1407,N_3666);
xnor U7845 (N_7845,N_1113,N_3576);
or U7846 (N_7846,N_1656,N_4609);
xnor U7847 (N_7847,N_1361,N_2116);
or U7848 (N_7848,N_149,N_967);
or U7849 (N_7849,N_3085,N_3568);
nor U7850 (N_7850,N_4930,N_1513);
or U7851 (N_7851,N_4371,N_232);
nand U7852 (N_7852,N_1112,N_4626);
nand U7853 (N_7853,N_141,N_1011);
nor U7854 (N_7854,N_1721,N_3047);
and U7855 (N_7855,N_2505,N_2086);
or U7856 (N_7856,N_2878,N_3895);
nand U7857 (N_7857,N_1606,N_506);
and U7858 (N_7858,N_2309,N_1001);
xor U7859 (N_7859,N_19,N_351);
or U7860 (N_7860,N_1341,N_471);
or U7861 (N_7861,N_4156,N_1671);
nor U7862 (N_7862,N_2840,N_2286);
nand U7863 (N_7863,N_2335,N_815);
and U7864 (N_7864,N_1555,N_2771);
xor U7865 (N_7865,N_4682,N_2367);
or U7866 (N_7866,N_4478,N_660);
and U7867 (N_7867,N_3960,N_2916);
or U7868 (N_7868,N_2730,N_3393);
nand U7869 (N_7869,N_678,N_2032);
nand U7870 (N_7870,N_1110,N_4198);
and U7871 (N_7871,N_2209,N_3189);
and U7872 (N_7872,N_281,N_3658);
nand U7873 (N_7873,N_538,N_3232);
xor U7874 (N_7874,N_4306,N_3901);
or U7875 (N_7875,N_3988,N_3095);
and U7876 (N_7876,N_1177,N_3291);
nand U7877 (N_7877,N_1386,N_4303);
nand U7878 (N_7878,N_3670,N_1484);
and U7879 (N_7879,N_896,N_4064);
and U7880 (N_7880,N_1643,N_754);
nand U7881 (N_7881,N_613,N_457);
nor U7882 (N_7882,N_2299,N_2649);
and U7883 (N_7883,N_4607,N_184);
or U7884 (N_7884,N_3403,N_3885);
xor U7885 (N_7885,N_1090,N_2576);
or U7886 (N_7886,N_1744,N_188);
or U7887 (N_7887,N_2538,N_4093);
nand U7888 (N_7888,N_1322,N_4460);
and U7889 (N_7889,N_2289,N_3787);
xor U7890 (N_7890,N_1635,N_2995);
nand U7891 (N_7891,N_3406,N_1537);
and U7892 (N_7892,N_1128,N_2606);
nor U7893 (N_7893,N_2592,N_3255);
nor U7894 (N_7894,N_43,N_1774);
nand U7895 (N_7895,N_2191,N_3396);
nor U7896 (N_7896,N_2039,N_4724);
nor U7897 (N_7897,N_3062,N_1037);
nand U7898 (N_7898,N_3389,N_2386);
and U7899 (N_7899,N_183,N_3366);
and U7900 (N_7900,N_4606,N_2243);
nand U7901 (N_7901,N_416,N_847);
xnor U7902 (N_7902,N_1724,N_3593);
and U7903 (N_7903,N_227,N_2705);
nand U7904 (N_7904,N_3606,N_2458);
nand U7905 (N_7905,N_2304,N_4925);
and U7906 (N_7906,N_2561,N_1252);
nand U7907 (N_7907,N_1215,N_4320);
nand U7908 (N_7908,N_2853,N_3566);
xnor U7909 (N_7909,N_2086,N_4275);
or U7910 (N_7910,N_2201,N_2482);
nor U7911 (N_7911,N_4357,N_1133);
and U7912 (N_7912,N_4412,N_2479);
xnor U7913 (N_7913,N_4849,N_2445);
and U7914 (N_7914,N_4865,N_784);
xnor U7915 (N_7915,N_3830,N_2142);
nor U7916 (N_7916,N_3324,N_535);
xor U7917 (N_7917,N_3839,N_4209);
nor U7918 (N_7918,N_2843,N_2862);
or U7919 (N_7919,N_3829,N_58);
or U7920 (N_7920,N_3886,N_1602);
xnor U7921 (N_7921,N_4776,N_4538);
nand U7922 (N_7922,N_3138,N_725);
nor U7923 (N_7923,N_660,N_3926);
xnor U7924 (N_7924,N_3428,N_3905);
nor U7925 (N_7925,N_4012,N_2674);
and U7926 (N_7926,N_248,N_3993);
nor U7927 (N_7927,N_1317,N_3629);
or U7928 (N_7928,N_1914,N_4799);
nor U7929 (N_7929,N_1544,N_634);
xnor U7930 (N_7930,N_3679,N_835);
nor U7931 (N_7931,N_3629,N_851);
nand U7932 (N_7932,N_3854,N_4353);
and U7933 (N_7933,N_3643,N_2323);
or U7934 (N_7934,N_312,N_1461);
nand U7935 (N_7935,N_2640,N_2532);
xnor U7936 (N_7936,N_692,N_3911);
and U7937 (N_7937,N_4376,N_1401);
xnor U7938 (N_7938,N_943,N_3051);
nand U7939 (N_7939,N_3992,N_973);
xor U7940 (N_7940,N_2119,N_2189);
xnor U7941 (N_7941,N_634,N_2900);
or U7942 (N_7942,N_4901,N_4011);
nor U7943 (N_7943,N_2674,N_3005);
or U7944 (N_7944,N_270,N_2668);
and U7945 (N_7945,N_1836,N_4067);
and U7946 (N_7946,N_2320,N_2050);
xnor U7947 (N_7947,N_3490,N_3631);
nor U7948 (N_7948,N_1300,N_4669);
xor U7949 (N_7949,N_2855,N_2946);
nor U7950 (N_7950,N_3356,N_3239);
xor U7951 (N_7951,N_667,N_1487);
nand U7952 (N_7952,N_1255,N_1942);
and U7953 (N_7953,N_3064,N_2304);
nand U7954 (N_7954,N_4159,N_470);
or U7955 (N_7955,N_3010,N_3909);
xnor U7956 (N_7956,N_1721,N_2446);
and U7957 (N_7957,N_4986,N_845);
xnor U7958 (N_7958,N_1493,N_4002);
or U7959 (N_7959,N_1714,N_1125);
nor U7960 (N_7960,N_58,N_4482);
and U7961 (N_7961,N_3624,N_4364);
xor U7962 (N_7962,N_2268,N_1123);
nand U7963 (N_7963,N_4870,N_3649);
nor U7964 (N_7964,N_1393,N_4118);
and U7965 (N_7965,N_3236,N_619);
nor U7966 (N_7966,N_2748,N_2802);
nor U7967 (N_7967,N_3587,N_382);
and U7968 (N_7968,N_3113,N_4081);
nand U7969 (N_7969,N_49,N_796);
or U7970 (N_7970,N_1850,N_3200);
nand U7971 (N_7971,N_1448,N_928);
nor U7972 (N_7972,N_3410,N_1951);
nor U7973 (N_7973,N_446,N_4051);
xor U7974 (N_7974,N_4238,N_4131);
or U7975 (N_7975,N_3851,N_4568);
nor U7976 (N_7976,N_321,N_4064);
or U7977 (N_7977,N_4808,N_2937);
nor U7978 (N_7978,N_4968,N_4003);
xor U7979 (N_7979,N_3648,N_929);
or U7980 (N_7980,N_4728,N_3744);
nand U7981 (N_7981,N_1490,N_1237);
and U7982 (N_7982,N_2431,N_1203);
xor U7983 (N_7983,N_4804,N_2743);
nand U7984 (N_7984,N_4169,N_2574);
nor U7985 (N_7985,N_4949,N_4287);
xor U7986 (N_7986,N_397,N_571);
or U7987 (N_7987,N_1675,N_4375);
nor U7988 (N_7988,N_1031,N_4981);
xnor U7989 (N_7989,N_3593,N_3798);
xor U7990 (N_7990,N_285,N_3493);
nand U7991 (N_7991,N_1983,N_1710);
or U7992 (N_7992,N_4912,N_379);
nand U7993 (N_7993,N_4569,N_2463);
nand U7994 (N_7994,N_1235,N_1338);
or U7995 (N_7995,N_2017,N_949);
nor U7996 (N_7996,N_4274,N_2716);
or U7997 (N_7997,N_1662,N_4200);
xnor U7998 (N_7998,N_3297,N_1270);
nand U7999 (N_7999,N_1489,N_3380);
nand U8000 (N_8000,N_1978,N_261);
and U8001 (N_8001,N_4014,N_2929);
xnor U8002 (N_8002,N_3819,N_3941);
nand U8003 (N_8003,N_3480,N_4226);
nand U8004 (N_8004,N_565,N_3862);
nor U8005 (N_8005,N_65,N_3445);
xnor U8006 (N_8006,N_3416,N_4508);
nand U8007 (N_8007,N_4236,N_3553);
nor U8008 (N_8008,N_1518,N_3402);
and U8009 (N_8009,N_2888,N_1371);
xor U8010 (N_8010,N_1895,N_4255);
or U8011 (N_8011,N_4960,N_3649);
and U8012 (N_8012,N_1191,N_4353);
and U8013 (N_8013,N_637,N_2113);
or U8014 (N_8014,N_636,N_2519);
and U8015 (N_8015,N_4613,N_1645);
and U8016 (N_8016,N_2589,N_681);
nand U8017 (N_8017,N_2405,N_1558);
xor U8018 (N_8018,N_742,N_245);
and U8019 (N_8019,N_2551,N_2697);
and U8020 (N_8020,N_353,N_2782);
nor U8021 (N_8021,N_3681,N_2470);
or U8022 (N_8022,N_2691,N_3968);
and U8023 (N_8023,N_21,N_4529);
and U8024 (N_8024,N_3220,N_4746);
and U8025 (N_8025,N_678,N_2580);
or U8026 (N_8026,N_2805,N_1488);
xnor U8027 (N_8027,N_1550,N_1109);
xor U8028 (N_8028,N_3709,N_2095);
and U8029 (N_8029,N_2880,N_2596);
xnor U8030 (N_8030,N_210,N_4745);
nor U8031 (N_8031,N_4807,N_3889);
nor U8032 (N_8032,N_3950,N_3790);
or U8033 (N_8033,N_215,N_50);
and U8034 (N_8034,N_1563,N_1811);
xnor U8035 (N_8035,N_2936,N_4256);
and U8036 (N_8036,N_2730,N_4363);
nand U8037 (N_8037,N_1635,N_4423);
and U8038 (N_8038,N_2811,N_721);
or U8039 (N_8039,N_2910,N_2859);
xor U8040 (N_8040,N_588,N_2026);
nor U8041 (N_8041,N_960,N_1886);
or U8042 (N_8042,N_5,N_3325);
or U8043 (N_8043,N_319,N_4005);
and U8044 (N_8044,N_3025,N_3647);
or U8045 (N_8045,N_294,N_1632);
xor U8046 (N_8046,N_4427,N_870);
nand U8047 (N_8047,N_4604,N_834);
or U8048 (N_8048,N_4786,N_1213);
nor U8049 (N_8049,N_4207,N_874);
xnor U8050 (N_8050,N_1736,N_741);
nand U8051 (N_8051,N_1484,N_4429);
and U8052 (N_8052,N_1639,N_555);
xor U8053 (N_8053,N_554,N_1748);
nor U8054 (N_8054,N_2534,N_865);
nor U8055 (N_8055,N_3617,N_3801);
or U8056 (N_8056,N_4173,N_2329);
xor U8057 (N_8057,N_4815,N_4859);
or U8058 (N_8058,N_4434,N_2116);
or U8059 (N_8059,N_2524,N_3770);
nor U8060 (N_8060,N_4914,N_368);
nand U8061 (N_8061,N_2733,N_2477);
nand U8062 (N_8062,N_4894,N_3685);
and U8063 (N_8063,N_4185,N_141);
nand U8064 (N_8064,N_162,N_1307);
nand U8065 (N_8065,N_4162,N_1679);
nand U8066 (N_8066,N_2396,N_2066);
nand U8067 (N_8067,N_1431,N_3837);
nand U8068 (N_8068,N_18,N_4990);
nand U8069 (N_8069,N_4739,N_3500);
xnor U8070 (N_8070,N_929,N_622);
xor U8071 (N_8071,N_3619,N_4317);
xnor U8072 (N_8072,N_4222,N_3920);
nor U8073 (N_8073,N_44,N_3642);
or U8074 (N_8074,N_3127,N_152);
nor U8075 (N_8075,N_826,N_1595);
nand U8076 (N_8076,N_1962,N_3655);
or U8077 (N_8077,N_1953,N_2151);
nor U8078 (N_8078,N_3111,N_4379);
and U8079 (N_8079,N_1054,N_351);
nor U8080 (N_8080,N_3268,N_2815);
and U8081 (N_8081,N_1035,N_2671);
xnor U8082 (N_8082,N_3886,N_3860);
and U8083 (N_8083,N_825,N_2307);
and U8084 (N_8084,N_1032,N_4002);
nand U8085 (N_8085,N_1596,N_3241);
or U8086 (N_8086,N_1711,N_2588);
and U8087 (N_8087,N_942,N_4201);
nor U8088 (N_8088,N_986,N_1004);
and U8089 (N_8089,N_928,N_2794);
and U8090 (N_8090,N_3407,N_4669);
or U8091 (N_8091,N_819,N_957);
and U8092 (N_8092,N_2388,N_1531);
and U8093 (N_8093,N_2453,N_1869);
xor U8094 (N_8094,N_3711,N_4972);
or U8095 (N_8095,N_1455,N_1828);
xnor U8096 (N_8096,N_4528,N_4578);
nor U8097 (N_8097,N_50,N_1599);
xor U8098 (N_8098,N_2661,N_3012);
and U8099 (N_8099,N_690,N_4722);
or U8100 (N_8100,N_4428,N_898);
nor U8101 (N_8101,N_1047,N_190);
nand U8102 (N_8102,N_4177,N_4133);
and U8103 (N_8103,N_3254,N_1);
or U8104 (N_8104,N_1569,N_4633);
and U8105 (N_8105,N_4610,N_2564);
nand U8106 (N_8106,N_2998,N_3819);
xor U8107 (N_8107,N_2581,N_815);
nor U8108 (N_8108,N_655,N_1468);
or U8109 (N_8109,N_1012,N_2348);
xnor U8110 (N_8110,N_920,N_964);
xor U8111 (N_8111,N_1975,N_2103);
nand U8112 (N_8112,N_1512,N_1923);
or U8113 (N_8113,N_4967,N_2660);
and U8114 (N_8114,N_4676,N_2594);
and U8115 (N_8115,N_1837,N_3152);
nand U8116 (N_8116,N_246,N_3033);
nand U8117 (N_8117,N_644,N_4964);
xnor U8118 (N_8118,N_1228,N_2088);
xor U8119 (N_8119,N_3743,N_4899);
or U8120 (N_8120,N_1824,N_385);
and U8121 (N_8121,N_443,N_4072);
or U8122 (N_8122,N_1946,N_3624);
nand U8123 (N_8123,N_463,N_4948);
nor U8124 (N_8124,N_3389,N_2208);
xor U8125 (N_8125,N_860,N_3845);
or U8126 (N_8126,N_585,N_2968);
xor U8127 (N_8127,N_87,N_1902);
or U8128 (N_8128,N_897,N_3985);
nand U8129 (N_8129,N_4669,N_2842);
nand U8130 (N_8130,N_1484,N_3382);
and U8131 (N_8131,N_53,N_4457);
xnor U8132 (N_8132,N_1902,N_626);
and U8133 (N_8133,N_2501,N_3955);
or U8134 (N_8134,N_308,N_1055);
or U8135 (N_8135,N_4653,N_2302);
xnor U8136 (N_8136,N_1438,N_4846);
xor U8137 (N_8137,N_2627,N_4500);
nor U8138 (N_8138,N_3306,N_3482);
nor U8139 (N_8139,N_2280,N_4627);
and U8140 (N_8140,N_745,N_1517);
and U8141 (N_8141,N_809,N_1591);
or U8142 (N_8142,N_1001,N_1210);
xor U8143 (N_8143,N_624,N_2741);
nand U8144 (N_8144,N_2152,N_492);
or U8145 (N_8145,N_625,N_1792);
nor U8146 (N_8146,N_4281,N_3487);
nor U8147 (N_8147,N_1059,N_942);
and U8148 (N_8148,N_2929,N_929);
or U8149 (N_8149,N_4207,N_2477);
and U8150 (N_8150,N_4628,N_3555);
nand U8151 (N_8151,N_144,N_612);
nor U8152 (N_8152,N_4013,N_86);
nor U8153 (N_8153,N_1917,N_2314);
and U8154 (N_8154,N_1522,N_2039);
xnor U8155 (N_8155,N_4276,N_617);
or U8156 (N_8156,N_2505,N_187);
xnor U8157 (N_8157,N_4356,N_148);
and U8158 (N_8158,N_3631,N_1250);
nor U8159 (N_8159,N_1826,N_4670);
xnor U8160 (N_8160,N_3996,N_4289);
and U8161 (N_8161,N_3597,N_39);
nor U8162 (N_8162,N_1530,N_873);
xor U8163 (N_8163,N_706,N_4250);
or U8164 (N_8164,N_4119,N_1394);
nand U8165 (N_8165,N_3139,N_1859);
or U8166 (N_8166,N_621,N_3561);
nand U8167 (N_8167,N_2747,N_935);
and U8168 (N_8168,N_1721,N_831);
nand U8169 (N_8169,N_4864,N_2636);
xnor U8170 (N_8170,N_4377,N_3052);
nor U8171 (N_8171,N_58,N_4710);
and U8172 (N_8172,N_2762,N_3076);
xor U8173 (N_8173,N_119,N_3597);
and U8174 (N_8174,N_2549,N_3492);
and U8175 (N_8175,N_699,N_3260);
nand U8176 (N_8176,N_2193,N_259);
nand U8177 (N_8177,N_1183,N_2730);
and U8178 (N_8178,N_3133,N_1267);
xor U8179 (N_8179,N_544,N_3732);
nor U8180 (N_8180,N_3356,N_960);
xnor U8181 (N_8181,N_2829,N_934);
or U8182 (N_8182,N_3052,N_4661);
xor U8183 (N_8183,N_2420,N_1656);
or U8184 (N_8184,N_2459,N_4153);
and U8185 (N_8185,N_1833,N_1665);
xor U8186 (N_8186,N_1712,N_467);
xor U8187 (N_8187,N_932,N_3266);
nor U8188 (N_8188,N_2164,N_2212);
and U8189 (N_8189,N_4641,N_4453);
and U8190 (N_8190,N_2083,N_830);
nor U8191 (N_8191,N_1538,N_2739);
xor U8192 (N_8192,N_4412,N_123);
xor U8193 (N_8193,N_383,N_265);
nor U8194 (N_8194,N_4667,N_2059);
nand U8195 (N_8195,N_1376,N_2067);
or U8196 (N_8196,N_4325,N_3879);
nor U8197 (N_8197,N_3751,N_1937);
xnor U8198 (N_8198,N_1017,N_974);
nand U8199 (N_8199,N_1412,N_1690);
xnor U8200 (N_8200,N_3204,N_4683);
nor U8201 (N_8201,N_3007,N_2594);
nor U8202 (N_8202,N_1890,N_2564);
xnor U8203 (N_8203,N_2193,N_1812);
xnor U8204 (N_8204,N_1467,N_4982);
nand U8205 (N_8205,N_4218,N_2463);
xor U8206 (N_8206,N_380,N_737);
and U8207 (N_8207,N_4560,N_184);
and U8208 (N_8208,N_3580,N_949);
nand U8209 (N_8209,N_4013,N_3818);
or U8210 (N_8210,N_2107,N_4481);
nand U8211 (N_8211,N_2437,N_275);
and U8212 (N_8212,N_1056,N_2415);
nand U8213 (N_8213,N_4263,N_2696);
or U8214 (N_8214,N_1794,N_973);
or U8215 (N_8215,N_4467,N_2036);
or U8216 (N_8216,N_4346,N_1829);
or U8217 (N_8217,N_2805,N_2981);
nor U8218 (N_8218,N_1620,N_4115);
and U8219 (N_8219,N_4652,N_1517);
or U8220 (N_8220,N_809,N_3463);
nand U8221 (N_8221,N_2671,N_2457);
and U8222 (N_8222,N_1849,N_892);
nand U8223 (N_8223,N_4169,N_2908);
xnor U8224 (N_8224,N_2228,N_1622);
and U8225 (N_8225,N_530,N_4103);
and U8226 (N_8226,N_3213,N_182);
or U8227 (N_8227,N_788,N_3720);
nor U8228 (N_8228,N_1363,N_0);
xnor U8229 (N_8229,N_1454,N_1233);
or U8230 (N_8230,N_234,N_223);
and U8231 (N_8231,N_449,N_4152);
and U8232 (N_8232,N_2083,N_4618);
and U8233 (N_8233,N_3415,N_4984);
and U8234 (N_8234,N_1010,N_4804);
or U8235 (N_8235,N_2420,N_3729);
xnor U8236 (N_8236,N_1496,N_2385);
or U8237 (N_8237,N_2879,N_4544);
or U8238 (N_8238,N_1316,N_1383);
nor U8239 (N_8239,N_4135,N_4912);
and U8240 (N_8240,N_74,N_4624);
nand U8241 (N_8241,N_4902,N_3902);
xor U8242 (N_8242,N_2869,N_4883);
and U8243 (N_8243,N_1322,N_4257);
and U8244 (N_8244,N_4917,N_2647);
nand U8245 (N_8245,N_2470,N_4453);
xnor U8246 (N_8246,N_3915,N_590);
nand U8247 (N_8247,N_4625,N_837);
xor U8248 (N_8248,N_1156,N_635);
and U8249 (N_8249,N_3909,N_427);
or U8250 (N_8250,N_719,N_1614);
nor U8251 (N_8251,N_4164,N_2780);
and U8252 (N_8252,N_3849,N_2737);
nor U8253 (N_8253,N_2241,N_3436);
and U8254 (N_8254,N_427,N_2542);
nand U8255 (N_8255,N_1430,N_4548);
and U8256 (N_8256,N_149,N_3113);
nor U8257 (N_8257,N_1443,N_547);
or U8258 (N_8258,N_1752,N_2815);
nand U8259 (N_8259,N_644,N_3529);
nand U8260 (N_8260,N_382,N_4262);
xor U8261 (N_8261,N_1130,N_384);
nand U8262 (N_8262,N_2782,N_4749);
nand U8263 (N_8263,N_4381,N_3255);
nor U8264 (N_8264,N_4071,N_4479);
nor U8265 (N_8265,N_2642,N_4080);
nand U8266 (N_8266,N_3151,N_643);
nand U8267 (N_8267,N_3548,N_1595);
and U8268 (N_8268,N_3539,N_3267);
nor U8269 (N_8269,N_3442,N_1378);
nor U8270 (N_8270,N_4165,N_2821);
xnor U8271 (N_8271,N_1192,N_3219);
or U8272 (N_8272,N_4450,N_4494);
or U8273 (N_8273,N_3234,N_848);
and U8274 (N_8274,N_3043,N_898);
or U8275 (N_8275,N_2317,N_1185);
nand U8276 (N_8276,N_1427,N_3671);
nor U8277 (N_8277,N_1612,N_3779);
or U8278 (N_8278,N_3336,N_1557);
and U8279 (N_8279,N_2476,N_4407);
nor U8280 (N_8280,N_1214,N_29);
nor U8281 (N_8281,N_4237,N_4923);
nor U8282 (N_8282,N_1840,N_811);
xor U8283 (N_8283,N_4994,N_3478);
xnor U8284 (N_8284,N_2531,N_4815);
or U8285 (N_8285,N_2661,N_1399);
xnor U8286 (N_8286,N_4389,N_568);
and U8287 (N_8287,N_2039,N_1345);
and U8288 (N_8288,N_3388,N_2191);
and U8289 (N_8289,N_1347,N_1744);
nor U8290 (N_8290,N_4649,N_1176);
nor U8291 (N_8291,N_1925,N_2616);
nand U8292 (N_8292,N_3829,N_4567);
and U8293 (N_8293,N_818,N_3369);
nor U8294 (N_8294,N_600,N_3211);
xor U8295 (N_8295,N_1364,N_1696);
xnor U8296 (N_8296,N_3976,N_4212);
or U8297 (N_8297,N_59,N_4315);
nor U8298 (N_8298,N_3735,N_623);
and U8299 (N_8299,N_1172,N_2652);
nand U8300 (N_8300,N_1462,N_1334);
and U8301 (N_8301,N_1472,N_794);
and U8302 (N_8302,N_2167,N_1403);
or U8303 (N_8303,N_608,N_4967);
xor U8304 (N_8304,N_2663,N_3472);
nor U8305 (N_8305,N_2645,N_3579);
nor U8306 (N_8306,N_4194,N_1301);
or U8307 (N_8307,N_1855,N_2143);
xnor U8308 (N_8308,N_221,N_291);
xor U8309 (N_8309,N_3005,N_4327);
nor U8310 (N_8310,N_4939,N_2101);
nor U8311 (N_8311,N_3801,N_4588);
or U8312 (N_8312,N_617,N_655);
or U8313 (N_8313,N_2383,N_578);
nand U8314 (N_8314,N_2607,N_1503);
or U8315 (N_8315,N_2866,N_3887);
xnor U8316 (N_8316,N_1023,N_537);
and U8317 (N_8317,N_997,N_3906);
nand U8318 (N_8318,N_234,N_1160);
and U8319 (N_8319,N_2081,N_2986);
or U8320 (N_8320,N_679,N_1195);
or U8321 (N_8321,N_1668,N_1857);
and U8322 (N_8322,N_4156,N_2470);
nand U8323 (N_8323,N_293,N_706);
nand U8324 (N_8324,N_1780,N_3302);
or U8325 (N_8325,N_2819,N_2057);
nand U8326 (N_8326,N_1218,N_4812);
and U8327 (N_8327,N_2391,N_3830);
xnor U8328 (N_8328,N_2436,N_182);
or U8329 (N_8329,N_2402,N_279);
xnor U8330 (N_8330,N_3529,N_2065);
nor U8331 (N_8331,N_2066,N_2579);
or U8332 (N_8332,N_3192,N_880);
xor U8333 (N_8333,N_3960,N_1771);
and U8334 (N_8334,N_1631,N_3837);
nor U8335 (N_8335,N_3405,N_2769);
nand U8336 (N_8336,N_3732,N_3885);
nand U8337 (N_8337,N_3593,N_2260);
nor U8338 (N_8338,N_4230,N_307);
xor U8339 (N_8339,N_13,N_2774);
nand U8340 (N_8340,N_4862,N_4451);
and U8341 (N_8341,N_2545,N_3718);
nand U8342 (N_8342,N_2816,N_4019);
nand U8343 (N_8343,N_3007,N_1028);
or U8344 (N_8344,N_4762,N_4688);
and U8345 (N_8345,N_1452,N_350);
xnor U8346 (N_8346,N_2970,N_1471);
xor U8347 (N_8347,N_2619,N_260);
nor U8348 (N_8348,N_733,N_4974);
xor U8349 (N_8349,N_843,N_3125);
nor U8350 (N_8350,N_4295,N_954);
nor U8351 (N_8351,N_2319,N_2307);
xnor U8352 (N_8352,N_2442,N_4620);
xnor U8353 (N_8353,N_1732,N_328);
and U8354 (N_8354,N_2172,N_4257);
nor U8355 (N_8355,N_1396,N_727);
nand U8356 (N_8356,N_1569,N_3294);
nand U8357 (N_8357,N_1050,N_4898);
or U8358 (N_8358,N_3242,N_4917);
xor U8359 (N_8359,N_2538,N_1254);
or U8360 (N_8360,N_977,N_1306);
or U8361 (N_8361,N_1632,N_2062);
or U8362 (N_8362,N_3128,N_1221);
nand U8363 (N_8363,N_2844,N_4909);
nand U8364 (N_8364,N_464,N_1005);
nand U8365 (N_8365,N_274,N_2854);
and U8366 (N_8366,N_3568,N_3215);
nor U8367 (N_8367,N_4500,N_2976);
and U8368 (N_8368,N_4655,N_4294);
xor U8369 (N_8369,N_1524,N_1020);
and U8370 (N_8370,N_2398,N_461);
or U8371 (N_8371,N_339,N_3048);
xnor U8372 (N_8372,N_2805,N_212);
nand U8373 (N_8373,N_2866,N_2506);
xor U8374 (N_8374,N_2478,N_3829);
nand U8375 (N_8375,N_3754,N_17);
xor U8376 (N_8376,N_785,N_3632);
and U8377 (N_8377,N_313,N_4372);
nand U8378 (N_8378,N_3231,N_110);
nand U8379 (N_8379,N_2396,N_2576);
xnor U8380 (N_8380,N_1383,N_2282);
and U8381 (N_8381,N_2277,N_994);
or U8382 (N_8382,N_2581,N_3110);
and U8383 (N_8383,N_3815,N_2482);
xor U8384 (N_8384,N_3639,N_4517);
xor U8385 (N_8385,N_1641,N_926);
nor U8386 (N_8386,N_1520,N_3802);
nor U8387 (N_8387,N_3558,N_2930);
or U8388 (N_8388,N_1054,N_3157);
and U8389 (N_8389,N_3239,N_1034);
nand U8390 (N_8390,N_4272,N_2931);
nor U8391 (N_8391,N_1246,N_321);
nor U8392 (N_8392,N_1348,N_990);
nand U8393 (N_8393,N_1859,N_4904);
nand U8394 (N_8394,N_1591,N_642);
xnor U8395 (N_8395,N_2315,N_3385);
and U8396 (N_8396,N_4571,N_3575);
nand U8397 (N_8397,N_913,N_434);
nand U8398 (N_8398,N_4043,N_71);
xnor U8399 (N_8399,N_4934,N_1840);
xor U8400 (N_8400,N_2677,N_1045);
or U8401 (N_8401,N_2141,N_2986);
nor U8402 (N_8402,N_3992,N_2855);
and U8403 (N_8403,N_1386,N_3549);
or U8404 (N_8404,N_3200,N_1921);
nor U8405 (N_8405,N_1993,N_138);
and U8406 (N_8406,N_2306,N_2161);
nand U8407 (N_8407,N_4121,N_3627);
or U8408 (N_8408,N_4316,N_290);
or U8409 (N_8409,N_3280,N_1138);
nand U8410 (N_8410,N_82,N_4961);
xnor U8411 (N_8411,N_3718,N_1540);
nor U8412 (N_8412,N_2661,N_161);
nor U8413 (N_8413,N_117,N_4807);
xor U8414 (N_8414,N_2907,N_3985);
nor U8415 (N_8415,N_2863,N_2621);
nand U8416 (N_8416,N_3174,N_2242);
and U8417 (N_8417,N_93,N_3048);
xnor U8418 (N_8418,N_2142,N_3852);
and U8419 (N_8419,N_431,N_269);
or U8420 (N_8420,N_1783,N_1678);
nand U8421 (N_8421,N_962,N_1314);
nor U8422 (N_8422,N_3574,N_4389);
or U8423 (N_8423,N_1914,N_204);
nor U8424 (N_8424,N_3220,N_573);
xnor U8425 (N_8425,N_334,N_4230);
xnor U8426 (N_8426,N_1324,N_2097);
or U8427 (N_8427,N_2161,N_673);
xnor U8428 (N_8428,N_4929,N_385);
or U8429 (N_8429,N_2771,N_37);
or U8430 (N_8430,N_1852,N_2823);
nand U8431 (N_8431,N_50,N_1737);
or U8432 (N_8432,N_4762,N_3165);
nand U8433 (N_8433,N_3004,N_3912);
nor U8434 (N_8434,N_4212,N_2392);
xnor U8435 (N_8435,N_2391,N_3139);
and U8436 (N_8436,N_1547,N_249);
nor U8437 (N_8437,N_383,N_2313);
xor U8438 (N_8438,N_3578,N_2738);
and U8439 (N_8439,N_4085,N_158);
xnor U8440 (N_8440,N_3577,N_4285);
xor U8441 (N_8441,N_600,N_1209);
and U8442 (N_8442,N_4548,N_228);
nand U8443 (N_8443,N_4579,N_1440);
xor U8444 (N_8444,N_2483,N_242);
or U8445 (N_8445,N_3523,N_3283);
and U8446 (N_8446,N_3803,N_4978);
nor U8447 (N_8447,N_950,N_1621);
and U8448 (N_8448,N_1990,N_3751);
nor U8449 (N_8449,N_3738,N_156);
nor U8450 (N_8450,N_1368,N_3358);
nor U8451 (N_8451,N_547,N_392);
nor U8452 (N_8452,N_2921,N_4729);
or U8453 (N_8453,N_4325,N_4725);
xnor U8454 (N_8454,N_3332,N_1323);
or U8455 (N_8455,N_3386,N_2738);
nand U8456 (N_8456,N_2562,N_1250);
nand U8457 (N_8457,N_3168,N_2263);
nor U8458 (N_8458,N_2064,N_970);
xnor U8459 (N_8459,N_2329,N_255);
and U8460 (N_8460,N_1228,N_3349);
and U8461 (N_8461,N_2547,N_1321);
nand U8462 (N_8462,N_2428,N_2842);
xnor U8463 (N_8463,N_110,N_2578);
and U8464 (N_8464,N_700,N_2728);
or U8465 (N_8465,N_3909,N_3174);
and U8466 (N_8466,N_2835,N_669);
xnor U8467 (N_8467,N_1934,N_3028);
nor U8468 (N_8468,N_3257,N_4651);
nand U8469 (N_8469,N_4014,N_1464);
and U8470 (N_8470,N_1998,N_683);
xor U8471 (N_8471,N_4002,N_4526);
nand U8472 (N_8472,N_2497,N_4969);
or U8473 (N_8473,N_2522,N_3435);
and U8474 (N_8474,N_3177,N_1530);
or U8475 (N_8475,N_221,N_163);
xnor U8476 (N_8476,N_2559,N_664);
nand U8477 (N_8477,N_3922,N_3571);
xnor U8478 (N_8478,N_1210,N_3034);
or U8479 (N_8479,N_80,N_376);
nand U8480 (N_8480,N_63,N_4896);
xnor U8481 (N_8481,N_4183,N_2403);
and U8482 (N_8482,N_2642,N_1858);
and U8483 (N_8483,N_145,N_2659);
nand U8484 (N_8484,N_1910,N_1022);
xor U8485 (N_8485,N_2971,N_2542);
nor U8486 (N_8486,N_1212,N_2415);
nand U8487 (N_8487,N_4036,N_4599);
nor U8488 (N_8488,N_4294,N_4182);
nand U8489 (N_8489,N_1178,N_3441);
nand U8490 (N_8490,N_1051,N_764);
and U8491 (N_8491,N_1311,N_3774);
xnor U8492 (N_8492,N_3246,N_576);
and U8493 (N_8493,N_3645,N_3130);
xor U8494 (N_8494,N_579,N_4247);
xnor U8495 (N_8495,N_4025,N_1030);
xor U8496 (N_8496,N_3589,N_2737);
or U8497 (N_8497,N_2113,N_1073);
nand U8498 (N_8498,N_4234,N_4123);
xnor U8499 (N_8499,N_2205,N_2063);
and U8500 (N_8500,N_1304,N_2444);
nor U8501 (N_8501,N_4162,N_3568);
or U8502 (N_8502,N_2863,N_3309);
and U8503 (N_8503,N_3034,N_2217);
xnor U8504 (N_8504,N_3878,N_1356);
nor U8505 (N_8505,N_4227,N_1405);
nor U8506 (N_8506,N_235,N_3509);
nor U8507 (N_8507,N_4466,N_1420);
or U8508 (N_8508,N_367,N_3231);
or U8509 (N_8509,N_3667,N_3687);
or U8510 (N_8510,N_2192,N_4819);
or U8511 (N_8511,N_2286,N_1477);
nor U8512 (N_8512,N_2808,N_278);
nand U8513 (N_8513,N_2517,N_3100);
nor U8514 (N_8514,N_4495,N_2326);
and U8515 (N_8515,N_1897,N_887);
or U8516 (N_8516,N_2299,N_2585);
or U8517 (N_8517,N_4318,N_184);
and U8518 (N_8518,N_4635,N_1233);
nor U8519 (N_8519,N_4303,N_4);
and U8520 (N_8520,N_417,N_3679);
nor U8521 (N_8521,N_596,N_4967);
nand U8522 (N_8522,N_4298,N_4609);
nand U8523 (N_8523,N_1173,N_2286);
and U8524 (N_8524,N_1236,N_2676);
nor U8525 (N_8525,N_673,N_2670);
and U8526 (N_8526,N_4242,N_3944);
xor U8527 (N_8527,N_3030,N_2230);
nand U8528 (N_8528,N_4191,N_4149);
or U8529 (N_8529,N_4912,N_3549);
xnor U8530 (N_8530,N_183,N_4885);
nor U8531 (N_8531,N_2596,N_3533);
xor U8532 (N_8532,N_3871,N_2565);
xnor U8533 (N_8533,N_504,N_3829);
nor U8534 (N_8534,N_4443,N_2986);
and U8535 (N_8535,N_4934,N_1148);
or U8536 (N_8536,N_595,N_3600);
and U8537 (N_8537,N_2670,N_3716);
or U8538 (N_8538,N_1522,N_4541);
and U8539 (N_8539,N_4102,N_2820);
or U8540 (N_8540,N_1196,N_4195);
or U8541 (N_8541,N_111,N_502);
nand U8542 (N_8542,N_3446,N_3847);
and U8543 (N_8543,N_4625,N_1278);
and U8544 (N_8544,N_788,N_4377);
xnor U8545 (N_8545,N_2039,N_2718);
and U8546 (N_8546,N_3279,N_1001);
nand U8547 (N_8547,N_2543,N_682);
and U8548 (N_8548,N_1933,N_3799);
nand U8549 (N_8549,N_3641,N_3336);
and U8550 (N_8550,N_217,N_2775);
xor U8551 (N_8551,N_907,N_2992);
nor U8552 (N_8552,N_2610,N_3055);
or U8553 (N_8553,N_2420,N_938);
or U8554 (N_8554,N_964,N_3016);
or U8555 (N_8555,N_360,N_4254);
and U8556 (N_8556,N_2191,N_2522);
nor U8557 (N_8557,N_4442,N_3769);
nand U8558 (N_8558,N_3529,N_1751);
nand U8559 (N_8559,N_2538,N_4380);
xnor U8560 (N_8560,N_1139,N_4845);
nand U8561 (N_8561,N_4070,N_2323);
xor U8562 (N_8562,N_2536,N_3246);
nor U8563 (N_8563,N_3703,N_1887);
xnor U8564 (N_8564,N_3262,N_2635);
and U8565 (N_8565,N_36,N_1087);
and U8566 (N_8566,N_3422,N_4665);
nand U8567 (N_8567,N_178,N_1534);
or U8568 (N_8568,N_130,N_4331);
and U8569 (N_8569,N_4729,N_4163);
and U8570 (N_8570,N_1905,N_2297);
xnor U8571 (N_8571,N_3286,N_3078);
nor U8572 (N_8572,N_2045,N_2168);
and U8573 (N_8573,N_1582,N_3500);
nor U8574 (N_8574,N_2795,N_2752);
nor U8575 (N_8575,N_835,N_1804);
nor U8576 (N_8576,N_1383,N_3218);
xnor U8577 (N_8577,N_128,N_1690);
nand U8578 (N_8578,N_2916,N_1486);
nand U8579 (N_8579,N_393,N_1030);
xor U8580 (N_8580,N_46,N_4364);
nand U8581 (N_8581,N_2049,N_1875);
and U8582 (N_8582,N_2285,N_3254);
nor U8583 (N_8583,N_1822,N_85);
or U8584 (N_8584,N_1334,N_831);
nand U8585 (N_8585,N_4854,N_2909);
or U8586 (N_8586,N_1454,N_626);
nand U8587 (N_8587,N_4958,N_561);
xnor U8588 (N_8588,N_2854,N_4904);
and U8589 (N_8589,N_2241,N_4693);
xor U8590 (N_8590,N_1517,N_2962);
nor U8591 (N_8591,N_2038,N_321);
xor U8592 (N_8592,N_2480,N_4137);
nand U8593 (N_8593,N_1320,N_4825);
and U8594 (N_8594,N_3339,N_3479);
xor U8595 (N_8595,N_728,N_1275);
nor U8596 (N_8596,N_4092,N_2809);
nor U8597 (N_8597,N_3657,N_1326);
or U8598 (N_8598,N_1066,N_2588);
xor U8599 (N_8599,N_1270,N_1138);
nor U8600 (N_8600,N_2522,N_2486);
nand U8601 (N_8601,N_138,N_4112);
or U8602 (N_8602,N_166,N_854);
nor U8603 (N_8603,N_4555,N_1155);
nor U8604 (N_8604,N_869,N_2136);
or U8605 (N_8605,N_4632,N_739);
nand U8606 (N_8606,N_3986,N_1044);
and U8607 (N_8607,N_890,N_3241);
nand U8608 (N_8608,N_1968,N_1176);
or U8609 (N_8609,N_3051,N_2946);
nor U8610 (N_8610,N_191,N_2951);
and U8611 (N_8611,N_1894,N_864);
or U8612 (N_8612,N_1429,N_1953);
or U8613 (N_8613,N_4194,N_3535);
and U8614 (N_8614,N_453,N_1335);
nor U8615 (N_8615,N_1260,N_521);
xnor U8616 (N_8616,N_3490,N_2033);
or U8617 (N_8617,N_2642,N_4607);
and U8618 (N_8618,N_4849,N_2310);
or U8619 (N_8619,N_2882,N_2832);
xnor U8620 (N_8620,N_3567,N_4538);
xnor U8621 (N_8621,N_844,N_3858);
nand U8622 (N_8622,N_3617,N_4738);
nand U8623 (N_8623,N_3949,N_3784);
nor U8624 (N_8624,N_3847,N_598);
nor U8625 (N_8625,N_898,N_445);
and U8626 (N_8626,N_4438,N_1626);
or U8627 (N_8627,N_2313,N_4440);
nand U8628 (N_8628,N_830,N_1192);
or U8629 (N_8629,N_714,N_3482);
or U8630 (N_8630,N_1066,N_375);
nor U8631 (N_8631,N_2076,N_143);
nor U8632 (N_8632,N_2015,N_4165);
or U8633 (N_8633,N_3226,N_3952);
nor U8634 (N_8634,N_1609,N_4235);
or U8635 (N_8635,N_4634,N_153);
and U8636 (N_8636,N_581,N_4338);
and U8637 (N_8637,N_3487,N_4192);
and U8638 (N_8638,N_2374,N_3567);
xnor U8639 (N_8639,N_2859,N_2575);
nand U8640 (N_8640,N_612,N_3782);
xor U8641 (N_8641,N_1073,N_499);
or U8642 (N_8642,N_204,N_2091);
and U8643 (N_8643,N_45,N_947);
nand U8644 (N_8644,N_3306,N_477);
xor U8645 (N_8645,N_2256,N_3306);
nor U8646 (N_8646,N_1157,N_3678);
or U8647 (N_8647,N_429,N_2173);
nor U8648 (N_8648,N_848,N_2815);
nor U8649 (N_8649,N_4435,N_1060);
and U8650 (N_8650,N_565,N_2231);
nand U8651 (N_8651,N_3339,N_2141);
xnor U8652 (N_8652,N_418,N_4992);
nand U8653 (N_8653,N_80,N_561);
nor U8654 (N_8654,N_3835,N_3031);
xnor U8655 (N_8655,N_1796,N_4605);
and U8656 (N_8656,N_3399,N_4962);
nor U8657 (N_8657,N_3078,N_312);
or U8658 (N_8658,N_3459,N_4285);
or U8659 (N_8659,N_3465,N_2185);
and U8660 (N_8660,N_1831,N_3417);
or U8661 (N_8661,N_749,N_892);
or U8662 (N_8662,N_1981,N_574);
nor U8663 (N_8663,N_4350,N_2715);
xor U8664 (N_8664,N_4327,N_4630);
and U8665 (N_8665,N_793,N_3194);
or U8666 (N_8666,N_2331,N_2624);
nand U8667 (N_8667,N_692,N_987);
or U8668 (N_8668,N_298,N_1776);
and U8669 (N_8669,N_3939,N_2702);
and U8670 (N_8670,N_404,N_4888);
and U8671 (N_8671,N_4147,N_2000);
and U8672 (N_8672,N_2618,N_4924);
and U8673 (N_8673,N_3820,N_3246);
nor U8674 (N_8674,N_166,N_4412);
nand U8675 (N_8675,N_4514,N_4638);
or U8676 (N_8676,N_1316,N_3743);
nand U8677 (N_8677,N_4674,N_4634);
xor U8678 (N_8678,N_4854,N_3790);
nor U8679 (N_8679,N_4694,N_498);
nand U8680 (N_8680,N_2469,N_766);
and U8681 (N_8681,N_1818,N_2742);
and U8682 (N_8682,N_2137,N_1006);
and U8683 (N_8683,N_3229,N_2399);
nor U8684 (N_8684,N_4090,N_3696);
nor U8685 (N_8685,N_3882,N_1312);
or U8686 (N_8686,N_1896,N_3201);
or U8687 (N_8687,N_3530,N_2962);
or U8688 (N_8688,N_1738,N_392);
xnor U8689 (N_8689,N_3944,N_2135);
and U8690 (N_8690,N_4332,N_4902);
xnor U8691 (N_8691,N_893,N_1231);
or U8692 (N_8692,N_2262,N_2776);
xnor U8693 (N_8693,N_4205,N_1115);
and U8694 (N_8694,N_962,N_2007);
nor U8695 (N_8695,N_2860,N_3442);
xnor U8696 (N_8696,N_4241,N_1102);
nor U8697 (N_8697,N_1662,N_86);
nor U8698 (N_8698,N_4054,N_1290);
nand U8699 (N_8699,N_4984,N_2139);
or U8700 (N_8700,N_3753,N_3746);
xnor U8701 (N_8701,N_1158,N_1876);
nor U8702 (N_8702,N_2369,N_4907);
nand U8703 (N_8703,N_4308,N_2411);
and U8704 (N_8704,N_3155,N_2042);
nor U8705 (N_8705,N_2122,N_595);
nand U8706 (N_8706,N_2365,N_309);
nor U8707 (N_8707,N_3446,N_4308);
or U8708 (N_8708,N_870,N_232);
nand U8709 (N_8709,N_4729,N_101);
xor U8710 (N_8710,N_2563,N_4421);
or U8711 (N_8711,N_112,N_2305);
nand U8712 (N_8712,N_2259,N_2919);
nor U8713 (N_8713,N_4531,N_1699);
xor U8714 (N_8714,N_3658,N_3116);
nor U8715 (N_8715,N_956,N_885);
nor U8716 (N_8716,N_180,N_4280);
xnor U8717 (N_8717,N_2807,N_304);
nand U8718 (N_8718,N_1675,N_952);
nor U8719 (N_8719,N_2500,N_1682);
xnor U8720 (N_8720,N_1219,N_2751);
or U8721 (N_8721,N_1183,N_3402);
nor U8722 (N_8722,N_4379,N_2793);
or U8723 (N_8723,N_3265,N_271);
or U8724 (N_8724,N_1916,N_4343);
or U8725 (N_8725,N_1024,N_4119);
nand U8726 (N_8726,N_4879,N_309);
nor U8727 (N_8727,N_3253,N_4977);
xnor U8728 (N_8728,N_4439,N_315);
nor U8729 (N_8729,N_4480,N_2782);
nand U8730 (N_8730,N_2148,N_3788);
nor U8731 (N_8731,N_2826,N_4096);
or U8732 (N_8732,N_1097,N_4431);
or U8733 (N_8733,N_1769,N_4302);
nand U8734 (N_8734,N_1087,N_2749);
or U8735 (N_8735,N_2668,N_3669);
and U8736 (N_8736,N_3212,N_570);
or U8737 (N_8737,N_4022,N_2287);
or U8738 (N_8738,N_1977,N_1203);
nand U8739 (N_8739,N_1639,N_4723);
nand U8740 (N_8740,N_720,N_3401);
and U8741 (N_8741,N_4198,N_4068);
nand U8742 (N_8742,N_4275,N_119);
xnor U8743 (N_8743,N_3692,N_4040);
nor U8744 (N_8744,N_4809,N_4252);
xor U8745 (N_8745,N_2419,N_2999);
nand U8746 (N_8746,N_4191,N_3652);
xnor U8747 (N_8747,N_2513,N_2682);
or U8748 (N_8748,N_2795,N_4353);
xnor U8749 (N_8749,N_2421,N_3811);
or U8750 (N_8750,N_1767,N_2403);
nand U8751 (N_8751,N_4741,N_2730);
xor U8752 (N_8752,N_4354,N_1704);
nor U8753 (N_8753,N_1761,N_4818);
nand U8754 (N_8754,N_267,N_777);
nor U8755 (N_8755,N_2600,N_4563);
and U8756 (N_8756,N_3755,N_967);
nand U8757 (N_8757,N_4379,N_2277);
xor U8758 (N_8758,N_2462,N_3153);
and U8759 (N_8759,N_355,N_4502);
nand U8760 (N_8760,N_819,N_737);
and U8761 (N_8761,N_114,N_2981);
or U8762 (N_8762,N_3278,N_1903);
xor U8763 (N_8763,N_4374,N_2389);
or U8764 (N_8764,N_4078,N_2323);
nand U8765 (N_8765,N_2082,N_4763);
nor U8766 (N_8766,N_3090,N_4858);
nand U8767 (N_8767,N_1761,N_3529);
xor U8768 (N_8768,N_2743,N_1901);
nand U8769 (N_8769,N_1347,N_1790);
and U8770 (N_8770,N_156,N_1187);
xor U8771 (N_8771,N_3375,N_1624);
xnor U8772 (N_8772,N_4500,N_2487);
nand U8773 (N_8773,N_2203,N_1660);
xnor U8774 (N_8774,N_1384,N_3614);
or U8775 (N_8775,N_836,N_2714);
and U8776 (N_8776,N_1298,N_2356);
nor U8777 (N_8777,N_4882,N_4932);
nor U8778 (N_8778,N_650,N_255);
xnor U8779 (N_8779,N_1620,N_3263);
or U8780 (N_8780,N_3678,N_2848);
xnor U8781 (N_8781,N_4885,N_3521);
xnor U8782 (N_8782,N_1591,N_714);
nand U8783 (N_8783,N_2013,N_3602);
and U8784 (N_8784,N_2913,N_1094);
nor U8785 (N_8785,N_1448,N_4565);
nand U8786 (N_8786,N_46,N_1238);
xnor U8787 (N_8787,N_2646,N_3303);
and U8788 (N_8788,N_4718,N_1923);
and U8789 (N_8789,N_1314,N_2600);
and U8790 (N_8790,N_2172,N_7);
nor U8791 (N_8791,N_2701,N_1962);
xnor U8792 (N_8792,N_3550,N_1671);
or U8793 (N_8793,N_2137,N_4964);
nand U8794 (N_8794,N_3829,N_3741);
and U8795 (N_8795,N_3107,N_2489);
xor U8796 (N_8796,N_1039,N_4981);
nand U8797 (N_8797,N_3107,N_1130);
nor U8798 (N_8798,N_1872,N_1195);
xor U8799 (N_8799,N_1414,N_3720);
xor U8800 (N_8800,N_3211,N_1092);
nand U8801 (N_8801,N_2936,N_3334);
nand U8802 (N_8802,N_2125,N_1328);
or U8803 (N_8803,N_1137,N_225);
nor U8804 (N_8804,N_2166,N_60);
and U8805 (N_8805,N_619,N_938);
xor U8806 (N_8806,N_220,N_3571);
nand U8807 (N_8807,N_1583,N_719);
nor U8808 (N_8808,N_71,N_1185);
nand U8809 (N_8809,N_2109,N_1546);
xor U8810 (N_8810,N_1549,N_3421);
nor U8811 (N_8811,N_1483,N_2536);
nor U8812 (N_8812,N_1729,N_227);
nand U8813 (N_8813,N_2923,N_2193);
or U8814 (N_8814,N_1680,N_4365);
and U8815 (N_8815,N_4198,N_146);
and U8816 (N_8816,N_1569,N_3727);
nand U8817 (N_8817,N_4008,N_2277);
or U8818 (N_8818,N_144,N_4846);
or U8819 (N_8819,N_1225,N_3860);
xor U8820 (N_8820,N_1429,N_2210);
or U8821 (N_8821,N_60,N_4245);
or U8822 (N_8822,N_1857,N_651);
or U8823 (N_8823,N_4131,N_2507);
or U8824 (N_8824,N_2869,N_3867);
or U8825 (N_8825,N_591,N_3721);
nor U8826 (N_8826,N_929,N_1921);
nand U8827 (N_8827,N_3298,N_2966);
and U8828 (N_8828,N_3742,N_2979);
nor U8829 (N_8829,N_2601,N_4757);
xnor U8830 (N_8830,N_1854,N_193);
nand U8831 (N_8831,N_228,N_4737);
nor U8832 (N_8832,N_2116,N_3574);
nor U8833 (N_8833,N_3609,N_2731);
nand U8834 (N_8834,N_4598,N_4711);
nor U8835 (N_8835,N_3357,N_2244);
or U8836 (N_8836,N_2506,N_3350);
and U8837 (N_8837,N_845,N_355);
nor U8838 (N_8838,N_2773,N_587);
and U8839 (N_8839,N_3148,N_2935);
and U8840 (N_8840,N_3366,N_1889);
nand U8841 (N_8841,N_3059,N_2568);
xor U8842 (N_8842,N_4491,N_1829);
nand U8843 (N_8843,N_1344,N_3883);
nand U8844 (N_8844,N_2811,N_1913);
nor U8845 (N_8845,N_4110,N_2008);
or U8846 (N_8846,N_2910,N_3594);
or U8847 (N_8847,N_970,N_3032);
nand U8848 (N_8848,N_3501,N_2537);
and U8849 (N_8849,N_4803,N_683);
nand U8850 (N_8850,N_719,N_2172);
nand U8851 (N_8851,N_3167,N_4193);
nand U8852 (N_8852,N_4131,N_2235);
xor U8853 (N_8853,N_3891,N_4368);
and U8854 (N_8854,N_4810,N_485);
nand U8855 (N_8855,N_2850,N_2236);
xor U8856 (N_8856,N_1965,N_948);
or U8857 (N_8857,N_3770,N_4895);
or U8858 (N_8858,N_203,N_495);
nor U8859 (N_8859,N_4648,N_2668);
and U8860 (N_8860,N_4451,N_1134);
or U8861 (N_8861,N_1879,N_2442);
nor U8862 (N_8862,N_271,N_4858);
nand U8863 (N_8863,N_3818,N_4959);
nor U8864 (N_8864,N_4640,N_2245);
and U8865 (N_8865,N_4441,N_4418);
and U8866 (N_8866,N_3589,N_2590);
nor U8867 (N_8867,N_655,N_4843);
xor U8868 (N_8868,N_4262,N_3394);
nand U8869 (N_8869,N_1780,N_857);
nand U8870 (N_8870,N_3949,N_4218);
nand U8871 (N_8871,N_4758,N_310);
nor U8872 (N_8872,N_2263,N_753);
nand U8873 (N_8873,N_2129,N_3634);
nand U8874 (N_8874,N_721,N_4906);
and U8875 (N_8875,N_4244,N_979);
nand U8876 (N_8876,N_1441,N_2989);
xor U8877 (N_8877,N_196,N_4249);
nor U8878 (N_8878,N_713,N_709);
nor U8879 (N_8879,N_627,N_3028);
nand U8880 (N_8880,N_487,N_731);
xor U8881 (N_8881,N_886,N_1773);
xnor U8882 (N_8882,N_3644,N_115);
nor U8883 (N_8883,N_3356,N_2510);
and U8884 (N_8884,N_1543,N_1456);
xor U8885 (N_8885,N_2990,N_2842);
xor U8886 (N_8886,N_3337,N_4119);
and U8887 (N_8887,N_4657,N_4734);
nand U8888 (N_8888,N_1133,N_2282);
nor U8889 (N_8889,N_2795,N_3337);
nor U8890 (N_8890,N_782,N_3798);
nor U8891 (N_8891,N_4375,N_4636);
or U8892 (N_8892,N_4897,N_4058);
nand U8893 (N_8893,N_740,N_2272);
or U8894 (N_8894,N_3332,N_1134);
and U8895 (N_8895,N_2367,N_3156);
nor U8896 (N_8896,N_4473,N_2092);
nand U8897 (N_8897,N_1357,N_849);
nand U8898 (N_8898,N_2367,N_4649);
nand U8899 (N_8899,N_4657,N_3917);
or U8900 (N_8900,N_3221,N_1442);
nor U8901 (N_8901,N_4962,N_3362);
and U8902 (N_8902,N_4948,N_4058);
nand U8903 (N_8903,N_370,N_2310);
xnor U8904 (N_8904,N_3068,N_2594);
and U8905 (N_8905,N_3835,N_1039);
and U8906 (N_8906,N_1767,N_4627);
and U8907 (N_8907,N_3368,N_3409);
nor U8908 (N_8908,N_173,N_4032);
nand U8909 (N_8909,N_1166,N_3979);
nand U8910 (N_8910,N_255,N_3813);
xnor U8911 (N_8911,N_1037,N_1198);
nor U8912 (N_8912,N_443,N_4788);
nor U8913 (N_8913,N_3348,N_2345);
nand U8914 (N_8914,N_3115,N_3242);
nor U8915 (N_8915,N_1721,N_1863);
xnor U8916 (N_8916,N_4151,N_3527);
xor U8917 (N_8917,N_492,N_4607);
nor U8918 (N_8918,N_167,N_57);
or U8919 (N_8919,N_2799,N_4271);
or U8920 (N_8920,N_3370,N_187);
xnor U8921 (N_8921,N_719,N_1178);
nor U8922 (N_8922,N_4700,N_2249);
xor U8923 (N_8923,N_3986,N_976);
xor U8924 (N_8924,N_3541,N_3597);
xor U8925 (N_8925,N_2117,N_1418);
or U8926 (N_8926,N_460,N_4400);
or U8927 (N_8927,N_766,N_3835);
and U8928 (N_8928,N_1205,N_2703);
xor U8929 (N_8929,N_2907,N_4475);
or U8930 (N_8930,N_4011,N_1215);
and U8931 (N_8931,N_543,N_2912);
and U8932 (N_8932,N_4005,N_3352);
or U8933 (N_8933,N_2694,N_3742);
or U8934 (N_8934,N_2741,N_2422);
or U8935 (N_8935,N_3249,N_1772);
nor U8936 (N_8936,N_3977,N_2502);
xor U8937 (N_8937,N_1491,N_1591);
or U8938 (N_8938,N_3714,N_3874);
and U8939 (N_8939,N_4226,N_407);
and U8940 (N_8940,N_1145,N_29);
nor U8941 (N_8941,N_3134,N_4700);
or U8942 (N_8942,N_2221,N_2397);
or U8943 (N_8943,N_4196,N_4905);
nand U8944 (N_8944,N_2688,N_28);
or U8945 (N_8945,N_3865,N_973);
nor U8946 (N_8946,N_714,N_1779);
xor U8947 (N_8947,N_4808,N_3988);
and U8948 (N_8948,N_329,N_3184);
or U8949 (N_8949,N_2425,N_1006);
and U8950 (N_8950,N_4617,N_3660);
nand U8951 (N_8951,N_2103,N_655);
xnor U8952 (N_8952,N_698,N_940);
nor U8953 (N_8953,N_2155,N_666);
or U8954 (N_8954,N_1755,N_202);
xnor U8955 (N_8955,N_2017,N_1641);
nor U8956 (N_8956,N_112,N_4338);
nor U8957 (N_8957,N_4780,N_3526);
nand U8958 (N_8958,N_2734,N_1199);
xor U8959 (N_8959,N_3102,N_4159);
nand U8960 (N_8960,N_2170,N_1705);
nor U8961 (N_8961,N_2362,N_4559);
nor U8962 (N_8962,N_3599,N_1138);
nand U8963 (N_8963,N_1244,N_4807);
and U8964 (N_8964,N_1801,N_4548);
nor U8965 (N_8965,N_4184,N_708);
and U8966 (N_8966,N_697,N_4732);
nor U8967 (N_8967,N_1126,N_3817);
or U8968 (N_8968,N_2393,N_655);
or U8969 (N_8969,N_2229,N_4698);
xnor U8970 (N_8970,N_2988,N_4557);
and U8971 (N_8971,N_860,N_1930);
nor U8972 (N_8972,N_516,N_64);
or U8973 (N_8973,N_321,N_373);
nor U8974 (N_8974,N_330,N_2668);
or U8975 (N_8975,N_4475,N_4356);
nand U8976 (N_8976,N_4703,N_2829);
and U8977 (N_8977,N_1693,N_4913);
nand U8978 (N_8978,N_2768,N_4058);
xnor U8979 (N_8979,N_824,N_1744);
nand U8980 (N_8980,N_2670,N_3123);
or U8981 (N_8981,N_1305,N_3142);
and U8982 (N_8982,N_2000,N_4920);
nor U8983 (N_8983,N_1279,N_2996);
or U8984 (N_8984,N_1357,N_2468);
and U8985 (N_8985,N_4754,N_4278);
nand U8986 (N_8986,N_3343,N_2280);
nand U8987 (N_8987,N_3272,N_3423);
or U8988 (N_8988,N_2262,N_2810);
nand U8989 (N_8989,N_523,N_3869);
xor U8990 (N_8990,N_839,N_209);
nand U8991 (N_8991,N_529,N_135);
nor U8992 (N_8992,N_390,N_2965);
nor U8993 (N_8993,N_3705,N_4164);
or U8994 (N_8994,N_1348,N_3548);
xor U8995 (N_8995,N_4909,N_4035);
nor U8996 (N_8996,N_574,N_3508);
and U8997 (N_8997,N_969,N_2591);
xnor U8998 (N_8998,N_1014,N_1356);
nand U8999 (N_8999,N_3081,N_4987);
xor U9000 (N_9000,N_500,N_3872);
and U9001 (N_9001,N_4615,N_4745);
nand U9002 (N_9002,N_3358,N_1640);
xnor U9003 (N_9003,N_376,N_3448);
nor U9004 (N_9004,N_3670,N_1190);
xor U9005 (N_9005,N_4882,N_374);
and U9006 (N_9006,N_2779,N_459);
nor U9007 (N_9007,N_4984,N_777);
nand U9008 (N_9008,N_2717,N_2486);
or U9009 (N_9009,N_2793,N_699);
and U9010 (N_9010,N_4228,N_3086);
or U9011 (N_9011,N_2163,N_4994);
nor U9012 (N_9012,N_3919,N_813);
and U9013 (N_9013,N_1170,N_4879);
and U9014 (N_9014,N_3086,N_1786);
xor U9015 (N_9015,N_1328,N_606);
nor U9016 (N_9016,N_196,N_882);
xor U9017 (N_9017,N_2629,N_1409);
nor U9018 (N_9018,N_682,N_3387);
nand U9019 (N_9019,N_634,N_1327);
nand U9020 (N_9020,N_3210,N_2560);
and U9021 (N_9021,N_2883,N_2431);
xor U9022 (N_9022,N_3900,N_4886);
nor U9023 (N_9023,N_3733,N_2731);
or U9024 (N_9024,N_3908,N_539);
nor U9025 (N_9025,N_2849,N_4037);
xnor U9026 (N_9026,N_2244,N_344);
nand U9027 (N_9027,N_4990,N_761);
or U9028 (N_9028,N_543,N_4270);
or U9029 (N_9029,N_3854,N_964);
and U9030 (N_9030,N_1365,N_2830);
or U9031 (N_9031,N_4418,N_2011);
and U9032 (N_9032,N_2536,N_1856);
xnor U9033 (N_9033,N_995,N_2879);
or U9034 (N_9034,N_659,N_4283);
xnor U9035 (N_9035,N_3454,N_147);
and U9036 (N_9036,N_95,N_2749);
nor U9037 (N_9037,N_4309,N_1213);
and U9038 (N_9038,N_2009,N_3821);
or U9039 (N_9039,N_354,N_4070);
xnor U9040 (N_9040,N_1331,N_4329);
nand U9041 (N_9041,N_4803,N_1481);
nand U9042 (N_9042,N_4828,N_2378);
or U9043 (N_9043,N_3259,N_1720);
and U9044 (N_9044,N_973,N_3160);
or U9045 (N_9045,N_2117,N_4779);
and U9046 (N_9046,N_1385,N_2883);
or U9047 (N_9047,N_2609,N_2851);
or U9048 (N_9048,N_50,N_2966);
or U9049 (N_9049,N_2759,N_250);
nand U9050 (N_9050,N_3942,N_3320);
nor U9051 (N_9051,N_1897,N_3428);
or U9052 (N_9052,N_368,N_1108);
nand U9053 (N_9053,N_2043,N_31);
or U9054 (N_9054,N_1459,N_4065);
xor U9055 (N_9055,N_3320,N_243);
and U9056 (N_9056,N_2081,N_3267);
nor U9057 (N_9057,N_463,N_326);
nor U9058 (N_9058,N_2470,N_3183);
or U9059 (N_9059,N_4651,N_4460);
or U9060 (N_9060,N_575,N_3269);
and U9061 (N_9061,N_2522,N_3921);
and U9062 (N_9062,N_782,N_2821);
xnor U9063 (N_9063,N_4955,N_261);
nand U9064 (N_9064,N_3396,N_2589);
and U9065 (N_9065,N_2876,N_3125);
and U9066 (N_9066,N_4411,N_415);
nor U9067 (N_9067,N_606,N_3182);
nor U9068 (N_9068,N_1672,N_3949);
nand U9069 (N_9069,N_340,N_176);
or U9070 (N_9070,N_608,N_4395);
xnor U9071 (N_9071,N_2306,N_4401);
nor U9072 (N_9072,N_3600,N_4359);
and U9073 (N_9073,N_3432,N_163);
and U9074 (N_9074,N_2634,N_399);
nor U9075 (N_9075,N_896,N_1787);
or U9076 (N_9076,N_1902,N_4367);
nand U9077 (N_9077,N_3607,N_4127);
xor U9078 (N_9078,N_1209,N_3995);
and U9079 (N_9079,N_2441,N_2247);
or U9080 (N_9080,N_4499,N_1304);
xnor U9081 (N_9081,N_3031,N_3233);
or U9082 (N_9082,N_3422,N_67);
nand U9083 (N_9083,N_2885,N_2063);
xnor U9084 (N_9084,N_1265,N_285);
nor U9085 (N_9085,N_1877,N_1214);
or U9086 (N_9086,N_2700,N_548);
or U9087 (N_9087,N_1593,N_522);
or U9088 (N_9088,N_1542,N_551);
nor U9089 (N_9089,N_4050,N_1679);
nor U9090 (N_9090,N_3042,N_4721);
nand U9091 (N_9091,N_4377,N_4488);
or U9092 (N_9092,N_3536,N_3362);
or U9093 (N_9093,N_1209,N_2634);
nor U9094 (N_9094,N_4599,N_4987);
nand U9095 (N_9095,N_4162,N_3187);
or U9096 (N_9096,N_1877,N_1946);
xor U9097 (N_9097,N_3398,N_4127);
and U9098 (N_9098,N_1907,N_4524);
nand U9099 (N_9099,N_1280,N_2424);
nand U9100 (N_9100,N_4970,N_852);
and U9101 (N_9101,N_4469,N_1570);
and U9102 (N_9102,N_3325,N_678);
nand U9103 (N_9103,N_2061,N_3202);
or U9104 (N_9104,N_4564,N_809);
nor U9105 (N_9105,N_4245,N_3916);
nand U9106 (N_9106,N_4289,N_4337);
xor U9107 (N_9107,N_2718,N_1162);
and U9108 (N_9108,N_2599,N_4636);
and U9109 (N_9109,N_404,N_4995);
or U9110 (N_9110,N_4127,N_787);
nand U9111 (N_9111,N_956,N_4989);
xnor U9112 (N_9112,N_2452,N_1295);
xnor U9113 (N_9113,N_2105,N_1922);
nor U9114 (N_9114,N_1749,N_2295);
xor U9115 (N_9115,N_1928,N_1347);
nand U9116 (N_9116,N_675,N_1837);
and U9117 (N_9117,N_3216,N_3912);
nand U9118 (N_9118,N_3321,N_3774);
or U9119 (N_9119,N_2386,N_4583);
nor U9120 (N_9120,N_4936,N_1245);
or U9121 (N_9121,N_1331,N_4941);
nand U9122 (N_9122,N_1623,N_4019);
nand U9123 (N_9123,N_292,N_1130);
nand U9124 (N_9124,N_1671,N_50);
or U9125 (N_9125,N_2141,N_2958);
nor U9126 (N_9126,N_2346,N_498);
xor U9127 (N_9127,N_107,N_458);
xnor U9128 (N_9128,N_1950,N_2682);
or U9129 (N_9129,N_1537,N_3422);
and U9130 (N_9130,N_1628,N_2357);
nand U9131 (N_9131,N_4401,N_3217);
nand U9132 (N_9132,N_3209,N_3003);
or U9133 (N_9133,N_4389,N_2603);
and U9134 (N_9134,N_2885,N_1162);
and U9135 (N_9135,N_1799,N_3891);
xor U9136 (N_9136,N_654,N_56);
and U9137 (N_9137,N_3214,N_2023);
or U9138 (N_9138,N_3300,N_2361);
xnor U9139 (N_9139,N_3925,N_1543);
and U9140 (N_9140,N_273,N_441);
nand U9141 (N_9141,N_1941,N_895);
xor U9142 (N_9142,N_2514,N_2531);
nand U9143 (N_9143,N_1229,N_4288);
and U9144 (N_9144,N_2353,N_1508);
or U9145 (N_9145,N_1736,N_2760);
nor U9146 (N_9146,N_4533,N_863);
nor U9147 (N_9147,N_3438,N_3657);
nor U9148 (N_9148,N_4588,N_1101);
nand U9149 (N_9149,N_4680,N_3257);
xor U9150 (N_9150,N_1435,N_4547);
and U9151 (N_9151,N_4903,N_3033);
nand U9152 (N_9152,N_1588,N_3486);
xor U9153 (N_9153,N_2266,N_200);
nand U9154 (N_9154,N_2095,N_370);
nand U9155 (N_9155,N_3556,N_4663);
nor U9156 (N_9156,N_4896,N_2571);
nand U9157 (N_9157,N_3246,N_2240);
xnor U9158 (N_9158,N_848,N_4380);
and U9159 (N_9159,N_2199,N_3753);
xnor U9160 (N_9160,N_1518,N_4385);
and U9161 (N_9161,N_227,N_4560);
and U9162 (N_9162,N_4469,N_3085);
nor U9163 (N_9163,N_3093,N_4700);
or U9164 (N_9164,N_2577,N_4729);
nand U9165 (N_9165,N_3005,N_4921);
nand U9166 (N_9166,N_2087,N_2606);
nor U9167 (N_9167,N_1835,N_1083);
and U9168 (N_9168,N_554,N_1335);
and U9169 (N_9169,N_4110,N_2103);
xor U9170 (N_9170,N_4881,N_3971);
xnor U9171 (N_9171,N_4365,N_3423);
nor U9172 (N_9172,N_402,N_3238);
and U9173 (N_9173,N_801,N_4042);
and U9174 (N_9174,N_3030,N_2149);
xor U9175 (N_9175,N_2802,N_3879);
and U9176 (N_9176,N_2965,N_4626);
nand U9177 (N_9177,N_3145,N_3452);
nor U9178 (N_9178,N_3352,N_1283);
and U9179 (N_9179,N_1800,N_155);
nor U9180 (N_9180,N_726,N_3928);
or U9181 (N_9181,N_2700,N_3346);
nor U9182 (N_9182,N_3537,N_673);
or U9183 (N_9183,N_1024,N_1888);
or U9184 (N_9184,N_2332,N_3486);
or U9185 (N_9185,N_3590,N_167);
or U9186 (N_9186,N_1242,N_4788);
nand U9187 (N_9187,N_3362,N_3843);
or U9188 (N_9188,N_3868,N_2059);
nor U9189 (N_9189,N_2742,N_2020);
or U9190 (N_9190,N_52,N_2545);
nor U9191 (N_9191,N_3072,N_3527);
xor U9192 (N_9192,N_4945,N_711);
nor U9193 (N_9193,N_2409,N_2965);
or U9194 (N_9194,N_383,N_916);
or U9195 (N_9195,N_2872,N_408);
and U9196 (N_9196,N_951,N_1932);
or U9197 (N_9197,N_3665,N_4655);
nand U9198 (N_9198,N_1910,N_1803);
nor U9199 (N_9199,N_1080,N_4001);
xnor U9200 (N_9200,N_513,N_4944);
xor U9201 (N_9201,N_2841,N_2759);
nand U9202 (N_9202,N_3789,N_4009);
xnor U9203 (N_9203,N_2409,N_3959);
nand U9204 (N_9204,N_433,N_2264);
nor U9205 (N_9205,N_1854,N_2381);
nor U9206 (N_9206,N_2905,N_4458);
and U9207 (N_9207,N_3066,N_1326);
and U9208 (N_9208,N_4002,N_4998);
or U9209 (N_9209,N_3870,N_4379);
nand U9210 (N_9210,N_2003,N_903);
nand U9211 (N_9211,N_2687,N_1437);
or U9212 (N_9212,N_3772,N_1363);
nand U9213 (N_9213,N_3498,N_2467);
nand U9214 (N_9214,N_377,N_2216);
nand U9215 (N_9215,N_3222,N_4396);
and U9216 (N_9216,N_3578,N_2258);
and U9217 (N_9217,N_1419,N_1567);
nand U9218 (N_9218,N_2062,N_2233);
and U9219 (N_9219,N_3078,N_502);
or U9220 (N_9220,N_464,N_2948);
and U9221 (N_9221,N_3081,N_15);
xnor U9222 (N_9222,N_977,N_1250);
xnor U9223 (N_9223,N_2324,N_3698);
and U9224 (N_9224,N_4244,N_2711);
or U9225 (N_9225,N_2375,N_3227);
nor U9226 (N_9226,N_599,N_1785);
and U9227 (N_9227,N_106,N_1540);
nor U9228 (N_9228,N_4474,N_3885);
and U9229 (N_9229,N_1688,N_600);
nor U9230 (N_9230,N_686,N_2991);
nand U9231 (N_9231,N_3407,N_4165);
and U9232 (N_9232,N_329,N_3225);
and U9233 (N_9233,N_664,N_969);
nor U9234 (N_9234,N_2484,N_0);
nand U9235 (N_9235,N_1633,N_3240);
nor U9236 (N_9236,N_2988,N_2149);
and U9237 (N_9237,N_844,N_1713);
nor U9238 (N_9238,N_3782,N_167);
xnor U9239 (N_9239,N_2182,N_3019);
nor U9240 (N_9240,N_1502,N_3047);
nor U9241 (N_9241,N_1432,N_4105);
nor U9242 (N_9242,N_1507,N_4732);
or U9243 (N_9243,N_4010,N_368);
xor U9244 (N_9244,N_2829,N_3745);
nand U9245 (N_9245,N_3090,N_2207);
nor U9246 (N_9246,N_4035,N_4995);
and U9247 (N_9247,N_3931,N_2157);
xor U9248 (N_9248,N_528,N_3940);
nand U9249 (N_9249,N_1865,N_1325);
nor U9250 (N_9250,N_4241,N_654);
nor U9251 (N_9251,N_2530,N_461);
or U9252 (N_9252,N_988,N_4245);
and U9253 (N_9253,N_3014,N_1721);
xor U9254 (N_9254,N_3777,N_3194);
nor U9255 (N_9255,N_1201,N_4283);
xor U9256 (N_9256,N_3280,N_2519);
nand U9257 (N_9257,N_4289,N_4954);
nor U9258 (N_9258,N_2784,N_4562);
nand U9259 (N_9259,N_553,N_1469);
nand U9260 (N_9260,N_1421,N_2714);
xor U9261 (N_9261,N_3083,N_1948);
or U9262 (N_9262,N_3976,N_437);
nand U9263 (N_9263,N_65,N_4964);
or U9264 (N_9264,N_2993,N_3580);
nor U9265 (N_9265,N_3569,N_2141);
nor U9266 (N_9266,N_1842,N_4670);
xor U9267 (N_9267,N_4597,N_3883);
nor U9268 (N_9268,N_4123,N_4441);
and U9269 (N_9269,N_4313,N_527);
nor U9270 (N_9270,N_4078,N_4331);
and U9271 (N_9271,N_2351,N_1907);
nor U9272 (N_9272,N_1386,N_3334);
or U9273 (N_9273,N_1102,N_1490);
nor U9274 (N_9274,N_4713,N_3538);
nor U9275 (N_9275,N_4555,N_840);
nor U9276 (N_9276,N_3856,N_1545);
and U9277 (N_9277,N_4244,N_4367);
nor U9278 (N_9278,N_3146,N_4057);
nor U9279 (N_9279,N_1449,N_1175);
nor U9280 (N_9280,N_1059,N_4605);
xor U9281 (N_9281,N_3907,N_2507);
nand U9282 (N_9282,N_1778,N_4010);
or U9283 (N_9283,N_1630,N_1571);
and U9284 (N_9284,N_4345,N_2513);
and U9285 (N_9285,N_4472,N_4210);
nor U9286 (N_9286,N_3637,N_3243);
nand U9287 (N_9287,N_115,N_2517);
xor U9288 (N_9288,N_849,N_2984);
and U9289 (N_9289,N_3488,N_2317);
xor U9290 (N_9290,N_1474,N_2368);
nor U9291 (N_9291,N_3450,N_333);
nor U9292 (N_9292,N_882,N_2727);
nand U9293 (N_9293,N_2819,N_1401);
nor U9294 (N_9294,N_3354,N_3702);
nand U9295 (N_9295,N_2757,N_3979);
and U9296 (N_9296,N_749,N_3400);
and U9297 (N_9297,N_1422,N_2254);
or U9298 (N_9298,N_2495,N_1405);
nand U9299 (N_9299,N_2382,N_4667);
and U9300 (N_9300,N_99,N_3306);
and U9301 (N_9301,N_3907,N_493);
nand U9302 (N_9302,N_1571,N_4435);
nor U9303 (N_9303,N_4940,N_4601);
and U9304 (N_9304,N_336,N_4938);
nand U9305 (N_9305,N_2429,N_2569);
nand U9306 (N_9306,N_3126,N_1375);
nand U9307 (N_9307,N_1278,N_4482);
xnor U9308 (N_9308,N_1803,N_3142);
or U9309 (N_9309,N_843,N_3642);
nand U9310 (N_9310,N_4258,N_968);
and U9311 (N_9311,N_1293,N_316);
xor U9312 (N_9312,N_260,N_2694);
xnor U9313 (N_9313,N_2973,N_2100);
and U9314 (N_9314,N_4965,N_3493);
and U9315 (N_9315,N_2792,N_4765);
nor U9316 (N_9316,N_85,N_3375);
nor U9317 (N_9317,N_3663,N_1829);
and U9318 (N_9318,N_853,N_2903);
nand U9319 (N_9319,N_18,N_3398);
nand U9320 (N_9320,N_1873,N_4501);
and U9321 (N_9321,N_3453,N_284);
or U9322 (N_9322,N_3560,N_4916);
or U9323 (N_9323,N_1867,N_2922);
and U9324 (N_9324,N_1589,N_4278);
and U9325 (N_9325,N_228,N_2644);
xnor U9326 (N_9326,N_4463,N_1621);
and U9327 (N_9327,N_708,N_1615);
and U9328 (N_9328,N_4619,N_1236);
nor U9329 (N_9329,N_3728,N_4404);
nor U9330 (N_9330,N_747,N_3793);
nor U9331 (N_9331,N_1618,N_2153);
xnor U9332 (N_9332,N_2507,N_1119);
nand U9333 (N_9333,N_3631,N_35);
and U9334 (N_9334,N_1227,N_2893);
or U9335 (N_9335,N_666,N_1006);
nand U9336 (N_9336,N_4291,N_2912);
or U9337 (N_9337,N_3818,N_3152);
xnor U9338 (N_9338,N_2096,N_1680);
nand U9339 (N_9339,N_2548,N_3652);
nor U9340 (N_9340,N_2691,N_2393);
or U9341 (N_9341,N_2819,N_3275);
nor U9342 (N_9342,N_2098,N_4610);
nand U9343 (N_9343,N_287,N_597);
or U9344 (N_9344,N_4034,N_3393);
and U9345 (N_9345,N_1152,N_2814);
nand U9346 (N_9346,N_2617,N_3021);
and U9347 (N_9347,N_3917,N_1968);
nor U9348 (N_9348,N_812,N_3533);
nor U9349 (N_9349,N_3924,N_2960);
or U9350 (N_9350,N_845,N_2500);
and U9351 (N_9351,N_661,N_2990);
nand U9352 (N_9352,N_4354,N_4335);
or U9353 (N_9353,N_4107,N_3081);
nand U9354 (N_9354,N_477,N_3648);
nand U9355 (N_9355,N_1932,N_1146);
nor U9356 (N_9356,N_4525,N_372);
nor U9357 (N_9357,N_3293,N_2832);
nor U9358 (N_9358,N_252,N_819);
or U9359 (N_9359,N_3506,N_2644);
and U9360 (N_9360,N_2867,N_3202);
nand U9361 (N_9361,N_377,N_3648);
xor U9362 (N_9362,N_2099,N_684);
nand U9363 (N_9363,N_4976,N_3776);
nor U9364 (N_9364,N_2636,N_509);
nand U9365 (N_9365,N_2388,N_3160);
and U9366 (N_9366,N_3990,N_3161);
nand U9367 (N_9367,N_2277,N_4178);
nor U9368 (N_9368,N_4949,N_4182);
or U9369 (N_9369,N_837,N_4638);
nand U9370 (N_9370,N_618,N_1788);
nand U9371 (N_9371,N_4459,N_3526);
nor U9372 (N_9372,N_2599,N_726);
and U9373 (N_9373,N_1318,N_767);
and U9374 (N_9374,N_1697,N_4672);
and U9375 (N_9375,N_1840,N_3652);
nor U9376 (N_9376,N_1064,N_598);
nor U9377 (N_9377,N_2154,N_1513);
or U9378 (N_9378,N_443,N_2369);
or U9379 (N_9379,N_2087,N_3944);
xnor U9380 (N_9380,N_1108,N_2112);
nand U9381 (N_9381,N_1960,N_4958);
nor U9382 (N_9382,N_3005,N_4990);
nand U9383 (N_9383,N_535,N_914);
or U9384 (N_9384,N_1624,N_507);
xnor U9385 (N_9385,N_1502,N_2687);
and U9386 (N_9386,N_2784,N_3399);
nand U9387 (N_9387,N_995,N_3976);
nand U9388 (N_9388,N_1832,N_789);
or U9389 (N_9389,N_2895,N_100);
xnor U9390 (N_9390,N_4694,N_2792);
nor U9391 (N_9391,N_3611,N_4385);
or U9392 (N_9392,N_4310,N_3572);
or U9393 (N_9393,N_4210,N_1061);
and U9394 (N_9394,N_2671,N_917);
xor U9395 (N_9395,N_1529,N_4935);
xnor U9396 (N_9396,N_3447,N_1391);
and U9397 (N_9397,N_4568,N_2207);
and U9398 (N_9398,N_1320,N_4359);
and U9399 (N_9399,N_3023,N_2237);
or U9400 (N_9400,N_2032,N_4422);
nand U9401 (N_9401,N_3171,N_878);
or U9402 (N_9402,N_766,N_3496);
nor U9403 (N_9403,N_3224,N_2012);
or U9404 (N_9404,N_1951,N_2323);
and U9405 (N_9405,N_4386,N_2482);
nand U9406 (N_9406,N_740,N_1813);
xor U9407 (N_9407,N_3105,N_4411);
xor U9408 (N_9408,N_2510,N_3754);
or U9409 (N_9409,N_2878,N_1682);
nor U9410 (N_9410,N_4045,N_2477);
nand U9411 (N_9411,N_1083,N_2976);
nand U9412 (N_9412,N_4243,N_2422);
and U9413 (N_9413,N_2580,N_3538);
or U9414 (N_9414,N_1651,N_3583);
nand U9415 (N_9415,N_739,N_223);
and U9416 (N_9416,N_711,N_4935);
xor U9417 (N_9417,N_866,N_1509);
or U9418 (N_9418,N_3252,N_3612);
or U9419 (N_9419,N_1426,N_4592);
xnor U9420 (N_9420,N_3035,N_2868);
xor U9421 (N_9421,N_1637,N_2377);
nand U9422 (N_9422,N_620,N_1208);
nor U9423 (N_9423,N_486,N_4252);
and U9424 (N_9424,N_166,N_4347);
or U9425 (N_9425,N_4825,N_1360);
nand U9426 (N_9426,N_1467,N_4931);
xnor U9427 (N_9427,N_3763,N_4290);
nor U9428 (N_9428,N_1195,N_1175);
nand U9429 (N_9429,N_758,N_2856);
xnor U9430 (N_9430,N_2136,N_1886);
xnor U9431 (N_9431,N_149,N_4759);
xor U9432 (N_9432,N_240,N_1993);
and U9433 (N_9433,N_4476,N_1058);
and U9434 (N_9434,N_151,N_347);
nor U9435 (N_9435,N_2903,N_4423);
and U9436 (N_9436,N_2818,N_1218);
or U9437 (N_9437,N_3166,N_3680);
or U9438 (N_9438,N_941,N_3597);
nor U9439 (N_9439,N_2987,N_3352);
nor U9440 (N_9440,N_2320,N_2940);
nand U9441 (N_9441,N_1540,N_4279);
nor U9442 (N_9442,N_357,N_2602);
nand U9443 (N_9443,N_4234,N_4902);
nand U9444 (N_9444,N_3905,N_462);
xnor U9445 (N_9445,N_2638,N_301);
and U9446 (N_9446,N_4789,N_4215);
nor U9447 (N_9447,N_4713,N_77);
nand U9448 (N_9448,N_1146,N_3235);
and U9449 (N_9449,N_4737,N_4244);
nor U9450 (N_9450,N_3939,N_3150);
or U9451 (N_9451,N_279,N_1921);
xnor U9452 (N_9452,N_3828,N_4126);
nand U9453 (N_9453,N_1510,N_616);
nor U9454 (N_9454,N_859,N_648);
or U9455 (N_9455,N_2508,N_1914);
or U9456 (N_9456,N_448,N_410);
nand U9457 (N_9457,N_1125,N_3552);
nand U9458 (N_9458,N_2352,N_4582);
xnor U9459 (N_9459,N_2047,N_419);
or U9460 (N_9460,N_1757,N_4189);
xor U9461 (N_9461,N_2258,N_347);
nor U9462 (N_9462,N_4111,N_3360);
nand U9463 (N_9463,N_4368,N_3064);
nand U9464 (N_9464,N_1081,N_2598);
nor U9465 (N_9465,N_4449,N_3163);
and U9466 (N_9466,N_2991,N_352);
or U9467 (N_9467,N_800,N_3059);
nor U9468 (N_9468,N_3404,N_4683);
xnor U9469 (N_9469,N_2003,N_410);
nor U9470 (N_9470,N_36,N_2233);
or U9471 (N_9471,N_2021,N_3669);
nand U9472 (N_9472,N_4277,N_2769);
and U9473 (N_9473,N_1383,N_4523);
xnor U9474 (N_9474,N_1739,N_2203);
nand U9475 (N_9475,N_3509,N_3101);
nand U9476 (N_9476,N_4527,N_1077);
and U9477 (N_9477,N_1795,N_2528);
and U9478 (N_9478,N_4608,N_4154);
xor U9479 (N_9479,N_450,N_596);
nor U9480 (N_9480,N_2121,N_3878);
nor U9481 (N_9481,N_3669,N_4143);
xor U9482 (N_9482,N_925,N_3890);
or U9483 (N_9483,N_1935,N_3663);
and U9484 (N_9484,N_390,N_1345);
nand U9485 (N_9485,N_3205,N_1776);
nor U9486 (N_9486,N_4798,N_4434);
xnor U9487 (N_9487,N_1252,N_4593);
nand U9488 (N_9488,N_4154,N_1896);
nand U9489 (N_9489,N_682,N_4893);
or U9490 (N_9490,N_3220,N_908);
or U9491 (N_9491,N_21,N_396);
or U9492 (N_9492,N_4347,N_2360);
nor U9493 (N_9493,N_1128,N_144);
or U9494 (N_9494,N_4875,N_902);
and U9495 (N_9495,N_1447,N_4207);
or U9496 (N_9496,N_654,N_2066);
nand U9497 (N_9497,N_4049,N_565);
nor U9498 (N_9498,N_2569,N_2769);
or U9499 (N_9499,N_1080,N_4972);
nand U9500 (N_9500,N_4329,N_1280);
xor U9501 (N_9501,N_1186,N_1397);
and U9502 (N_9502,N_633,N_2363);
and U9503 (N_9503,N_1125,N_3977);
or U9504 (N_9504,N_4078,N_2229);
xnor U9505 (N_9505,N_1880,N_4308);
nor U9506 (N_9506,N_3155,N_2511);
or U9507 (N_9507,N_1305,N_4342);
and U9508 (N_9508,N_1560,N_3106);
nor U9509 (N_9509,N_972,N_935);
nand U9510 (N_9510,N_2375,N_3144);
nand U9511 (N_9511,N_4778,N_1472);
and U9512 (N_9512,N_3344,N_4314);
nand U9513 (N_9513,N_3520,N_2164);
xnor U9514 (N_9514,N_3181,N_1154);
nand U9515 (N_9515,N_4698,N_2698);
and U9516 (N_9516,N_4934,N_2151);
xor U9517 (N_9517,N_2249,N_689);
and U9518 (N_9518,N_4361,N_4028);
or U9519 (N_9519,N_2017,N_1813);
nand U9520 (N_9520,N_1093,N_2117);
and U9521 (N_9521,N_122,N_1600);
nand U9522 (N_9522,N_550,N_2610);
xor U9523 (N_9523,N_4972,N_753);
or U9524 (N_9524,N_1294,N_1363);
xnor U9525 (N_9525,N_768,N_4139);
or U9526 (N_9526,N_1400,N_4064);
nor U9527 (N_9527,N_4113,N_1797);
nand U9528 (N_9528,N_1722,N_4246);
xor U9529 (N_9529,N_645,N_3143);
and U9530 (N_9530,N_1287,N_873);
xnor U9531 (N_9531,N_2546,N_423);
nor U9532 (N_9532,N_145,N_1654);
xor U9533 (N_9533,N_677,N_3920);
or U9534 (N_9534,N_1128,N_2944);
nand U9535 (N_9535,N_2526,N_2635);
xnor U9536 (N_9536,N_118,N_1847);
nor U9537 (N_9537,N_4986,N_296);
or U9538 (N_9538,N_4332,N_477);
xor U9539 (N_9539,N_1990,N_3547);
nor U9540 (N_9540,N_1196,N_4124);
nand U9541 (N_9541,N_4985,N_4276);
xnor U9542 (N_9542,N_1569,N_2142);
xor U9543 (N_9543,N_3736,N_2492);
and U9544 (N_9544,N_4380,N_896);
or U9545 (N_9545,N_2821,N_151);
or U9546 (N_9546,N_429,N_3844);
and U9547 (N_9547,N_1568,N_3783);
or U9548 (N_9548,N_1743,N_3660);
and U9549 (N_9549,N_3246,N_1314);
xor U9550 (N_9550,N_1642,N_1500);
or U9551 (N_9551,N_3947,N_3419);
and U9552 (N_9552,N_4853,N_4805);
and U9553 (N_9553,N_4820,N_1368);
or U9554 (N_9554,N_3156,N_3250);
xor U9555 (N_9555,N_2150,N_817);
xnor U9556 (N_9556,N_1863,N_4866);
nand U9557 (N_9557,N_1704,N_4404);
and U9558 (N_9558,N_950,N_3866);
or U9559 (N_9559,N_536,N_2410);
or U9560 (N_9560,N_2897,N_4827);
or U9561 (N_9561,N_1155,N_2491);
or U9562 (N_9562,N_867,N_1843);
and U9563 (N_9563,N_232,N_2702);
xnor U9564 (N_9564,N_38,N_1756);
nand U9565 (N_9565,N_4672,N_3989);
xor U9566 (N_9566,N_2392,N_4880);
nor U9567 (N_9567,N_4518,N_417);
nor U9568 (N_9568,N_4770,N_1999);
nor U9569 (N_9569,N_3780,N_3586);
or U9570 (N_9570,N_3442,N_706);
nand U9571 (N_9571,N_3279,N_4473);
nand U9572 (N_9572,N_237,N_391);
xor U9573 (N_9573,N_4950,N_1793);
or U9574 (N_9574,N_4358,N_3057);
nand U9575 (N_9575,N_2280,N_3371);
or U9576 (N_9576,N_3286,N_3390);
nand U9577 (N_9577,N_3535,N_3047);
nor U9578 (N_9578,N_3670,N_1756);
or U9579 (N_9579,N_478,N_3272);
and U9580 (N_9580,N_2984,N_4165);
nand U9581 (N_9581,N_4186,N_869);
or U9582 (N_9582,N_578,N_3114);
nand U9583 (N_9583,N_1555,N_1874);
nand U9584 (N_9584,N_184,N_3929);
xor U9585 (N_9585,N_1475,N_4771);
nand U9586 (N_9586,N_1211,N_981);
nor U9587 (N_9587,N_1352,N_2402);
nor U9588 (N_9588,N_330,N_3326);
xor U9589 (N_9589,N_1274,N_287);
nor U9590 (N_9590,N_3961,N_4710);
xnor U9591 (N_9591,N_90,N_1219);
nor U9592 (N_9592,N_929,N_4426);
nand U9593 (N_9593,N_1608,N_4176);
xnor U9594 (N_9594,N_1540,N_2077);
xnor U9595 (N_9595,N_4337,N_513);
or U9596 (N_9596,N_2984,N_4392);
nor U9597 (N_9597,N_2919,N_1121);
nor U9598 (N_9598,N_3859,N_4611);
nand U9599 (N_9599,N_3238,N_3834);
xnor U9600 (N_9600,N_270,N_436);
or U9601 (N_9601,N_3272,N_1311);
xor U9602 (N_9602,N_657,N_3856);
nand U9603 (N_9603,N_4910,N_4897);
or U9604 (N_9604,N_1750,N_1904);
nand U9605 (N_9605,N_4734,N_872);
nor U9606 (N_9606,N_1351,N_70);
or U9607 (N_9607,N_379,N_3271);
xnor U9608 (N_9608,N_1078,N_1343);
nor U9609 (N_9609,N_552,N_85);
or U9610 (N_9610,N_1247,N_409);
or U9611 (N_9611,N_4251,N_1174);
nor U9612 (N_9612,N_4824,N_4490);
nand U9613 (N_9613,N_1897,N_4939);
nand U9614 (N_9614,N_4229,N_1457);
or U9615 (N_9615,N_823,N_4327);
xor U9616 (N_9616,N_1503,N_2494);
nand U9617 (N_9617,N_1450,N_2064);
xnor U9618 (N_9618,N_3727,N_931);
xor U9619 (N_9619,N_4912,N_1708);
and U9620 (N_9620,N_2150,N_4584);
nor U9621 (N_9621,N_2318,N_3740);
and U9622 (N_9622,N_4407,N_937);
nand U9623 (N_9623,N_3674,N_2005);
and U9624 (N_9624,N_3295,N_1335);
nor U9625 (N_9625,N_93,N_601);
nand U9626 (N_9626,N_3964,N_4583);
nor U9627 (N_9627,N_3635,N_3897);
nor U9628 (N_9628,N_2152,N_4382);
and U9629 (N_9629,N_3414,N_1700);
nor U9630 (N_9630,N_2600,N_3409);
and U9631 (N_9631,N_4750,N_2972);
xnor U9632 (N_9632,N_1032,N_1429);
and U9633 (N_9633,N_1559,N_1062);
xor U9634 (N_9634,N_686,N_2714);
nand U9635 (N_9635,N_391,N_797);
and U9636 (N_9636,N_3892,N_3547);
nor U9637 (N_9637,N_3415,N_1344);
or U9638 (N_9638,N_37,N_4211);
or U9639 (N_9639,N_541,N_988);
or U9640 (N_9640,N_1768,N_2404);
nand U9641 (N_9641,N_2954,N_3953);
nand U9642 (N_9642,N_2840,N_3755);
nor U9643 (N_9643,N_3356,N_4303);
or U9644 (N_9644,N_404,N_3200);
nand U9645 (N_9645,N_4754,N_4782);
nand U9646 (N_9646,N_293,N_2235);
xnor U9647 (N_9647,N_2788,N_4388);
or U9648 (N_9648,N_4062,N_2511);
nor U9649 (N_9649,N_1009,N_1727);
xnor U9650 (N_9650,N_1385,N_2402);
xnor U9651 (N_9651,N_1764,N_1466);
and U9652 (N_9652,N_3594,N_695);
xor U9653 (N_9653,N_4231,N_357);
nor U9654 (N_9654,N_4910,N_4250);
and U9655 (N_9655,N_500,N_2461);
or U9656 (N_9656,N_2419,N_2937);
nor U9657 (N_9657,N_4735,N_127);
or U9658 (N_9658,N_1431,N_2080);
nor U9659 (N_9659,N_3468,N_4131);
and U9660 (N_9660,N_27,N_3516);
nor U9661 (N_9661,N_631,N_1968);
nand U9662 (N_9662,N_2181,N_420);
and U9663 (N_9663,N_1716,N_2720);
nand U9664 (N_9664,N_3886,N_1818);
or U9665 (N_9665,N_4804,N_4252);
nand U9666 (N_9666,N_3817,N_733);
or U9667 (N_9667,N_1809,N_4654);
and U9668 (N_9668,N_4222,N_2645);
or U9669 (N_9669,N_2441,N_4036);
nor U9670 (N_9670,N_625,N_2439);
xor U9671 (N_9671,N_2153,N_1343);
or U9672 (N_9672,N_2312,N_2646);
or U9673 (N_9673,N_3617,N_3896);
xnor U9674 (N_9674,N_1765,N_659);
nor U9675 (N_9675,N_3317,N_1416);
nand U9676 (N_9676,N_239,N_4197);
or U9677 (N_9677,N_3069,N_4332);
and U9678 (N_9678,N_1119,N_931);
or U9679 (N_9679,N_4427,N_2714);
xor U9680 (N_9680,N_3393,N_594);
or U9681 (N_9681,N_773,N_3450);
nor U9682 (N_9682,N_833,N_4382);
nand U9683 (N_9683,N_1257,N_4081);
xor U9684 (N_9684,N_547,N_1742);
nand U9685 (N_9685,N_954,N_218);
or U9686 (N_9686,N_370,N_661);
and U9687 (N_9687,N_4459,N_2448);
nand U9688 (N_9688,N_3742,N_2029);
nand U9689 (N_9689,N_1996,N_3647);
nand U9690 (N_9690,N_3897,N_3369);
xor U9691 (N_9691,N_2361,N_223);
or U9692 (N_9692,N_2846,N_4788);
and U9693 (N_9693,N_1383,N_2908);
nand U9694 (N_9694,N_4791,N_636);
xor U9695 (N_9695,N_1081,N_981);
nand U9696 (N_9696,N_858,N_1792);
nor U9697 (N_9697,N_1563,N_1762);
nor U9698 (N_9698,N_3976,N_2879);
nor U9699 (N_9699,N_1166,N_1275);
and U9700 (N_9700,N_4297,N_464);
nand U9701 (N_9701,N_3156,N_1230);
nand U9702 (N_9702,N_1242,N_4776);
nand U9703 (N_9703,N_3200,N_3887);
and U9704 (N_9704,N_3449,N_1418);
and U9705 (N_9705,N_3098,N_730);
xor U9706 (N_9706,N_1460,N_2279);
nand U9707 (N_9707,N_2243,N_224);
and U9708 (N_9708,N_1704,N_1595);
and U9709 (N_9709,N_1781,N_1243);
or U9710 (N_9710,N_1415,N_2378);
and U9711 (N_9711,N_1359,N_144);
nand U9712 (N_9712,N_1123,N_2525);
and U9713 (N_9713,N_994,N_4413);
nor U9714 (N_9714,N_3700,N_1258);
and U9715 (N_9715,N_3250,N_1378);
nand U9716 (N_9716,N_1954,N_4371);
nand U9717 (N_9717,N_636,N_3901);
xor U9718 (N_9718,N_3036,N_425);
and U9719 (N_9719,N_1313,N_4878);
and U9720 (N_9720,N_1233,N_1762);
and U9721 (N_9721,N_33,N_2425);
and U9722 (N_9722,N_4169,N_3233);
nand U9723 (N_9723,N_4612,N_2113);
nand U9724 (N_9724,N_1987,N_2127);
nor U9725 (N_9725,N_905,N_3922);
nand U9726 (N_9726,N_4709,N_103);
nor U9727 (N_9727,N_1602,N_478);
and U9728 (N_9728,N_2340,N_51);
nand U9729 (N_9729,N_162,N_69);
or U9730 (N_9730,N_4425,N_2732);
or U9731 (N_9731,N_1683,N_3177);
or U9732 (N_9732,N_4769,N_2746);
or U9733 (N_9733,N_4635,N_1946);
or U9734 (N_9734,N_2875,N_1654);
and U9735 (N_9735,N_3439,N_3425);
or U9736 (N_9736,N_924,N_2612);
or U9737 (N_9737,N_3991,N_1463);
nor U9738 (N_9738,N_1533,N_4955);
nor U9739 (N_9739,N_1970,N_4670);
and U9740 (N_9740,N_4229,N_1469);
or U9741 (N_9741,N_549,N_3160);
xor U9742 (N_9742,N_1331,N_4875);
nand U9743 (N_9743,N_3374,N_1447);
or U9744 (N_9744,N_628,N_2961);
nor U9745 (N_9745,N_3800,N_189);
xnor U9746 (N_9746,N_2531,N_1062);
and U9747 (N_9747,N_1276,N_4062);
and U9748 (N_9748,N_4986,N_4894);
or U9749 (N_9749,N_627,N_2764);
xor U9750 (N_9750,N_4151,N_3537);
or U9751 (N_9751,N_4540,N_391);
or U9752 (N_9752,N_4271,N_2455);
xnor U9753 (N_9753,N_1204,N_2033);
and U9754 (N_9754,N_175,N_4800);
xnor U9755 (N_9755,N_3867,N_1483);
and U9756 (N_9756,N_3107,N_385);
and U9757 (N_9757,N_4682,N_4194);
or U9758 (N_9758,N_1589,N_1381);
or U9759 (N_9759,N_4757,N_774);
nand U9760 (N_9760,N_2225,N_657);
nor U9761 (N_9761,N_1270,N_485);
nand U9762 (N_9762,N_4559,N_1720);
and U9763 (N_9763,N_996,N_4950);
nor U9764 (N_9764,N_96,N_152);
and U9765 (N_9765,N_1478,N_4412);
xnor U9766 (N_9766,N_3180,N_3265);
nor U9767 (N_9767,N_3558,N_528);
xor U9768 (N_9768,N_960,N_4418);
nor U9769 (N_9769,N_1050,N_2807);
nor U9770 (N_9770,N_3985,N_1769);
or U9771 (N_9771,N_3228,N_2579);
or U9772 (N_9772,N_4398,N_3496);
nand U9773 (N_9773,N_2928,N_2079);
nand U9774 (N_9774,N_4418,N_2470);
nand U9775 (N_9775,N_253,N_887);
or U9776 (N_9776,N_1430,N_1735);
or U9777 (N_9777,N_4510,N_2204);
xor U9778 (N_9778,N_2062,N_4831);
or U9779 (N_9779,N_919,N_1337);
nand U9780 (N_9780,N_4016,N_3044);
nand U9781 (N_9781,N_3735,N_1813);
or U9782 (N_9782,N_4561,N_4023);
xor U9783 (N_9783,N_3565,N_4303);
and U9784 (N_9784,N_3411,N_2183);
or U9785 (N_9785,N_3575,N_524);
nor U9786 (N_9786,N_3246,N_1275);
and U9787 (N_9787,N_4175,N_4679);
nor U9788 (N_9788,N_2344,N_3322);
xor U9789 (N_9789,N_1668,N_3465);
xnor U9790 (N_9790,N_3858,N_859);
nand U9791 (N_9791,N_3548,N_2667);
or U9792 (N_9792,N_2646,N_1509);
xor U9793 (N_9793,N_2393,N_1505);
or U9794 (N_9794,N_2472,N_2901);
and U9795 (N_9795,N_203,N_281);
nor U9796 (N_9796,N_2746,N_2269);
or U9797 (N_9797,N_3190,N_1852);
and U9798 (N_9798,N_433,N_4997);
and U9799 (N_9799,N_2365,N_2230);
xor U9800 (N_9800,N_4356,N_1655);
xor U9801 (N_9801,N_1821,N_3334);
nand U9802 (N_9802,N_542,N_4459);
nor U9803 (N_9803,N_1302,N_998);
nor U9804 (N_9804,N_1527,N_1515);
nor U9805 (N_9805,N_1205,N_316);
and U9806 (N_9806,N_3625,N_4164);
xnor U9807 (N_9807,N_922,N_4262);
and U9808 (N_9808,N_2035,N_1269);
and U9809 (N_9809,N_1035,N_4096);
nand U9810 (N_9810,N_1856,N_825);
and U9811 (N_9811,N_3008,N_1323);
or U9812 (N_9812,N_2712,N_719);
xnor U9813 (N_9813,N_2206,N_4926);
nand U9814 (N_9814,N_4210,N_1643);
or U9815 (N_9815,N_178,N_4476);
or U9816 (N_9816,N_324,N_885);
nor U9817 (N_9817,N_212,N_1808);
nor U9818 (N_9818,N_3454,N_1636);
or U9819 (N_9819,N_430,N_2030);
and U9820 (N_9820,N_3421,N_4713);
nor U9821 (N_9821,N_3911,N_444);
or U9822 (N_9822,N_844,N_2865);
xor U9823 (N_9823,N_3766,N_931);
nor U9824 (N_9824,N_4944,N_446);
or U9825 (N_9825,N_2769,N_1779);
nor U9826 (N_9826,N_1162,N_987);
xnor U9827 (N_9827,N_3533,N_4799);
nor U9828 (N_9828,N_1748,N_579);
or U9829 (N_9829,N_4626,N_4596);
or U9830 (N_9830,N_309,N_4579);
xnor U9831 (N_9831,N_4175,N_2672);
and U9832 (N_9832,N_942,N_534);
or U9833 (N_9833,N_4880,N_4706);
nor U9834 (N_9834,N_2440,N_3964);
nand U9835 (N_9835,N_1951,N_3064);
or U9836 (N_9836,N_3080,N_873);
or U9837 (N_9837,N_2750,N_492);
xor U9838 (N_9838,N_3049,N_1808);
or U9839 (N_9839,N_4240,N_2159);
nand U9840 (N_9840,N_2902,N_1382);
or U9841 (N_9841,N_3465,N_1576);
and U9842 (N_9842,N_2523,N_1372);
nand U9843 (N_9843,N_3984,N_2565);
or U9844 (N_9844,N_765,N_3294);
nor U9845 (N_9845,N_625,N_1150);
or U9846 (N_9846,N_657,N_3626);
nor U9847 (N_9847,N_565,N_3701);
xnor U9848 (N_9848,N_2414,N_2022);
nand U9849 (N_9849,N_4834,N_3913);
xor U9850 (N_9850,N_50,N_4372);
nand U9851 (N_9851,N_4253,N_1700);
xor U9852 (N_9852,N_1156,N_306);
or U9853 (N_9853,N_1610,N_4681);
nand U9854 (N_9854,N_1236,N_1150);
or U9855 (N_9855,N_2908,N_2754);
nand U9856 (N_9856,N_1023,N_2931);
nor U9857 (N_9857,N_146,N_2835);
and U9858 (N_9858,N_2091,N_3153);
or U9859 (N_9859,N_2558,N_577);
xor U9860 (N_9860,N_1583,N_2696);
or U9861 (N_9861,N_2517,N_2371);
xnor U9862 (N_9862,N_514,N_145);
or U9863 (N_9863,N_4134,N_4002);
nor U9864 (N_9864,N_1020,N_4644);
xor U9865 (N_9865,N_429,N_1652);
and U9866 (N_9866,N_2272,N_565);
and U9867 (N_9867,N_3214,N_3477);
nand U9868 (N_9868,N_400,N_4240);
xnor U9869 (N_9869,N_3874,N_4742);
and U9870 (N_9870,N_3806,N_4887);
nor U9871 (N_9871,N_2463,N_3090);
nor U9872 (N_9872,N_1360,N_1121);
xnor U9873 (N_9873,N_1500,N_2989);
and U9874 (N_9874,N_4660,N_2710);
and U9875 (N_9875,N_274,N_1929);
and U9876 (N_9876,N_2534,N_3819);
or U9877 (N_9877,N_1006,N_1113);
and U9878 (N_9878,N_1967,N_2536);
nor U9879 (N_9879,N_3196,N_267);
nand U9880 (N_9880,N_844,N_2035);
nand U9881 (N_9881,N_1476,N_3950);
and U9882 (N_9882,N_4338,N_1490);
nand U9883 (N_9883,N_3317,N_1066);
or U9884 (N_9884,N_4515,N_4848);
xor U9885 (N_9885,N_3698,N_1608);
and U9886 (N_9886,N_4626,N_835);
or U9887 (N_9887,N_1998,N_4404);
and U9888 (N_9888,N_3724,N_2594);
or U9889 (N_9889,N_2159,N_1982);
xnor U9890 (N_9890,N_1078,N_1602);
and U9891 (N_9891,N_3466,N_1372);
or U9892 (N_9892,N_1331,N_2718);
or U9893 (N_9893,N_4929,N_372);
or U9894 (N_9894,N_2784,N_3095);
or U9895 (N_9895,N_3157,N_4594);
xnor U9896 (N_9896,N_2000,N_2820);
nand U9897 (N_9897,N_3000,N_2613);
xor U9898 (N_9898,N_4916,N_2712);
nor U9899 (N_9899,N_1157,N_658);
nand U9900 (N_9900,N_3807,N_3426);
nand U9901 (N_9901,N_3907,N_397);
or U9902 (N_9902,N_2267,N_665);
nor U9903 (N_9903,N_4644,N_3660);
and U9904 (N_9904,N_2341,N_4796);
nor U9905 (N_9905,N_1687,N_4314);
and U9906 (N_9906,N_4655,N_2059);
nor U9907 (N_9907,N_429,N_52);
and U9908 (N_9908,N_4233,N_1056);
or U9909 (N_9909,N_727,N_2825);
nand U9910 (N_9910,N_4684,N_3705);
and U9911 (N_9911,N_374,N_2338);
or U9912 (N_9912,N_2978,N_377);
nor U9913 (N_9913,N_1046,N_2839);
or U9914 (N_9914,N_4907,N_1941);
and U9915 (N_9915,N_2698,N_1589);
and U9916 (N_9916,N_4133,N_945);
and U9917 (N_9917,N_1954,N_1188);
nor U9918 (N_9918,N_2195,N_1786);
or U9919 (N_9919,N_2753,N_1714);
or U9920 (N_9920,N_145,N_3210);
or U9921 (N_9921,N_187,N_565);
and U9922 (N_9922,N_3250,N_2812);
or U9923 (N_9923,N_225,N_2899);
xnor U9924 (N_9924,N_2559,N_754);
and U9925 (N_9925,N_404,N_2561);
xor U9926 (N_9926,N_4973,N_524);
nor U9927 (N_9927,N_2804,N_4802);
nand U9928 (N_9928,N_3381,N_2488);
nand U9929 (N_9929,N_4823,N_3385);
or U9930 (N_9930,N_4348,N_1428);
nand U9931 (N_9931,N_217,N_2267);
and U9932 (N_9932,N_729,N_4205);
or U9933 (N_9933,N_4433,N_1060);
or U9934 (N_9934,N_4940,N_342);
xor U9935 (N_9935,N_4343,N_721);
and U9936 (N_9936,N_1436,N_4627);
nor U9937 (N_9937,N_2397,N_1729);
nor U9938 (N_9938,N_2416,N_1905);
and U9939 (N_9939,N_2205,N_3993);
nand U9940 (N_9940,N_3810,N_1130);
xor U9941 (N_9941,N_4568,N_3761);
xor U9942 (N_9942,N_4974,N_4130);
and U9943 (N_9943,N_4083,N_1487);
or U9944 (N_9944,N_1489,N_1260);
and U9945 (N_9945,N_4588,N_2382);
xor U9946 (N_9946,N_3853,N_2292);
xor U9947 (N_9947,N_4529,N_4284);
xnor U9948 (N_9948,N_4200,N_4913);
and U9949 (N_9949,N_2529,N_3610);
and U9950 (N_9950,N_275,N_1011);
or U9951 (N_9951,N_426,N_3076);
nand U9952 (N_9952,N_169,N_2918);
nand U9953 (N_9953,N_2887,N_4656);
and U9954 (N_9954,N_2901,N_2180);
and U9955 (N_9955,N_3817,N_3756);
nand U9956 (N_9956,N_714,N_937);
and U9957 (N_9957,N_1796,N_1650);
or U9958 (N_9958,N_4181,N_3700);
or U9959 (N_9959,N_2792,N_3325);
nand U9960 (N_9960,N_609,N_1300);
xor U9961 (N_9961,N_2727,N_2257);
or U9962 (N_9962,N_3286,N_46);
or U9963 (N_9963,N_1518,N_1746);
or U9964 (N_9964,N_2044,N_886);
or U9965 (N_9965,N_1213,N_4351);
nand U9966 (N_9966,N_2162,N_3970);
and U9967 (N_9967,N_3212,N_3188);
nor U9968 (N_9968,N_2816,N_4459);
or U9969 (N_9969,N_2509,N_140);
or U9970 (N_9970,N_3432,N_2398);
and U9971 (N_9971,N_3125,N_4293);
nor U9972 (N_9972,N_4569,N_4178);
and U9973 (N_9973,N_3321,N_4003);
or U9974 (N_9974,N_2426,N_2787);
and U9975 (N_9975,N_2049,N_3043);
xnor U9976 (N_9976,N_3905,N_4213);
or U9977 (N_9977,N_1599,N_4921);
nand U9978 (N_9978,N_3046,N_4904);
and U9979 (N_9979,N_4411,N_825);
and U9980 (N_9980,N_165,N_1168);
and U9981 (N_9981,N_24,N_3434);
or U9982 (N_9982,N_1564,N_2869);
and U9983 (N_9983,N_3598,N_4488);
xnor U9984 (N_9984,N_1367,N_1994);
and U9985 (N_9985,N_1552,N_3923);
xor U9986 (N_9986,N_1128,N_2437);
or U9987 (N_9987,N_105,N_807);
nand U9988 (N_9988,N_2902,N_4814);
xnor U9989 (N_9989,N_2310,N_1136);
or U9990 (N_9990,N_150,N_2376);
nand U9991 (N_9991,N_551,N_201);
xnor U9992 (N_9992,N_3420,N_2696);
or U9993 (N_9993,N_4661,N_4711);
and U9994 (N_9994,N_3416,N_4273);
nand U9995 (N_9995,N_476,N_1424);
xor U9996 (N_9996,N_2714,N_2500);
and U9997 (N_9997,N_2803,N_2974);
xor U9998 (N_9998,N_2358,N_3725);
or U9999 (N_9999,N_2145,N_881);
xor U10000 (N_10000,N_6034,N_8171);
nand U10001 (N_10001,N_9580,N_5713);
and U10002 (N_10002,N_6015,N_7108);
and U10003 (N_10003,N_7881,N_9729);
or U10004 (N_10004,N_7262,N_8022);
and U10005 (N_10005,N_5773,N_6858);
nand U10006 (N_10006,N_6025,N_7258);
and U10007 (N_10007,N_6926,N_6701);
nand U10008 (N_10008,N_7979,N_6692);
xnor U10009 (N_10009,N_9868,N_6117);
nand U10010 (N_10010,N_5948,N_6866);
or U10011 (N_10011,N_7410,N_8867);
xnor U10012 (N_10012,N_7550,N_5987);
nor U10013 (N_10013,N_5405,N_5960);
nor U10014 (N_10014,N_8449,N_5208);
xnor U10015 (N_10015,N_5609,N_8840);
and U10016 (N_10016,N_9944,N_8365);
xor U10017 (N_10017,N_7787,N_9299);
and U10018 (N_10018,N_6419,N_6439);
nand U10019 (N_10019,N_6870,N_8961);
nor U10020 (N_10020,N_9077,N_6791);
nor U10021 (N_10021,N_6982,N_7929);
and U10022 (N_10022,N_7765,N_8709);
nand U10023 (N_10023,N_9328,N_8037);
nand U10024 (N_10024,N_5651,N_9276);
and U10025 (N_10025,N_6835,N_6722);
or U10026 (N_10026,N_8686,N_5168);
xor U10027 (N_10027,N_8297,N_9024);
xor U10028 (N_10028,N_8580,N_6972);
or U10029 (N_10029,N_6007,N_5240);
nand U10030 (N_10030,N_7464,N_7894);
nand U10031 (N_10031,N_9466,N_5607);
nand U10032 (N_10032,N_5281,N_9091);
and U10033 (N_10033,N_6712,N_6113);
nand U10034 (N_10034,N_5867,N_9740);
or U10035 (N_10035,N_6407,N_9681);
or U10036 (N_10036,N_7887,N_9732);
or U10037 (N_10037,N_9346,N_8148);
or U10038 (N_10038,N_8200,N_9217);
nor U10039 (N_10039,N_9799,N_9436);
nor U10040 (N_10040,N_6328,N_8450);
xnor U10041 (N_10041,N_7481,N_6843);
nor U10042 (N_10042,N_9356,N_5827);
nor U10043 (N_10043,N_6275,N_5107);
or U10044 (N_10044,N_8787,N_9618);
nand U10045 (N_10045,N_9686,N_7083);
nand U10046 (N_10046,N_9080,N_9408);
nor U10047 (N_10047,N_7255,N_5047);
nand U10048 (N_10048,N_6104,N_7378);
nand U10049 (N_10049,N_5579,N_8878);
nand U10050 (N_10050,N_5089,N_8361);
and U10051 (N_10051,N_9019,N_8298);
and U10052 (N_10052,N_6687,N_5066);
nand U10053 (N_10053,N_8705,N_9338);
or U10054 (N_10054,N_8154,N_9782);
and U10055 (N_10055,N_6698,N_6608);
and U10056 (N_10056,N_9544,N_6251);
and U10057 (N_10057,N_6285,N_5660);
nand U10058 (N_10058,N_9099,N_5812);
nand U10059 (N_10059,N_5043,N_6013);
or U10060 (N_10060,N_8494,N_8672);
and U10061 (N_10061,N_8875,N_9243);
and U10062 (N_10062,N_9362,N_9143);
or U10063 (N_10063,N_9701,N_6740);
nor U10064 (N_10064,N_6081,N_9929);
and U10065 (N_10065,N_8809,N_6356);
nand U10066 (N_10066,N_9988,N_7143);
xnor U10067 (N_10067,N_9115,N_8452);
nor U10068 (N_10068,N_5144,N_7716);
nand U10069 (N_10069,N_5557,N_8668);
nand U10070 (N_10070,N_7019,N_8687);
nor U10071 (N_10071,N_5002,N_7189);
or U10072 (N_10072,N_6404,N_6484);
nor U10073 (N_10073,N_9590,N_5244);
nor U10074 (N_10074,N_7688,N_9357);
and U10075 (N_10075,N_5618,N_8507);
nand U10076 (N_10076,N_6165,N_7321);
xnor U10077 (N_10077,N_5622,N_7977);
xnor U10078 (N_10078,N_9969,N_9600);
nor U10079 (N_10079,N_8525,N_6560);
xor U10080 (N_10080,N_5554,N_5856);
nor U10081 (N_10081,N_5269,N_8420);
nand U10082 (N_10082,N_9985,N_7988);
and U10083 (N_10083,N_8123,N_5217);
nand U10084 (N_10084,N_6916,N_9971);
and U10085 (N_10085,N_9164,N_5008);
and U10086 (N_10086,N_9364,N_9620);
xnor U10087 (N_10087,N_5359,N_7735);
and U10088 (N_10088,N_7400,N_8654);
nor U10089 (N_10089,N_8491,N_5226);
or U10090 (N_10090,N_9124,N_5709);
or U10091 (N_10091,N_7657,N_8575);
nand U10092 (N_10092,N_6848,N_5594);
or U10093 (N_10093,N_7107,N_7561);
nand U10094 (N_10094,N_6445,N_5369);
nand U10095 (N_10095,N_7014,N_8890);
nor U10096 (N_10096,N_7905,N_7487);
nand U10097 (N_10097,N_6547,N_5355);
or U10098 (N_10098,N_9384,N_8874);
nor U10099 (N_10099,N_8052,N_7222);
or U10100 (N_10100,N_5791,N_8489);
xor U10101 (N_10101,N_5422,N_9591);
nor U10102 (N_10102,N_8985,N_6959);
nand U10103 (N_10103,N_8457,N_8090);
nand U10104 (N_10104,N_8158,N_7034);
or U10105 (N_10105,N_9032,N_5239);
or U10106 (N_10106,N_7411,N_7655);
or U10107 (N_10107,N_9864,N_5210);
or U10108 (N_10108,N_7516,N_9222);
xor U10109 (N_10109,N_6453,N_9035);
or U10110 (N_10110,N_8830,N_8376);
or U10111 (N_10111,N_5693,N_8739);
nand U10112 (N_10112,N_8071,N_6323);
nand U10113 (N_10113,N_7354,N_8488);
xor U10114 (N_10114,N_7144,N_5711);
xor U10115 (N_10115,N_9020,N_5521);
nand U10116 (N_10116,N_7599,N_6781);
or U10117 (N_10117,N_6999,N_5677);
and U10118 (N_10118,N_6599,N_7597);
xor U10119 (N_10119,N_8326,N_7250);
nand U10120 (N_10120,N_8124,N_6097);
nand U10121 (N_10121,N_6246,N_9915);
nor U10122 (N_10122,N_7797,N_8898);
nand U10123 (N_10123,N_9284,N_8292);
and U10124 (N_10124,N_9279,N_6896);
xor U10125 (N_10125,N_9201,N_9768);
nor U10126 (N_10126,N_9285,N_5057);
xor U10127 (N_10127,N_8370,N_9050);
xnor U10128 (N_10128,N_9769,N_9885);
xnor U10129 (N_10129,N_8864,N_8577);
or U10130 (N_10130,N_5112,N_7126);
nand U10131 (N_10131,N_6646,N_7745);
nor U10132 (N_10132,N_5808,N_7188);
and U10133 (N_10133,N_8939,N_6772);
xnor U10134 (N_10134,N_8938,N_6925);
or U10135 (N_10135,N_7035,N_5058);
and U10136 (N_10136,N_5337,N_9826);
or U10137 (N_10137,N_5067,N_5558);
and U10138 (N_10138,N_7240,N_8400);
xnor U10139 (N_10139,N_6195,N_5407);
or U10140 (N_10140,N_6253,N_5481);
nor U10141 (N_10141,N_6659,N_6054);
or U10142 (N_10142,N_6934,N_5354);
and U10143 (N_10143,N_7071,N_6052);
or U10144 (N_10144,N_6262,N_6942);
nand U10145 (N_10145,N_8418,N_6640);
nor U10146 (N_10146,N_7123,N_7814);
nand U10147 (N_10147,N_8613,N_5023);
nor U10148 (N_10148,N_7159,N_7016);
nand U10149 (N_10149,N_8551,N_7678);
or U10150 (N_10150,N_9633,N_5434);
or U10151 (N_10151,N_8044,N_8793);
nor U10152 (N_10152,N_6331,N_8646);
nor U10153 (N_10153,N_8925,N_9387);
or U10154 (N_10154,N_6428,N_7635);
or U10155 (N_10155,N_8547,N_6048);
or U10156 (N_10156,N_6639,N_7946);
or U10157 (N_10157,N_8426,N_8333);
or U10158 (N_10158,N_5266,N_6416);
nand U10159 (N_10159,N_7566,N_8283);
nor U10160 (N_10160,N_8579,N_5010);
xor U10161 (N_10161,N_7059,N_8529);
nand U10162 (N_10162,N_5599,N_7552);
xnor U10163 (N_10163,N_6948,N_7295);
nand U10164 (N_10164,N_6927,N_5194);
nor U10165 (N_10165,N_5859,N_5631);
nand U10166 (N_10166,N_5961,N_7010);
nor U10167 (N_10167,N_9809,N_8560);
and U10168 (N_10168,N_8541,N_8702);
nand U10169 (N_10169,N_6035,N_9957);
xnor U10170 (N_10170,N_8942,N_9529);
xor U10171 (N_10171,N_5687,N_8582);
nor U10172 (N_10172,N_5953,N_6402);
or U10173 (N_10173,N_9961,N_7466);
xnor U10174 (N_10174,N_5251,N_9872);
nor U10175 (N_10175,N_9937,N_9053);
xnor U10176 (N_10176,N_7268,N_7095);
nor U10177 (N_10177,N_5092,N_8315);
or U10178 (N_10178,N_8358,N_5674);
and U10179 (N_10179,N_5811,N_7551);
xor U10180 (N_10180,N_5854,N_6456);
xnor U10181 (N_10181,N_7406,N_6799);
nor U10182 (N_10182,N_7547,N_7828);
or U10183 (N_10183,N_9000,N_8909);
nand U10184 (N_10184,N_5012,N_5587);
and U10185 (N_10185,N_7491,N_7362);
nand U10186 (N_10186,N_8980,N_8596);
or U10187 (N_10187,N_7984,N_9555);
nand U10188 (N_10188,N_9948,N_5573);
xor U10189 (N_10189,N_8098,N_5024);
or U10190 (N_10190,N_5486,N_9398);
or U10191 (N_10191,N_5446,N_5629);
nor U10192 (N_10192,N_7831,N_6418);
or U10193 (N_10193,N_8534,N_6759);
or U10194 (N_10194,N_7766,N_9608);
and U10195 (N_10195,N_7184,N_7176);
nand U10196 (N_10196,N_8873,N_6968);
nor U10197 (N_10197,N_9386,N_7585);
nor U10198 (N_10198,N_8199,N_7981);
nand U10199 (N_10199,N_7665,N_5007);
xnor U10200 (N_10200,N_6248,N_8632);
xor U10201 (N_10201,N_8605,N_6429);
nor U10202 (N_10202,N_8462,N_6297);
or U10203 (N_10203,N_8771,N_5155);
nor U10204 (N_10204,N_8643,N_9031);
and U10205 (N_10205,N_6780,N_7571);
nand U10206 (N_10206,N_7293,N_9865);
nor U10207 (N_10207,N_8362,N_9946);
nor U10208 (N_10208,N_5899,N_7274);
nor U10209 (N_10209,N_5431,N_5881);
nand U10210 (N_10210,N_8801,N_7600);
and U10211 (N_10211,N_5996,N_7077);
xor U10212 (N_10212,N_8369,N_7621);
and U10213 (N_10213,N_7965,N_7649);
nor U10214 (N_10214,N_7748,N_7799);
or U10215 (N_10215,N_7524,N_9349);
and U10216 (N_10216,N_7767,N_9882);
and U10217 (N_10217,N_6040,N_7468);
or U10218 (N_10218,N_9756,N_6758);
xor U10219 (N_10219,N_9315,N_7368);
or U10220 (N_10220,N_5983,N_6338);
and U10221 (N_10221,N_8195,N_9564);
xnor U10222 (N_10222,N_9623,N_7111);
nand U10223 (N_10223,N_9294,N_6309);
xor U10224 (N_10224,N_5596,N_7542);
xnor U10225 (N_10225,N_9712,N_6715);
xnor U10226 (N_10226,N_9901,N_8190);
nor U10227 (N_10227,N_9573,N_9136);
nor U10228 (N_10228,N_8975,N_5616);
and U10229 (N_10229,N_9216,N_8557);
xnor U10230 (N_10230,N_8730,N_6793);
or U10231 (N_10231,N_7336,N_5873);
or U10232 (N_10232,N_8626,N_8759);
nor U10233 (N_10233,N_8307,N_9309);
nor U10234 (N_10234,N_5230,N_8395);
nand U10235 (N_10235,N_8153,N_5177);
and U10236 (N_10236,N_8849,N_8314);
xnor U10237 (N_10237,N_5030,N_7838);
xnor U10238 (N_10238,N_7922,N_9463);
or U10239 (N_10239,N_5371,N_9435);
xor U10240 (N_10240,N_6466,N_9639);
xnor U10241 (N_10241,N_6977,N_5744);
and U10242 (N_10242,N_8140,N_8847);
xor U10243 (N_10243,N_5982,N_7795);
or U10244 (N_10244,N_7478,N_7777);
xnor U10245 (N_10245,N_9481,N_7427);
nand U10246 (N_10246,N_9705,N_7584);
xor U10247 (N_10247,N_5655,N_9895);
nor U10248 (N_10248,N_9247,N_5879);
xor U10249 (N_10249,N_8947,N_9416);
nand U10250 (N_10250,N_8761,N_6280);
nand U10251 (N_10251,N_5658,N_5588);
nor U10252 (N_10252,N_9456,N_8366);
xnor U10253 (N_10253,N_9537,N_7985);
nor U10254 (N_10254,N_8956,N_7398);
and U10255 (N_10255,N_5906,N_9366);
nor U10256 (N_10256,N_6124,N_7328);
nand U10257 (N_10257,N_8993,N_9494);
xnor U10258 (N_10258,N_7673,N_8576);
or U10259 (N_10259,N_5895,N_9001);
and U10260 (N_10260,N_7619,N_8998);
xor U10261 (N_10261,N_7507,N_7574);
xor U10262 (N_10262,N_8253,N_6160);
xnor U10263 (N_10263,N_5094,N_6457);
xor U10264 (N_10264,N_6810,N_5746);
or U10265 (N_10265,N_9601,N_5307);
or U10266 (N_10266,N_6293,N_6359);
nand U10267 (N_10267,N_5356,N_9714);
or U10268 (N_10268,N_7200,N_8642);
or U10269 (N_10269,N_5525,N_5743);
nor U10270 (N_10270,N_9310,N_9381);
nor U10271 (N_10271,N_5957,N_9794);
or U10272 (N_10272,N_7241,N_9958);
xor U10273 (N_10273,N_6489,N_8069);
nor U10274 (N_10274,N_5507,N_6600);
xor U10275 (N_10275,N_8727,N_5690);
or U10276 (N_10276,N_8080,N_6783);
nor U10277 (N_10277,N_9818,N_8631);
nand U10278 (N_10278,N_5470,N_6964);
or U10279 (N_10279,N_8715,N_9440);
xor U10280 (N_10280,N_5575,N_8198);
and U10281 (N_10281,N_6764,N_6992);
or U10282 (N_10282,N_5148,N_8012);
xnor U10283 (N_10283,N_7672,N_9272);
and U10284 (N_10284,N_8937,N_6534);
xor U10285 (N_10285,N_5626,N_5528);
nor U10286 (N_10286,N_6296,N_7102);
or U10287 (N_10287,N_7567,N_8664);
nor U10288 (N_10288,N_6522,N_8807);
or U10289 (N_10289,N_7538,N_6244);
nand U10290 (N_10290,N_6973,N_5352);
nor U10291 (N_10291,N_7072,N_8306);
nor U10292 (N_10292,N_7429,N_9760);
nand U10293 (N_10293,N_7634,N_8581);
and U10294 (N_10294,N_9420,N_7667);
nand U10295 (N_10295,N_7757,N_8619);
nor U10296 (N_10296,N_6350,N_5102);
xor U10297 (N_10297,N_6235,N_5125);
nor U10298 (N_10298,N_5967,N_7177);
and U10299 (N_10299,N_6194,N_9635);
xor U10300 (N_10300,N_5219,N_5167);
and U10301 (N_10301,N_6876,N_9018);
nor U10302 (N_10302,N_6766,N_9999);
xnor U10303 (N_10303,N_5615,N_6314);
or U10304 (N_10304,N_6514,N_5817);
nand U10305 (N_10305,N_7025,N_5072);
nand U10306 (N_10306,N_6087,N_8542);
xnor U10307 (N_10307,N_5461,N_6443);
or U10308 (N_10308,N_6967,N_9188);
and U10309 (N_10309,N_5831,N_9910);
or U10310 (N_10310,N_6240,N_5071);
nor U10311 (N_10311,N_8146,N_9779);
xor U10312 (N_10312,N_9371,N_9327);
nor U10313 (N_10313,N_9606,N_5333);
and U10314 (N_10314,N_6474,N_6311);
nand U10315 (N_10315,N_9827,N_9121);
or U10316 (N_10316,N_9215,N_6465);
nor U10317 (N_10317,N_5706,N_7972);
and U10318 (N_10318,N_8299,N_5886);
nand U10319 (N_10319,N_6879,N_5474);
xor U10320 (N_10320,N_8456,N_7685);
xor U10321 (N_10321,N_5719,N_9158);
xor U10322 (N_10322,N_7385,N_7853);
nand U10323 (N_10323,N_9627,N_6621);
nand U10324 (N_10324,N_7002,N_9908);
or U10325 (N_10325,N_8110,N_5601);
and U10326 (N_10326,N_6133,N_8588);
xor U10327 (N_10327,N_9218,N_6539);
and U10328 (N_10328,N_8568,N_8960);
or U10329 (N_10329,N_8217,N_8437);
nand U10330 (N_10330,N_7172,N_8322);
xnor U10331 (N_10331,N_5046,N_6581);
nand U10332 (N_10332,N_5574,N_6614);
nor U10333 (N_10333,N_6819,N_9855);
nand U10334 (N_10334,N_9202,N_8442);
nand U10335 (N_10335,N_9670,N_6778);
or U10336 (N_10336,N_9127,N_7991);
nand U10337 (N_10337,N_5274,N_8764);
nor U10338 (N_10338,N_5098,N_6475);
nand U10339 (N_10339,N_6824,N_9241);
nor U10340 (N_10340,N_9875,N_6568);
and U10341 (N_10341,N_8417,N_7197);
nor U10342 (N_10342,N_5504,N_5918);
nor U10343 (N_10343,N_5025,N_7437);
xor U10344 (N_10344,N_8500,N_9772);
or U10345 (N_10345,N_5611,N_7053);
xor U10346 (N_10346,N_7903,N_9229);
xnor U10347 (N_10347,N_8530,N_8732);
nor U10348 (N_10348,N_9005,N_6066);
and U10349 (N_10349,N_8286,N_8122);
nand U10350 (N_10350,N_5584,N_8966);
or U10351 (N_10351,N_6910,N_5055);
and U10352 (N_10352,N_8453,N_5862);
nor U10353 (N_10353,N_6367,N_6752);
nand U10354 (N_10354,N_9689,N_5756);
nand U10355 (N_10355,N_7650,N_6952);
xnor U10356 (N_10356,N_6271,N_9622);
and U10357 (N_10357,N_6928,N_7289);
and U10358 (N_10358,N_9046,N_8471);
nand U10359 (N_10359,N_9058,N_9187);
and U10360 (N_10360,N_8443,N_7587);
nor U10361 (N_10361,N_7381,N_8341);
and U10362 (N_10362,N_7983,N_7245);
and U10363 (N_10363,N_6526,N_5464);
nand U10364 (N_10364,N_8692,N_9129);
xor U10365 (N_10365,N_8440,N_5749);
nor U10366 (N_10366,N_6143,N_7580);
nor U10367 (N_10367,N_9238,N_5174);
nor U10368 (N_10368,N_6004,N_7801);
or U10369 (N_10369,N_7577,N_8389);
and U10370 (N_10370,N_7224,N_9509);
nor U10371 (N_10371,N_6272,N_7724);
and U10372 (N_10372,N_5797,N_6880);
nor U10373 (N_10373,N_8347,N_5828);
xnor U10374 (N_10374,N_6016,N_9292);
xor U10375 (N_10375,N_6317,N_5530);
and U10376 (N_10376,N_6136,N_8081);
and U10377 (N_10377,N_9097,N_9615);
nand U10378 (N_10378,N_5518,N_7517);
nand U10379 (N_10379,N_7998,N_5400);
nor U10380 (N_10380,N_5546,N_8927);
xnor U10381 (N_10381,N_8302,N_6472);
nand U10382 (N_10382,N_6989,N_7068);
and U10383 (N_10383,N_9715,N_8435);
and U10384 (N_10384,N_8816,N_8811);
and U10385 (N_10385,N_9792,N_8378);
or U10386 (N_10386,N_8691,N_6689);
nor U10387 (N_10387,N_6017,N_5737);
or U10388 (N_10388,N_5727,N_7909);
nand U10389 (N_10389,N_8742,N_9967);
and U10390 (N_10390,N_9313,N_9087);
and U10391 (N_10391,N_7952,N_5496);
nor U10392 (N_10392,N_9459,N_6508);
xor U10393 (N_10393,N_9609,N_5130);
and U10394 (N_10394,N_8061,N_6622);
and U10395 (N_10395,N_5318,N_8774);
or U10396 (N_10396,N_8870,N_8424);
xnor U10397 (N_10397,N_6471,N_7100);
or U10398 (N_10398,N_9566,N_9388);
or U10399 (N_10399,N_5225,N_5198);
nor U10400 (N_10400,N_6111,N_9673);
xnor U10401 (N_10401,N_8892,N_7730);
nand U10402 (N_10402,N_5998,N_9663);
or U10403 (N_10403,N_6763,N_5816);
nand U10404 (N_10404,N_9425,N_6287);
and U10405 (N_10405,N_5196,N_9932);
nand U10406 (N_10406,N_7434,N_7279);
nand U10407 (N_10407,N_8272,N_6050);
nand U10408 (N_10408,N_7915,N_8377);
and U10409 (N_10409,N_6201,N_7682);
nand U10410 (N_10410,N_6965,N_7088);
nor U10411 (N_10411,N_6373,N_6979);
nor U10412 (N_10412,N_8015,N_6458);
and U10413 (N_10413,N_5294,N_9628);
and U10414 (N_10414,N_8229,N_5218);
and U10415 (N_10415,N_6653,N_8587);
or U10416 (N_10416,N_9814,N_9180);
and U10417 (N_10417,N_8103,N_9541);
and U10418 (N_10418,N_5748,N_9744);
nor U10419 (N_10419,N_8428,N_8114);
xor U10420 (N_10420,N_8120,N_7705);
and U10421 (N_10421,N_9848,N_9407);
or U10422 (N_10422,N_6812,N_6361);
and U10423 (N_10423,N_8160,N_9711);
nor U10424 (N_10424,N_7578,N_9232);
or U10425 (N_10425,N_8652,N_8992);
and U10426 (N_10426,N_8591,N_7927);
nor U10427 (N_10427,N_5624,N_5765);
nand U10428 (N_10428,N_6088,N_8329);
nand U10429 (N_10429,N_7135,N_8928);
nor U10430 (N_10430,N_7555,N_6446);
nand U10431 (N_10431,N_9900,N_9036);
or U10432 (N_10432,N_7340,N_9506);
nand U10433 (N_10433,N_7738,N_6396);
nand U10434 (N_10434,N_7302,N_6545);
or U10435 (N_10435,N_6538,N_8725);
xnor U10436 (N_10436,N_8214,N_5848);
nand U10437 (N_10437,N_8111,N_8002);
or U10438 (N_10438,N_7579,N_6389);
or U10439 (N_10439,N_7346,N_9293);
nand U10440 (N_10440,N_6158,N_5424);
nand U10441 (N_10441,N_5454,N_5835);
nand U10442 (N_10442,N_9153,N_5820);
xor U10443 (N_10443,N_9656,N_8622);
nor U10444 (N_10444,N_6288,N_6413);
xnor U10445 (N_10445,N_5166,N_8043);
and U10446 (N_10446,N_7768,N_9479);
nand U10447 (N_10447,N_6938,N_8330);
nor U10448 (N_10448,N_8295,N_7148);
nor U10449 (N_10449,N_5551,N_7811);
or U10450 (N_10450,N_6559,N_9448);
xnor U10451 (N_10451,N_5245,N_9708);
xnor U10452 (N_10452,N_8791,N_7353);
xnor U10453 (N_10453,N_6658,N_9249);
or U10454 (N_10454,N_6383,N_6326);
and U10455 (N_10455,N_9282,N_5206);
nor U10456 (N_10456,N_9360,N_9184);
xnor U10457 (N_10457,N_7690,N_6227);
nand U10458 (N_10458,N_7223,N_5221);
nand U10459 (N_10459,N_5292,N_9921);
and U10460 (N_10460,N_5087,N_8018);
nor U10461 (N_10461,N_6237,N_5988);
or U10462 (N_10462,N_8829,N_6612);
and U10463 (N_10463,N_9086,N_9054);
nand U10464 (N_10464,N_6354,N_6092);
and U10465 (N_10465,N_7775,N_6865);
xor U10466 (N_10466,N_5235,N_6767);
nand U10467 (N_10467,N_7749,N_9075);
nand U10468 (N_10468,N_8549,N_8846);
and U10469 (N_10469,N_8615,N_7926);
nand U10470 (N_10470,N_9197,N_8321);
or U10471 (N_10471,N_7618,N_7511);
or U10472 (N_10472,N_5567,N_9781);
nand U10473 (N_10473,N_6186,N_9662);
and U10474 (N_10474,N_9951,N_6332);
and U10475 (N_10475,N_9010,N_6209);
and U10476 (N_10476,N_7919,N_6028);
nor U10477 (N_10477,N_8678,N_7638);
or U10478 (N_10478,N_7115,N_8554);
nor U10479 (N_10479,N_6177,N_6479);
or U10480 (N_10480,N_6541,N_9329);
nand U10481 (N_10481,N_9755,N_7397);
and U10482 (N_10482,N_5522,N_5493);
and U10483 (N_10483,N_9592,N_6266);
xnor U10484 (N_10484,N_5542,N_5059);
and U10485 (N_10485,N_8499,N_8483);
nor U10486 (N_10486,N_5710,N_5430);
and U10487 (N_10487,N_7616,N_9795);
nor U10488 (N_10488,N_8567,N_7700);
nor U10489 (N_10489,N_9341,N_7254);
and U10490 (N_10490,N_5038,N_7769);
xnor U10491 (N_10491,N_5261,N_7931);
xor U10492 (N_10492,N_9936,N_6208);
nor U10493 (N_10493,N_7548,N_7532);
or U10494 (N_10494,N_6966,N_5312);
xor U10495 (N_10495,N_6482,N_5015);
nand U10496 (N_10496,N_6694,N_8216);
and U10497 (N_10497,N_5362,N_7272);
nand U10498 (N_10498,N_5954,N_5804);
or U10499 (N_10499,N_6613,N_8657);
or U10500 (N_10500,N_5379,N_9568);
nand U10501 (N_10501,N_8915,N_7425);
nand U10502 (N_10502,N_9495,N_9454);
xor U10503 (N_10503,N_8074,N_9178);
xor U10504 (N_10504,N_9862,N_9068);
xnor U10505 (N_10505,N_9009,N_7615);
and U10506 (N_10506,N_7388,N_9752);
xor U10507 (N_10507,N_8179,N_5394);
nor U10508 (N_10508,N_5195,N_7661);
xnor U10509 (N_10509,N_6468,N_5807);
and U10510 (N_10510,N_7997,N_5277);
or U10511 (N_10511,N_7743,N_9759);
nand U10512 (N_10512,N_8282,N_5884);
xnor U10513 (N_10513,N_6995,N_8508);
or U10514 (N_10514,N_9359,N_5149);
xnor U10515 (N_10515,N_9903,N_7049);
nor U10516 (N_10516,N_5268,N_8502);
or U10517 (N_10517,N_8354,N_5770);
nor U10518 (N_10518,N_8930,N_5783);
or U10519 (N_10519,N_5845,N_5722);
nor U10520 (N_10520,N_6957,N_8439);
xnor U10521 (N_10521,N_6286,N_7453);
nand U10522 (N_10522,N_7780,N_5282);
xor U10523 (N_10523,N_9444,N_5774);
nand U10524 (N_10524,N_9913,N_6243);
and U10525 (N_10525,N_5220,N_5000);
nand U10526 (N_10526,N_7277,N_8584);
or U10527 (N_10527,N_7396,N_8480);
or U10528 (N_10528,N_9559,N_8106);
and U10529 (N_10529,N_7598,N_5056);
and U10530 (N_10530,N_5823,N_9645);
xor U10531 (N_10531,N_6076,N_7320);
xnor U10532 (N_10532,N_6461,N_5069);
nor U10533 (N_10533,N_6207,N_6029);
nor U10534 (N_10534,N_7329,N_5045);
nor U10535 (N_10535,N_8446,N_5386);
xnor U10536 (N_10536,N_7231,N_8288);
nand U10537 (N_10537,N_5154,N_8275);
nor U10538 (N_10538,N_9028,N_7956);
or U10539 (N_10539,N_5535,N_8940);
xor U10540 (N_10540,N_7215,N_6574);
and U10541 (N_10541,N_5593,N_5539);
and U10542 (N_10542,N_9939,N_7850);
xor U10543 (N_10543,N_7960,N_5246);
or U10544 (N_10544,N_8023,N_6023);
xor U10545 (N_10545,N_8734,N_5570);
and U10546 (N_10546,N_7654,N_9916);
and U10547 (N_10547,N_7570,N_7726);
nor U10548 (N_10548,N_8385,N_8419);
nand U10549 (N_10549,N_7348,N_9278);
nor U10550 (N_10550,N_9395,N_5039);
nand U10551 (N_10551,N_6563,N_5779);
and U10552 (N_10552,N_5843,N_6065);
nand U10553 (N_10553,N_5922,N_9863);
or U10554 (N_10554,N_8232,N_7029);
nand U10555 (N_10555,N_9918,N_8030);
nor U10556 (N_10556,N_6503,N_8228);
nor U10557 (N_10557,N_7658,N_5286);
xnor U10558 (N_10558,N_5484,N_7916);
or U10559 (N_10559,N_7018,N_9942);
and U10560 (N_10560,N_6036,N_8411);
nor U10561 (N_10561,N_5662,N_5678);
xor U10562 (N_10562,N_8781,N_6424);
and U10563 (N_10563,N_5295,N_5494);
xor U10564 (N_10564,N_5945,N_7414);
or U10565 (N_10565,N_8344,N_7392);
or U10566 (N_10566,N_7859,N_9339);
or U10567 (N_10567,N_6512,N_5329);
and U10568 (N_10568,N_6987,N_9631);
or U10569 (N_10569,N_5133,N_9472);
xnor U10570 (N_10570,N_6231,N_9403);
or U10571 (N_10571,N_7564,N_5760);
xor U10572 (N_10572,N_7201,N_8812);
and U10573 (N_10573,N_8912,N_9478);
or U10574 (N_10574,N_8599,N_7475);
and U10575 (N_10575,N_5947,N_6652);
and U10576 (N_10576,N_8057,N_8072);
nor U10577 (N_10577,N_8540,N_7889);
xnor U10578 (N_10578,N_7356,N_7380);
xor U10579 (N_10579,N_9057,N_9676);
nand U10580 (N_10580,N_9017,N_9935);
xnor U10581 (N_10581,N_5353,N_6583);
nor U10582 (N_10582,N_9482,N_5806);
and U10583 (N_10583,N_9492,N_6099);
nand U10584 (N_10584,N_8648,N_9584);
and U10585 (N_10585,N_8285,N_5520);
nand U10586 (N_10586,N_5639,N_7030);
xnor U10587 (N_10587,N_6825,N_8161);
and U10588 (N_10588,N_5364,N_7306);
nand U10589 (N_10589,N_5316,N_8410);
and U10590 (N_10590,N_6905,N_8150);
xor U10591 (N_10591,N_8403,N_9445);
nand U10592 (N_10592,N_8845,N_8176);
xnor U10593 (N_10593,N_7036,N_9949);
nor U10594 (N_10594,N_8222,N_5620);
and U10595 (N_10595,N_9980,N_6582);
and U10596 (N_10596,N_8373,N_8033);
xnor U10597 (N_10597,N_6665,N_9954);
and U10598 (N_10598,N_8941,N_5630);
and U10599 (N_10599,N_7472,N_7365);
nor U10600 (N_10600,N_8237,N_8486);
and U10601 (N_10601,N_9267,N_6058);
nand U10602 (N_10602,N_8931,N_8796);
nand U10603 (N_10603,N_9757,N_9225);
and U10604 (N_10604,N_8035,N_8303);
nor U10605 (N_10605,N_5439,N_9259);
and U10606 (N_10606,N_5176,N_9607);
and U10607 (N_10607,N_6126,N_5541);
or U10608 (N_10608,N_5483,N_7097);
and U10609 (N_10609,N_5729,N_7951);
and U10610 (N_10610,N_5785,N_9065);
xnor U10611 (N_10611,N_8661,N_8854);
or U10612 (N_10612,N_6702,N_6832);
nand U10613 (N_10613,N_7180,N_7932);
xnor U10614 (N_10614,N_5432,N_9557);
nor U10615 (N_10615,N_6787,N_8905);
xor U10616 (N_10616,N_6026,N_8383);
or U10617 (N_10617,N_8139,N_7914);
nor U10618 (N_10618,N_7504,N_5363);
xnor U10619 (N_10619,N_7146,N_9095);
xor U10620 (N_10620,N_5392,N_7407);
xor U10621 (N_10621,N_5741,N_6277);
and U10622 (N_10622,N_5663,N_9483);
or U10623 (N_10623,N_6333,N_8233);
nor U10624 (N_10624,N_7590,N_6078);
xnor U10625 (N_10625,N_6442,N_6693);
or U10626 (N_10626,N_9098,N_7796);
xor U10627 (N_10627,N_8922,N_5258);
nor U10628 (N_10628,N_8425,N_6704);
nor U10629 (N_10629,N_6595,N_9647);
or U10630 (N_10630,N_5952,N_7457);
or U10631 (N_10631,N_7198,N_7785);
nand U10632 (N_10632,N_9599,N_6869);
nor U10633 (N_10633,N_6696,N_8094);
or U10634 (N_10634,N_6501,N_8105);
and U10635 (N_10635,N_9355,N_6803);
and U10636 (N_10636,N_9470,N_7063);
and U10637 (N_10637,N_8371,N_6360);
xnor U10638 (N_10638,N_7936,N_8733);
xnor U10639 (N_10639,N_9819,N_5236);
or U10640 (N_10640,N_5936,N_6806);
xor U10641 (N_10641,N_7496,N_6757);
and U10642 (N_10642,N_6161,N_6249);
and U10643 (N_10643,N_8461,N_7052);
xnor U10644 (N_10644,N_7244,N_6312);
nor U10645 (N_10645,N_8065,N_5249);
xnor U10646 (N_10646,N_7281,N_6644);
or U10647 (N_10647,N_7298,N_7819);
nor U10648 (N_10648,N_9519,N_8757);
nor U10649 (N_10649,N_7609,N_8536);
nand U10650 (N_10650,N_7686,N_6922);
nand U10651 (N_10651,N_6100,N_6135);
or U10652 (N_10652,N_6346,N_7588);
and U10653 (N_10653,N_9784,N_6018);
or U10654 (N_10654,N_9962,N_9641);
or U10655 (N_10655,N_5141,N_6833);
nor U10656 (N_10656,N_6064,N_9887);
or U10657 (N_10657,N_9905,N_5825);
nor U10658 (N_10658,N_6184,N_8408);
or U10659 (N_10659,N_6523,N_5040);
or U10660 (N_10660,N_7242,N_5457);
nor U10661 (N_10661,N_5247,N_9802);
nor U10662 (N_10662,N_5401,N_6455);
nor U10663 (N_10663,N_8136,N_9177);
nand U10664 (N_10664,N_7737,N_7430);
and U10665 (N_10665,N_8876,N_7046);
xor U10666 (N_10666,N_9090,N_9735);
nor U10667 (N_10667,N_9982,N_8280);
and U10668 (N_10668,N_5723,N_7221);
and U10669 (N_10669,N_9402,N_5140);
and U10670 (N_10670,N_5048,N_6543);
nor U10671 (N_10671,N_6861,N_5035);
nand U10672 (N_10672,N_8144,N_5547);
xor U10673 (N_10673,N_9023,N_7162);
or U10674 (N_10674,N_8995,N_7497);
xor U10675 (N_10675,N_5068,N_9333);
and U10676 (N_10676,N_8503,N_5423);
and U10677 (N_10677,N_8634,N_6552);
and U10678 (N_10678,N_7163,N_7800);
xor U10679 (N_10679,N_7450,N_5681);
nor U10680 (N_10680,N_5169,N_8005);
and U10681 (N_10681,N_5619,N_8647);
nor U10682 (N_10682,N_8563,N_9335);
nor U10683 (N_10683,N_7057,N_7470);
xor U10684 (N_10684,N_9542,N_9101);
or U10685 (N_10685,N_7728,N_7500);
and U10686 (N_10686,N_7236,N_9476);
and U10687 (N_10687,N_8349,N_6857);
nor U10688 (N_10688,N_6902,N_7982);
nor U10689 (N_10689,N_6688,N_6719);
nor U10690 (N_10690,N_7228,N_7349);
and U10691 (N_10691,N_5465,N_7595);
and U10692 (N_10692,N_8031,N_7213);
xor U10693 (N_10693,N_9854,N_7278);
xnor U10694 (N_10694,N_5914,N_9941);
xor U10695 (N_10695,N_7080,N_9849);
nand U10696 (N_10696,N_9014,N_7518);
or U10697 (N_10697,N_6291,N_5684);
nand U10698 (N_10698,N_5365,N_9350);
nor U10699 (N_10699,N_8182,N_8082);
or U10700 (N_10700,N_8552,N_5001);
and U10701 (N_10701,N_8852,N_9651);
or U10702 (N_10702,N_8143,N_7535);
or U10703 (N_10703,N_5145,N_7286);
nand U10704 (N_10704,N_6032,N_5088);
and U10705 (N_10705,N_7129,N_7081);
or U10706 (N_10706,N_7490,N_6854);
and U10707 (N_10707,N_9262,N_8755);
nor U10708 (N_10708,N_5623,N_9893);
nand U10709 (N_10709,N_9596,N_6840);
xor U10710 (N_10710,N_9727,N_6348);
xnor U10711 (N_10711,N_7986,N_8175);
nand U10712 (N_10712,N_6045,N_9323);
or U10713 (N_10713,N_9361,N_6447);
and U10714 (N_10714,N_7545,N_8372);
nand U10715 (N_10715,N_9268,N_8987);
xnor U10716 (N_10716,N_9611,N_9733);
nor U10717 (N_10717,N_5120,N_8404);
and U10718 (N_10718,N_8189,N_9521);
or U10719 (N_10719,N_7352,N_6451);
nand U10720 (N_10720,N_9660,N_8312);
and U10721 (N_10721,N_7543,N_5019);
nand U10722 (N_10722,N_5752,N_8009);
and U10723 (N_10723,N_5849,N_9007);
or U10724 (N_10724,N_6821,N_6478);
or U10725 (N_10725,N_9824,N_6198);
nor U10726 (N_10726,N_9255,N_6737);
and U10727 (N_10727,N_5657,N_9617);
xnor U10728 (N_10728,N_5271,N_9189);
or U10729 (N_10729,N_5935,N_8630);
xor U10730 (N_10730,N_5993,N_8553);
xor U10731 (N_10731,N_6921,N_8024);
nor U10732 (N_10732,N_7601,N_9423);
or U10733 (N_10733,N_6258,N_8463);
xnor U10734 (N_10734,N_6394,N_7238);
or U10735 (N_10735,N_5850,N_7456);
nand U10736 (N_10736,N_6557,N_7602);
or U10737 (N_10737,N_6770,N_7893);
and U10738 (N_10738,N_5234,N_6006);
xor U10739 (N_10739,N_5654,N_6814);
nand U10740 (N_10740,N_5085,N_7314);
or U10741 (N_10741,N_9861,N_5193);
xnor U10742 (N_10742,N_7674,N_8901);
or U10743 (N_10743,N_5991,N_9382);
nand U10744 (N_10744,N_5156,N_9646);
or U10745 (N_10745,N_9286,N_8969);
or U10746 (N_10746,N_6839,N_6216);
and U10747 (N_10747,N_8748,N_7605);
nor U10748 (N_10748,N_6435,N_7386);
or U10749 (N_10749,N_5688,N_6884);
xnor U10750 (N_10750,N_5420,N_7844);
and U10751 (N_10751,N_8826,N_8797);
and U10752 (N_10752,N_6929,N_7546);
nor U10753 (N_10753,N_9437,N_7666);
or U10754 (N_10754,N_9517,N_7541);
and U10755 (N_10755,N_5326,N_7044);
and U10756 (N_10756,N_9228,N_7539);
nand U10757 (N_10757,N_6256,N_8328);
or U10758 (N_10758,N_8535,N_7676);
nor U10759 (N_10759,N_6107,N_6388);
xor U10760 (N_10760,N_6889,N_8208);
and U10761 (N_10761,N_5200,N_8977);
nor U10762 (N_10762,N_8821,N_7441);
xor U10763 (N_10763,N_8550,N_5115);
nor U10764 (N_10764,N_8914,N_9264);
nand U10765 (N_10765,N_6594,N_9801);
nor U10766 (N_10766,N_5384,N_8837);
and U10767 (N_10767,N_6860,N_9842);
nand U10768 (N_10768,N_9242,N_9271);
xnor U10769 (N_10769,N_9828,N_8946);
or U10770 (N_10770,N_5490,N_7645);
and U10771 (N_10771,N_5257,N_5143);
nand U10772 (N_10772,N_9312,N_8244);
nor U10773 (N_10773,N_6790,N_5348);
and U10774 (N_10774,N_8433,N_8751);
or U10775 (N_10775,N_6185,N_5372);
nand U10776 (N_10776,N_5815,N_7058);
or U10777 (N_10777,N_8775,N_8227);
nor U10778 (N_10778,N_8573,N_8291);
and U10779 (N_10779,N_5028,N_7744);
nor U10780 (N_10780,N_6318,N_9467);
and U10781 (N_10781,N_6410,N_6024);
nor U10782 (N_10782,N_7786,N_9100);
or U10783 (N_10783,N_6144,N_9043);
and U10784 (N_10784,N_8628,N_7357);
or U10785 (N_10785,N_7195,N_9535);
nand U10786 (N_10786,N_9850,N_5437);
nor U10787 (N_10787,N_6798,N_9434);
or U10788 (N_10788,N_9514,N_7670);
nor U10789 (N_10789,N_9741,N_9354);
nor U10790 (N_10790,N_9142,N_5419);
nand U10791 (N_10791,N_6263,N_9816);
nand U10792 (N_10792,N_6020,N_8872);
or U10793 (N_10793,N_5358,N_9311);
nand U10794 (N_10794,N_7161,N_7925);
xor U10795 (N_10795,N_9523,N_7704);
xor U10796 (N_10796,N_8178,N_5595);
or U10797 (N_10797,N_7642,N_8406);
and U10798 (N_10798,N_9365,N_9975);
and U10799 (N_10799,N_7008,N_7498);
and U10800 (N_10800,N_6863,N_9083);
nor U10801 (N_10801,N_6173,N_8644);
nor U10802 (N_10802,N_8434,N_5801);
xor U10803 (N_10803,N_7699,N_7824);
and U10804 (N_10804,N_7055,N_9890);
nor U10805 (N_10805,N_6578,N_9516);
xor U10806 (N_10806,N_6168,N_7489);
xnor U10807 (N_10807,N_9273,N_9152);
and U10808 (N_10808,N_6071,N_5931);
nand U10809 (N_10809,N_7446,N_9103);
or U10810 (N_10810,N_9079,N_5304);
xor U10811 (N_10811,N_8802,N_6381);
or U10812 (N_10812,N_5421,N_5398);
nand U10813 (N_10813,N_8239,N_8025);
xnor U10814 (N_10814,N_9579,N_8902);
and U10815 (N_10815,N_7124,N_5635);
nor U10816 (N_10816,N_5842,N_5925);
and U10817 (N_10817,N_7257,N_7752);
or U10818 (N_10818,N_5417,N_6729);
nand U10819 (N_10819,N_9060,N_8028);
and U10820 (N_10820,N_8827,N_5776);
nand U10821 (N_10821,N_8988,N_7890);
or U10822 (N_10822,N_7839,N_6012);
nor U10823 (N_10823,N_8880,N_6362);
xnor U10824 (N_10824,N_7338,N_7283);
nor U10825 (N_10825,N_5833,N_5382);
nor U10826 (N_10826,N_8409,N_6182);
or U10827 (N_10827,N_6935,N_8085);
or U10828 (N_10828,N_7271,N_8497);
or U10829 (N_10829,N_8250,N_8564);
or U10830 (N_10830,N_7312,N_8756);
and U10831 (N_10831,N_6630,N_9843);
and U10832 (N_10832,N_7867,N_8162);
xnor U10833 (N_10833,N_6316,N_5642);
and U10834 (N_10834,N_8210,N_9358);
nand U10835 (N_10835,N_6507,N_8270);
xnor U10836 (N_10836,N_6436,N_5553);
or U10837 (N_10837,N_5137,N_5275);
nand U10838 (N_10838,N_6009,N_8958);
xor U10839 (N_10839,N_5091,N_5844);
nor U10840 (N_10840,N_5839,N_7419);
or U10841 (N_10841,N_8650,N_7643);
nand U10842 (N_10842,N_8255,N_5018);
nor U10843 (N_10843,N_6219,N_9991);
xor U10844 (N_10844,N_8800,N_7880);
and U10845 (N_10845,N_9305,N_9439);
and U10846 (N_10846,N_6425,N_8531);
nor U10847 (N_10847,N_9525,N_7062);
xor U10848 (N_10848,N_9834,N_9724);
xor U10849 (N_10849,N_8659,N_7395);
xnor U10850 (N_10850,N_9140,N_5475);
and U10851 (N_10851,N_9693,N_5426);
and U10852 (N_10852,N_6196,N_7235);
nand U10853 (N_10853,N_6923,N_8570);
and U10854 (N_10854,N_9150,N_9161);
or U10855 (N_10855,N_6105,N_5150);
xor U10856 (N_10856,N_6281,N_7471);
or U10857 (N_10857,N_5278,N_8064);
nand U10858 (N_10858,N_9165,N_7461);
nand U10859 (N_10859,N_6218,N_6751);
nor U10860 (N_10860,N_6463,N_6498);
xor U10861 (N_10861,N_6377,N_7917);
or U10862 (N_10862,N_7740,N_8917);
xnor U10863 (N_10863,N_9055,N_5076);
or U10864 (N_10864,N_8528,N_5758);
or U10865 (N_10865,N_7267,N_9737);
nor U10866 (N_10866,N_7402,N_5604);
nand U10867 (N_10867,N_8595,N_8235);
nor U10868 (N_10868,N_8475,N_8436);
and U10869 (N_10869,N_8444,N_6571);
nor U10870 (N_10870,N_7734,N_8060);
nand U10871 (N_10871,N_7679,N_5049);
xor U10872 (N_10872,N_9166,N_6802);
nand U10873 (N_10873,N_7203,N_5302);
nor U10874 (N_10874,N_6811,N_7680);
xor U10875 (N_10875,N_6898,N_8364);
or U10876 (N_10876,N_7810,N_5301);
xnor U10877 (N_10877,N_7762,N_9373);
or U10878 (N_10878,N_7164,N_5070);
or U10879 (N_10879,N_8224,N_9135);
nor U10880 (N_10880,N_6049,N_7379);
nor U10881 (N_10881,N_6878,N_6075);
or U10882 (N_10882,N_6635,N_7586);
and U10883 (N_10883,N_7361,N_8145);
xor U10884 (N_10884,N_5077,N_7741);
xnor U10885 (N_10885,N_5940,N_5877);
nor U10886 (N_10886,N_8695,N_6939);
nor U10887 (N_10887,N_9089,N_6553);
or U10888 (N_10888,N_5297,N_7739);
nand U10889 (N_10889,N_5129,N_5963);
nor U10890 (N_10890,N_9959,N_8526);
xor U10891 (N_10891,N_6852,N_5583);
or U10892 (N_10892,N_6645,N_7924);
xnor U10893 (N_10893,N_7073,N_6467);
or U10894 (N_10894,N_7297,N_6121);
and U10895 (N_10895,N_8590,N_7276);
xor U10896 (N_10896,N_9841,N_8351);
and U10897 (N_10897,N_9548,N_7121);
nand U10898 (N_10898,N_9806,N_6808);
or U10899 (N_10899,N_9912,N_7280);
or U10900 (N_10900,N_5924,N_6519);
nand U10901 (N_10901,N_6871,N_9515);
or U10902 (N_10902,N_5179,N_5861);
or U10903 (N_10903,N_6486,N_6749);
nor U10904 (N_10904,N_7418,N_9934);
xnor U10905 (N_10905,N_6090,N_7694);
and U10906 (N_10906,N_6887,N_6970);
nand U10907 (N_10907,N_7563,N_5463);
xnor U10908 (N_10908,N_8157,N_5736);
and U10909 (N_10909,N_6163,N_7721);
xor U10910 (N_10910,N_5313,N_7715);
nor U10911 (N_10911,N_5915,N_7310);
nor U10912 (N_10912,N_9839,N_7196);
nand U10913 (N_10913,N_8147,N_8518);
nor U10914 (N_10914,N_7253,N_5874);
and U10915 (N_10915,N_6313,N_9846);
nor U10916 (N_10916,N_9914,N_6535);
xnor U10917 (N_10917,N_9504,N_7776);
xor U10918 (N_10918,N_9671,N_5248);
xnor U10919 (N_10919,N_5733,N_8414);
nor U10920 (N_10920,N_9507,N_7825);
xor U10921 (N_10921,N_5109,N_8639);
and U10922 (N_10922,N_9902,N_9629);
xnor U10923 (N_10923,N_5772,N_5207);
xnor U10924 (N_10924,N_7751,N_6069);
and U10925 (N_10925,N_6001,N_9112);
xnor U10926 (N_10926,N_5223,N_5566);
and U10927 (N_10927,N_5767,N_6518);
nor U10928 (N_10928,N_8238,N_9938);
and U10929 (N_10929,N_8045,N_6485);
xnor U10930 (N_10930,N_8116,N_6667);
or U10931 (N_10931,N_8948,N_5738);
nor U10932 (N_10932,N_9269,N_6671);
nor U10933 (N_10933,N_7261,N_7166);
or U10934 (N_10934,N_7404,N_8290);
and U10935 (N_10935,N_9239,N_5834);
xor U10936 (N_10936,N_6068,N_6505);
nand U10937 (N_10937,N_9248,N_9205);
xnor U10938 (N_10938,N_6877,N_6607);
xor U10939 (N_10939,N_6083,N_5488);
xor U10940 (N_10940,N_7848,N_8511);
xnor U10941 (N_10941,N_7405,N_9696);
nor U10942 (N_10942,N_6953,N_6788);
or U10943 (N_10943,N_6960,N_6936);
xnor U10944 (N_10944,N_6564,N_8056);
nand U10945 (N_10945,N_9840,N_6797);
nor U10946 (N_10946,N_9137,N_8010);
or U10947 (N_10947,N_5044,N_9296);
xor U10948 (N_10948,N_9726,N_5830);
or U10949 (N_10949,N_9405,N_5704);
or U10950 (N_10950,N_9460,N_8000);
xnor U10951 (N_10951,N_6913,N_7079);
nand U10952 (N_10952,N_6221,N_8627);
nor U10953 (N_10953,N_6951,N_7173);
or U10954 (N_10954,N_9983,N_5980);
and U10955 (N_10955,N_7950,N_5503);
xnor U10956 (N_10956,N_6153,N_9774);
nand U10957 (N_10957,N_8910,N_7488);
nor U10958 (N_10958,N_9989,N_7836);
xor U10959 (N_10959,N_5965,N_8916);
and U10960 (N_10960,N_8495,N_5533);
nand U10961 (N_10961,N_9505,N_6422);
nand U10962 (N_10962,N_6947,N_5184);
and U10963 (N_10963,N_6983,N_5777);
nand U10964 (N_10964,N_5121,N_6912);
and U10965 (N_10965,N_5096,N_5443);
xnor U10966 (N_10966,N_5888,N_9786);
nor U10967 (N_10967,N_6755,N_7995);
nand U10968 (N_10968,N_5511,N_6282);
or U10969 (N_10969,N_5290,N_9539);
or U10970 (N_10970,N_5289,N_7636);
xnor U10971 (N_10971,N_9442,N_8096);
and U10972 (N_10972,N_5471,N_8156);
and U10973 (N_10973,N_6606,N_5078);
nand U10974 (N_10974,N_8810,N_6849);
xnor U10975 (N_10975,N_9891,N_9697);
xor U10976 (N_10976,N_5063,N_6801);
or U10977 (N_10977,N_9261,N_9758);
or U10978 (N_10978,N_7559,N_7957);
nor U10979 (N_10979,N_9652,N_5682);
xnor U10980 (N_10980,N_6592,N_9672);
or U10981 (N_10981,N_6171,N_7829);
or U10982 (N_10982,N_8331,N_5472);
nor U10983 (N_10983,N_6002,N_7150);
nor U10984 (N_10984,N_9195,N_6883);
nand U10985 (N_10985,N_7269,N_7589);
and U10986 (N_10986,N_6395,N_9037);
nor U10987 (N_10987,N_5079,N_7736);
xor U10988 (N_10988,N_6845,N_7117);
xor U10989 (N_10989,N_7692,N_9621);
nor U10990 (N_10990,N_7576,N_7971);
xnor U10991 (N_10991,N_9556,N_7761);
and U10992 (N_10992,N_7192,N_5523);
or U10993 (N_10993,N_5725,N_9093);
or U10994 (N_10994,N_9322,N_6956);
and U10995 (N_10995,N_6299,N_9379);
nand U10996 (N_10996,N_7613,N_8844);
xnor U10997 (N_10997,N_9522,N_5939);
xor U10998 (N_10998,N_9823,N_5502);
nor U10999 (N_10999,N_7534,N_5605);
or U11000 (N_11000,N_8886,N_8267);
nor U11001 (N_11001,N_5676,N_7876);
or U11002 (N_11002,N_6164,N_9219);
nand U11003 (N_11003,N_8076,N_7773);
or U11004 (N_11004,N_8174,N_8684);
nand U11005 (N_11005,N_6134,N_9027);
nand U11006 (N_11006,N_9833,N_9457);
xor U11007 (N_11007,N_5985,N_8688);
nor U11008 (N_11008,N_5667,N_7194);
nor U11009 (N_11009,N_5373,N_9290);
nand U11010 (N_11010,N_5602,N_6349);
or U11011 (N_11011,N_9220,N_6340);
and U11012 (N_11012,N_8135,N_7103);
or U11013 (N_11013,N_5122,N_8308);
and U11014 (N_11014,N_6566,N_7802);
and U11015 (N_11015,N_9307,N_5135);
or U11016 (N_11016,N_7845,N_9040);
nor U11017 (N_11017,N_9061,N_7084);
nand U11018 (N_11018,N_7695,N_9750);
or U11019 (N_11019,N_9528,N_6357);
nor U11020 (N_11020,N_7644,N_8566);
nor U11021 (N_11021,N_7315,N_6513);
or U11022 (N_11022,N_6238,N_8608);
or U11023 (N_11023,N_7784,N_8167);
or U11024 (N_11024,N_7843,N_9453);
nor U11025 (N_11025,N_9734,N_9297);
nand U11026 (N_11026,N_7399,N_5668);
nand U11027 (N_11027,N_8164,N_6335);
or U11028 (N_11028,N_6411,N_8336);
nor U11029 (N_11029,N_9904,N_5592);
and U11030 (N_11030,N_9510,N_8700);
nor U11031 (N_11031,N_6154,N_7401);
and U11032 (N_11032,N_7554,N_8460);
nor U11033 (N_11033,N_5907,N_7611);
or U11034 (N_11034,N_5042,N_9553);
nand U11035 (N_11035,N_6546,N_6874);
xor U11036 (N_11036,N_7809,N_9762);
or U11037 (N_11037,N_5645,N_8048);
nand U11038 (N_11038,N_8629,N_6649);
nand U11039 (N_11039,N_9943,N_6632);
nand U11040 (N_11040,N_7375,N_7993);
or U11041 (N_11041,N_5097,N_9979);
xor U11042 (N_11042,N_8125,N_9907);
or U11043 (N_11043,N_8477,N_7753);
nand U11044 (N_11044,N_9598,N_7701);
or U11045 (N_11045,N_6174,N_6823);
and U11046 (N_11046,N_7334,N_8268);
xnor U11047 (N_11047,N_9275,N_9619);
and U11048 (N_11048,N_6731,N_7116);
and U11049 (N_11049,N_8660,N_5860);
xnor U11050 (N_11050,N_6604,N_6086);
or U11051 (N_11051,N_5582,N_6986);
xor U11052 (N_11052,N_8482,N_7610);
xnor U11053 (N_11053,N_8773,N_7011);
or U11054 (N_11054,N_7964,N_6572);
nand U11055 (N_11055,N_9753,N_8316);
nand U11056 (N_11056,N_6703,N_6298);
xnor U11057 (N_11057,N_6903,N_8851);
or U11058 (N_11058,N_6888,N_7384);
xor U11059 (N_11059,N_8206,N_8472);
and U11060 (N_11060,N_5739,N_5116);
nor U11061 (N_11061,N_5183,N_7335);
nand U11062 (N_11062,N_6765,N_7422);
nand U11063 (N_11063,N_5666,N_6690);
and U11064 (N_11064,N_6483,N_5074);
and U11065 (N_11065,N_5053,N_8959);
nor U11066 (N_11066,N_9867,N_9817);
and U11067 (N_11067,N_9940,N_6039);
nor U11068 (N_11068,N_5142,N_6351);
nor U11069 (N_11069,N_6616,N_6680);
or U11070 (N_11070,N_7681,N_9344);
xor U11071 (N_11071,N_6233,N_6996);
nor U11072 (N_11072,N_6415,N_9692);
nor U11073 (N_11073,N_6551,N_6532);
nand U11074 (N_11074,N_9223,N_7920);
xor U11075 (N_11075,N_5203,N_9586);
and U11076 (N_11076,N_6720,N_8219);
and U11077 (N_11077,N_6700,N_9116);
nor U11078 (N_11078,N_6855,N_7033);
and U11079 (N_11079,N_9721,N_6591);
xnor U11080 (N_11080,N_9450,N_5182);
and U11081 (N_11081,N_8651,N_8487);
and U11082 (N_11082,N_5438,N_9512);
nor U11083 (N_11083,N_9390,N_7424);
or U11084 (N_11084,N_7945,N_9154);
xor U11085 (N_11085,N_6742,N_5872);
or U11086 (N_11086,N_8817,N_7251);
and U11087 (N_11087,N_5101,N_6358);
nand U11088 (N_11088,N_7067,N_9899);
or U11089 (N_11089,N_9430,N_9657);
nor U11090 (N_11090,N_9070,N_8427);
xor U11091 (N_11091,N_5410,N_8032);
nor U11092 (N_11092,N_6754,N_8274);
or U11093 (N_11093,N_6284,N_6080);
or U11094 (N_11094,N_7624,N_7710);
nor U11095 (N_11095,N_8900,N_6382);
nand U11096 (N_11096,N_9612,N_9871);
nor U11097 (N_11097,N_6499,N_5026);
xnor U11098 (N_11098,N_5591,N_8957);
nor U11099 (N_11099,N_7026,N_8026);
xor U11100 (N_11100,N_5878,N_7746);
and U11101 (N_11101,N_5250,N_9073);
xor U11102 (N_11102,N_6386,N_6473);
and U11103 (N_11103,N_7005,N_7003);
xnor U11104 (N_11104,N_6500,N_5720);
and U11105 (N_11105,N_5299,N_9224);
xnor U11106 (N_11106,N_9319,N_5803);
and U11107 (N_11107,N_9022,N_6245);
nand U11108 (N_11108,N_8848,N_9141);
xor U11109 (N_11109,N_8118,N_7864);
nand U11110 (N_11110,N_5351,N_7856);
nor U11111 (N_11111,N_8151,N_9383);
nor U11112 (N_11112,N_5428,N_5855);
or U11113 (N_11113,N_6030,N_6744);
nand U11114 (N_11114,N_5919,N_5865);
xor U11115 (N_11115,N_5625,N_6641);
or U11116 (N_11116,N_8075,N_5315);
xnor U11117 (N_11117,N_9417,N_8945);
and U11118 (N_11118,N_9775,N_6063);
xnor U11119 (N_11119,N_8888,N_5036);
or U11120 (N_11120,N_7623,N_9709);
nand U11121 (N_11121,N_9374,N_5255);
or U11122 (N_11122,N_5891,N_7112);
and U11123 (N_11123,N_8823,N_6320);
xor U11124 (N_11124,N_9301,N_6847);
and U11125 (N_11125,N_9798,N_5726);
nand U11126 (N_11126,N_5202,N_6730);
or U11127 (N_11127,N_8783,N_7606);
nor U11128 (N_11128,N_8399,N_8230);
nand U11129 (N_11129,N_6250,N_5686);
or U11130 (N_11130,N_5598,N_7522);
xor U11131 (N_11131,N_8375,N_6232);
nor U11132 (N_11132,N_9678,N_5340);
and U11133 (N_11133,N_8429,N_7821);
nand U11134 (N_11134,N_7813,N_8729);
xnor U11135 (N_11135,N_9283,N_8640);
nand U11136 (N_11136,N_6661,N_5968);
or U11137 (N_11137,N_6370,N_7641);
and U11138 (N_11138,N_9597,N_8412);
nand U11139 (N_11139,N_6390,N_7006);
or U11140 (N_11140,N_7139,N_9162);
and U11141 (N_11141,N_7506,N_5322);
nor U11142 (N_11142,N_5597,N_8520);
xor U11143 (N_11143,N_6991,N_7847);
and U11144 (N_11144,N_9730,N_7485);
xor U11145 (N_11145,N_8093,N_7754);
nand U11146 (N_11146,N_9280,N_7499);
xor U11147 (N_11147,N_8868,N_5532);
nand U11148 (N_11148,N_7549,N_6775);
and U11149 (N_11149,N_6189,N_7358);
or U11150 (N_11150,N_9084,N_5173);
and U11151 (N_11151,N_7296,N_5228);
and U11152 (N_11152,N_9465,N_8728);
xor U11153 (N_11153,N_5452,N_9706);
xnor U11154 (N_11154,N_9587,N_8726);
and U11155 (N_11155,N_7830,N_6837);
nor U11156 (N_11156,N_9830,N_8269);
nand U11157 (N_11157,N_6962,N_7907);
and U11158 (N_11158,N_5476,N_7553);
or U11159 (N_11159,N_7963,N_9847);
nand U11160 (N_11160,N_7061,N_8263);
nor U11161 (N_11161,N_7042,N_7041);
or U11162 (N_11162,N_8084,N_7999);
xnor U11163 (N_11163,N_7219,N_7628);
nor U11164 (N_11164,N_6116,N_9447);
xor U11165 (N_11165,N_6057,N_7514);
or U11166 (N_11166,N_5325,N_5989);
and U11167 (N_11167,N_6981,N_5871);
nand U11168 (N_11168,N_5259,N_8266);
xnor U11169 (N_11169,N_7849,N_7342);
nor U11170 (N_11170,N_5160,N_9530);
xor U11171 (N_11171,N_7436,N_5568);
and U11172 (N_11172,N_6110,N_7855);
and U11173 (N_11173,N_7509,N_8402);
xor U11174 (N_11174,N_7558,N_5664);
or U11175 (N_11175,N_6450,N_9526);
nand U11176 (N_11176,N_5022,N_7698);
or U11177 (N_11177,N_8698,N_8658);
and U11178 (N_11178,N_9745,N_5050);
or U11179 (N_11179,N_9569,N_5904);
and U11180 (N_11180,N_7371,N_9108);
nor U11181 (N_11181,N_5508,N_7770);
nor U11182 (N_11182,N_7232,N_5451);
and U11183 (N_11183,N_7660,N_7966);
or U11184 (N_11184,N_8046,N_5890);
xnor U11185 (N_11185,N_6343,N_6807);
and U11186 (N_11186,N_8506,N_7817);
xor U11187 (N_11187,N_8934,N_5131);
xnor U11188 (N_11188,N_5798,N_6709);
xnor U11189 (N_11189,N_9118,N_6059);
and U11190 (N_11190,N_9953,N_5636);
xor U11191 (N_11191,N_9791,N_9451);
nand U11192 (N_11192,N_6283,N_7732);
nand U11193 (N_11193,N_8313,N_7130);
and U11194 (N_11194,N_6524,N_5699);
and U11195 (N_11195,N_8895,N_6336);
xnor U11196 (N_11196,N_5778,N_9498);
nand U11197 (N_11197,N_9175,N_6344);
or U11198 (N_11198,N_9490,N_9392);
nor U11199 (N_11199,N_5928,N_9110);
nand U11200 (N_11200,N_5480,N_5921);
and U11201 (N_11201,N_5659,N_7841);
nand U11202 (N_11202,N_5273,N_9630);
nor U11203 (N_11203,N_8236,N_6454);
or U11204 (N_11204,N_9074,N_9920);
nor U11205 (N_11205,N_5242,N_7167);
nand U11206 (N_11206,N_8884,N_6214);
and U11207 (N_11207,N_6602,N_8234);
nor U11208 (N_11208,N_9289,N_7512);
or U11209 (N_11209,N_5128,N_5732);
or U11210 (N_11210,N_7996,N_8614);
nand U11211 (N_11211,N_6834,N_9156);
xnor U11212 (N_11212,N_8908,N_6303);
nand U11213 (N_11213,N_7793,N_5238);
or U11214 (N_11214,N_5455,N_9837);
nand U11215 (N_11215,N_8991,N_9739);
or U11216 (N_11216,N_9011,N_7479);
and U11217 (N_11217,N_9171,N_6139);
nor U11218 (N_11218,N_6226,N_9015);
or U11219 (N_11219,N_8638,N_8343);
or U11220 (N_11220,N_7959,N_5755);
nand U11221 (N_11221,N_9480,N_8871);
xor U11222 (N_11222,N_5606,N_8398);
nand U11223 (N_11223,N_7170,N_7403);
and U11224 (N_11224,N_8401,N_9897);
and U11225 (N_11225,N_8616,N_6399);
or U11226 (N_11226,N_9497,N_9675);
and U11227 (N_11227,N_7878,N_7182);
nand U11228 (N_11228,N_5321,N_7789);
nand U11229 (N_11229,N_9092,N_6706);
or U11230 (N_11230,N_7529,N_7137);
nand U11231 (N_11231,N_6259,N_5802);
nand U11232 (N_11232,N_9345,N_5014);
nor U11233 (N_11233,N_5912,N_6188);
or U11234 (N_11234,N_5449,N_9085);
nand U11235 (N_11235,N_6710,N_6091);
xor U11236 (N_11236,N_8353,N_9493);
nor U11237 (N_11237,N_5973,N_7782);
nand U11238 (N_11238,N_6496,N_6192);
xor U11239 (N_11239,N_7930,N_8183);
and U11240 (N_11240,N_6528,N_5296);
xor U11241 (N_11241,N_7962,N_9500);
nand U11242 (N_11242,N_5903,N_5393);
or U11243 (N_11243,N_7693,N_7382);
nand U11244 (N_11244,N_7941,N_9518);
xnor U11245 (N_11245,N_7285,N_8565);
nor U11246 (N_11246,N_6374,N_9638);
nand U11247 (N_11247,N_5634,N_8392);
or U11248 (N_11248,N_8166,N_5841);
nand U11249 (N_11249,N_5190,N_7593);
nor U11250 (N_11250,N_6181,N_8186);
nor U11251 (N_11251,N_6257,N_9815);
xor U11252 (N_11252,N_7039,N_5864);
nand U11253 (N_11253,N_7647,N_5108);
nor U11254 (N_11254,N_6598,N_9399);
nand U11255 (N_11255,N_6904,N_6421);
nor U11256 (N_11256,N_9879,N_8714);
xnor U11257 (N_11257,N_6850,N_8974);
nand U11258 (N_11258,N_5347,N_7208);
nand U11259 (N_11259,N_8346,N_8633);
and U11260 (N_11260,N_9973,N_8662);
nand U11261 (N_11261,N_8745,N_6391);
and U11262 (N_11262,N_6554,N_6084);
nand U11263 (N_11263,N_8097,N_7263);
nand U11264 (N_11264,N_8690,N_7884);
nand U11265 (N_11265,N_5162,N_5665);
xnor U11266 (N_11266,N_5396,N_8305);
xnor U11267 (N_11267,N_7778,N_9805);
xnor U11268 (N_11268,N_9877,N_9081);
xnor U11269 (N_11269,N_5950,N_6140);
nand U11270 (N_11270,N_7439,N_8036);
or U11271 (N_11271,N_9534,N_7872);
and U11272 (N_11272,N_8350,N_9302);
nand U11273 (N_11273,N_7703,N_8131);
nand U11274 (N_11274,N_9683,N_5436);
nor U11275 (N_11275,N_8666,N_7408);
nor U11276 (N_11276,N_9771,N_7747);
or U11277 (N_11277,N_6853,N_5641);
xor U11278 (N_11278,N_9400,N_5889);
and U11279 (N_11279,N_6321,N_7217);
nand U11280 (N_11280,N_8782,N_5211);
or U11281 (N_11281,N_5824,N_8091);
or U11282 (N_11282,N_5846,N_9972);
nor U11283 (N_11283,N_6617,N_9570);
nor U11284 (N_11284,N_8724,N_6495);
and U11285 (N_11285,N_7347,N_8770);
nor U11286 (N_11286,N_7933,N_5707);
nand U11287 (N_11287,N_7742,N_8780);
nand U11288 (N_11288,N_9667,N_7815);
nand U11289 (N_11289,N_8964,N_6516);
nand U11290 (N_11290,N_8719,N_6376);
or U11291 (N_11291,N_7662,N_6521);
or U11292 (N_11292,N_5516,N_6971);
or U11293 (N_11293,N_6707,N_9351);
nor U11294 (N_11294,N_9252,N_6044);
and U11295 (N_11295,N_6176,N_5308);
or U11296 (N_11296,N_6112,N_5851);
and U11297 (N_11297,N_9807,N_8262);
or U11298 (N_11298,N_8562,N_9369);
or U11299 (N_11299,N_6998,N_6264);
xor U11300 (N_11300,N_9183,N_9870);
xnor U11301 (N_11301,N_5216,N_8155);
and U11302 (N_11302,N_6576,N_7323);
nand U11303 (N_11303,N_9742,N_6037);
or U11304 (N_11304,N_8514,N_9533);
and U11305 (N_11305,N_5763,N_7082);
and U11306 (N_11306,N_9574,N_6931);
xor U11307 (N_11307,N_8623,N_9687);
nor U11308 (N_11308,N_9473,N_6527);
nand U11309 (N_11309,N_5395,N_7113);
and U11310 (N_11310,N_5505,N_5309);
or U11311 (N_11311,N_5781,N_9661);
nor U11312 (N_11312,N_7031,N_9613);
xnor U11313 (N_11313,N_5435,N_8997);
nand U11314 (N_11314,N_7804,N_7975);
and U11315 (N_11315,N_9616,N_7389);
xor U11316 (N_11316,N_6738,N_7772);
xor U11317 (N_11317,N_6220,N_6363);
nor U11318 (N_11318,N_8247,N_9977);
and U11319 (N_11319,N_8641,N_5852);
xor U11320 (N_11320,N_9226,N_9669);
nand U11321 (N_11321,N_9172,N_6041);
nor U11322 (N_11322,N_5442,N_6533);
xnor U11323 (N_11323,N_9603,N_5153);
xor U11324 (N_11324,N_9761,N_7027);
xnor U11325 (N_11325,N_5264,N_6403);
nand U11326 (N_11326,N_6241,N_5932);
nand U11327 (N_11327,N_9052,N_8704);
or U11328 (N_11328,N_5252,N_8356);
nor U11329 (N_11329,N_9945,N_5689);
xnor U11330 (N_11330,N_5787,N_8762);
and U11331 (N_11331,N_6993,N_8132);
xnor U11332 (N_11332,N_6342,N_9308);
xnor U11333 (N_11333,N_7544,N_7540);
xnor U11334 (N_11334,N_9094,N_6555);
or U11335 (N_11335,N_5111,N_8655);
or U11336 (N_11336,N_8944,N_6627);
or U11337 (N_11337,N_9707,N_5715);
nor U11338 (N_11338,N_9353,N_8310);
or U11339 (N_11339,N_9560,N_9788);
nor U11340 (N_11340,N_9894,N_7992);
nor U11341 (N_11341,N_7794,N_8881);
nand U11342 (N_11342,N_5562,N_5585);
nor U11343 (N_11343,N_9277,N_6836);
nor U11344 (N_11344,N_7990,N_5771);
or U11345 (N_11345,N_9109,N_7259);
and U11346 (N_11346,N_8379,N_7935);
nor U11347 (N_11347,N_6897,N_9776);
and U11348 (N_11348,N_9291,N_6205);
or U11349 (N_11349,N_9130,N_9777);
xor U11350 (N_11350,N_9898,N_8459);
and U11351 (N_11351,N_9469,N_9477);
nor U11352 (N_11352,N_8223,N_9221);
nor U11353 (N_11353,N_7953,N_8338);
nor U11354 (N_11354,N_5338,N_8653);
and U11355 (N_11355,N_9428,N_6372);
xor U11356 (N_11356,N_5569,N_6255);
nand U11357 (N_11357,N_9213,N_5724);
or U11358 (N_11358,N_6155,N_5813);
or U11359 (N_11359,N_7949,N_7874);
nor U11360 (N_11360,N_7442,N_5847);
xnor U11361 (N_11361,N_8904,N_8561);
nand U11362 (N_11362,N_6380,N_7423);
and U11363 (N_11363,N_6115,N_5956);
or U11364 (N_11364,N_9532,N_7022);
nand U11365 (N_11365,N_6809,N_8697);
nor U11366 (N_11366,N_6469,N_5425);
xor U11367 (N_11367,N_7750,N_9665);
xnor U11368 (N_11368,N_6067,N_6191);
xor U11369 (N_11369,N_5714,N_5712);
nor U11370 (N_11370,N_5730,N_6517);
xnor U11371 (N_11371,N_8521,N_9571);
xnor U11372 (N_11372,N_8332,N_9409);
xor U11373 (N_11373,N_9394,N_8731);
xor U11374 (N_11374,N_7938,N_7980);
nand U11375 (N_11375,N_9589,N_5479);
nor U11376 (N_11376,N_8976,N_6123);
nand U11377 (N_11377,N_6047,N_5747);
and U11378 (N_11378,N_5440,N_7131);
xor U11379 (N_11379,N_7648,N_5564);
or U11380 (N_11380,N_7592,N_8753);
xor U11381 (N_11381,N_6727,N_7273);
nor U11382 (N_11382,N_9527,N_9748);
nor U11383 (N_11383,N_7906,N_8926);
nand U11384 (N_11384,N_8447,N_7206);
nand U11385 (N_11385,N_5126,N_9499);
nand U11386 (N_11386,N_7474,N_8965);
nand U11387 (N_11387,N_8468,N_8095);
or U11388 (N_11388,N_6625,N_9725);
xor U11389 (N_11389,N_8548,N_5971);
nor U11390 (N_11390,N_5124,N_5810);
or U11391 (N_11391,N_5669,N_8879);
nor U11392 (N_11392,N_5083,N_5986);
nor U11393 (N_11393,N_5383,N_7074);
xor U11394 (N_11394,N_8006,N_6974);
or U11395 (N_11395,N_6678,N_8451);
xnor U11396 (N_11396,N_8598,N_7243);
nor U11397 (N_11397,N_9790,N_8099);
nand U11398 (N_11398,N_6322,N_7515);
nand U11399 (N_11399,N_8187,N_5671);
or U11400 (N_11400,N_9078,N_5628);
xnor U11401 (N_11401,N_5955,N_7835);
nand U11402 (N_11402,N_6750,N_6405);
xnor U11403 (N_11403,N_7136,N_9933);
nor U11404 (N_11404,N_5224,N_5159);
and U11405 (N_11405,N_8126,N_5334);
or U11406 (N_11406,N_6743,N_6393);
and U11407 (N_11407,N_8718,N_5118);
nor U11408 (N_11408,N_6202,N_7013);
xnor U11409 (N_11409,N_5291,N_5692);
and U11410 (N_11410,N_7360,N_7367);
or U11411 (N_11411,N_9324,N_8201);
xor U11412 (N_11412,N_8079,N_9738);
nor U11413 (N_11413,N_7341,N_7708);
nor U11414 (N_11414,N_7834,N_7369);
nor U11415 (N_11415,N_5685,N_5032);
nand U11416 (N_11416,N_7758,N_6179);
and U11417 (N_11417,N_8933,N_7114);
or U11418 (N_11418,N_5306,N_8117);
nand U11419 (N_11419,N_9064,N_9102);
and U11420 (N_11420,N_7098,N_8706);
nor U11421 (N_11421,N_9265,N_7707);
nand U11422 (N_11422,N_5172,N_7857);
or U11423 (N_11423,N_6650,N_8519);
and U11424 (N_11424,N_8574,N_7781);
and U11425 (N_11425,N_5344,N_6119);
nor U11426 (N_11426,N_5805,N_8612);
nor U11427 (N_11427,N_5653,N_5984);
nor U11428 (N_11428,N_7152,N_7961);
or U11429 (N_11429,N_6724,N_9659);
nand U11430 (N_11430,N_5081,N_9254);
nor U11431 (N_11431,N_5123,N_8304);
and U11432 (N_11432,N_7885,N_5673);
nor U11433 (N_11433,N_7771,N_9567);
xor U11434 (N_11434,N_6924,N_5799);
and U11435 (N_11435,N_9071,N_6891);
and U11436 (N_11436,N_8464,N_5113);
nor U11437 (N_11437,N_5556,N_6549);
nand U11438 (N_11438,N_7702,N_7774);
xor U11439 (N_11439,N_5387,N_5284);
xnor U11440 (N_11440,N_9995,N_7449);
and U11441 (N_11441,N_5199,N_9718);
nand U11442 (N_11442,N_8393,N_9858);
and U11443 (N_11443,N_7806,N_9203);
and U11444 (N_11444,N_9924,N_7205);
nor U11445 (N_11445,N_8068,N_8984);
nand U11446 (N_11446,N_8220,N_8544);
and U11447 (N_11447,N_7178,N_8749);
nor U11448 (N_11448,N_6675,N_7677);
or U11449 (N_11449,N_5485,N_9415);
xor U11450 (N_11450,N_8481,N_5029);
or U11451 (N_11451,N_6094,N_8699);
nor U11452 (N_11452,N_9207,N_6053);
xor U11453 (N_11453,N_9391,N_6785);
nor U11454 (N_11454,N_7175,N_7663);
or U11455 (N_11455,N_9256,N_6631);
nand U11456 (N_11456,N_6072,N_6894);
nor U11457 (N_11457,N_8454,N_5643);
xor U11458 (N_11458,N_6315,N_9780);
xnor U11459 (N_11459,N_9688,N_5084);
nand U11460 (N_11460,N_9986,N_5456);
xor U11461 (N_11461,N_8474,N_7871);
and U11462 (N_11462,N_6642,N_8712);
xnor U11463 (N_11463,N_7572,N_6488);
xor U11464 (N_11464,N_6122,N_9960);
and U11465 (N_11465,N_9174,N_7640);
nand U11466 (N_11466,N_5409,N_5110);
and U11467 (N_11467,N_9426,N_7581);
xor U11468 (N_11468,N_8134,N_5938);
xnor U11469 (N_11469,N_5650,N_7614);
nand U11470 (N_11470,N_8185,N_6494);
xor U11471 (N_11471,N_6937,N_8086);
nor U11472 (N_11472,N_7248,N_5367);
nor U11473 (N_11473,N_6490,N_8041);
nor U11474 (N_11474,N_8016,N_9429);
nand U11475 (N_11475,N_9583,N_6021);
nand U11476 (N_11476,N_5189,N_8955);
or U11477 (N_11477,N_7093,N_9821);
nor U11478 (N_11478,N_9554,N_9367);
nand U11479 (N_11479,N_9044,N_6375);
nor U11480 (N_11480,N_5613,N_7591);
nand U11481 (N_11481,N_6736,N_8767);
and U11482 (N_11482,N_9159,N_8078);
or U11483 (N_11483,N_5800,N_5158);
nand U11484 (N_11484,N_8885,N_6816);
or U11485 (N_11485,N_9930,N_5073);
nand U11486 (N_11486,N_7808,N_5656);
nor U11487 (N_11487,N_9513,N_6082);
xnor U11488 (N_11488,N_9471,N_8604);
nand U11489 (N_11489,N_9042,N_6120);
xor U11490 (N_11490,N_9048,N_7020);
nor U11491 (N_11491,N_6864,N_9926);
or U11492 (N_11492,N_6239,N_7717);
and U11493 (N_11493,N_9056,N_9911);
and U11494 (N_11494,N_5370,N_6379);
or U11495 (N_11495,N_8484,N_8772);
xor U11496 (N_11496,N_6784,N_9263);
nor U11497 (N_11497,N_6655,N_6873);
nand U11498 (N_11498,N_7333,N_7473);
nand U11499 (N_11499,N_8092,N_6345);
or U11500 (N_11500,N_5679,N_6804);
xor U11501 (N_11501,N_6815,N_8671);
nand U11502 (N_11502,N_7503,N_5885);
nor U11503 (N_11503,N_9334,N_6462);
nand U11504 (N_11504,N_6368,N_6941);
and U11505 (N_11505,N_6125,N_7435);
nor U11506 (N_11506,N_7455,N_8899);
or U11507 (N_11507,N_9385,N_5041);
or U11508 (N_11508,N_9300,N_9928);
nand U11509 (N_11509,N_5552,N_9602);
or U11510 (N_11510,N_5397,N_5796);
nor U11511 (N_11511,N_7954,N_7266);
xnor U11512 (N_11512,N_6529,N_9963);
nor U11513 (N_11513,N_8194,N_5869);
or U11514 (N_11514,N_8319,N_7391);
and U11515 (N_11515,N_7028,N_9258);
and U11516 (N_11516,N_6637,N_7140);
and U11517 (N_11517,N_7594,N_6224);
and U11518 (N_11518,N_6206,N_5253);
and U11519 (N_11519,N_5563,N_9006);
xnor U11520 (N_11520,N_8492,N_7803);
and U11521 (N_11521,N_6817,N_8891);
nor U11522 (N_11522,N_6846,N_7858);
xor U11523 (N_11523,N_7284,N_8180);
xor U11524 (N_11524,N_7669,N_6398);
nor U11525 (N_11525,N_7133,N_7651);
nand U11526 (N_11526,N_9474,N_7021);
nor U11527 (N_11527,N_7978,N_9114);
nand U11528 (N_11528,N_7923,N_7939);
nand U11529 (N_11529,N_8986,N_9200);
xor U11530 (N_11530,N_7417,N_8163);
nor U11531 (N_11531,N_7928,N_8172);
and U11532 (N_11532,N_5981,N_7573);
xnor U11533 (N_11533,N_7989,N_7119);
xnor U11534 (N_11534,N_7165,N_5838);
xnor U11535 (N_11535,N_7154,N_7426);
nor U11536 (N_11536,N_6151,N_8248);
nand U11537 (N_11537,N_5578,N_6636);
nor U11538 (N_11538,N_9925,N_8808);
and U11539 (N_11539,N_8141,N_6859);
xnor U11540 (N_11540,N_7185,N_8231);
nor U11541 (N_11541,N_7445,N_8696);
xor U11542 (N_11542,N_6152,N_9145);
xor U11543 (N_11543,N_7788,N_7718);
and U11544 (N_11544,N_9746,N_7818);
nor U11545 (N_11545,N_7664,N_6610);
or U11546 (N_11546,N_5897,N_7204);
nand U11547 (N_11547,N_8289,N_6149);
or U11548 (N_11548,N_7763,N_6401);
nand U11549 (N_11549,N_5962,N_7656);
and U11550 (N_11550,N_9484,N_9892);
and U11551 (N_11551,N_8203,N_5780);
nand U11552 (N_11552,N_9666,N_9133);
xor U11553 (N_11553,N_7092,N_8109);
or U11554 (N_11554,N_8978,N_9803);
nor U11555 (N_11555,N_5205,N_7157);
or U11556 (N_11556,N_9021,N_6822);
nand U11557 (N_11557,N_8768,N_8458);
xor U11558 (N_11558,N_8246,N_7727);
and U11559 (N_11559,N_6423,N_6180);
xor U11560 (N_11560,N_5933,N_7421);
or U11561 (N_11561,N_9632,N_6055);
or U11562 (N_11562,N_5378,N_5644);
and U11563 (N_11563,N_8225,N_9524);
nor U11564 (N_11564,N_7520,N_6725);
nor U11565 (N_11565,N_8670,N_6520);
nand U11566 (N_11566,N_8710,N_9462);
or U11567 (N_11567,N_6914,N_8431);
and U11568 (N_11568,N_7968,N_5916);
and U11569 (N_11569,N_9605,N_9185);
or U11570 (N_11570,N_5004,N_8819);
nand U11571 (N_11571,N_6984,N_5448);
or U11572 (N_11572,N_6200,N_7755);
nand U11573 (N_11573,N_5826,N_7343);
and U11574 (N_11574,N_9461,N_7901);
and U11575 (N_11575,N_5942,N_9702);
nor U11576 (N_11576,N_8813,N_7104);
and U11577 (N_11577,N_9438,N_5821);
nor U11578 (N_11578,N_5883,N_9642);
nor U11579 (N_11579,N_9186,N_5537);
xor U11580 (N_11580,N_5549,N_7723);
nor U11581 (N_11581,N_9343,N_5065);
or U11582 (N_11582,N_7060,N_7311);
nor U11583 (N_11583,N_9722,N_9919);
xnor U11584 (N_11584,N_8001,N_5262);
and U11585 (N_11585,N_8264,N_6098);
and U11586 (N_11586,N_8243,N_6795);
and U11587 (N_11587,N_8776,N_7096);
nor U11588 (N_11588,N_9487,N_8722);
or U11589 (N_11589,N_6011,N_8027);
nor U11590 (N_11590,N_6813,N_9684);
nand U11591 (N_11591,N_8861,N_6392);
xnor U11592 (N_11592,N_8825,N_7387);
nand U11593 (N_11593,N_8967,N_8242);
and U11594 (N_11594,N_9107,N_8994);
and U11595 (N_11595,N_9051,N_8169);
xnor U11596 (N_11596,N_9169,N_6565);
nor U11597 (N_11597,N_9884,N_8133);
nand U11598 (N_11598,N_8102,N_7846);
xor U11599 (N_11599,N_6302,N_7486);
nor U11600 (N_11600,N_6027,N_7608);
xnor U11601 (N_11601,N_7009,N_6247);
xnor U11602 (N_11602,N_7181,N_8055);
nand U11603 (N_11603,N_8963,N_5702);
or U11604 (N_11604,N_5402,N_9653);
xnor U11605 (N_11605,N_8388,N_7779);
or U11606 (N_11606,N_6677,N_8445);
xnor U11607 (N_11607,N_6341,N_7832);
xnor U11608 (N_11608,N_5740,N_8856);
nand U11609 (N_11609,N_8610,N_9572);
xor U11610 (N_11610,N_8979,N_5469);
xor U11611 (N_11611,N_5694,N_5009);
nor U11612 (N_11612,N_6769,N_6900);
or U11613 (N_11613,N_7713,N_5652);
xor U11614 (N_11614,N_9076,N_7252);
nand U11615 (N_11615,N_5052,N_7896);
nor U11616 (N_11616,N_5896,N_8493);
xnor U11617 (N_11617,N_5514,N_9139);
nand U11618 (N_11618,N_7467,N_8087);
nand U11619 (N_11619,N_8301,N_8467);
nor U11620 (N_11620,N_5638,N_6603);
or U11621 (N_11621,N_9968,N_5197);
xor U11622 (N_11622,N_5543,N_7332);
or U11623 (N_11623,N_9778,N_6487);
xnor U11624 (N_11624,N_5489,N_6142);
or U11625 (N_11625,N_6963,N_8973);
xnor U11626 (N_11626,N_6502,N_8083);
nand U11627 (N_11627,N_8159,N_6334);
nand U11628 (N_11628,N_6716,N_9853);
nand U11629 (N_11629,N_7183,N_8192);
or U11630 (N_11630,N_6570,N_9030);
xor U11631 (N_11631,N_9820,N_5550);
or U11632 (N_11632,N_5768,N_6994);
xor U11633 (N_11633,N_9874,N_5614);
xor U11634 (N_11634,N_8317,N_7275);
nor U11635 (N_11635,N_6760,N_7331);
or U11636 (N_11636,N_5911,N_6460);
xor U11637 (N_11637,N_9041,N_8173);
nor U11638 (N_11638,N_7304,N_8716);
nor U11639 (N_11639,N_5213,N_6211);
xor U11640 (N_11640,N_6544,N_9909);
xnor U11641 (N_11641,N_8020,N_6930);
nand U11642 (N_11642,N_5054,N_7798);
nand U11643 (N_11643,N_8413,N_5680);
nor U11644 (N_11644,N_8760,N_9966);
xnor U11645 (N_11645,N_6141,N_7783);
xor U11646 (N_11646,N_9787,N_6958);
nand U11647 (N_11647,N_6019,N_7637);
nand U11648 (N_11648,N_5117,N_7443);
and U11649 (N_11649,N_7330,N_6378);
and U11650 (N_11650,N_6711,N_6329);
nor U11651 (N_11651,N_8594,N_6254);
and U11652 (N_11652,N_6290,N_7290);
xnor U11653 (N_11653,N_9881,N_5293);
nand U11654 (N_11654,N_8889,N_8713);
or U11655 (N_11655,N_9531,N_9640);
and U11656 (N_11656,N_6756,N_8805);
nand U11657 (N_11657,N_9713,N_8906);
xnor U11658 (N_11658,N_9990,N_9690);
nand U11659 (N_11659,N_9763,N_5062);
and U11660 (N_11660,N_8603,N_6267);
nand U11661 (N_11661,N_7282,N_5703);
nand U11662 (N_11662,N_8188,N_9896);
and U11663 (N_11663,N_8981,N_7895);
xor U11664 (N_11664,N_8003,N_9190);
nor U11665 (N_11665,N_6620,N_5633);
nand U11666 (N_11666,N_7326,N_9413);
nand U11667 (N_11667,N_5590,N_7458);
xnor U11668 (N_11668,N_6400,N_7142);
nor U11669 (N_11669,N_5979,N_8935);
nand U11670 (N_11670,N_7696,N_7045);
nand U11671 (N_11671,N_8971,N_5672);
nand U11672 (N_11672,N_8894,N_5571);
xnor U11673 (N_11673,N_5524,N_6102);
xor U11674 (N_11674,N_9998,N_9033);
xor U11675 (N_11675,N_5818,N_9976);
nor U11676 (N_11676,N_6872,N_5473);
and U11677 (N_11677,N_5728,N_5265);
and U11678 (N_11678,N_7604,N_7218);
and U11679 (N_11679,N_8327,N_5646);
xnor U11680 (N_11680,N_6162,N_8953);
xnor U11681 (N_11681,N_7625,N_7612);
xor U11682 (N_11682,N_9314,N_7875);
xor U11683 (N_11683,N_6118,N_5882);
nand U11684 (N_11684,N_8240,N_5132);
and U11685 (N_11685,N_8735,N_8887);
and U11686 (N_11686,N_6234,N_9209);
or U11687 (N_11687,N_5538,N_8636);
nand U11688 (N_11688,N_8391,N_8752);
nand U11689 (N_11689,N_8168,N_8606);
nor U11690 (N_11690,N_8077,N_9581);
nand U11691 (N_11691,N_9151,N_5237);
nand U11692 (N_11692,N_8804,N_6426);
xor U11693 (N_11693,N_5381,N_5769);
or U11694 (N_11694,N_7729,N_9126);
nand U11695 (N_11695,N_5970,N_6510);
or U11696 (N_11696,N_7075,N_8949);
xor U11697 (N_11697,N_8152,N_9236);
or U11698 (N_11698,N_8924,N_5926);
nor U11699 (N_11699,N_8850,N_6217);
or U11700 (N_11700,N_7722,N_6175);
nor U11701 (N_11701,N_8386,N_9576);
nand U11702 (N_11702,N_5951,N_7861);
xnor U11703 (N_11703,N_6449,N_5447);
nor U11704 (N_11704,N_5905,N_5501);
xnor U11705 (N_11705,N_6387,N_8794);
xor U11706 (N_11706,N_8390,N_7720);
nor U11707 (N_11707,N_9443,N_9812);
nor U11708 (N_11708,N_6000,N_6190);
or U11709 (N_11709,N_5389,N_9636);
nand U11710 (N_11710,N_8919,N_6955);
and U11711 (N_11711,N_6308,N_6010);
nand U11712 (N_11712,N_6619,N_5902);
nor U11713 (N_11713,N_6691,N_6629);
xor U11714 (N_11714,N_7377,N_6638);
and U11715 (N_11715,N_5399,N_6573);
and U11716 (N_11716,N_8063,N_9655);
nand U11717 (N_11717,N_7047,N_7687);
nand U11718 (N_11718,N_8509,N_6585);
nor U11719 (N_11719,N_6666,N_7711);
and U11720 (N_11720,N_8505,N_9800);
and U11721 (N_11721,N_5976,N_7050);
xor U11722 (N_11722,N_7390,N_6548);
or U11723 (N_11723,N_5608,N_6212);
and U11724 (N_11724,N_8211,N_9168);
nand U11725 (N_11725,N_9368,N_6491);
nor U11726 (N_11726,N_6626,N_6830);
xnor U11727 (N_11727,N_7596,N_7288);
and U11728 (N_11728,N_8611,N_9468);
or U11729 (N_11729,N_8923,N_5146);
xor U11730 (N_11730,N_5675,N_9295);
or U11731 (N_11731,N_8260,N_5341);
or U11732 (N_11732,N_8824,N_8720);
and U11733 (N_11733,N_5320,N_7900);
nor U11734 (N_11734,N_7065,N_5222);
and U11735 (N_11735,N_8736,N_8601);
or U11736 (N_11736,N_7327,N_5229);
nor U11737 (N_11737,N_6796,N_5328);
and U11738 (N_11738,N_7345,N_7969);
nor U11739 (N_11739,N_5270,N_9062);
nor U11740 (N_11740,N_9829,N_6558);
nand U11741 (N_11741,N_5691,N_6717);
xor U11742 (N_11742,N_9682,N_7671);
or U11743 (N_11743,N_8501,N_8070);
or U11744 (N_11744,N_6648,N_5388);
nor U11745 (N_11745,N_8309,N_7568);
nand U11746 (N_11746,N_5790,N_9731);
nor U11747 (N_11747,N_5186,N_8256);
nor U11748 (N_11748,N_9831,N_6949);
nand U11749 (N_11749,N_5836,N_8680);
nor U11750 (N_11750,N_9208,N_7066);
and U11751 (N_11751,N_9231,N_5336);
nand U11752 (N_11752,N_5718,N_5958);
nand U11753 (N_11753,N_8968,N_8838);
and U11754 (N_11754,N_6103,N_9227);
or U11755 (N_11755,N_6761,N_7852);
or U11756 (N_11756,N_8758,N_6129);
xor U11757 (N_11757,N_9648,N_8558);
xor U11758 (N_11758,N_7363,N_5374);
or U11759 (N_11759,N_6236,N_8004);
or U11760 (N_11760,N_6300,N_9501);
nand U11761 (N_11761,N_5171,N_5444);
nor U11762 (N_11762,N_7040,N_6670);
xnor U11763 (N_11763,N_6022,N_7199);
xnor U11764 (N_11764,N_9970,N_5170);
and U11765 (N_11765,N_7691,N_9770);
xnor U11766 (N_11766,N_8999,N_7764);
nand U11767 (N_11767,N_6985,N_9736);
nor U11768 (N_11768,N_8545,N_6961);
xnor U11769 (N_11769,N_6203,N_8050);
or U11770 (N_11770,N_6440,N_8104);
nor U11771 (N_11771,N_6786,N_5034);
nand U11772 (N_11772,N_5531,N_8273);
and U11773 (N_11773,N_8747,N_8962);
nand U11774 (N_11774,N_8465,N_9650);
or U11775 (N_11775,N_6268,N_6274);
and U11776 (N_11776,N_7409,N_6556);
or U11777 (N_11777,N_7064,N_7632);
and U11778 (N_11778,N_7463,N_9765);
xor U11779 (N_11779,N_5734,N_6682);
nor U11780 (N_11780,N_6940,N_8496);
xor U11781 (N_11781,N_7226,N_8278);
nand U11782 (N_11782,N_7955,N_6714);
nand U11783 (N_11783,N_8355,N_7023);
or U11784 (N_11784,N_6908,N_5165);
and U11785 (N_11785,N_5366,N_6157);
and U11786 (N_11786,N_5106,N_6008);
or U11787 (N_11787,N_9270,N_5795);
and U11788 (N_11788,N_5317,N_9698);
nor U11789 (N_11789,N_9410,N_8621);
nor U11790 (N_11790,N_6774,N_6242);
or U11791 (N_11791,N_9191,N_5311);
nand U11792 (N_11792,N_5529,N_9397);
and U11793 (N_11793,N_6292,N_7530);
and U11794 (N_11794,N_8721,N_7171);
nand U11795 (N_11795,N_9182,N_7265);
or U11796 (N_11796,N_5610,N_7873);
nor U11797 (N_11797,N_9720,N_8913);
xnor U11798 (N_11798,N_7174,N_5944);
and U11799 (N_11799,N_7452,N_5188);
and U11800 (N_11800,N_5941,N_9886);
and U11801 (N_11801,N_5789,N_5283);
and U11802 (N_11802,N_6537,N_6867);
and U11803 (N_11803,N_8384,N_7428);
and U11804 (N_11804,N_7260,N_5458);
and U11805 (N_11805,N_5515,N_7169);
nand U11806 (N_11806,N_9917,N_9025);
and U11807 (N_11807,N_7094,N_9838);
xor U11808 (N_11808,N_6325,N_5519);
and U11809 (N_11809,N_7460,N_8479);
nor U11810 (N_11810,N_5784,N_6260);
or U11811 (N_11811,N_7569,N_5134);
xor U11812 (N_11812,N_9326,N_7631);
and U11813 (N_11813,N_6826,N_7158);
and U11814 (N_11814,N_7480,N_9923);
or U11815 (N_11815,N_5560,N_7109);
xor U11816 (N_11816,N_8113,N_9422);
and U11817 (N_11817,N_7294,N_7683);
or U11818 (N_11818,N_9674,N_7760);
and U11819 (N_11819,N_5946,N_6831);
or U11820 (N_11820,N_8624,N_8177);
nor U11821 (N_11821,N_5346,N_6768);
or U11822 (N_11822,N_5151,N_6169);
nor U11823 (N_11823,N_9578,N_6448);
xor U11824 (N_11824,N_7214,N_9134);
or U11825 (N_11825,N_7127,N_5880);
nand U11826 (N_11826,N_9432,N_5376);
nor U11827 (N_11827,N_8637,N_7629);
nand U11828 (N_11828,N_5793,N_8943);
or U11829 (N_11829,N_5978,N_6397);
and U11830 (N_11830,N_8839,N_5500);
xnor U11831 (N_11831,N_8669,N_6371);
and U11832 (N_11832,N_6550,N_7160);
and U11833 (N_11833,N_6172,N_5698);
or U11834 (N_11834,N_8572,N_6723);
nand U11835 (N_11835,N_8271,N_9204);
and U11836 (N_11836,N_7319,N_9122);
or U11837 (N_11837,N_7151,N_5164);
nand U11838 (N_11838,N_6170,N_8693);
nand U11839 (N_11839,N_7212,N_5959);
xor U11840 (N_11840,N_9878,N_6589);
or U11841 (N_11841,N_6369,N_8089);
nand U11842 (N_11842,N_8405,N_8512);
and U11843 (N_11843,N_5377,N_6304);
nor U11844 (N_11844,N_6732,N_5648);
or U11845 (N_11845,N_9562,N_7351);
nand U11846 (N_11846,N_9049,N_5509);
nand U11847 (N_11847,N_7653,N_7291);
nand U11848 (N_11848,N_5995,N_7202);
and U11849 (N_11849,N_8300,N_7712);
nand U11850 (N_11850,N_6590,N_5339);
and U11851 (N_11851,N_6885,N_9536);
and U11852 (N_11852,N_7000,N_5964);
nor U11853 (N_11853,N_8795,N_6147);
or U11854 (N_11854,N_9233,N_8951);
nor U11855 (N_11855,N_9700,N_9540);
or U11856 (N_11856,N_8858,N_9766);
nand U11857 (N_11857,N_9246,N_5006);
and U11858 (N_11858,N_7469,N_9455);
and U11859 (N_11859,N_8197,N_8524);
or U11860 (N_11860,N_6492,N_8820);
nand U11861 (N_11861,N_6079,N_5460);
xnor U11862 (N_11862,N_6509,N_8863);
or U11863 (N_11863,N_8592,N_9717);
and U11864 (N_11864,N_8284,N_8970);
nand U11865 (N_11865,N_8600,N_7493);
nand U11866 (N_11866,N_6676,N_8803);
nor U11867 (N_11867,N_6511,N_9974);
xnor U11868 (N_11868,N_8121,N_6856);
and U11869 (N_11869,N_9585,N_9489);
nand U11870 (N_11870,N_6493,N_6384);
or U11871 (N_11871,N_5233,N_7851);
xor U11872 (N_11872,N_8877,N_7709);
xnor U11873 (N_11873,N_5403,N_9120);
or U11874 (N_11874,N_9317,N_9375);
xnor U11875 (N_11875,N_8276,N_5637);
and U11876 (N_11876,N_5241,N_7527);
nand U11877 (N_11877,N_8181,N_6355);
xnor U11878 (N_11878,N_5943,N_9170);
and U11879 (N_11879,N_8202,N_5214);
and U11880 (N_11880,N_5201,N_5670);
xor U11881 (N_11881,N_9260,N_5477);
xor U11882 (N_11882,N_6586,N_7583);
or U11883 (N_11883,N_8207,N_9575);
and U11884 (N_11884,N_8743,N_5753);
nor U11885 (N_11885,N_8663,N_5466);
nand U11886 (N_11886,N_7125,N_6319);
or U11887 (N_11887,N_9588,N_7322);
and U11888 (N_11888,N_5335,N_8130);
and U11889 (N_11889,N_9804,N_6261);
and U11890 (N_11890,N_6684,N_9685);
or U11891 (N_11891,N_8907,N_8323);
and U11892 (N_11892,N_8137,N_7216);
nor U11893 (N_11893,N_7156,N_7866);
and U11894 (N_11894,N_7210,N_7492);
or U11895 (N_11895,N_7308,N_7307);
or U11896 (N_11896,N_7303,N_5361);
nand U11897 (N_11897,N_9393,N_5330);
nor U11898 (N_11898,N_5966,N_7451);
nand U11899 (N_11899,N_7138,N_6433);
nand U11900 (N_11900,N_7870,N_7147);
and U11901 (N_11901,N_5192,N_7444);
and U11902 (N_11902,N_6420,N_7627);
nor U11903 (N_11903,N_6975,N_6672);
nor U11904 (N_11904,N_7862,N_9340);
and U11905 (N_11905,N_9196,N_5870);
nor U11906 (N_11906,N_8883,N_7822);
or U11907 (N_11907,N_7339,N_6915);
and U11908 (N_11908,N_6093,N_5027);
nor U11909 (N_11909,N_7032,N_8455);
nand U11910 (N_11910,N_9337,N_8318);
or U11911 (N_11911,N_6279,N_5003);
or U11912 (N_11912,N_9104,N_7562);
nor U11913 (N_11913,N_6215,N_8415);
xnor U11914 (N_11914,N_8831,N_8287);
xor U11915 (N_11915,N_9582,N_5260);
nor U11916 (N_11916,N_8490,N_5415);
nand U11917 (N_11917,N_5147,N_6497);
or U11918 (N_11918,N_6624,N_9637);
and U11919 (N_11919,N_5300,N_9836);
and U11920 (N_11920,N_9703,N_9274);
or U11921 (N_11921,N_8073,N_9026);
or U11922 (N_11922,N_9176,N_6596);
xor U11923 (N_11923,N_9047,N_9321);
xor U11924 (N_11924,N_5212,N_7287);
or U11925 (N_11925,N_8360,N_8814);
and U11926 (N_11926,N_9691,N_9237);
or U11927 (N_11927,N_7842,N_8335);
nand U11928 (N_11928,N_8191,N_8381);
nor U11929 (N_11929,N_5209,N_8741);
nor U11930 (N_11930,N_7239,N_6969);
xnor U11931 (N_11931,N_7521,N_8067);
or U11932 (N_11932,N_5927,N_9625);
nor U11933 (N_11933,N_9593,N_8701);
and U11934 (N_11934,N_7209,N_7438);
nor U11935 (N_11935,N_7833,N_5095);
nor U11936 (N_11936,N_8042,N_5180);
or U11937 (N_11937,N_6634,N_9013);
and U11938 (N_11938,N_5716,N_6337);
or U11939 (N_11939,N_8555,N_8533);
or U11940 (N_11940,N_8860,N_9876);
nand U11941 (N_11941,N_9996,N_9214);
or U11942 (N_11942,N_5999,N_8261);
nor U11943 (N_11943,N_8708,N_9563);
or U11944 (N_11944,N_9694,N_6101);
nand U11945 (N_11945,N_6628,N_6726);
nor U11946 (N_11946,N_6718,N_5910);
xor U11947 (N_11947,N_7085,N_9710);
nand U11948 (N_11948,N_7526,N_7626);
nand U11949 (N_11949,N_5412,N_5427);
or U11950 (N_11950,N_8367,N_8766);
and U11951 (N_11951,N_6782,N_6920);
nand U11952 (N_11952,N_8515,N_6741);
and U11953 (N_11953,N_7122,N_6046);
and U11954 (N_11954,N_5649,N_8204);
nand U11955 (N_11955,N_6588,N_9992);
nand U11956 (N_11956,N_8259,N_7533);
and U11957 (N_11957,N_6932,N_6862);
xnor U11958 (N_11958,N_7433,N_9266);
nand U11959 (N_11959,N_9981,N_6651);
nand U11960 (N_11960,N_9997,N_8620);
and U11961 (N_11961,N_6669,N_7706);
nor U11962 (N_11962,N_9004,N_8510);
nand U11963 (N_11963,N_9206,N_8556);
nand U11964 (N_11964,N_6228,N_9464);
nor U11965 (N_11965,N_7105,N_6265);
xnor U11966 (N_11966,N_5323,N_8387);
nand U11967 (N_11967,N_9927,N_8990);
or U11968 (N_11968,N_7264,N_7247);
nand U11969 (N_11969,N_8478,N_7054);
or U11970 (N_11970,N_9304,N_6933);
nor U11971 (N_11971,N_8784,N_7118);
and U11972 (N_11972,N_5757,N_6579);
and U11973 (N_11973,N_6530,N_8469);
nand U11974 (N_11974,N_5104,N_9511);
or U11975 (N_11975,N_7337,N_8165);
nand U11976 (N_11976,N_5343,N_6365);
nand U11977 (N_11977,N_5822,N_6777);
or U11978 (N_11978,N_5627,N_9546);
or U11979 (N_11979,N_7947,N_8473);
xnor U11980 (N_11980,N_9716,N_7313);
and U11981 (N_11981,N_9604,N_5064);
nand U11982 (N_11982,N_8017,N_6138);
nor U11983 (N_11983,N_6584,N_7659);
xor U11984 (N_11984,N_9008,N_7837);
and U11985 (N_11985,N_8348,N_6210);
nor U11986 (N_11986,N_8252,N_9320);
nand U11987 (N_11987,N_8281,N_9034);
or U11988 (N_11988,N_7101,N_6269);
nand U11989 (N_11989,N_9244,N_7697);
nor U11990 (N_11990,N_6306,N_6734);
and U11991 (N_11991,N_6990,N_6183);
xnor U11992 (N_11992,N_5683,N_9889);
nand U11993 (N_11993,N_8517,N_8049);
xnor U11994 (N_11994,N_6464,N_8853);
or U11995 (N_11995,N_6721,N_8422);
and U11996 (N_11996,N_8324,N_6907);
xor U11997 (N_11997,N_5545,N_5972);
xor U11998 (N_11998,N_8193,N_9488);
nor U11999 (N_11999,N_5231,N_7921);
nand U12000 (N_12000,N_8869,N_8293);
nor U12001 (N_12001,N_8088,N_6434);
or U12002 (N_12002,N_5853,N_9431);
xnor U12003 (N_12003,N_5544,N_5254);
or U12004 (N_12004,N_9538,N_5332);
and U12005 (N_12005,N_7805,N_7620);
xnor U12006 (N_12006,N_9160,N_8835);
and U12007 (N_12007,N_7944,N_8649);
or U12008 (N_12008,N_6204,N_9719);
xor U12009 (N_12009,N_6647,N_7883);
nor U12010 (N_12010,N_7913,N_6699);
or U12011 (N_12011,N_7091,N_5303);
xnor U12012 (N_12012,N_5974,N_6166);
or U12013 (N_12013,N_6310,N_7622);
and U12014 (N_12014,N_7495,N_7299);
or U12015 (N_12015,N_6156,N_6827);
xor U12016 (N_12016,N_5499,N_9866);
xor U12017 (N_12017,N_8008,N_6137);
nor U12018 (N_12018,N_6199,N_8345);
and U12019 (N_12019,N_9424,N_8053);
nor U12020 (N_12020,N_6893,N_8209);
and U12021 (N_12021,N_6431,N_9552);
xnor U12022 (N_12022,N_5792,N_6597);
nand U12023 (N_12023,N_7918,N_5759);
and U12024 (N_12024,N_8040,N_7970);
and U12025 (N_12025,N_8676,N_7001);
nor U12026 (N_12026,N_8936,N_5385);
xnor U12027 (N_12027,N_8790,N_8618);
or U12028 (N_12028,N_8828,N_5513);
nand U12029 (N_12029,N_9565,N_9123);
xor U12030 (N_12030,N_7393,N_7416);
nor U12031 (N_12031,N_6307,N_9396);
nand U12032 (N_12032,N_6587,N_8226);
xnor U12033 (N_12033,N_6618,N_8921);
xnor U12034 (N_12034,N_5809,N_5181);
nor U12035 (N_12035,N_9192,N_5413);
xor U12036 (N_12036,N_6146,N_7432);
nand U12037 (N_12037,N_5445,N_6735);
and U12038 (N_12038,N_8007,N_7557);
and U12039 (N_12039,N_9230,N_5920);
xnor U12040 (N_12040,N_7725,N_6061);
or U12041 (N_12041,N_8740,N_5031);
and U12042 (N_12042,N_5324,N_7897);
nor U12043 (N_12043,N_7477,N_5949);
or U12044 (N_12044,N_7943,N_5161);
nand U12045 (N_12045,N_7812,N_5287);
or U12046 (N_12046,N_8932,N_7256);
xor U12047 (N_12047,N_9066,N_5814);
nand U12048 (N_12048,N_9235,N_6776);
or U12049 (N_12049,N_6145,N_9325);
nand U12050 (N_12050,N_6441,N_9372);
or U12051 (N_12051,N_5548,N_6844);
xor U12052 (N_12052,N_8470,N_6892);
or U12053 (N_12053,N_9984,N_9508);
nand U12054 (N_12054,N_7531,N_7132);
or U12055 (N_12055,N_9723,N_8138);
xor U12056 (N_12056,N_5342,N_8340);
nand U12057 (N_12057,N_7792,N_9704);
nor U12058 (N_12058,N_8363,N_5467);
and U12059 (N_12059,N_7911,N_5565);
nor U12060 (N_12060,N_5263,N_8432);
nor U12061 (N_12061,N_9045,N_7128);
and U12062 (N_12062,N_6159,N_8723);
nand U12063 (N_12063,N_8394,N_7523);
nand U12064 (N_12064,N_9888,N_9987);
nand U12065 (N_12065,N_6353,N_7807);
nand U12066 (N_12066,N_7513,N_9298);
nand U12067 (N_12067,N_6945,N_7099);
nor U12068 (N_12068,N_7089,N_5786);
xnor U12069 (N_12069,N_9234,N_9811);
and U12070 (N_12070,N_6789,N_7575);
and U12071 (N_12071,N_9485,N_9644);
and U12072 (N_12072,N_5977,N_6056);
or U12073 (N_12073,N_5487,N_8059);
nor U12074 (N_12074,N_7325,N_8212);
nand U12075 (N_12075,N_5232,N_9412);
nand U12076 (N_12076,N_9198,N_5892);
or U12077 (N_12077,N_5695,N_8769);
and U12078 (N_12078,N_9105,N_8785);
or U12079 (N_12079,N_7603,N_8342);
nand U12080 (N_12080,N_5647,N_5764);
or U12081 (N_12081,N_5586,N_5898);
nand U12082 (N_12082,N_6073,N_9767);
xnor U12083 (N_12083,N_6096,N_5462);
nand U12084 (N_12084,N_8857,N_7816);
and U12085 (N_12085,N_5411,N_7344);
and U12086 (N_12086,N_5731,N_6663);
nand U12087 (N_12087,N_6773,N_6042);
or U12088 (N_12088,N_8421,N_6733);
and U12089 (N_12089,N_7865,N_9550);
xnor U12090 (N_12090,N_8021,N_8792);
and U12091 (N_12091,N_8589,N_7494);
xor U12092 (N_12092,N_9376,N_6950);
and U12093 (N_12093,N_7229,N_7087);
and U12094 (N_12094,N_8578,N_8504);
nor U12095 (N_12095,N_6536,N_9952);
and U12096 (N_12096,N_9950,N_8779);
nor U12097 (N_12097,N_8374,N_5506);
nand U12098 (N_12098,N_6060,N_6954);
xor U12099 (N_12099,N_9965,N_7012);
and U12100 (N_12100,N_9002,N_5536);
nand U12101 (N_12101,N_7508,N_7179);
xor U12102 (N_12102,N_6679,N_8170);
nand U12103 (N_12103,N_7015,N_5272);
xnor U12104 (N_12104,N_7994,N_6459);
xnor U12105 (N_12105,N_9808,N_6033);
and U12106 (N_12106,N_9797,N_8441);
nand U12107 (N_12107,N_7412,N_6230);
xnor U12108 (N_12108,N_8834,N_8694);
nand U12109 (N_12109,N_6601,N_7617);
and U12110 (N_12110,N_5298,N_9199);
or U12111 (N_12111,N_6673,N_9654);
nor U12112 (N_12112,N_8382,N_6946);
or U12113 (N_12113,N_5331,N_5581);
xor U12114 (N_12114,N_6225,N_8047);
nor U12115 (N_12115,N_9789,N_6697);
and U12116 (N_12116,N_9649,N_7537);
nand U12117 (N_12117,N_7607,N_5576);
or U12118 (N_12118,N_9543,N_8128);
nor U12119 (N_12119,N_6577,N_5701);
xor U12120 (N_12120,N_5099,N_7237);
or U12121 (N_12121,N_6127,N_5913);
xnor U12122 (N_12122,N_8777,N_8221);
or U12123 (N_12123,N_7141,N_6444);
or U12124 (N_12124,N_6906,N_6427);
or U12125 (N_12125,N_5406,N_6739);
xnor U12126 (N_12126,N_8265,N_9251);
and U12127 (N_12127,N_6531,N_7190);
xor U12128 (N_12128,N_8127,N_6051);
or U12129 (N_12129,N_8882,N_7431);
or U12130 (N_12130,N_5875,N_6728);
nor U12131 (N_12131,N_5721,N_9491);
nor U12132 (N_12132,N_9342,N_6132);
or U12133 (N_12133,N_9149,N_5893);
xnor U12134 (N_12134,N_8983,N_9695);
xnor U12135 (N_12135,N_9626,N_8754);
xor U12136 (N_12136,N_9082,N_5794);
xor U12137 (N_12137,N_6911,N_7719);
nand U12138 (N_12138,N_7004,N_7525);
xnor U12139 (N_12139,N_9125,N_8396);
and U12140 (N_12140,N_7317,N_5414);
or U12141 (N_12141,N_8911,N_8039);
and U12142 (N_12142,N_5350,N_6713);
and U12143 (N_12143,N_6276,N_7891);
or U12144 (N_12144,N_9796,N_5540);
or U12145 (N_12145,N_9677,N_9978);
and U12146 (N_12146,N_6875,N_7582);
nand U12147 (N_12147,N_6504,N_8744);
xor U12148 (N_12148,N_5766,N_6364);
or U12149 (N_12149,N_6792,N_6657);
and U12150 (N_12150,N_5450,N_7448);
and U12151 (N_12151,N_6820,N_8397);
nand U12152 (N_12152,N_5152,N_5894);
and U12153 (N_12153,N_7292,N_7376);
xnor U12154 (N_12154,N_7689,N_5705);
xor U12155 (N_12155,N_9547,N_6593);
nand U12156 (N_12156,N_7465,N_7145);
nand U12157 (N_12157,N_7233,N_7976);
nand U12158 (N_12158,N_7501,N_6944);
nand U12159 (N_12159,N_8066,N_6430);
nand U12160 (N_12160,N_7415,N_8656);
or U12161 (N_12161,N_7886,N_8833);
nor U12162 (N_12162,N_7854,N_8786);
or U12163 (N_12163,N_5175,N_6525);
and U12164 (N_12164,N_5762,N_8667);
or U12165 (N_12165,N_7168,N_8539);
nand U12166 (N_12166,N_8989,N_8681);
nor U12167 (N_12167,N_8119,N_9401);
xnor U12168 (N_12168,N_5314,N_6481);
or U12169 (N_12169,N_9851,N_7790);
and U12170 (N_12170,N_6605,N_6409);
xnor U12171 (N_12171,N_9728,N_8778);
nand U12172 (N_12172,N_8516,N_9418);
or U12173 (N_12173,N_8818,N_5478);
xor U12174 (N_12174,N_7912,N_6229);
nand U12175 (N_12175,N_5700,N_9179);
nand U12176 (N_12176,N_6708,N_9003);
nor U12177 (N_12177,N_9549,N_7668);
and U12178 (N_12178,N_6038,N_7633);
or U12179 (N_12179,N_9822,N_7230);
nor U12180 (N_12180,N_7249,N_6899);
and U12181 (N_12181,N_6417,N_5923);
nor U12182 (N_12182,N_8523,N_5990);
nor U12183 (N_12183,N_7868,N_5082);
or U12184 (N_12184,N_8527,N_7910);
nand U12185 (N_12185,N_5086,N_6167);
nand U12186 (N_12186,N_9181,N_8205);
xnor U12187 (N_12187,N_7902,N_8855);
nand U12188 (N_12188,N_7823,N_9111);
nand U12189 (N_12189,N_9845,N_6366);
xor U12190 (N_12190,N_8029,N_6695);
and U12191 (N_12191,N_8438,N_9743);
and U12192 (N_12192,N_5391,N_8750);
nand U12193 (N_12193,N_7370,N_5517);
nand U12194 (N_12194,N_8789,N_8862);
nand U12195 (N_12195,N_7904,N_9212);
or U12196 (N_12196,N_9486,N_8635);
or U12197 (N_12197,N_9352,N_7155);
or U12198 (N_12198,N_9852,N_8893);
xnor U12199 (N_12199,N_8368,N_5280);
nor U12200 (N_12200,N_9857,N_7270);
nor U12201 (N_12201,N_5900,N_8034);
xor U12202 (N_12202,N_6615,N_8679);
and U12203 (N_12203,N_7860,N_8674);
and U12204 (N_12204,N_9558,N_5418);
nor U12205 (N_12205,N_7211,N_8101);
or U12206 (N_12206,N_5612,N_8062);
xor U12207 (N_12207,N_9063,N_9993);
and U12208 (N_12208,N_5937,N_8296);
xnor U12209 (N_12209,N_5433,N_5887);
or U12210 (N_12210,N_6868,N_5969);
nand U12211 (N_12211,N_7937,N_7359);
nor U12212 (N_12212,N_9883,N_8929);
or U12213 (N_12213,N_7350,N_5139);
or U12214 (N_12214,N_6567,N_5051);
and U12215 (N_12215,N_6470,N_5975);
nand U12216 (N_12216,N_9922,N_6569);
nor U12217 (N_12217,N_9668,N_9303);
or U12218 (N_12218,N_5603,N_5555);
xor U12219 (N_12219,N_5404,N_8339);
nor U12220 (N_12220,N_6223,N_6406);
and U12221 (N_12221,N_6432,N_6408);
nand U12222 (N_12222,N_9363,N_5368);
xnor U12223 (N_12223,N_5319,N_6278);
xor U12224 (N_12224,N_8920,N_8569);
xor U12225 (N_12225,N_5782,N_9832);
or U12226 (N_12226,N_6062,N_5459);
or U12227 (N_12227,N_8609,N_7110);
nand U12228 (N_12228,N_7459,N_6095);
nand U12229 (N_12229,N_8954,N_8241);
nor U12230 (N_12230,N_5482,N_6074);
or U12231 (N_12231,N_8054,N_7372);
nand U12232 (N_12232,N_5178,N_5256);
nand U12233 (N_12233,N_5577,N_7187);
nor U12234 (N_12234,N_9193,N_8602);
nor U12235 (N_12235,N_5495,N_7899);
or U12236 (N_12236,N_9316,N_5441);
and U12237 (N_12237,N_5185,N_6330);
or U12238 (N_12238,N_7908,N_5157);
xnor U12239 (N_12239,N_9016,N_9088);
nand U12240 (N_12240,N_7974,N_8788);
xnor U12241 (N_12241,N_8673,N_7898);
nand U12242 (N_12242,N_9148,N_6686);
nor U12243 (N_12243,N_9793,N_8311);
xnor U12244 (N_12244,N_9835,N_6480);
or U12245 (N_12245,N_9419,N_5279);
nor U12246 (N_12246,N_6385,N_5929);
or U12247 (N_12247,N_8513,N_6609);
nand U12248 (N_12248,N_9427,N_8149);
nand U12249 (N_12249,N_8866,N_9551);
or U12250 (N_12250,N_6881,N_7840);
nand U12251 (N_12251,N_7652,N_5819);
xnor U12252 (N_12252,N_5011,N_5100);
and U12253 (N_12253,N_7502,N_9306);
and U12254 (N_12254,N_9747,N_8215);
nor U12255 (N_12255,N_5138,N_6327);
nand U12256 (N_12256,N_7394,N_7106);
or U12257 (N_12257,N_6580,N_5640);
and U12258 (N_12258,N_9783,N_9072);
or U12259 (N_12259,N_8675,N_6818);
or U12260 (N_12260,N_6089,N_8822);
or U12261 (N_12261,N_7675,N_7374);
nor U12262 (N_12262,N_7967,N_8625);
xnor U12263 (N_12263,N_8258,N_9764);
nor U12264 (N_12264,N_7560,N_6252);
and U12265 (N_12265,N_7043,N_6668);
nand U12266 (N_12266,N_9561,N_9113);
nor U12267 (N_12267,N_7869,N_5305);
nor U12268 (N_12268,N_8665,N_9680);
or U12269 (N_12269,N_5243,N_6779);
xor U12270 (N_12270,N_6014,N_9810);
nand U12271 (N_12271,N_6654,N_9813);
and U12272 (N_12272,N_9240,N_8746);
nor U12273 (N_12273,N_9380,N_6890);
nand U12274 (N_12274,N_9955,N_7484);
and U12275 (N_12275,N_5866,N_5013);
and U12276 (N_12276,N_6918,N_7505);
xor U12277 (N_12277,N_5697,N_9614);
nor U12278 (N_12278,N_8357,N_8896);
and U12279 (N_12279,N_9873,N_7364);
and U12280 (N_12280,N_5497,N_8842);
nand U12281 (N_12281,N_6753,N_6506);
or U12282 (N_12282,N_7454,N_7756);
nand U12283 (N_12283,N_9449,N_8677);
nand U12284 (N_12284,N_7153,N_5453);
nor U12285 (N_12285,N_8466,N_7934);
nand U12286 (N_12286,N_7528,N_8683);
nor U12287 (N_12287,N_6746,N_8543);
nor U12288 (N_12288,N_6003,N_9751);
or U12289 (N_12289,N_5075,N_9059);
or U12290 (N_12290,N_8430,N_7958);
nand U12291 (N_12291,N_9956,N_7038);
nand U12292 (N_12292,N_5093,N_8689);
nand U12293 (N_12293,N_5717,N_7826);
nand U12294 (N_12294,N_7948,N_8011);
xor U12295 (N_12295,N_6222,N_9931);
xnor U12296 (N_12296,N_7220,N_8218);
nor U12297 (N_12297,N_5191,N_7207);
xnor U12298 (N_12298,N_6828,N_8950);
and U12299 (N_12299,N_7536,N_7879);
nand U12300 (N_12300,N_5621,N_7639);
xnor U12301 (N_12301,N_8448,N_7731);
xnor U12302 (N_12302,N_6476,N_6477);
and U12303 (N_12303,N_9106,N_6980);
or U12304 (N_12304,N_7759,N_6294);
nand U12305 (N_12305,N_8583,N_6851);
nor U12306 (N_12306,N_5016,N_6805);
xor U12307 (N_12307,N_5408,N_7440);
nand U12308 (N_12308,N_8815,N_7076);
or U12309 (N_12309,N_5745,N_6193);
and U12310 (N_12310,N_7227,N_6289);
nand U12311 (N_12311,N_9699,N_8836);
nand U12312 (N_12312,N_9378,N_5632);
or U12313 (N_12313,N_7714,N_8352);
or U12314 (N_12314,N_5037,N_6623);
or U12315 (N_12315,N_5661,N_5561);
nand U12316 (N_12316,N_9520,N_8585);
nor U12317 (N_12317,N_6943,N_9859);
and U12318 (N_12318,N_6542,N_7051);
and U12319 (N_12319,N_5187,N_5788);
and U12320 (N_12320,N_6683,N_7684);
xnor U12321 (N_12321,N_9138,N_7309);
and U12322 (N_12322,N_8707,N_9288);
xor U12323 (N_12323,N_8765,N_6213);
or U12324 (N_12324,N_9147,N_5357);
xnor U12325 (N_12325,N_9994,N_7942);
xnor U12326 (N_12326,N_6909,N_9194);
xnor U12327 (N_12327,N_9825,N_6643);
nand U12328 (N_12328,N_6109,N_6414);
xor U12329 (N_12329,N_6611,N_9257);
nand U12330 (N_12330,N_9128,N_7037);
or U12331 (N_12331,N_5510,N_5080);
and U12332 (N_12332,N_6339,N_6919);
and U12333 (N_12333,N_8019,N_8597);
nor U12334 (N_12334,N_7186,N_6575);
or U12335 (N_12335,N_8337,N_6771);
or U12336 (N_12336,N_7888,N_8607);
or U12337 (N_12337,N_5021,N_6656);
xnor U12338 (N_12338,N_9624,N_5735);
xnor U12339 (N_12339,N_9785,N_5761);
or U12340 (N_12340,N_9577,N_5017);
xnor U12341 (N_12341,N_8196,N_9446);
xnor U12342 (N_12342,N_9245,N_7646);
nand U12343 (N_12343,N_8142,N_8013);
nand U12344 (N_12344,N_6662,N_6895);
nand U12345 (N_12345,N_7820,N_8859);
nor U12346 (N_12346,N_8108,N_8832);
or U12347 (N_12347,N_8100,N_5580);
nor U12348 (N_12348,N_9173,N_5285);
nand U12349 (N_12349,N_6295,N_9856);
or U12350 (N_12350,N_9860,N_6347);
and U12351 (N_12351,N_8996,N_7069);
nor U12352 (N_12352,N_9634,N_7462);
nand U12353 (N_12353,N_5840,N_5857);
nor U12354 (N_12354,N_8423,N_9117);
xor U12355 (N_12355,N_7476,N_6043);
nor U12356 (N_12356,N_6437,N_6681);
xnor U12357 (N_12357,N_6917,N_5127);
and U12358 (N_12358,N_7318,N_9119);
and U12359 (N_12359,N_5491,N_9210);
and U12360 (N_12360,N_8593,N_5060);
and U12361 (N_12361,N_8982,N_7413);
or U12362 (N_12362,N_6685,N_9096);
and U12363 (N_12363,N_6794,N_8537);
nand U12364 (N_12364,N_6270,N_9250);
or U12365 (N_12365,N_9167,N_9039);
xor U12366 (N_12366,N_6976,N_8559);
or U12367 (N_12367,N_7420,N_7300);
nand U12368 (N_12368,N_7791,N_5512);
nand U12369 (N_12369,N_8717,N_5288);
nand U12370 (N_12370,N_6762,N_5215);
nand U12371 (N_12371,N_7225,N_8294);
and U12372 (N_12372,N_8532,N_5429);
nor U12373 (N_12373,N_6838,N_8359);
xor U12374 (N_12374,N_8586,N_8320);
nor U12375 (N_12375,N_6882,N_8277);
or U12376 (N_12376,N_7086,N_8972);
nor U12377 (N_12377,N_8245,N_8380);
and U12378 (N_12378,N_9643,N_6988);
nor U12379 (N_12379,N_5600,N_7234);
xor U12380 (N_12380,N_7120,N_6085);
nor U12381 (N_12381,N_8711,N_9679);
nor U12382 (N_12382,N_8738,N_7519);
and U12383 (N_12383,N_7827,N_9069);
xnor U12384 (N_12384,N_7316,N_5163);
nor U12385 (N_12385,N_9377,N_9594);
nor U12386 (N_12386,N_7024,N_5994);
nand U12387 (N_12387,N_7733,N_6800);
and U12388 (N_12388,N_9664,N_6660);
and U12389 (N_12389,N_5837,N_7246);
nand U12390 (N_12390,N_8107,N_9146);
and U12391 (N_12391,N_6352,N_8546);
xnor U12392 (N_12392,N_6674,N_6128);
and U12393 (N_12393,N_9773,N_9132);
nor U12394 (N_12394,N_6305,N_7193);
nand U12395 (N_12395,N_8251,N_9067);
or U12396 (N_12396,N_6515,N_6130);
nor U12397 (N_12397,N_7373,N_8058);
and U12398 (N_12398,N_9414,N_5227);
nand U12399 (N_12399,N_9332,N_5696);
or U12400 (N_12400,N_6561,N_8112);
xnor U12401 (N_12401,N_5534,N_5090);
nand U12402 (N_12402,N_8129,N_9330);
nand U12403 (N_12403,N_6301,N_5934);
nor U12404 (N_12404,N_8841,N_5917);
xnor U12405 (N_12405,N_8799,N_9211);
nor U12406 (N_12406,N_6901,N_7383);
or U12407 (N_12407,N_5310,N_9475);
and U12408 (N_12408,N_8763,N_5114);
or U12409 (N_12409,N_8685,N_9503);
nand U12410 (N_12410,N_5909,N_8249);
or U12411 (N_12411,N_9754,N_7510);
or U12412 (N_12412,N_5858,N_7007);
nand U12413 (N_12413,N_6562,N_5708);
xnor U12414 (N_12414,N_8279,N_9880);
xnor U12415 (N_12415,N_6412,N_6540);
and U12416 (N_12416,N_5868,N_8798);
or U12417 (N_12417,N_7882,N_7078);
or U12418 (N_12418,N_7987,N_5930);
and U12419 (N_12419,N_8257,N_8737);
nor U12420 (N_12420,N_6324,N_8538);
or U12421 (N_12421,N_5276,N_9318);
xnor U12422 (N_12422,N_6178,N_7305);
nor U12423 (N_12423,N_5390,N_6633);
or U12424 (N_12424,N_7090,N_9844);
or U12425 (N_12425,N_9012,N_9496);
xor U12426 (N_12426,N_5020,N_5204);
xor U12427 (N_12427,N_8865,N_5105);
and U12428 (N_12428,N_5751,N_8682);
or U12429 (N_12429,N_5498,N_6452);
nand U12430 (N_12430,N_5267,N_7565);
or U12431 (N_12431,N_8645,N_7863);
nor U12432 (N_12432,N_5527,N_9411);
xnor U12433 (N_12433,N_6438,N_9947);
nand U12434 (N_12434,N_6077,N_5901);
xnor U12435 (N_12435,N_6273,N_9595);
and U12436 (N_12436,N_5750,N_9502);
nor U12437 (N_12437,N_9157,N_6841);
nand U12438 (N_12438,N_6829,N_5468);
or U12439 (N_12439,N_7070,N_5492);
xnor U12440 (N_12440,N_8213,N_6070);
nor U12441 (N_12441,N_9452,N_5863);
or U12442 (N_12442,N_9545,N_7191);
or U12443 (N_12443,N_6842,N_6997);
or U12444 (N_12444,N_8416,N_9336);
xnor U12445 (N_12445,N_8476,N_9404);
nor U12446 (N_12446,N_8334,N_6150);
or U12447 (N_12447,N_6106,N_9749);
nand U12448 (N_12448,N_5589,N_8703);
nand U12449 (N_12449,N_8485,N_9389);
nand U12450 (N_12450,N_8325,N_6664);
or U12451 (N_12451,N_6108,N_6005);
nor U12452 (N_12452,N_9406,N_6031);
nor U12453 (N_12453,N_7556,N_9131);
or U12454 (N_12454,N_7482,N_8806);
nand U12455 (N_12455,N_9287,N_5005);
or U12456 (N_12456,N_6978,N_9869);
xnor U12457 (N_12457,N_6114,N_9348);
and U12458 (N_12458,N_5033,N_5775);
xor U12459 (N_12459,N_8952,N_5136);
xnor U12460 (N_12460,N_5375,N_8903);
nor U12461 (N_12461,N_8843,N_5416);
or U12462 (N_12462,N_5992,N_7056);
nand U12463 (N_12463,N_9347,N_6148);
or U12464 (N_12464,N_8254,N_5349);
xor U12465 (N_12465,N_5103,N_8014);
nor U12466 (N_12466,N_8522,N_6747);
nand U12467 (N_12467,N_5754,N_5559);
nor U12468 (N_12468,N_5832,N_6187);
nor U12469 (N_12469,N_9331,N_9155);
and U12470 (N_12470,N_8115,N_8897);
xor U12471 (N_12471,N_6197,N_8407);
nor U12472 (N_12472,N_9441,N_7447);
nand U12473 (N_12473,N_7149,N_7048);
xor U12474 (N_12474,N_7877,N_5617);
or U12475 (N_12475,N_8498,N_8038);
or U12476 (N_12476,N_5345,N_5526);
xnor U12477 (N_12477,N_9144,N_7973);
and U12478 (N_12478,N_8918,N_9964);
and U12479 (N_12479,N_5327,N_8184);
or U12480 (N_12480,N_7940,N_9421);
xor U12481 (N_12481,N_5742,N_8571);
and U12482 (N_12482,N_6131,N_5360);
xnor U12483 (N_12483,N_5829,N_7630);
xnor U12484 (N_12484,N_7483,N_7017);
nand U12485 (N_12485,N_7892,N_6886);
nor U12486 (N_12486,N_9281,N_8617);
nand U12487 (N_12487,N_9370,N_9029);
xor U12488 (N_12488,N_9433,N_6705);
or U12489 (N_12489,N_5997,N_7134);
xnor U12490 (N_12490,N_7301,N_9253);
or U12491 (N_12491,N_9610,N_7366);
or U12492 (N_12492,N_9163,N_5061);
and U12493 (N_12493,N_5908,N_9038);
or U12494 (N_12494,N_8051,N_5380);
nor U12495 (N_12495,N_9458,N_6745);
nor U12496 (N_12496,N_9906,N_7355);
and U12497 (N_12497,N_5572,N_5119);
and U12498 (N_12498,N_9658,N_7324);
nor U12499 (N_12499,N_5876,N_6748);
nor U12500 (N_12500,N_7404,N_9429);
nor U12501 (N_12501,N_7508,N_8381);
and U12502 (N_12502,N_8181,N_5873);
nand U12503 (N_12503,N_6602,N_7656);
and U12504 (N_12504,N_6484,N_6731);
and U12505 (N_12505,N_6393,N_9899);
nor U12506 (N_12506,N_8617,N_9624);
nor U12507 (N_12507,N_7972,N_8101);
and U12508 (N_12508,N_8037,N_7035);
xnor U12509 (N_12509,N_8978,N_6071);
and U12510 (N_12510,N_9434,N_6215);
or U12511 (N_12511,N_9496,N_6015);
nand U12512 (N_12512,N_6821,N_6745);
nand U12513 (N_12513,N_7807,N_6936);
and U12514 (N_12514,N_8614,N_6406);
or U12515 (N_12515,N_9612,N_7878);
nor U12516 (N_12516,N_5745,N_8653);
nand U12517 (N_12517,N_6344,N_5559);
and U12518 (N_12518,N_7487,N_5501);
xnor U12519 (N_12519,N_7064,N_6775);
nor U12520 (N_12520,N_6184,N_9131);
nand U12521 (N_12521,N_8407,N_7811);
nand U12522 (N_12522,N_9148,N_9700);
nor U12523 (N_12523,N_5627,N_8871);
nor U12524 (N_12524,N_6085,N_5194);
nand U12525 (N_12525,N_9188,N_8265);
and U12526 (N_12526,N_5506,N_9586);
and U12527 (N_12527,N_7295,N_9850);
and U12528 (N_12528,N_9939,N_5785);
nand U12529 (N_12529,N_7344,N_5318);
nand U12530 (N_12530,N_9128,N_7649);
or U12531 (N_12531,N_5123,N_9814);
nand U12532 (N_12532,N_9944,N_7390);
and U12533 (N_12533,N_5849,N_6419);
or U12534 (N_12534,N_6077,N_9991);
or U12535 (N_12535,N_8324,N_5711);
or U12536 (N_12536,N_6554,N_8685);
nor U12537 (N_12537,N_5765,N_8972);
nand U12538 (N_12538,N_5949,N_8555);
nand U12539 (N_12539,N_6448,N_7075);
or U12540 (N_12540,N_6549,N_6372);
and U12541 (N_12541,N_6253,N_6143);
or U12542 (N_12542,N_8367,N_9874);
and U12543 (N_12543,N_8452,N_6666);
and U12544 (N_12544,N_7186,N_9397);
nor U12545 (N_12545,N_9623,N_8117);
and U12546 (N_12546,N_8365,N_9930);
and U12547 (N_12547,N_7598,N_9265);
xor U12548 (N_12548,N_5706,N_6978);
xnor U12549 (N_12549,N_5169,N_6652);
nor U12550 (N_12550,N_5150,N_9183);
nand U12551 (N_12551,N_9178,N_5045);
nor U12552 (N_12552,N_6651,N_9052);
and U12553 (N_12553,N_7752,N_5563);
nand U12554 (N_12554,N_7702,N_6258);
nor U12555 (N_12555,N_9111,N_6832);
xnor U12556 (N_12556,N_7319,N_6108);
nand U12557 (N_12557,N_7136,N_7998);
xor U12558 (N_12558,N_9735,N_6028);
xor U12559 (N_12559,N_7733,N_6111);
xor U12560 (N_12560,N_6926,N_6993);
and U12561 (N_12561,N_8290,N_7392);
and U12562 (N_12562,N_6303,N_5118);
and U12563 (N_12563,N_6695,N_9034);
or U12564 (N_12564,N_5285,N_8879);
nand U12565 (N_12565,N_5382,N_5728);
or U12566 (N_12566,N_9221,N_7597);
nand U12567 (N_12567,N_8834,N_7507);
xor U12568 (N_12568,N_6637,N_6588);
or U12569 (N_12569,N_5301,N_8755);
or U12570 (N_12570,N_9578,N_8839);
nor U12571 (N_12571,N_8706,N_6594);
xnor U12572 (N_12572,N_5833,N_6694);
and U12573 (N_12573,N_6961,N_6188);
xor U12574 (N_12574,N_5363,N_9718);
and U12575 (N_12575,N_5606,N_8610);
xor U12576 (N_12576,N_9966,N_9821);
xor U12577 (N_12577,N_6695,N_7691);
or U12578 (N_12578,N_6802,N_7479);
xnor U12579 (N_12579,N_5533,N_8381);
or U12580 (N_12580,N_6185,N_5426);
and U12581 (N_12581,N_7491,N_9987);
xnor U12582 (N_12582,N_6918,N_7068);
and U12583 (N_12583,N_6706,N_8431);
or U12584 (N_12584,N_8739,N_6135);
and U12585 (N_12585,N_7252,N_5998);
nand U12586 (N_12586,N_6298,N_8265);
nor U12587 (N_12587,N_9239,N_5255);
nand U12588 (N_12588,N_5739,N_9505);
xnor U12589 (N_12589,N_7993,N_5445);
nand U12590 (N_12590,N_8477,N_5961);
nand U12591 (N_12591,N_7110,N_8441);
nand U12592 (N_12592,N_8562,N_7916);
or U12593 (N_12593,N_5228,N_7162);
xnor U12594 (N_12594,N_9988,N_5430);
or U12595 (N_12595,N_9133,N_9171);
nand U12596 (N_12596,N_8038,N_8591);
and U12597 (N_12597,N_6731,N_8021);
nand U12598 (N_12598,N_6685,N_6139);
nor U12599 (N_12599,N_6764,N_8083);
nor U12600 (N_12600,N_7749,N_8035);
or U12601 (N_12601,N_8311,N_7137);
xnor U12602 (N_12602,N_9445,N_5925);
nor U12603 (N_12603,N_6901,N_6734);
and U12604 (N_12604,N_5946,N_6584);
or U12605 (N_12605,N_7751,N_9142);
xor U12606 (N_12606,N_9246,N_5448);
nor U12607 (N_12607,N_6963,N_5477);
and U12608 (N_12608,N_8173,N_9865);
xor U12609 (N_12609,N_8132,N_5589);
xnor U12610 (N_12610,N_5355,N_7081);
nand U12611 (N_12611,N_5993,N_5785);
nand U12612 (N_12612,N_9479,N_9365);
and U12613 (N_12613,N_8097,N_6098);
xor U12614 (N_12614,N_7305,N_8756);
nor U12615 (N_12615,N_5119,N_7281);
nor U12616 (N_12616,N_6617,N_9550);
xnor U12617 (N_12617,N_5488,N_7973);
nand U12618 (N_12618,N_7926,N_9011);
or U12619 (N_12619,N_5836,N_6081);
xor U12620 (N_12620,N_9132,N_9500);
or U12621 (N_12621,N_9889,N_9908);
or U12622 (N_12622,N_8895,N_8273);
and U12623 (N_12623,N_7457,N_6646);
and U12624 (N_12624,N_6333,N_7260);
or U12625 (N_12625,N_6761,N_5607);
or U12626 (N_12626,N_5974,N_5458);
xor U12627 (N_12627,N_8951,N_9821);
or U12628 (N_12628,N_9120,N_7852);
and U12629 (N_12629,N_9861,N_9626);
nor U12630 (N_12630,N_6476,N_8453);
xnor U12631 (N_12631,N_7508,N_8197);
xor U12632 (N_12632,N_8013,N_9054);
nand U12633 (N_12633,N_9905,N_6096);
and U12634 (N_12634,N_5177,N_9653);
nand U12635 (N_12635,N_8211,N_9937);
and U12636 (N_12636,N_8748,N_6791);
nor U12637 (N_12637,N_8663,N_9578);
and U12638 (N_12638,N_7425,N_8848);
nand U12639 (N_12639,N_6631,N_9910);
xnor U12640 (N_12640,N_7133,N_7239);
xnor U12641 (N_12641,N_6681,N_9194);
nand U12642 (N_12642,N_7430,N_9557);
nand U12643 (N_12643,N_9637,N_5291);
xnor U12644 (N_12644,N_7786,N_6366);
nor U12645 (N_12645,N_5949,N_7070);
or U12646 (N_12646,N_9666,N_8320);
or U12647 (N_12647,N_6260,N_8383);
nand U12648 (N_12648,N_8786,N_7081);
and U12649 (N_12649,N_6148,N_6634);
nor U12650 (N_12650,N_9814,N_5491);
and U12651 (N_12651,N_9831,N_6527);
nand U12652 (N_12652,N_5346,N_9332);
nor U12653 (N_12653,N_9935,N_8772);
nand U12654 (N_12654,N_6617,N_9113);
xor U12655 (N_12655,N_7967,N_9097);
xor U12656 (N_12656,N_6878,N_5007);
or U12657 (N_12657,N_7478,N_5843);
xor U12658 (N_12658,N_7552,N_5408);
xor U12659 (N_12659,N_6774,N_6469);
nor U12660 (N_12660,N_5133,N_6845);
xor U12661 (N_12661,N_6527,N_6928);
nor U12662 (N_12662,N_5943,N_5904);
nand U12663 (N_12663,N_8386,N_8738);
nor U12664 (N_12664,N_6855,N_7485);
xor U12665 (N_12665,N_5261,N_8344);
nand U12666 (N_12666,N_6597,N_9609);
nor U12667 (N_12667,N_8419,N_9618);
xnor U12668 (N_12668,N_9940,N_6323);
and U12669 (N_12669,N_6138,N_7453);
xnor U12670 (N_12670,N_8625,N_6334);
or U12671 (N_12671,N_5174,N_6018);
or U12672 (N_12672,N_6643,N_5840);
and U12673 (N_12673,N_8148,N_6702);
or U12674 (N_12674,N_9126,N_9366);
nand U12675 (N_12675,N_6269,N_6626);
nor U12676 (N_12676,N_9896,N_8433);
and U12677 (N_12677,N_8266,N_8184);
nand U12678 (N_12678,N_9131,N_7473);
nand U12679 (N_12679,N_8596,N_9840);
nand U12680 (N_12680,N_7561,N_8065);
nor U12681 (N_12681,N_9170,N_9828);
and U12682 (N_12682,N_6531,N_5325);
or U12683 (N_12683,N_5675,N_5477);
or U12684 (N_12684,N_6546,N_5716);
nor U12685 (N_12685,N_8985,N_9063);
nor U12686 (N_12686,N_7734,N_6752);
or U12687 (N_12687,N_7461,N_9831);
xnor U12688 (N_12688,N_9306,N_6261);
or U12689 (N_12689,N_9362,N_7992);
nand U12690 (N_12690,N_6600,N_9695);
xor U12691 (N_12691,N_8370,N_6071);
and U12692 (N_12692,N_8771,N_5597);
and U12693 (N_12693,N_8725,N_9053);
and U12694 (N_12694,N_9967,N_7267);
and U12695 (N_12695,N_8108,N_7789);
xor U12696 (N_12696,N_8319,N_8250);
xor U12697 (N_12697,N_6941,N_5040);
nor U12698 (N_12698,N_8544,N_8048);
nand U12699 (N_12699,N_6868,N_5602);
xor U12700 (N_12700,N_5101,N_6206);
nand U12701 (N_12701,N_6486,N_8543);
nor U12702 (N_12702,N_5340,N_5360);
xnor U12703 (N_12703,N_9241,N_8641);
and U12704 (N_12704,N_5007,N_7208);
xor U12705 (N_12705,N_5046,N_5969);
and U12706 (N_12706,N_7597,N_5031);
nor U12707 (N_12707,N_6812,N_9117);
or U12708 (N_12708,N_8410,N_9732);
nand U12709 (N_12709,N_8392,N_7832);
xor U12710 (N_12710,N_7279,N_8581);
nand U12711 (N_12711,N_5400,N_6940);
and U12712 (N_12712,N_5934,N_5844);
or U12713 (N_12713,N_9229,N_6360);
nor U12714 (N_12714,N_6861,N_5495);
or U12715 (N_12715,N_8167,N_6840);
nand U12716 (N_12716,N_6346,N_6576);
xor U12717 (N_12717,N_5156,N_9602);
nor U12718 (N_12718,N_5476,N_9885);
or U12719 (N_12719,N_9575,N_7516);
nand U12720 (N_12720,N_8162,N_7835);
nor U12721 (N_12721,N_7927,N_5990);
nor U12722 (N_12722,N_7788,N_7317);
and U12723 (N_12723,N_9867,N_5340);
or U12724 (N_12724,N_9548,N_5032);
or U12725 (N_12725,N_6288,N_7718);
and U12726 (N_12726,N_9935,N_8896);
nand U12727 (N_12727,N_9146,N_9859);
and U12728 (N_12728,N_8165,N_9929);
nand U12729 (N_12729,N_8757,N_8606);
nand U12730 (N_12730,N_5070,N_8670);
nand U12731 (N_12731,N_6524,N_7946);
xnor U12732 (N_12732,N_6583,N_7755);
or U12733 (N_12733,N_8455,N_8129);
xor U12734 (N_12734,N_8571,N_5964);
xnor U12735 (N_12735,N_8135,N_9116);
nor U12736 (N_12736,N_6086,N_7452);
xnor U12737 (N_12737,N_8939,N_7031);
xnor U12738 (N_12738,N_9962,N_8929);
or U12739 (N_12739,N_7642,N_5000);
xnor U12740 (N_12740,N_8318,N_5186);
xnor U12741 (N_12741,N_5061,N_6874);
xnor U12742 (N_12742,N_9557,N_8639);
and U12743 (N_12743,N_9765,N_7325);
nand U12744 (N_12744,N_6272,N_6710);
nor U12745 (N_12745,N_6265,N_8413);
nand U12746 (N_12746,N_9464,N_8012);
xor U12747 (N_12747,N_7144,N_7275);
xor U12748 (N_12748,N_8491,N_8253);
xnor U12749 (N_12749,N_8669,N_8956);
xor U12750 (N_12750,N_6291,N_9038);
xnor U12751 (N_12751,N_9483,N_6110);
xnor U12752 (N_12752,N_8730,N_9975);
and U12753 (N_12753,N_7753,N_7032);
or U12754 (N_12754,N_7315,N_7178);
or U12755 (N_12755,N_9751,N_6143);
nor U12756 (N_12756,N_6886,N_7771);
nor U12757 (N_12757,N_6561,N_6821);
nand U12758 (N_12758,N_5193,N_7299);
or U12759 (N_12759,N_6230,N_9690);
nand U12760 (N_12760,N_9087,N_5974);
or U12761 (N_12761,N_7682,N_8273);
nand U12762 (N_12762,N_8897,N_6922);
xor U12763 (N_12763,N_9737,N_7956);
nand U12764 (N_12764,N_5098,N_8243);
and U12765 (N_12765,N_6791,N_6064);
and U12766 (N_12766,N_7836,N_6811);
nor U12767 (N_12767,N_7404,N_9293);
or U12768 (N_12768,N_7256,N_6251);
nand U12769 (N_12769,N_6136,N_8692);
xnor U12770 (N_12770,N_7305,N_9136);
xnor U12771 (N_12771,N_6457,N_8245);
and U12772 (N_12772,N_9573,N_9966);
or U12773 (N_12773,N_8123,N_7959);
nand U12774 (N_12774,N_8870,N_7756);
nand U12775 (N_12775,N_8813,N_7199);
nor U12776 (N_12776,N_9101,N_7386);
or U12777 (N_12777,N_8512,N_8959);
and U12778 (N_12778,N_6147,N_6143);
nand U12779 (N_12779,N_5529,N_9571);
nand U12780 (N_12780,N_6519,N_7761);
or U12781 (N_12781,N_5660,N_9272);
nand U12782 (N_12782,N_9507,N_5433);
xnor U12783 (N_12783,N_8300,N_6606);
and U12784 (N_12784,N_7267,N_5449);
nor U12785 (N_12785,N_6256,N_6021);
nand U12786 (N_12786,N_7023,N_9621);
or U12787 (N_12787,N_9827,N_8898);
and U12788 (N_12788,N_5105,N_8395);
xor U12789 (N_12789,N_9705,N_9756);
nor U12790 (N_12790,N_5178,N_7416);
nand U12791 (N_12791,N_8386,N_7808);
xnor U12792 (N_12792,N_5925,N_7081);
xor U12793 (N_12793,N_9784,N_7904);
xor U12794 (N_12794,N_7661,N_5964);
nand U12795 (N_12795,N_5827,N_6339);
xnor U12796 (N_12796,N_8069,N_7875);
or U12797 (N_12797,N_5113,N_9250);
and U12798 (N_12798,N_6799,N_6407);
xor U12799 (N_12799,N_7353,N_6435);
nand U12800 (N_12800,N_8621,N_8794);
nand U12801 (N_12801,N_8968,N_5758);
nor U12802 (N_12802,N_7232,N_7673);
xnor U12803 (N_12803,N_5963,N_8507);
or U12804 (N_12804,N_5851,N_8670);
nand U12805 (N_12805,N_6930,N_6487);
or U12806 (N_12806,N_5067,N_6519);
nor U12807 (N_12807,N_6831,N_7771);
nor U12808 (N_12808,N_9112,N_7487);
xor U12809 (N_12809,N_9574,N_7575);
xnor U12810 (N_12810,N_7151,N_5667);
or U12811 (N_12811,N_7746,N_9195);
and U12812 (N_12812,N_5106,N_6431);
nor U12813 (N_12813,N_7466,N_7011);
nand U12814 (N_12814,N_7723,N_6516);
or U12815 (N_12815,N_9336,N_7532);
nor U12816 (N_12816,N_6238,N_5606);
xnor U12817 (N_12817,N_7376,N_9438);
xor U12818 (N_12818,N_9376,N_6424);
xor U12819 (N_12819,N_7337,N_8111);
or U12820 (N_12820,N_8824,N_9150);
and U12821 (N_12821,N_5897,N_5646);
xnor U12822 (N_12822,N_8555,N_5675);
or U12823 (N_12823,N_5333,N_9873);
xor U12824 (N_12824,N_9204,N_9230);
or U12825 (N_12825,N_8475,N_9804);
xor U12826 (N_12826,N_5330,N_9179);
nor U12827 (N_12827,N_9643,N_9227);
nor U12828 (N_12828,N_8058,N_7262);
nand U12829 (N_12829,N_8214,N_8856);
or U12830 (N_12830,N_6598,N_5098);
and U12831 (N_12831,N_6836,N_6114);
nand U12832 (N_12832,N_5947,N_6021);
xnor U12833 (N_12833,N_7099,N_9945);
nand U12834 (N_12834,N_5581,N_7019);
nand U12835 (N_12835,N_7495,N_9434);
nand U12836 (N_12836,N_7750,N_5141);
nand U12837 (N_12837,N_5118,N_7070);
nand U12838 (N_12838,N_9255,N_8339);
or U12839 (N_12839,N_8070,N_5045);
xnor U12840 (N_12840,N_9048,N_6485);
and U12841 (N_12841,N_5789,N_6364);
xor U12842 (N_12842,N_9308,N_6781);
or U12843 (N_12843,N_8605,N_9733);
nor U12844 (N_12844,N_5674,N_8557);
nand U12845 (N_12845,N_7914,N_7588);
xor U12846 (N_12846,N_9058,N_9878);
nor U12847 (N_12847,N_9516,N_5208);
nand U12848 (N_12848,N_9290,N_9983);
and U12849 (N_12849,N_6796,N_6167);
and U12850 (N_12850,N_7319,N_6418);
and U12851 (N_12851,N_6988,N_6422);
and U12852 (N_12852,N_9884,N_5979);
xnor U12853 (N_12853,N_9871,N_7886);
nand U12854 (N_12854,N_8547,N_7701);
and U12855 (N_12855,N_9543,N_6900);
xor U12856 (N_12856,N_7555,N_5482);
and U12857 (N_12857,N_7371,N_6425);
and U12858 (N_12858,N_6082,N_6250);
or U12859 (N_12859,N_5714,N_6091);
and U12860 (N_12860,N_8712,N_8476);
nand U12861 (N_12861,N_5800,N_6026);
or U12862 (N_12862,N_5878,N_6975);
and U12863 (N_12863,N_9102,N_6368);
nor U12864 (N_12864,N_8426,N_6179);
nor U12865 (N_12865,N_6902,N_6310);
or U12866 (N_12866,N_9527,N_7287);
or U12867 (N_12867,N_8041,N_5062);
and U12868 (N_12868,N_9798,N_8458);
or U12869 (N_12869,N_9186,N_5323);
nor U12870 (N_12870,N_6299,N_9349);
or U12871 (N_12871,N_6646,N_9317);
xor U12872 (N_12872,N_7506,N_9840);
xor U12873 (N_12873,N_7486,N_9299);
nor U12874 (N_12874,N_6805,N_6747);
xor U12875 (N_12875,N_7567,N_6169);
or U12876 (N_12876,N_6501,N_8539);
nor U12877 (N_12877,N_8746,N_7785);
xor U12878 (N_12878,N_7153,N_8397);
and U12879 (N_12879,N_8980,N_5314);
and U12880 (N_12880,N_8874,N_7972);
or U12881 (N_12881,N_6754,N_8756);
xor U12882 (N_12882,N_5626,N_6562);
and U12883 (N_12883,N_5173,N_7004);
or U12884 (N_12884,N_5624,N_7770);
or U12885 (N_12885,N_6136,N_8163);
and U12886 (N_12886,N_5029,N_5372);
or U12887 (N_12887,N_7259,N_8857);
nand U12888 (N_12888,N_7367,N_8151);
nor U12889 (N_12889,N_7338,N_9843);
nand U12890 (N_12890,N_6390,N_6771);
xnor U12891 (N_12891,N_8677,N_8443);
nor U12892 (N_12892,N_5488,N_7005);
and U12893 (N_12893,N_6071,N_8199);
or U12894 (N_12894,N_8762,N_6333);
and U12895 (N_12895,N_5507,N_6900);
nor U12896 (N_12896,N_8653,N_5281);
or U12897 (N_12897,N_8585,N_5976);
or U12898 (N_12898,N_7373,N_6842);
and U12899 (N_12899,N_7631,N_6794);
and U12900 (N_12900,N_7570,N_8162);
and U12901 (N_12901,N_7516,N_8640);
xor U12902 (N_12902,N_5018,N_5734);
and U12903 (N_12903,N_9184,N_9022);
xnor U12904 (N_12904,N_6923,N_7508);
nand U12905 (N_12905,N_8681,N_7809);
and U12906 (N_12906,N_9427,N_5227);
and U12907 (N_12907,N_9573,N_7250);
nand U12908 (N_12908,N_8054,N_9925);
nor U12909 (N_12909,N_7392,N_5289);
xor U12910 (N_12910,N_7817,N_7653);
xor U12911 (N_12911,N_7239,N_9005);
nand U12912 (N_12912,N_7405,N_6084);
or U12913 (N_12913,N_8984,N_5064);
xor U12914 (N_12914,N_6666,N_8636);
nand U12915 (N_12915,N_6814,N_9815);
xnor U12916 (N_12916,N_9671,N_5709);
or U12917 (N_12917,N_7044,N_6622);
xor U12918 (N_12918,N_7236,N_5674);
and U12919 (N_12919,N_7749,N_8952);
nor U12920 (N_12920,N_7548,N_9684);
nand U12921 (N_12921,N_5158,N_7366);
xnor U12922 (N_12922,N_7578,N_6457);
and U12923 (N_12923,N_5028,N_8991);
and U12924 (N_12924,N_6137,N_8863);
or U12925 (N_12925,N_5782,N_6537);
xor U12926 (N_12926,N_5166,N_5818);
nand U12927 (N_12927,N_6089,N_9070);
nand U12928 (N_12928,N_9644,N_6867);
or U12929 (N_12929,N_6912,N_9498);
nor U12930 (N_12930,N_8886,N_8477);
xor U12931 (N_12931,N_8671,N_5062);
nor U12932 (N_12932,N_6468,N_8521);
and U12933 (N_12933,N_7834,N_5882);
xor U12934 (N_12934,N_5942,N_5569);
and U12935 (N_12935,N_8029,N_9040);
xor U12936 (N_12936,N_8297,N_6657);
and U12937 (N_12937,N_8590,N_5949);
nand U12938 (N_12938,N_6928,N_8708);
or U12939 (N_12939,N_6493,N_6092);
and U12940 (N_12940,N_5178,N_8602);
or U12941 (N_12941,N_8621,N_9352);
and U12942 (N_12942,N_6956,N_9357);
nor U12943 (N_12943,N_7564,N_5862);
xor U12944 (N_12944,N_7390,N_8870);
xnor U12945 (N_12945,N_5889,N_6656);
xor U12946 (N_12946,N_5641,N_9994);
or U12947 (N_12947,N_7315,N_7397);
xor U12948 (N_12948,N_9519,N_9163);
nor U12949 (N_12949,N_8136,N_5429);
or U12950 (N_12950,N_9335,N_6610);
nand U12951 (N_12951,N_5885,N_8178);
or U12952 (N_12952,N_7509,N_7996);
and U12953 (N_12953,N_5768,N_8664);
xor U12954 (N_12954,N_6329,N_5120);
xor U12955 (N_12955,N_6298,N_8740);
nand U12956 (N_12956,N_6009,N_6086);
nand U12957 (N_12957,N_9498,N_5953);
xor U12958 (N_12958,N_7325,N_7582);
and U12959 (N_12959,N_9274,N_8153);
xor U12960 (N_12960,N_8600,N_7522);
nand U12961 (N_12961,N_7649,N_9291);
nand U12962 (N_12962,N_8441,N_8599);
xor U12963 (N_12963,N_5361,N_9551);
and U12964 (N_12964,N_9230,N_8911);
and U12965 (N_12965,N_9897,N_5285);
and U12966 (N_12966,N_7526,N_7098);
or U12967 (N_12967,N_5304,N_9435);
or U12968 (N_12968,N_6197,N_6271);
or U12969 (N_12969,N_7469,N_9725);
xnor U12970 (N_12970,N_7858,N_7025);
and U12971 (N_12971,N_9895,N_5809);
or U12972 (N_12972,N_6339,N_7722);
xnor U12973 (N_12973,N_5990,N_8455);
nor U12974 (N_12974,N_5482,N_9706);
nor U12975 (N_12975,N_8476,N_5593);
xor U12976 (N_12976,N_9292,N_9437);
xor U12977 (N_12977,N_5279,N_5045);
or U12978 (N_12978,N_5659,N_8967);
nor U12979 (N_12979,N_9089,N_7457);
nand U12980 (N_12980,N_7512,N_9438);
xor U12981 (N_12981,N_7292,N_9179);
nand U12982 (N_12982,N_7349,N_9231);
nor U12983 (N_12983,N_8451,N_9885);
and U12984 (N_12984,N_6440,N_5172);
nor U12985 (N_12985,N_9003,N_9417);
or U12986 (N_12986,N_7323,N_8745);
or U12987 (N_12987,N_6582,N_5454);
nor U12988 (N_12988,N_9900,N_8317);
xor U12989 (N_12989,N_6220,N_9430);
nand U12990 (N_12990,N_7049,N_7236);
or U12991 (N_12991,N_7518,N_5791);
xor U12992 (N_12992,N_8591,N_8081);
or U12993 (N_12993,N_9464,N_8473);
nor U12994 (N_12994,N_8798,N_8827);
nor U12995 (N_12995,N_5116,N_5158);
xor U12996 (N_12996,N_6046,N_8928);
or U12997 (N_12997,N_9353,N_6973);
xor U12998 (N_12998,N_9529,N_5546);
or U12999 (N_12999,N_5676,N_6628);
nor U13000 (N_13000,N_5176,N_6094);
xor U13001 (N_13001,N_7969,N_7184);
nand U13002 (N_13002,N_6425,N_7193);
or U13003 (N_13003,N_8312,N_6039);
nand U13004 (N_13004,N_8442,N_7212);
nand U13005 (N_13005,N_7795,N_7239);
and U13006 (N_13006,N_8528,N_7721);
and U13007 (N_13007,N_7994,N_9084);
and U13008 (N_13008,N_9440,N_6046);
or U13009 (N_13009,N_5761,N_5921);
nand U13010 (N_13010,N_7872,N_5360);
xor U13011 (N_13011,N_8421,N_9285);
and U13012 (N_13012,N_9233,N_5529);
or U13013 (N_13013,N_9101,N_8503);
or U13014 (N_13014,N_9419,N_7023);
nand U13015 (N_13015,N_7738,N_6411);
nand U13016 (N_13016,N_5490,N_8052);
nand U13017 (N_13017,N_8127,N_6997);
or U13018 (N_13018,N_8916,N_8737);
nand U13019 (N_13019,N_6552,N_7060);
nor U13020 (N_13020,N_5325,N_9102);
nor U13021 (N_13021,N_8155,N_6763);
nor U13022 (N_13022,N_9223,N_7675);
xor U13023 (N_13023,N_9235,N_8785);
nand U13024 (N_13024,N_8399,N_6134);
nand U13025 (N_13025,N_6557,N_9203);
or U13026 (N_13026,N_9232,N_5137);
and U13027 (N_13027,N_6651,N_8862);
or U13028 (N_13028,N_9472,N_7710);
or U13029 (N_13029,N_8038,N_6071);
nor U13030 (N_13030,N_7032,N_5750);
or U13031 (N_13031,N_5910,N_8546);
xnor U13032 (N_13032,N_6945,N_8638);
xnor U13033 (N_13033,N_7380,N_6925);
and U13034 (N_13034,N_9660,N_6179);
and U13035 (N_13035,N_5313,N_8328);
xor U13036 (N_13036,N_6838,N_8244);
and U13037 (N_13037,N_7959,N_9287);
nor U13038 (N_13038,N_6867,N_6801);
or U13039 (N_13039,N_8305,N_6864);
nor U13040 (N_13040,N_7918,N_6396);
xnor U13041 (N_13041,N_9755,N_8110);
xnor U13042 (N_13042,N_7959,N_8868);
and U13043 (N_13043,N_8251,N_8512);
or U13044 (N_13044,N_7895,N_9904);
xnor U13045 (N_13045,N_6580,N_8541);
or U13046 (N_13046,N_5658,N_7632);
or U13047 (N_13047,N_7245,N_6886);
nand U13048 (N_13048,N_6043,N_6613);
xor U13049 (N_13049,N_9165,N_9086);
nor U13050 (N_13050,N_5295,N_6487);
xor U13051 (N_13051,N_7090,N_5665);
nor U13052 (N_13052,N_6878,N_9177);
nand U13053 (N_13053,N_5142,N_6788);
nand U13054 (N_13054,N_7280,N_5081);
xnor U13055 (N_13055,N_9101,N_7377);
xor U13056 (N_13056,N_6776,N_7968);
xnor U13057 (N_13057,N_5846,N_7125);
and U13058 (N_13058,N_6335,N_5895);
xnor U13059 (N_13059,N_6538,N_9357);
nor U13060 (N_13060,N_8856,N_6064);
and U13061 (N_13061,N_6629,N_6364);
xor U13062 (N_13062,N_6244,N_6972);
nand U13063 (N_13063,N_8449,N_8872);
and U13064 (N_13064,N_9245,N_8489);
nand U13065 (N_13065,N_6489,N_9729);
or U13066 (N_13066,N_5522,N_8249);
xnor U13067 (N_13067,N_9508,N_5900);
nand U13068 (N_13068,N_8779,N_9673);
or U13069 (N_13069,N_8250,N_6638);
xnor U13070 (N_13070,N_7476,N_9308);
nor U13071 (N_13071,N_9635,N_6438);
nor U13072 (N_13072,N_8427,N_5237);
nand U13073 (N_13073,N_5510,N_6157);
and U13074 (N_13074,N_7633,N_6782);
xnor U13075 (N_13075,N_8935,N_9672);
xor U13076 (N_13076,N_7288,N_5634);
nand U13077 (N_13077,N_6911,N_9817);
and U13078 (N_13078,N_7206,N_8849);
xnor U13079 (N_13079,N_6683,N_5009);
nor U13080 (N_13080,N_8188,N_7843);
xnor U13081 (N_13081,N_7055,N_6728);
or U13082 (N_13082,N_6509,N_8954);
and U13083 (N_13083,N_5330,N_9588);
xnor U13084 (N_13084,N_9369,N_9007);
or U13085 (N_13085,N_5524,N_7219);
nand U13086 (N_13086,N_5578,N_6673);
nand U13087 (N_13087,N_8597,N_6134);
or U13088 (N_13088,N_8683,N_9141);
or U13089 (N_13089,N_6004,N_7985);
nand U13090 (N_13090,N_6432,N_6559);
nand U13091 (N_13091,N_7389,N_7878);
nand U13092 (N_13092,N_5756,N_5623);
or U13093 (N_13093,N_5932,N_5444);
nor U13094 (N_13094,N_5562,N_9893);
nand U13095 (N_13095,N_5414,N_5752);
xor U13096 (N_13096,N_7303,N_6300);
nor U13097 (N_13097,N_6632,N_9614);
nand U13098 (N_13098,N_9313,N_8335);
xor U13099 (N_13099,N_8721,N_8655);
nor U13100 (N_13100,N_5066,N_8906);
xor U13101 (N_13101,N_8398,N_6127);
nor U13102 (N_13102,N_8741,N_8536);
nand U13103 (N_13103,N_7011,N_9271);
and U13104 (N_13104,N_9496,N_9835);
or U13105 (N_13105,N_7673,N_9499);
nand U13106 (N_13106,N_8206,N_5496);
nor U13107 (N_13107,N_8994,N_9641);
xor U13108 (N_13108,N_8640,N_8894);
or U13109 (N_13109,N_5044,N_7386);
nand U13110 (N_13110,N_9643,N_8496);
xor U13111 (N_13111,N_6954,N_9711);
or U13112 (N_13112,N_6296,N_5098);
xor U13113 (N_13113,N_8350,N_6486);
nor U13114 (N_13114,N_8326,N_6055);
nor U13115 (N_13115,N_8419,N_7849);
xor U13116 (N_13116,N_7165,N_7347);
and U13117 (N_13117,N_7824,N_9891);
xnor U13118 (N_13118,N_5701,N_5035);
nand U13119 (N_13119,N_7802,N_5184);
nor U13120 (N_13120,N_5074,N_8384);
or U13121 (N_13121,N_9973,N_8375);
or U13122 (N_13122,N_7920,N_8243);
nand U13123 (N_13123,N_9490,N_7715);
or U13124 (N_13124,N_6012,N_8244);
or U13125 (N_13125,N_7566,N_6215);
nand U13126 (N_13126,N_8353,N_8596);
xnor U13127 (N_13127,N_5539,N_8940);
nand U13128 (N_13128,N_8443,N_5484);
nand U13129 (N_13129,N_7176,N_6484);
and U13130 (N_13130,N_7956,N_9286);
nor U13131 (N_13131,N_8428,N_7233);
or U13132 (N_13132,N_9317,N_8013);
xnor U13133 (N_13133,N_7694,N_7998);
and U13134 (N_13134,N_5557,N_6386);
and U13135 (N_13135,N_6577,N_5785);
or U13136 (N_13136,N_8561,N_7289);
xor U13137 (N_13137,N_8765,N_6478);
xor U13138 (N_13138,N_6067,N_5247);
nand U13139 (N_13139,N_5704,N_6633);
and U13140 (N_13140,N_5711,N_6755);
and U13141 (N_13141,N_5288,N_8622);
and U13142 (N_13142,N_5542,N_6418);
or U13143 (N_13143,N_8390,N_7312);
or U13144 (N_13144,N_7073,N_8480);
or U13145 (N_13145,N_7741,N_6341);
nor U13146 (N_13146,N_9519,N_7365);
or U13147 (N_13147,N_6026,N_7257);
or U13148 (N_13148,N_9279,N_8889);
nor U13149 (N_13149,N_9136,N_8640);
nor U13150 (N_13150,N_7947,N_8348);
nor U13151 (N_13151,N_6659,N_9739);
or U13152 (N_13152,N_9580,N_5742);
nor U13153 (N_13153,N_5531,N_6732);
nand U13154 (N_13154,N_6055,N_7825);
or U13155 (N_13155,N_8791,N_8263);
or U13156 (N_13156,N_9765,N_9129);
and U13157 (N_13157,N_7840,N_8159);
and U13158 (N_13158,N_9615,N_9319);
and U13159 (N_13159,N_7482,N_6408);
and U13160 (N_13160,N_5661,N_5507);
nand U13161 (N_13161,N_8135,N_7712);
nor U13162 (N_13162,N_5350,N_7745);
and U13163 (N_13163,N_6132,N_5357);
xnor U13164 (N_13164,N_7982,N_8620);
and U13165 (N_13165,N_7720,N_6608);
nand U13166 (N_13166,N_9994,N_6595);
nand U13167 (N_13167,N_8244,N_5911);
or U13168 (N_13168,N_6157,N_9877);
xor U13169 (N_13169,N_5170,N_9299);
or U13170 (N_13170,N_7719,N_5673);
nand U13171 (N_13171,N_7029,N_9733);
or U13172 (N_13172,N_9701,N_8380);
xor U13173 (N_13173,N_8001,N_9383);
and U13174 (N_13174,N_6546,N_7784);
and U13175 (N_13175,N_5682,N_7872);
and U13176 (N_13176,N_8347,N_8613);
and U13177 (N_13177,N_5114,N_8431);
nor U13178 (N_13178,N_6957,N_8254);
or U13179 (N_13179,N_7635,N_7604);
or U13180 (N_13180,N_6397,N_9861);
nor U13181 (N_13181,N_8254,N_9716);
or U13182 (N_13182,N_9898,N_5439);
and U13183 (N_13183,N_9606,N_5184);
and U13184 (N_13184,N_5822,N_8991);
and U13185 (N_13185,N_8780,N_5429);
nand U13186 (N_13186,N_7437,N_7585);
or U13187 (N_13187,N_8607,N_6221);
or U13188 (N_13188,N_6127,N_5008);
xor U13189 (N_13189,N_7528,N_8611);
xor U13190 (N_13190,N_9310,N_5510);
and U13191 (N_13191,N_5475,N_6741);
xnor U13192 (N_13192,N_8784,N_6225);
xor U13193 (N_13193,N_5042,N_7423);
xnor U13194 (N_13194,N_8967,N_9923);
nor U13195 (N_13195,N_8016,N_8921);
and U13196 (N_13196,N_7411,N_7326);
xor U13197 (N_13197,N_7755,N_8139);
nand U13198 (N_13198,N_8268,N_9677);
and U13199 (N_13199,N_7273,N_7096);
or U13200 (N_13200,N_6568,N_8912);
xnor U13201 (N_13201,N_9478,N_7510);
or U13202 (N_13202,N_7017,N_8338);
nor U13203 (N_13203,N_7495,N_5774);
or U13204 (N_13204,N_9835,N_5540);
or U13205 (N_13205,N_6719,N_6119);
nand U13206 (N_13206,N_6179,N_6918);
nand U13207 (N_13207,N_6236,N_5132);
and U13208 (N_13208,N_9543,N_7477);
and U13209 (N_13209,N_5185,N_5580);
nand U13210 (N_13210,N_5033,N_6585);
nand U13211 (N_13211,N_8305,N_7317);
nor U13212 (N_13212,N_7869,N_7266);
nand U13213 (N_13213,N_7687,N_6220);
nor U13214 (N_13214,N_9247,N_6994);
nand U13215 (N_13215,N_8972,N_6936);
xnor U13216 (N_13216,N_7519,N_9850);
and U13217 (N_13217,N_9898,N_7246);
or U13218 (N_13218,N_6135,N_5883);
xnor U13219 (N_13219,N_5608,N_9028);
xnor U13220 (N_13220,N_6845,N_8543);
xnor U13221 (N_13221,N_7250,N_5973);
nand U13222 (N_13222,N_9558,N_5738);
nand U13223 (N_13223,N_6955,N_5449);
or U13224 (N_13224,N_8180,N_7045);
nand U13225 (N_13225,N_7652,N_7820);
nand U13226 (N_13226,N_7451,N_9371);
nand U13227 (N_13227,N_6230,N_8795);
nand U13228 (N_13228,N_6157,N_5652);
or U13229 (N_13229,N_5173,N_6561);
xnor U13230 (N_13230,N_6709,N_9016);
xnor U13231 (N_13231,N_5981,N_7679);
nor U13232 (N_13232,N_6058,N_6457);
nor U13233 (N_13233,N_6633,N_8335);
nor U13234 (N_13234,N_9515,N_8493);
and U13235 (N_13235,N_8663,N_6240);
and U13236 (N_13236,N_7036,N_6871);
or U13237 (N_13237,N_8770,N_9653);
nand U13238 (N_13238,N_5348,N_9420);
xnor U13239 (N_13239,N_7058,N_5471);
nand U13240 (N_13240,N_5663,N_7945);
xor U13241 (N_13241,N_7106,N_5959);
xor U13242 (N_13242,N_5703,N_7962);
or U13243 (N_13243,N_6400,N_9713);
xnor U13244 (N_13244,N_6517,N_9996);
nand U13245 (N_13245,N_9820,N_6108);
xnor U13246 (N_13246,N_5618,N_7155);
nor U13247 (N_13247,N_8138,N_5650);
and U13248 (N_13248,N_6940,N_6867);
or U13249 (N_13249,N_7306,N_5151);
nor U13250 (N_13250,N_8597,N_5826);
nand U13251 (N_13251,N_5229,N_5445);
nor U13252 (N_13252,N_8752,N_9986);
nor U13253 (N_13253,N_6173,N_9397);
nand U13254 (N_13254,N_9694,N_7698);
nor U13255 (N_13255,N_8601,N_5829);
nand U13256 (N_13256,N_9099,N_6281);
or U13257 (N_13257,N_8016,N_8763);
and U13258 (N_13258,N_8732,N_7361);
nand U13259 (N_13259,N_6128,N_8873);
or U13260 (N_13260,N_8135,N_7978);
nor U13261 (N_13261,N_9365,N_7769);
xnor U13262 (N_13262,N_7045,N_9637);
and U13263 (N_13263,N_5265,N_6325);
or U13264 (N_13264,N_9359,N_9420);
xor U13265 (N_13265,N_6055,N_8618);
nor U13266 (N_13266,N_8654,N_9850);
or U13267 (N_13267,N_9471,N_7243);
xor U13268 (N_13268,N_9978,N_7202);
xor U13269 (N_13269,N_7471,N_5590);
and U13270 (N_13270,N_7026,N_6928);
and U13271 (N_13271,N_5203,N_6492);
nor U13272 (N_13272,N_9691,N_6662);
or U13273 (N_13273,N_8903,N_9594);
or U13274 (N_13274,N_8567,N_6602);
xnor U13275 (N_13275,N_7972,N_6411);
nor U13276 (N_13276,N_5156,N_6786);
or U13277 (N_13277,N_7472,N_8644);
nand U13278 (N_13278,N_6763,N_7744);
nand U13279 (N_13279,N_7103,N_5671);
or U13280 (N_13280,N_7938,N_9359);
or U13281 (N_13281,N_7444,N_5449);
nor U13282 (N_13282,N_7518,N_5646);
and U13283 (N_13283,N_6333,N_6407);
or U13284 (N_13284,N_6978,N_7471);
nor U13285 (N_13285,N_6234,N_8679);
and U13286 (N_13286,N_6342,N_7087);
or U13287 (N_13287,N_8983,N_6669);
nand U13288 (N_13288,N_8653,N_6535);
nand U13289 (N_13289,N_8468,N_9950);
nor U13290 (N_13290,N_5542,N_5842);
or U13291 (N_13291,N_6130,N_6650);
xnor U13292 (N_13292,N_5887,N_6746);
or U13293 (N_13293,N_9903,N_8031);
or U13294 (N_13294,N_7361,N_7235);
or U13295 (N_13295,N_7066,N_9301);
xnor U13296 (N_13296,N_5278,N_7932);
nand U13297 (N_13297,N_8808,N_9542);
xor U13298 (N_13298,N_5644,N_5397);
nand U13299 (N_13299,N_5834,N_8125);
xnor U13300 (N_13300,N_9389,N_7842);
nand U13301 (N_13301,N_8316,N_5133);
xor U13302 (N_13302,N_7612,N_6617);
xor U13303 (N_13303,N_6626,N_9826);
nor U13304 (N_13304,N_7482,N_8468);
xnor U13305 (N_13305,N_6191,N_9783);
and U13306 (N_13306,N_9911,N_5742);
xor U13307 (N_13307,N_6648,N_9412);
nor U13308 (N_13308,N_7032,N_9751);
and U13309 (N_13309,N_6784,N_7480);
nor U13310 (N_13310,N_7599,N_8594);
nor U13311 (N_13311,N_7632,N_5712);
or U13312 (N_13312,N_5000,N_6755);
and U13313 (N_13313,N_5864,N_5002);
and U13314 (N_13314,N_8724,N_9642);
xnor U13315 (N_13315,N_5474,N_7325);
nand U13316 (N_13316,N_6286,N_9069);
nor U13317 (N_13317,N_6623,N_9839);
nor U13318 (N_13318,N_6273,N_9354);
xnor U13319 (N_13319,N_9592,N_6944);
nand U13320 (N_13320,N_6273,N_8405);
or U13321 (N_13321,N_5944,N_9577);
nand U13322 (N_13322,N_5546,N_6260);
or U13323 (N_13323,N_7923,N_9975);
nand U13324 (N_13324,N_8042,N_7091);
or U13325 (N_13325,N_6378,N_8517);
xnor U13326 (N_13326,N_9455,N_6973);
nor U13327 (N_13327,N_6771,N_5764);
xnor U13328 (N_13328,N_6497,N_5330);
and U13329 (N_13329,N_9122,N_9993);
nand U13330 (N_13330,N_7618,N_8606);
and U13331 (N_13331,N_6024,N_8742);
and U13332 (N_13332,N_6747,N_6849);
nor U13333 (N_13333,N_6441,N_6798);
nor U13334 (N_13334,N_9650,N_5323);
xor U13335 (N_13335,N_9595,N_9426);
nor U13336 (N_13336,N_6247,N_6044);
xor U13337 (N_13337,N_5185,N_6899);
nand U13338 (N_13338,N_7738,N_6755);
and U13339 (N_13339,N_5282,N_6402);
and U13340 (N_13340,N_7158,N_7177);
nor U13341 (N_13341,N_9479,N_6955);
xor U13342 (N_13342,N_7258,N_5502);
and U13343 (N_13343,N_8384,N_7744);
nor U13344 (N_13344,N_7842,N_6231);
nor U13345 (N_13345,N_5993,N_5862);
nand U13346 (N_13346,N_9280,N_6406);
nor U13347 (N_13347,N_6095,N_6032);
nor U13348 (N_13348,N_7033,N_5504);
nand U13349 (N_13349,N_5392,N_9343);
nand U13350 (N_13350,N_6130,N_8654);
or U13351 (N_13351,N_8626,N_5887);
nor U13352 (N_13352,N_9664,N_6834);
nand U13353 (N_13353,N_5009,N_6393);
or U13354 (N_13354,N_5683,N_6676);
nor U13355 (N_13355,N_7387,N_5447);
xnor U13356 (N_13356,N_5765,N_9418);
nand U13357 (N_13357,N_7416,N_6252);
nand U13358 (N_13358,N_9898,N_7728);
or U13359 (N_13359,N_9637,N_8653);
or U13360 (N_13360,N_8421,N_7865);
or U13361 (N_13361,N_9183,N_7889);
and U13362 (N_13362,N_8494,N_8647);
nor U13363 (N_13363,N_5392,N_5594);
nor U13364 (N_13364,N_9997,N_7586);
nand U13365 (N_13365,N_5238,N_8027);
or U13366 (N_13366,N_6035,N_9080);
xnor U13367 (N_13367,N_9251,N_5028);
and U13368 (N_13368,N_5874,N_6427);
and U13369 (N_13369,N_5493,N_7637);
nand U13370 (N_13370,N_6374,N_7612);
and U13371 (N_13371,N_8624,N_9815);
or U13372 (N_13372,N_6309,N_7582);
or U13373 (N_13373,N_8239,N_5174);
nor U13374 (N_13374,N_8925,N_9197);
or U13375 (N_13375,N_5253,N_7728);
or U13376 (N_13376,N_7726,N_6506);
or U13377 (N_13377,N_7490,N_9628);
and U13378 (N_13378,N_6027,N_8799);
nor U13379 (N_13379,N_8361,N_6793);
nand U13380 (N_13380,N_8393,N_7591);
nor U13381 (N_13381,N_5557,N_8757);
nor U13382 (N_13382,N_5312,N_7165);
xor U13383 (N_13383,N_8337,N_9992);
and U13384 (N_13384,N_6301,N_9307);
nand U13385 (N_13385,N_5989,N_5247);
and U13386 (N_13386,N_7736,N_7058);
nor U13387 (N_13387,N_8379,N_8299);
nor U13388 (N_13388,N_5446,N_8596);
xor U13389 (N_13389,N_8784,N_7389);
and U13390 (N_13390,N_7933,N_8620);
and U13391 (N_13391,N_7239,N_9271);
and U13392 (N_13392,N_8113,N_5515);
xor U13393 (N_13393,N_9208,N_6226);
or U13394 (N_13394,N_8974,N_6536);
or U13395 (N_13395,N_7670,N_9368);
and U13396 (N_13396,N_7597,N_6488);
nand U13397 (N_13397,N_5044,N_5463);
xor U13398 (N_13398,N_6861,N_8864);
xnor U13399 (N_13399,N_9473,N_7590);
xor U13400 (N_13400,N_9075,N_5631);
or U13401 (N_13401,N_8015,N_6482);
nand U13402 (N_13402,N_8023,N_8757);
xor U13403 (N_13403,N_8732,N_8794);
xnor U13404 (N_13404,N_8189,N_6362);
nand U13405 (N_13405,N_8668,N_7804);
nor U13406 (N_13406,N_8816,N_5508);
nand U13407 (N_13407,N_7638,N_6789);
and U13408 (N_13408,N_8439,N_8960);
and U13409 (N_13409,N_8089,N_8420);
xnor U13410 (N_13410,N_9370,N_8794);
or U13411 (N_13411,N_9505,N_8279);
and U13412 (N_13412,N_6684,N_5372);
and U13413 (N_13413,N_9944,N_8555);
or U13414 (N_13414,N_6988,N_7848);
or U13415 (N_13415,N_6942,N_9474);
nor U13416 (N_13416,N_8954,N_5824);
nor U13417 (N_13417,N_8012,N_7939);
nand U13418 (N_13418,N_5795,N_7682);
and U13419 (N_13419,N_9300,N_8986);
or U13420 (N_13420,N_8270,N_9296);
nand U13421 (N_13421,N_6603,N_5481);
nor U13422 (N_13422,N_9312,N_9191);
or U13423 (N_13423,N_7195,N_5506);
xnor U13424 (N_13424,N_6230,N_7921);
or U13425 (N_13425,N_8403,N_6645);
nor U13426 (N_13426,N_8071,N_8663);
xor U13427 (N_13427,N_8465,N_7846);
xor U13428 (N_13428,N_7771,N_9026);
nor U13429 (N_13429,N_6454,N_8842);
and U13430 (N_13430,N_9452,N_8222);
or U13431 (N_13431,N_5418,N_8623);
nor U13432 (N_13432,N_8221,N_6114);
nand U13433 (N_13433,N_9147,N_9610);
nand U13434 (N_13434,N_5514,N_8290);
nand U13435 (N_13435,N_8849,N_7409);
or U13436 (N_13436,N_5768,N_5624);
nand U13437 (N_13437,N_5929,N_6661);
nand U13438 (N_13438,N_9415,N_6849);
nand U13439 (N_13439,N_7514,N_6112);
and U13440 (N_13440,N_7668,N_7909);
nand U13441 (N_13441,N_8449,N_8178);
nand U13442 (N_13442,N_5863,N_8167);
or U13443 (N_13443,N_5713,N_8460);
and U13444 (N_13444,N_8834,N_7378);
xnor U13445 (N_13445,N_8884,N_8734);
or U13446 (N_13446,N_7421,N_9805);
nor U13447 (N_13447,N_7752,N_7119);
nand U13448 (N_13448,N_5616,N_8268);
and U13449 (N_13449,N_7436,N_7545);
xnor U13450 (N_13450,N_5729,N_7103);
or U13451 (N_13451,N_6330,N_9825);
nand U13452 (N_13452,N_7068,N_7603);
and U13453 (N_13453,N_9735,N_9742);
or U13454 (N_13454,N_9589,N_7004);
or U13455 (N_13455,N_8202,N_5938);
nor U13456 (N_13456,N_9326,N_8238);
xnor U13457 (N_13457,N_6790,N_8682);
nor U13458 (N_13458,N_8502,N_6871);
xor U13459 (N_13459,N_7575,N_7794);
and U13460 (N_13460,N_9088,N_6646);
nand U13461 (N_13461,N_9357,N_6178);
or U13462 (N_13462,N_8076,N_9797);
nor U13463 (N_13463,N_9710,N_9049);
xnor U13464 (N_13464,N_9422,N_6691);
or U13465 (N_13465,N_5291,N_5614);
nor U13466 (N_13466,N_6774,N_6679);
xor U13467 (N_13467,N_9133,N_8168);
nor U13468 (N_13468,N_5104,N_8023);
or U13469 (N_13469,N_8386,N_7340);
or U13470 (N_13470,N_9771,N_7193);
xnor U13471 (N_13471,N_7515,N_7815);
and U13472 (N_13472,N_8716,N_6080);
nand U13473 (N_13473,N_7387,N_9734);
nor U13474 (N_13474,N_7260,N_8699);
and U13475 (N_13475,N_9689,N_6381);
nor U13476 (N_13476,N_6087,N_7872);
nand U13477 (N_13477,N_7551,N_7331);
nor U13478 (N_13478,N_5666,N_9809);
xnor U13479 (N_13479,N_8121,N_8672);
and U13480 (N_13480,N_7387,N_5518);
xnor U13481 (N_13481,N_6094,N_9316);
and U13482 (N_13482,N_8155,N_9999);
nor U13483 (N_13483,N_8461,N_5680);
xor U13484 (N_13484,N_5498,N_9597);
or U13485 (N_13485,N_7678,N_6037);
or U13486 (N_13486,N_6693,N_9153);
and U13487 (N_13487,N_7259,N_7798);
and U13488 (N_13488,N_7816,N_8237);
xnor U13489 (N_13489,N_5511,N_6101);
nor U13490 (N_13490,N_6581,N_6091);
and U13491 (N_13491,N_5637,N_7828);
xor U13492 (N_13492,N_5756,N_5843);
nor U13493 (N_13493,N_6539,N_5499);
xnor U13494 (N_13494,N_5847,N_8460);
or U13495 (N_13495,N_7807,N_7941);
nor U13496 (N_13496,N_7161,N_9062);
nor U13497 (N_13497,N_9383,N_7679);
or U13498 (N_13498,N_6003,N_9071);
xor U13499 (N_13499,N_7627,N_6805);
nor U13500 (N_13500,N_8360,N_8370);
nor U13501 (N_13501,N_6422,N_7479);
or U13502 (N_13502,N_9212,N_8326);
or U13503 (N_13503,N_7680,N_6287);
and U13504 (N_13504,N_9631,N_5462);
nand U13505 (N_13505,N_6944,N_5380);
nor U13506 (N_13506,N_9547,N_8551);
nand U13507 (N_13507,N_7666,N_8335);
or U13508 (N_13508,N_7524,N_6455);
nand U13509 (N_13509,N_7738,N_5127);
or U13510 (N_13510,N_9314,N_6878);
and U13511 (N_13511,N_6059,N_6705);
nor U13512 (N_13512,N_5775,N_7301);
xor U13513 (N_13513,N_8654,N_7214);
xnor U13514 (N_13514,N_8314,N_5170);
nand U13515 (N_13515,N_8592,N_7988);
or U13516 (N_13516,N_7084,N_5287);
xnor U13517 (N_13517,N_5605,N_5211);
nand U13518 (N_13518,N_9281,N_8056);
and U13519 (N_13519,N_6849,N_5256);
xor U13520 (N_13520,N_9879,N_6345);
or U13521 (N_13521,N_7016,N_7497);
or U13522 (N_13522,N_6683,N_8948);
or U13523 (N_13523,N_9875,N_7365);
xor U13524 (N_13524,N_9236,N_5801);
nand U13525 (N_13525,N_5673,N_5205);
and U13526 (N_13526,N_6341,N_7216);
and U13527 (N_13527,N_9814,N_8628);
nor U13528 (N_13528,N_7138,N_9800);
xor U13529 (N_13529,N_5767,N_6344);
xnor U13530 (N_13530,N_7602,N_7499);
nand U13531 (N_13531,N_7114,N_9660);
xor U13532 (N_13532,N_8675,N_7297);
nand U13533 (N_13533,N_7510,N_7784);
xor U13534 (N_13534,N_8362,N_7061);
and U13535 (N_13535,N_9580,N_5291);
nand U13536 (N_13536,N_6730,N_8816);
nand U13537 (N_13537,N_8054,N_9992);
nor U13538 (N_13538,N_9614,N_6047);
xor U13539 (N_13539,N_5129,N_8636);
or U13540 (N_13540,N_5601,N_5318);
xor U13541 (N_13541,N_8345,N_5506);
or U13542 (N_13542,N_8771,N_6411);
nor U13543 (N_13543,N_6411,N_6909);
or U13544 (N_13544,N_8866,N_6983);
and U13545 (N_13545,N_7285,N_9772);
nor U13546 (N_13546,N_9026,N_9574);
nand U13547 (N_13547,N_5702,N_7119);
nand U13548 (N_13548,N_9177,N_9883);
or U13549 (N_13549,N_9698,N_9910);
and U13550 (N_13550,N_9592,N_8670);
nand U13551 (N_13551,N_8841,N_7711);
xor U13552 (N_13552,N_8984,N_7714);
nand U13553 (N_13553,N_7985,N_5633);
xor U13554 (N_13554,N_5089,N_7610);
xor U13555 (N_13555,N_5185,N_9506);
xnor U13556 (N_13556,N_7575,N_9629);
nor U13557 (N_13557,N_8540,N_5655);
nor U13558 (N_13558,N_6987,N_5052);
or U13559 (N_13559,N_6216,N_9767);
and U13560 (N_13560,N_8125,N_8498);
nand U13561 (N_13561,N_9108,N_5023);
xor U13562 (N_13562,N_8797,N_7697);
nor U13563 (N_13563,N_7368,N_9095);
xnor U13564 (N_13564,N_8647,N_8255);
xnor U13565 (N_13565,N_7910,N_9466);
nor U13566 (N_13566,N_5754,N_9507);
nor U13567 (N_13567,N_8814,N_5325);
nor U13568 (N_13568,N_8080,N_7102);
nor U13569 (N_13569,N_5691,N_6191);
and U13570 (N_13570,N_9150,N_8567);
and U13571 (N_13571,N_7127,N_5010);
and U13572 (N_13572,N_7081,N_5349);
nor U13573 (N_13573,N_7485,N_5855);
and U13574 (N_13574,N_9813,N_9212);
nand U13575 (N_13575,N_7205,N_7095);
or U13576 (N_13576,N_6304,N_8081);
xnor U13577 (N_13577,N_7436,N_7358);
or U13578 (N_13578,N_8617,N_7762);
or U13579 (N_13579,N_8611,N_5980);
xnor U13580 (N_13580,N_5612,N_6231);
xor U13581 (N_13581,N_9769,N_9210);
nand U13582 (N_13582,N_7519,N_8043);
nand U13583 (N_13583,N_8411,N_9953);
nor U13584 (N_13584,N_6741,N_8840);
nor U13585 (N_13585,N_8164,N_5554);
and U13586 (N_13586,N_7565,N_8651);
and U13587 (N_13587,N_5026,N_6519);
nor U13588 (N_13588,N_9142,N_6161);
nor U13589 (N_13589,N_5493,N_8706);
or U13590 (N_13590,N_9231,N_9987);
nand U13591 (N_13591,N_6207,N_8280);
nand U13592 (N_13592,N_5675,N_7811);
and U13593 (N_13593,N_8171,N_5583);
nand U13594 (N_13594,N_6212,N_7897);
nand U13595 (N_13595,N_5390,N_7792);
nor U13596 (N_13596,N_6608,N_9310);
xnor U13597 (N_13597,N_5511,N_7114);
or U13598 (N_13598,N_5833,N_5471);
or U13599 (N_13599,N_5735,N_7416);
or U13600 (N_13600,N_8865,N_9830);
and U13601 (N_13601,N_8165,N_9345);
xor U13602 (N_13602,N_5736,N_8479);
or U13603 (N_13603,N_6622,N_6102);
nor U13604 (N_13604,N_7281,N_9752);
nor U13605 (N_13605,N_7948,N_9504);
xnor U13606 (N_13606,N_6270,N_5432);
nor U13607 (N_13607,N_9153,N_6742);
nand U13608 (N_13608,N_5738,N_6135);
or U13609 (N_13609,N_7930,N_6424);
nand U13610 (N_13610,N_7799,N_6093);
nor U13611 (N_13611,N_6647,N_7896);
xnor U13612 (N_13612,N_7502,N_7490);
xor U13613 (N_13613,N_8883,N_8790);
xor U13614 (N_13614,N_7678,N_6067);
or U13615 (N_13615,N_8361,N_6914);
nand U13616 (N_13616,N_9263,N_9515);
and U13617 (N_13617,N_7895,N_7494);
nor U13618 (N_13618,N_9887,N_9000);
and U13619 (N_13619,N_7190,N_8689);
and U13620 (N_13620,N_9294,N_7296);
nor U13621 (N_13621,N_5385,N_5221);
xnor U13622 (N_13622,N_6716,N_6162);
and U13623 (N_13623,N_5666,N_8854);
nand U13624 (N_13624,N_8781,N_9964);
xor U13625 (N_13625,N_9961,N_9564);
and U13626 (N_13626,N_5080,N_5470);
and U13627 (N_13627,N_7544,N_7331);
or U13628 (N_13628,N_9086,N_9109);
nand U13629 (N_13629,N_9307,N_9489);
or U13630 (N_13630,N_7450,N_6832);
xnor U13631 (N_13631,N_5583,N_6095);
or U13632 (N_13632,N_9096,N_7456);
xnor U13633 (N_13633,N_8319,N_6424);
xor U13634 (N_13634,N_8676,N_9131);
nand U13635 (N_13635,N_9748,N_5326);
nor U13636 (N_13636,N_7610,N_8396);
nand U13637 (N_13637,N_7542,N_8908);
xnor U13638 (N_13638,N_5979,N_8761);
xnor U13639 (N_13639,N_6479,N_8786);
nand U13640 (N_13640,N_5397,N_5918);
xnor U13641 (N_13641,N_9327,N_9906);
and U13642 (N_13642,N_5438,N_9799);
nor U13643 (N_13643,N_6377,N_5439);
nor U13644 (N_13644,N_9173,N_5886);
nor U13645 (N_13645,N_9041,N_8482);
xor U13646 (N_13646,N_6591,N_8045);
nor U13647 (N_13647,N_9285,N_6296);
and U13648 (N_13648,N_6274,N_6987);
nand U13649 (N_13649,N_6625,N_7785);
nor U13650 (N_13650,N_9160,N_9413);
nor U13651 (N_13651,N_8036,N_5863);
and U13652 (N_13652,N_8423,N_7445);
xnor U13653 (N_13653,N_9293,N_9725);
nand U13654 (N_13654,N_8620,N_6269);
or U13655 (N_13655,N_6172,N_9033);
and U13656 (N_13656,N_6439,N_8915);
xnor U13657 (N_13657,N_5823,N_9124);
nand U13658 (N_13658,N_6420,N_8333);
and U13659 (N_13659,N_5705,N_8550);
or U13660 (N_13660,N_8145,N_7117);
nand U13661 (N_13661,N_7376,N_8175);
nor U13662 (N_13662,N_6970,N_7466);
or U13663 (N_13663,N_5529,N_6757);
or U13664 (N_13664,N_8643,N_5674);
nor U13665 (N_13665,N_8514,N_8850);
xor U13666 (N_13666,N_7379,N_9441);
and U13667 (N_13667,N_6848,N_9061);
or U13668 (N_13668,N_5731,N_7737);
and U13669 (N_13669,N_6112,N_8021);
xor U13670 (N_13670,N_5983,N_7039);
nor U13671 (N_13671,N_6217,N_8241);
nand U13672 (N_13672,N_5987,N_7046);
nor U13673 (N_13673,N_8992,N_9615);
xor U13674 (N_13674,N_6672,N_6750);
nand U13675 (N_13675,N_8762,N_8871);
xnor U13676 (N_13676,N_6382,N_9993);
xnor U13677 (N_13677,N_8427,N_8568);
xor U13678 (N_13678,N_6483,N_9407);
nor U13679 (N_13679,N_6650,N_7953);
and U13680 (N_13680,N_9054,N_5299);
and U13681 (N_13681,N_8050,N_7583);
xor U13682 (N_13682,N_9541,N_5721);
and U13683 (N_13683,N_9152,N_7989);
nor U13684 (N_13684,N_5165,N_5051);
and U13685 (N_13685,N_5696,N_9100);
or U13686 (N_13686,N_5506,N_8974);
xor U13687 (N_13687,N_6595,N_8965);
and U13688 (N_13688,N_9710,N_9971);
xnor U13689 (N_13689,N_5873,N_6534);
nand U13690 (N_13690,N_7737,N_8873);
or U13691 (N_13691,N_8942,N_5134);
and U13692 (N_13692,N_8171,N_5329);
xnor U13693 (N_13693,N_8800,N_6346);
nor U13694 (N_13694,N_5876,N_8210);
nand U13695 (N_13695,N_9051,N_7441);
nand U13696 (N_13696,N_5091,N_6105);
nand U13697 (N_13697,N_9886,N_7597);
or U13698 (N_13698,N_9223,N_6774);
xnor U13699 (N_13699,N_5421,N_6385);
xor U13700 (N_13700,N_8926,N_9662);
nor U13701 (N_13701,N_7482,N_5513);
or U13702 (N_13702,N_7890,N_5843);
xor U13703 (N_13703,N_8077,N_9009);
or U13704 (N_13704,N_5510,N_5943);
xnor U13705 (N_13705,N_7094,N_8318);
nand U13706 (N_13706,N_9055,N_6025);
nor U13707 (N_13707,N_6615,N_9499);
or U13708 (N_13708,N_6496,N_5087);
nor U13709 (N_13709,N_5044,N_6913);
or U13710 (N_13710,N_9604,N_6689);
nand U13711 (N_13711,N_8989,N_8851);
xor U13712 (N_13712,N_9017,N_8582);
xnor U13713 (N_13713,N_6679,N_5839);
xor U13714 (N_13714,N_9143,N_7666);
nor U13715 (N_13715,N_7720,N_6943);
xnor U13716 (N_13716,N_9402,N_7258);
nor U13717 (N_13717,N_6796,N_9513);
or U13718 (N_13718,N_5399,N_5908);
or U13719 (N_13719,N_7467,N_6256);
and U13720 (N_13720,N_9620,N_5194);
and U13721 (N_13721,N_9988,N_6178);
or U13722 (N_13722,N_6506,N_5114);
or U13723 (N_13723,N_7238,N_7409);
or U13724 (N_13724,N_5474,N_7277);
nand U13725 (N_13725,N_5977,N_8353);
nand U13726 (N_13726,N_9038,N_5793);
xor U13727 (N_13727,N_6301,N_5436);
and U13728 (N_13728,N_5704,N_8676);
or U13729 (N_13729,N_9743,N_9097);
nor U13730 (N_13730,N_7340,N_5877);
or U13731 (N_13731,N_7150,N_9330);
nor U13732 (N_13732,N_6593,N_5798);
nand U13733 (N_13733,N_8802,N_6279);
or U13734 (N_13734,N_9525,N_9217);
nor U13735 (N_13735,N_9254,N_9218);
and U13736 (N_13736,N_8954,N_9766);
nor U13737 (N_13737,N_8885,N_8155);
xor U13738 (N_13738,N_5347,N_9682);
or U13739 (N_13739,N_6160,N_7537);
nor U13740 (N_13740,N_5841,N_7840);
xnor U13741 (N_13741,N_7530,N_5886);
or U13742 (N_13742,N_6866,N_9317);
nor U13743 (N_13743,N_9236,N_7614);
nand U13744 (N_13744,N_5675,N_6073);
nor U13745 (N_13745,N_6551,N_8987);
nand U13746 (N_13746,N_8019,N_7777);
or U13747 (N_13747,N_9905,N_9532);
xnor U13748 (N_13748,N_8880,N_9735);
nor U13749 (N_13749,N_9081,N_7697);
or U13750 (N_13750,N_7808,N_9110);
nand U13751 (N_13751,N_5212,N_9926);
and U13752 (N_13752,N_8076,N_8381);
or U13753 (N_13753,N_6596,N_6018);
or U13754 (N_13754,N_6429,N_5438);
nor U13755 (N_13755,N_6657,N_7838);
xor U13756 (N_13756,N_6382,N_5920);
and U13757 (N_13757,N_5612,N_9304);
xnor U13758 (N_13758,N_5689,N_8900);
or U13759 (N_13759,N_5174,N_9789);
xor U13760 (N_13760,N_9308,N_7082);
or U13761 (N_13761,N_9692,N_6796);
nand U13762 (N_13762,N_6018,N_9511);
and U13763 (N_13763,N_9990,N_8372);
nor U13764 (N_13764,N_6994,N_5259);
or U13765 (N_13765,N_5930,N_5997);
and U13766 (N_13766,N_7781,N_8201);
nor U13767 (N_13767,N_7912,N_9205);
or U13768 (N_13768,N_7686,N_5704);
xnor U13769 (N_13769,N_8344,N_5516);
or U13770 (N_13770,N_8033,N_5887);
nor U13771 (N_13771,N_7370,N_8779);
nand U13772 (N_13772,N_6298,N_6495);
and U13773 (N_13773,N_5798,N_5744);
or U13774 (N_13774,N_8513,N_5627);
and U13775 (N_13775,N_5200,N_5821);
and U13776 (N_13776,N_6025,N_9916);
xor U13777 (N_13777,N_7612,N_8534);
nand U13778 (N_13778,N_6457,N_5435);
nor U13779 (N_13779,N_5399,N_7116);
and U13780 (N_13780,N_6653,N_7780);
xor U13781 (N_13781,N_9851,N_5696);
or U13782 (N_13782,N_8254,N_7120);
nand U13783 (N_13783,N_8382,N_5637);
xor U13784 (N_13784,N_9887,N_8112);
or U13785 (N_13785,N_7999,N_5378);
or U13786 (N_13786,N_5452,N_7276);
xnor U13787 (N_13787,N_7340,N_5774);
nand U13788 (N_13788,N_5659,N_7742);
or U13789 (N_13789,N_6786,N_5508);
or U13790 (N_13790,N_9684,N_8463);
and U13791 (N_13791,N_6784,N_8222);
or U13792 (N_13792,N_5197,N_8936);
and U13793 (N_13793,N_7706,N_5987);
or U13794 (N_13794,N_6325,N_5330);
xnor U13795 (N_13795,N_9998,N_9619);
nand U13796 (N_13796,N_5173,N_7870);
or U13797 (N_13797,N_8374,N_8031);
and U13798 (N_13798,N_9468,N_6118);
xnor U13799 (N_13799,N_5883,N_9810);
nand U13800 (N_13800,N_7619,N_6114);
nand U13801 (N_13801,N_5609,N_7269);
nand U13802 (N_13802,N_6050,N_5213);
nand U13803 (N_13803,N_9486,N_6751);
xnor U13804 (N_13804,N_7655,N_5347);
nand U13805 (N_13805,N_9856,N_5975);
and U13806 (N_13806,N_8582,N_6618);
nor U13807 (N_13807,N_7847,N_9883);
or U13808 (N_13808,N_9850,N_6982);
xnor U13809 (N_13809,N_9198,N_7980);
nand U13810 (N_13810,N_7492,N_7447);
xnor U13811 (N_13811,N_9607,N_8230);
nor U13812 (N_13812,N_5605,N_9736);
nor U13813 (N_13813,N_5851,N_8832);
nand U13814 (N_13814,N_9069,N_6129);
nor U13815 (N_13815,N_8203,N_5539);
and U13816 (N_13816,N_7378,N_6429);
xnor U13817 (N_13817,N_8175,N_8905);
nor U13818 (N_13818,N_6959,N_6565);
nor U13819 (N_13819,N_7402,N_8021);
xor U13820 (N_13820,N_6305,N_8209);
nand U13821 (N_13821,N_5014,N_7112);
nor U13822 (N_13822,N_5464,N_6007);
and U13823 (N_13823,N_6804,N_5091);
nor U13824 (N_13824,N_5570,N_6724);
nand U13825 (N_13825,N_5047,N_5462);
xor U13826 (N_13826,N_8063,N_7175);
and U13827 (N_13827,N_5718,N_8182);
nor U13828 (N_13828,N_5141,N_8519);
or U13829 (N_13829,N_5747,N_5492);
nor U13830 (N_13830,N_9724,N_7182);
nor U13831 (N_13831,N_6713,N_5665);
nor U13832 (N_13832,N_9673,N_5151);
nand U13833 (N_13833,N_7886,N_7929);
or U13834 (N_13834,N_8782,N_8911);
nand U13835 (N_13835,N_9951,N_6579);
or U13836 (N_13836,N_7868,N_6790);
and U13837 (N_13837,N_8169,N_8635);
xnor U13838 (N_13838,N_8401,N_5236);
nor U13839 (N_13839,N_9537,N_6302);
or U13840 (N_13840,N_9442,N_5370);
nor U13841 (N_13841,N_5811,N_7240);
and U13842 (N_13842,N_8221,N_7945);
nor U13843 (N_13843,N_7878,N_6036);
or U13844 (N_13844,N_7864,N_9361);
and U13845 (N_13845,N_6289,N_5716);
nand U13846 (N_13846,N_5586,N_5800);
or U13847 (N_13847,N_8308,N_9174);
nand U13848 (N_13848,N_7819,N_9446);
nand U13849 (N_13849,N_7854,N_8768);
nor U13850 (N_13850,N_8357,N_7803);
xor U13851 (N_13851,N_8823,N_8046);
nand U13852 (N_13852,N_5317,N_9624);
or U13853 (N_13853,N_7886,N_6493);
and U13854 (N_13854,N_7319,N_9813);
xor U13855 (N_13855,N_5732,N_7030);
or U13856 (N_13856,N_5280,N_5120);
nor U13857 (N_13857,N_8538,N_6041);
nand U13858 (N_13858,N_7708,N_8484);
xor U13859 (N_13859,N_5696,N_7066);
nand U13860 (N_13860,N_9150,N_6139);
nand U13861 (N_13861,N_5833,N_5500);
and U13862 (N_13862,N_8886,N_7708);
xnor U13863 (N_13863,N_7316,N_5038);
nand U13864 (N_13864,N_7445,N_8764);
xor U13865 (N_13865,N_5429,N_9309);
and U13866 (N_13866,N_7914,N_7651);
or U13867 (N_13867,N_6514,N_8514);
nor U13868 (N_13868,N_5538,N_7334);
or U13869 (N_13869,N_8107,N_6267);
nand U13870 (N_13870,N_7795,N_9561);
and U13871 (N_13871,N_5952,N_5550);
and U13872 (N_13872,N_5914,N_8064);
xor U13873 (N_13873,N_8369,N_9707);
or U13874 (N_13874,N_5351,N_6700);
and U13875 (N_13875,N_8536,N_8687);
and U13876 (N_13876,N_5795,N_7661);
nand U13877 (N_13877,N_5344,N_9332);
and U13878 (N_13878,N_9738,N_9723);
and U13879 (N_13879,N_5782,N_6701);
xor U13880 (N_13880,N_5971,N_6747);
and U13881 (N_13881,N_6448,N_7567);
and U13882 (N_13882,N_6212,N_5675);
nor U13883 (N_13883,N_5993,N_5766);
or U13884 (N_13884,N_6655,N_8033);
or U13885 (N_13885,N_7732,N_9330);
nor U13886 (N_13886,N_5736,N_5551);
or U13887 (N_13887,N_5327,N_6120);
nor U13888 (N_13888,N_5025,N_9632);
nor U13889 (N_13889,N_9700,N_5035);
or U13890 (N_13890,N_9281,N_7653);
and U13891 (N_13891,N_7983,N_9476);
nor U13892 (N_13892,N_6994,N_8033);
xor U13893 (N_13893,N_6557,N_7775);
xor U13894 (N_13894,N_5091,N_7280);
nor U13895 (N_13895,N_8996,N_8603);
and U13896 (N_13896,N_5184,N_5440);
nor U13897 (N_13897,N_6801,N_9831);
and U13898 (N_13898,N_7029,N_8017);
nand U13899 (N_13899,N_6316,N_8022);
xor U13900 (N_13900,N_9900,N_5845);
and U13901 (N_13901,N_7175,N_7471);
and U13902 (N_13902,N_9405,N_6044);
nor U13903 (N_13903,N_9814,N_7730);
xnor U13904 (N_13904,N_7828,N_5973);
xnor U13905 (N_13905,N_6170,N_6123);
xor U13906 (N_13906,N_8411,N_8962);
or U13907 (N_13907,N_6602,N_5910);
nor U13908 (N_13908,N_9850,N_6839);
xor U13909 (N_13909,N_6023,N_5552);
nand U13910 (N_13910,N_6534,N_5502);
nand U13911 (N_13911,N_9174,N_5607);
nand U13912 (N_13912,N_5570,N_8924);
or U13913 (N_13913,N_6855,N_9614);
nor U13914 (N_13914,N_9464,N_6403);
xnor U13915 (N_13915,N_7537,N_5074);
nand U13916 (N_13916,N_6444,N_9289);
or U13917 (N_13917,N_7333,N_7700);
nand U13918 (N_13918,N_6590,N_6571);
nor U13919 (N_13919,N_6455,N_5378);
xor U13920 (N_13920,N_9443,N_6483);
nor U13921 (N_13921,N_6613,N_7302);
and U13922 (N_13922,N_5208,N_8246);
nor U13923 (N_13923,N_8292,N_9859);
and U13924 (N_13924,N_8684,N_5264);
or U13925 (N_13925,N_8610,N_9224);
and U13926 (N_13926,N_8749,N_5663);
nor U13927 (N_13927,N_8060,N_5792);
nor U13928 (N_13928,N_6676,N_9071);
xnor U13929 (N_13929,N_7395,N_5142);
or U13930 (N_13930,N_5585,N_5089);
nor U13931 (N_13931,N_6105,N_5973);
xnor U13932 (N_13932,N_7829,N_6547);
nand U13933 (N_13933,N_9472,N_5737);
xnor U13934 (N_13934,N_6751,N_8725);
nand U13935 (N_13935,N_6182,N_9131);
nor U13936 (N_13936,N_6098,N_7837);
xor U13937 (N_13937,N_9299,N_5661);
nor U13938 (N_13938,N_5022,N_7423);
or U13939 (N_13939,N_6904,N_6205);
or U13940 (N_13940,N_5103,N_9279);
and U13941 (N_13941,N_6872,N_8614);
nor U13942 (N_13942,N_7636,N_6449);
xnor U13943 (N_13943,N_5019,N_7859);
or U13944 (N_13944,N_9292,N_6825);
nand U13945 (N_13945,N_9827,N_7716);
or U13946 (N_13946,N_5069,N_7265);
nand U13947 (N_13947,N_9751,N_7093);
nand U13948 (N_13948,N_9959,N_6536);
nor U13949 (N_13949,N_9454,N_8682);
xnor U13950 (N_13950,N_9216,N_5605);
or U13951 (N_13951,N_5822,N_9987);
nand U13952 (N_13952,N_9326,N_5768);
nor U13953 (N_13953,N_6233,N_9828);
nand U13954 (N_13954,N_8208,N_5852);
or U13955 (N_13955,N_7220,N_7459);
or U13956 (N_13956,N_5780,N_7238);
and U13957 (N_13957,N_9224,N_5036);
xor U13958 (N_13958,N_6909,N_7652);
and U13959 (N_13959,N_7502,N_7063);
xor U13960 (N_13960,N_6581,N_6697);
and U13961 (N_13961,N_9818,N_7841);
nor U13962 (N_13962,N_6411,N_5098);
nor U13963 (N_13963,N_9313,N_8201);
or U13964 (N_13964,N_7542,N_5948);
or U13965 (N_13965,N_8590,N_9391);
nand U13966 (N_13966,N_8173,N_5140);
nand U13967 (N_13967,N_9284,N_5243);
xor U13968 (N_13968,N_8891,N_8397);
nand U13969 (N_13969,N_7144,N_8069);
and U13970 (N_13970,N_7892,N_6056);
xor U13971 (N_13971,N_9721,N_6669);
or U13972 (N_13972,N_5995,N_9410);
or U13973 (N_13973,N_6659,N_9655);
nor U13974 (N_13974,N_6942,N_7628);
and U13975 (N_13975,N_8849,N_5975);
nor U13976 (N_13976,N_5418,N_9114);
nor U13977 (N_13977,N_6257,N_7971);
nand U13978 (N_13978,N_5667,N_5566);
nand U13979 (N_13979,N_7844,N_9213);
xnor U13980 (N_13980,N_6969,N_8137);
or U13981 (N_13981,N_9826,N_5099);
or U13982 (N_13982,N_6811,N_6145);
nand U13983 (N_13983,N_7232,N_9231);
nand U13984 (N_13984,N_7721,N_7472);
and U13985 (N_13985,N_5257,N_9591);
xor U13986 (N_13986,N_5547,N_8482);
nand U13987 (N_13987,N_5977,N_6136);
nand U13988 (N_13988,N_6781,N_6099);
nor U13989 (N_13989,N_8274,N_7945);
or U13990 (N_13990,N_6181,N_8732);
or U13991 (N_13991,N_6501,N_9190);
or U13992 (N_13992,N_9798,N_9077);
xor U13993 (N_13993,N_9322,N_9245);
or U13994 (N_13994,N_5765,N_5867);
or U13995 (N_13995,N_7911,N_8007);
nand U13996 (N_13996,N_5321,N_5123);
or U13997 (N_13997,N_7299,N_6024);
and U13998 (N_13998,N_9436,N_9646);
xor U13999 (N_13999,N_8838,N_5588);
xnor U14000 (N_14000,N_5882,N_6047);
or U14001 (N_14001,N_9960,N_9082);
and U14002 (N_14002,N_8213,N_6375);
xor U14003 (N_14003,N_8511,N_6393);
xnor U14004 (N_14004,N_8960,N_5042);
nand U14005 (N_14005,N_7530,N_6990);
or U14006 (N_14006,N_8786,N_6651);
nor U14007 (N_14007,N_7073,N_6338);
nand U14008 (N_14008,N_9917,N_7010);
and U14009 (N_14009,N_9514,N_6437);
nand U14010 (N_14010,N_8527,N_9322);
nor U14011 (N_14011,N_6712,N_9465);
nand U14012 (N_14012,N_5345,N_9849);
xor U14013 (N_14013,N_9810,N_6324);
and U14014 (N_14014,N_5078,N_8391);
nor U14015 (N_14015,N_9828,N_5066);
nand U14016 (N_14016,N_8194,N_7706);
or U14017 (N_14017,N_9674,N_7712);
nand U14018 (N_14018,N_7157,N_7646);
nor U14019 (N_14019,N_5265,N_7613);
or U14020 (N_14020,N_7213,N_8488);
nand U14021 (N_14021,N_8392,N_9875);
and U14022 (N_14022,N_8713,N_9773);
xor U14023 (N_14023,N_8773,N_5545);
and U14024 (N_14024,N_7857,N_8608);
or U14025 (N_14025,N_6130,N_6303);
nand U14026 (N_14026,N_8347,N_8717);
or U14027 (N_14027,N_9080,N_6919);
nand U14028 (N_14028,N_5419,N_6799);
and U14029 (N_14029,N_8469,N_6624);
nand U14030 (N_14030,N_5209,N_7269);
or U14031 (N_14031,N_8146,N_8238);
nand U14032 (N_14032,N_9309,N_5766);
nor U14033 (N_14033,N_7942,N_5553);
nand U14034 (N_14034,N_6750,N_9163);
xor U14035 (N_14035,N_9704,N_8118);
nand U14036 (N_14036,N_7285,N_9038);
xor U14037 (N_14037,N_7189,N_6711);
or U14038 (N_14038,N_5597,N_8734);
xnor U14039 (N_14039,N_8173,N_6334);
or U14040 (N_14040,N_5575,N_6536);
xor U14041 (N_14041,N_5806,N_8407);
or U14042 (N_14042,N_5240,N_5408);
nand U14043 (N_14043,N_9979,N_6756);
nand U14044 (N_14044,N_7018,N_9822);
nor U14045 (N_14045,N_8343,N_6713);
nor U14046 (N_14046,N_5798,N_6959);
nor U14047 (N_14047,N_8423,N_7789);
or U14048 (N_14048,N_8848,N_6213);
and U14049 (N_14049,N_6440,N_9751);
nand U14050 (N_14050,N_9421,N_5019);
xnor U14051 (N_14051,N_6941,N_7795);
nor U14052 (N_14052,N_7256,N_6954);
or U14053 (N_14053,N_7631,N_6031);
nor U14054 (N_14054,N_6095,N_7553);
or U14055 (N_14055,N_9707,N_9514);
nor U14056 (N_14056,N_8684,N_7506);
or U14057 (N_14057,N_6966,N_8379);
nor U14058 (N_14058,N_9139,N_5981);
xnor U14059 (N_14059,N_8997,N_5852);
nor U14060 (N_14060,N_8617,N_9797);
nor U14061 (N_14061,N_6786,N_8149);
and U14062 (N_14062,N_7043,N_6907);
and U14063 (N_14063,N_9968,N_7305);
nor U14064 (N_14064,N_7816,N_9858);
nor U14065 (N_14065,N_7396,N_5663);
and U14066 (N_14066,N_9058,N_6509);
nand U14067 (N_14067,N_8808,N_5769);
and U14068 (N_14068,N_8450,N_9277);
xor U14069 (N_14069,N_6273,N_9018);
nor U14070 (N_14070,N_8951,N_9842);
nor U14071 (N_14071,N_7626,N_5243);
xor U14072 (N_14072,N_7153,N_7879);
or U14073 (N_14073,N_8876,N_6725);
nand U14074 (N_14074,N_8593,N_7440);
nand U14075 (N_14075,N_8436,N_7957);
or U14076 (N_14076,N_7687,N_7486);
nor U14077 (N_14077,N_6712,N_7995);
nand U14078 (N_14078,N_8487,N_8965);
or U14079 (N_14079,N_6698,N_6049);
xor U14080 (N_14080,N_9599,N_7626);
and U14081 (N_14081,N_5081,N_5302);
and U14082 (N_14082,N_7116,N_7871);
nor U14083 (N_14083,N_7237,N_6071);
and U14084 (N_14084,N_9861,N_6586);
xor U14085 (N_14085,N_5088,N_7876);
and U14086 (N_14086,N_5218,N_8701);
nand U14087 (N_14087,N_8192,N_6525);
and U14088 (N_14088,N_9134,N_8921);
or U14089 (N_14089,N_5619,N_7637);
nand U14090 (N_14090,N_9262,N_9769);
or U14091 (N_14091,N_6089,N_9819);
nor U14092 (N_14092,N_8163,N_5971);
or U14093 (N_14093,N_8140,N_8349);
nand U14094 (N_14094,N_7250,N_6387);
and U14095 (N_14095,N_9901,N_5049);
or U14096 (N_14096,N_9753,N_6186);
nand U14097 (N_14097,N_5143,N_7718);
nor U14098 (N_14098,N_8017,N_5678);
nor U14099 (N_14099,N_6721,N_5652);
xnor U14100 (N_14100,N_7904,N_9502);
nand U14101 (N_14101,N_6389,N_7132);
nor U14102 (N_14102,N_5174,N_6527);
xor U14103 (N_14103,N_7538,N_8550);
nand U14104 (N_14104,N_7537,N_5495);
nand U14105 (N_14105,N_8096,N_7051);
or U14106 (N_14106,N_9109,N_7014);
nand U14107 (N_14107,N_5445,N_6003);
nand U14108 (N_14108,N_6541,N_9310);
nor U14109 (N_14109,N_8535,N_5894);
nor U14110 (N_14110,N_5820,N_7039);
or U14111 (N_14111,N_5678,N_6587);
or U14112 (N_14112,N_7595,N_6754);
xnor U14113 (N_14113,N_7428,N_6611);
nand U14114 (N_14114,N_7436,N_9846);
or U14115 (N_14115,N_5320,N_9519);
nor U14116 (N_14116,N_6432,N_9095);
or U14117 (N_14117,N_6830,N_9559);
and U14118 (N_14118,N_6634,N_6550);
xnor U14119 (N_14119,N_5675,N_9564);
and U14120 (N_14120,N_5086,N_7102);
nor U14121 (N_14121,N_6941,N_9621);
and U14122 (N_14122,N_6606,N_7831);
nor U14123 (N_14123,N_5763,N_5482);
xnor U14124 (N_14124,N_6022,N_5373);
nor U14125 (N_14125,N_8034,N_6703);
xnor U14126 (N_14126,N_7697,N_6063);
or U14127 (N_14127,N_9892,N_6093);
or U14128 (N_14128,N_9339,N_8990);
xor U14129 (N_14129,N_9524,N_6168);
xor U14130 (N_14130,N_5533,N_6233);
nand U14131 (N_14131,N_6211,N_9062);
nor U14132 (N_14132,N_7822,N_9920);
and U14133 (N_14133,N_9606,N_7410);
nor U14134 (N_14134,N_5762,N_9694);
nor U14135 (N_14135,N_6081,N_8278);
and U14136 (N_14136,N_6522,N_7523);
or U14137 (N_14137,N_5835,N_7021);
xor U14138 (N_14138,N_7556,N_6473);
nand U14139 (N_14139,N_5751,N_5990);
or U14140 (N_14140,N_9646,N_9381);
nand U14141 (N_14141,N_9289,N_6941);
or U14142 (N_14142,N_9645,N_6675);
or U14143 (N_14143,N_7521,N_8793);
xor U14144 (N_14144,N_9938,N_6555);
xnor U14145 (N_14145,N_9826,N_7584);
or U14146 (N_14146,N_5111,N_7090);
and U14147 (N_14147,N_6496,N_6461);
or U14148 (N_14148,N_6091,N_7072);
and U14149 (N_14149,N_8961,N_8461);
xnor U14150 (N_14150,N_6534,N_7835);
xor U14151 (N_14151,N_6421,N_8153);
and U14152 (N_14152,N_5142,N_8361);
nand U14153 (N_14153,N_8481,N_9152);
or U14154 (N_14154,N_9159,N_8313);
nor U14155 (N_14155,N_9853,N_8620);
xnor U14156 (N_14156,N_9061,N_8683);
nor U14157 (N_14157,N_6731,N_6378);
or U14158 (N_14158,N_8275,N_8289);
or U14159 (N_14159,N_5029,N_5689);
and U14160 (N_14160,N_9144,N_5537);
nand U14161 (N_14161,N_8579,N_7562);
nand U14162 (N_14162,N_5390,N_7304);
xor U14163 (N_14163,N_6170,N_8681);
or U14164 (N_14164,N_9227,N_9857);
and U14165 (N_14165,N_9580,N_9028);
and U14166 (N_14166,N_7020,N_6931);
or U14167 (N_14167,N_9022,N_6401);
xor U14168 (N_14168,N_7987,N_8798);
nand U14169 (N_14169,N_8204,N_9158);
nand U14170 (N_14170,N_5115,N_6039);
nand U14171 (N_14171,N_9018,N_5341);
xnor U14172 (N_14172,N_9805,N_5718);
or U14173 (N_14173,N_9095,N_8528);
nor U14174 (N_14174,N_9822,N_9624);
nor U14175 (N_14175,N_9709,N_8615);
nor U14176 (N_14176,N_6343,N_5191);
and U14177 (N_14177,N_9889,N_8561);
nor U14178 (N_14178,N_5352,N_9092);
and U14179 (N_14179,N_9116,N_6926);
or U14180 (N_14180,N_8004,N_5362);
xnor U14181 (N_14181,N_9375,N_9903);
nand U14182 (N_14182,N_7900,N_7886);
nand U14183 (N_14183,N_7584,N_6943);
and U14184 (N_14184,N_9312,N_8720);
xnor U14185 (N_14185,N_9386,N_8054);
or U14186 (N_14186,N_7793,N_8872);
or U14187 (N_14187,N_8281,N_9362);
nand U14188 (N_14188,N_6419,N_9209);
nand U14189 (N_14189,N_5703,N_7228);
xor U14190 (N_14190,N_6966,N_6273);
nand U14191 (N_14191,N_9940,N_6510);
xnor U14192 (N_14192,N_5217,N_6051);
and U14193 (N_14193,N_8810,N_6145);
and U14194 (N_14194,N_9821,N_5298);
nor U14195 (N_14195,N_5798,N_6166);
and U14196 (N_14196,N_9274,N_7068);
or U14197 (N_14197,N_6405,N_8981);
nand U14198 (N_14198,N_8069,N_9519);
nor U14199 (N_14199,N_9041,N_5698);
nand U14200 (N_14200,N_9712,N_5233);
xor U14201 (N_14201,N_9827,N_8031);
and U14202 (N_14202,N_7650,N_6599);
or U14203 (N_14203,N_5222,N_7265);
or U14204 (N_14204,N_5586,N_5848);
nand U14205 (N_14205,N_8703,N_8682);
xnor U14206 (N_14206,N_7440,N_5969);
and U14207 (N_14207,N_7206,N_8284);
nand U14208 (N_14208,N_5707,N_7651);
nor U14209 (N_14209,N_9748,N_9463);
nand U14210 (N_14210,N_9405,N_8928);
and U14211 (N_14211,N_8252,N_8434);
nor U14212 (N_14212,N_6472,N_7233);
nand U14213 (N_14213,N_9927,N_6800);
or U14214 (N_14214,N_9198,N_9563);
or U14215 (N_14215,N_8173,N_7893);
nor U14216 (N_14216,N_7516,N_5470);
nor U14217 (N_14217,N_5951,N_9622);
or U14218 (N_14218,N_5694,N_5803);
and U14219 (N_14219,N_7629,N_5128);
or U14220 (N_14220,N_6679,N_8819);
nor U14221 (N_14221,N_8120,N_9098);
and U14222 (N_14222,N_9276,N_8721);
nor U14223 (N_14223,N_9633,N_8362);
xnor U14224 (N_14224,N_5713,N_5224);
nor U14225 (N_14225,N_5913,N_6593);
xnor U14226 (N_14226,N_9780,N_6520);
xor U14227 (N_14227,N_6257,N_8186);
nand U14228 (N_14228,N_8648,N_8007);
or U14229 (N_14229,N_9448,N_7317);
nand U14230 (N_14230,N_8105,N_9456);
or U14231 (N_14231,N_5645,N_9709);
or U14232 (N_14232,N_7133,N_7346);
nor U14233 (N_14233,N_6659,N_9171);
nand U14234 (N_14234,N_6412,N_5860);
or U14235 (N_14235,N_6167,N_9832);
xnor U14236 (N_14236,N_9510,N_5035);
nor U14237 (N_14237,N_6612,N_8279);
and U14238 (N_14238,N_8729,N_8917);
and U14239 (N_14239,N_5442,N_6260);
and U14240 (N_14240,N_6831,N_5583);
nand U14241 (N_14241,N_8217,N_5709);
nand U14242 (N_14242,N_8939,N_6569);
or U14243 (N_14243,N_5361,N_6268);
xor U14244 (N_14244,N_7601,N_5829);
or U14245 (N_14245,N_7366,N_6811);
or U14246 (N_14246,N_9363,N_5365);
and U14247 (N_14247,N_8704,N_7713);
or U14248 (N_14248,N_7970,N_9973);
nand U14249 (N_14249,N_9010,N_9618);
xnor U14250 (N_14250,N_6609,N_7174);
nand U14251 (N_14251,N_8269,N_6796);
or U14252 (N_14252,N_9271,N_9487);
xnor U14253 (N_14253,N_7159,N_9189);
or U14254 (N_14254,N_5791,N_5740);
nand U14255 (N_14255,N_8039,N_5899);
and U14256 (N_14256,N_6282,N_8742);
xnor U14257 (N_14257,N_7894,N_8615);
or U14258 (N_14258,N_9091,N_6468);
nand U14259 (N_14259,N_9682,N_8229);
and U14260 (N_14260,N_6081,N_8072);
and U14261 (N_14261,N_6366,N_7087);
nor U14262 (N_14262,N_5519,N_5491);
and U14263 (N_14263,N_9422,N_8131);
nor U14264 (N_14264,N_8139,N_8592);
and U14265 (N_14265,N_9793,N_6721);
nor U14266 (N_14266,N_8354,N_8118);
nand U14267 (N_14267,N_8803,N_7450);
or U14268 (N_14268,N_8602,N_8701);
or U14269 (N_14269,N_5851,N_6101);
xnor U14270 (N_14270,N_9712,N_6535);
nand U14271 (N_14271,N_9958,N_5805);
and U14272 (N_14272,N_6195,N_8873);
nand U14273 (N_14273,N_6534,N_5528);
nor U14274 (N_14274,N_7321,N_5069);
or U14275 (N_14275,N_9751,N_8982);
nand U14276 (N_14276,N_7806,N_6755);
xor U14277 (N_14277,N_9400,N_6211);
and U14278 (N_14278,N_8092,N_7850);
xor U14279 (N_14279,N_5011,N_7784);
xor U14280 (N_14280,N_5026,N_9971);
nor U14281 (N_14281,N_5413,N_7143);
nor U14282 (N_14282,N_8361,N_5024);
or U14283 (N_14283,N_5126,N_7280);
nor U14284 (N_14284,N_9346,N_8290);
and U14285 (N_14285,N_7531,N_8328);
and U14286 (N_14286,N_6456,N_6465);
nand U14287 (N_14287,N_5356,N_6955);
or U14288 (N_14288,N_6804,N_9859);
xnor U14289 (N_14289,N_5509,N_7983);
or U14290 (N_14290,N_7123,N_6435);
and U14291 (N_14291,N_8359,N_5592);
nor U14292 (N_14292,N_8096,N_7481);
nor U14293 (N_14293,N_7897,N_9046);
nand U14294 (N_14294,N_8102,N_6666);
xor U14295 (N_14295,N_8466,N_5578);
nand U14296 (N_14296,N_7540,N_8180);
or U14297 (N_14297,N_7638,N_5968);
and U14298 (N_14298,N_5394,N_5389);
and U14299 (N_14299,N_5186,N_7519);
and U14300 (N_14300,N_8611,N_6459);
xor U14301 (N_14301,N_8637,N_5151);
or U14302 (N_14302,N_6068,N_9248);
nor U14303 (N_14303,N_8571,N_8650);
nor U14304 (N_14304,N_9850,N_9207);
or U14305 (N_14305,N_8636,N_7268);
xnor U14306 (N_14306,N_6240,N_8638);
nand U14307 (N_14307,N_9358,N_7637);
xnor U14308 (N_14308,N_5980,N_9056);
or U14309 (N_14309,N_8650,N_5727);
or U14310 (N_14310,N_5100,N_5527);
nand U14311 (N_14311,N_9962,N_7713);
nand U14312 (N_14312,N_9314,N_6667);
nand U14313 (N_14313,N_6735,N_6015);
nor U14314 (N_14314,N_7578,N_5799);
or U14315 (N_14315,N_5241,N_6419);
and U14316 (N_14316,N_6346,N_8123);
and U14317 (N_14317,N_7505,N_5810);
nand U14318 (N_14318,N_5866,N_7589);
xor U14319 (N_14319,N_8054,N_7050);
nor U14320 (N_14320,N_8215,N_5674);
and U14321 (N_14321,N_8236,N_6941);
nor U14322 (N_14322,N_8519,N_5372);
and U14323 (N_14323,N_7144,N_6011);
nor U14324 (N_14324,N_8525,N_8190);
nand U14325 (N_14325,N_8903,N_7667);
nand U14326 (N_14326,N_9241,N_8979);
nand U14327 (N_14327,N_5797,N_6348);
xor U14328 (N_14328,N_9762,N_7166);
nand U14329 (N_14329,N_8465,N_7221);
xor U14330 (N_14330,N_7644,N_6509);
nor U14331 (N_14331,N_9759,N_7681);
and U14332 (N_14332,N_8515,N_6192);
nor U14333 (N_14333,N_6970,N_6984);
nor U14334 (N_14334,N_9081,N_8891);
nor U14335 (N_14335,N_8428,N_9855);
nor U14336 (N_14336,N_5269,N_8301);
xor U14337 (N_14337,N_7858,N_7043);
and U14338 (N_14338,N_5975,N_6679);
xnor U14339 (N_14339,N_5907,N_8116);
xor U14340 (N_14340,N_5772,N_8834);
or U14341 (N_14341,N_6085,N_8585);
nand U14342 (N_14342,N_8685,N_6608);
xnor U14343 (N_14343,N_5113,N_6297);
nor U14344 (N_14344,N_6204,N_6604);
and U14345 (N_14345,N_5616,N_6766);
or U14346 (N_14346,N_6617,N_6685);
xnor U14347 (N_14347,N_8645,N_7462);
nand U14348 (N_14348,N_7085,N_6565);
or U14349 (N_14349,N_8998,N_9919);
nand U14350 (N_14350,N_7215,N_5851);
or U14351 (N_14351,N_7145,N_8856);
or U14352 (N_14352,N_7896,N_7247);
nand U14353 (N_14353,N_7393,N_6123);
and U14354 (N_14354,N_7309,N_5858);
and U14355 (N_14355,N_9595,N_6841);
nor U14356 (N_14356,N_5142,N_7331);
nor U14357 (N_14357,N_9649,N_7096);
or U14358 (N_14358,N_8086,N_5206);
nand U14359 (N_14359,N_7150,N_9895);
nor U14360 (N_14360,N_9374,N_9577);
nand U14361 (N_14361,N_9928,N_7664);
or U14362 (N_14362,N_5008,N_9587);
nor U14363 (N_14363,N_5108,N_6839);
or U14364 (N_14364,N_7596,N_6604);
xnor U14365 (N_14365,N_7223,N_9203);
xnor U14366 (N_14366,N_9952,N_5739);
nand U14367 (N_14367,N_8668,N_7733);
nand U14368 (N_14368,N_7987,N_6671);
xor U14369 (N_14369,N_8221,N_5604);
nor U14370 (N_14370,N_8388,N_7808);
nand U14371 (N_14371,N_9338,N_8793);
nor U14372 (N_14372,N_9423,N_6449);
nor U14373 (N_14373,N_9663,N_5209);
xor U14374 (N_14374,N_5730,N_7840);
nor U14375 (N_14375,N_5990,N_6244);
nor U14376 (N_14376,N_6183,N_5832);
xnor U14377 (N_14377,N_5888,N_6901);
nand U14378 (N_14378,N_5735,N_7863);
and U14379 (N_14379,N_6653,N_7032);
nor U14380 (N_14380,N_9150,N_7618);
and U14381 (N_14381,N_9783,N_5804);
nand U14382 (N_14382,N_8450,N_7658);
xor U14383 (N_14383,N_6997,N_8813);
or U14384 (N_14384,N_5533,N_9156);
and U14385 (N_14385,N_5719,N_5703);
nand U14386 (N_14386,N_7537,N_8037);
nor U14387 (N_14387,N_6466,N_7710);
nor U14388 (N_14388,N_6133,N_9702);
or U14389 (N_14389,N_9997,N_6165);
nor U14390 (N_14390,N_6477,N_8749);
nand U14391 (N_14391,N_9368,N_7451);
and U14392 (N_14392,N_5489,N_8682);
or U14393 (N_14393,N_9565,N_9079);
nor U14394 (N_14394,N_7853,N_5058);
nand U14395 (N_14395,N_8352,N_7584);
nand U14396 (N_14396,N_6587,N_9534);
xor U14397 (N_14397,N_6120,N_8496);
or U14398 (N_14398,N_6706,N_9194);
xnor U14399 (N_14399,N_9336,N_9079);
nand U14400 (N_14400,N_7722,N_8747);
and U14401 (N_14401,N_9399,N_6393);
nor U14402 (N_14402,N_5952,N_6261);
nand U14403 (N_14403,N_7170,N_8852);
nor U14404 (N_14404,N_5712,N_5925);
or U14405 (N_14405,N_9452,N_5044);
xnor U14406 (N_14406,N_6679,N_7622);
nor U14407 (N_14407,N_9836,N_6196);
nor U14408 (N_14408,N_6144,N_5029);
and U14409 (N_14409,N_8419,N_8596);
xnor U14410 (N_14410,N_8484,N_7646);
nand U14411 (N_14411,N_9485,N_8212);
nor U14412 (N_14412,N_9217,N_6185);
nand U14413 (N_14413,N_6737,N_5804);
xnor U14414 (N_14414,N_8540,N_6650);
and U14415 (N_14415,N_5045,N_6583);
or U14416 (N_14416,N_5403,N_7156);
and U14417 (N_14417,N_7595,N_7345);
xnor U14418 (N_14418,N_8544,N_8998);
xnor U14419 (N_14419,N_5709,N_9335);
xor U14420 (N_14420,N_7565,N_8582);
xor U14421 (N_14421,N_5891,N_6547);
or U14422 (N_14422,N_9997,N_8172);
or U14423 (N_14423,N_6187,N_8830);
xor U14424 (N_14424,N_9118,N_5038);
nand U14425 (N_14425,N_8791,N_5856);
nand U14426 (N_14426,N_6285,N_6820);
xnor U14427 (N_14427,N_6983,N_9669);
nand U14428 (N_14428,N_7960,N_7166);
or U14429 (N_14429,N_5582,N_7300);
nor U14430 (N_14430,N_7354,N_5131);
nor U14431 (N_14431,N_5437,N_8944);
xor U14432 (N_14432,N_9690,N_5952);
nand U14433 (N_14433,N_9341,N_5703);
or U14434 (N_14434,N_9250,N_7879);
or U14435 (N_14435,N_8400,N_9915);
nor U14436 (N_14436,N_7001,N_9605);
nor U14437 (N_14437,N_6670,N_6498);
nand U14438 (N_14438,N_5742,N_7897);
xor U14439 (N_14439,N_9198,N_9319);
nand U14440 (N_14440,N_9613,N_5513);
or U14441 (N_14441,N_5702,N_9723);
nor U14442 (N_14442,N_8916,N_5052);
nand U14443 (N_14443,N_7446,N_5770);
xor U14444 (N_14444,N_5583,N_7494);
or U14445 (N_14445,N_7162,N_5230);
xnor U14446 (N_14446,N_6830,N_9285);
nand U14447 (N_14447,N_6350,N_9880);
and U14448 (N_14448,N_7126,N_9785);
nor U14449 (N_14449,N_5889,N_8442);
or U14450 (N_14450,N_7068,N_8405);
nand U14451 (N_14451,N_9891,N_6717);
nor U14452 (N_14452,N_7181,N_9158);
xor U14453 (N_14453,N_7741,N_6523);
and U14454 (N_14454,N_8578,N_6277);
xor U14455 (N_14455,N_8118,N_7536);
and U14456 (N_14456,N_7021,N_6893);
nand U14457 (N_14457,N_9831,N_9430);
nand U14458 (N_14458,N_7156,N_6155);
xnor U14459 (N_14459,N_5787,N_6439);
xnor U14460 (N_14460,N_5636,N_7938);
xor U14461 (N_14461,N_9096,N_5245);
nor U14462 (N_14462,N_5258,N_9997);
or U14463 (N_14463,N_6301,N_8574);
nand U14464 (N_14464,N_6751,N_8968);
nand U14465 (N_14465,N_6234,N_7537);
and U14466 (N_14466,N_7029,N_7389);
and U14467 (N_14467,N_8387,N_6789);
or U14468 (N_14468,N_6560,N_5840);
nor U14469 (N_14469,N_5153,N_6118);
xnor U14470 (N_14470,N_8159,N_7666);
nand U14471 (N_14471,N_9036,N_6632);
xor U14472 (N_14472,N_6084,N_7171);
and U14473 (N_14473,N_7192,N_7957);
and U14474 (N_14474,N_9305,N_8561);
nor U14475 (N_14475,N_5196,N_7141);
nand U14476 (N_14476,N_8094,N_5419);
and U14477 (N_14477,N_5615,N_9063);
nor U14478 (N_14478,N_5904,N_6856);
nor U14479 (N_14479,N_6416,N_5040);
xnor U14480 (N_14480,N_6431,N_8184);
nor U14481 (N_14481,N_7607,N_9332);
nand U14482 (N_14482,N_9770,N_5739);
nor U14483 (N_14483,N_7518,N_6006);
or U14484 (N_14484,N_9926,N_5077);
or U14485 (N_14485,N_8426,N_6995);
nor U14486 (N_14486,N_8278,N_5495);
xor U14487 (N_14487,N_6741,N_9977);
or U14488 (N_14488,N_5189,N_6040);
nand U14489 (N_14489,N_8013,N_5977);
nand U14490 (N_14490,N_8222,N_6599);
or U14491 (N_14491,N_9454,N_9412);
xor U14492 (N_14492,N_9167,N_7950);
xnor U14493 (N_14493,N_9823,N_9927);
xor U14494 (N_14494,N_9945,N_5134);
nand U14495 (N_14495,N_9231,N_8908);
nor U14496 (N_14496,N_9215,N_5008);
or U14497 (N_14497,N_5791,N_7230);
or U14498 (N_14498,N_7849,N_9972);
nand U14499 (N_14499,N_6533,N_5263);
nor U14500 (N_14500,N_6916,N_8079);
nor U14501 (N_14501,N_5032,N_6163);
nor U14502 (N_14502,N_8841,N_9104);
or U14503 (N_14503,N_7056,N_8193);
and U14504 (N_14504,N_5759,N_7966);
nand U14505 (N_14505,N_8378,N_7133);
nand U14506 (N_14506,N_9105,N_9339);
or U14507 (N_14507,N_9100,N_8982);
nand U14508 (N_14508,N_8630,N_7798);
nand U14509 (N_14509,N_7617,N_5713);
nand U14510 (N_14510,N_5553,N_9093);
xor U14511 (N_14511,N_9006,N_8825);
nor U14512 (N_14512,N_5192,N_9497);
and U14513 (N_14513,N_5740,N_6194);
or U14514 (N_14514,N_9683,N_7069);
or U14515 (N_14515,N_7975,N_9584);
nand U14516 (N_14516,N_7276,N_6807);
nand U14517 (N_14517,N_8860,N_8065);
or U14518 (N_14518,N_6373,N_8117);
or U14519 (N_14519,N_5023,N_6416);
or U14520 (N_14520,N_7247,N_9302);
xor U14521 (N_14521,N_6978,N_7301);
nor U14522 (N_14522,N_7042,N_6519);
or U14523 (N_14523,N_5563,N_8482);
or U14524 (N_14524,N_8702,N_7783);
and U14525 (N_14525,N_6213,N_8628);
nor U14526 (N_14526,N_8067,N_9718);
nand U14527 (N_14527,N_9993,N_9189);
nand U14528 (N_14528,N_5312,N_5648);
and U14529 (N_14529,N_6136,N_5011);
xnor U14530 (N_14530,N_7014,N_5347);
xnor U14531 (N_14531,N_8565,N_7279);
nor U14532 (N_14532,N_7532,N_7246);
or U14533 (N_14533,N_5706,N_9128);
xnor U14534 (N_14534,N_8463,N_6379);
nor U14535 (N_14535,N_7604,N_6122);
nor U14536 (N_14536,N_8361,N_8334);
nor U14537 (N_14537,N_7260,N_5413);
or U14538 (N_14538,N_7521,N_9276);
nor U14539 (N_14539,N_8694,N_7438);
nor U14540 (N_14540,N_6660,N_8015);
and U14541 (N_14541,N_5815,N_8446);
nand U14542 (N_14542,N_9936,N_7267);
or U14543 (N_14543,N_7733,N_5892);
nor U14544 (N_14544,N_9441,N_8597);
xnor U14545 (N_14545,N_6345,N_6542);
and U14546 (N_14546,N_9273,N_5829);
xor U14547 (N_14547,N_8764,N_6851);
nand U14548 (N_14548,N_5762,N_8147);
nand U14549 (N_14549,N_6595,N_7083);
nand U14550 (N_14550,N_8569,N_9434);
nand U14551 (N_14551,N_8862,N_9006);
or U14552 (N_14552,N_5331,N_8874);
nand U14553 (N_14553,N_9751,N_6653);
nand U14554 (N_14554,N_5079,N_6346);
nand U14555 (N_14555,N_8829,N_5615);
and U14556 (N_14556,N_5972,N_6450);
or U14557 (N_14557,N_9301,N_9228);
nor U14558 (N_14558,N_7860,N_7897);
or U14559 (N_14559,N_9386,N_5400);
nand U14560 (N_14560,N_5950,N_7731);
nand U14561 (N_14561,N_7164,N_9150);
and U14562 (N_14562,N_7349,N_7861);
nor U14563 (N_14563,N_8781,N_8601);
and U14564 (N_14564,N_5003,N_9132);
nand U14565 (N_14565,N_7114,N_6475);
or U14566 (N_14566,N_7286,N_7591);
or U14567 (N_14567,N_9579,N_6469);
nand U14568 (N_14568,N_6512,N_7348);
or U14569 (N_14569,N_6338,N_8428);
and U14570 (N_14570,N_5354,N_8395);
and U14571 (N_14571,N_6249,N_6985);
and U14572 (N_14572,N_9081,N_9411);
xor U14573 (N_14573,N_9735,N_9873);
nor U14574 (N_14574,N_5775,N_5896);
and U14575 (N_14575,N_8981,N_5050);
or U14576 (N_14576,N_8151,N_8495);
nor U14577 (N_14577,N_9550,N_7999);
xor U14578 (N_14578,N_6848,N_7890);
xor U14579 (N_14579,N_9880,N_6511);
or U14580 (N_14580,N_8992,N_8166);
nor U14581 (N_14581,N_6982,N_6572);
xnor U14582 (N_14582,N_8912,N_6569);
and U14583 (N_14583,N_9148,N_8655);
and U14584 (N_14584,N_5485,N_9671);
or U14585 (N_14585,N_5653,N_8052);
and U14586 (N_14586,N_8964,N_6020);
nor U14587 (N_14587,N_6462,N_6452);
xor U14588 (N_14588,N_8992,N_5606);
nand U14589 (N_14589,N_8467,N_7888);
or U14590 (N_14590,N_5872,N_7430);
or U14591 (N_14591,N_7792,N_6152);
nand U14592 (N_14592,N_9397,N_9157);
and U14593 (N_14593,N_6045,N_5306);
and U14594 (N_14594,N_5837,N_5895);
and U14595 (N_14595,N_8195,N_6396);
xor U14596 (N_14596,N_9970,N_9483);
xnor U14597 (N_14597,N_5471,N_8797);
or U14598 (N_14598,N_9384,N_9899);
xnor U14599 (N_14599,N_5714,N_9019);
or U14600 (N_14600,N_8595,N_9528);
nor U14601 (N_14601,N_7534,N_8682);
nand U14602 (N_14602,N_9665,N_5248);
xor U14603 (N_14603,N_8183,N_6922);
or U14604 (N_14604,N_7034,N_6338);
and U14605 (N_14605,N_6255,N_9746);
and U14606 (N_14606,N_6155,N_5553);
and U14607 (N_14607,N_9174,N_6876);
or U14608 (N_14608,N_6527,N_8149);
or U14609 (N_14609,N_8527,N_9794);
xor U14610 (N_14610,N_6866,N_6578);
and U14611 (N_14611,N_6061,N_5743);
nor U14612 (N_14612,N_6011,N_6848);
and U14613 (N_14613,N_5524,N_9350);
and U14614 (N_14614,N_6661,N_8355);
and U14615 (N_14615,N_6649,N_7934);
xnor U14616 (N_14616,N_8012,N_5533);
or U14617 (N_14617,N_6132,N_8122);
and U14618 (N_14618,N_9685,N_9249);
or U14619 (N_14619,N_9734,N_5408);
nand U14620 (N_14620,N_8265,N_8637);
xnor U14621 (N_14621,N_6994,N_7692);
xnor U14622 (N_14622,N_7354,N_7598);
or U14623 (N_14623,N_5076,N_7501);
xnor U14624 (N_14624,N_7041,N_8071);
nand U14625 (N_14625,N_5658,N_9412);
xor U14626 (N_14626,N_7381,N_8607);
nand U14627 (N_14627,N_6199,N_8047);
or U14628 (N_14628,N_6392,N_9359);
nand U14629 (N_14629,N_5881,N_9465);
nand U14630 (N_14630,N_7369,N_6971);
nor U14631 (N_14631,N_6729,N_6415);
nor U14632 (N_14632,N_9041,N_9542);
nor U14633 (N_14633,N_6051,N_5288);
and U14634 (N_14634,N_7744,N_9754);
nand U14635 (N_14635,N_9478,N_8328);
xor U14636 (N_14636,N_8782,N_6042);
xnor U14637 (N_14637,N_7952,N_6450);
nor U14638 (N_14638,N_9975,N_8557);
and U14639 (N_14639,N_7971,N_5424);
nand U14640 (N_14640,N_7738,N_8256);
and U14641 (N_14641,N_8968,N_6171);
and U14642 (N_14642,N_8916,N_5458);
or U14643 (N_14643,N_5729,N_5557);
nor U14644 (N_14644,N_7658,N_8326);
nor U14645 (N_14645,N_5529,N_6990);
nor U14646 (N_14646,N_7836,N_8780);
nor U14647 (N_14647,N_9535,N_7838);
nand U14648 (N_14648,N_6497,N_7806);
xor U14649 (N_14649,N_9295,N_8226);
xnor U14650 (N_14650,N_7214,N_5867);
or U14651 (N_14651,N_6887,N_9810);
nand U14652 (N_14652,N_9385,N_8947);
or U14653 (N_14653,N_5352,N_7991);
nor U14654 (N_14654,N_6322,N_7178);
xnor U14655 (N_14655,N_6347,N_7219);
nand U14656 (N_14656,N_8478,N_6966);
or U14657 (N_14657,N_5739,N_9677);
nand U14658 (N_14658,N_9133,N_6048);
or U14659 (N_14659,N_9211,N_7646);
and U14660 (N_14660,N_5498,N_5279);
and U14661 (N_14661,N_7462,N_9796);
and U14662 (N_14662,N_8992,N_6908);
nand U14663 (N_14663,N_6885,N_8738);
or U14664 (N_14664,N_6607,N_9430);
nor U14665 (N_14665,N_5417,N_7455);
nand U14666 (N_14666,N_5130,N_7260);
or U14667 (N_14667,N_5667,N_8738);
nor U14668 (N_14668,N_6270,N_9085);
nand U14669 (N_14669,N_9972,N_9214);
nor U14670 (N_14670,N_9922,N_8431);
nand U14671 (N_14671,N_8490,N_8349);
or U14672 (N_14672,N_5507,N_9733);
nand U14673 (N_14673,N_8538,N_6234);
xnor U14674 (N_14674,N_5601,N_7639);
xnor U14675 (N_14675,N_5499,N_5438);
nor U14676 (N_14676,N_6677,N_9434);
nor U14677 (N_14677,N_8591,N_8066);
nor U14678 (N_14678,N_9172,N_9691);
xnor U14679 (N_14679,N_8336,N_8000);
nor U14680 (N_14680,N_9932,N_8604);
nor U14681 (N_14681,N_8593,N_6146);
nor U14682 (N_14682,N_8321,N_5342);
nand U14683 (N_14683,N_5446,N_6622);
nor U14684 (N_14684,N_7893,N_9803);
and U14685 (N_14685,N_7569,N_8918);
or U14686 (N_14686,N_7322,N_6549);
and U14687 (N_14687,N_7152,N_9985);
xor U14688 (N_14688,N_8452,N_6298);
and U14689 (N_14689,N_5612,N_9785);
xnor U14690 (N_14690,N_6814,N_5208);
nor U14691 (N_14691,N_9011,N_9440);
nor U14692 (N_14692,N_8302,N_9323);
or U14693 (N_14693,N_9107,N_6136);
nand U14694 (N_14694,N_5331,N_9862);
nand U14695 (N_14695,N_9062,N_6182);
or U14696 (N_14696,N_5015,N_9689);
xor U14697 (N_14697,N_6127,N_7282);
xnor U14698 (N_14698,N_6925,N_6969);
nor U14699 (N_14699,N_6502,N_6100);
xnor U14700 (N_14700,N_8258,N_8901);
xor U14701 (N_14701,N_5283,N_5712);
and U14702 (N_14702,N_5027,N_6328);
xor U14703 (N_14703,N_9413,N_5161);
nand U14704 (N_14704,N_7009,N_8662);
nand U14705 (N_14705,N_7056,N_7836);
nand U14706 (N_14706,N_5276,N_7813);
or U14707 (N_14707,N_5318,N_8624);
nor U14708 (N_14708,N_7013,N_8804);
nor U14709 (N_14709,N_5254,N_8221);
nor U14710 (N_14710,N_8178,N_6015);
nand U14711 (N_14711,N_5218,N_7380);
or U14712 (N_14712,N_9939,N_5630);
or U14713 (N_14713,N_9511,N_6010);
xnor U14714 (N_14714,N_8960,N_7305);
nor U14715 (N_14715,N_7468,N_9963);
nor U14716 (N_14716,N_6029,N_8168);
xor U14717 (N_14717,N_6787,N_6311);
or U14718 (N_14718,N_5693,N_7189);
or U14719 (N_14719,N_5269,N_6028);
nand U14720 (N_14720,N_9953,N_9943);
and U14721 (N_14721,N_6760,N_6158);
nand U14722 (N_14722,N_5394,N_5403);
xnor U14723 (N_14723,N_8627,N_6062);
xnor U14724 (N_14724,N_8880,N_7380);
or U14725 (N_14725,N_7596,N_9236);
or U14726 (N_14726,N_7706,N_6692);
nor U14727 (N_14727,N_8297,N_7267);
or U14728 (N_14728,N_6709,N_5854);
nor U14729 (N_14729,N_6570,N_6721);
and U14730 (N_14730,N_8351,N_9350);
xnor U14731 (N_14731,N_7670,N_6546);
nand U14732 (N_14732,N_7460,N_6187);
and U14733 (N_14733,N_6871,N_9482);
or U14734 (N_14734,N_9280,N_7626);
and U14735 (N_14735,N_7610,N_5900);
xor U14736 (N_14736,N_6319,N_5519);
nor U14737 (N_14737,N_6883,N_7693);
nor U14738 (N_14738,N_9903,N_6609);
or U14739 (N_14739,N_5365,N_9907);
or U14740 (N_14740,N_8604,N_9125);
or U14741 (N_14741,N_6384,N_9026);
nor U14742 (N_14742,N_8845,N_8561);
nor U14743 (N_14743,N_7961,N_8521);
or U14744 (N_14744,N_9258,N_5409);
nand U14745 (N_14745,N_5392,N_6962);
xor U14746 (N_14746,N_8605,N_8671);
xnor U14747 (N_14747,N_8316,N_9710);
and U14748 (N_14748,N_8799,N_9497);
and U14749 (N_14749,N_8242,N_8585);
nand U14750 (N_14750,N_6515,N_7923);
nand U14751 (N_14751,N_8855,N_6350);
or U14752 (N_14752,N_6864,N_8002);
nor U14753 (N_14753,N_6884,N_7028);
xor U14754 (N_14754,N_6335,N_8697);
xor U14755 (N_14755,N_5084,N_5256);
nand U14756 (N_14756,N_6960,N_7719);
xnor U14757 (N_14757,N_9659,N_8369);
nor U14758 (N_14758,N_5218,N_9732);
and U14759 (N_14759,N_6177,N_8533);
nand U14760 (N_14760,N_7447,N_6315);
or U14761 (N_14761,N_5945,N_8572);
nand U14762 (N_14762,N_9136,N_6830);
or U14763 (N_14763,N_7378,N_9784);
nor U14764 (N_14764,N_9462,N_7016);
nor U14765 (N_14765,N_9352,N_5705);
or U14766 (N_14766,N_8826,N_7823);
xor U14767 (N_14767,N_9831,N_6764);
xor U14768 (N_14768,N_6267,N_8172);
or U14769 (N_14769,N_9251,N_6301);
nor U14770 (N_14770,N_8491,N_8427);
and U14771 (N_14771,N_5433,N_5997);
xnor U14772 (N_14772,N_9408,N_6403);
or U14773 (N_14773,N_9957,N_7071);
or U14774 (N_14774,N_6227,N_7409);
xnor U14775 (N_14775,N_6146,N_7053);
xor U14776 (N_14776,N_6274,N_7335);
xnor U14777 (N_14777,N_6273,N_6313);
nand U14778 (N_14778,N_6086,N_5301);
nor U14779 (N_14779,N_8905,N_7048);
or U14780 (N_14780,N_6176,N_9672);
nand U14781 (N_14781,N_7193,N_8261);
or U14782 (N_14782,N_8865,N_8077);
nand U14783 (N_14783,N_5917,N_9378);
nor U14784 (N_14784,N_5624,N_7244);
xor U14785 (N_14785,N_9807,N_8639);
and U14786 (N_14786,N_8277,N_9545);
xnor U14787 (N_14787,N_8911,N_6578);
xor U14788 (N_14788,N_8825,N_5778);
and U14789 (N_14789,N_7328,N_9653);
and U14790 (N_14790,N_9805,N_5789);
or U14791 (N_14791,N_7706,N_8790);
nor U14792 (N_14792,N_5703,N_5471);
nand U14793 (N_14793,N_9154,N_8159);
xor U14794 (N_14794,N_5418,N_8566);
and U14795 (N_14795,N_7753,N_8557);
or U14796 (N_14796,N_5962,N_9078);
nand U14797 (N_14797,N_6003,N_8614);
or U14798 (N_14798,N_5961,N_5976);
nand U14799 (N_14799,N_6628,N_5400);
nor U14800 (N_14800,N_7442,N_6333);
nand U14801 (N_14801,N_9764,N_8696);
and U14802 (N_14802,N_7314,N_6078);
nand U14803 (N_14803,N_7585,N_7475);
and U14804 (N_14804,N_8106,N_6828);
and U14805 (N_14805,N_9332,N_6265);
or U14806 (N_14806,N_7639,N_7985);
xor U14807 (N_14807,N_5277,N_7347);
xor U14808 (N_14808,N_9426,N_6591);
or U14809 (N_14809,N_5475,N_8579);
xor U14810 (N_14810,N_7573,N_8356);
or U14811 (N_14811,N_9057,N_6542);
nor U14812 (N_14812,N_5501,N_7043);
and U14813 (N_14813,N_7041,N_7297);
nor U14814 (N_14814,N_6288,N_6294);
xor U14815 (N_14815,N_9756,N_5513);
nor U14816 (N_14816,N_9640,N_9259);
nand U14817 (N_14817,N_8499,N_5630);
or U14818 (N_14818,N_5350,N_8924);
nor U14819 (N_14819,N_9836,N_6132);
nor U14820 (N_14820,N_5584,N_7620);
nand U14821 (N_14821,N_5897,N_8800);
nand U14822 (N_14822,N_8714,N_7856);
or U14823 (N_14823,N_8607,N_5657);
and U14824 (N_14824,N_5228,N_7481);
xor U14825 (N_14825,N_8508,N_5524);
and U14826 (N_14826,N_5503,N_6733);
nor U14827 (N_14827,N_7465,N_9061);
xor U14828 (N_14828,N_7982,N_7359);
or U14829 (N_14829,N_7565,N_7589);
nand U14830 (N_14830,N_8543,N_9389);
nor U14831 (N_14831,N_6644,N_5954);
or U14832 (N_14832,N_8848,N_5014);
and U14833 (N_14833,N_9678,N_6054);
xnor U14834 (N_14834,N_8277,N_7044);
or U14835 (N_14835,N_7070,N_6926);
xor U14836 (N_14836,N_7678,N_8288);
nor U14837 (N_14837,N_9707,N_8540);
xnor U14838 (N_14838,N_8695,N_6254);
and U14839 (N_14839,N_5610,N_5162);
or U14840 (N_14840,N_5500,N_8868);
and U14841 (N_14841,N_9101,N_5203);
or U14842 (N_14842,N_7405,N_5145);
nand U14843 (N_14843,N_6098,N_5032);
xor U14844 (N_14844,N_8365,N_9536);
nand U14845 (N_14845,N_8751,N_9859);
and U14846 (N_14846,N_9340,N_8506);
and U14847 (N_14847,N_8383,N_9973);
nand U14848 (N_14848,N_7711,N_9944);
nor U14849 (N_14849,N_7498,N_7370);
nor U14850 (N_14850,N_8225,N_9194);
nor U14851 (N_14851,N_7098,N_5821);
or U14852 (N_14852,N_9266,N_6907);
or U14853 (N_14853,N_9872,N_8314);
xor U14854 (N_14854,N_8405,N_5335);
nand U14855 (N_14855,N_8383,N_6841);
or U14856 (N_14856,N_8688,N_6573);
nand U14857 (N_14857,N_8528,N_6986);
nand U14858 (N_14858,N_9166,N_5722);
and U14859 (N_14859,N_7082,N_8015);
xnor U14860 (N_14860,N_5993,N_9645);
nor U14861 (N_14861,N_9394,N_5407);
and U14862 (N_14862,N_5496,N_6376);
nand U14863 (N_14863,N_6014,N_9729);
nand U14864 (N_14864,N_5071,N_6882);
and U14865 (N_14865,N_8317,N_5224);
and U14866 (N_14866,N_8006,N_8992);
xnor U14867 (N_14867,N_6333,N_8692);
or U14868 (N_14868,N_5285,N_9631);
nand U14869 (N_14869,N_8902,N_7971);
nand U14870 (N_14870,N_7042,N_5056);
nor U14871 (N_14871,N_5879,N_8998);
xnor U14872 (N_14872,N_9055,N_7598);
or U14873 (N_14873,N_7500,N_8480);
or U14874 (N_14874,N_6795,N_6885);
nand U14875 (N_14875,N_9151,N_6027);
nor U14876 (N_14876,N_6062,N_7802);
nand U14877 (N_14877,N_8163,N_9421);
nand U14878 (N_14878,N_5958,N_6128);
xor U14879 (N_14879,N_8660,N_5972);
nand U14880 (N_14880,N_9965,N_5111);
nor U14881 (N_14881,N_5057,N_5168);
nor U14882 (N_14882,N_5451,N_6866);
xnor U14883 (N_14883,N_6066,N_8194);
nor U14884 (N_14884,N_7520,N_9084);
nand U14885 (N_14885,N_9037,N_6798);
or U14886 (N_14886,N_7851,N_6565);
and U14887 (N_14887,N_6725,N_8485);
nor U14888 (N_14888,N_8963,N_6939);
or U14889 (N_14889,N_8514,N_8552);
nand U14890 (N_14890,N_5990,N_6008);
or U14891 (N_14891,N_5895,N_7957);
nor U14892 (N_14892,N_7363,N_5343);
nand U14893 (N_14893,N_8665,N_5199);
or U14894 (N_14894,N_9679,N_7947);
nor U14895 (N_14895,N_6878,N_5925);
xnor U14896 (N_14896,N_9341,N_6965);
xnor U14897 (N_14897,N_5373,N_9759);
and U14898 (N_14898,N_5850,N_5145);
nand U14899 (N_14899,N_8932,N_5776);
or U14900 (N_14900,N_6372,N_8986);
and U14901 (N_14901,N_9389,N_6994);
nor U14902 (N_14902,N_5971,N_6637);
nand U14903 (N_14903,N_6326,N_6310);
and U14904 (N_14904,N_5863,N_8940);
xor U14905 (N_14905,N_7712,N_9411);
and U14906 (N_14906,N_5701,N_7297);
xor U14907 (N_14907,N_8082,N_9886);
or U14908 (N_14908,N_5035,N_5746);
xor U14909 (N_14909,N_9158,N_6292);
and U14910 (N_14910,N_8630,N_7577);
or U14911 (N_14911,N_9046,N_8899);
or U14912 (N_14912,N_7890,N_8108);
nand U14913 (N_14913,N_7094,N_5577);
or U14914 (N_14914,N_7227,N_7888);
or U14915 (N_14915,N_9005,N_9742);
xor U14916 (N_14916,N_5251,N_8492);
or U14917 (N_14917,N_5886,N_6275);
nand U14918 (N_14918,N_6636,N_7578);
nor U14919 (N_14919,N_9448,N_5495);
nand U14920 (N_14920,N_7638,N_7068);
or U14921 (N_14921,N_9272,N_9923);
xnor U14922 (N_14922,N_9459,N_7533);
or U14923 (N_14923,N_6673,N_8077);
nor U14924 (N_14924,N_5683,N_6986);
nor U14925 (N_14925,N_6515,N_5697);
or U14926 (N_14926,N_7266,N_9737);
xor U14927 (N_14927,N_5256,N_6792);
and U14928 (N_14928,N_6619,N_6608);
or U14929 (N_14929,N_5663,N_8603);
nor U14930 (N_14930,N_6769,N_7577);
or U14931 (N_14931,N_8899,N_8668);
nand U14932 (N_14932,N_5315,N_8719);
or U14933 (N_14933,N_9773,N_7278);
or U14934 (N_14934,N_7024,N_7967);
or U14935 (N_14935,N_7963,N_8299);
or U14936 (N_14936,N_8743,N_9794);
nor U14937 (N_14937,N_8650,N_6445);
and U14938 (N_14938,N_8344,N_5421);
and U14939 (N_14939,N_6013,N_7718);
or U14940 (N_14940,N_9115,N_7557);
nand U14941 (N_14941,N_7136,N_9635);
and U14942 (N_14942,N_7709,N_7822);
or U14943 (N_14943,N_7168,N_5382);
or U14944 (N_14944,N_6141,N_8939);
nand U14945 (N_14945,N_8333,N_8788);
nand U14946 (N_14946,N_5714,N_7480);
or U14947 (N_14947,N_6053,N_9269);
nor U14948 (N_14948,N_5686,N_8325);
nor U14949 (N_14949,N_7837,N_9243);
or U14950 (N_14950,N_9049,N_7771);
nor U14951 (N_14951,N_9301,N_9344);
nand U14952 (N_14952,N_5890,N_5195);
xor U14953 (N_14953,N_8280,N_6898);
nor U14954 (N_14954,N_9816,N_5142);
xnor U14955 (N_14955,N_5426,N_5920);
xnor U14956 (N_14956,N_9598,N_6946);
or U14957 (N_14957,N_6421,N_6733);
and U14958 (N_14958,N_9986,N_9754);
nor U14959 (N_14959,N_8867,N_9568);
or U14960 (N_14960,N_5577,N_7546);
or U14961 (N_14961,N_5329,N_5463);
nand U14962 (N_14962,N_7254,N_5491);
nand U14963 (N_14963,N_6898,N_8939);
or U14964 (N_14964,N_7627,N_5678);
nand U14965 (N_14965,N_6610,N_6412);
and U14966 (N_14966,N_5029,N_5625);
nor U14967 (N_14967,N_6634,N_9561);
and U14968 (N_14968,N_6322,N_5266);
xnor U14969 (N_14969,N_7324,N_7464);
or U14970 (N_14970,N_7241,N_5036);
or U14971 (N_14971,N_6715,N_9080);
xnor U14972 (N_14972,N_6657,N_6689);
nand U14973 (N_14973,N_8338,N_5089);
nand U14974 (N_14974,N_5367,N_7132);
nor U14975 (N_14975,N_7852,N_8413);
nor U14976 (N_14976,N_8203,N_6480);
and U14977 (N_14977,N_6118,N_9230);
nor U14978 (N_14978,N_8736,N_9181);
and U14979 (N_14979,N_6915,N_5229);
and U14980 (N_14980,N_5896,N_5072);
or U14981 (N_14981,N_8923,N_8635);
and U14982 (N_14982,N_9751,N_8002);
nand U14983 (N_14983,N_7131,N_8445);
nand U14984 (N_14984,N_8972,N_6899);
and U14985 (N_14985,N_7286,N_5749);
nor U14986 (N_14986,N_5730,N_7454);
and U14987 (N_14987,N_8280,N_8606);
or U14988 (N_14988,N_9077,N_6511);
nand U14989 (N_14989,N_9272,N_6314);
nor U14990 (N_14990,N_7680,N_6745);
nor U14991 (N_14991,N_7487,N_8323);
and U14992 (N_14992,N_7048,N_5953);
or U14993 (N_14993,N_6450,N_7117);
nand U14994 (N_14994,N_7501,N_8232);
nor U14995 (N_14995,N_9077,N_6979);
nor U14996 (N_14996,N_7149,N_8958);
nor U14997 (N_14997,N_8974,N_5777);
nor U14998 (N_14998,N_7407,N_9345);
nand U14999 (N_14999,N_6093,N_6337);
nor U15000 (N_15000,N_12589,N_12524);
nand U15001 (N_15001,N_10111,N_12088);
nor U15002 (N_15002,N_10551,N_10530);
nor U15003 (N_15003,N_10554,N_10402);
and U15004 (N_15004,N_14652,N_10003);
and U15005 (N_15005,N_14844,N_11379);
or U15006 (N_15006,N_11158,N_11226);
xor U15007 (N_15007,N_13183,N_10997);
or U15008 (N_15008,N_10299,N_10694);
or U15009 (N_15009,N_13314,N_13977);
xor U15010 (N_15010,N_12207,N_14591);
nand U15011 (N_15011,N_13248,N_13493);
nor U15012 (N_15012,N_11326,N_12371);
and U15013 (N_15013,N_12213,N_14115);
nor U15014 (N_15014,N_13892,N_14690);
nor U15015 (N_15015,N_12457,N_12868);
xnor U15016 (N_15016,N_11919,N_10103);
and U15017 (N_15017,N_14354,N_10595);
or U15018 (N_15018,N_13974,N_10398);
and U15019 (N_15019,N_13007,N_12197);
or U15020 (N_15020,N_10696,N_10466);
nor U15021 (N_15021,N_11712,N_13025);
xor U15022 (N_15022,N_14696,N_14407);
nand U15023 (N_15023,N_11605,N_10698);
or U15024 (N_15024,N_11902,N_10203);
nand U15025 (N_15025,N_14944,N_13843);
nor U15026 (N_15026,N_11537,N_10913);
nand U15027 (N_15027,N_14484,N_13794);
nor U15028 (N_15028,N_13517,N_10056);
xor U15029 (N_15029,N_11133,N_14956);
nor U15030 (N_15030,N_10049,N_13366);
nor U15031 (N_15031,N_14868,N_12859);
xnor U15032 (N_15032,N_11492,N_14141);
and U15033 (N_15033,N_10993,N_10173);
nor U15034 (N_15034,N_11907,N_11152);
nor U15035 (N_15035,N_13222,N_10209);
nand U15036 (N_15036,N_11650,N_14098);
and U15037 (N_15037,N_12609,N_11238);
nor U15038 (N_15038,N_11791,N_13901);
xnor U15039 (N_15039,N_14434,N_13484);
nor U15040 (N_15040,N_14140,N_14843);
xor U15041 (N_15041,N_12908,N_11365);
nor U15042 (N_15042,N_10855,N_10545);
xor U15043 (N_15043,N_10083,N_13175);
nand U15044 (N_15044,N_12316,N_12560);
or U15045 (N_15045,N_10628,N_12607);
xnor U15046 (N_15046,N_13562,N_10377);
nand U15047 (N_15047,N_14074,N_11215);
and U15048 (N_15048,N_13301,N_14532);
or U15049 (N_15049,N_14220,N_11825);
nand U15050 (N_15050,N_14025,N_12720);
or U15051 (N_15051,N_11896,N_12285);
nor U15052 (N_15052,N_11937,N_13016);
nor U15053 (N_15053,N_10784,N_11534);
and U15054 (N_15054,N_10620,N_13757);
xnor U15055 (N_15055,N_14110,N_13940);
nor U15056 (N_15056,N_12564,N_13859);
nor U15057 (N_15057,N_12296,N_14465);
nand U15058 (N_15058,N_10290,N_13755);
nand U15059 (N_15059,N_12901,N_10124);
xnor U15060 (N_15060,N_14886,N_14488);
xnor U15061 (N_15061,N_14983,N_10890);
or U15062 (N_15062,N_12271,N_12969);
or U15063 (N_15063,N_11736,N_10077);
xnor U15064 (N_15064,N_14863,N_11583);
nand U15065 (N_15065,N_14778,N_10165);
and U15066 (N_15066,N_12604,N_12716);
xnor U15067 (N_15067,N_12391,N_11439);
nor U15068 (N_15068,N_11608,N_13272);
and U15069 (N_15069,N_12401,N_12826);
or U15070 (N_15070,N_13832,N_14460);
nand U15071 (N_15071,N_11125,N_11097);
or U15072 (N_15072,N_12225,N_12576);
nand U15073 (N_15073,N_12506,N_13996);
xor U15074 (N_15074,N_10104,N_10505);
nand U15075 (N_15075,N_12193,N_14806);
or U15076 (N_15076,N_10518,N_14125);
and U15077 (N_15077,N_11885,N_12143);
and U15078 (N_15078,N_11661,N_10683);
xor U15079 (N_15079,N_12038,N_12516);
nor U15080 (N_15080,N_12893,N_11422);
nand U15081 (N_15081,N_12542,N_10803);
xor U15082 (N_15082,N_13191,N_14749);
nand U15083 (N_15083,N_12164,N_11994);
and U15084 (N_15084,N_10725,N_12327);
nor U15085 (N_15085,N_13262,N_14583);
nor U15086 (N_15086,N_11690,N_14038);
nand U15087 (N_15087,N_13982,N_11281);
and U15088 (N_15088,N_11444,N_12109);
nor U15089 (N_15089,N_11855,N_11074);
nand U15090 (N_15090,N_11739,N_13850);
nor U15091 (N_15091,N_14709,N_12334);
nor U15092 (N_15092,N_11732,N_10719);
or U15093 (N_15093,N_14901,N_10221);
or U15094 (N_15094,N_12768,N_13657);
and U15095 (N_15095,N_12873,N_13779);
and U15096 (N_15096,N_10632,N_11665);
and U15097 (N_15097,N_12237,N_10503);
nand U15098 (N_15098,N_10019,N_13825);
and U15099 (N_15099,N_13478,N_10871);
xor U15100 (N_15100,N_10968,N_11938);
nand U15101 (N_15101,N_10831,N_10260);
xor U15102 (N_15102,N_13156,N_10668);
nor U15103 (N_15103,N_10034,N_13720);
nand U15104 (N_15104,N_10571,N_12219);
or U15105 (N_15105,N_10592,N_10043);
nor U15106 (N_15106,N_14784,N_10159);
and U15107 (N_15107,N_14129,N_11904);
xor U15108 (N_15108,N_12106,N_11785);
and U15109 (N_15109,N_14100,N_13253);
nand U15110 (N_15110,N_14547,N_11331);
nor U15111 (N_15111,N_14528,N_11005);
or U15112 (N_15112,N_10622,N_14296);
nor U15113 (N_15113,N_11059,N_12111);
xnor U15114 (N_15114,N_14351,N_14383);
and U15115 (N_15115,N_13769,N_10058);
nand U15116 (N_15116,N_14582,N_13044);
nor U15117 (N_15117,N_12120,N_13775);
xor U15118 (N_15118,N_10889,N_13090);
or U15119 (N_15119,N_10629,N_13851);
xnor U15120 (N_15120,N_11556,N_10129);
xor U15121 (N_15121,N_11272,N_13506);
nand U15122 (N_15122,N_14378,N_10869);
and U15123 (N_15123,N_11911,N_10097);
and U15124 (N_15124,N_14737,N_13275);
or U15125 (N_15125,N_14523,N_14231);
nor U15126 (N_15126,N_13030,N_13626);
nor U15127 (N_15127,N_10477,N_14720);
nand U15128 (N_15128,N_12422,N_10938);
nand U15129 (N_15129,N_12860,N_12137);
nor U15130 (N_15130,N_14119,N_13322);
nor U15131 (N_15131,N_13316,N_14040);
or U15132 (N_15132,N_14243,N_12572);
or U15133 (N_15133,N_10788,N_10712);
nor U15134 (N_15134,N_13710,N_13689);
nor U15135 (N_15135,N_11871,N_14406);
or U15136 (N_15136,N_14469,N_11597);
and U15137 (N_15137,N_12466,N_11347);
xor U15138 (N_15138,N_11166,N_13283);
nand U15139 (N_15139,N_11830,N_10279);
xor U15140 (N_15140,N_10678,N_14173);
nor U15141 (N_15141,N_10186,N_10036);
or U15142 (N_15142,N_10969,N_14062);
nand U15143 (N_15143,N_13210,N_11063);
nor U15144 (N_15144,N_14021,N_11763);
nor U15145 (N_15145,N_10846,N_14216);
xnor U15146 (N_15146,N_13497,N_13541);
or U15147 (N_15147,N_10047,N_14888);
nand U15148 (N_15148,N_14486,N_12640);
and U15149 (N_15149,N_11689,N_12973);
and U15150 (N_15150,N_14933,N_11749);
nor U15151 (N_15151,N_10114,N_13266);
or U15152 (N_15152,N_12886,N_12956);
nor U15153 (N_15153,N_13670,N_12698);
and U15154 (N_15154,N_13797,N_11124);
and U15155 (N_15155,N_12399,N_12658);
nor U15156 (N_15156,N_12686,N_13966);
nand U15157 (N_15157,N_11956,N_12739);
nor U15158 (N_15158,N_12963,N_13711);
nor U15159 (N_15159,N_13535,N_11382);
xor U15160 (N_15160,N_12622,N_10387);
nor U15161 (N_15161,N_13043,N_10747);
xor U15162 (N_15162,N_13856,N_11046);
xnor U15163 (N_15163,N_10858,N_13189);
and U15164 (N_15164,N_10705,N_10736);
nor U15165 (N_15165,N_14360,N_10270);
xor U15166 (N_15166,N_10359,N_12481);
or U15167 (N_15167,N_12508,N_13992);
nor U15168 (N_15168,N_13129,N_11566);
or U15169 (N_15169,N_12728,N_14197);
and U15170 (N_15170,N_14050,N_10222);
xnor U15171 (N_15171,N_14157,N_14626);
and U15172 (N_15172,N_13629,N_14028);
xnor U15173 (N_15173,N_13390,N_14345);
or U15174 (N_15174,N_10676,N_14061);
or U15175 (N_15175,N_10364,N_11954);
and U15176 (N_15176,N_12014,N_12488);
nand U15177 (N_15177,N_10610,N_14938);
or U15178 (N_15178,N_10671,N_13865);
and U15179 (N_15179,N_13807,N_13782);
xor U15180 (N_15180,N_10125,N_13527);
or U15181 (N_15181,N_10147,N_12676);
nand U15182 (N_15182,N_12256,N_11231);
xor U15183 (N_15183,N_14271,N_13231);
or U15184 (N_15184,N_13987,N_11115);
nand U15185 (N_15185,N_13890,N_14907);
nor U15186 (N_15186,N_14043,N_11880);
nor U15187 (N_15187,N_14550,N_13834);
or U15188 (N_15188,N_11768,N_11870);
nor U15189 (N_15189,N_12212,N_10010);
and U15190 (N_15190,N_12816,N_14819);
or U15191 (N_15191,N_10985,N_10630);
or U15192 (N_15192,N_14879,N_10488);
and U15193 (N_15193,N_11606,N_11789);
xnor U15194 (N_15194,N_12112,N_12030);
xor U15195 (N_15195,N_14909,N_12865);
xnor U15196 (N_15196,N_14000,N_11582);
xor U15197 (N_15197,N_11230,N_11245);
nand U15198 (N_15198,N_10236,N_10272);
nand U15199 (N_15199,N_11104,N_11864);
nor U15200 (N_15200,N_14498,N_12458);
or U15201 (N_15201,N_12100,N_13830);
or U15202 (N_15202,N_14796,N_12923);
nor U15203 (N_15203,N_14916,N_10623);
and U15204 (N_15204,N_12389,N_13200);
xnor U15205 (N_15205,N_12898,N_14587);
or U15206 (N_15206,N_10394,N_11729);
xnor U15207 (N_15207,N_12682,N_14116);
xnor U15208 (N_15208,N_13296,N_12707);
or U15209 (N_15209,N_14966,N_13544);
nand U15210 (N_15210,N_11834,N_13192);
nor U15211 (N_15211,N_14272,N_14153);
nand U15212 (N_15212,N_11519,N_11394);
and U15213 (N_15213,N_13298,N_14152);
and U15214 (N_15214,N_10506,N_11558);
xnor U15215 (N_15215,N_12402,N_12862);
and U15216 (N_15216,N_12058,N_14945);
xnor U15217 (N_15217,N_11531,N_12210);
nand U15218 (N_15218,N_14836,N_11090);
or U15219 (N_15219,N_10136,N_14396);
nor U15220 (N_15220,N_12759,N_13781);
or U15221 (N_15221,N_12804,N_12001);
nor U15222 (N_15222,N_14769,N_10312);
nand U15223 (N_15223,N_13078,N_14385);
and U15224 (N_15224,N_12734,N_10142);
and U15225 (N_15225,N_10230,N_12730);
nor U15226 (N_15226,N_14952,N_10320);
and U15227 (N_15227,N_12735,N_13023);
or U15228 (N_15228,N_11053,N_14555);
nand U15229 (N_15229,N_12671,N_12127);
nor U15230 (N_15230,N_14177,N_13060);
nand U15231 (N_15231,N_12861,N_12061);
or U15232 (N_15232,N_10662,N_13736);
xnor U15233 (N_15233,N_10112,N_10025);
nand U15234 (N_15234,N_10562,N_11214);
xor U15235 (N_15235,N_10957,N_10489);
nand U15236 (N_15236,N_11021,N_10762);
or U15237 (N_15237,N_13798,N_13516);
xnor U15238 (N_15238,N_13494,N_12568);
nand U15239 (N_15239,N_12055,N_10565);
or U15240 (N_15240,N_10075,N_12944);
or U15241 (N_15241,N_11551,N_13328);
and U15242 (N_15242,N_12927,N_13767);
nand U15243 (N_15243,N_13473,N_12298);
and U15244 (N_15244,N_10037,N_13559);
xor U15245 (N_15245,N_14618,N_10318);
and U15246 (N_15246,N_14592,N_12043);
and U15247 (N_15247,N_14978,N_12342);
and U15248 (N_15248,N_13435,N_12113);
nor U15249 (N_15249,N_13162,N_11332);
nor U15250 (N_15250,N_13219,N_10130);
nor U15251 (N_15251,N_14093,N_10443);
nand U15252 (N_15252,N_12179,N_13127);
xor U15253 (N_15253,N_14448,N_14715);
or U15254 (N_15254,N_12477,N_14973);
nor U15255 (N_15255,N_12654,N_14756);
nand U15256 (N_15256,N_13028,N_12482);
and U15257 (N_15257,N_10117,N_10816);
or U15258 (N_15258,N_13905,N_11888);
nor U15259 (N_15259,N_11643,N_12957);
nand U15260 (N_15260,N_14067,N_11378);
nor U15261 (N_15261,N_12544,N_14828);
or U15262 (N_15262,N_10432,N_14455);
nand U15263 (N_15263,N_14075,N_14232);
xor U15264 (N_15264,N_13004,N_12585);
xor U15265 (N_15265,N_11777,N_13876);
xor U15266 (N_15266,N_11620,N_12417);
and U15267 (N_15267,N_12273,N_13914);
xor U15268 (N_15268,N_10746,N_11488);
nand U15269 (N_15269,N_13627,N_14492);
nor U15270 (N_15270,N_14946,N_11111);
or U15271 (N_15271,N_10480,N_11547);
and U15272 (N_15272,N_13730,N_12383);
nand U15273 (N_15273,N_13533,N_14403);
nor U15274 (N_15274,N_13228,N_13567);
nand U15275 (N_15275,N_13079,N_12530);
nand U15276 (N_15276,N_12400,N_14188);
or U15277 (N_15277,N_11452,N_13102);
nor U15278 (N_15278,N_12360,N_11892);
nor U15279 (N_15279,N_11928,N_11939);
nor U15280 (N_15280,N_10135,N_10431);
nor U15281 (N_15281,N_14953,N_12577);
or U15282 (N_15282,N_14341,N_11812);
and U15283 (N_15283,N_10338,N_11336);
nand U15284 (N_15284,N_10315,N_11664);
nor U15285 (N_15285,N_13835,N_14068);
and U15286 (N_15286,N_13001,N_10153);
and U15287 (N_15287,N_12307,N_11100);
and U15288 (N_15288,N_13695,N_14304);
xor U15289 (N_15289,N_14285,N_11048);
xor U15290 (N_15290,N_10637,N_10041);
xor U15291 (N_15291,N_11499,N_10617);
and U15292 (N_15292,N_11634,N_13218);
or U15293 (N_15293,N_10335,N_14728);
or U15294 (N_15294,N_10640,N_12373);
nand U15295 (N_15295,N_13572,N_11248);
and U15296 (N_15296,N_10681,N_11150);
nor U15297 (N_15297,N_13561,N_11039);
nor U15298 (N_15298,N_12000,N_14979);
or U15299 (N_15299,N_12117,N_13667);
or U15300 (N_15300,N_12292,N_12461);
nand U15301 (N_15301,N_13161,N_10649);
and U15302 (N_15302,N_10673,N_13613);
xnor U15303 (N_15303,N_12738,N_14390);
and U15304 (N_15304,N_11972,N_11656);
and U15305 (N_15305,N_11561,N_13457);
and U15306 (N_15306,N_11599,N_13003);
nor U15307 (N_15307,N_11254,N_10675);
xor U15308 (N_15308,N_10799,N_13615);
nor U15309 (N_15309,N_14792,N_11208);
nor U15310 (N_15310,N_14072,N_14073);
or U15311 (N_15311,N_12810,N_12136);
and U15312 (N_15312,N_13868,N_13197);
or U15313 (N_15313,N_14384,N_14156);
or U15314 (N_15314,N_10152,N_13915);
xnor U15315 (N_15315,N_12900,N_14568);
nor U15316 (N_15316,N_10040,N_13594);
xor U15317 (N_15317,N_12470,N_10511);
nor U15318 (N_15318,N_14107,N_13837);
or U15319 (N_15319,N_10928,N_13240);
xor U15320 (N_15320,N_13976,N_10996);
xnor U15321 (N_15321,N_13566,N_10175);
and U15322 (N_15322,N_10192,N_10689);
nor U15323 (N_15323,N_11700,N_10949);
nand U15324 (N_15324,N_13076,N_13988);
nor U15325 (N_15325,N_10426,N_13554);
nand U15326 (N_15326,N_10252,N_12044);
or U15327 (N_15327,N_13088,N_11621);
and U15328 (N_15328,N_10569,N_13871);
or U15329 (N_15329,N_10907,N_10864);
nand U15330 (N_15330,N_11589,N_14866);
xor U15331 (N_15331,N_13729,N_10851);
or U15332 (N_15332,N_14027,N_13768);
xor U15333 (N_15333,N_13522,N_10718);
xor U15334 (N_15334,N_12982,N_10524);
and U15335 (N_15335,N_11970,N_14112);
nand U15336 (N_15336,N_13867,N_14142);
nand U15337 (N_15337,N_12964,N_10570);
nor U15338 (N_15338,N_10919,N_11814);
xnor U15339 (N_15339,N_13268,N_14770);
or U15340 (N_15340,N_11741,N_13848);
nor U15341 (N_15341,N_12758,N_11542);
xor U15342 (N_15342,N_12536,N_11623);
and U15343 (N_15343,N_13972,N_13679);
nand U15344 (N_15344,N_10709,N_10614);
or U15345 (N_15345,N_14544,N_11300);
and U15346 (N_15346,N_12131,N_14309);
and U15347 (N_15347,N_11529,N_10661);
and U15348 (N_15348,N_10391,N_14343);
nor U15349 (N_15349,N_12523,N_11258);
nand U15350 (N_15350,N_11188,N_14848);
nor U15351 (N_15351,N_12526,N_11734);
and U15352 (N_15352,N_13120,N_10115);
xor U15353 (N_15353,N_11957,N_12016);
and U15354 (N_15354,N_10943,N_11831);
nor U15355 (N_15355,N_14619,N_14194);
xor U15356 (N_15356,N_11895,N_11550);
and U15357 (N_15357,N_10193,N_14942);
nor U15358 (N_15358,N_13326,N_14624);
and U15359 (N_15359,N_11363,N_10361);
nor U15360 (N_15360,N_14039,N_11651);
or U15361 (N_15361,N_14521,N_12166);
nand U15362 (N_15362,N_13654,N_11387);
nand U15363 (N_15363,N_14706,N_13292);
nor U15364 (N_15364,N_11602,N_13748);
and U15365 (N_15365,N_14765,N_14847);
xnor U15366 (N_15366,N_13303,N_13889);
nor U15367 (N_15367,N_10925,N_10801);
nor U15368 (N_15368,N_13121,N_12007);
xnor U15369 (N_15369,N_12541,N_12772);
nand U15370 (N_15370,N_14563,N_12918);
nor U15371 (N_15371,N_13181,N_13059);
nand U15372 (N_15372,N_13587,N_14411);
and U15373 (N_15373,N_12569,N_11278);
or U15374 (N_15374,N_11515,N_14999);
or U15375 (N_15375,N_11816,N_10714);
nand U15376 (N_15376,N_14052,N_13632);
nand U15377 (N_15377,N_14215,N_12203);
xor U15378 (N_15378,N_14059,N_12566);
nand U15379 (N_15379,N_13605,N_11813);
or U15380 (N_15380,N_13735,N_10150);
or U15381 (N_15381,N_11370,N_14036);
and U15382 (N_15382,N_14421,N_10206);
xnor U15383 (N_15383,N_13857,N_12076);
xnor U15384 (N_15384,N_11506,N_11434);
and U15385 (N_15385,N_12657,N_14258);
xor U15386 (N_15386,N_10806,N_12895);
nor U15387 (N_15387,N_10885,N_10383);
or U15388 (N_15388,N_12156,N_14695);
and U15389 (N_15389,N_14372,N_11503);
nand U15390 (N_15390,N_13575,N_13339);
nand U15391 (N_15391,N_13368,N_11291);
nand U15392 (N_15392,N_13531,N_14841);
xor U15393 (N_15393,N_11032,N_13250);
and U15394 (N_15394,N_11316,N_13928);
xnor U15395 (N_15395,N_13937,N_11947);
xor U15396 (N_15396,N_14562,N_12983);
nand U15397 (N_15397,N_13655,N_14008);
nand U15398 (N_15398,N_14604,N_11004);
or U15399 (N_15399,N_13873,N_13713);
xnor U15400 (N_15400,N_10319,N_10261);
nand U15401 (N_15401,N_13367,N_11836);
nor U15402 (N_15402,N_13944,N_11731);
or U15403 (N_15403,N_14698,N_10128);
and U15404 (N_15404,N_10340,N_14884);
nand U15405 (N_15405,N_10693,N_11696);
nand U15406 (N_15406,N_13583,N_12601);
and U15407 (N_15407,N_10903,N_13789);
nor U15408 (N_15408,N_10009,N_10909);
or U15409 (N_15409,N_12811,N_10734);
and U15410 (N_15410,N_14430,N_14374);
and U15411 (N_15411,N_11415,N_10374);
nor U15412 (N_15412,N_14234,N_13696);
xnor U15413 (N_15413,N_13415,N_12934);
and U15414 (N_15414,N_11701,N_10048);
and U15415 (N_15415,N_14323,N_13285);
xor U15416 (N_15416,N_12899,N_11116);
nor U15417 (N_15417,N_11507,N_12801);
nand U15418 (N_15418,N_14009,N_11356);
or U15419 (N_15419,N_12659,N_13681);
nor U15420 (N_15420,N_11820,N_11019);
or U15421 (N_15421,N_12891,N_13190);
or U15422 (N_15422,N_11174,N_13866);
or U15423 (N_15423,N_12303,N_14511);
nor U15424 (N_15424,N_12040,N_13440);
and U15425 (N_15425,N_14809,N_11835);
or U15426 (N_15426,N_14889,N_14837);
nor U15427 (N_15427,N_10962,N_10959);
and U15428 (N_15428,N_12069,N_10633);
nor U15429 (N_15429,N_14615,N_10292);
and U15430 (N_15430,N_10350,N_10183);
xor U15431 (N_15431,N_13780,N_14755);
nand U15432 (N_15432,N_12093,N_14635);
nand U15433 (N_15433,N_14569,N_11203);
xnor U15434 (N_15434,N_11112,N_10830);
nor U15435 (N_15435,N_10763,N_12062);
or U15436 (N_15436,N_12504,N_13331);
nor U15437 (N_15437,N_14005,N_12883);
nor U15438 (N_15438,N_11709,N_14481);
or U15439 (N_15439,N_13749,N_11129);
or U15440 (N_15440,N_13180,N_11107);
and U15441 (N_15441,N_11012,N_13194);
and U15442 (N_15442,N_13092,N_12719);
nor U15443 (N_15443,N_12475,N_11960);
or U15444 (N_15444,N_12190,N_14510);
or U15445 (N_15445,N_10857,N_10686);
nand U15446 (N_15446,N_14661,N_13501);
or U15447 (N_15447,N_14517,N_10370);
or U15448 (N_15448,N_11857,N_13365);
xnor U15449 (N_15449,N_14244,N_13433);
and U15450 (N_15450,N_10081,N_12940);
nand U15451 (N_15451,N_10815,N_10706);
nor U15452 (N_15452,N_11171,N_12755);
or U15453 (N_15453,N_11965,N_13448);
or U15454 (N_15454,N_14601,N_13113);
nand U15455 (N_15455,N_10579,N_10464);
nor U15456 (N_15456,N_13542,N_12362);
xnor U15457 (N_15457,N_13416,N_10276);
nor U15458 (N_15458,N_14949,N_13659);
or U15459 (N_15459,N_14239,N_14146);
nand U15460 (N_15460,N_11799,N_13578);
and U15461 (N_15461,N_13754,N_10005);
xnor U15462 (N_15462,N_12877,N_12588);
or U15463 (N_15463,N_11458,N_14801);
and U15464 (N_15464,N_10544,N_12777);
nand U15465 (N_15465,N_12280,N_11851);
xor U15466 (N_15466,N_12896,N_14717);
nand U15467 (N_15467,N_10158,N_12794);
or U15468 (N_15468,N_11873,N_11156);
nand U15469 (N_15469,N_11983,N_11553);
or U15470 (N_15470,N_10311,N_12757);
nand U15471 (N_15471,N_11724,N_10491);
nand U15472 (N_15472,N_10866,N_11819);
xnor U15473 (N_15473,N_10650,N_13978);
or U15474 (N_15474,N_12003,N_14369);
and U15475 (N_15475,N_14085,N_14988);
nor U15476 (N_15476,N_10022,N_14995);
nand U15477 (N_15477,N_11290,N_14890);
or U15478 (N_15478,N_11635,N_11809);
xor U15479 (N_15479,N_11775,N_11630);
nor U15480 (N_15480,N_13177,N_10704);
nand U15481 (N_15481,N_14402,N_12775);
nor U15482 (N_15482,N_10844,N_13128);
nand U15483 (N_15483,N_10467,N_13833);
nand U15484 (N_15484,N_11838,N_11437);
or U15485 (N_15485,N_13662,N_14376);
nand U15486 (N_15486,N_10860,N_10468);
nand U15487 (N_15487,N_10283,N_13690);
and U15488 (N_15488,N_13293,N_11270);
nand U15489 (N_15489,N_10429,N_11334);
and U15490 (N_15490,N_12502,N_12115);
xor U15491 (N_15491,N_12835,N_11009);
nor U15492 (N_15492,N_10828,N_13716);
and U15493 (N_15493,N_10669,N_14287);
and U15494 (N_15494,N_13875,N_13214);
or U15495 (N_15495,N_14162,N_13481);
nor U15496 (N_15496,N_13510,N_10358);
xnor U15497 (N_15497,N_11277,N_11592);
and U15498 (N_15498,N_14795,N_13595);
nand U15499 (N_15499,N_11793,N_14353);
nor U15500 (N_15500,N_13953,N_12008);
nand U15501 (N_15501,N_12539,N_14094);
nor U15502 (N_15502,N_14464,N_11669);
or U15503 (N_15503,N_10099,N_10098);
nor U15504 (N_15504,N_10007,N_14219);
nor U15505 (N_15505,N_12699,N_13348);
xor U15506 (N_15506,N_10791,N_14284);
xnor U15507 (N_15507,N_14876,N_11041);
and U15508 (N_15508,N_12315,N_11253);
or U15509 (N_15509,N_12178,N_10018);
nand U15510 (N_15510,N_10872,N_11184);
nor U15511 (N_15511,N_10819,N_14947);
xor U15512 (N_15512,N_14738,N_13340);
nor U15513 (N_15513,N_12513,N_13089);
or U15514 (N_15514,N_14803,N_10499);
and U15515 (N_15515,N_14056,N_10137);
xnor U15516 (N_15516,N_11189,N_12805);
nand U15517 (N_15517,N_10045,N_14893);
nor U15518 (N_15518,N_11521,N_11475);
xor U15519 (N_15519,N_10249,N_13269);
xnor U15520 (N_15520,N_11884,N_12462);
xnor U15521 (N_15521,N_11134,N_12533);
xnor U15522 (N_15522,N_12145,N_13722);
or U15523 (N_15523,N_14468,N_12472);
nand U15524 (N_15524,N_13279,N_13565);
or U15525 (N_15525,N_14589,N_10039);
nor U15526 (N_15526,N_14810,N_11343);
nor U15527 (N_15527,N_14920,N_11038);
nand U15528 (N_15528,N_13377,N_14887);
nor U15529 (N_15529,N_13235,N_11850);
and U15530 (N_15530,N_11017,N_10105);
and U15531 (N_15531,N_10741,N_14035);
xor U15532 (N_15532,N_11935,N_10707);
and U15533 (N_15533,N_11246,N_13199);
xnor U15534 (N_15534,N_12253,N_14404);
nand U15535 (N_15535,N_11752,N_12455);
nand U15536 (N_15536,N_12988,N_13398);
nor U15537 (N_15537,N_14501,N_10541);
xnor U15538 (N_15538,N_11874,N_10224);
xor U15539 (N_15539,N_14996,N_10684);
nor U15540 (N_15540,N_13631,N_12184);
and U15541 (N_15541,N_11671,N_12435);
nor U15542 (N_15542,N_13135,N_14969);
xnor U15543 (N_15543,N_13518,N_12929);
nand U15544 (N_15544,N_12252,N_10014);
nand U15545 (N_15545,N_14856,N_11425);
xor U15546 (N_15546,N_12428,N_11843);
xnor U15547 (N_15547,N_10455,N_11192);
or U15548 (N_15548,N_13139,N_12224);
nor U15549 (N_15549,N_12871,N_11468);
nor U15550 (N_15550,N_13008,N_10867);
xnor U15551 (N_15551,N_10345,N_11395);
and U15552 (N_15552,N_13421,N_10893);
and U15553 (N_15553,N_10325,N_13664);
or U15554 (N_15554,N_14700,N_12217);
xor U15555 (N_15555,N_12855,N_14721);
xor U15556 (N_15556,N_10134,N_12104);
or U15557 (N_15557,N_11249,N_11504);
xnor U15558 (N_15558,N_10008,N_10231);
nand U15559 (N_15559,N_13342,N_11501);
nor U15560 (N_15560,N_12932,N_11427);
xnor U15561 (N_15561,N_13418,N_13480);
nand U15562 (N_15562,N_10409,N_12912);
or U15563 (N_15563,N_14977,N_12884);
xnor U15564 (N_15564,N_12602,N_12495);
nor U15565 (N_15565,N_10643,N_11497);
and U15566 (N_15566,N_10289,N_10028);
nor U15567 (N_15567,N_14045,N_12836);
or U15568 (N_15568,N_11526,N_13459);
and U15569 (N_15569,N_13141,N_12047);
or U15570 (N_15570,N_11966,N_13136);
and U15571 (N_15571,N_13727,N_11196);
xor U15572 (N_15572,N_14497,N_13759);
and U15573 (N_15573,N_14833,N_14476);
and U15574 (N_15574,N_13529,N_10138);
nor U15575 (N_15575,N_11193,N_14334);
xor U15576 (N_15576,N_12753,N_13840);
xor U15577 (N_15577,N_12765,N_12424);
nand U15578 (N_15578,N_12460,N_14646);
nor U15579 (N_15579,N_13762,N_13788);
and U15580 (N_15580,N_11847,N_12736);
nor U15581 (N_15581,N_12072,N_12991);
or U15582 (N_15582,N_10106,N_13683);
xor U15583 (N_15583,N_13855,N_12555);
and U15584 (N_15584,N_14377,N_10948);
nor U15585 (N_15585,N_14266,N_14041);
xnor U15586 (N_15586,N_11137,N_10448);
and U15587 (N_15587,N_13171,N_10862);
nor U15588 (N_15588,N_11996,N_12625);
xnor U15589 (N_15589,N_13563,N_11241);
xnor U15590 (N_15590,N_13942,N_13795);
nor U15591 (N_15591,N_11323,N_13827);
xnor U15592 (N_15592,N_11461,N_12845);
nor U15593 (N_15593,N_13744,N_10642);
and U15594 (N_15594,N_10133,N_13699);
nand U15595 (N_15595,N_14222,N_12480);
nand U15596 (N_15596,N_11182,N_13732);
and U15597 (N_15597,N_12254,N_11298);
xor U15598 (N_15598,N_13052,N_14829);
nand U15599 (N_15599,N_11841,N_11743);
nand U15600 (N_15600,N_13617,N_10110);
nor U15601 (N_15601,N_10991,N_13081);
nor U15602 (N_15602,N_14237,N_12797);
xor U15603 (N_15603,N_11217,N_12170);
xnor U15604 (N_15604,N_12238,N_13980);
or U15605 (N_15605,N_10755,N_12086);
and U15606 (N_15606,N_13085,N_11595);
xor U15607 (N_15607,N_11436,N_13665);
nor U15608 (N_15608,N_13356,N_12974);
nand U15609 (N_15609,N_13256,N_11933);
or U15610 (N_15610,N_14462,N_14734);
nand U15611 (N_15611,N_14785,N_12194);
xor U15612 (N_15612,N_12525,N_11273);
nand U15613 (N_15613,N_12453,N_13954);
xnor U15614 (N_15614,N_14854,N_10168);
and U15615 (N_15615,N_11200,N_12750);
or U15616 (N_15616,N_12665,N_10092);
and U15617 (N_15617,N_10328,N_12168);
and U15618 (N_15618,N_10140,N_14250);
nor U15619 (N_15619,N_11518,N_14775);
nand U15620 (N_15620,N_14816,N_12540);
or U15621 (N_15621,N_13046,N_12711);
nand U15622 (N_15622,N_11968,N_10685);
or U15623 (N_15623,N_12331,N_10457);
xnor U15624 (N_15624,N_11910,N_14263);
or U15625 (N_15625,N_14598,N_12856);
xnor U15626 (N_15626,N_11473,N_14166);
or U15627 (N_15627,N_10566,N_14559);
xor U15628 (N_15628,N_13343,N_11072);
xnor U15629 (N_15629,N_11029,N_14827);
xnor U15630 (N_15630,N_10636,N_13329);
or U15631 (N_15631,N_10266,N_11146);
or U15632 (N_15632,N_13639,N_12591);
xor U15633 (N_15633,N_12205,N_13860);
xnor U15634 (N_15634,N_12187,N_13006);
nand U15635 (N_15635,N_11990,N_12656);
nor U15636 (N_15636,N_14182,N_12330);
and U15637 (N_15637,N_10062,N_10465);
nand U15638 (N_15638,N_12059,N_13887);
and U15639 (N_15639,N_13579,N_13226);
xor U15640 (N_15640,N_13929,N_13178);
nand U15641 (N_15641,N_14034,N_11546);
nor U15642 (N_15642,N_12632,N_13813);
or U15643 (N_15643,N_14480,N_13187);
xnor U15644 (N_15644,N_12563,N_13149);
or U15645 (N_15645,N_11969,N_14633);
nor U15646 (N_15646,N_12595,N_11126);
and U15647 (N_15647,N_12384,N_14923);
nand U15648 (N_15648,N_10768,N_13599);
and U15649 (N_15649,N_11554,N_13100);
and U15650 (N_15650,N_11037,N_13492);
or U15651 (N_15651,N_11413,N_11209);
or U15652 (N_15652,N_14208,N_11711);
xnor U15653 (N_15653,N_11716,N_13360);
xnor U15654 (N_15654,N_12629,N_13157);
or U15655 (N_15655,N_13051,N_12894);
xnor U15656 (N_15656,N_10013,N_10939);
nand U15657 (N_15657,N_13108,N_10548);
or U15658 (N_15658,N_10744,N_12198);
and U15659 (N_15659,N_13521,N_13400);
nand U15660 (N_15660,N_10156,N_13734);
nor U15661 (N_15661,N_11920,N_12905);
xnor U15662 (N_15662,N_10581,N_12911);
and U15663 (N_15663,N_14984,N_12505);
xnor U15664 (N_15664,N_14001,N_14066);
xnor U15665 (N_15665,N_10563,N_14415);
xnor U15666 (N_15666,N_12163,N_10456);
nand U15667 (N_15667,N_12837,N_10501);
xor U15668 (N_15668,N_14688,N_11084);
and U15669 (N_15669,N_13962,N_13756);
nor U15670 (N_15670,N_14181,N_10875);
xnor U15671 (N_15671,N_12438,N_10386);
nand U15672 (N_15672,N_10244,N_12653);
xnor U15673 (N_15673,N_12840,N_14623);
xnor U15674 (N_15674,N_12608,N_13406);
nor U15675 (N_15675,N_13345,N_11806);
or U15676 (N_15676,N_14622,N_13959);
or U15677 (N_15677,N_14982,N_11201);
and U15678 (N_15678,N_10888,N_14880);
and U15679 (N_15679,N_11367,N_11697);
or U15680 (N_15680,N_11802,N_13381);
xor U15681 (N_15681,N_13054,N_14303);
nor U15682 (N_15682,N_11893,N_11760);
or U15683 (N_15683,N_13574,N_14726);
or U15684 (N_15684,N_12534,N_11527);
xor U15685 (N_15685,N_12729,N_11438);
xor U15686 (N_15686,N_10327,N_14588);
nor U15687 (N_15687,N_14405,N_12718);
xor U15688 (N_15688,N_14963,N_12531);
nor U15689 (N_15689,N_14813,N_11068);
xnor U15690 (N_15690,N_14233,N_12301);
xor U15691 (N_15691,N_12761,N_10415);
or U15692 (N_15692,N_12175,N_10458);
xor U15693 (N_15693,N_13387,N_13885);
nand U15694 (N_15694,N_13142,N_13464);
and U15695 (N_15695,N_14147,N_14518);
xnor U15696 (N_15696,N_13511,N_14307);
nand U15697 (N_15697,N_11381,N_14409);
xor U15698 (N_15698,N_13792,N_12537);
or U15699 (N_15699,N_11329,N_10892);
and U15700 (N_15700,N_11110,N_11748);
nand U15701 (N_15701,N_12955,N_12839);
and U15702 (N_15702,N_13998,N_12514);
or U15703 (N_15703,N_10776,N_12597);
and U15704 (N_15704,N_14579,N_11432);
nand U15705 (N_15705,N_14449,N_12611);
nand U15706 (N_15706,N_13082,N_10742);
nor U15707 (N_15707,N_14644,N_12245);
nor U15708 (N_15708,N_10724,N_14851);
or U15709 (N_15709,N_14500,N_12049);
nand U15710 (N_15710,N_14329,N_11243);
or U15711 (N_15711,N_12732,N_10608);
and U15712 (N_15712,N_13697,N_11860);
nor U15713 (N_15713,N_10601,N_14097);
and U15714 (N_15714,N_14295,N_13297);
xor U15715 (N_15715,N_14349,N_10988);
and U15716 (N_15716,N_12812,N_13422);
xnor U15717 (N_15717,N_11462,N_12990);
and U15718 (N_15718,N_14331,N_13682);
xor U15719 (N_15719,N_12078,N_13383);
nor U15720 (N_15720,N_13853,N_10421);
nand U15721 (N_15721,N_11699,N_14613);
nor U15722 (N_15722,N_12954,N_10513);
xor U15723 (N_15723,N_13165,N_12666);
or U15724 (N_15724,N_14252,N_10779);
and U15725 (N_15725,N_12798,N_13224);
and U15726 (N_15726,N_14132,N_12249);
and U15727 (N_15727,N_14727,N_13470);
or U15728 (N_15728,N_10583,N_10641);
xor U15729 (N_15729,N_12571,N_13881);
and U15730 (N_15730,N_13965,N_14595);
nor U15731 (N_15731,N_11626,N_14748);
xor U15732 (N_15732,N_12689,N_12624);
or U15733 (N_15733,N_11878,N_11001);
nand U15734 (N_15734,N_11216,N_14505);
and U15735 (N_15735,N_14545,N_10486);
and U15736 (N_15736,N_14750,N_13960);
and U15737 (N_15737,N_10580,N_10657);
nand U15738 (N_15738,N_11817,N_14362);
nor U15739 (N_15739,N_13894,N_13245);
nor U15740 (N_15740,N_14418,N_10248);
xor U15741 (N_15741,N_10323,N_11829);
or U15742 (N_15742,N_12419,N_14096);
nand U15743 (N_15743,N_11538,N_11311);
nor U15744 (N_15744,N_12414,N_12356);
and U15745 (N_15745,N_10995,N_12680);
nor U15746 (N_15746,N_11549,N_14026);
xor U15747 (N_15747,N_12227,N_12806);
and U15748 (N_15748,N_10635,N_10805);
or U15749 (N_15749,N_13252,N_14143);
and U15750 (N_15750,N_12107,N_14226);
nor U15751 (N_15751,N_13230,N_11989);
nand U15752 (N_15752,N_11536,N_10258);
nand U15753 (N_15753,N_12297,N_10543);
and U15754 (N_15754,N_14433,N_14735);
xnor U15755 (N_15755,N_14541,N_11149);
nand U15756 (N_15756,N_10838,N_14692);
xor U15757 (N_15757,N_10896,N_10802);
xor U15758 (N_15758,N_11915,N_14669);
nor U15759 (N_15759,N_13118,N_11510);
or U15760 (N_15760,N_14210,N_10473);
xor U15761 (N_15761,N_14145,N_12679);
and U15762 (N_15762,N_10030,N_12188);
xnor U15763 (N_15763,N_14007,N_11143);
and U15764 (N_15764,N_13761,N_12870);
nand U15765 (N_15765,N_10564,N_13673);
or U15766 (N_15766,N_14761,N_10979);
nor U15767 (N_15767,N_13163,N_10647);
xnor U15768 (N_15768,N_13126,N_11639);
nand U15769 (N_15769,N_13515,N_14131);
or U15770 (N_15770,N_11096,N_14594);
or U15771 (N_15771,N_12485,N_10476);
nand U15772 (N_15772,N_13741,N_11346);
and U15773 (N_15773,N_10061,N_14857);
and U15774 (N_15774,N_12353,N_11694);
nand U15775 (N_15775,N_11980,N_10381);
and U15776 (N_15776,N_10773,N_11198);
nor U15777 (N_15777,N_12950,N_11377);
xor U15778 (N_15778,N_10535,N_12028);
nor U15779 (N_15779,N_10257,N_14292);
nor U15780 (N_15780,N_10652,N_10870);
or U15781 (N_15781,N_13454,N_10121);
and U15782 (N_15782,N_12325,N_10035);
nor U15783 (N_15783,N_14060,N_11926);
or U15784 (N_15784,N_12468,N_11640);
or U15785 (N_15785,N_13712,N_10575);
nand U15786 (N_15786,N_14612,N_11991);
xor U15787 (N_15787,N_11454,N_11511);
and U15788 (N_15788,N_11351,N_12029);
and U15789 (N_15789,N_10384,N_12103);
or U15790 (N_15790,N_10677,N_14205);
xor U15791 (N_15791,N_10895,N_11315);
or U15792 (N_15792,N_14954,N_10001);
or U15793 (N_15793,N_11355,N_11839);
nand U15794 (N_15794,N_11257,N_11087);
nor U15795 (N_15795,N_14919,N_14903);
xor U15796 (N_15796,N_14175,N_13476);
or U15797 (N_15797,N_12489,N_12764);
nand U15798 (N_15798,N_13642,N_13396);
or U15799 (N_15799,N_14912,N_14425);
nor U15800 (N_15800,N_12299,N_14660);
and U15801 (N_15801,N_10967,N_13705);
and U15802 (N_15802,N_11963,N_11707);
or U15803 (N_15803,N_11051,N_12878);
nand U15804 (N_15804,N_10445,N_14054);
or U15805 (N_15805,N_13074,N_14990);
xor U15806 (N_15806,N_10309,N_14014);
xor U15807 (N_15807,N_10495,N_13384);
and U15808 (N_15808,N_11899,N_10420);
xnor U15809 (N_15809,N_13700,N_12023);
and U15810 (N_15810,N_14636,N_14873);
and U15811 (N_15811,N_13133,N_10095);
or U15812 (N_15812,N_13300,N_14316);
nand U15813 (N_15813,N_13568,N_11530);
and U15814 (N_15814,N_12792,N_11686);
xnor U15815 (N_15815,N_10250,N_14332);
and U15816 (N_15816,N_12791,N_13549);
nand U15817 (N_15817,N_13397,N_10116);
xor U15818 (N_15818,N_12052,N_14400);
xnor U15819 (N_15819,N_11719,N_14229);
xnor U15820 (N_15820,N_11474,N_11476);
nor U15821 (N_15821,N_12420,N_14273);
and U15822 (N_15822,N_13592,N_12057);
nand U15823 (N_15823,N_14519,N_13571);
xor U15824 (N_15824,N_10659,N_10089);
nor U15825 (N_15825,N_14350,N_12409);
xnor U15826 (N_15826,N_11795,N_14230);
xnor U15827 (N_15827,N_14149,N_13370);
nand U15828 (N_15828,N_10485,N_14551);
nor U15829 (N_15829,N_12829,N_10813);
or U15830 (N_15830,N_13437,N_14668);
xor U15831 (N_15831,N_11823,N_11088);
or U15832 (N_15832,N_13675,N_13154);
nor U15833 (N_15833,N_10804,N_14800);
and U15834 (N_15834,N_13143,N_10606);
or U15835 (N_15835,N_14849,N_13763);
nor U15836 (N_15836,N_14424,N_13751);
nor U15837 (N_15837,N_11282,N_13307);
nand U15838 (N_15838,N_12744,N_13035);
or U15839 (N_15839,N_13071,N_12636);
nand U15840 (N_15840,N_11797,N_14716);
nor U15841 (N_15841,N_10720,N_10716);
or U15842 (N_15842,N_14470,N_14659);
xor U15843 (N_15843,N_14317,N_13900);
xnor U15844 (N_15844,N_14254,N_13598);
or U15845 (N_15845,N_12808,N_11962);
and U15846 (N_15846,N_14291,N_10972);
xor U15847 (N_15847,N_14102,N_14018);
or U15848 (N_15848,N_12821,N_12116);
nand U15849 (N_15849,N_14764,N_10330);
and U15850 (N_15850,N_12010,N_11299);
and U15851 (N_15851,N_11237,N_12452);
nor U15852 (N_15852,N_12579,N_14399);
or U15853 (N_15853,N_13678,N_13973);
or U15854 (N_15854,N_13116,N_13361);
and U15855 (N_15855,N_11268,N_10416);
and U15856 (N_15856,N_14566,N_10310);
nor U15857 (N_15857,N_12250,N_10638);
or U15858 (N_15858,N_14223,N_13820);
nand U15859 (N_15859,N_12009,N_13941);
nand U15860 (N_15860,N_13355,N_13130);
or U15861 (N_15861,N_12814,N_14438);
xnor U15862 (N_15862,N_12819,N_11659);
or U15863 (N_15863,N_10366,N_13553);
or U15864 (N_15864,N_10085,N_12673);
nor U15865 (N_15865,N_14365,N_13803);
nor U15866 (N_15866,N_11177,N_13507);
nand U15867 (N_15867,N_13024,N_11105);
xor U15868 (N_15868,N_11858,N_10932);
nor U15869 (N_15869,N_10171,N_11693);
and U15870 (N_15870,N_11881,N_10120);
and U15871 (N_15871,N_14321,N_14053);
or U15872 (N_15872,N_12183,N_13907);
or U15873 (N_15873,N_10131,N_10951);
or U15874 (N_15874,N_14852,N_14192);
and U15875 (N_15875,N_13564,N_14414);
nand U15876 (N_15876,N_10771,N_10371);
nor U15877 (N_15877,N_11026,N_10887);
or U15878 (N_15878,N_14802,N_11898);
nor U15879 (N_15879,N_14487,N_11417);
xnor U15880 (N_15880,N_10873,N_10484);
nand U15881 (N_15881,N_10863,N_14642);
nand U15882 (N_15882,N_13055,N_14729);
nor U15883 (N_15883,N_11094,N_13672);
or U15884 (N_15884,N_10717,N_12130);
or U15885 (N_15885,N_12967,N_10956);
xor U15886 (N_15886,N_11441,N_13921);
or U15887 (N_15887,N_14571,N_11349);
nor U15888 (N_15888,N_13545,N_10729);
xnor U15889 (N_15889,N_13923,N_14122);
xnor U15890 (N_15890,N_10336,N_14322);
or U15891 (N_15891,N_11265,N_13056);
and U15892 (N_15892,N_10539,N_14363);
or U15893 (N_15893,N_11212,N_14213);
nand U15894 (N_15894,N_14639,N_10278);
xor U15895 (N_15895,N_10847,N_11197);
nor U15896 (N_15896,N_11992,N_12073);
and U15897 (N_15897,N_10052,N_14398);
or U15898 (N_15898,N_10731,N_13717);
and U15899 (N_15899,N_11421,N_14280);
xnor U15900 (N_15900,N_10710,N_12463);
and U15901 (N_15901,N_10407,N_12916);
xnor U15902 (N_15902,N_10759,N_12741);
or U15903 (N_15903,N_13095,N_10378);
or U15904 (N_15904,N_10918,N_13801);
nand U15905 (N_15905,N_14092,N_14941);
or U15906 (N_15906,N_14895,N_13968);
xor U15907 (N_15907,N_13123,N_11383);
and U15908 (N_15908,N_12522,N_10624);
xnor U15909 (N_15909,N_11384,N_10066);
and U15910 (N_15910,N_10645,N_10989);
and U15911 (N_15911,N_11755,N_14312);
or U15912 (N_15912,N_12972,N_13439);
nand U15913 (N_15913,N_12852,N_13282);
and U15914 (N_15914,N_13261,N_14256);
xnor U15915 (N_15915,N_13993,N_13358);
and U15916 (N_15916,N_13743,N_14478);
nand U15917 (N_15917,N_13694,N_11981);
nor U15918 (N_15918,N_13306,N_10042);
xor U15919 (N_15919,N_10930,N_11943);
nor U15920 (N_15920,N_12026,N_10699);
or U15921 (N_15921,N_14930,N_11572);
xnor U15922 (N_15922,N_12407,N_10777);
nor U15923 (N_15923,N_11557,N_11959);
nand U15924 (N_15924,N_10700,N_14917);
or U15925 (N_15925,N_10164,N_13669);
nand U15926 (N_15926,N_11663,N_12364);
nand U15927 (N_15927,N_14649,N_10785);
xnor U15928 (N_15928,N_11588,N_13290);
or U15929 (N_15929,N_10672,N_11040);
nand U15930 (N_15930,N_11988,N_14047);
nand U15931 (N_15931,N_14348,N_13336);
nor U15932 (N_15932,N_12570,N_10406);
and U15933 (N_15933,N_14811,N_14416);
nor U15934 (N_15934,N_14913,N_14236);
nor U15935 (N_15935,N_10911,N_10395);
nand U15936 (N_15936,N_12922,N_10020);
and U15937 (N_15937,N_12300,N_13332);
and U15938 (N_15938,N_14989,N_12358);
nor U15939 (N_15939,N_12386,N_14629);
nor U15940 (N_15940,N_14357,N_13709);
and U15941 (N_15941,N_13469,N_11679);
nand U15942 (N_15942,N_12639,N_13963);
nand U15943 (N_15943,N_13374,N_11704);
xnor U15944 (N_15944,N_10202,N_12557);
nor U15945 (N_15945,N_10078,N_11405);
and U15946 (N_15946,N_13220,N_13246);
or U15947 (N_15947,N_11714,N_10349);
and U15948 (N_15948,N_10964,N_10096);
or U15949 (N_15949,N_13552,N_13758);
nand U15950 (N_15950,N_11371,N_11168);
nor U15951 (N_15951,N_11085,N_12432);
and U15952 (N_15952,N_12779,N_10333);
and U15953 (N_15953,N_13600,N_12456);
or U15954 (N_15954,N_10832,N_11867);
nand U15955 (N_15955,N_14058,N_10839);
or U15956 (N_15956,N_10599,N_11767);
nand U15957 (N_15957,N_11614,N_10229);
nor U15958 (N_15958,N_14974,N_12981);
nand U15959 (N_15959,N_11138,N_14029);
xnor U15960 (N_15960,N_14076,N_13774);
xor U15961 (N_15961,N_13550,N_12051);
nor U15962 (N_15962,N_11043,N_11842);
and U15963 (N_15963,N_10765,N_11154);
or U15964 (N_15964,N_10481,N_12842);
xor U15965 (N_15965,N_10064,N_11190);
nand U15966 (N_15966,N_12142,N_11054);
and U15967 (N_15967,N_13242,N_12341);
xnor U15968 (N_15968,N_11207,N_14114);
xor U15969 (N_15969,N_13447,N_12672);
nand U15970 (N_15970,N_14012,N_12279);
nand U15971 (N_15971,N_13818,N_10187);
or U15972 (N_15972,N_10953,N_12405);
and U15973 (N_15973,N_13543,N_10334);
or U15974 (N_15974,N_11545,N_12710);
xor U15975 (N_15975,N_12697,N_12242);
xor U15976 (N_15976,N_14685,N_10372);
and U15977 (N_15977,N_10615,N_10170);
or U15978 (N_15978,N_13938,N_10247);
and U15979 (N_15979,N_10587,N_10935);
xor U15980 (N_15980,N_14440,N_10305);
nor U15981 (N_15981,N_14838,N_13101);
nor U15982 (N_15982,N_13548,N_11971);
nor U15983 (N_15983,N_14772,N_13350);
xnor U15984 (N_15984,N_11532,N_12946);
and U15985 (N_15985,N_12257,N_14621);
nor U15986 (N_15986,N_12221,N_13576);
xor U15987 (N_15987,N_12854,N_13070);
xor U15988 (N_15988,N_12647,N_14364);
or U15989 (N_15989,N_10177,N_13111);
nor U15990 (N_15990,N_13750,N_12074);
xnor U15991 (N_15991,N_11502,N_14109);
nand U15992 (N_15992,N_11442,N_10690);
nand U15993 (N_15993,N_11250,N_11339);
or U15994 (N_15994,N_12308,N_11161);
or U15995 (N_15995,N_12265,N_12907);
nand U15996 (N_15996,N_11695,N_11162);
and U15997 (N_15997,N_12612,N_14964);
and U15998 (N_15998,N_12295,N_12079);
and U15999 (N_15999,N_11826,N_10393);
or U16000 (N_16000,N_10526,N_11872);
and U16001 (N_16001,N_12914,N_14083);
xor U16002 (N_16002,N_10738,N_11974);
and U16003 (N_16003,N_13225,N_13251);
xor U16004 (N_16004,N_10691,N_12547);
nor U16005 (N_16005,N_14991,N_13064);
nand U16006 (N_16006,N_10460,N_13703);
nor U16007 (N_16007,N_12941,N_12247);
or U16008 (N_16008,N_14902,N_14751);
nand U16009 (N_16009,N_13495,N_13317);
or U16010 (N_16010,N_14697,N_11995);
or U16011 (N_16011,N_10882,N_11082);
nor U16012 (N_16012,N_14789,N_10602);
or U16013 (N_16013,N_10767,N_10191);
and U16014 (N_16014,N_13068,N_13349);
nor U16015 (N_16015,N_10796,N_10540);
or U16016 (N_16016,N_12095,N_11318);
xor U16017 (N_16017,N_12176,N_10057);
or U16018 (N_16018,N_10354,N_14534);
xnor U16019 (N_16019,N_14878,N_13103);
nor U16020 (N_16020,N_10306,N_10487);
or U16021 (N_16021,N_12961,N_14163);
xnor U16022 (N_16022,N_13861,N_10695);
nand U16023 (N_16023,N_12182,N_13558);
nand U16024 (N_16024,N_12583,N_12674);
nand U16025 (N_16025,N_13488,N_12783);
and U16026 (N_16026,N_13686,N_10452);
or U16027 (N_16027,N_13882,N_13431);
or U16028 (N_16028,N_11598,N_11263);
and U16029 (N_16029,N_11373,N_12124);
or U16030 (N_16030,N_11304,N_14020);
xor U16031 (N_16031,N_10462,N_14278);
nor U16032 (N_16032,N_10754,N_10735);
and U16033 (N_16033,N_13386,N_10363);
or U16034 (N_16034,N_10342,N_12366);
or U16035 (N_16035,N_12952,N_11067);
xor U16036 (N_16036,N_10787,N_14389);
or U16037 (N_16037,N_12092,N_12196);
nand U16038 (N_16038,N_14195,N_14937);
nand U16039 (N_16039,N_13913,N_11358);
nand U16040 (N_16040,N_10537,N_13083);
or U16041 (N_16041,N_13468,N_11805);
nand U16042 (N_16042,N_13426,N_12830);
xor U16043 (N_16043,N_10520,N_11252);
nor U16044 (N_16044,N_10877,N_14779);
and U16045 (N_16045,N_14495,N_10027);
nor U16046 (N_16046,N_12437,N_11593);
nand U16047 (N_16047,N_14301,N_14381);
xor U16048 (N_16048,N_13624,N_13265);
and U16049 (N_16049,N_10618,N_11940);
nand U16050 (N_16050,N_10380,N_11164);
nor U16051 (N_16051,N_10963,N_13432);
xnor U16052 (N_16052,N_13170,N_13456);
nor U16053 (N_16053,N_13581,N_12264);
or U16054 (N_16054,N_14257,N_12024);
and U16055 (N_16055,N_12321,N_12275);
nand U16056 (N_16056,N_14394,N_11260);
and U16057 (N_16057,N_12230,N_10288);
or U16058 (N_16058,N_13814,N_12920);
or U16059 (N_16059,N_12945,N_12345);
xnor U16060 (N_16060,N_11240,N_14262);
nor U16061 (N_16061,N_13022,N_13255);
nand U16062 (N_16062,N_14820,N_11487);
nand U16063 (N_16063,N_14643,N_13498);
or U16064 (N_16064,N_14474,N_12752);
xor U16065 (N_16065,N_14686,N_10341);
or U16066 (N_16066,N_10405,N_13159);
nor U16067 (N_16067,N_11027,N_13312);
xnor U16068 (N_16068,N_12161,N_14095);
or U16069 (N_16069,N_11117,N_13217);
xnor U16070 (N_16070,N_13948,N_10952);
nor U16071 (N_16071,N_11181,N_13491);
nor U16072 (N_16072,N_14453,N_11913);
nand U16073 (N_16073,N_12742,N_12846);
nor U16074 (N_16074,N_11658,N_12787);
nand U16075 (N_16075,N_12688,N_12068);
nand U16076 (N_16076,N_12512,N_12132);
and U16077 (N_16077,N_13193,N_11853);
and U16078 (N_16078,N_12857,N_10576);
or U16079 (N_16079,N_14355,N_11416);
or U16080 (N_16080,N_11157,N_10836);
xnor U16081 (N_16081,N_11187,N_13184);
or U16082 (N_16082,N_11368,N_11571);
xor U16083 (N_16083,N_13614,N_11862);
or U16084 (N_16084,N_10145,N_12314);
xor U16085 (N_16085,N_14118,N_13391);
nand U16086 (N_16086,N_11204,N_13984);
nor U16087 (N_16087,N_10469,N_14872);
nor U16088 (N_16088,N_12749,N_13573);
and U16089 (N_16089,N_13237,N_12204);
and U16090 (N_16090,N_12151,N_12251);
or U16091 (N_16091,N_14245,N_13707);
nor U16092 (N_16092,N_10917,N_11771);
or U16093 (N_16093,N_11828,N_13733);
xor U16094 (N_16094,N_10255,N_13728);
or U16095 (N_16095,N_13375,N_10263);
or U16096 (N_16096,N_11683,N_12592);
or U16097 (N_16097,N_14993,N_14922);
and U16098 (N_16098,N_10073,N_14766);
xor U16099 (N_16099,N_14951,N_12822);
and U16100 (N_16100,N_12562,N_10625);
nor U16101 (N_16101,N_12169,N_11705);
nand U16102 (N_16102,N_14379,N_12959);
xor U16103 (N_16103,N_14269,N_12693);
or U16104 (N_16104,N_13289,N_11590);
and U16105 (N_16105,N_11324,N_12620);
nand U16106 (N_16106,N_12487,N_11080);
nand U16107 (N_16107,N_12628,N_10444);
xnor U16108 (N_16108,N_12616,N_10181);
xnor U16109 (N_16109,N_14674,N_13922);
and U16110 (N_16110,N_13701,N_12374);
nor U16111 (N_16111,N_11498,N_14539);
nor U16112 (N_16112,N_14900,N_10852);
xnor U16113 (N_16113,N_14003,N_13172);
nand U16114 (N_16114,N_14288,N_14687);
xnor U16115 (N_16115,N_13423,N_10748);
nor U16116 (N_16116,N_13482,N_13504);
nand U16117 (N_16117,N_13318,N_13649);
and U16118 (N_16118,N_10475,N_13933);
nand U16119 (N_16119,N_12215,N_13376);
or U16120 (N_16120,N_10586,N_13309);
xor U16121 (N_16121,N_12976,N_12395);
nor U16122 (N_16122,N_12382,N_13286);
nand U16123 (N_16123,N_14422,N_14683);
nor U16124 (N_16124,N_13304,N_13593);
nand U16125 (N_16125,N_12439,N_14689);
or U16126 (N_16126,N_14522,N_12192);
nor U16127 (N_16127,N_14392,N_13321);
and U16128 (N_16128,N_11480,N_11455);
nor U16129 (N_16129,N_12553,N_12494);
nand U16130 (N_16130,N_11242,N_12065);
or U16131 (N_16131,N_12291,N_12105);
xnor U16132 (N_16132,N_10853,N_12800);
nand U16133 (N_16133,N_10529,N_10966);
xor U16134 (N_16134,N_13666,N_10954);
nand U16135 (N_16135,N_11917,N_11543);
xor U16136 (N_16136,N_10825,N_14777);
nand U16137 (N_16137,N_13086,N_10591);
and U16138 (N_16138,N_12933,N_11091);
or U16139 (N_16139,N_14393,N_10226);
nand U16140 (N_16140,N_14452,N_12232);
or U16141 (N_16141,N_13425,N_12248);
and U16142 (N_16142,N_12121,N_11408);
or U16143 (N_16143,N_14707,N_13970);
xor U16144 (N_16144,N_14883,N_14300);
nand U16145 (N_16145,N_10067,N_11423);
or U16146 (N_16146,N_13485,N_10304);
xnor U16147 (N_16147,N_11706,N_13021);
and U16148 (N_16148,N_10437,N_11276);
nor U16149 (N_16149,N_10590,N_13392);
or U16150 (N_16150,N_12148,N_12067);
or U16151 (N_16151,N_10582,N_13802);
and U16152 (N_16152,N_13831,N_11228);
or U16153 (N_16153,N_12917,N_12427);
xnor U16154 (N_16154,N_11617,N_10438);
or U16155 (N_16155,N_14456,N_11218);
or U16156 (N_16156,N_10978,N_12266);
or U16157 (N_16157,N_10916,N_11568);
xnor U16158 (N_16158,N_14224,N_13241);
or U16159 (N_16159,N_11607,N_14443);
nor U16160 (N_16160,N_14499,N_10840);
nand U16161 (N_16161,N_12388,N_10958);
xor U16162 (N_16162,N_12089,N_10408);
nor U16163 (N_16163,N_11139,N_10102);
nand U16164 (N_16164,N_13719,N_10376);
and U16165 (N_16165,N_14105,N_11118);
xor U16166 (N_16166,N_11674,N_14896);
and U16167 (N_16167,N_10271,N_11108);
nand U16168 (N_16168,N_14437,N_12333);
nand U16169 (N_16169,N_11262,N_11742);
or U16170 (N_16170,N_12473,N_11745);
and U16171 (N_16171,N_11148,N_12368);
and U16172 (N_16172,N_11987,N_14877);
or U16173 (N_16173,N_11677,N_11478);
and U16174 (N_16174,N_13597,N_13151);
and U16175 (N_16175,N_14136,N_12773);
nand U16176 (N_16176,N_13364,N_11852);
or U16177 (N_16177,N_14961,N_10126);
nor U16178 (N_16178,N_14576,N_14211);
nor U16179 (N_16179,N_14533,N_10215);
or U16180 (N_16180,N_11906,N_10811);
and U16181 (N_16181,N_10859,N_11758);
nand U16182 (N_16182,N_11644,N_10425);
and U16183 (N_16183,N_10365,N_13428);
and U16184 (N_16184,N_11773,N_11065);
nor U16185 (N_16185,N_13042,N_14420);
and U16186 (N_16186,N_12748,N_14023);
nor U16187 (N_16187,N_14679,N_13125);
nor U16188 (N_16188,N_14975,N_14299);
nand U16189 (N_16189,N_10143,N_11020);
or U16190 (N_16190,N_14051,N_10403);
xor U16191 (N_16191,N_14641,N_14898);
and U16192 (N_16192,N_14826,N_12731);
or U16193 (N_16193,N_11132,N_14033);
nand U16194 (N_16194,N_10547,N_10849);
nor U16195 (N_16195,N_13032,N_13047);
xor U16196 (N_16196,N_14180,N_13630);
or U16197 (N_16197,N_13207,N_12712);
nor U16198 (N_16198,N_12309,N_14441);
or U16199 (N_16199,N_12290,N_11386);
xor U16200 (N_16200,N_10603,N_10653);
and U16201 (N_16201,N_14675,N_11975);
nor U16202 (N_16202,N_14314,N_11628);
nand U16203 (N_16203,N_13808,N_10015);
nor U16204 (N_16204,N_14368,N_11052);
and U16205 (N_16205,N_11389,N_13946);
xor U16206 (N_16206,N_11101,N_12393);
or U16207 (N_16207,N_10983,N_13206);
nand U16208 (N_16208,N_14773,N_11725);
xor U16209 (N_16209,N_11113,N_14603);
and U16210 (N_16210,N_11310,N_10207);
and U16211 (N_16211,N_14693,N_11654);
and U16212 (N_16212,N_13660,N_10308);
xnor U16213 (N_16213,N_11433,N_11513);
or U16214 (N_16214,N_12546,N_13952);
and U16215 (N_16215,N_10217,N_10297);
or U16216 (N_16216,N_10904,N_10723);
and U16217 (N_16217,N_12174,N_14493);
and U16218 (N_16218,N_14359,N_10282);
and U16219 (N_16219,N_14787,N_12191);
or U16220 (N_16220,N_12651,N_11317);
nor U16221 (N_16221,N_10080,N_11750);
xnor U16222 (N_16222,N_10531,N_14665);
and U16223 (N_16223,N_14283,N_13596);
and U16224 (N_16224,N_11875,N_11631);
nor U16225 (N_16225,N_10194,N_14268);
nor U16226 (N_16226,N_14135,N_13852);
or U16227 (N_16227,N_10076,N_13896);
and U16228 (N_16228,N_14277,N_12747);
and U16229 (N_16229,N_12496,N_10267);
and U16230 (N_16230,N_10498,N_13650);
or U16231 (N_16231,N_11400,N_11471);
or U16232 (N_16232,N_12338,N_12885);
nor U16233 (N_16233,N_12630,N_14086);
xnor U16234 (N_16234,N_14270,N_11737);
xnor U16235 (N_16235,N_13621,N_14184);
nand U16236 (N_16236,N_11914,N_13434);
nand U16237 (N_16237,N_11720,N_10154);
nor U16238 (N_16238,N_11713,N_10369);
xor U16239 (N_16239,N_13990,N_14958);
nand U16240 (N_16240,N_10195,N_10389);
nand U16241 (N_16241,N_11908,N_14313);
and U16242 (N_16242,N_11759,N_10122);
xnor U16243 (N_16243,N_11440,N_13017);
or U16244 (N_16244,N_10510,N_11868);
and U16245 (N_16245,N_14620,N_13212);
nor U16246 (N_16246,N_11629,N_14821);
and U16247 (N_16247,N_12520,N_12032);
nand U16248 (N_16248,N_12033,N_13027);
and U16249 (N_16249,N_10546,N_10646);
nand U16250 (N_16250,N_10810,N_10430);
nor U16251 (N_16251,N_13590,N_12598);
or U16252 (N_16252,N_14730,N_10329);
or U16253 (N_16253,N_11845,N_13806);
xnor U16254 (N_16254,N_13158,N_10974);
nor U16255 (N_16255,N_10946,N_11647);
nand U16256 (N_16256,N_14261,N_12827);
xnor U16257 (N_16257,N_12149,N_12627);
and U16258 (N_16258,N_14631,N_13747);
nor U16259 (N_16259,N_13499,N_13604);
nand U16260 (N_16260,N_10346,N_14429);
and U16261 (N_16261,N_10219,N_13883);
nor U16262 (N_16262,N_11392,N_12863);
or U16263 (N_16263,N_10730,N_11636);
nand U16264 (N_16264,N_10878,N_13724);
nor U16265 (N_16265,N_10084,N_11682);
xnor U16266 (N_16266,N_14927,N_11465);
xor U16267 (N_16267,N_14319,N_12662);
or U16268 (N_16268,N_13445,N_14514);
nand U16269 (N_16269,N_10418,N_14164);
xnor U16270 (N_16270,N_12754,N_10225);
nor U16271 (N_16271,N_12118,N_14148);
and U16272 (N_16272,N_14672,N_13277);
or U16273 (N_16273,N_12150,N_11698);
and U16274 (N_16274,N_14338,N_13508);
nand U16275 (N_16275,N_11717,N_10931);
nor U16276 (N_16276,N_10204,N_10897);
nor U16277 (N_16277,N_11360,N_12440);
xor U16278 (N_16278,N_13786,N_13692);
or U16279 (N_16279,N_12090,N_12042);
or U16280 (N_16280,N_14106,N_13073);
xor U16281 (N_16281,N_13451,N_12708);
xor U16282 (N_16282,N_14144,N_12709);
and U16283 (N_16283,N_12352,N_14967);
or U16284 (N_16284,N_14178,N_10692);
or U16285 (N_16285,N_14987,N_12155);
or U16286 (N_16286,N_12084,N_12996);
nand U16287 (N_16287,N_13243,N_14281);
and U16288 (N_16288,N_10536,N_11361);
and U16289 (N_16289,N_12471,N_13957);
and U16290 (N_16290,N_14607,N_10069);
and U16291 (N_16291,N_10141,N_11662);
and U16292 (N_16292,N_13512,N_13847);
or U16293 (N_16293,N_13644,N_11325);
or U16294 (N_16294,N_12685,N_10924);
nor U16295 (N_16295,N_12517,N_11520);
and U16296 (N_16296,N_14091,N_11195);
or U16297 (N_16297,N_10210,N_13405);
xnor U16298 (N_16298,N_12403,N_14960);
or U16299 (N_16299,N_12987,N_11613);
or U16300 (N_16300,N_12655,N_11083);
nand U16301 (N_16301,N_13394,N_13132);
nand U16302 (N_16302,N_14600,N_12005);
nand U16303 (N_16303,N_12556,N_11469);
nand U16304 (N_16304,N_13354,N_13505);
or U16305 (N_16305,N_12152,N_11211);
nor U16306 (N_16306,N_10268,N_12935);
nand U16307 (N_16307,N_11467,N_10023);
nand U16308 (N_16308,N_11266,N_10792);
xor U16309 (N_16309,N_11036,N_11302);
or U16310 (N_16310,N_13836,N_10245);
xor U16311 (N_16311,N_11256,N_12123);
nor U16312 (N_16312,N_13643,N_12041);
xnor U16313 (N_16313,N_12206,N_14320);
nor U16314 (N_16314,N_11927,N_12381);
and U16315 (N_16315,N_13080,N_12498);
nor U16316 (N_16316,N_13817,N_11840);
nor U16317 (N_16317,N_14768,N_13442);
xnor U16318 (N_16318,N_11997,N_14310);
nor U16319 (N_16319,N_10351,N_13096);
or U16320 (N_16320,N_10301,N_11569);
or U16321 (N_16321,N_10790,N_11581);
and U16322 (N_16322,N_11456,N_10502);
or U16323 (N_16323,N_14431,N_10507);
nand U16324 (N_16324,N_13438,N_10605);
nand U16325 (N_16325,N_11746,N_11221);
or U16326 (N_16326,N_11655,N_12965);
xnor U16327 (N_16327,N_14527,N_12387);
nand U16328 (N_16328,N_13877,N_14782);
or U16329 (N_16329,N_12144,N_14461);
xor U16330 (N_16330,N_14055,N_13812);
and U16331 (N_16331,N_13069,N_13773);
xor U16332 (N_16332,N_12305,N_14932);
nand U16333 (N_16333,N_14708,N_12449);
nand U16334 (N_16334,N_12701,N_10185);
nor U16335 (N_16335,N_10362,N_11509);
or U16336 (N_16336,N_11886,N_10285);
or U16337 (N_16337,N_14531,N_13087);
or U16338 (N_16338,N_12441,N_13752);
nor U16339 (N_16339,N_12906,N_12529);
and U16340 (N_16340,N_10451,N_14482);
or U16341 (N_16341,N_10920,N_14723);
nand U16342 (N_16342,N_10883,N_10021);
xnor U16343 (N_16343,N_13609,N_11863);
or U16344 (N_16344,N_14315,N_13067);
or U16345 (N_16345,N_12670,N_11342);
xor U16346 (N_16346,N_12992,N_14200);
xor U16347 (N_16347,N_10929,N_14855);
or U16348 (N_16348,N_14308,N_13647);
nor U16349 (N_16349,N_12915,N_12216);
nor U16350 (N_16350,N_14808,N_10990);
nor U16351 (N_16351,N_11837,N_10293);
and U16352 (N_16352,N_11109,N_13075);
or U16353 (N_16353,N_11122,N_10054);
or U16354 (N_16354,N_13026,N_13839);
xor U16355 (N_16355,N_12423,N_14426);
nor U16356 (N_16356,N_10424,N_12287);
or U16357 (N_16357,N_10321,N_10596);
xor U16358 (N_16358,N_14294,N_14581);
nor U16359 (N_16359,N_11751,N_11393);
or U16360 (N_16360,N_13271,N_10269);
and U16361 (N_16361,N_12351,N_10343);
and U16362 (N_16362,N_11013,N_12324);
nand U16363 (N_16363,N_10482,N_13898);
and U16364 (N_16364,N_10999,N_14992);
or U16365 (N_16365,N_11093,N_11251);
and U16366 (N_16366,N_14134,N_11064);
or U16367 (N_16367,N_10732,N_14962);
or U16368 (N_16368,N_13633,N_13569);
or U16369 (N_16369,N_14935,N_10348);
nor U16370 (N_16370,N_12200,N_12066);
xnor U16371 (N_16371,N_13939,N_11735);
nor U16372 (N_16372,N_11587,N_10884);
xnor U16373 (N_16373,N_14714,N_10390);
xor U16374 (N_16374,N_13315,N_13114);
xor U16375 (N_16375,N_10127,N_11464);
nand U16376 (N_16376,N_12778,N_10971);
xnor U16377 (N_16377,N_12953,N_14084);
or U16378 (N_16378,N_13971,N_14980);
or U16379 (N_16379,N_14193,N_10399);
and U16380 (N_16380,N_12501,N_12312);
nand U16381 (N_16381,N_12046,N_13528);
nand U16382 (N_16382,N_12363,N_11702);
nor U16383 (N_16383,N_12108,N_13646);
xor U16384 (N_16384,N_12634,N_11727);
or U16385 (N_16385,N_14170,N_14733);
xor U16386 (N_16386,N_11321,N_13726);
nor U16387 (N_16387,N_11202,N_11832);
or U16388 (N_16388,N_11016,N_14297);
and U16389 (N_16389,N_13411,N_12283);
nor U16390 (N_16390,N_14457,N_10397);
xor U16391 (N_16391,N_11766,N_13862);
nor U16392 (N_16392,N_12022,N_13740);
or U16393 (N_16393,N_10302,N_14921);
nor U16394 (N_16394,N_12491,N_12970);
nand U16395 (N_16395,N_14832,N_10922);
or U16396 (N_16396,N_12788,N_10071);
xor U16397 (N_16397,N_11403,N_13465);
and U16398 (N_16398,N_10253,N_13099);
or U16399 (N_16399,N_13164,N_13955);
and U16400 (N_16400,N_11472,N_13205);
nand U16401 (N_16401,N_12229,N_13540);
nor U16402 (N_16402,N_11151,N_14503);
or U16403 (N_16403,N_13844,N_12763);
and U16404 (N_16404,N_10558,N_12146);
xnor U16405 (N_16405,N_10588,N_12406);
nor U16406 (N_16406,N_10533,N_10757);
nand U16407 (N_16407,N_11944,N_13232);
and U16408 (N_16408,N_13063,N_14871);
xnor U16409 (N_16409,N_13072,N_10385);
nor U16410 (N_16410,N_10517,N_10557);
xor U16411 (N_16411,N_14255,N_10317);
nand U16412 (N_16412,N_13634,N_14824);
nand U16413 (N_16413,N_12284,N_13140);
nor U16414 (N_16414,N_12558,N_11225);
xor U16415 (N_16415,N_13213,N_13842);
nand U16416 (N_16416,N_10634,N_11901);
or U16417 (N_16417,N_13449,N_10146);
xor U16418 (N_16418,N_13869,N_12039);
nor U16419 (N_16419,N_12600,N_13765);
nor U16420 (N_16420,N_11042,N_12234);
nand U16421 (N_16421,N_11484,N_11784);
nand U16422 (N_16422,N_14063,N_12828);
xnor U16423 (N_16423,N_14071,N_14915);
and U16424 (N_16424,N_13620,N_13975);
or U16425 (N_16425,N_11335,N_11179);
nand U16426 (N_16426,N_12807,N_10068);
nor U16427 (N_16427,N_11376,N_14077);
and U16428 (N_16428,N_11131,N_14206);
and U16429 (N_16429,N_12318,N_13410);
or U16430 (N_16430,N_10905,N_14894);
or U16431 (N_16431,N_10574,N_10313);
or U16432 (N_16432,N_11578,N_12745);
xor U16433 (N_16433,N_10478,N_10463);
and U16434 (N_16434,N_12274,N_13999);
and U16435 (N_16435,N_14804,N_10616);
xnor U16436 (N_16436,N_13403,N_11942);
or U16437 (N_16437,N_11900,N_14451);
nand U16438 (N_16438,N_14477,N_10392);
nor U16439 (N_16439,N_12080,N_11398);
nand U16440 (N_16440,N_14585,N_11958);
or U16441 (N_16441,N_11567,N_12559);
and U16442 (N_16442,N_12347,N_11641);
and U16443 (N_16443,N_11429,N_14968);
nor U16444 (N_16444,N_14017,N_12337);
xnor U16445 (N_16445,N_14540,N_12722);
nor U16446 (N_16446,N_10604,N_10942);
xnor U16447 (N_16447,N_12669,N_12705);
xnor U16448 (N_16448,N_13636,N_12767);
and U16449 (N_16449,N_11123,N_14183);
xnor U16450 (N_16450,N_13209,N_12278);
nand U16451 (N_16451,N_12243,N_12581);
or U16452 (N_16452,N_11279,N_12054);
and U16453 (N_16453,N_12101,N_10139);
nand U16454 (N_16454,N_11297,N_12926);
xnor U16455 (N_16455,N_11338,N_11618);
or U16456 (N_16456,N_10865,N_14647);
xnor U16457 (N_16457,N_13557,N_12263);
nor U16458 (N_16458,N_14169,N_10568);
or U16459 (N_16459,N_12645,N_13215);
and U16460 (N_16460,N_14651,N_13038);
nor U16461 (N_16461,N_14957,N_11095);
xnor U16462 (N_16462,N_12385,N_13057);
and U16463 (N_16463,N_10986,N_11887);
or U16464 (N_16464,N_11865,N_12447);
nor U16465 (N_16465,N_14670,N_11103);
or U16466 (N_16466,N_11909,N_13084);
and U16467 (N_16467,N_14627,N_14617);
and U16468 (N_16468,N_10169,N_11998);
nand U16469 (N_16469,N_13688,N_13280);
nor U16470 (N_16470,N_11950,N_11333);
xnor U16471 (N_16471,N_11035,N_11185);
nand U16472 (N_16472,N_10235,N_10428);
or U16473 (N_16473,N_11078,N_10441);
xnor U16474 (N_16474,N_11525,N_10621);
xor U16475 (N_16475,N_11780,N_14925);
nor U16476 (N_16476,N_13429,N_12493);
xor U16477 (N_16477,N_13346,N_11402);
and U16478 (N_16478,N_13378,N_10188);
nor U16479 (N_16479,N_11153,N_12050);
nand U16480 (N_16480,N_12649,N_14805);
nor U16481 (N_16481,N_10739,N_13049);
nor U16482 (N_16482,N_11610,N_14088);
and U16483 (N_16483,N_11293,N_12246);
and U16484 (N_16484,N_14228,N_11756);
nand U16485 (N_16485,N_10002,N_14926);
xnor U16486 (N_16486,N_10086,N_10727);
and U16487 (N_16487,N_10552,N_10375);
nor U16488 (N_16488,N_12511,N_14549);
nand U16489 (N_16489,N_11047,N_13742);
and U16490 (N_16490,N_14609,N_13311);
and U16491 (N_16491,N_11859,N_14502);
nor U16492 (N_16492,N_14276,N_13783);
nor U16493 (N_16493,N_11517,N_11494);
xor U16494 (N_16494,N_11070,N_14346);
xnor U16495 (N_16495,N_12354,N_14758);
xor U16496 (N_16496,N_14694,N_14186);
nor U16497 (N_16497,N_10749,N_12771);
and U16498 (N_16498,N_13640,N_13816);
and U16499 (N_16499,N_10955,N_10184);
or U16500 (N_16500,N_11721,N_14799);
or U16501 (N_16501,N_13458,N_13606);
xor U16502 (N_16502,N_12949,N_11450);
nand U16503 (N_16503,N_14742,N_10322);
xor U16504 (N_16504,N_13496,N_13065);
or U16505 (N_16505,N_11601,N_10947);
nor U16506 (N_16506,N_10316,N_14371);
xnor U16507 (N_16507,N_11319,N_12503);
and U16508 (N_16508,N_14022,N_12336);
or U16509 (N_16509,N_13910,N_10975);
xnor U16510 (N_16510,N_10166,N_14823);
nand U16511 (N_16511,N_13382,N_12140);
xor U16512 (N_16512,N_13532,N_14302);
nor U16513 (N_16513,N_11114,N_14423);
and U16514 (N_16514,N_13947,N_10471);
and U16515 (N_16515,N_14247,N_13770);
or U16516 (N_16516,N_10298,N_14575);
and U16517 (N_16517,N_12740,N_10032);
nor U16518 (N_16518,N_12426,N_11006);
or U16519 (N_16519,N_12431,N_13211);
nand U16520 (N_16520,N_14471,N_12700);
nor U16521 (N_16521,N_14530,N_10910);
or U16522 (N_16522,N_14358,N_10927);
xnor U16523 (N_16523,N_11406,N_14506);
or U16524 (N_16524,N_11312,N_12879);
nand U16525 (N_16525,N_12824,N_14691);
nor U16526 (N_16526,N_11505,N_11163);
or U16527 (N_16527,N_14536,N_13288);
nand U16528 (N_16528,N_12638,N_12937);
nand U16529 (N_16529,N_13033,N_13327);
nor U16530 (N_16530,N_13359,N_14557);
xor U16531 (N_16531,N_12853,N_14577);
nor U16532 (N_16532,N_12085,N_10808);
nor U16533 (N_16533,N_12635,N_13179);
nor U16534 (N_16534,N_11205,N_10213);
and U16535 (N_16535,N_11014,N_11594);
and U16536 (N_16536,N_11060,N_10980);
or U16537 (N_16537,N_11496,N_11180);
nor U16538 (N_16538,N_12813,N_10412);
or U16539 (N_16539,N_12186,N_11710);
xor U16540 (N_16540,N_12864,N_13622);
nand U16541 (N_16541,N_13254,N_11500);
and U16542 (N_16542,N_14976,N_14891);
nand U16543 (N_16543,N_12584,N_10419);
nand U16544 (N_16544,N_11524,N_14473);
and U16545 (N_16545,N_14016,N_13260);
and U16546 (N_16546,N_13702,N_10525);
nor U16547 (N_16547,N_11160,N_10521);
xnor U16548 (N_16548,N_10493,N_14099);
nor U16549 (N_16549,N_13828,N_13201);
or U16550 (N_16550,N_14006,N_14573);
and U16551 (N_16551,N_14599,N_13299);
nor U16552 (N_16552,N_11866,N_13611);
and U16553 (N_16553,N_11089,N_12302);
xor U16554 (N_16554,N_12500,N_10199);
or U16555 (N_16555,N_14435,N_13117);
and U16556 (N_16556,N_12015,N_14760);
nand U16557 (N_16557,N_14667,N_14653);
and U16558 (N_16558,N_12412,N_11222);
or U16559 (N_16559,N_13287,N_12139);
xnor U16560 (N_16560,N_10664,N_11652);
or U16561 (N_16561,N_10921,N_13152);
nor U16562 (N_16562,N_13257,N_10619);
nand U16563 (N_16563,N_11399,N_14699);
and U16564 (N_16564,N_14830,N_11391);
xnor U16565 (N_16565,N_12081,N_10347);
nand U16566 (N_16566,N_11305,N_12782);
xor U16567 (N_16567,N_11512,N_13041);
xnor U16568 (N_16568,N_10132,N_10793);
nor U16569 (N_16569,N_14225,N_11577);
nand U16570 (N_16570,N_12180,N_14227);
and U16571 (N_16571,N_11023,N_14108);
nor U16572 (N_16572,N_11576,N_12099);
and U16573 (N_16573,N_13115,N_11691);
and U16574 (N_16574,N_13500,N_14914);
and U16575 (N_16575,N_12231,N_13951);
xor U16576 (N_16576,N_12165,N_14366);
and U16577 (N_16577,N_13436,N_13404);
nand U16578 (N_16578,N_10234,N_13413);
nor U16579 (N_16579,N_12064,N_13906);
and U16580 (N_16580,N_10841,N_12002);
nand U16581 (N_16581,N_13284,N_14746);
xor U16582 (N_16582,N_13486,N_13341);
nor U16583 (N_16583,N_11993,N_12378);
nand U16584 (N_16584,N_12226,N_13169);
xor U16585 (N_16585,N_10881,N_11322);
or U16586 (N_16586,N_13295,N_12606);
or U16587 (N_16587,N_13000,N_10823);
xnor U16588 (N_16588,N_11573,N_11815);
and U16589 (N_16589,N_12919,N_11848);
nand U16590 (N_16590,N_13353,N_14908);
nand U16591 (N_16591,N_14367,N_12997);
nand U16592 (N_16592,N_13841,N_11348);
and U16593 (N_16593,N_11774,N_12157);
xnor U16594 (N_16594,N_11460,N_12832);
and U16595 (N_16595,N_12454,N_13994);
nand U16596 (N_16596,N_12444,N_14905);
nor U16597 (N_16597,N_10807,N_11827);
nor U16598 (N_16598,N_12695,N_14031);
xor U16599 (N_16599,N_12268,N_13460);
or U16600 (N_16600,N_12098,N_11555);
nor U16601 (N_16601,N_11769,N_12269);
and U16602 (N_16602,N_13979,N_14121);
nand U16603 (N_16603,N_14712,N_14496);
xnor U16604 (N_16604,N_11007,N_10051);
xnor U16605 (N_16605,N_12619,N_11443);
xnor U16606 (N_16606,N_11533,N_14155);
or U16607 (N_16607,N_10945,N_13503);
and U16608 (N_16608,N_13138,N_12304);
xnor U16609 (N_16609,N_12421,N_14187);
nand U16610 (N_16610,N_12394,N_11159);
nand U16611 (N_16611,N_14682,N_14525);
nand U16612 (N_16612,N_11233,N_12392);
xor U16613 (N_16613,N_14490,N_11024);
or U16614 (N_16614,N_13784,N_12938);
or U16615 (N_16615,N_11645,N_14235);
nand U16616 (N_16616,N_13969,N_13879);
and U16617 (N_16617,N_13053,N_14904);
xor U16618 (N_16618,N_13020,N_11565);
nor U16619 (N_16619,N_14634,N_13623);
nand U16620 (N_16620,N_10050,N_14137);
and U16621 (N_16621,N_13991,N_12134);
nand U16622 (N_16622,N_14489,N_14203);
nand U16623 (N_16623,N_12715,N_14762);
and U16624 (N_16624,N_12091,N_12561);
and U16625 (N_16625,N_10733,N_11925);
and U16626 (N_16626,N_11619,N_14165);
xor U16627 (N_16627,N_11570,N_13811);
xor U16628 (N_16628,N_14336,N_11128);
xnor U16629 (N_16629,N_14934,N_14199);
or U16630 (N_16630,N_14447,N_12346);
nor U16631 (N_16631,N_11445,N_12097);
nand U16632 (N_16632,N_12928,N_12841);
and U16633 (N_16633,N_13785,N_10514);
nor U16634 (N_16634,N_11144,N_14611);
or U16635 (N_16635,N_10845,N_12096);
and U16636 (N_16636,N_12966,N_11022);
or U16637 (N_16637,N_13725,N_10711);
nor U16638 (N_16638,N_13917,N_10423);
nor U16639 (N_16639,N_12858,N_12233);
or U16640 (N_16640,N_12379,N_14267);
and U16641 (N_16641,N_11579,N_12866);
nor U16642 (N_16642,N_14259,N_11194);
or U16643 (N_16643,N_11142,N_13324);
and U16644 (N_16644,N_10214,N_11340);
xnor U16645 (N_16645,N_12692,N_12869);
nand U16646 (N_16646,N_10775,N_13247);
nand U16647 (N_16647,N_14724,N_11344);
nor U16648 (N_16648,N_13586,N_10291);
or U16649 (N_16649,N_12527,N_12904);
nor U16650 (N_16650,N_14950,N_12311);
and U16651 (N_16651,N_12998,N_10809);
or U16652 (N_16652,N_13414,N_10072);
nor U16653 (N_16653,N_12702,N_12037);
nand U16654 (N_16654,N_13772,N_11967);
or U16655 (N_16655,N_12138,N_10795);
and U16656 (N_16656,N_14011,N_14538);
xor U16657 (N_16657,N_14875,N_12596);
nor U16658 (N_16658,N_14853,N_14710);
nand U16659 (N_16659,N_10665,N_14101);
or U16660 (N_16660,N_14387,N_11637);
nand U16661 (N_16661,N_12785,N_12448);
and U16662 (N_16662,N_14788,N_11612);
and U16663 (N_16663,N_13584,N_14442);
nor U16664 (N_16664,N_10038,N_13389);
nand U16665 (N_16665,N_10934,N_12848);
nand U16666 (N_16666,N_13676,N_13147);
or U16667 (N_16667,N_13489,N_12006);
xor U16668 (N_16668,N_11932,N_10055);
nor U16669 (N_16669,N_14616,N_11660);
and U16670 (N_16670,N_10396,N_12897);
or U16671 (N_16671,N_11239,N_11788);
and U16672 (N_16672,N_14845,N_10240);
xnor U16673 (N_16673,N_11982,N_14780);
xor U16674 (N_16674,N_11330,N_14124);
and U16675 (N_16675,N_14892,N_10981);
nand U16676 (N_16676,N_10519,N_11178);
xnor U16677 (N_16677,N_14069,N_12549);
xnor U16678 (N_16678,N_13824,N_13412);
or U16679 (N_16679,N_12211,N_12817);
and U16680 (N_16680,N_10496,N_13691);
nand U16681 (N_16681,N_10820,N_12684);
nor U16682 (N_16682,N_13417,N_10172);
and U16683 (N_16683,N_14342,N_12218);
and U16684 (N_16684,N_10835,N_10550);
and U16685 (N_16685,N_13145,N_11854);
nand U16686 (N_16686,N_12642,N_13393);
and U16687 (N_16687,N_11186,N_14113);
xnor U16688 (N_16688,N_13407,N_13680);
nor U16689 (N_16689,N_12497,N_10516);
nand U16690 (N_16690,N_13281,N_10256);
or U16691 (N_16691,N_11435,N_13144);
or U16692 (N_16692,N_11985,N_13487);
xor U16693 (N_16693,N_13536,N_11889);
and U16694 (N_16694,N_10556,N_10880);
or U16695 (N_16695,N_11535,N_13244);
xor U16696 (N_16696,N_13534,N_12329);
and U16697 (N_16697,N_12746,N_11430);
nor U16698 (N_16698,N_13628,N_10016);
nor U16699 (N_16699,N_10254,N_12056);
and U16700 (N_16700,N_13002,N_12451);
nor U16701 (N_16701,N_10745,N_11362);
and U16702 (N_16702,N_13174,N_12129);
nor U16703 (N_16703,N_10766,N_10612);
nand U16704 (N_16704,N_13173,N_14253);
nand U16705 (N_16705,N_14542,N_11313);
or U16706 (N_16706,N_14718,N_11544);
nor U16707 (N_16707,N_12721,N_10237);
xor U16708 (N_16708,N_14574,N_12535);
nand U16709 (N_16709,N_10440,N_10446);
or U16710 (N_16710,N_12413,N_11978);
xor U16711 (N_16711,N_13018,N_12889);
and U16712 (N_16712,N_14032,N_12372);
and U16713 (N_16713,N_13344,N_12552);
nor U16714 (N_16714,N_10822,N_14614);
or U16715 (N_16715,N_14128,N_10891);
nor U16716 (N_16716,N_10567,N_13745);
and U16717 (N_16717,N_12762,N_14564);
xnor U16718 (N_16718,N_12348,N_13880);
and U16719 (N_16719,N_11003,N_10899);
nand U16720 (N_16720,N_12126,N_12011);
xor U16721 (N_16721,N_13714,N_11420);
nand U16722 (N_16722,N_12924,N_11428);
nand U16723 (N_16723,N_13805,N_14373);
or U16724 (N_16724,N_10091,N_12844);
and U16725 (N_16725,N_10561,N_12255);
xnor U16726 (N_16726,N_13239,N_14260);
nand U16727 (N_16727,N_12171,N_11856);
xor U16728 (N_16728,N_10000,N_10490);
nor U16729 (N_16729,N_10243,N_12980);
nand U16730 (N_16730,N_11058,N_13523);
nor U16731 (N_16731,N_12521,N_11670);
nand U16732 (N_16732,N_11076,N_14630);
nand U16733 (N_16733,N_14899,N_13793);
nor U16734 (N_16734,N_14397,N_12189);
nor U16735 (N_16735,N_14572,N_10886);
nor U16736 (N_16736,N_13608,N_10101);
or U16737 (N_16737,N_14013,N_12661);
nor U16738 (N_16738,N_12486,N_10914);
nor U16739 (N_16739,N_13997,N_10818);
and U16740 (N_16740,N_13904,N_13551);
and U16741 (N_16741,N_10902,N_14218);
nor U16742 (N_16742,N_14986,N_12060);
nand U16743 (N_16743,N_11604,N_12962);
and U16744 (N_16744,N_13663,N_12793);
or U16745 (N_16745,N_11611,N_13778);
and U16746 (N_16746,N_11401,N_13270);
or U16747 (N_16747,N_10770,N_11801);
nand U16748 (N_16748,N_14757,N_11385);
nor U16749 (N_16749,N_12683,N_13313);
nand U16750 (N_16750,N_12328,N_11463);
xor U16751 (N_16751,N_14526,N_13539);
nor U16752 (N_16752,N_13591,N_11165);
xor U16753 (N_16753,N_10182,N_13723);
nor U16754 (N_16754,N_11964,N_13893);
nor U16755 (N_16755,N_14747,N_12013);
and U16756 (N_16756,N_14793,N_13249);
or U16757 (N_16757,N_14817,N_13294);
or U16758 (N_16758,N_13379,N_11485);
nand U16759 (N_16759,N_13653,N_11286);
nor U16760 (N_16760,N_13911,N_11726);
nor U16761 (N_16761,N_14552,N_13259);
and U16762 (N_16762,N_12989,N_10233);
or U16763 (N_16763,N_14202,N_13308);
or U16764 (N_16764,N_12369,N_10281);
and U16765 (N_16765,N_10167,N_14347);
nor U16766 (N_16766,N_13034,N_11341);
and U16767 (N_16767,N_12675,N_14554);
xnor U16768 (N_16768,N_13094,N_12567);
xnor U16769 (N_16769,N_10006,N_10197);
nand U16770 (N_16770,N_13182,N_11575);
xor U16771 (N_16771,N_14567,N_13635);
nor U16772 (N_16772,N_12208,N_10631);
xnor U16773 (N_16773,N_12119,N_14509);
nand U16774 (N_16774,N_13186,N_11625);
nor U16775 (N_16775,N_10353,N_13097);
xnor U16776 (N_16776,N_12847,N_12361);
nand U16777 (N_16777,N_13927,N_14786);
or U16778 (N_16778,N_11369,N_10401);
or U16779 (N_16779,N_14596,N_14638);
nor U16780 (N_16780,N_10439,N_13264);
nor U16781 (N_16781,N_12717,N_14910);
xnor U16782 (N_16782,N_10584,N_14580);
and U16783 (N_16783,N_12947,N_14767);
or U16784 (N_16784,N_12469,N_14274);
and U16785 (N_16785,N_13483,N_12359);
nor U16786 (N_16786,N_14133,N_10284);
xnor U16787 (N_16787,N_11062,N_12236);
xnor U16788 (N_16788,N_11879,N_13753);
and U16789 (N_16789,N_14701,N_10087);
nand U16790 (N_16790,N_14798,N_14656);
and U16791 (N_16791,N_10205,N_11803);
xnor U16792 (N_16792,N_12272,N_13471);
nor U16793 (N_16793,N_12045,N_10817);
nor U16794 (N_16794,N_14897,N_14794);
nand U16795 (N_16795,N_13845,N_12510);
or U16796 (N_16796,N_13799,N_14711);
nor U16797 (N_16797,N_12921,N_11765);
nand U16798 (N_16798,N_10031,N_11431);
or U16799 (N_16799,N_14282,N_10470);
or U16800 (N_16800,N_11477,N_11229);
or U16801 (N_16801,N_13822,N_13895);
xnor U16802 (N_16802,N_12110,N_14459);
nand U16803 (N_16803,N_10427,N_12450);
nor U16804 (N_16804,N_12410,N_10833);
or U16805 (N_16805,N_12641,N_11320);
and U16806 (N_16806,N_13490,N_12160);
nor U16807 (N_16807,N_10609,N_10065);
or U16808 (N_16808,N_11183,N_13455);
xor U16809 (N_16809,N_10294,N_14251);
xor U16810 (N_16810,N_12545,N_13738);
nor U16811 (N_16811,N_12396,N_11296);
nor U16812 (N_16812,N_14732,N_14535);
xnor U16813 (N_16813,N_14556,N_12135);
nor U16814 (N_16814,N_12349,N_10814);
nor U16815 (N_16815,N_12888,N_12643);
and U16816 (N_16816,N_12436,N_10287);
and U16817 (N_16817,N_11936,N_13335);
xnor U16818 (N_16818,N_10912,N_11876);
or U16819 (N_16819,N_10837,N_10663);
nor U16820 (N_16820,N_11364,N_14797);
and U16821 (N_16821,N_14375,N_14207);
nor U16822 (N_16822,N_13062,N_14264);
or U16823 (N_16823,N_12483,N_11483);
nor U16824 (N_16824,N_12790,N_12874);
and U16825 (N_16825,N_11976,N_14042);
and U16826 (N_16826,N_14548,N_12593);
nor U16827 (N_16827,N_11563,N_13908);
nor U16828 (N_16828,N_14965,N_14835);
xnor U16829 (N_16829,N_11280,N_14867);
and U16830 (N_16830,N_11034,N_11390);
nand U16831 (N_16831,N_10987,N_10232);
xnor U16832 (N_16832,N_10726,N_14561);
and U16833 (N_16833,N_10326,N_13153);
nand U16834 (N_16834,N_14064,N_13854);
nand U16835 (N_16835,N_14082,N_12743);
xor U16836 (N_16836,N_14161,N_12618);
and U16837 (N_16837,N_11247,N_12262);
and U16838 (N_16838,N_10937,N_14361);
nand U16839 (N_16839,N_10821,N_11479);
or U16840 (N_16840,N_13119,N_12415);
and U16841 (N_16841,N_11539,N_11220);
nand U16842 (N_16842,N_14850,N_11622);
and U16843 (N_16843,N_13369,N_13441);
or U16844 (N_16844,N_10433,N_13015);
or U16845 (N_16845,N_10965,N_11271);
nor U16846 (N_16846,N_13556,N_11061);
nand U16847 (N_16847,N_13645,N_14655);
or U16848 (N_16848,N_13874,N_14472);
nand U16849 (N_16849,N_11285,N_10627);
nor U16850 (N_16850,N_13371,N_10190);
and U16851 (N_16851,N_11409,N_13607);
nand U16852 (N_16852,N_12880,N_12650);
nand U16853 (N_16853,N_11264,N_14520);
nor U16854 (N_16854,N_14154,N_14515);
xor U16855 (N_16855,N_13012,N_10300);
nand U16856 (N_16856,N_12704,N_13746);
nor U16857 (N_16857,N_10876,N_13160);
or U16858 (N_16858,N_10201,N_13330);
nand U16859 (N_16859,N_13619,N_14417);
or U16860 (N_16860,N_11008,N_13427);
nor U16861 (N_16861,N_10626,N_14678);
or U16862 (N_16862,N_12724,N_13185);
xnor U16863 (N_16863,N_10450,N_12532);
or U16864 (N_16864,N_12958,N_13109);
nand U16865 (N_16865,N_10400,N_10750);
or U16866 (N_16866,N_10651,N_14330);
nor U16867 (N_16867,N_10196,N_14204);
xor U16868 (N_16868,N_11267,N_10017);
or U16869 (N_16869,N_11418,N_11657);
and U16870 (N_16870,N_11287,N_11653);
xor U16871 (N_16871,N_12339,N_14558);
nand U16872 (N_16872,N_13603,N_13912);
and U16873 (N_16873,N_12082,N_11796);
nor U16874 (N_16874,N_12094,N_10950);
nor U16875 (N_16875,N_10436,N_13864);
xnor U16876 (N_16876,N_14943,N_12614);
or U16877 (N_16877,N_14606,N_11424);
nor U16878 (N_16878,N_11632,N_11744);
xnor U16879 (N_16879,N_14238,N_14512);
and U16880 (N_16880,N_11495,N_12021);
xor U16881 (N_16881,N_11821,N_11692);
or U16882 (N_16882,N_11986,N_11984);
or U16883 (N_16883,N_10295,N_14705);
or U16884 (N_16884,N_11234,N_14928);
and U16885 (N_16885,N_11761,N_12587);
nand U16886 (N_16886,N_13888,N_10280);
nor U16887 (N_16887,N_13380,N_13932);
nor U16888 (N_16888,N_12177,N_10666);
nand U16889 (N_16889,N_11781,N_11491);
or U16890 (N_16890,N_11616,N_14597);
nor U16891 (N_16891,N_13870,N_11800);
nor U16892 (N_16892,N_12554,N_12815);
xnor U16893 (N_16893,N_12313,N_11470);
nor U16894 (N_16894,N_10708,N_10373);
and U16895 (N_16895,N_13513,N_11776);
and U16896 (N_16896,N_12053,N_11447);
and U16897 (N_16897,N_12276,N_10764);
xnor U16898 (N_16898,N_13520,N_10100);
or U16899 (N_16899,N_11708,N_11922);
nand U16900 (N_16900,N_10703,N_11350);
and U16901 (N_16901,N_11269,N_13777);
nor U16902 (N_16902,N_13302,N_12465);
nand U16903 (N_16903,N_12986,N_12948);
and U16904 (N_16904,N_13721,N_14176);
nand U16905 (N_16905,N_12960,N_14246);
or U16906 (N_16906,N_13323,N_11798);
or U16907 (N_16907,N_11050,N_11102);
nor U16908 (N_16908,N_14924,N_14861);
nand U16909 (N_16909,N_12209,N_10915);
nor U16910 (N_16910,N_10760,N_14386);
or U16911 (N_16911,N_10453,N_12220);
nor U16912 (N_16912,N_14752,N_13131);
xor U16913 (N_16913,N_12603,N_13013);
or U16914 (N_16914,N_13924,N_11849);
or U16915 (N_16915,N_13166,N_12756);
or U16916 (N_16916,N_14918,N_11591);
nor U16917 (N_16917,N_13019,N_10474);
nand U16918 (N_16918,N_13320,N_13530);
nand U16919 (N_16919,N_13227,N_13589);
nand U16920 (N_16920,N_10611,N_13014);
nor U16921 (N_16921,N_10118,N_14475);
nand U16922 (N_16922,N_14658,N_11754);
or U16923 (N_16923,N_14159,N_14111);
or U16924 (N_16924,N_10155,N_13305);
nand U16925 (N_16925,N_13651,N_11523);
nor U16926 (N_16926,N_12199,N_10218);
and U16927 (N_16927,N_14344,N_13325);
nor U16928 (N_16928,N_11811,N_10239);
and U16929 (N_16929,N_10713,N_12147);
nand U16930 (N_16930,N_13985,N_13446);
xor U16931 (N_16931,N_10559,N_13124);
or U16932 (N_16932,N_13444,N_13903);
nand U16933 (N_16933,N_11675,N_12913);
or U16934 (N_16934,N_10655,N_13547);
nand U16935 (N_16935,N_12499,N_12706);
and U16936 (N_16936,N_12995,N_11411);
and U16937 (N_16937,N_10761,N_11905);
nand U16938 (N_16938,N_12433,N_12890);
or U16939 (N_16939,N_14939,N_13525);
xnor U16940 (N_16940,N_10578,N_12442);
or U16941 (N_16941,N_12425,N_13236);
or U16942 (N_16942,N_12979,N_11930);
nand U16943 (N_16943,N_12548,N_10585);
and U16944 (N_16944,N_14981,N_11140);
nand U16945 (N_16945,N_13037,N_10223);
nor U16946 (N_16946,N_11934,N_10379);
and U16947 (N_16947,N_12235,N_13846);
xnor U16948 (N_16948,N_11667,N_12430);
nand U16949 (N_16949,N_13829,N_13731);
nor U16950 (N_16950,N_12723,N_12833);
or U16951 (N_16951,N_10781,N_12696);
xor U16952 (N_16952,N_14382,N_14906);
nand U16953 (N_16953,N_12411,N_14676);
and U16954 (N_16954,N_10728,N_11057);
and U16955 (N_16955,N_13519,N_12621);
nor U16956 (N_16956,N_11353,N_14719);
or U16957 (N_16957,N_14713,N_10961);
nand U16958 (N_16958,N_10238,N_10894);
xnor U16959 (N_16959,N_12228,N_11457);
xor U16960 (N_16960,N_10542,N_14570);
and U16961 (N_16961,N_14822,N_12071);
or U16962 (N_16962,N_10800,N_11357);
nor U16963 (N_16963,N_14089,N_10176);
or U16964 (N_16964,N_13472,N_11075);
nand U16965 (N_16965,N_10898,N_10594);
or U16966 (N_16966,N_14120,N_10701);
xor U16967 (N_16967,N_11649,N_11818);
xor U16968 (N_16968,N_14671,N_11564);
xnor U16969 (N_16969,N_14814,N_13616);
xnor U16970 (N_16970,N_11923,N_13450);
nand U16971 (N_16971,N_14654,N_11449);
or U16972 (N_16972,N_11912,N_11045);
xor U16973 (N_16973,N_13202,N_12925);
xor U16974 (N_16974,N_12518,N_14327);
nand U16975 (N_16975,N_12875,N_12125);
and U16976 (N_16976,N_14185,N_14352);
and U16977 (N_16977,N_10555,N_11289);
nand U16978 (N_16978,N_13005,N_13849);
and U16979 (N_16979,N_14807,N_14862);
nand U16980 (N_16980,N_14560,N_13509);
nand U16981 (N_16981,N_13234,N_10461);
or U16982 (N_16982,N_11086,N_11446);
and U16983 (N_16983,N_13039,N_13267);
nand U16984 (N_16984,N_11120,N_13029);
nand U16985 (N_16985,N_11372,N_10046);
and U16986 (N_16986,N_11055,N_12615);
and U16987 (N_16987,N_13693,N_14024);
or U16988 (N_16988,N_13949,N_12843);
nand U16989 (N_16989,N_14972,N_14818);
nor U16990 (N_16990,N_14664,N_12971);
xor U16991 (N_16991,N_11703,N_14628);
xnor U16992 (N_16992,N_11552,N_10033);
nand U16993 (N_16993,N_12850,N_14139);
and U16994 (N_16994,N_11135,N_14340);
or U16995 (N_16995,N_12172,N_11548);
nand U16996 (N_16996,N_12799,N_11121);
nand U16997 (N_16997,N_10752,N_11127);
nor U16998 (N_16998,N_14771,N_14831);
xnor U16999 (N_16999,N_10721,N_14412);
nor U17000 (N_17000,N_14305,N_10411);
nor U17001 (N_17001,N_12083,N_14610);
nand U17002 (N_17002,N_12167,N_11973);
nand U17003 (N_17003,N_12528,N_14167);
nand U17004 (N_17004,N_12398,N_13385);
nor U17005 (N_17005,N_10275,N_12478);
nor U17006 (N_17006,N_13671,N_12678);
and U17007 (N_17007,N_13766,N_13931);
or U17008 (N_17008,N_12825,N_12975);
nor U17009 (N_17009,N_11175,N_11945);
nor U17010 (N_17010,N_10674,N_13926);
or U17011 (N_17011,N_10063,N_10352);
nor U17012 (N_17012,N_13229,N_10246);
nand U17013 (N_17013,N_14171,N_13176);
and U17014 (N_17014,N_14479,N_14994);
or U17015 (N_17015,N_14662,N_13706);
nor U17016 (N_17016,N_14010,N_13809);
nor U17017 (N_17017,N_10906,N_11638);
and U17018 (N_17018,N_12936,N_14681);
and U17019 (N_17019,N_11833,N_13995);
nor U17020 (N_17020,N_13066,N_10331);
and U17021 (N_17021,N_10508,N_12259);
or U17022 (N_17022,N_11869,N_12838);
nand U17023 (N_17023,N_13424,N_14395);
nand U17024 (N_17024,N_10715,N_13983);
xor U17025 (N_17025,N_14439,N_12019);
or U17026 (N_17026,N_13610,N_14191);
and U17027 (N_17027,N_13637,N_14546);
or U17028 (N_17028,N_12214,N_14858);
or U17029 (N_17029,N_14815,N_12574);
and U17030 (N_17030,N_13216,N_10241);
xnor U17031 (N_17031,N_10593,N_11459);
and U17032 (N_17032,N_12677,N_11056);
nor U17033 (N_17033,N_10515,N_11952);
nor U17034 (N_17034,N_11810,N_13357);
xor U17035 (N_17035,N_11099,N_14677);
and U17036 (N_17036,N_10512,N_12703);
or U17037 (N_17037,N_12930,N_10998);
nor U17038 (N_17038,N_13443,N_12994);
nand U17039 (N_17039,N_11227,N_10644);
or U17040 (N_17040,N_12942,N_10264);
nor U17041 (N_17041,N_11516,N_10296);
nand U17042 (N_17042,N_14401,N_11941);
and U17043 (N_17043,N_11540,N_12025);
nand U17044 (N_17044,N_13502,N_13148);
xor U17045 (N_17045,N_14741,N_12586);
xor U17046 (N_17046,N_14286,N_12397);
and U17047 (N_17047,N_12760,N_13958);
nand U17048 (N_17048,N_13580,N_14408);
nand U17049 (N_17049,N_12968,N_12202);
nand U17050 (N_17050,N_12288,N_11359);
xor U17051 (N_17051,N_11033,N_13045);
nor U17052 (N_17052,N_14326,N_14002);
xor U17053 (N_17053,N_12774,N_13310);
or U17054 (N_17054,N_12613,N_13886);
or U17055 (N_17055,N_11071,N_14997);
nor U17056 (N_17056,N_14249,N_12004);
xor U17057 (N_17057,N_12978,N_13462);
nand U17058 (N_17058,N_12515,N_12770);
and U17059 (N_17059,N_11130,N_13684);
and U17060 (N_17060,N_14645,N_11757);
nor U17061 (N_17061,N_11596,N_14212);
nor U17062 (N_17062,N_11308,N_14483);
nand U17063 (N_17063,N_13363,N_12780);
or U17064 (N_17064,N_10483,N_14078);
xnor U17065 (N_17065,N_12575,N_10090);
or U17066 (N_17066,N_10688,N_14201);
or U17067 (N_17067,N_13338,N_10189);
nor U17068 (N_17068,N_14745,N_14882);
and U17069 (N_17069,N_13514,N_13167);
nor U17070 (N_17070,N_10944,N_14648);
nor U17071 (N_17071,N_13674,N_10410);
nor U17072 (N_17072,N_14151,N_10824);
or U17073 (N_17073,N_11559,N_14080);
nand U17074 (N_17074,N_13800,N_14445);
and U17075 (N_17075,N_12344,N_13945);
and U17076 (N_17076,N_12332,N_10600);
nor U17077 (N_17077,N_11787,N_14885);
nand U17078 (N_17078,N_11314,N_13196);
nor U17079 (N_17079,N_11740,N_10573);
or U17080 (N_17080,N_11730,N_12751);
or U17081 (N_17081,N_10148,N_14104);
and U17082 (N_17082,N_11804,N_14860);
nand U17083 (N_17083,N_13943,N_13058);
nand U17084 (N_17084,N_12648,N_14444);
and U17085 (N_17085,N_13278,N_11448);
nor U17086 (N_17086,N_12222,N_14241);
or U17087 (N_17087,N_14168,N_11337);
xnor U17088 (N_17088,N_14666,N_13372);
xor U17089 (N_17089,N_11903,N_14955);
and U17090 (N_17090,N_14130,N_13585);
nand U17091 (N_17091,N_11284,N_12789);
xnor U17092 (N_17092,N_10339,N_12594);
and U17093 (N_17093,N_14776,N_10856);
or U17094 (N_17094,N_12931,N_10174);
xor U17095 (N_17095,N_13137,N_12223);
nor U17096 (N_17096,N_14306,N_12543);
nand U17097 (N_17097,N_11627,N_10108);
or U17098 (N_17098,N_14736,N_10151);
or U17099 (N_17099,N_14673,N_11486);
and U17100 (N_17100,N_11681,N_13276);
and U17101 (N_17101,N_11792,N_11999);
nand U17102 (N_17102,N_12018,N_10367);
nand U17103 (N_17103,N_12727,N_12294);
nor U17104 (N_17104,N_14275,N_11786);
and U17105 (N_17105,N_11609,N_14625);
and U17106 (N_17106,N_14485,N_11883);
and U17107 (N_17107,N_12573,N_12681);
nor U17108 (N_17108,N_11301,N_13704);
and U17109 (N_17109,N_11098,N_10492);
and U17110 (N_17110,N_11015,N_14743);
nor U17111 (N_17111,N_14911,N_12017);
nor U17112 (N_17112,N_10751,N_10388);
nor U17113 (N_17113,N_11232,N_12367);
xor U17114 (N_17114,N_11688,N_14513);
nor U17115 (N_17115,N_12776,N_10532);
nand U17116 (N_17116,N_13461,N_13920);
nand U17117 (N_17117,N_11600,N_12820);
xnor U17118 (N_17118,N_13698,N_11489);
nand U17119 (N_17119,N_11772,N_10123);
or U17120 (N_17120,N_13098,N_12270);
nand U17121 (N_17121,N_13362,N_14044);
and U17122 (N_17122,N_12668,N_13430);
nor U17123 (N_17123,N_10494,N_11170);
nand U17124 (N_17124,N_11642,N_11807);
nand U17125 (N_17125,N_11025,N_13347);
and U17126 (N_17126,N_10743,N_12490);
and U17127 (N_17127,N_11414,N_12831);
or U17128 (N_17128,N_13989,N_10834);
xnor U17129 (N_17129,N_11528,N_11782);
xnor U17130 (N_17130,N_10667,N_13638);
xor U17131 (N_17131,N_11374,N_12623);
xor U17132 (N_17132,N_12694,N_10509);
nor U17133 (N_17133,N_11235,N_12737);
nor U17134 (N_17134,N_12162,N_12578);
nor U17135 (N_17135,N_14446,N_11916);
nand U17136 (N_17136,N_12102,N_14057);
xnor U17137 (N_17137,N_10180,N_13373);
or U17138 (N_17138,N_10012,N_10843);
and U17139 (N_17139,N_14702,N_12114);
nor U17140 (N_17140,N_12909,N_12350);
xor U17141 (N_17141,N_11303,N_10417);
or U17142 (N_17142,N_13916,N_10528);
nor U17143 (N_17143,N_11522,N_11328);
or U17144 (N_17144,N_13582,N_13155);
nand U17145 (N_17145,N_11327,N_14494);
xor U17146 (N_17146,N_10697,N_10029);
or U17147 (N_17147,N_13899,N_12474);
or U17148 (N_17148,N_14279,N_11294);
nand U17149 (N_17149,N_13203,N_10682);
xor U17150 (N_17150,N_10307,N_13134);
xnor U17151 (N_17151,N_13291,N_11715);
and U17152 (N_17152,N_11213,N_12795);
nand U17153 (N_17153,N_12322,N_10093);
xor U17154 (N_17154,N_11354,N_13687);
and U17155 (N_17155,N_10597,N_11136);
nand U17156 (N_17156,N_10082,N_12289);
or U17157 (N_17157,N_12335,N_10679);
nand U17158 (N_17158,N_11049,N_12951);
nor U17159 (N_17159,N_14214,N_13715);
or U17160 (N_17160,N_10829,N_10786);
or U17161 (N_17161,N_12985,N_11508);
or U17162 (N_17162,N_10088,N_12310);
and U17163 (N_17163,N_14419,N_12550);
xor U17164 (N_17164,N_10178,N_13337);
and U17165 (N_17165,N_14834,N_10926);
nor U17166 (N_17166,N_10355,N_11979);
nand U17167 (N_17167,N_12713,N_12244);
xor U17168 (N_17168,N_12357,N_12882);
nand U17169 (N_17169,N_14593,N_12031);
or U17170 (N_17170,N_11844,N_14328);
or U17171 (N_17171,N_11210,N_13223);
and U17172 (N_17172,N_13195,N_12876);
nor U17173 (N_17173,N_12551,N_11077);
and U17174 (N_17174,N_11921,N_12631);
and U17175 (N_17175,N_14543,N_10522);
and U17176 (N_17176,N_14650,N_14774);
or U17177 (N_17177,N_10160,N_11687);
xnor U17178 (N_17178,N_14087,N_11861);
nor U17179 (N_17179,N_11894,N_14739);
nor U17180 (N_17180,N_12507,N_13112);
xnor U17181 (N_17181,N_12459,N_13930);
nand U17182 (N_17182,N_14507,N_10162);
nand U17183 (N_17183,N_10560,N_11779);
or U17184 (N_17184,N_11808,N_11541);
nand U17185 (N_17185,N_14290,N_10874);
and U17186 (N_17186,N_12637,N_10639);
and U17187 (N_17187,N_12154,N_10324);
or U17188 (N_17188,N_13150,N_12484);
and U17189 (N_17189,N_12902,N_13601);
nor U17190 (N_17190,N_13821,N_12446);
and U17191 (N_17191,N_13618,N_12984);
nor U17192 (N_17192,N_13718,N_14864);
or U17193 (N_17193,N_11069,N_10854);
nand U17194 (N_17194,N_12887,N_10538);
or U17195 (N_17195,N_14333,N_14450);
nand U17196 (N_17196,N_10332,N_10994);
or U17197 (N_17197,N_14463,N_12939);
or U17198 (N_17198,N_12610,N_11295);
nand U17199 (N_17199,N_10908,N_13475);
nor U17200 (N_17200,N_11481,N_13061);
and U17201 (N_17201,N_14491,N_12370);
nor U17202 (N_17202,N_13935,N_10442);
nor U17203 (N_17203,N_11562,N_14335);
or U17204 (N_17204,N_11747,N_13986);
nor U17205 (N_17205,N_14929,N_11236);
nand U17206 (N_17206,N_12158,N_11397);
or U17207 (N_17207,N_12241,N_12786);
and U17208 (N_17208,N_13588,N_11666);
or U17209 (N_17209,N_13652,N_10753);
and U17210 (N_17210,N_10251,N_11824);
nor U17211 (N_17211,N_10161,N_12286);
nand U17212 (N_17212,N_11028,N_10079);
xnor U17213 (N_17213,N_14725,N_13538);
nand U17214 (N_17214,N_14127,N_11081);
or U17215 (N_17215,N_13526,N_12690);
and U17216 (N_17216,N_13188,N_11718);
nand U17217 (N_17217,N_11274,N_14265);
or U17218 (N_17218,N_10004,N_10778);
nand U17219 (N_17219,N_13819,N_10827);
nor U17220 (N_17220,N_12261,N_11466);
nor U17221 (N_17221,N_11147,N_13555);
or U17222 (N_17222,N_14529,N_10242);
or U17223 (N_17223,N_14632,N_10940);
nor U17224 (N_17224,N_14174,N_10680);
nor U17225 (N_17225,N_10337,N_14870);
nand U17226 (N_17226,N_11890,N_13333);
and U17227 (N_17227,N_12492,N_14248);
or U17228 (N_17228,N_12652,N_10303);
or U17229 (N_17229,N_14019,N_14046);
nand U17230 (N_17230,N_11307,N_11206);
or U17231 (N_17231,N_13474,N_12802);
and U17232 (N_17232,N_10737,N_14160);
xnor U17233 (N_17233,N_14289,N_12599);
or U17234 (N_17234,N_11770,N_11380);
and U17235 (N_17235,N_10368,N_12479);
or U17236 (N_17236,N_11723,N_12867);
nor U17237 (N_17237,N_10879,N_12733);
nor U17238 (N_17238,N_12133,N_14586);
xnor U17239 (N_17239,N_12429,N_11410);
and U17240 (N_17240,N_10977,N_14410);
nand U17241 (N_17241,N_13739,N_11490);
or U17242 (N_17242,N_11762,N_13048);
nor U17243 (N_17243,N_10523,N_12027);
xnor U17244 (N_17244,N_11219,N_10670);
nor U17245 (N_17245,N_13106,N_11822);
xnor U17246 (N_17246,N_12509,N_11309);
nand U17247 (N_17247,N_10936,N_11396);
nor U17248 (N_17248,N_11261,N_11388);
xnor U17249 (N_17249,N_10572,N_14015);
or U17250 (N_17250,N_10598,N_14081);
nand U17251 (N_17251,N_14722,N_10527);
nor U17252 (N_17252,N_10702,N_12340);
xnor U17253 (N_17253,N_14117,N_12443);
nand U17254 (N_17254,N_14030,N_12633);
nand U17255 (N_17255,N_12173,N_10992);
nand U17256 (N_17256,N_12070,N_11412);
nand U17257 (N_17257,N_14605,N_13011);
or U17258 (N_17258,N_11141,N_14427);
nand U17259 (N_17259,N_10549,N_10259);
nand U17260 (N_17260,N_10901,N_11684);
nand U17261 (N_17261,N_12796,N_10842);
xnor U17262 (N_17262,N_10722,N_13077);
or U17263 (N_17263,N_12153,N_13708);
and U17264 (N_17264,N_11668,N_14537);
and U17265 (N_17265,N_13107,N_12277);
nand U17266 (N_17266,N_13909,N_14874);
xor U17267 (N_17267,N_13685,N_11173);
and U17268 (N_17268,N_12644,N_13010);
and U17269 (N_17269,N_11764,N_12293);
nand U17270 (N_17270,N_12646,N_10656);
nand U17271 (N_17271,N_10654,N_13110);
xor U17272 (N_17272,N_12663,N_14242);
nor U17273 (N_17273,N_11931,N_10449);
nor U17274 (N_17274,N_12977,N_14049);
and U17275 (N_17275,N_14126,N_12781);
xor U17276 (N_17276,N_14948,N_13274);
and U17277 (N_17277,N_14869,N_12260);
nor U17278 (N_17278,N_10783,N_11951);
and U17279 (N_17279,N_14759,N_10216);
xor U17280 (N_17280,N_13791,N_13477);
xor U17281 (N_17281,N_11924,N_12565);
nor U17282 (N_17282,N_13950,N_13826);
xor U17283 (N_17283,N_14865,N_12519);
xor U17284 (N_17284,N_10772,N_13395);
xnor U17285 (N_17285,N_11259,N_10447);
and U17286 (N_17286,N_14467,N_12159);
xnor U17287 (N_17287,N_11603,N_14436);
nor U17288 (N_17288,N_10607,N_13677);
xnor U17289 (N_17289,N_12185,N_11092);
nand U17290 (N_17290,N_13104,N_11167);
nor U17291 (N_17291,N_13823,N_14198);
and U17292 (N_17292,N_11244,N_11753);
nor U17293 (N_17293,N_14881,N_14602);
and U17294 (N_17294,N_10382,N_13036);
nor U17295 (N_17295,N_10434,N_13956);
or U17296 (N_17296,N_12892,N_14590);
nor U17297 (N_17297,N_14840,N_11407);
xor U17298 (N_17298,N_13796,N_10198);
and U17299 (N_17299,N_10826,N_14428);
nor U17300 (N_17300,N_11119,N_10277);
nor U17301 (N_17301,N_13577,N_13934);
xnor U17302 (N_17302,N_13258,N_14753);
nor U17303 (N_17303,N_12416,N_12365);
nand U17304 (N_17304,N_11846,N_10740);
nand U17305 (N_17305,N_10577,N_12020);
nor U17306 (N_17306,N_13964,N_13815);
nor U17307 (N_17307,N_14458,N_12034);
or U17308 (N_17308,N_13787,N_13453);
nand U17309 (N_17309,N_11948,N_11366);
or U17310 (N_17310,N_10782,N_14079);
nor U17311 (N_17311,N_14070,N_14744);
nand U17312 (N_17312,N_10648,N_13537);
xnor U17313 (N_17313,N_13656,N_13981);
nor U17314 (N_17314,N_14339,N_13625);
xnor U17315 (N_17315,N_12687,N_11073);
or U17316 (N_17316,N_10687,N_11955);
nand U17317 (N_17317,N_10265,N_10107);
nand U17318 (N_17318,N_13648,N_11977);
or U17319 (N_17319,N_14138,N_13884);
nor U17320 (N_17320,N_10026,N_14842);
or U17321 (N_17321,N_14048,N_11961);
and U17322 (N_17322,N_13408,N_13961);
or U17323 (N_17323,N_12258,N_13463);
or U17324 (N_17324,N_10422,N_11011);
or U17325 (N_17325,N_13602,N_10984);
nand U17326 (N_17326,N_12267,N_11031);
xor U17327 (N_17327,N_14680,N_10868);
nor U17328 (N_17328,N_10789,N_10976);
and U17329 (N_17329,N_11482,N_10113);
xnor U17330 (N_17330,N_14970,N_13466);
nor U17331 (N_17331,N_11882,N_14370);
and U17332 (N_17332,N_14859,N_14103);
nand U17333 (N_17333,N_12725,N_10060);
nor U17334 (N_17334,N_10144,N_10459);
xor U17335 (N_17335,N_14311,N_10211);
nand U17336 (N_17336,N_13351,N_14209);
or U17337 (N_17337,N_13902,N_10413);
nand U17338 (N_17338,N_12626,N_10613);
nand U17339 (N_17339,N_10769,N_11283);
or U17340 (N_17340,N_12664,N_11648);
xnor U17341 (N_17341,N_14179,N_11079);
nand U17342 (N_17342,N_11728,N_13452);
xor U17343 (N_17343,N_12910,N_14740);
and U17344 (N_17344,N_13409,N_14217);
nor U17345 (N_17345,N_13402,N_12077);
xor U17346 (N_17346,N_14971,N_14190);
xnor U17347 (N_17347,N_12036,N_14791);
or U17348 (N_17348,N_12201,N_11680);
and U17349 (N_17349,N_13967,N_12380);
nand U17350 (N_17350,N_11733,N_10848);
nand U17351 (N_17351,N_11918,N_13918);
nor U17352 (N_17352,N_13546,N_12691);
nor U17353 (N_17353,N_10024,N_13838);
nor U17354 (N_17354,N_13661,N_12605);
and U17355 (N_17355,N_14037,N_10933);
nor U17356 (N_17356,N_10794,N_13612);
nand U17357 (N_17357,N_11722,N_11929);
nand U17358 (N_17358,N_11678,N_12408);
or U17359 (N_17359,N_13668,N_13273);
nand U17360 (N_17360,N_11560,N_12834);
xor U17361 (N_17361,N_12390,N_14356);
or U17362 (N_17362,N_11030,N_14158);
nand U17363 (N_17363,N_14380,N_12714);
nand U17364 (N_17364,N_11172,N_13146);
xnor U17365 (N_17365,N_12784,N_13641);
or U17366 (N_17366,N_14325,N_14754);
and U17367 (N_17367,N_10497,N_10414);
nor U17368 (N_17368,N_12538,N_14846);
nand U17369 (N_17369,N_13420,N_10982);
and U17370 (N_17370,N_14240,N_12803);
xor U17371 (N_17371,N_13810,N_12320);
or U17372 (N_17372,N_12726,N_10454);
or U17373 (N_17373,N_11176,N_14959);
nor U17374 (N_17374,N_11352,N_12326);
xnor U17375 (N_17375,N_12376,N_13658);
nor U17376 (N_17376,N_12239,N_12590);
or U17377 (N_17377,N_11106,N_10286);
or U17378 (N_17378,N_12355,N_14998);
nor U17379 (N_17379,N_13804,N_13737);
nand U17380 (N_17380,N_10973,N_11672);
or U17381 (N_17381,N_13198,N_10053);
nand U17382 (N_17382,N_14812,N_11292);
and U17383 (N_17383,N_12404,N_13031);
xor U17384 (N_17384,N_11453,N_13319);
nor U17385 (N_17385,N_14516,N_11066);
or U17386 (N_17386,N_10861,N_14318);
or U17387 (N_17387,N_10356,N_13858);
nand U17388 (N_17388,N_11615,N_12377);
nor U17389 (N_17389,N_10435,N_10850);
nor U17390 (N_17390,N_13352,N_14790);
or U17391 (N_17391,N_12281,N_10094);
nor U17392 (N_17392,N_14684,N_10344);
or U17393 (N_17393,N_12818,N_11574);
xnor U17394 (N_17394,N_10109,N_14985);
xor U17395 (N_17395,N_10479,N_14123);
nand U17396 (N_17396,N_12872,N_14388);
or U17397 (N_17397,N_11790,N_11002);
or U17398 (N_17398,N_11224,N_13208);
xor U17399 (N_17399,N_11306,N_12476);
or U17400 (N_17400,N_14150,N_12993);
or U17401 (N_17401,N_10059,N_12617);
and U17402 (N_17402,N_11000,N_14763);
nor U17403 (N_17403,N_12660,N_14663);
or U17404 (N_17404,N_14504,N_13891);
and U17405 (N_17405,N_11010,N_10208);
nand U17406 (N_17406,N_12282,N_12317);
nand U17407 (N_17407,N_14196,N_12667);
xnor U17408 (N_17408,N_12849,N_11891);
nand U17409 (N_17409,N_10500,N_10200);
or U17410 (N_17410,N_12181,N_12012);
or U17411 (N_17411,N_14466,N_12418);
or U17412 (N_17412,N_12582,N_14640);
xor U17413 (N_17413,N_12903,N_12769);
xor U17414 (N_17414,N_13863,N_10812);
or U17415 (N_17415,N_13168,N_13105);
and U17416 (N_17416,N_13790,N_12823);
or U17417 (N_17417,N_11345,N_12467);
nand U17418 (N_17418,N_10660,N_14578);
xor U17419 (N_17419,N_14189,N_10658);
and U17420 (N_17420,N_10163,N_14004);
nor U17421 (N_17421,N_10774,N_13091);
or U17422 (N_17422,N_11953,N_14293);
xnor U17423 (N_17423,N_14298,N_12580);
nor U17424 (N_17424,N_10798,N_11624);
and U17425 (N_17425,N_12128,N_12195);
nor U17426 (N_17426,N_13560,N_14637);
xor U17427 (N_17427,N_10070,N_13040);
xor U17428 (N_17428,N_13221,N_12999);
xnor U17429 (N_17429,N_14940,N_12943);
nor U17430 (N_17430,N_10212,N_14839);
nand U17431 (N_17431,N_11044,N_13524);
xnor U17432 (N_17432,N_14703,N_13388);
xnor U17433 (N_17433,N_14172,N_11493);
xor U17434 (N_17434,N_14413,N_10273);
nor U17435 (N_17435,N_14731,N_10758);
xor U17436 (N_17436,N_10970,N_14931);
or U17437 (N_17437,N_10534,N_14565);
nor U17438 (N_17438,N_10504,N_13263);
nand U17439 (N_17439,N_11419,N_10119);
or U17440 (N_17440,N_10923,N_10756);
or U17441 (N_17441,N_12343,N_11404);
xor U17442 (N_17442,N_13419,N_10157);
nand U17443 (N_17443,N_13122,N_12434);
or U17444 (N_17444,N_14090,N_11676);
or U17445 (N_17445,N_13776,N_12035);
and U17446 (N_17446,N_12851,N_14825);
or U17447 (N_17447,N_13233,N_10179);
xnor U17448 (N_17448,N_14524,N_14508);
xnor U17449 (N_17449,N_11451,N_14781);
nor U17450 (N_17450,N_13764,N_12375);
or U17451 (N_17451,N_13872,N_13399);
nand U17452 (N_17452,N_14454,N_12319);
or U17453 (N_17453,N_10227,N_11145);
xor U17454 (N_17454,N_10228,N_12306);
xnor U17455 (N_17455,N_10472,N_11794);
and U17456 (N_17456,N_12445,N_13467);
and U17457 (N_17457,N_11946,N_13479);
xnor U17458 (N_17458,N_12048,N_11584);
xnor U17459 (N_17459,N_14065,N_12141);
and U17460 (N_17460,N_10780,N_10011);
nor U17461 (N_17461,N_12881,N_12809);
nand U17462 (N_17462,N_10553,N_11897);
xor U17463 (N_17463,N_12122,N_11275);
xnor U17464 (N_17464,N_10357,N_12766);
and U17465 (N_17465,N_11738,N_11426);
and U17466 (N_17466,N_11778,N_10360);
xor U17467 (N_17467,N_14783,N_13760);
or U17468 (N_17468,N_12087,N_14337);
nand U17469 (N_17469,N_11633,N_10404);
or U17470 (N_17470,N_13771,N_13936);
nand U17471 (N_17471,N_11673,N_13878);
xnor U17472 (N_17472,N_11255,N_14391);
and U17473 (N_17473,N_11018,N_11783);
xor U17474 (N_17474,N_10220,N_11646);
nor U17475 (N_17475,N_11155,N_14584);
nand U17476 (N_17476,N_14936,N_13009);
or U17477 (N_17477,N_11191,N_10314);
and U17478 (N_17478,N_11877,N_13050);
nor U17479 (N_17479,N_14553,N_12464);
nor U17480 (N_17480,N_11685,N_11580);
nand U17481 (N_17481,N_11375,N_11288);
nand U17482 (N_17482,N_10589,N_10941);
or U17483 (N_17483,N_11223,N_11199);
xor U17484 (N_17484,N_12063,N_14432);
nor U17485 (N_17485,N_10960,N_14704);
or U17486 (N_17486,N_13334,N_11586);
nand U17487 (N_17487,N_10797,N_13204);
xnor U17488 (N_17488,N_14221,N_14657);
nand U17489 (N_17489,N_12075,N_10262);
nand U17490 (N_17490,N_13401,N_14324);
nor U17491 (N_17491,N_11169,N_11514);
nor U17492 (N_17492,N_10274,N_13925);
nor U17493 (N_17493,N_10074,N_13897);
xor U17494 (N_17494,N_13093,N_13919);
nor U17495 (N_17495,N_10149,N_13238);
and U17496 (N_17496,N_12323,N_11949);
and U17497 (N_17497,N_10900,N_14608);
nor U17498 (N_17498,N_11585,N_12240);
nor U17499 (N_17499,N_13570,N_10044);
or U17500 (N_17500,N_14210,N_13433);
xor U17501 (N_17501,N_13537,N_10988);
nand U17502 (N_17502,N_11026,N_12828);
or U17503 (N_17503,N_12929,N_12893);
or U17504 (N_17504,N_13682,N_10860);
nand U17505 (N_17505,N_10789,N_13953);
nor U17506 (N_17506,N_10239,N_13893);
nor U17507 (N_17507,N_10894,N_12834);
nand U17508 (N_17508,N_12110,N_14643);
nand U17509 (N_17509,N_13678,N_10984);
and U17510 (N_17510,N_11264,N_13609);
nand U17511 (N_17511,N_12460,N_13984);
or U17512 (N_17512,N_11797,N_12139);
xnor U17513 (N_17513,N_11304,N_14667);
nor U17514 (N_17514,N_11696,N_13514);
nand U17515 (N_17515,N_11083,N_12176);
nand U17516 (N_17516,N_13847,N_13091);
xor U17517 (N_17517,N_10875,N_12950);
nand U17518 (N_17518,N_10055,N_14085);
or U17519 (N_17519,N_11754,N_12390);
nand U17520 (N_17520,N_12897,N_11279);
nand U17521 (N_17521,N_11453,N_12777);
and U17522 (N_17522,N_12243,N_14729);
nand U17523 (N_17523,N_12564,N_10415);
xor U17524 (N_17524,N_12027,N_10722);
and U17525 (N_17525,N_13287,N_12609);
or U17526 (N_17526,N_10472,N_10621);
nor U17527 (N_17527,N_13194,N_14931);
nand U17528 (N_17528,N_12267,N_10945);
or U17529 (N_17529,N_11042,N_11117);
nand U17530 (N_17530,N_13505,N_14994);
or U17531 (N_17531,N_13572,N_10049);
and U17532 (N_17532,N_12310,N_10702);
nor U17533 (N_17533,N_13236,N_10970);
xnor U17534 (N_17534,N_12920,N_10516);
and U17535 (N_17535,N_10752,N_12164);
nand U17536 (N_17536,N_13268,N_12538);
and U17537 (N_17537,N_12797,N_14003);
or U17538 (N_17538,N_12653,N_13373);
nor U17539 (N_17539,N_11602,N_10733);
and U17540 (N_17540,N_14756,N_12704);
nor U17541 (N_17541,N_14833,N_10855);
or U17542 (N_17542,N_13356,N_14774);
and U17543 (N_17543,N_12121,N_11943);
xnor U17544 (N_17544,N_13770,N_10874);
xor U17545 (N_17545,N_13353,N_12415);
xnor U17546 (N_17546,N_10391,N_10248);
nand U17547 (N_17547,N_14868,N_12909);
and U17548 (N_17548,N_13632,N_12187);
nand U17549 (N_17549,N_11541,N_13312);
and U17550 (N_17550,N_12214,N_13419);
and U17551 (N_17551,N_10315,N_10639);
or U17552 (N_17552,N_13113,N_13495);
nor U17553 (N_17553,N_11259,N_11627);
or U17554 (N_17554,N_14732,N_10829);
xor U17555 (N_17555,N_10167,N_11245);
or U17556 (N_17556,N_10916,N_12197);
and U17557 (N_17557,N_11130,N_13017);
or U17558 (N_17558,N_13244,N_12991);
or U17559 (N_17559,N_10855,N_13497);
nor U17560 (N_17560,N_10052,N_13240);
or U17561 (N_17561,N_10143,N_14431);
nand U17562 (N_17562,N_11792,N_12610);
xnor U17563 (N_17563,N_14135,N_10004);
nor U17564 (N_17564,N_10962,N_10476);
and U17565 (N_17565,N_11034,N_12520);
or U17566 (N_17566,N_14363,N_11549);
or U17567 (N_17567,N_10294,N_10320);
or U17568 (N_17568,N_11462,N_13563);
and U17569 (N_17569,N_12110,N_12767);
nor U17570 (N_17570,N_13954,N_11726);
nor U17571 (N_17571,N_11525,N_11083);
and U17572 (N_17572,N_12264,N_10790);
or U17573 (N_17573,N_12259,N_12013);
or U17574 (N_17574,N_13743,N_14959);
nand U17575 (N_17575,N_10220,N_10495);
nor U17576 (N_17576,N_11787,N_14410);
xor U17577 (N_17577,N_11402,N_11318);
or U17578 (N_17578,N_14229,N_10728);
nand U17579 (N_17579,N_11598,N_11847);
nand U17580 (N_17580,N_11103,N_13436);
xnor U17581 (N_17581,N_11066,N_10816);
nor U17582 (N_17582,N_10417,N_14706);
nand U17583 (N_17583,N_13303,N_14910);
or U17584 (N_17584,N_12613,N_13723);
and U17585 (N_17585,N_10412,N_10690);
and U17586 (N_17586,N_12489,N_13952);
xor U17587 (N_17587,N_13268,N_11753);
or U17588 (N_17588,N_10690,N_11605);
or U17589 (N_17589,N_13604,N_14201);
or U17590 (N_17590,N_11169,N_12095);
nand U17591 (N_17591,N_11625,N_11111);
and U17592 (N_17592,N_14871,N_10230);
or U17593 (N_17593,N_13542,N_12682);
nor U17594 (N_17594,N_12840,N_14113);
or U17595 (N_17595,N_12288,N_12114);
nor U17596 (N_17596,N_11996,N_12398);
xnor U17597 (N_17597,N_10042,N_11649);
or U17598 (N_17598,N_14630,N_12177);
nand U17599 (N_17599,N_13346,N_13927);
or U17600 (N_17600,N_12547,N_12534);
nor U17601 (N_17601,N_11080,N_13405);
xor U17602 (N_17602,N_14760,N_14287);
nand U17603 (N_17603,N_11984,N_12040);
or U17604 (N_17604,N_13690,N_14217);
nor U17605 (N_17605,N_11956,N_13902);
nor U17606 (N_17606,N_12641,N_10419);
nor U17607 (N_17607,N_14544,N_14584);
nand U17608 (N_17608,N_13167,N_13184);
nand U17609 (N_17609,N_11310,N_11806);
nor U17610 (N_17610,N_13439,N_14702);
and U17611 (N_17611,N_11941,N_13005);
nor U17612 (N_17612,N_12247,N_14987);
xor U17613 (N_17613,N_11989,N_14498);
nand U17614 (N_17614,N_11486,N_12623);
nand U17615 (N_17615,N_11486,N_13779);
nor U17616 (N_17616,N_12727,N_10430);
nor U17617 (N_17617,N_14897,N_14987);
nand U17618 (N_17618,N_14065,N_11397);
xor U17619 (N_17619,N_14780,N_10103);
nand U17620 (N_17620,N_12600,N_13634);
nand U17621 (N_17621,N_10457,N_11105);
nand U17622 (N_17622,N_11922,N_10697);
and U17623 (N_17623,N_14025,N_14342);
or U17624 (N_17624,N_14023,N_10549);
nor U17625 (N_17625,N_11224,N_12100);
and U17626 (N_17626,N_10915,N_10496);
nand U17627 (N_17627,N_11557,N_10985);
and U17628 (N_17628,N_14900,N_12938);
or U17629 (N_17629,N_13028,N_13777);
nand U17630 (N_17630,N_12784,N_12671);
nor U17631 (N_17631,N_14483,N_13111);
nor U17632 (N_17632,N_12682,N_10613);
xnor U17633 (N_17633,N_11208,N_10046);
nand U17634 (N_17634,N_14140,N_10920);
or U17635 (N_17635,N_13207,N_10462);
and U17636 (N_17636,N_11606,N_12055);
nor U17637 (N_17637,N_11555,N_10730);
nor U17638 (N_17638,N_11590,N_13576);
nand U17639 (N_17639,N_11184,N_12433);
xnor U17640 (N_17640,N_13087,N_11693);
or U17641 (N_17641,N_12075,N_10349);
nand U17642 (N_17642,N_10326,N_12830);
nor U17643 (N_17643,N_14435,N_10558);
nand U17644 (N_17644,N_11331,N_11967);
xor U17645 (N_17645,N_12535,N_13055);
or U17646 (N_17646,N_11427,N_14540);
or U17647 (N_17647,N_12516,N_12258);
xnor U17648 (N_17648,N_10057,N_10878);
or U17649 (N_17649,N_14566,N_11050);
xor U17650 (N_17650,N_13354,N_12844);
and U17651 (N_17651,N_10639,N_11261);
or U17652 (N_17652,N_13561,N_10704);
nor U17653 (N_17653,N_14964,N_10893);
nand U17654 (N_17654,N_11983,N_10009);
and U17655 (N_17655,N_14309,N_14370);
and U17656 (N_17656,N_11630,N_14100);
xnor U17657 (N_17657,N_12316,N_11798);
nor U17658 (N_17658,N_10428,N_10804);
or U17659 (N_17659,N_10035,N_14424);
xnor U17660 (N_17660,N_13920,N_13660);
nor U17661 (N_17661,N_10438,N_12524);
and U17662 (N_17662,N_12906,N_13496);
nand U17663 (N_17663,N_10014,N_14706);
or U17664 (N_17664,N_11880,N_13482);
and U17665 (N_17665,N_14350,N_14048);
nor U17666 (N_17666,N_10965,N_13276);
and U17667 (N_17667,N_10374,N_12909);
or U17668 (N_17668,N_13955,N_12725);
or U17669 (N_17669,N_11840,N_10325);
xor U17670 (N_17670,N_10093,N_13526);
nand U17671 (N_17671,N_13998,N_14492);
nand U17672 (N_17672,N_10648,N_13130);
nor U17673 (N_17673,N_11951,N_13755);
xnor U17674 (N_17674,N_14555,N_12494);
xnor U17675 (N_17675,N_13672,N_11262);
nor U17676 (N_17676,N_10127,N_12093);
nand U17677 (N_17677,N_12662,N_14206);
nor U17678 (N_17678,N_12683,N_11863);
xnor U17679 (N_17679,N_14483,N_13200);
and U17680 (N_17680,N_13743,N_13667);
nor U17681 (N_17681,N_10888,N_10808);
and U17682 (N_17682,N_13598,N_14103);
xnor U17683 (N_17683,N_10221,N_12422);
or U17684 (N_17684,N_11153,N_11926);
xor U17685 (N_17685,N_14432,N_12023);
nor U17686 (N_17686,N_10653,N_11933);
nand U17687 (N_17687,N_11831,N_14945);
and U17688 (N_17688,N_12834,N_11251);
and U17689 (N_17689,N_14231,N_10832);
nand U17690 (N_17690,N_12457,N_10671);
xor U17691 (N_17691,N_14640,N_10142);
and U17692 (N_17692,N_13734,N_10280);
nand U17693 (N_17693,N_13354,N_13612);
nand U17694 (N_17694,N_11211,N_13156);
nor U17695 (N_17695,N_13729,N_11092);
and U17696 (N_17696,N_13306,N_14568);
nand U17697 (N_17697,N_11427,N_12680);
nand U17698 (N_17698,N_14012,N_11272);
and U17699 (N_17699,N_10918,N_14113);
nor U17700 (N_17700,N_12270,N_13587);
nand U17701 (N_17701,N_10665,N_14280);
xor U17702 (N_17702,N_11621,N_12065);
nand U17703 (N_17703,N_14451,N_13471);
xor U17704 (N_17704,N_11054,N_14705);
nand U17705 (N_17705,N_14630,N_11135);
or U17706 (N_17706,N_12078,N_14775);
nand U17707 (N_17707,N_12170,N_14513);
nor U17708 (N_17708,N_13111,N_10867);
and U17709 (N_17709,N_10654,N_14388);
and U17710 (N_17710,N_13198,N_13232);
nor U17711 (N_17711,N_14476,N_14273);
or U17712 (N_17712,N_10261,N_14782);
and U17713 (N_17713,N_11211,N_11529);
or U17714 (N_17714,N_14324,N_13513);
or U17715 (N_17715,N_10193,N_11809);
nor U17716 (N_17716,N_10213,N_13595);
and U17717 (N_17717,N_13548,N_10698);
and U17718 (N_17718,N_12736,N_11174);
xor U17719 (N_17719,N_13460,N_10463);
nand U17720 (N_17720,N_14000,N_11740);
or U17721 (N_17721,N_12228,N_14758);
or U17722 (N_17722,N_11320,N_14932);
and U17723 (N_17723,N_14751,N_12813);
or U17724 (N_17724,N_14755,N_12947);
and U17725 (N_17725,N_13405,N_10642);
or U17726 (N_17726,N_11813,N_13026);
or U17727 (N_17727,N_11581,N_13911);
nand U17728 (N_17728,N_14934,N_13861);
or U17729 (N_17729,N_10821,N_10316);
or U17730 (N_17730,N_14639,N_10838);
nand U17731 (N_17731,N_10915,N_14426);
xor U17732 (N_17732,N_13230,N_10461);
nor U17733 (N_17733,N_13166,N_10091);
xor U17734 (N_17734,N_13006,N_11453);
nand U17735 (N_17735,N_14879,N_12545);
nor U17736 (N_17736,N_12580,N_13359);
xnor U17737 (N_17737,N_11796,N_10530);
xnor U17738 (N_17738,N_10210,N_13736);
nand U17739 (N_17739,N_11866,N_11799);
or U17740 (N_17740,N_14226,N_10377);
nand U17741 (N_17741,N_14705,N_14780);
or U17742 (N_17742,N_12574,N_14823);
xnor U17743 (N_17743,N_11186,N_13928);
or U17744 (N_17744,N_13721,N_10643);
xnor U17745 (N_17745,N_11831,N_12978);
xnor U17746 (N_17746,N_14502,N_14999);
nor U17747 (N_17747,N_10578,N_14697);
and U17748 (N_17748,N_13992,N_12433);
nand U17749 (N_17749,N_13710,N_10806);
nor U17750 (N_17750,N_10540,N_12888);
or U17751 (N_17751,N_12639,N_14570);
nor U17752 (N_17752,N_13498,N_11590);
nor U17753 (N_17753,N_13871,N_11674);
and U17754 (N_17754,N_14109,N_10864);
or U17755 (N_17755,N_10448,N_10579);
nor U17756 (N_17756,N_14296,N_14687);
nand U17757 (N_17757,N_10838,N_13821);
or U17758 (N_17758,N_10207,N_10680);
nand U17759 (N_17759,N_10511,N_13369);
and U17760 (N_17760,N_13977,N_11887);
nor U17761 (N_17761,N_10838,N_12473);
or U17762 (N_17762,N_11956,N_12848);
and U17763 (N_17763,N_12686,N_14539);
or U17764 (N_17764,N_14758,N_11972);
and U17765 (N_17765,N_13357,N_13232);
or U17766 (N_17766,N_13338,N_14829);
nor U17767 (N_17767,N_11743,N_14388);
and U17768 (N_17768,N_12023,N_13596);
or U17769 (N_17769,N_13642,N_13284);
xor U17770 (N_17770,N_10659,N_14158);
and U17771 (N_17771,N_14124,N_10049);
xnor U17772 (N_17772,N_12219,N_14798);
nor U17773 (N_17773,N_10116,N_14599);
and U17774 (N_17774,N_14390,N_11025);
nor U17775 (N_17775,N_12548,N_12309);
and U17776 (N_17776,N_11442,N_14921);
or U17777 (N_17777,N_13965,N_14143);
xor U17778 (N_17778,N_11660,N_12228);
nand U17779 (N_17779,N_11109,N_11488);
nand U17780 (N_17780,N_13219,N_10713);
xor U17781 (N_17781,N_13272,N_10467);
nand U17782 (N_17782,N_10386,N_12284);
nand U17783 (N_17783,N_10017,N_14355);
nor U17784 (N_17784,N_12032,N_12584);
nand U17785 (N_17785,N_10758,N_10780);
or U17786 (N_17786,N_13843,N_10249);
xor U17787 (N_17787,N_12999,N_10719);
nand U17788 (N_17788,N_14588,N_12463);
and U17789 (N_17789,N_12293,N_12742);
and U17790 (N_17790,N_10807,N_14443);
nor U17791 (N_17791,N_10022,N_11155);
nand U17792 (N_17792,N_11462,N_11574);
or U17793 (N_17793,N_11152,N_12024);
and U17794 (N_17794,N_11796,N_14969);
nor U17795 (N_17795,N_13897,N_13028);
or U17796 (N_17796,N_13691,N_13791);
nand U17797 (N_17797,N_10808,N_10366);
and U17798 (N_17798,N_13252,N_11596);
and U17799 (N_17799,N_13211,N_13646);
nand U17800 (N_17800,N_11034,N_12758);
nor U17801 (N_17801,N_14657,N_11350);
and U17802 (N_17802,N_14873,N_12121);
and U17803 (N_17803,N_13645,N_14913);
xor U17804 (N_17804,N_14082,N_13195);
and U17805 (N_17805,N_13631,N_11588);
nor U17806 (N_17806,N_14743,N_12872);
xor U17807 (N_17807,N_10370,N_10252);
xor U17808 (N_17808,N_11642,N_14643);
or U17809 (N_17809,N_14909,N_11665);
or U17810 (N_17810,N_11917,N_12513);
nor U17811 (N_17811,N_13642,N_12876);
xor U17812 (N_17812,N_11981,N_14102);
xor U17813 (N_17813,N_11306,N_12944);
or U17814 (N_17814,N_12605,N_11501);
xnor U17815 (N_17815,N_13655,N_10697);
or U17816 (N_17816,N_13428,N_13255);
or U17817 (N_17817,N_14630,N_10661);
xor U17818 (N_17818,N_13220,N_13384);
and U17819 (N_17819,N_13883,N_14284);
xnor U17820 (N_17820,N_10104,N_11932);
xnor U17821 (N_17821,N_14913,N_13815);
nand U17822 (N_17822,N_11390,N_13725);
xor U17823 (N_17823,N_12739,N_12857);
nand U17824 (N_17824,N_10659,N_13046);
nand U17825 (N_17825,N_10944,N_13810);
nor U17826 (N_17826,N_13290,N_12959);
or U17827 (N_17827,N_12576,N_12882);
nor U17828 (N_17828,N_12822,N_11971);
or U17829 (N_17829,N_13546,N_14425);
nor U17830 (N_17830,N_10044,N_13522);
nand U17831 (N_17831,N_14966,N_11302);
nand U17832 (N_17832,N_12979,N_11908);
nand U17833 (N_17833,N_11548,N_11044);
nand U17834 (N_17834,N_10280,N_12674);
and U17835 (N_17835,N_10747,N_14914);
nor U17836 (N_17836,N_13190,N_14474);
and U17837 (N_17837,N_14361,N_13254);
and U17838 (N_17838,N_14278,N_11996);
and U17839 (N_17839,N_11086,N_14161);
or U17840 (N_17840,N_12746,N_11839);
and U17841 (N_17841,N_11599,N_14045);
nor U17842 (N_17842,N_12606,N_12086);
nand U17843 (N_17843,N_12009,N_12950);
or U17844 (N_17844,N_12663,N_11295);
and U17845 (N_17845,N_10782,N_10434);
and U17846 (N_17846,N_10284,N_14413);
xnor U17847 (N_17847,N_12077,N_11771);
nand U17848 (N_17848,N_12903,N_10643);
or U17849 (N_17849,N_12858,N_13590);
nand U17850 (N_17850,N_11533,N_11866);
nor U17851 (N_17851,N_14269,N_12350);
and U17852 (N_17852,N_12980,N_10671);
nand U17853 (N_17853,N_13915,N_12845);
nor U17854 (N_17854,N_14887,N_10680);
xor U17855 (N_17855,N_11208,N_10405);
and U17856 (N_17856,N_12539,N_10102);
or U17857 (N_17857,N_13284,N_13241);
and U17858 (N_17858,N_13394,N_13715);
or U17859 (N_17859,N_10880,N_10399);
and U17860 (N_17860,N_12213,N_11118);
xor U17861 (N_17861,N_13101,N_14628);
nand U17862 (N_17862,N_14725,N_11711);
or U17863 (N_17863,N_10734,N_12522);
nor U17864 (N_17864,N_13157,N_13104);
and U17865 (N_17865,N_14951,N_12770);
and U17866 (N_17866,N_14285,N_12369);
nand U17867 (N_17867,N_14450,N_11402);
nor U17868 (N_17868,N_11982,N_13450);
xor U17869 (N_17869,N_11821,N_11090);
xnor U17870 (N_17870,N_11446,N_10129);
and U17871 (N_17871,N_13233,N_10949);
nand U17872 (N_17872,N_13477,N_10487);
and U17873 (N_17873,N_14172,N_11861);
and U17874 (N_17874,N_14095,N_11218);
and U17875 (N_17875,N_10029,N_13024);
nor U17876 (N_17876,N_12223,N_13425);
and U17877 (N_17877,N_11186,N_13810);
nand U17878 (N_17878,N_12219,N_11521);
nand U17879 (N_17879,N_13002,N_14441);
xnor U17880 (N_17880,N_11905,N_12807);
nand U17881 (N_17881,N_14426,N_12894);
nor U17882 (N_17882,N_12311,N_14819);
nor U17883 (N_17883,N_12900,N_11203);
or U17884 (N_17884,N_11231,N_14152);
or U17885 (N_17885,N_14418,N_10377);
xor U17886 (N_17886,N_10011,N_13350);
nor U17887 (N_17887,N_14506,N_12706);
and U17888 (N_17888,N_12040,N_14332);
or U17889 (N_17889,N_14919,N_14376);
or U17890 (N_17890,N_13935,N_14447);
or U17891 (N_17891,N_11052,N_10610);
and U17892 (N_17892,N_11737,N_14317);
nand U17893 (N_17893,N_13399,N_11667);
and U17894 (N_17894,N_12051,N_10530);
or U17895 (N_17895,N_13161,N_12716);
or U17896 (N_17896,N_11350,N_14433);
nand U17897 (N_17897,N_10044,N_13477);
xnor U17898 (N_17898,N_14777,N_10573);
nand U17899 (N_17899,N_11848,N_10743);
nand U17900 (N_17900,N_14183,N_10495);
nand U17901 (N_17901,N_14671,N_10039);
and U17902 (N_17902,N_11189,N_14477);
nor U17903 (N_17903,N_14414,N_10486);
xnor U17904 (N_17904,N_11677,N_10857);
or U17905 (N_17905,N_11083,N_10702);
nor U17906 (N_17906,N_13440,N_14359);
xnor U17907 (N_17907,N_11104,N_10658);
or U17908 (N_17908,N_13380,N_11488);
and U17909 (N_17909,N_11367,N_12882);
nand U17910 (N_17910,N_10260,N_12210);
nand U17911 (N_17911,N_13063,N_14815);
nand U17912 (N_17912,N_10330,N_14481);
nand U17913 (N_17913,N_11649,N_14947);
nor U17914 (N_17914,N_14387,N_13410);
or U17915 (N_17915,N_11423,N_10292);
nor U17916 (N_17916,N_10099,N_12734);
nor U17917 (N_17917,N_10617,N_10826);
nor U17918 (N_17918,N_11386,N_11047);
or U17919 (N_17919,N_14773,N_13190);
nand U17920 (N_17920,N_13774,N_14283);
nand U17921 (N_17921,N_13455,N_11808);
nor U17922 (N_17922,N_10684,N_12854);
nor U17923 (N_17923,N_10517,N_11278);
xor U17924 (N_17924,N_10599,N_14217);
nor U17925 (N_17925,N_13420,N_14762);
or U17926 (N_17926,N_12765,N_13289);
nand U17927 (N_17927,N_12667,N_12396);
nand U17928 (N_17928,N_13008,N_11230);
or U17929 (N_17929,N_13317,N_14680);
xor U17930 (N_17930,N_10530,N_14568);
and U17931 (N_17931,N_10756,N_14906);
and U17932 (N_17932,N_13753,N_13420);
and U17933 (N_17933,N_10691,N_10433);
and U17934 (N_17934,N_12655,N_10296);
xor U17935 (N_17935,N_10166,N_10836);
and U17936 (N_17936,N_13842,N_12895);
or U17937 (N_17937,N_11748,N_12686);
nand U17938 (N_17938,N_13165,N_10863);
xnor U17939 (N_17939,N_11232,N_13787);
nor U17940 (N_17940,N_14790,N_13779);
or U17941 (N_17941,N_12242,N_12275);
xor U17942 (N_17942,N_11740,N_12014);
xor U17943 (N_17943,N_13461,N_14598);
nand U17944 (N_17944,N_14499,N_12536);
and U17945 (N_17945,N_10529,N_14550);
or U17946 (N_17946,N_13669,N_14049);
nor U17947 (N_17947,N_11420,N_10898);
or U17948 (N_17948,N_14679,N_13209);
nor U17949 (N_17949,N_13743,N_14906);
nor U17950 (N_17950,N_11742,N_10826);
and U17951 (N_17951,N_10845,N_12494);
or U17952 (N_17952,N_14683,N_12116);
nand U17953 (N_17953,N_14028,N_12696);
and U17954 (N_17954,N_14504,N_13896);
nor U17955 (N_17955,N_12394,N_14858);
or U17956 (N_17956,N_11839,N_14098);
nand U17957 (N_17957,N_14838,N_12374);
xor U17958 (N_17958,N_11890,N_14651);
and U17959 (N_17959,N_11690,N_14410);
nor U17960 (N_17960,N_13380,N_11485);
and U17961 (N_17961,N_11920,N_14513);
or U17962 (N_17962,N_11348,N_12867);
xnor U17963 (N_17963,N_13859,N_14845);
and U17964 (N_17964,N_13660,N_12574);
and U17965 (N_17965,N_14287,N_11082);
nand U17966 (N_17966,N_11926,N_13671);
and U17967 (N_17967,N_11793,N_11373);
xnor U17968 (N_17968,N_12213,N_12251);
xor U17969 (N_17969,N_11561,N_10085);
nor U17970 (N_17970,N_12661,N_14853);
and U17971 (N_17971,N_13356,N_11226);
nor U17972 (N_17972,N_14239,N_13934);
nor U17973 (N_17973,N_13747,N_11111);
nand U17974 (N_17974,N_11325,N_13295);
or U17975 (N_17975,N_11230,N_13816);
nand U17976 (N_17976,N_11248,N_12022);
nand U17977 (N_17977,N_13836,N_14634);
nor U17978 (N_17978,N_12153,N_14218);
xnor U17979 (N_17979,N_13966,N_14745);
and U17980 (N_17980,N_14743,N_11603);
and U17981 (N_17981,N_14892,N_12256);
xnor U17982 (N_17982,N_11641,N_11339);
nor U17983 (N_17983,N_10307,N_14836);
xor U17984 (N_17984,N_11301,N_11752);
nand U17985 (N_17985,N_11097,N_12456);
or U17986 (N_17986,N_11736,N_10970);
or U17987 (N_17987,N_10362,N_11176);
nand U17988 (N_17988,N_14434,N_13856);
and U17989 (N_17989,N_14143,N_14816);
and U17990 (N_17990,N_11888,N_14354);
and U17991 (N_17991,N_11653,N_12641);
xnor U17992 (N_17992,N_12305,N_12532);
or U17993 (N_17993,N_12301,N_12346);
nor U17994 (N_17994,N_10502,N_13428);
xor U17995 (N_17995,N_14664,N_10848);
or U17996 (N_17996,N_10019,N_12938);
and U17997 (N_17997,N_12977,N_11244);
xnor U17998 (N_17998,N_12827,N_13428);
and U17999 (N_17999,N_12467,N_12120);
nand U18000 (N_18000,N_10709,N_10641);
and U18001 (N_18001,N_12868,N_10488);
or U18002 (N_18002,N_11770,N_13757);
nor U18003 (N_18003,N_12690,N_14677);
xnor U18004 (N_18004,N_12592,N_13950);
nand U18005 (N_18005,N_14766,N_13652);
or U18006 (N_18006,N_12010,N_13307);
or U18007 (N_18007,N_14621,N_12162);
or U18008 (N_18008,N_14852,N_12550);
or U18009 (N_18009,N_12341,N_10363);
nor U18010 (N_18010,N_11338,N_12114);
xnor U18011 (N_18011,N_10091,N_13198);
and U18012 (N_18012,N_14670,N_14008);
nor U18013 (N_18013,N_11400,N_12778);
nand U18014 (N_18014,N_10461,N_12600);
nand U18015 (N_18015,N_11157,N_11899);
xnor U18016 (N_18016,N_10159,N_12250);
xor U18017 (N_18017,N_13920,N_12238);
nand U18018 (N_18018,N_12111,N_12295);
xnor U18019 (N_18019,N_11540,N_12978);
or U18020 (N_18020,N_10263,N_13905);
nand U18021 (N_18021,N_12222,N_13436);
or U18022 (N_18022,N_14145,N_13933);
nor U18023 (N_18023,N_13764,N_13682);
or U18024 (N_18024,N_10369,N_12010);
and U18025 (N_18025,N_12675,N_14885);
xnor U18026 (N_18026,N_11323,N_13016);
and U18027 (N_18027,N_14830,N_14172);
or U18028 (N_18028,N_11690,N_10511);
and U18029 (N_18029,N_12562,N_10396);
and U18030 (N_18030,N_10058,N_12368);
nor U18031 (N_18031,N_13220,N_10878);
and U18032 (N_18032,N_13141,N_10488);
nor U18033 (N_18033,N_13804,N_11768);
nand U18034 (N_18034,N_12247,N_11686);
xnor U18035 (N_18035,N_10967,N_12146);
xor U18036 (N_18036,N_14960,N_12459);
nor U18037 (N_18037,N_11978,N_12150);
nor U18038 (N_18038,N_13689,N_11851);
nand U18039 (N_18039,N_12735,N_14851);
or U18040 (N_18040,N_11808,N_14571);
xnor U18041 (N_18041,N_10199,N_12857);
nor U18042 (N_18042,N_10227,N_10242);
and U18043 (N_18043,N_12505,N_13377);
or U18044 (N_18044,N_12093,N_10810);
and U18045 (N_18045,N_10192,N_12608);
nand U18046 (N_18046,N_11076,N_11366);
xor U18047 (N_18047,N_14979,N_11187);
and U18048 (N_18048,N_11465,N_10862);
or U18049 (N_18049,N_10253,N_12976);
xnor U18050 (N_18050,N_12056,N_13200);
nor U18051 (N_18051,N_14737,N_13298);
or U18052 (N_18052,N_12724,N_11085);
or U18053 (N_18053,N_10863,N_11648);
nand U18054 (N_18054,N_10927,N_12630);
xnor U18055 (N_18055,N_13774,N_14358);
and U18056 (N_18056,N_10046,N_14859);
and U18057 (N_18057,N_10253,N_11496);
and U18058 (N_18058,N_13318,N_14146);
and U18059 (N_18059,N_14136,N_12399);
or U18060 (N_18060,N_14895,N_14152);
nand U18061 (N_18061,N_12873,N_14569);
and U18062 (N_18062,N_10762,N_11428);
nand U18063 (N_18063,N_10513,N_13338);
or U18064 (N_18064,N_12690,N_12596);
nand U18065 (N_18065,N_12376,N_14697);
xor U18066 (N_18066,N_13248,N_11728);
and U18067 (N_18067,N_11976,N_14509);
or U18068 (N_18068,N_10151,N_12158);
and U18069 (N_18069,N_13829,N_10907);
nor U18070 (N_18070,N_11716,N_13086);
nand U18071 (N_18071,N_14770,N_12650);
nand U18072 (N_18072,N_13277,N_11389);
xor U18073 (N_18073,N_12246,N_14208);
xor U18074 (N_18074,N_10411,N_10594);
and U18075 (N_18075,N_13445,N_13645);
nor U18076 (N_18076,N_10786,N_11294);
or U18077 (N_18077,N_13568,N_12281);
and U18078 (N_18078,N_12913,N_13989);
nand U18079 (N_18079,N_11855,N_12633);
xnor U18080 (N_18080,N_13911,N_13148);
xor U18081 (N_18081,N_13030,N_14199);
nor U18082 (N_18082,N_14647,N_11210);
or U18083 (N_18083,N_13562,N_10127);
nand U18084 (N_18084,N_11746,N_13597);
or U18085 (N_18085,N_11272,N_11924);
nor U18086 (N_18086,N_14208,N_13260);
nand U18087 (N_18087,N_11112,N_11982);
and U18088 (N_18088,N_11692,N_12175);
xnor U18089 (N_18089,N_10057,N_11938);
nor U18090 (N_18090,N_11317,N_12519);
nand U18091 (N_18091,N_13188,N_11379);
or U18092 (N_18092,N_10430,N_10249);
nand U18093 (N_18093,N_14678,N_10460);
xor U18094 (N_18094,N_13506,N_12272);
or U18095 (N_18095,N_10037,N_11009);
or U18096 (N_18096,N_13863,N_10697);
xor U18097 (N_18097,N_14695,N_13252);
nor U18098 (N_18098,N_10337,N_12136);
nor U18099 (N_18099,N_14976,N_12256);
or U18100 (N_18100,N_12011,N_12190);
or U18101 (N_18101,N_11653,N_10414);
nand U18102 (N_18102,N_14317,N_11003);
xnor U18103 (N_18103,N_11766,N_12273);
or U18104 (N_18104,N_14034,N_10348);
xor U18105 (N_18105,N_14848,N_13237);
and U18106 (N_18106,N_13187,N_11431);
or U18107 (N_18107,N_11678,N_10254);
nand U18108 (N_18108,N_14959,N_13783);
and U18109 (N_18109,N_10920,N_10552);
nor U18110 (N_18110,N_13362,N_12625);
and U18111 (N_18111,N_12715,N_11635);
nor U18112 (N_18112,N_11502,N_12328);
nand U18113 (N_18113,N_14122,N_14698);
nor U18114 (N_18114,N_10371,N_12374);
nor U18115 (N_18115,N_10003,N_14162);
xor U18116 (N_18116,N_13901,N_14698);
nor U18117 (N_18117,N_13489,N_13070);
or U18118 (N_18118,N_14217,N_11279);
or U18119 (N_18119,N_12242,N_14220);
and U18120 (N_18120,N_14742,N_12819);
nand U18121 (N_18121,N_10807,N_14871);
xnor U18122 (N_18122,N_11573,N_12526);
nor U18123 (N_18123,N_10930,N_13869);
or U18124 (N_18124,N_14437,N_12535);
and U18125 (N_18125,N_11711,N_14736);
and U18126 (N_18126,N_11975,N_10425);
or U18127 (N_18127,N_12222,N_12624);
or U18128 (N_18128,N_11863,N_11565);
and U18129 (N_18129,N_11676,N_14601);
and U18130 (N_18130,N_13889,N_13143);
or U18131 (N_18131,N_13516,N_12464);
or U18132 (N_18132,N_11770,N_14678);
nor U18133 (N_18133,N_10664,N_14558);
nand U18134 (N_18134,N_10324,N_12947);
and U18135 (N_18135,N_14401,N_14586);
or U18136 (N_18136,N_10978,N_13277);
nor U18137 (N_18137,N_12152,N_13448);
or U18138 (N_18138,N_10751,N_13191);
nor U18139 (N_18139,N_14365,N_13079);
nand U18140 (N_18140,N_12155,N_12965);
xnor U18141 (N_18141,N_11073,N_13409);
nand U18142 (N_18142,N_14304,N_14679);
nor U18143 (N_18143,N_13468,N_14595);
and U18144 (N_18144,N_13121,N_13925);
nand U18145 (N_18145,N_11029,N_14525);
nand U18146 (N_18146,N_10256,N_12984);
and U18147 (N_18147,N_13817,N_14428);
nand U18148 (N_18148,N_10231,N_14659);
and U18149 (N_18149,N_14092,N_13417);
nand U18150 (N_18150,N_11762,N_12540);
and U18151 (N_18151,N_14867,N_13327);
and U18152 (N_18152,N_12314,N_11707);
xor U18153 (N_18153,N_11884,N_14571);
or U18154 (N_18154,N_12837,N_11851);
and U18155 (N_18155,N_14682,N_12158);
and U18156 (N_18156,N_11966,N_13844);
nand U18157 (N_18157,N_14070,N_14255);
and U18158 (N_18158,N_14322,N_11588);
nor U18159 (N_18159,N_10573,N_14213);
or U18160 (N_18160,N_10964,N_13998);
and U18161 (N_18161,N_12852,N_14693);
or U18162 (N_18162,N_10446,N_13140);
nor U18163 (N_18163,N_12568,N_14333);
xor U18164 (N_18164,N_12651,N_12518);
and U18165 (N_18165,N_14157,N_10123);
xor U18166 (N_18166,N_12224,N_11128);
or U18167 (N_18167,N_10200,N_10220);
and U18168 (N_18168,N_13755,N_10170);
nand U18169 (N_18169,N_12913,N_12321);
and U18170 (N_18170,N_10434,N_14887);
xnor U18171 (N_18171,N_11556,N_10739);
nand U18172 (N_18172,N_10961,N_14145);
nand U18173 (N_18173,N_14534,N_10233);
nor U18174 (N_18174,N_10293,N_14180);
or U18175 (N_18175,N_13348,N_11555);
or U18176 (N_18176,N_10341,N_14623);
nor U18177 (N_18177,N_14216,N_13047);
and U18178 (N_18178,N_13230,N_14728);
xor U18179 (N_18179,N_11756,N_11628);
nor U18180 (N_18180,N_11041,N_14442);
nor U18181 (N_18181,N_13883,N_13588);
nor U18182 (N_18182,N_10102,N_12163);
nor U18183 (N_18183,N_10375,N_12485);
or U18184 (N_18184,N_11354,N_14599);
xor U18185 (N_18185,N_12445,N_12241);
or U18186 (N_18186,N_10655,N_11252);
and U18187 (N_18187,N_12529,N_12415);
or U18188 (N_18188,N_10747,N_13398);
and U18189 (N_18189,N_11779,N_14731);
and U18190 (N_18190,N_12650,N_11329);
nor U18191 (N_18191,N_11301,N_14081);
or U18192 (N_18192,N_13120,N_10161);
nor U18193 (N_18193,N_13448,N_10182);
or U18194 (N_18194,N_14274,N_11102);
or U18195 (N_18195,N_11085,N_10822);
and U18196 (N_18196,N_13184,N_14550);
and U18197 (N_18197,N_10827,N_10323);
and U18198 (N_18198,N_14582,N_14437);
nor U18199 (N_18199,N_11725,N_11319);
or U18200 (N_18200,N_13761,N_11691);
xor U18201 (N_18201,N_10546,N_13024);
or U18202 (N_18202,N_11255,N_12039);
xor U18203 (N_18203,N_13493,N_13298);
nor U18204 (N_18204,N_14818,N_14354);
and U18205 (N_18205,N_10516,N_10205);
xor U18206 (N_18206,N_11487,N_12949);
or U18207 (N_18207,N_13223,N_11616);
or U18208 (N_18208,N_13774,N_10079);
nor U18209 (N_18209,N_10200,N_14741);
nor U18210 (N_18210,N_10733,N_11536);
xnor U18211 (N_18211,N_13898,N_12505);
nand U18212 (N_18212,N_11206,N_13207);
nor U18213 (N_18213,N_13458,N_12740);
or U18214 (N_18214,N_14045,N_11896);
nor U18215 (N_18215,N_12324,N_12505);
and U18216 (N_18216,N_10244,N_13241);
or U18217 (N_18217,N_11123,N_10820);
and U18218 (N_18218,N_12934,N_10081);
xor U18219 (N_18219,N_14004,N_12933);
nand U18220 (N_18220,N_14560,N_14075);
nor U18221 (N_18221,N_11060,N_10414);
nand U18222 (N_18222,N_13831,N_11725);
nor U18223 (N_18223,N_12314,N_10121);
nor U18224 (N_18224,N_10843,N_11083);
and U18225 (N_18225,N_10137,N_12605);
and U18226 (N_18226,N_11680,N_11981);
or U18227 (N_18227,N_14737,N_12380);
nor U18228 (N_18228,N_11813,N_14227);
nor U18229 (N_18229,N_13174,N_12590);
xor U18230 (N_18230,N_12408,N_14926);
nor U18231 (N_18231,N_13839,N_10316);
or U18232 (N_18232,N_14469,N_12982);
nor U18233 (N_18233,N_12743,N_12745);
nand U18234 (N_18234,N_13389,N_10165);
and U18235 (N_18235,N_11773,N_11873);
and U18236 (N_18236,N_10197,N_13933);
xor U18237 (N_18237,N_12901,N_13081);
xnor U18238 (N_18238,N_12940,N_13896);
or U18239 (N_18239,N_12970,N_12190);
nand U18240 (N_18240,N_12725,N_14173);
xnor U18241 (N_18241,N_10671,N_12267);
nand U18242 (N_18242,N_13419,N_13361);
nand U18243 (N_18243,N_11027,N_10534);
xor U18244 (N_18244,N_12405,N_11665);
and U18245 (N_18245,N_11285,N_14723);
xor U18246 (N_18246,N_14585,N_14109);
or U18247 (N_18247,N_10257,N_13079);
xnor U18248 (N_18248,N_12433,N_11930);
and U18249 (N_18249,N_12851,N_10878);
nor U18250 (N_18250,N_12919,N_12737);
and U18251 (N_18251,N_13404,N_10303);
xor U18252 (N_18252,N_13758,N_14125);
and U18253 (N_18253,N_12790,N_12523);
xor U18254 (N_18254,N_13065,N_13572);
nor U18255 (N_18255,N_14205,N_12568);
nor U18256 (N_18256,N_13717,N_12407);
and U18257 (N_18257,N_13012,N_13859);
nand U18258 (N_18258,N_11784,N_10653);
nand U18259 (N_18259,N_12091,N_13686);
xor U18260 (N_18260,N_12537,N_11222);
and U18261 (N_18261,N_14348,N_12709);
and U18262 (N_18262,N_11591,N_11507);
nor U18263 (N_18263,N_10254,N_14442);
nor U18264 (N_18264,N_10464,N_11058);
or U18265 (N_18265,N_11111,N_10199);
and U18266 (N_18266,N_13411,N_14616);
or U18267 (N_18267,N_13282,N_12101);
nor U18268 (N_18268,N_14418,N_10787);
and U18269 (N_18269,N_12236,N_12889);
xor U18270 (N_18270,N_14059,N_12660);
xnor U18271 (N_18271,N_11707,N_13998);
xnor U18272 (N_18272,N_14190,N_11003);
nor U18273 (N_18273,N_11203,N_11265);
or U18274 (N_18274,N_14722,N_13584);
nor U18275 (N_18275,N_10904,N_10493);
and U18276 (N_18276,N_12012,N_13978);
nor U18277 (N_18277,N_14325,N_10418);
and U18278 (N_18278,N_13639,N_12826);
nand U18279 (N_18279,N_12173,N_12541);
or U18280 (N_18280,N_12024,N_14959);
or U18281 (N_18281,N_10070,N_12672);
xor U18282 (N_18282,N_14907,N_12596);
xor U18283 (N_18283,N_12025,N_13727);
xor U18284 (N_18284,N_10286,N_10126);
nor U18285 (N_18285,N_10634,N_14607);
nand U18286 (N_18286,N_10591,N_10993);
nor U18287 (N_18287,N_11274,N_10549);
xnor U18288 (N_18288,N_13473,N_10228);
and U18289 (N_18289,N_11515,N_14882);
nand U18290 (N_18290,N_11697,N_13687);
nor U18291 (N_18291,N_12108,N_12988);
xor U18292 (N_18292,N_11499,N_11899);
or U18293 (N_18293,N_10474,N_11453);
and U18294 (N_18294,N_13488,N_11380);
or U18295 (N_18295,N_14668,N_14525);
nor U18296 (N_18296,N_10884,N_11045);
nand U18297 (N_18297,N_11948,N_14312);
nand U18298 (N_18298,N_14620,N_13167);
nand U18299 (N_18299,N_14135,N_12541);
nand U18300 (N_18300,N_13624,N_13248);
xnor U18301 (N_18301,N_14325,N_14706);
and U18302 (N_18302,N_10097,N_10137);
nor U18303 (N_18303,N_12077,N_14995);
nand U18304 (N_18304,N_11362,N_13542);
xnor U18305 (N_18305,N_12045,N_10181);
nand U18306 (N_18306,N_10865,N_11294);
xor U18307 (N_18307,N_12834,N_11995);
xnor U18308 (N_18308,N_14608,N_11876);
and U18309 (N_18309,N_12534,N_13097);
and U18310 (N_18310,N_11575,N_11033);
and U18311 (N_18311,N_14999,N_13639);
nand U18312 (N_18312,N_14443,N_13557);
or U18313 (N_18313,N_11055,N_10906);
nand U18314 (N_18314,N_12425,N_10085);
or U18315 (N_18315,N_12877,N_11970);
and U18316 (N_18316,N_11275,N_14334);
or U18317 (N_18317,N_11315,N_14075);
nand U18318 (N_18318,N_14801,N_10004);
and U18319 (N_18319,N_14628,N_12646);
nor U18320 (N_18320,N_10107,N_14379);
nor U18321 (N_18321,N_13647,N_12195);
or U18322 (N_18322,N_11495,N_11625);
nor U18323 (N_18323,N_11829,N_11878);
and U18324 (N_18324,N_12360,N_13403);
nand U18325 (N_18325,N_14065,N_13238);
nor U18326 (N_18326,N_10923,N_12795);
nor U18327 (N_18327,N_11965,N_11873);
nand U18328 (N_18328,N_12873,N_11918);
or U18329 (N_18329,N_11611,N_13124);
nor U18330 (N_18330,N_10146,N_13347);
and U18331 (N_18331,N_13444,N_10191);
nand U18332 (N_18332,N_11323,N_11769);
or U18333 (N_18333,N_13126,N_14332);
and U18334 (N_18334,N_12886,N_10992);
xor U18335 (N_18335,N_13712,N_14857);
and U18336 (N_18336,N_12521,N_10764);
nor U18337 (N_18337,N_10302,N_12231);
nor U18338 (N_18338,N_10494,N_13591);
xor U18339 (N_18339,N_13309,N_12780);
xnor U18340 (N_18340,N_14422,N_13695);
and U18341 (N_18341,N_11257,N_11038);
nand U18342 (N_18342,N_13451,N_13982);
nor U18343 (N_18343,N_10157,N_11886);
xnor U18344 (N_18344,N_11489,N_12666);
nor U18345 (N_18345,N_11646,N_10512);
and U18346 (N_18346,N_10083,N_10111);
and U18347 (N_18347,N_10358,N_13426);
xnor U18348 (N_18348,N_11647,N_11835);
and U18349 (N_18349,N_13681,N_12625);
xnor U18350 (N_18350,N_14219,N_11958);
nand U18351 (N_18351,N_13053,N_12821);
xor U18352 (N_18352,N_14248,N_11562);
and U18353 (N_18353,N_12975,N_14043);
xnor U18354 (N_18354,N_10959,N_11592);
nand U18355 (N_18355,N_11340,N_12376);
nor U18356 (N_18356,N_12754,N_13326);
nor U18357 (N_18357,N_13417,N_10664);
or U18358 (N_18358,N_12938,N_10274);
nor U18359 (N_18359,N_14510,N_13420);
and U18360 (N_18360,N_14482,N_12883);
nor U18361 (N_18361,N_13348,N_13057);
xnor U18362 (N_18362,N_12455,N_12018);
and U18363 (N_18363,N_11777,N_11121);
and U18364 (N_18364,N_11874,N_12584);
or U18365 (N_18365,N_12494,N_12119);
xor U18366 (N_18366,N_12278,N_12346);
xnor U18367 (N_18367,N_12606,N_10827);
and U18368 (N_18368,N_14393,N_14661);
or U18369 (N_18369,N_14610,N_10223);
xor U18370 (N_18370,N_12773,N_14655);
nor U18371 (N_18371,N_14576,N_11645);
nand U18372 (N_18372,N_10300,N_10285);
or U18373 (N_18373,N_14159,N_10714);
nand U18374 (N_18374,N_14682,N_12583);
or U18375 (N_18375,N_14139,N_11150);
nand U18376 (N_18376,N_14418,N_12438);
xnor U18377 (N_18377,N_12783,N_14287);
nor U18378 (N_18378,N_11636,N_10619);
xor U18379 (N_18379,N_13478,N_14878);
or U18380 (N_18380,N_13893,N_11972);
nor U18381 (N_18381,N_13694,N_12474);
or U18382 (N_18382,N_14941,N_11971);
nand U18383 (N_18383,N_14862,N_14283);
nor U18384 (N_18384,N_12942,N_10388);
or U18385 (N_18385,N_10723,N_12592);
and U18386 (N_18386,N_12031,N_11974);
xnor U18387 (N_18387,N_11073,N_14682);
xor U18388 (N_18388,N_14227,N_12315);
nand U18389 (N_18389,N_14543,N_14310);
and U18390 (N_18390,N_12789,N_12234);
or U18391 (N_18391,N_14287,N_13424);
and U18392 (N_18392,N_13285,N_14411);
nor U18393 (N_18393,N_13193,N_13743);
or U18394 (N_18394,N_14763,N_14342);
and U18395 (N_18395,N_11358,N_12892);
nand U18396 (N_18396,N_12735,N_12742);
nand U18397 (N_18397,N_10451,N_10547);
nor U18398 (N_18398,N_10125,N_14722);
nor U18399 (N_18399,N_13940,N_10228);
and U18400 (N_18400,N_12584,N_10561);
nor U18401 (N_18401,N_10613,N_11029);
and U18402 (N_18402,N_12629,N_12003);
nand U18403 (N_18403,N_12837,N_13612);
nor U18404 (N_18404,N_14789,N_13003);
and U18405 (N_18405,N_12938,N_14517);
xor U18406 (N_18406,N_11849,N_14898);
and U18407 (N_18407,N_13453,N_12744);
xnor U18408 (N_18408,N_10477,N_12790);
xor U18409 (N_18409,N_11699,N_13418);
and U18410 (N_18410,N_12160,N_13020);
xnor U18411 (N_18411,N_10120,N_11893);
nand U18412 (N_18412,N_13613,N_12840);
or U18413 (N_18413,N_14179,N_10861);
nor U18414 (N_18414,N_14419,N_12072);
and U18415 (N_18415,N_11452,N_14168);
and U18416 (N_18416,N_11303,N_10889);
nand U18417 (N_18417,N_14989,N_14200);
xor U18418 (N_18418,N_10772,N_13011);
or U18419 (N_18419,N_12126,N_12480);
and U18420 (N_18420,N_13385,N_14157);
and U18421 (N_18421,N_12825,N_11774);
and U18422 (N_18422,N_11618,N_12846);
xnor U18423 (N_18423,N_13465,N_10248);
nand U18424 (N_18424,N_13449,N_10085);
and U18425 (N_18425,N_11379,N_12300);
or U18426 (N_18426,N_11308,N_13369);
xor U18427 (N_18427,N_13207,N_10148);
xnor U18428 (N_18428,N_13458,N_11790);
nor U18429 (N_18429,N_10309,N_10876);
nor U18430 (N_18430,N_12642,N_11991);
and U18431 (N_18431,N_12794,N_12148);
nor U18432 (N_18432,N_14672,N_12845);
or U18433 (N_18433,N_13485,N_12002);
nor U18434 (N_18434,N_12615,N_14701);
nand U18435 (N_18435,N_14385,N_10652);
and U18436 (N_18436,N_12967,N_10626);
nor U18437 (N_18437,N_14044,N_14973);
and U18438 (N_18438,N_14438,N_14198);
or U18439 (N_18439,N_11378,N_11317);
or U18440 (N_18440,N_14902,N_10218);
and U18441 (N_18441,N_13344,N_11122);
nor U18442 (N_18442,N_14955,N_12871);
nor U18443 (N_18443,N_11443,N_10256);
xor U18444 (N_18444,N_13415,N_10332);
nand U18445 (N_18445,N_13643,N_11518);
or U18446 (N_18446,N_12273,N_11702);
nor U18447 (N_18447,N_10051,N_14869);
and U18448 (N_18448,N_13823,N_11657);
and U18449 (N_18449,N_14043,N_12049);
and U18450 (N_18450,N_10223,N_11953);
nand U18451 (N_18451,N_14706,N_12399);
nand U18452 (N_18452,N_10639,N_12192);
and U18453 (N_18453,N_12075,N_14810);
nor U18454 (N_18454,N_10402,N_14169);
nor U18455 (N_18455,N_13301,N_10889);
nand U18456 (N_18456,N_11201,N_11577);
nand U18457 (N_18457,N_12876,N_11536);
nor U18458 (N_18458,N_14602,N_13303);
nand U18459 (N_18459,N_12380,N_14244);
nor U18460 (N_18460,N_11752,N_14132);
or U18461 (N_18461,N_10170,N_13076);
or U18462 (N_18462,N_12743,N_11708);
and U18463 (N_18463,N_12892,N_12447);
or U18464 (N_18464,N_10504,N_10456);
nand U18465 (N_18465,N_11917,N_12501);
nand U18466 (N_18466,N_13741,N_13060);
nor U18467 (N_18467,N_14734,N_14831);
nor U18468 (N_18468,N_12492,N_12307);
nor U18469 (N_18469,N_13760,N_14112);
nand U18470 (N_18470,N_10826,N_10494);
and U18471 (N_18471,N_14997,N_13367);
nand U18472 (N_18472,N_10501,N_12679);
nand U18473 (N_18473,N_10914,N_11615);
and U18474 (N_18474,N_11639,N_13903);
and U18475 (N_18475,N_13195,N_11796);
and U18476 (N_18476,N_12289,N_13228);
and U18477 (N_18477,N_10384,N_14046);
xor U18478 (N_18478,N_14295,N_11384);
and U18479 (N_18479,N_13682,N_13228);
and U18480 (N_18480,N_11502,N_14962);
nor U18481 (N_18481,N_13764,N_13672);
and U18482 (N_18482,N_13887,N_13484);
or U18483 (N_18483,N_11268,N_12709);
xnor U18484 (N_18484,N_14235,N_13672);
and U18485 (N_18485,N_14265,N_13621);
nand U18486 (N_18486,N_10592,N_14209);
or U18487 (N_18487,N_11561,N_11633);
or U18488 (N_18488,N_10564,N_11233);
and U18489 (N_18489,N_13965,N_13407);
and U18490 (N_18490,N_11910,N_10860);
and U18491 (N_18491,N_12621,N_11268);
xnor U18492 (N_18492,N_10255,N_13146);
nor U18493 (N_18493,N_14579,N_10653);
or U18494 (N_18494,N_10747,N_13591);
nor U18495 (N_18495,N_11220,N_12808);
xnor U18496 (N_18496,N_11774,N_14466);
and U18497 (N_18497,N_14190,N_14976);
nand U18498 (N_18498,N_13405,N_12517);
and U18499 (N_18499,N_11673,N_14094);
nor U18500 (N_18500,N_10012,N_10990);
and U18501 (N_18501,N_14271,N_14742);
or U18502 (N_18502,N_14093,N_13541);
or U18503 (N_18503,N_12925,N_10044);
and U18504 (N_18504,N_14693,N_13051);
xnor U18505 (N_18505,N_12305,N_10880);
xnor U18506 (N_18506,N_14390,N_14822);
nor U18507 (N_18507,N_14596,N_12484);
or U18508 (N_18508,N_14937,N_11962);
xor U18509 (N_18509,N_11266,N_12651);
nand U18510 (N_18510,N_11224,N_10252);
xnor U18511 (N_18511,N_14268,N_11559);
or U18512 (N_18512,N_11505,N_12264);
and U18513 (N_18513,N_10722,N_12095);
or U18514 (N_18514,N_10001,N_12672);
or U18515 (N_18515,N_12525,N_11198);
or U18516 (N_18516,N_11743,N_10342);
xnor U18517 (N_18517,N_12497,N_13110);
nor U18518 (N_18518,N_11228,N_12236);
nor U18519 (N_18519,N_11869,N_14052);
and U18520 (N_18520,N_14736,N_11674);
nand U18521 (N_18521,N_14903,N_10973);
and U18522 (N_18522,N_10140,N_10868);
nor U18523 (N_18523,N_12983,N_13266);
and U18524 (N_18524,N_10202,N_13738);
and U18525 (N_18525,N_14150,N_14432);
xor U18526 (N_18526,N_13671,N_14922);
and U18527 (N_18527,N_13409,N_12622);
nor U18528 (N_18528,N_12293,N_10666);
nand U18529 (N_18529,N_12169,N_11750);
or U18530 (N_18530,N_12343,N_13646);
or U18531 (N_18531,N_14936,N_10440);
nor U18532 (N_18532,N_13645,N_14753);
nand U18533 (N_18533,N_10150,N_13314);
xor U18534 (N_18534,N_12433,N_12623);
nand U18535 (N_18535,N_12087,N_10302);
and U18536 (N_18536,N_13113,N_11277);
and U18537 (N_18537,N_14417,N_12205);
nand U18538 (N_18538,N_12020,N_14616);
nor U18539 (N_18539,N_14246,N_12488);
xnor U18540 (N_18540,N_12997,N_14478);
or U18541 (N_18541,N_11088,N_11400);
nor U18542 (N_18542,N_12841,N_13649);
nand U18543 (N_18543,N_11245,N_12459);
xor U18544 (N_18544,N_13483,N_11872);
and U18545 (N_18545,N_11040,N_10632);
or U18546 (N_18546,N_13081,N_12786);
xnor U18547 (N_18547,N_10470,N_12918);
and U18548 (N_18548,N_13724,N_10747);
xor U18549 (N_18549,N_10125,N_10052);
or U18550 (N_18550,N_14893,N_13020);
xor U18551 (N_18551,N_10125,N_14533);
or U18552 (N_18552,N_13965,N_11338);
and U18553 (N_18553,N_13603,N_10625);
or U18554 (N_18554,N_14141,N_14156);
xor U18555 (N_18555,N_14083,N_14819);
nand U18556 (N_18556,N_13368,N_14365);
or U18557 (N_18557,N_13017,N_14491);
and U18558 (N_18558,N_13316,N_14817);
xor U18559 (N_18559,N_10514,N_13354);
and U18560 (N_18560,N_11993,N_12980);
or U18561 (N_18561,N_10868,N_14372);
nor U18562 (N_18562,N_11366,N_10238);
nand U18563 (N_18563,N_11176,N_12463);
nor U18564 (N_18564,N_10144,N_10394);
xnor U18565 (N_18565,N_10213,N_11189);
or U18566 (N_18566,N_12357,N_14319);
nand U18567 (N_18567,N_12191,N_11953);
or U18568 (N_18568,N_14776,N_12887);
and U18569 (N_18569,N_11101,N_13129);
and U18570 (N_18570,N_14168,N_12813);
and U18571 (N_18571,N_12210,N_12134);
nand U18572 (N_18572,N_13186,N_13691);
nor U18573 (N_18573,N_10970,N_14444);
or U18574 (N_18574,N_12768,N_14073);
and U18575 (N_18575,N_13440,N_14819);
and U18576 (N_18576,N_10897,N_12517);
nand U18577 (N_18577,N_12048,N_13593);
or U18578 (N_18578,N_14168,N_14818);
nand U18579 (N_18579,N_11471,N_11603);
nand U18580 (N_18580,N_12943,N_12038);
xor U18581 (N_18581,N_14160,N_11648);
nor U18582 (N_18582,N_11442,N_13232);
or U18583 (N_18583,N_13684,N_11019);
nor U18584 (N_18584,N_11718,N_14590);
and U18585 (N_18585,N_14615,N_10553);
nand U18586 (N_18586,N_11615,N_11568);
xor U18587 (N_18587,N_13402,N_10991);
nor U18588 (N_18588,N_10850,N_10202);
or U18589 (N_18589,N_14146,N_14376);
or U18590 (N_18590,N_11826,N_13971);
and U18591 (N_18591,N_13372,N_11593);
xor U18592 (N_18592,N_11534,N_12912);
nand U18593 (N_18593,N_12795,N_11175);
nor U18594 (N_18594,N_10275,N_10435);
and U18595 (N_18595,N_10347,N_14104);
and U18596 (N_18596,N_11694,N_14435);
and U18597 (N_18597,N_14316,N_12553);
and U18598 (N_18598,N_12288,N_11150);
nor U18599 (N_18599,N_10990,N_14457);
xor U18600 (N_18600,N_10880,N_10016);
or U18601 (N_18601,N_12695,N_13309);
or U18602 (N_18602,N_14896,N_10974);
nor U18603 (N_18603,N_11353,N_10375);
nor U18604 (N_18604,N_12779,N_14909);
nand U18605 (N_18605,N_12473,N_14521);
nand U18606 (N_18606,N_14064,N_10256);
xnor U18607 (N_18607,N_11043,N_13886);
nand U18608 (N_18608,N_10472,N_10077);
xor U18609 (N_18609,N_10385,N_11308);
nand U18610 (N_18610,N_12755,N_10112);
and U18611 (N_18611,N_13745,N_14465);
nor U18612 (N_18612,N_12241,N_10981);
nand U18613 (N_18613,N_11860,N_13929);
and U18614 (N_18614,N_13015,N_10643);
xor U18615 (N_18615,N_11344,N_12340);
or U18616 (N_18616,N_11946,N_10903);
and U18617 (N_18617,N_10945,N_14656);
nand U18618 (N_18618,N_10284,N_13412);
and U18619 (N_18619,N_12796,N_13999);
nor U18620 (N_18620,N_11560,N_11084);
or U18621 (N_18621,N_12363,N_13405);
and U18622 (N_18622,N_11629,N_10577);
nor U18623 (N_18623,N_13639,N_11123);
and U18624 (N_18624,N_14072,N_11220);
nor U18625 (N_18625,N_12635,N_10164);
nand U18626 (N_18626,N_12441,N_12563);
xnor U18627 (N_18627,N_14414,N_11888);
xnor U18628 (N_18628,N_10250,N_12729);
nor U18629 (N_18629,N_13897,N_12345);
or U18630 (N_18630,N_13218,N_14718);
or U18631 (N_18631,N_14376,N_14546);
nand U18632 (N_18632,N_10682,N_12934);
and U18633 (N_18633,N_12012,N_13773);
and U18634 (N_18634,N_10443,N_11306);
and U18635 (N_18635,N_14027,N_14844);
and U18636 (N_18636,N_13500,N_12237);
or U18637 (N_18637,N_14265,N_10283);
or U18638 (N_18638,N_13109,N_14631);
and U18639 (N_18639,N_11726,N_11447);
and U18640 (N_18640,N_13804,N_10861);
or U18641 (N_18641,N_11909,N_14939);
and U18642 (N_18642,N_12709,N_14811);
or U18643 (N_18643,N_12369,N_12730);
and U18644 (N_18644,N_11912,N_14779);
xnor U18645 (N_18645,N_12153,N_10306);
nand U18646 (N_18646,N_10185,N_12094);
nand U18647 (N_18647,N_10450,N_14581);
xor U18648 (N_18648,N_13873,N_11047);
xor U18649 (N_18649,N_13326,N_13241);
nand U18650 (N_18650,N_14678,N_14718);
nand U18651 (N_18651,N_12040,N_13302);
xor U18652 (N_18652,N_13876,N_11908);
nand U18653 (N_18653,N_10378,N_10235);
and U18654 (N_18654,N_14267,N_11664);
nand U18655 (N_18655,N_14273,N_10935);
or U18656 (N_18656,N_10836,N_13856);
nand U18657 (N_18657,N_13748,N_11512);
and U18658 (N_18658,N_13904,N_11055);
nand U18659 (N_18659,N_12286,N_14762);
xnor U18660 (N_18660,N_14169,N_11458);
and U18661 (N_18661,N_11115,N_13037);
or U18662 (N_18662,N_14575,N_10236);
nand U18663 (N_18663,N_12698,N_12158);
or U18664 (N_18664,N_11116,N_14693);
xor U18665 (N_18665,N_11895,N_13791);
nor U18666 (N_18666,N_14337,N_11453);
or U18667 (N_18667,N_10254,N_11895);
and U18668 (N_18668,N_10191,N_14150);
xnor U18669 (N_18669,N_14187,N_11786);
xnor U18670 (N_18670,N_12294,N_10443);
nor U18671 (N_18671,N_12293,N_13830);
nor U18672 (N_18672,N_14082,N_13217);
xor U18673 (N_18673,N_14391,N_10204);
xnor U18674 (N_18674,N_12006,N_14667);
nor U18675 (N_18675,N_14362,N_14058);
or U18676 (N_18676,N_14557,N_14127);
and U18677 (N_18677,N_10619,N_14615);
nand U18678 (N_18678,N_11995,N_12580);
nor U18679 (N_18679,N_11929,N_10321);
nand U18680 (N_18680,N_10497,N_12019);
and U18681 (N_18681,N_12778,N_13257);
nor U18682 (N_18682,N_10872,N_10630);
nand U18683 (N_18683,N_14159,N_10780);
xnor U18684 (N_18684,N_12496,N_12246);
nor U18685 (N_18685,N_12911,N_14012);
and U18686 (N_18686,N_12404,N_11289);
nand U18687 (N_18687,N_12686,N_13707);
or U18688 (N_18688,N_14554,N_14692);
nor U18689 (N_18689,N_10595,N_12389);
and U18690 (N_18690,N_10120,N_10366);
or U18691 (N_18691,N_11807,N_11995);
and U18692 (N_18692,N_13862,N_13035);
nor U18693 (N_18693,N_11384,N_10676);
nand U18694 (N_18694,N_12499,N_11795);
nand U18695 (N_18695,N_12239,N_10046);
xor U18696 (N_18696,N_10134,N_12368);
nor U18697 (N_18697,N_13684,N_14523);
xnor U18698 (N_18698,N_10022,N_13206);
or U18699 (N_18699,N_12267,N_10760);
or U18700 (N_18700,N_13981,N_13336);
or U18701 (N_18701,N_10239,N_11393);
nor U18702 (N_18702,N_11712,N_11321);
xnor U18703 (N_18703,N_11635,N_12890);
nand U18704 (N_18704,N_13779,N_11469);
nand U18705 (N_18705,N_10684,N_13792);
nand U18706 (N_18706,N_14995,N_11835);
or U18707 (N_18707,N_13669,N_10975);
and U18708 (N_18708,N_14819,N_13460);
and U18709 (N_18709,N_14717,N_12910);
or U18710 (N_18710,N_13336,N_12242);
nand U18711 (N_18711,N_12598,N_11554);
nor U18712 (N_18712,N_11699,N_14494);
xnor U18713 (N_18713,N_11084,N_10192);
nor U18714 (N_18714,N_14244,N_12093);
nor U18715 (N_18715,N_10790,N_11367);
or U18716 (N_18716,N_13807,N_11040);
nor U18717 (N_18717,N_13942,N_12533);
nand U18718 (N_18718,N_10755,N_14133);
nand U18719 (N_18719,N_14987,N_13357);
and U18720 (N_18720,N_11927,N_11759);
or U18721 (N_18721,N_11958,N_11877);
and U18722 (N_18722,N_12461,N_13606);
nor U18723 (N_18723,N_13872,N_10631);
or U18724 (N_18724,N_12471,N_14849);
nor U18725 (N_18725,N_11935,N_13891);
nor U18726 (N_18726,N_14425,N_10550);
and U18727 (N_18727,N_14006,N_14585);
xor U18728 (N_18728,N_10921,N_12932);
xnor U18729 (N_18729,N_11487,N_13251);
nor U18730 (N_18730,N_14024,N_12065);
or U18731 (N_18731,N_11178,N_13431);
or U18732 (N_18732,N_14569,N_13420);
nor U18733 (N_18733,N_11686,N_13556);
nand U18734 (N_18734,N_12494,N_14907);
and U18735 (N_18735,N_13313,N_12766);
and U18736 (N_18736,N_14709,N_13450);
or U18737 (N_18737,N_12035,N_11432);
and U18738 (N_18738,N_10314,N_14288);
nand U18739 (N_18739,N_11130,N_12301);
nor U18740 (N_18740,N_11638,N_10940);
nor U18741 (N_18741,N_11773,N_11946);
nand U18742 (N_18742,N_13888,N_11317);
xor U18743 (N_18743,N_12587,N_10978);
and U18744 (N_18744,N_10060,N_12096);
xor U18745 (N_18745,N_14535,N_13903);
xor U18746 (N_18746,N_10175,N_14384);
or U18747 (N_18747,N_13552,N_10532);
or U18748 (N_18748,N_13623,N_13063);
nand U18749 (N_18749,N_13406,N_10228);
xor U18750 (N_18750,N_11508,N_14551);
xnor U18751 (N_18751,N_11674,N_13400);
or U18752 (N_18752,N_13678,N_11110);
nand U18753 (N_18753,N_13606,N_13428);
xnor U18754 (N_18754,N_13824,N_12854);
xnor U18755 (N_18755,N_13008,N_10205);
xor U18756 (N_18756,N_13386,N_11315);
or U18757 (N_18757,N_12921,N_10664);
or U18758 (N_18758,N_11369,N_12321);
nand U18759 (N_18759,N_14685,N_10254);
and U18760 (N_18760,N_12814,N_13241);
nor U18761 (N_18761,N_14585,N_13337);
nor U18762 (N_18762,N_13190,N_11709);
and U18763 (N_18763,N_12491,N_14462);
nor U18764 (N_18764,N_13532,N_10183);
and U18765 (N_18765,N_11986,N_13134);
nand U18766 (N_18766,N_12744,N_11426);
and U18767 (N_18767,N_10514,N_14155);
nor U18768 (N_18768,N_11182,N_10665);
nand U18769 (N_18769,N_10840,N_10830);
nor U18770 (N_18770,N_14490,N_11006);
nor U18771 (N_18771,N_13580,N_10570);
xor U18772 (N_18772,N_13937,N_14531);
nor U18773 (N_18773,N_12044,N_13052);
nand U18774 (N_18774,N_10072,N_12578);
xor U18775 (N_18775,N_11202,N_13659);
or U18776 (N_18776,N_10015,N_10860);
nand U18777 (N_18777,N_13015,N_12312);
and U18778 (N_18778,N_12573,N_11887);
nand U18779 (N_18779,N_14646,N_11194);
xnor U18780 (N_18780,N_12994,N_11397);
nor U18781 (N_18781,N_12223,N_10813);
nor U18782 (N_18782,N_11010,N_12028);
and U18783 (N_18783,N_12178,N_11623);
nand U18784 (N_18784,N_12640,N_10944);
nor U18785 (N_18785,N_13818,N_10647);
or U18786 (N_18786,N_14912,N_11040);
xor U18787 (N_18787,N_10669,N_11057);
and U18788 (N_18788,N_12211,N_14609);
and U18789 (N_18789,N_12934,N_11247);
and U18790 (N_18790,N_10123,N_13716);
and U18791 (N_18791,N_12950,N_13349);
or U18792 (N_18792,N_12116,N_14574);
nor U18793 (N_18793,N_14308,N_10969);
nand U18794 (N_18794,N_11895,N_12942);
nor U18795 (N_18795,N_11018,N_14495);
nand U18796 (N_18796,N_11896,N_12397);
nor U18797 (N_18797,N_12937,N_10566);
and U18798 (N_18798,N_11937,N_12268);
and U18799 (N_18799,N_14002,N_10961);
nor U18800 (N_18800,N_12149,N_13129);
nor U18801 (N_18801,N_10250,N_13126);
xnor U18802 (N_18802,N_13788,N_13385);
or U18803 (N_18803,N_14083,N_13750);
nand U18804 (N_18804,N_14850,N_10101);
xnor U18805 (N_18805,N_13103,N_13030);
or U18806 (N_18806,N_10354,N_14140);
nand U18807 (N_18807,N_13069,N_14104);
nand U18808 (N_18808,N_11754,N_13288);
and U18809 (N_18809,N_13149,N_14001);
nand U18810 (N_18810,N_14911,N_10141);
nor U18811 (N_18811,N_11291,N_11272);
and U18812 (N_18812,N_14741,N_12168);
and U18813 (N_18813,N_10462,N_14065);
nor U18814 (N_18814,N_13110,N_10794);
or U18815 (N_18815,N_11302,N_12254);
xnor U18816 (N_18816,N_13777,N_13673);
and U18817 (N_18817,N_14549,N_14716);
nor U18818 (N_18818,N_14273,N_14066);
or U18819 (N_18819,N_13108,N_14712);
or U18820 (N_18820,N_10130,N_11345);
xnor U18821 (N_18821,N_11764,N_14713);
nand U18822 (N_18822,N_13274,N_10979);
or U18823 (N_18823,N_13742,N_13038);
and U18824 (N_18824,N_12760,N_11901);
or U18825 (N_18825,N_10665,N_13207);
or U18826 (N_18826,N_10551,N_13649);
xor U18827 (N_18827,N_12175,N_12588);
nand U18828 (N_18828,N_12829,N_14864);
and U18829 (N_18829,N_10986,N_13340);
or U18830 (N_18830,N_11063,N_14089);
xor U18831 (N_18831,N_14356,N_10835);
nand U18832 (N_18832,N_12162,N_11622);
and U18833 (N_18833,N_14318,N_11403);
nor U18834 (N_18834,N_12325,N_11067);
and U18835 (N_18835,N_14639,N_10622);
nand U18836 (N_18836,N_13739,N_10076);
nand U18837 (N_18837,N_12862,N_10843);
and U18838 (N_18838,N_12805,N_13772);
xnor U18839 (N_18839,N_12256,N_13309);
nor U18840 (N_18840,N_10255,N_13261);
nor U18841 (N_18841,N_13576,N_13866);
xor U18842 (N_18842,N_12801,N_14131);
xnor U18843 (N_18843,N_14699,N_14945);
nor U18844 (N_18844,N_14657,N_11727);
nand U18845 (N_18845,N_12198,N_12492);
and U18846 (N_18846,N_11567,N_11781);
nand U18847 (N_18847,N_11213,N_11481);
or U18848 (N_18848,N_11150,N_10454);
nand U18849 (N_18849,N_14040,N_10426);
nor U18850 (N_18850,N_10864,N_12515);
nand U18851 (N_18851,N_10467,N_11664);
and U18852 (N_18852,N_14536,N_12037);
nor U18853 (N_18853,N_11202,N_14382);
xnor U18854 (N_18854,N_13148,N_11403);
xor U18855 (N_18855,N_14575,N_14555);
nand U18856 (N_18856,N_13040,N_13062);
and U18857 (N_18857,N_12573,N_13665);
or U18858 (N_18858,N_10120,N_14470);
or U18859 (N_18859,N_10704,N_11480);
nor U18860 (N_18860,N_10180,N_13595);
xnor U18861 (N_18861,N_10620,N_10812);
nand U18862 (N_18862,N_13304,N_12871);
or U18863 (N_18863,N_14632,N_12478);
xnor U18864 (N_18864,N_13020,N_12445);
nor U18865 (N_18865,N_14648,N_14751);
xor U18866 (N_18866,N_13021,N_13035);
nand U18867 (N_18867,N_14911,N_13043);
nor U18868 (N_18868,N_10531,N_10021);
or U18869 (N_18869,N_14182,N_14848);
or U18870 (N_18870,N_11494,N_12926);
and U18871 (N_18871,N_11655,N_14092);
or U18872 (N_18872,N_13711,N_11533);
nand U18873 (N_18873,N_14377,N_11953);
and U18874 (N_18874,N_13890,N_11658);
nor U18875 (N_18875,N_10060,N_12308);
and U18876 (N_18876,N_11463,N_13631);
nor U18877 (N_18877,N_13453,N_12417);
and U18878 (N_18878,N_12331,N_13431);
nand U18879 (N_18879,N_11003,N_13344);
xnor U18880 (N_18880,N_10978,N_13111);
nand U18881 (N_18881,N_13065,N_14803);
nand U18882 (N_18882,N_14484,N_14704);
and U18883 (N_18883,N_11532,N_10348);
nor U18884 (N_18884,N_11706,N_14850);
nand U18885 (N_18885,N_11285,N_14679);
and U18886 (N_18886,N_10643,N_13913);
nor U18887 (N_18887,N_12741,N_13535);
or U18888 (N_18888,N_12796,N_13248);
and U18889 (N_18889,N_14357,N_10606);
or U18890 (N_18890,N_11845,N_10726);
xor U18891 (N_18891,N_13707,N_11943);
or U18892 (N_18892,N_10077,N_11840);
xor U18893 (N_18893,N_12968,N_12041);
xor U18894 (N_18894,N_12923,N_11027);
nor U18895 (N_18895,N_14822,N_10690);
or U18896 (N_18896,N_14547,N_13257);
and U18897 (N_18897,N_13073,N_14928);
xnor U18898 (N_18898,N_14725,N_11201);
nor U18899 (N_18899,N_12969,N_11665);
xor U18900 (N_18900,N_11590,N_10362);
nor U18901 (N_18901,N_10951,N_13633);
or U18902 (N_18902,N_14324,N_14395);
nand U18903 (N_18903,N_12896,N_12422);
nor U18904 (N_18904,N_10865,N_14490);
or U18905 (N_18905,N_12196,N_14430);
nand U18906 (N_18906,N_10177,N_10292);
nand U18907 (N_18907,N_10595,N_14350);
nand U18908 (N_18908,N_11982,N_11213);
nand U18909 (N_18909,N_11341,N_13780);
xor U18910 (N_18910,N_10900,N_13606);
nor U18911 (N_18911,N_14950,N_11514);
or U18912 (N_18912,N_14168,N_10626);
nor U18913 (N_18913,N_13421,N_14411);
and U18914 (N_18914,N_11241,N_11566);
nor U18915 (N_18915,N_14868,N_14699);
nor U18916 (N_18916,N_12648,N_11664);
or U18917 (N_18917,N_14026,N_11669);
or U18918 (N_18918,N_12343,N_12666);
or U18919 (N_18919,N_13361,N_10427);
nor U18920 (N_18920,N_10721,N_10256);
xnor U18921 (N_18921,N_11253,N_10737);
nand U18922 (N_18922,N_13089,N_13195);
nor U18923 (N_18923,N_11316,N_10247);
nand U18924 (N_18924,N_11045,N_11769);
xor U18925 (N_18925,N_13022,N_11945);
and U18926 (N_18926,N_11638,N_13470);
nor U18927 (N_18927,N_12775,N_10247);
nor U18928 (N_18928,N_14723,N_12414);
and U18929 (N_18929,N_11776,N_14964);
and U18930 (N_18930,N_14162,N_13350);
nand U18931 (N_18931,N_14692,N_14704);
nor U18932 (N_18932,N_13753,N_11449);
xnor U18933 (N_18933,N_10029,N_11405);
nand U18934 (N_18934,N_10590,N_14469);
nor U18935 (N_18935,N_10904,N_12792);
nor U18936 (N_18936,N_13970,N_12202);
nor U18937 (N_18937,N_11432,N_14828);
xnor U18938 (N_18938,N_11538,N_13792);
nand U18939 (N_18939,N_10799,N_10239);
nand U18940 (N_18940,N_10461,N_11261);
nor U18941 (N_18941,N_11312,N_13691);
and U18942 (N_18942,N_13984,N_12069);
xnor U18943 (N_18943,N_14306,N_12192);
or U18944 (N_18944,N_13023,N_10226);
or U18945 (N_18945,N_12720,N_11115);
xnor U18946 (N_18946,N_11717,N_11494);
nor U18947 (N_18947,N_10108,N_11616);
xnor U18948 (N_18948,N_13721,N_14249);
nor U18949 (N_18949,N_13527,N_14967);
and U18950 (N_18950,N_12713,N_11631);
nand U18951 (N_18951,N_13357,N_14980);
and U18952 (N_18952,N_11782,N_14118);
or U18953 (N_18953,N_11065,N_10527);
xnor U18954 (N_18954,N_12670,N_14862);
or U18955 (N_18955,N_12408,N_11407);
or U18956 (N_18956,N_14454,N_12387);
nor U18957 (N_18957,N_14025,N_11949);
nor U18958 (N_18958,N_10077,N_13420);
nand U18959 (N_18959,N_11484,N_13128);
xnor U18960 (N_18960,N_12223,N_12942);
nand U18961 (N_18961,N_13188,N_12005);
and U18962 (N_18962,N_14323,N_10761);
or U18963 (N_18963,N_11117,N_13652);
and U18964 (N_18964,N_13008,N_12018);
or U18965 (N_18965,N_11364,N_11944);
nor U18966 (N_18966,N_13979,N_13182);
nor U18967 (N_18967,N_13452,N_13065);
nand U18968 (N_18968,N_14536,N_14059);
and U18969 (N_18969,N_12064,N_11810);
xor U18970 (N_18970,N_12565,N_11586);
nor U18971 (N_18971,N_10147,N_10485);
nor U18972 (N_18972,N_14123,N_11570);
nand U18973 (N_18973,N_14831,N_12351);
nand U18974 (N_18974,N_13363,N_12572);
nor U18975 (N_18975,N_11327,N_13730);
and U18976 (N_18976,N_11093,N_11801);
or U18977 (N_18977,N_11812,N_14079);
or U18978 (N_18978,N_10244,N_10249);
xnor U18979 (N_18979,N_12732,N_11567);
nor U18980 (N_18980,N_10697,N_12833);
xnor U18981 (N_18981,N_12640,N_11947);
and U18982 (N_18982,N_11719,N_11567);
nor U18983 (N_18983,N_13074,N_11434);
nand U18984 (N_18984,N_13122,N_11667);
nor U18985 (N_18985,N_14375,N_12125);
or U18986 (N_18986,N_14494,N_11727);
nand U18987 (N_18987,N_11084,N_12195);
nand U18988 (N_18988,N_12956,N_11956);
nor U18989 (N_18989,N_14933,N_11680);
nor U18990 (N_18990,N_12590,N_12281);
nand U18991 (N_18991,N_14624,N_12538);
xor U18992 (N_18992,N_10214,N_12871);
or U18993 (N_18993,N_13628,N_11894);
or U18994 (N_18994,N_12839,N_11471);
xor U18995 (N_18995,N_13700,N_11644);
or U18996 (N_18996,N_12279,N_11120);
nand U18997 (N_18997,N_11632,N_12024);
nor U18998 (N_18998,N_12704,N_13583);
xor U18999 (N_18999,N_11506,N_12745);
xor U19000 (N_19000,N_12650,N_12967);
and U19001 (N_19001,N_12766,N_14059);
xor U19002 (N_19002,N_11792,N_13046);
and U19003 (N_19003,N_14902,N_11364);
xnor U19004 (N_19004,N_12414,N_12169);
or U19005 (N_19005,N_14895,N_14365);
and U19006 (N_19006,N_12662,N_12136);
or U19007 (N_19007,N_13388,N_12413);
and U19008 (N_19008,N_12192,N_14076);
or U19009 (N_19009,N_10897,N_14002);
or U19010 (N_19010,N_10594,N_13420);
nor U19011 (N_19011,N_10867,N_10634);
nand U19012 (N_19012,N_10496,N_12943);
nand U19013 (N_19013,N_14075,N_14766);
and U19014 (N_19014,N_13094,N_10749);
xor U19015 (N_19015,N_13374,N_12594);
or U19016 (N_19016,N_12367,N_12358);
nand U19017 (N_19017,N_14990,N_10681);
nand U19018 (N_19018,N_10076,N_13908);
nand U19019 (N_19019,N_10454,N_14029);
nor U19020 (N_19020,N_13803,N_10862);
xnor U19021 (N_19021,N_12163,N_13855);
nand U19022 (N_19022,N_11538,N_10123);
nor U19023 (N_19023,N_13040,N_14289);
xnor U19024 (N_19024,N_10445,N_13992);
and U19025 (N_19025,N_11228,N_10020);
and U19026 (N_19026,N_11897,N_14052);
or U19027 (N_19027,N_10199,N_13007);
nand U19028 (N_19028,N_13380,N_12555);
or U19029 (N_19029,N_10733,N_10430);
xor U19030 (N_19030,N_11169,N_10750);
nor U19031 (N_19031,N_11443,N_13769);
xor U19032 (N_19032,N_11449,N_14155);
nor U19033 (N_19033,N_12308,N_11636);
or U19034 (N_19034,N_10534,N_13302);
and U19035 (N_19035,N_10256,N_14019);
xnor U19036 (N_19036,N_11508,N_12870);
or U19037 (N_19037,N_13126,N_10605);
nand U19038 (N_19038,N_10292,N_12706);
and U19039 (N_19039,N_12014,N_13764);
xor U19040 (N_19040,N_11725,N_14782);
xnor U19041 (N_19041,N_12594,N_10576);
nand U19042 (N_19042,N_13426,N_11116);
nand U19043 (N_19043,N_13020,N_12121);
or U19044 (N_19044,N_11988,N_14996);
xor U19045 (N_19045,N_13067,N_13967);
nor U19046 (N_19046,N_12819,N_11539);
and U19047 (N_19047,N_11668,N_10896);
or U19048 (N_19048,N_12332,N_14205);
xnor U19049 (N_19049,N_12549,N_14353);
xor U19050 (N_19050,N_13515,N_11848);
nor U19051 (N_19051,N_14764,N_11231);
or U19052 (N_19052,N_12913,N_10415);
or U19053 (N_19053,N_10142,N_13574);
xor U19054 (N_19054,N_11191,N_11959);
or U19055 (N_19055,N_11894,N_14372);
nor U19056 (N_19056,N_14934,N_12473);
or U19057 (N_19057,N_11597,N_10568);
and U19058 (N_19058,N_10956,N_12646);
xor U19059 (N_19059,N_14771,N_12782);
nor U19060 (N_19060,N_13152,N_11438);
xnor U19061 (N_19061,N_12350,N_13239);
or U19062 (N_19062,N_13955,N_14156);
nor U19063 (N_19063,N_10953,N_13237);
nor U19064 (N_19064,N_10389,N_11420);
xnor U19065 (N_19065,N_13347,N_11076);
nor U19066 (N_19066,N_13817,N_13716);
nand U19067 (N_19067,N_14677,N_11058);
xor U19068 (N_19068,N_14751,N_12877);
or U19069 (N_19069,N_13166,N_11344);
nand U19070 (N_19070,N_13166,N_10923);
nor U19071 (N_19071,N_10715,N_13190);
nand U19072 (N_19072,N_13805,N_14066);
xnor U19073 (N_19073,N_13487,N_12033);
xor U19074 (N_19074,N_14884,N_10172);
nand U19075 (N_19075,N_12451,N_12915);
or U19076 (N_19076,N_12769,N_12056);
xnor U19077 (N_19077,N_14039,N_13281);
nor U19078 (N_19078,N_14808,N_11935);
nor U19079 (N_19079,N_11891,N_13161);
nor U19080 (N_19080,N_11108,N_13229);
nand U19081 (N_19081,N_11322,N_11225);
or U19082 (N_19082,N_12102,N_14922);
and U19083 (N_19083,N_10500,N_14753);
and U19084 (N_19084,N_10342,N_13018);
xor U19085 (N_19085,N_12401,N_14749);
nand U19086 (N_19086,N_10231,N_13799);
nand U19087 (N_19087,N_11340,N_13895);
xor U19088 (N_19088,N_14104,N_10618);
and U19089 (N_19089,N_13702,N_10294);
or U19090 (N_19090,N_10355,N_10273);
nand U19091 (N_19091,N_12578,N_14872);
or U19092 (N_19092,N_12400,N_12692);
xnor U19093 (N_19093,N_13183,N_14618);
and U19094 (N_19094,N_14336,N_10386);
nor U19095 (N_19095,N_11388,N_13536);
nand U19096 (N_19096,N_11074,N_10573);
nand U19097 (N_19097,N_10129,N_14534);
or U19098 (N_19098,N_11333,N_11695);
nand U19099 (N_19099,N_12836,N_11970);
and U19100 (N_19100,N_11139,N_14377);
nand U19101 (N_19101,N_10286,N_10238);
nor U19102 (N_19102,N_13902,N_14010);
nor U19103 (N_19103,N_13610,N_14949);
and U19104 (N_19104,N_13379,N_11155);
and U19105 (N_19105,N_12234,N_10095);
xor U19106 (N_19106,N_10475,N_13283);
xor U19107 (N_19107,N_14287,N_10550);
nand U19108 (N_19108,N_12808,N_10492);
xor U19109 (N_19109,N_14274,N_14540);
nand U19110 (N_19110,N_12326,N_13209);
nor U19111 (N_19111,N_11396,N_10279);
xor U19112 (N_19112,N_11577,N_14145);
or U19113 (N_19113,N_11128,N_11792);
and U19114 (N_19114,N_14386,N_13357);
nand U19115 (N_19115,N_13934,N_10950);
and U19116 (N_19116,N_12135,N_14686);
or U19117 (N_19117,N_13359,N_10857);
nand U19118 (N_19118,N_10883,N_10760);
nor U19119 (N_19119,N_11026,N_13512);
xor U19120 (N_19120,N_11976,N_11508);
nor U19121 (N_19121,N_14591,N_12059);
nand U19122 (N_19122,N_13767,N_13324);
and U19123 (N_19123,N_14233,N_14327);
xnor U19124 (N_19124,N_14425,N_13430);
nor U19125 (N_19125,N_14639,N_13456);
or U19126 (N_19126,N_12510,N_11367);
or U19127 (N_19127,N_12215,N_10233);
and U19128 (N_19128,N_11975,N_14802);
nor U19129 (N_19129,N_13668,N_14247);
or U19130 (N_19130,N_10928,N_14292);
nand U19131 (N_19131,N_11591,N_12588);
nand U19132 (N_19132,N_14830,N_11567);
and U19133 (N_19133,N_13937,N_13961);
or U19134 (N_19134,N_10829,N_12032);
nand U19135 (N_19135,N_14044,N_13419);
nor U19136 (N_19136,N_14132,N_14814);
or U19137 (N_19137,N_12171,N_12251);
and U19138 (N_19138,N_14465,N_11452);
or U19139 (N_19139,N_13191,N_11316);
nand U19140 (N_19140,N_12202,N_14028);
nor U19141 (N_19141,N_14134,N_14287);
or U19142 (N_19142,N_14961,N_13485);
or U19143 (N_19143,N_13983,N_10379);
nand U19144 (N_19144,N_14657,N_10377);
and U19145 (N_19145,N_14330,N_13333);
nand U19146 (N_19146,N_12933,N_14884);
xor U19147 (N_19147,N_11076,N_14280);
and U19148 (N_19148,N_13764,N_13378);
nand U19149 (N_19149,N_12686,N_10225);
or U19150 (N_19150,N_11726,N_14719);
or U19151 (N_19151,N_14517,N_11956);
nand U19152 (N_19152,N_14341,N_10544);
nand U19153 (N_19153,N_11996,N_12239);
and U19154 (N_19154,N_12543,N_13484);
nand U19155 (N_19155,N_13179,N_11343);
nand U19156 (N_19156,N_12283,N_14293);
nand U19157 (N_19157,N_13849,N_12450);
and U19158 (N_19158,N_11048,N_11853);
or U19159 (N_19159,N_10257,N_10492);
nor U19160 (N_19160,N_11095,N_11891);
xor U19161 (N_19161,N_12577,N_10615);
or U19162 (N_19162,N_11090,N_10219);
nor U19163 (N_19163,N_14536,N_11679);
nor U19164 (N_19164,N_14337,N_12545);
xnor U19165 (N_19165,N_10178,N_14515);
nand U19166 (N_19166,N_14177,N_10345);
nand U19167 (N_19167,N_10298,N_10237);
or U19168 (N_19168,N_14406,N_14009);
and U19169 (N_19169,N_11211,N_10976);
nand U19170 (N_19170,N_14109,N_10433);
nand U19171 (N_19171,N_11231,N_12849);
and U19172 (N_19172,N_14578,N_14293);
xnor U19173 (N_19173,N_11465,N_11373);
xor U19174 (N_19174,N_11170,N_12778);
or U19175 (N_19175,N_13445,N_11121);
or U19176 (N_19176,N_14419,N_12597);
nand U19177 (N_19177,N_12299,N_10986);
and U19178 (N_19178,N_12925,N_14141);
nand U19179 (N_19179,N_10057,N_12228);
and U19180 (N_19180,N_10966,N_14077);
and U19181 (N_19181,N_12379,N_13935);
and U19182 (N_19182,N_12124,N_14777);
nor U19183 (N_19183,N_11480,N_10878);
xor U19184 (N_19184,N_12973,N_12198);
and U19185 (N_19185,N_13765,N_14546);
or U19186 (N_19186,N_11000,N_10027);
and U19187 (N_19187,N_10438,N_12229);
or U19188 (N_19188,N_13173,N_12242);
or U19189 (N_19189,N_12218,N_10732);
and U19190 (N_19190,N_14052,N_12683);
or U19191 (N_19191,N_14256,N_12660);
nand U19192 (N_19192,N_10579,N_13452);
and U19193 (N_19193,N_14254,N_14750);
nand U19194 (N_19194,N_14015,N_10784);
xor U19195 (N_19195,N_11956,N_10911);
xnor U19196 (N_19196,N_10536,N_10899);
and U19197 (N_19197,N_11394,N_12396);
xor U19198 (N_19198,N_12272,N_13913);
nor U19199 (N_19199,N_10712,N_14687);
and U19200 (N_19200,N_14612,N_10684);
nor U19201 (N_19201,N_11214,N_12731);
nand U19202 (N_19202,N_10477,N_11935);
nand U19203 (N_19203,N_13179,N_14528);
nand U19204 (N_19204,N_12069,N_12765);
nand U19205 (N_19205,N_10239,N_14484);
and U19206 (N_19206,N_14341,N_11464);
nor U19207 (N_19207,N_11982,N_14282);
nor U19208 (N_19208,N_13379,N_10816);
xnor U19209 (N_19209,N_13823,N_11564);
xnor U19210 (N_19210,N_13113,N_11065);
or U19211 (N_19211,N_10608,N_11720);
or U19212 (N_19212,N_10273,N_12997);
or U19213 (N_19213,N_12766,N_12997);
and U19214 (N_19214,N_13100,N_13185);
xnor U19215 (N_19215,N_12019,N_14268);
nor U19216 (N_19216,N_14610,N_14520);
xnor U19217 (N_19217,N_13678,N_11206);
or U19218 (N_19218,N_13578,N_10095);
xor U19219 (N_19219,N_11747,N_14393);
xor U19220 (N_19220,N_10798,N_14762);
nor U19221 (N_19221,N_13309,N_12241);
xnor U19222 (N_19222,N_14551,N_12206);
nand U19223 (N_19223,N_14638,N_10675);
or U19224 (N_19224,N_10693,N_13119);
nand U19225 (N_19225,N_11214,N_11903);
nand U19226 (N_19226,N_11225,N_11478);
or U19227 (N_19227,N_12832,N_12154);
and U19228 (N_19228,N_13175,N_13858);
xor U19229 (N_19229,N_11323,N_14366);
nand U19230 (N_19230,N_13537,N_13491);
nand U19231 (N_19231,N_14004,N_11460);
nand U19232 (N_19232,N_10028,N_11362);
or U19233 (N_19233,N_10989,N_12754);
xor U19234 (N_19234,N_12535,N_14739);
nand U19235 (N_19235,N_10548,N_13449);
nor U19236 (N_19236,N_12956,N_12820);
nor U19237 (N_19237,N_13177,N_14166);
and U19238 (N_19238,N_11843,N_12277);
nor U19239 (N_19239,N_13234,N_10958);
and U19240 (N_19240,N_13416,N_12906);
or U19241 (N_19241,N_10709,N_12954);
nand U19242 (N_19242,N_14522,N_14776);
xnor U19243 (N_19243,N_11300,N_13788);
nand U19244 (N_19244,N_14283,N_11240);
or U19245 (N_19245,N_10794,N_11833);
and U19246 (N_19246,N_10579,N_14058);
nor U19247 (N_19247,N_14264,N_14247);
or U19248 (N_19248,N_13905,N_13097);
and U19249 (N_19249,N_14124,N_13842);
nor U19250 (N_19250,N_11913,N_11027);
nand U19251 (N_19251,N_14175,N_14242);
nand U19252 (N_19252,N_14575,N_13095);
nor U19253 (N_19253,N_10247,N_12613);
nand U19254 (N_19254,N_10998,N_10778);
nand U19255 (N_19255,N_13670,N_12292);
xor U19256 (N_19256,N_12030,N_13554);
and U19257 (N_19257,N_10131,N_13727);
nand U19258 (N_19258,N_14980,N_11198);
nand U19259 (N_19259,N_10210,N_13184);
and U19260 (N_19260,N_14155,N_14648);
nand U19261 (N_19261,N_10132,N_10644);
or U19262 (N_19262,N_11220,N_13980);
nand U19263 (N_19263,N_14369,N_10179);
nand U19264 (N_19264,N_12832,N_11016);
xor U19265 (N_19265,N_14398,N_14660);
and U19266 (N_19266,N_12260,N_10800);
nor U19267 (N_19267,N_11712,N_13501);
or U19268 (N_19268,N_10307,N_14618);
nor U19269 (N_19269,N_10075,N_10443);
and U19270 (N_19270,N_11751,N_13086);
nand U19271 (N_19271,N_12298,N_12584);
nor U19272 (N_19272,N_14956,N_10213);
xor U19273 (N_19273,N_11229,N_13482);
nand U19274 (N_19274,N_10100,N_12479);
nand U19275 (N_19275,N_11432,N_13263);
nand U19276 (N_19276,N_10029,N_12247);
nor U19277 (N_19277,N_12652,N_12886);
xor U19278 (N_19278,N_10449,N_14978);
and U19279 (N_19279,N_14950,N_14791);
nand U19280 (N_19280,N_13088,N_13834);
nand U19281 (N_19281,N_12661,N_14396);
xnor U19282 (N_19282,N_10925,N_13825);
xnor U19283 (N_19283,N_11278,N_13646);
nand U19284 (N_19284,N_11352,N_13123);
nand U19285 (N_19285,N_13422,N_14889);
or U19286 (N_19286,N_10120,N_12073);
or U19287 (N_19287,N_14310,N_10740);
nand U19288 (N_19288,N_12434,N_10885);
xor U19289 (N_19289,N_14895,N_13129);
nor U19290 (N_19290,N_12644,N_12485);
and U19291 (N_19291,N_11651,N_14730);
nor U19292 (N_19292,N_14918,N_14240);
xnor U19293 (N_19293,N_12709,N_13330);
and U19294 (N_19294,N_14075,N_12505);
nor U19295 (N_19295,N_12276,N_11152);
or U19296 (N_19296,N_13423,N_12138);
xor U19297 (N_19297,N_13246,N_12711);
and U19298 (N_19298,N_12381,N_13371);
and U19299 (N_19299,N_14831,N_11807);
nor U19300 (N_19300,N_10142,N_12622);
xor U19301 (N_19301,N_13488,N_11088);
and U19302 (N_19302,N_12377,N_14756);
nor U19303 (N_19303,N_11631,N_12499);
xor U19304 (N_19304,N_13256,N_12116);
nor U19305 (N_19305,N_13335,N_14661);
or U19306 (N_19306,N_10411,N_12359);
nor U19307 (N_19307,N_13318,N_11721);
xnor U19308 (N_19308,N_11333,N_11028);
nand U19309 (N_19309,N_10762,N_12457);
or U19310 (N_19310,N_14242,N_10863);
nand U19311 (N_19311,N_12638,N_10416);
and U19312 (N_19312,N_10748,N_13718);
xnor U19313 (N_19313,N_12884,N_10256);
or U19314 (N_19314,N_12539,N_13227);
and U19315 (N_19315,N_12652,N_10631);
and U19316 (N_19316,N_10008,N_10552);
and U19317 (N_19317,N_13834,N_10332);
xnor U19318 (N_19318,N_14882,N_11796);
xor U19319 (N_19319,N_10461,N_10892);
and U19320 (N_19320,N_12512,N_11549);
nor U19321 (N_19321,N_14165,N_10267);
xor U19322 (N_19322,N_11434,N_14071);
or U19323 (N_19323,N_14577,N_13013);
or U19324 (N_19324,N_14921,N_14299);
and U19325 (N_19325,N_12392,N_13122);
nand U19326 (N_19326,N_14902,N_10160);
nor U19327 (N_19327,N_10713,N_11506);
nor U19328 (N_19328,N_13884,N_10940);
xnor U19329 (N_19329,N_14858,N_10380);
or U19330 (N_19330,N_13878,N_10936);
xnor U19331 (N_19331,N_14344,N_12972);
xnor U19332 (N_19332,N_12034,N_11240);
and U19333 (N_19333,N_11538,N_11618);
or U19334 (N_19334,N_12214,N_11106);
and U19335 (N_19335,N_14397,N_12887);
and U19336 (N_19336,N_12572,N_13571);
and U19337 (N_19337,N_10688,N_12103);
and U19338 (N_19338,N_14845,N_10105);
or U19339 (N_19339,N_13537,N_12595);
nor U19340 (N_19340,N_14047,N_10637);
nor U19341 (N_19341,N_14145,N_13695);
xnor U19342 (N_19342,N_14362,N_11756);
or U19343 (N_19343,N_11831,N_12904);
xnor U19344 (N_19344,N_12246,N_14686);
xor U19345 (N_19345,N_12841,N_12664);
xor U19346 (N_19346,N_13301,N_14925);
or U19347 (N_19347,N_10632,N_10171);
xnor U19348 (N_19348,N_10275,N_11717);
nand U19349 (N_19349,N_14062,N_12153);
and U19350 (N_19350,N_10585,N_13966);
or U19351 (N_19351,N_10729,N_11777);
nor U19352 (N_19352,N_12709,N_14689);
or U19353 (N_19353,N_11858,N_11392);
nand U19354 (N_19354,N_11633,N_14900);
nor U19355 (N_19355,N_14176,N_10361);
nor U19356 (N_19356,N_14712,N_14280);
nand U19357 (N_19357,N_14558,N_10402);
nand U19358 (N_19358,N_11268,N_13840);
nand U19359 (N_19359,N_14880,N_10580);
nor U19360 (N_19360,N_13972,N_12852);
and U19361 (N_19361,N_14028,N_13295);
and U19362 (N_19362,N_10439,N_12419);
and U19363 (N_19363,N_14473,N_14066);
or U19364 (N_19364,N_11572,N_12426);
nor U19365 (N_19365,N_11396,N_11591);
or U19366 (N_19366,N_11668,N_11074);
nand U19367 (N_19367,N_13901,N_14120);
nor U19368 (N_19368,N_13759,N_14446);
and U19369 (N_19369,N_14219,N_13041);
or U19370 (N_19370,N_12471,N_13045);
nand U19371 (N_19371,N_11357,N_12372);
and U19372 (N_19372,N_11535,N_12747);
nand U19373 (N_19373,N_14221,N_13915);
and U19374 (N_19374,N_13660,N_13733);
nand U19375 (N_19375,N_10874,N_13006);
nor U19376 (N_19376,N_10584,N_13608);
and U19377 (N_19377,N_11365,N_11985);
or U19378 (N_19378,N_11471,N_12466);
xnor U19379 (N_19379,N_14721,N_13815);
xnor U19380 (N_19380,N_12389,N_10104);
and U19381 (N_19381,N_14483,N_14283);
or U19382 (N_19382,N_12488,N_10330);
or U19383 (N_19383,N_10739,N_10024);
and U19384 (N_19384,N_10046,N_12352);
xor U19385 (N_19385,N_10250,N_13612);
xor U19386 (N_19386,N_11444,N_13663);
xnor U19387 (N_19387,N_12014,N_12421);
nor U19388 (N_19388,N_12724,N_14851);
or U19389 (N_19389,N_11237,N_10842);
nor U19390 (N_19390,N_13150,N_10033);
and U19391 (N_19391,N_13291,N_13098);
or U19392 (N_19392,N_11055,N_12145);
xor U19393 (N_19393,N_13498,N_10027);
or U19394 (N_19394,N_12523,N_10385);
nand U19395 (N_19395,N_12828,N_11140);
or U19396 (N_19396,N_11705,N_12193);
and U19397 (N_19397,N_10665,N_13684);
xor U19398 (N_19398,N_11812,N_14756);
xor U19399 (N_19399,N_10694,N_14975);
nor U19400 (N_19400,N_12671,N_13037);
nor U19401 (N_19401,N_10703,N_13423);
xnor U19402 (N_19402,N_14522,N_12865);
xor U19403 (N_19403,N_14625,N_13924);
xnor U19404 (N_19404,N_14243,N_14739);
nor U19405 (N_19405,N_11844,N_13178);
or U19406 (N_19406,N_11896,N_12481);
or U19407 (N_19407,N_11173,N_12509);
nand U19408 (N_19408,N_11702,N_11267);
xor U19409 (N_19409,N_10754,N_13790);
nand U19410 (N_19410,N_14150,N_10363);
and U19411 (N_19411,N_13941,N_14269);
nor U19412 (N_19412,N_10863,N_14463);
and U19413 (N_19413,N_11412,N_14405);
nor U19414 (N_19414,N_14891,N_11538);
and U19415 (N_19415,N_14982,N_11515);
xnor U19416 (N_19416,N_10849,N_14927);
or U19417 (N_19417,N_13172,N_13248);
or U19418 (N_19418,N_12379,N_10535);
nand U19419 (N_19419,N_12993,N_10431);
or U19420 (N_19420,N_10690,N_10043);
and U19421 (N_19421,N_10838,N_14780);
and U19422 (N_19422,N_13318,N_14161);
nor U19423 (N_19423,N_10212,N_13831);
xnor U19424 (N_19424,N_12770,N_10986);
xnor U19425 (N_19425,N_11172,N_10471);
and U19426 (N_19426,N_10295,N_13557);
and U19427 (N_19427,N_14876,N_11138);
xor U19428 (N_19428,N_10390,N_10816);
xnor U19429 (N_19429,N_13193,N_11218);
and U19430 (N_19430,N_13687,N_14352);
and U19431 (N_19431,N_13337,N_11357);
nor U19432 (N_19432,N_12520,N_10478);
nor U19433 (N_19433,N_14582,N_12881);
or U19434 (N_19434,N_11059,N_10698);
or U19435 (N_19435,N_13519,N_10768);
and U19436 (N_19436,N_13730,N_10294);
nor U19437 (N_19437,N_14153,N_13746);
or U19438 (N_19438,N_11962,N_10645);
and U19439 (N_19439,N_14908,N_13422);
nand U19440 (N_19440,N_10331,N_13229);
nand U19441 (N_19441,N_11623,N_14612);
or U19442 (N_19442,N_11441,N_10076);
nor U19443 (N_19443,N_10407,N_12394);
or U19444 (N_19444,N_11989,N_14085);
or U19445 (N_19445,N_10700,N_14087);
nor U19446 (N_19446,N_11650,N_10500);
nor U19447 (N_19447,N_13641,N_11039);
nor U19448 (N_19448,N_14451,N_10643);
and U19449 (N_19449,N_11343,N_14639);
nor U19450 (N_19450,N_12363,N_14766);
or U19451 (N_19451,N_11573,N_12691);
and U19452 (N_19452,N_12290,N_13693);
nor U19453 (N_19453,N_10039,N_10896);
nand U19454 (N_19454,N_10856,N_13606);
and U19455 (N_19455,N_10464,N_10035);
nand U19456 (N_19456,N_13194,N_11669);
nand U19457 (N_19457,N_13171,N_11168);
xnor U19458 (N_19458,N_14826,N_11065);
or U19459 (N_19459,N_14520,N_14218);
nor U19460 (N_19460,N_11186,N_11531);
nor U19461 (N_19461,N_12437,N_13256);
nand U19462 (N_19462,N_12876,N_10002);
and U19463 (N_19463,N_10426,N_13836);
and U19464 (N_19464,N_12827,N_10509);
nand U19465 (N_19465,N_11000,N_11532);
nor U19466 (N_19466,N_10742,N_12797);
or U19467 (N_19467,N_11803,N_14915);
xor U19468 (N_19468,N_12253,N_11894);
nand U19469 (N_19469,N_10884,N_14333);
nand U19470 (N_19470,N_11928,N_12393);
and U19471 (N_19471,N_11884,N_12071);
nand U19472 (N_19472,N_10658,N_11790);
xnor U19473 (N_19473,N_10839,N_14928);
or U19474 (N_19474,N_11547,N_14491);
xor U19475 (N_19475,N_14761,N_12150);
and U19476 (N_19476,N_10471,N_13206);
nor U19477 (N_19477,N_10056,N_13727);
nand U19478 (N_19478,N_12015,N_14666);
and U19479 (N_19479,N_13977,N_12072);
or U19480 (N_19480,N_13274,N_12691);
or U19481 (N_19481,N_12624,N_10248);
nand U19482 (N_19482,N_11902,N_13629);
xor U19483 (N_19483,N_11220,N_14135);
and U19484 (N_19484,N_10683,N_14478);
nand U19485 (N_19485,N_14554,N_14043);
xor U19486 (N_19486,N_14664,N_13947);
nor U19487 (N_19487,N_13602,N_11854);
xor U19488 (N_19488,N_10711,N_11229);
nand U19489 (N_19489,N_12685,N_11724);
and U19490 (N_19490,N_14416,N_11404);
xnor U19491 (N_19491,N_10576,N_13207);
nand U19492 (N_19492,N_12623,N_13837);
nor U19493 (N_19493,N_10680,N_14244);
nor U19494 (N_19494,N_14579,N_13764);
nand U19495 (N_19495,N_12611,N_11494);
xor U19496 (N_19496,N_12725,N_12608);
or U19497 (N_19497,N_10566,N_13690);
and U19498 (N_19498,N_11387,N_10290);
nor U19499 (N_19499,N_11739,N_11066);
xor U19500 (N_19500,N_12931,N_13697);
and U19501 (N_19501,N_13067,N_12063);
and U19502 (N_19502,N_13245,N_10699);
nand U19503 (N_19503,N_11282,N_11800);
nor U19504 (N_19504,N_10100,N_14362);
nor U19505 (N_19505,N_11175,N_11185);
nand U19506 (N_19506,N_12779,N_14248);
and U19507 (N_19507,N_12883,N_14818);
nor U19508 (N_19508,N_14960,N_12421);
nand U19509 (N_19509,N_11013,N_12610);
xnor U19510 (N_19510,N_10674,N_14088);
and U19511 (N_19511,N_12648,N_11380);
nand U19512 (N_19512,N_11431,N_10156);
nor U19513 (N_19513,N_14698,N_14575);
xor U19514 (N_19514,N_12077,N_13015);
nor U19515 (N_19515,N_11988,N_11385);
or U19516 (N_19516,N_12604,N_13931);
and U19517 (N_19517,N_13595,N_12621);
or U19518 (N_19518,N_10342,N_11054);
nand U19519 (N_19519,N_10718,N_13455);
nor U19520 (N_19520,N_12402,N_14220);
nand U19521 (N_19521,N_10756,N_12357);
nand U19522 (N_19522,N_14285,N_13657);
or U19523 (N_19523,N_10653,N_13605);
and U19524 (N_19524,N_14474,N_10488);
xnor U19525 (N_19525,N_14279,N_11655);
or U19526 (N_19526,N_14953,N_14025);
xor U19527 (N_19527,N_14954,N_12013);
and U19528 (N_19528,N_13763,N_12419);
xor U19529 (N_19529,N_14612,N_11812);
nand U19530 (N_19530,N_14454,N_14456);
xor U19531 (N_19531,N_14540,N_10695);
xnor U19532 (N_19532,N_12286,N_12811);
and U19533 (N_19533,N_14764,N_13026);
and U19534 (N_19534,N_14254,N_11901);
nand U19535 (N_19535,N_10578,N_13882);
xor U19536 (N_19536,N_12159,N_10781);
or U19537 (N_19537,N_10401,N_10399);
nand U19538 (N_19538,N_10051,N_10370);
nand U19539 (N_19539,N_14605,N_12427);
nor U19540 (N_19540,N_11660,N_11761);
xnor U19541 (N_19541,N_14116,N_12662);
nand U19542 (N_19542,N_12832,N_11501);
and U19543 (N_19543,N_14130,N_10255);
nor U19544 (N_19544,N_13709,N_11823);
xnor U19545 (N_19545,N_11391,N_12164);
nor U19546 (N_19546,N_14206,N_14233);
xnor U19547 (N_19547,N_10606,N_14263);
xnor U19548 (N_19548,N_11157,N_12920);
or U19549 (N_19549,N_13323,N_14618);
or U19550 (N_19550,N_12105,N_13723);
nor U19551 (N_19551,N_11340,N_13024);
or U19552 (N_19552,N_10163,N_14741);
nand U19553 (N_19553,N_13336,N_10430);
nand U19554 (N_19554,N_14062,N_13506);
xnor U19555 (N_19555,N_12523,N_12578);
and U19556 (N_19556,N_14879,N_12297);
nor U19557 (N_19557,N_13033,N_14578);
xor U19558 (N_19558,N_13278,N_13291);
or U19559 (N_19559,N_13654,N_13033);
nor U19560 (N_19560,N_10781,N_11949);
nor U19561 (N_19561,N_11433,N_14924);
nor U19562 (N_19562,N_13338,N_11756);
and U19563 (N_19563,N_12716,N_13537);
or U19564 (N_19564,N_11696,N_14386);
nor U19565 (N_19565,N_12405,N_12695);
nand U19566 (N_19566,N_12552,N_14332);
or U19567 (N_19567,N_12575,N_10626);
and U19568 (N_19568,N_14640,N_10066);
or U19569 (N_19569,N_11278,N_14703);
nand U19570 (N_19570,N_11296,N_13973);
xnor U19571 (N_19571,N_14868,N_10372);
or U19572 (N_19572,N_11182,N_14050);
and U19573 (N_19573,N_10318,N_14667);
or U19574 (N_19574,N_12434,N_14528);
xnor U19575 (N_19575,N_14954,N_13178);
and U19576 (N_19576,N_13789,N_12290);
xor U19577 (N_19577,N_10976,N_12020);
nor U19578 (N_19578,N_12390,N_12185);
nand U19579 (N_19579,N_14140,N_14248);
xnor U19580 (N_19580,N_10930,N_14640);
nor U19581 (N_19581,N_11201,N_10043);
xnor U19582 (N_19582,N_13916,N_11520);
or U19583 (N_19583,N_10842,N_12898);
nor U19584 (N_19584,N_10525,N_14028);
nor U19585 (N_19585,N_12656,N_12509);
and U19586 (N_19586,N_10093,N_12042);
xnor U19587 (N_19587,N_11281,N_11471);
and U19588 (N_19588,N_13440,N_10477);
and U19589 (N_19589,N_14030,N_12550);
nor U19590 (N_19590,N_11711,N_10947);
nand U19591 (N_19591,N_14508,N_12949);
or U19592 (N_19592,N_13926,N_14610);
xor U19593 (N_19593,N_14172,N_12550);
nand U19594 (N_19594,N_12821,N_14512);
nand U19595 (N_19595,N_12618,N_13808);
and U19596 (N_19596,N_14667,N_14179);
nor U19597 (N_19597,N_13284,N_12008);
or U19598 (N_19598,N_11774,N_13257);
xnor U19599 (N_19599,N_11990,N_11047);
nand U19600 (N_19600,N_12851,N_11987);
and U19601 (N_19601,N_11009,N_13537);
nor U19602 (N_19602,N_12744,N_13546);
or U19603 (N_19603,N_13920,N_12701);
nor U19604 (N_19604,N_10679,N_13921);
and U19605 (N_19605,N_13251,N_11464);
xor U19606 (N_19606,N_14134,N_10418);
or U19607 (N_19607,N_10584,N_11508);
nand U19608 (N_19608,N_13010,N_10478);
and U19609 (N_19609,N_10501,N_10668);
and U19610 (N_19610,N_10962,N_14731);
or U19611 (N_19611,N_11912,N_13055);
nor U19612 (N_19612,N_14325,N_12329);
and U19613 (N_19613,N_11789,N_10463);
or U19614 (N_19614,N_12465,N_11681);
or U19615 (N_19615,N_11196,N_13645);
nor U19616 (N_19616,N_14826,N_12733);
nor U19617 (N_19617,N_12288,N_10358);
or U19618 (N_19618,N_13443,N_12921);
or U19619 (N_19619,N_10917,N_13703);
and U19620 (N_19620,N_10078,N_13821);
and U19621 (N_19621,N_10242,N_12673);
or U19622 (N_19622,N_12912,N_12299);
nand U19623 (N_19623,N_10545,N_13710);
nand U19624 (N_19624,N_10117,N_11475);
or U19625 (N_19625,N_12399,N_13792);
xnor U19626 (N_19626,N_11750,N_12825);
nor U19627 (N_19627,N_11213,N_14999);
and U19628 (N_19628,N_13761,N_14073);
xnor U19629 (N_19629,N_14036,N_14380);
nor U19630 (N_19630,N_10536,N_10803);
nand U19631 (N_19631,N_11356,N_14003);
nand U19632 (N_19632,N_14825,N_12400);
and U19633 (N_19633,N_10604,N_13148);
xnor U19634 (N_19634,N_14168,N_13264);
and U19635 (N_19635,N_14677,N_13359);
and U19636 (N_19636,N_12644,N_12627);
nor U19637 (N_19637,N_13520,N_11550);
and U19638 (N_19638,N_11924,N_10345);
or U19639 (N_19639,N_10784,N_11229);
nand U19640 (N_19640,N_14011,N_12879);
nand U19641 (N_19641,N_13159,N_11226);
xnor U19642 (N_19642,N_12755,N_11757);
xnor U19643 (N_19643,N_13905,N_14037);
xor U19644 (N_19644,N_10002,N_12631);
xor U19645 (N_19645,N_10566,N_12509);
nand U19646 (N_19646,N_10411,N_10325);
nor U19647 (N_19647,N_12842,N_14270);
xnor U19648 (N_19648,N_12919,N_13006);
nand U19649 (N_19649,N_12281,N_10577);
nand U19650 (N_19650,N_10911,N_13897);
xnor U19651 (N_19651,N_11616,N_14529);
xnor U19652 (N_19652,N_10664,N_11986);
nor U19653 (N_19653,N_12721,N_12326);
xor U19654 (N_19654,N_13568,N_11920);
and U19655 (N_19655,N_14876,N_10867);
or U19656 (N_19656,N_14836,N_11703);
or U19657 (N_19657,N_13192,N_14312);
nor U19658 (N_19658,N_13956,N_10074);
nor U19659 (N_19659,N_13664,N_14329);
and U19660 (N_19660,N_10467,N_12004);
nand U19661 (N_19661,N_10137,N_13887);
or U19662 (N_19662,N_13912,N_12775);
xnor U19663 (N_19663,N_12763,N_14236);
and U19664 (N_19664,N_14473,N_14451);
nor U19665 (N_19665,N_12909,N_13461);
or U19666 (N_19666,N_13169,N_10167);
nand U19667 (N_19667,N_13098,N_14509);
and U19668 (N_19668,N_11535,N_10660);
nor U19669 (N_19669,N_11682,N_11490);
nand U19670 (N_19670,N_12138,N_11543);
xnor U19671 (N_19671,N_12139,N_12687);
or U19672 (N_19672,N_10479,N_10089);
or U19673 (N_19673,N_13675,N_14529);
xor U19674 (N_19674,N_14407,N_13160);
and U19675 (N_19675,N_10503,N_13513);
xor U19676 (N_19676,N_10123,N_13213);
nand U19677 (N_19677,N_13143,N_11625);
and U19678 (N_19678,N_13480,N_12317);
and U19679 (N_19679,N_11200,N_10074);
and U19680 (N_19680,N_13761,N_13746);
nand U19681 (N_19681,N_12920,N_12877);
nor U19682 (N_19682,N_10501,N_11118);
nor U19683 (N_19683,N_14036,N_14732);
xnor U19684 (N_19684,N_13999,N_12079);
nor U19685 (N_19685,N_12133,N_14718);
or U19686 (N_19686,N_13482,N_12410);
nand U19687 (N_19687,N_12694,N_10984);
xor U19688 (N_19688,N_13303,N_12002);
or U19689 (N_19689,N_10368,N_12842);
nor U19690 (N_19690,N_11957,N_12714);
or U19691 (N_19691,N_14004,N_11860);
nand U19692 (N_19692,N_14537,N_10688);
nand U19693 (N_19693,N_13779,N_13632);
nor U19694 (N_19694,N_10353,N_12689);
or U19695 (N_19695,N_13692,N_14639);
or U19696 (N_19696,N_11499,N_10079);
or U19697 (N_19697,N_10040,N_10570);
and U19698 (N_19698,N_10957,N_10614);
or U19699 (N_19699,N_13953,N_12002);
and U19700 (N_19700,N_13032,N_13869);
nor U19701 (N_19701,N_14950,N_11142);
xor U19702 (N_19702,N_11799,N_11384);
or U19703 (N_19703,N_10793,N_13744);
nand U19704 (N_19704,N_12463,N_13095);
xor U19705 (N_19705,N_13950,N_12774);
xor U19706 (N_19706,N_14126,N_13022);
nor U19707 (N_19707,N_13781,N_10614);
nand U19708 (N_19708,N_13909,N_11377);
and U19709 (N_19709,N_13637,N_13203);
and U19710 (N_19710,N_13648,N_10564);
and U19711 (N_19711,N_12773,N_12126);
nor U19712 (N_19712,N_14304,N_10880);
xnor U19713 (N_19713,N_11154,N_12595);
or U19714 (N_19714,N_14442,N_14769);
nand U19715 (N_19715,N_13008,N_10824);
xnor U19716 (N_19716,N_13837,N_14918);
nor U19717 (N_19717,N_13647,N_13778);
nand U19718 (N_19718,N_12872,N_14123);
and U19719 (N_19719,N_12894,N_12426);
nor U19720 (N_19720,N_12471,N_13280);
nor U19721 (N_19721,N_10661,N_12100);
or U19722 (N_19722,N_11425,N_13966);
xnor U19723 (N_19723,N_13201,N_11185);
xnor U19724 (N_19724,N_13272,N_13405);
nand U19725 (N_19725,N_14662,N_13953);
nand U19726 (N_19726,N_13993,N_14356);
nand U19727 (N_19727,N_13506,N_10168);
nor U19728 (N_19728,N_12750,N_11137);
or U19729 (N_19729,N_13158,N_13480);
or U19730 (N_19730,N_14667,N_13568);
nor U19731 (N_19731,N_13493,N_11462);
and U19732 (N_19732,N_11707,N_10496);
nor U19733 (N_19733,N_11491,N_10760);
and U19734 (N_19734,N_12152,N_11090);
xor U19735 (N_19735,N_12805,N_11763);
nand U19736 (N_19736,N_13195,N_11214);
or U19737 (N_19737,N_11128,N_13849);
and U19738 (N_19738,N_10883,N_10499);
xnor U19739 (N_19739,N_11448,N_13015);
and U19740 (N_19740,N_10138,N_11048);
nand U19741 (N_19741,N_12214,N_13780);
nand U19742 (N_19742,N_13270,N_13423);
nand U19743 (N_19743,N_11291,N_14011);
or U19744 (N_19744,N_11267,N_14150);
xnor U19745 (N_19745,N_10928,N_12090);
nor U19746 (N_19746,N_11500,N_11623);
and U19747 (N_19747,N_12526,N_10743);
xor U19748 (N_19748,N_13099,N_11783);
or U19749 (N_19749,N_10310,N_12650);
xor U19750 (N_19750,N_14080,N_14704);
and U19751 (N_19751,N_11557,N_13447);
nand U19752 (N_19752,N_14274,N_11426);
nor U19753 (N_19753,N_13327,N_11012);
nand U19754 (N_19754,N_12071,N_10143);
and U19755 (N_19755,N_14171,N_12894);
xnor U19756 (N_19756,N_10449,N_13748);
nand U19757 (N_19757,N_11958,N_12777);
nor U19758 (N_19758,N_14415,N_11880);
or U19759 (N_19759,N_14409,N_14542);
nand U19760 (N_19760,N_12526,N_14234);
nor U19761 (N_19761,N_14271,N_13638);
xor U19762 (N_19762,N_10488,N_10007);
nor U19763 (N_19763,N_13207,N_13871);
nor U19764 (N_19764,N_10445,N_13609);
xnor U19765 (N_19765,N_13459,N_10463);
nand U19766 (N_19766,N_11036,N_12953);
nor U19767 (N_19767,N_10739,N_10346);
nand U19768 (N_19768,N_13022,N_11628);
and U19769 (N_19769,N_12131,N_13713);
or U19770 (N_19770,N_10101,N_11067);
or U19771 (N_19771,N_11523,N_11170);
or U19772 (N_19772,N_12508,N_10532);
xnor U19773 (N_19773,N_10527,N_13981);
or U19774 (N_19774,N_10897,N_10117);
or U19775 (N_19775,N_13353,N_10002);
nor U19776 (N_19776,N_12391,N_12420);
and U19777 (N_19777,N_12872,N_10454);
nor U19778 (N_19778,N_14730,N_10391);
and U19779 (N_19779,N_13357,N_10865);
nand U19780 (N_19780,N_12921,N_14528);
nor U19781 (N_19781,N_10944,N_10835);
or U19782 (N_19782,N_10296,N_11210);
xor U19783 (N_19783,N_10612,N_12036);
and U19784 (N_19784,N_13991,N_12828);
nand U19785 (N_19785,N_11578,N_13870);
nand U19786 (N_19786,N_14211,N_12783);
or U19787 (N_19787,N_14053,N_10901);
xnor U19788 (N_19788,N_14793,N_10180);
xor U19789 (N_19789,N_11302,N_12428);
nand U19790 (N_19790,N_10041,N_11689);
nand U19791 (N_19791,N_14055,N_10626);
or U19792 (N_19792,N_13419,N_12250);
and U19793 (N_19793,N_12090,N_11476);
xnor U19794 (N_19794,N_13059,N_11400);
or U19795 (N_19795,N_13466,N_13975);
xnor U19796 (N_19796,N_14158,N_10446);
xnor U19797 (N_19797,N_11728,N_10106);
and U19798 (N_19798,N_10962,N_13040);
nand U19799 (N_19799,N_12903,N_10228);
nor U19800 (N_19800,N_10343,N_11064);
xnor U19801 (N_19801,N_11735,N_13239);
and U19802 (N_19802,N_10232,N_14235);
nand U19803 (N_19803,N_10538,N_10592);
xnor U19804 (N_19804,N_10405,N_10134);
and U19805 (N_19805,N_11394,N_11008);
nor U19806 (N_19806,N_13755,N_14591);
or U19807 (N_19807,N_13065,N_12397);
xnor U19808 (N_19808,N_13952,N_12516);
xor U19809 (N_19809,N_12707,N_12778);
and U19810 (N_19810,N_14751,N_11168);
and U19811 (N_19811,N_13689,N_13918);
xor U19812 (N_19812,N_10737,N_12045);
nand U19813 (N_19813,N_10656,N_14166);
nand U19814 (N_19814,N_10434,N_11392);
or U19815 (N_19815,N_11078,N_14448);
or U19816 (N_19816,N_14428,N_11631);
nor U19817 (N_19817,N_12438,N_12244);
nand U19818 (N_19818,N_13756,N_13467);
or U19819 (N_19819,N_14926,N_11450);
xor U19820 (N_19820,N_12028,N_14929);
nand U19821 (N_19821,N_13814,N_10966);
or U19822 (N_19822,N_11776,N_10929);
nand U19823 (N_19823,N_14512,N_12116);
or U19824 (N_19824,N_12867,N_10116);
xnor U19825 (N_19825,N_13188,N_12098);
and U19826 (N_19826,N_12026,N_11992);
nand U19827 (N_19827,N_14571,N_13737);
xnor U19828 (N_19828,N_13590,N_12134);
or U19829 (N_19829,N_12643,N_13348);
or U19830 (N_19830,N_14942,N_11455);
or U19831 (N_19831,N_13575,N_14567);
xor U19832 (N_19832,N_10807,N_11023);
nor U19833 (N_19833,N_11799,N_10822);
nand U19834 (N_19834,N_10264,N_12117);
and U19835 (N_19835,N_10201,N_11515);
or U19836 (N_19836,N_12832,N_13444);
xnor U19837 (N_19837,N_12278,N_11671);
xor U19838 (N_19838,N_11960,N_13951);
nor U19839 (N_19839,N_10420,N_11474);
xor U19840 (N_19840,N_14292,N_14561);
or U19841 (N_19841,N_10875,N_10796);
xor U19842 (N_19842,N_13182,N_14921);
and U19843 (N_19843,N_10102,N_12030);
or U19844 (N_19844,N_11280,N_13775);
xor U19845 (N_19845,N_10625,N_14800);
xnor U19846 (N_19846,N_13507,N_12923);
nor U19847 (N_19847,N_13945,N_11136);
nand U19848 (N_19848,N_13970,N_12206);
xor U19849 (N_19849,N_14503,N_11500);
and U19850 (N_19850,N_13602,N_12559);
or U19851 (N_19851,N_13581,N_11268);
and U19852 (N_19852,N_12804,N_11647);
and U19853 (N_19853,N_10247,N_10623);
xnor U19854 (N_19854,N_11939,N_12073);
nand U19855 (N_19855,N_11493,N_11645);
and U19856 (N_19856,N_12813,N_11673);
and U19857 (N_19857,N_12301,N_10151);
nor U19858 (N_19858,N_13276,N_10277);
or U19859 (N_19859,N_12243,N_10314);
xor U19860 (N_19860,N_14698,N_12039);
nor U19861 (N_19861,N_12170,N_11589);
xnor U19862 (N_19862,N_13421,N_10348);
and U19863 (N_19863,N_10386,N_10390);
nor U19864 (N_19864,N_10314,N_14446);
and U19865 (N_19865,N_12883,N_10286);
xnor U19866 (N_19866,N_13211,N_13824);
xor U19867 (N_19867,N_11434,N_11507);
or U19868 (N_19868,N_14606,N_12015);
or U19869 (N_19869,N_10112,N_13281);
xnor U19870 (N_19870,N_11613,N_14609);
and U19871 (N_19871,N_13968,N_12912);
nand U19872 (N_19872,N_10709,N_14113);
or U19873 (N_19873,N_13169,N_11994);
and U19874 (N_19874,N_14063,N_11121);
xnor U19875 (N_19875,N_12581,N_12755);
nor U19876 (N_19876,N_13370,N_14310);
nor U19877 (N_19877,N_14300,N_11865);
nor U19878 (N_19878,N_12154,N_14702);
and U19879 (N_19879,N_14412,N_13292);
or U19880 (N_19880,N_12403,N_10985);
xor U19881 (N_19881,N_14660,N_12218);
and U19882 (N_19882,N_12420,N_13366);
nor U19883 (N_19883,N_14358,N_14469);
or U19884 (N_19884,N_11642,N_11430);
nand U19885 (N_19885,N_12825,N_12680);
xor U19886 (N_19886,N_13571,N_13202);
and U19887 (N_19887,N_14660,N_12746);
nand U19888 (N_19888,N_14821,N_11620);
or U19889 (N_19889,N_13895,N_13120);
xnor U19890 (N_19890,N_14285,N_14926);
nor U19891 (N_19891,N_12053,N_11535);
xor U19892 (N_19892,N_10389,N_11722);
and U19893 (N_19893,N_14961,N_13260);
or U19894 (N_19894,N_13869,N_10479);
xnor U19895 (N_19895,N_13379,N_10926);
xnor U19896 (N_19896,N_11037,N_12545);
xor U19897 (N_19897,N_12940,N_12610);
and U19898 (N_19898,N_13325,N_11159);
and U19899 (N_19899,N_11018,N_10189);
nand U19900 (N_19900,N_14658,N_11782);
and U19901 (N_19901,N_11444,N_10423);
nand U19902 (N_19902,N_13437,N_10156);
xnor U19903 (N_19903,N_10648,N_12380);
xnor U19904 (N_19904,N_14309,N_12504);
xnor U19905 (N_19905,N_11378,N_13262);
nand U19906 (N_19906,N_12880,N_11109);
and U19907 (N_19907,N_11025,N_12815);
nand U19908 (N_19908,N_10369,N_13843);
nand U19909 (N_19909,N_14165,N_10190);
nand U19910 (N_19910,N_12172,N_11738);
nand U19911 (N_19911,N_14625,N_11886);
nand U19912 (N_19912,N_13797,N_13297);
nor U19913 (N_19913,N_14503,N_10688);
nand U19914 (N_19914,N_13165,N_14958);
and U19915 (N_19915,N_11503,N_10805);
and U19916 (N_19916,N_13418,N_14329);
and U19917 (N_19917,N_14739,N_12467);
or U19918 (N_19918,N_12382,N_12340);
nor U19919 (N_19919,N_11054,N_11457);
or U19920 (N_19920,N_11316,N_13641);
or U19921 (N_19921,N_11117,N_11685);
xor U19922 (N_19922,N_14278,N_11997);
xnor U19923 (N_19923,N_12540,N_14209);
nor U19924 (N_19924,N_10049,N_11608);
nand U19925 (N_19925,N_12339,N_10536);
xor U19926 (N_19926,N_13875,N_12535);
nand U19927 (N_19927,N_14187,N_10216);
and U19928 (N_19928,N_13739,N_12920);
xor U19929 (N_19929,N_14451,N_13338);
nor U19930 (N_19930,N_13307,N_13526);
nor U19931 (N_19931,N_14551,N_14880);
and U19932 (N_19932,N_10280,N_11124);
or U19933 (N_19933,N_14528,N_10232);
nand U19934 (N_19934,N_14001,N_14974);
and U19935 (N_19935,N_12992,N_13135);
nor U19936 (N_19936,N_14807,N_11162);
or U19937 (N_19937,N_10381,N_14325);
xor U19938 (N_19938,N_14932,N_12733);
xnor U19939 (N_19939,N_14842,N_11954);
xnor U19940 (N_19940,N_13641,N_11756);
or U19941 (N_19941,N_11564,N_12885);
nand U19942 (N_19942,N_14085,N_10161);
and U19943 (N_19943,N_14269,N_10554);
nand U19944 (N_19944,N_11943,N_11703);
and U19945 (N_19945,N_12129,N_13249);
xnor U19946 (N_19946,N_14629,N_10290);
nor U19947 (N_19947,N_10143,N_13784);
nor U19948 (N_19948,N_10935,N_13993);
nand U19949 (N_19949,N_11437,N_10407);
nor U19950 (N_19950,N_12897,N_12798);
and U19951 (N_19951,N_13238,N_11820);
and U19952 (N_19952,N_13454,N_12034);
and U19953 (N_19953,N_14354,N_10504);
xor U19954 (N_19954,N_13684,N_13466);
or U19955 (N_19955,N_14041,N_14573);
nor U19956 (N_19956,N_13320,N_14593);
nor U19957 (N_19957,N_11300,N_13354);
and U19958 (N_19958,N_10987,N_11493);
nand U19959 (N_19959,N_14945,N_14853);
nor U19960 (N_19960,N_11074,N_14561);
nor U19961 (N_19961,N_10015,N_10698);
and U19962 (N_19962,N_10976,N_10247);
xor U19963 (N_19963,N_13714,N_10986);
or U19964 (N_19964,N_12355,N_12628);
and U19965 (N_19965,N_11610,N_12868);
xnor U19966 (N_19966,N_14948,N_13358);
or U19967 (N_19967,N_14869,N_12277);
and U19968 (N_19968,N_14085,N_14112);
nor U19969 (N_19969,N_13213,N_14729);
and U19970 (N_19970,N_11485,N_11554);
nand U19971 (N_19971,N_12275,N_12535);
xnor U19972 (N_19972,N_14516,N_12464);
or U19973 (N_19973,N_11691,N_14443);
or U19974 (N_19974,N_12119,N_10706);
nor U19975 (N_19975,N_10949,N_13976);
nand U19976 (N_19976,N_11638,N_14316);
nor U19977 (N_19977,N_12252,N_10883);
xor U19978 (N_19978,N_13429,N_13391);
and U19979 (N_19979,N_14437,N_12240);
or U19980 (N_19980,N_14114,N_14557);
or U19981 (N_19981,N_13568,N_13583);
nor U19982 (N_19982,N_11312,N_12582);
nand U19983 (N_19983,N_10477,N_10069);
nand U19984 (N_19984,N_12998,N_12654);
or U19985 (N_19985,N_13342,N_10332);
xor U19986 (N_19986,N_11766,N_13892);
and U19987 (N_19987,N_14325,N_13671);
xor U19988 (N_19988,N_11135,N_12240);
nor U19989 (N_19989,N_14303,N_11809);
and U19990 (N_19990,N_11538,N_12617);
nand U19991 (N_19991,N_12023,N_12723);
or U19992 (N_19992,N_14757,N_10699);
and U19993 (N_19993,N_14392,N_12127);
nor U19994 (N_19994,N_14371,N_10415);
nand U19995 (N_19995,N_12249,N_13489);
nand U19996 (N_19996,N_10607,N_13110);
nor U19997 (N_19997,N_12415,N_13436);
and U19998 (N_19998,N_11167,N_13174);
nand U19999 (N_19999,N_11993,N_14622);
or U20000 (N_20000,N_17321,N_15938);
and U20001 (N_20001,N_17541,N_16773);
or U20002 (N_20002,N_16224,N_15598);
or U20003 (N_20003,N_16971,N_15243);
or U20004 (N_20004,N_16799,N_17776);
or U20005 (N_20005,N_15226,N_15138);
and U20006 (N_20006,N_16766,N_16784);
nor U20007 (N_20007,N_19057,N_16745);
and U20008 (N_20008,N_16843,N_17311);
or U20009 (N_20009,N_18957,N_15410);
nor U20010 (N_20010,N_18910,N_18864);
xnor U20011 (N_20011,N_17026,N_19652);
xor U20012 (N_20012,N_15480,N_19931);
and U20013 (N_20013,N_15246,N_15450);
xor U20014 (N_20014,N_19139,N_18550);
or U20015 (N_20015,N_15016,N_15776);
nor U20016 (N_20016,N_15645,N_17338);
nor U20017 (N_20017,N_18646,N_15924);
and U20018 (N_20018,N_17930,N_18213);
or U20019 (N_20019,N_18435,N_15417);
xnor U20020 (N_20020,N_18282,N_15808);
xnor U20021 (N_20021,N_17487,N_17494);
nand U20022 (N_20022,N_15041,N_17211);
nand U20023 (N_20023,N_16925,N_15754);
and U20024 (N_20024,N_17962,N_17373);
nand U20025 (N_20025,N_17119,N_18670);
nor U20026 (N_20026,N_17611,N_17187);
nor U20027 (N_20027,N_15809,N_16802);
or U20028 (N_20028,N_18665,N_16083);
nand U20029 (N_20029,N_15520,N_19250);
nand U20030 (N_20030,N_17282,N_19428);
or U20031 (N_20031,N_16000,N_18112);
and U20032 (N_20032,N_18300,N_18445);
xnor U20033 (N_20033,N_15845,N_16994);
nand U20034 (N_20034,N_15735,N_15556);
or U20035 (N_20035,N_18531,N_16797);
nand U20036 (N_20036,N_18537,N_18442);
xnor U20037 (N_20037,N_16553,N_19806);
xor U20038 (N_20038,N_17569,N_17938);
and U20039 (N_20039,N_19510,N_18524);
and U20040 (N_20040,N_19655,N_16777);
and U20041 (N_20041,N_19046,N_15106);
or U20042 (N_20042,N_17379,N_15501);
or U20043 (N_20043,N_15842,N_17217);
or U20044 (N_20044,N_15033,N_16442);
nor U20045 (N_20045,N_16614,N_16241);
xor U20046 (N_20046,N_18610,N_19337);
nor U20047 (N_20047,N_19997,N_18629);
and U20048 (N_20048,N_16259,N_18750);
nand U20049 (N_20049,N_16926,N_19108);
xnor U20050 (N_20050,N_18838,N_15320);
nor U20051 (N_20051,N_16611,N_17572);
and U20052 (N_20052,N_17824,N_16390);
and U20053 (N_20053,N_19918,N_15839);
nand U20054 (N_20054,N_17326,N_18323);
nand U20055 (N_20055,N_19040,N_15683);
nor U20056 (N_20056,N_19444,N_19827);
xor U20057 (N_20057,N_19523,N_17994);
xnor U20058 (N_20058,N_19842,N_17452);
nand U20059 (N_20059,N_18911,N_16322);
or U20060 (N_20060,N_16425,N_16514);
nand U20061 (N_20061,N_19726,N_19230);
xnor U20062 (N_20062,N_15470,N_15336);
or U20063 (N_20063,N_18438,N_16552);
nand U20064 (N_20064,N_15230,N_18362);
or U20065 (N_20065,N_19625,N_17017);
or U20066 (N_20066,N_18286,N_17958);
nand U20067 (N_20067,N_19802,N_18225);
nand U20068 (N_20068,N_19304,N_16513);
nor U20069 (N_20069,N_15346,N_17702);
and U20070 (N_20070,N_15303,N_15180);
or U20071 (N_20071,N_15663,N_17421);
xnor U20072 (N_20072,N_18974,N_16833);
and U20073 (N_20073,N_15657,N_18803);
xor U20074 (N_20074,N_18771,N_18485);
nand U20075 (N_20075,N_18473,N_16407);
and U20076 (N_20076,N_16470,N_17432);
nor U20077 (N_20077,N_18860,N_15562);
nor U20078 (N_20078,N_18804,N_16010);
or U20079 (N_20079,N_18971,N_18726);
xnor U20080 (N_20080,N_17065,N_16751);
and U20081 (N_20081,N_16380,N_18760);
nor U20082 (N_20082,N_15884,N_17850);
xor U20083 (N_20083,N_19665,N_16385);
or U20084 (N_20084,N_17859,N_17021);
nand U20085 (N_20085,N_18951,N_15950);
or U20086 (N_20086,N_18317,N_15765);
nand U20087 (N_20087,N_17622,N_19168);
and U20088 (N_20088,N_16518,N_17526);
nor U20089 (N_20089,N_17503,N_19551);
and U20090 (N_20090,N_16836,N_15418);
nor U20091 (N_20091,N_18586,N_15555);
or U20092 (N_20092,N_15524,N_17351);
xnor U20093 (N_20093,N_18105,N_15902);
nor U20094 (N_20094,N_18378,N_17558);
and U20095 (N_20095,N_17359,N_16040);
and U20096 (N_20096,N_16557,N_16324);
and U20097 (N_20097,N_16675,N_15255);
xnor U20098 (N_20098,N_19882,N_16495);
nand U20099 (N_20099,N_18812,N_16504);
nor U20100 (N_20100,N_19533,N_15658);
nor U20101 (N_20101,N_16570,N_16317);
or U20102 (N_20102,N_17641,N_17290);
xor U20103 (N_20103,N_15932,N_19700);
xor U20104 (N_20104,N_19450,N_17616);
nor U20105 (N_20105,N_15630,N_15193);
xnor U20106 (N_20106,N_15881,N_19702);
nor U20107 (N_20107,N_16431,N_15828);
nor U20108 (N_20108,N_19147,N_18275);
or U20109 (N_20109,N_19078,N_19674);
and U20110 (N_20110,N_19870,N_17695);
xor U20111 (N_20111,N_16668,N_16353);
or U20112 (N_20112,N_15232,N_15566);
nand U20113 (N_20113,N_17058,N_19492);
xnor U20114 (N_20114,N_17443,N_19958);
nand U20115 (N_20115,N_16868,N_18732);
and U20116 (N_20116,N_19171,N_17714);
nor U20117 (N_20117,N_15622,N_18051);
and U20118 (N_20118,N_18019,N_17208);
xnor U20119 (N_20119,N_18143,N_16526);
nand U20120 (N_20120,N_17078,N_17816);
nor U20121 (N_20121,N_18628,N_16318);
xor U20122 (N_20122,N_19272,N_16869);
nand U20123 (N_20123,N_19769,N_16543);
xor U20124 (N_20124,N_15904,N_18977);
xor U20125 (N_20125,N_15305,N_15538);
nand U20126 (N_20126,N_19195,N_15741);
or U20127 (N_20127,N_16837,N_19379);
and U20128 (N_20128,N_17803,N_15901);
nor U20129 (N_20129,N_17857,N_17814);
nor U20130 (N_20130,N_17957,N_19395);
and U20131 (N_20131,N_17583,N_15025);
nor U20132 (N_20132,N_19602,N_18966);
xor U20133 (N_20133,N_18155,N_15406);
nor U20134 (N_20134,N_17689,N_17981);
nand U20135 (N_20135,N_18158,N_17447);
or U20136 (N_20136,N_15964,N_16962);
and U20137 (N_20137,N_18131,N_18061);
or U20138 (N_20138,N_17176,N_17895);
nand U20139 (N_20139,N_16633,N_18431);
nand U20140 (N_20140,N_17554,N_18727);
or U20141 (N_20141,N_15582,N_19595);
nand U20142 (N_20142,N_19154,N_19728);
and U20143 (N_20143,N_17810,N_18274);
xnor U20144 (N_20144,N_16612,N_16654);
nand U20145 (N_20145,N_15945,N_19857);
or U20146 (N_20146,N_15494,N_18941);
nand U20147 (N_20147,N_15662,N_19204);
or U20148 (N_20148,N_18847,N_18160);
and U20149 (N_20149,N_19408,N_15888);
or U20150 (N_20150,N_19292,N_18697);
xor U20151 (N_20151,N_17739,N_18677);
nand U20152 (N_20152,N_19926,N_17354);
and U20153 (N_20153,N_19540,N_18689);
xor U20154 (N_20154,N_17672,N_18873);
and U20155 (N_20155,N_17372,N_18126);
xnor U20156 (N_20156,N_19268,N_16575);
or U20157 (N_20157,N_19412,N_19748);
nand U20158 (N_20158,N_17592,N_15458);
nor U20159 (N_20159,N_15504,N_17086);
xnor U20160 (N_20160,N_17428,N_18942);
nand U20161 (N_20161,N_18059,N_19328);
nand U20162 (N_20162,N_17153,N_15135);
or U20163 (N_20163,N_16674,N_19105);
xnor U20164 (N_20164,N_18690,N_16043);
or U20165 (N_20165,N_16337,N_17157);
and U20166 (N_20166,N_16061,N_19356);
nor U20167 (N_20167,N_19805,N_19936);
or U20168 (N_20168,N_15838,N_17301);
or U20169 (N_20169,N_17697,N_19442);
nand U20170 (N_20170,N_18273,N_17075);
xnor U20171 (N_20171,N_17542,N_18602);
nor U20172 (N_20172,N_16138,N_19487);
xnor U20173 (N_20173,N_16860,N_15609);
nor U20174 (N_20174,N_15646,N_16024);
nor U20175 (N_20175,N_16983,N_15527);
nand U20176 (N_20176,N_18630,N_19079);
nor U20177 (N_20177,N_18523,N_19651);
xnor U20178 (N_20178,N_15251,N_17943);
or U20179 (N_20179,N_16591,N_17174);
nand U20180 (N_20180,N_18107,N_17263);
or U20181 (N_20181,N_18736,N_16260);
or U20182 (N_20182,N_16814,N_19446);
and U20183 (N_20183,N_19576,N_17927);
and U20184 (N_20184,N_17564,N_18662);
xnor U20185 (N_20185,N_16817,N_18195);
nor U20186 (N_20186,N_18111,N_15007);
xor U20187 (N_20187,N_18448,N_18405);
and U20188 (N_20188,N_16527,N_16792);
and U20189 (N_20189,N_17070,N_16579);
nor U20190 (N_20190,N_19513,N_17717);
xnor U20191 (N_20191,N_17360,N_19603);
nand U20192 (N_20192,N_15624,N_17020);
or U20193 (N_20193,N_18678,N_17870);
or U20194 (N_20194,N_18540,N_15618);
and U20195 (N_20195,N_16039,N_19839);
nor U20196 (N_20196,N_19344,N_18142);
or U20197 (N_20197,N_17254,N_17745);
nor U20198 (N_20198,N_19445,N_16300);
xnor U20199 (N_20199,N_18876,N_18130);
nand U20200 (N_20200,N_18253,N_16546);
nor U20201 (N_20201,N_17552,N_16199);
or U20202 (N_20202,N_16944,N_17606);
or U20203 (N_20203,N_16295,N_16999);
or U20204 (N_20204,N_16253,N_18350);
nand U20205 (N_20205,N_16605,N_15155);
or U20206 (N_20206,N_15413,N_17560);
xor U20207 (N_20207,N_18589,N_19366);
or U20208 (N_20208,N_18426,N_19759);
and U20209 (N_20209,N_15090,N_19508);
xnor U20210 (N_20210,N_15580,N_16947);
xor U20211 (N_20211,N_17120,N_15824);
or U20212 (N_20212,N_19766,N_17499);
or U20213 (N_20213,N_18809,N_15969);
or U20214 (N_20214,N_18014,N_17374);
nor U20215 (N_20215,N_17094,N_19989);
and U20216 (N_20216,N_16942,N_15100);
nand U20217 (N_20217,N_18724,N_19512);
xor U20218 (N_20218,N_15392,N_18177);
nand U20219 (N_20219,N_15471,N_18333);
and U20220 (N_20220,N_17821,N_17220);
nand U20221 (N_20221,N_18845,N_15134);
nor U20222 (N_20222,N_19479,N_17921);
nand U20223 (N_20223,N_19588,N_18912);
and U20224 (N_20224,N_16396,N_18731);
xnor U20225 (N_20225,N_18784,N_15581);
nor U20226 (N_20226,N_17313,N_18147);
xor U20227 (N_20227,N_16428,N_17645);
and U20228 (N_20228,N_15039,N_15165);
xor U20229 (N_20229,N_16443,N_18985);
or U20230 (N_20230,N_15862,N_16759);
nor U20231 (N_20231,N_17956,N_18358);
nor U20232 (N_20232,N_16195,N_16309);
and U20233 (N_20233,N_15182,N_17950);
nand U20234 (N_20234,N_19447,N_18250);
nand U20235 (N_20235,N_18679,N_15941);
nand U20236 (N_20236,N_16819,N_15907);
xnor U20237 (N_20237,N_16343,N_15981);
nand U20238 (N_20238,N_19488,N_17789);
and U20239 (N_20239,N_17225,N_15249);
and U20240 (N_20240,N_16519,N_19433);
or U20241 (N_20241,N_19593,N_18478);
xor U20242 (N_20242,N_19648,N_15145);
xnor U20243 (N_20243,N_15936,N_18163);
nor U20244 (N_20244,N_19768,N_17330);
nor U20245 (N_20245,N_18790,N_19003);
xor U20246 (N_20246,N_19247,N_15472);
or U20247 (N_20247,N_18616,N_18507);
or U20248 (N_20248,N_15891,N_19861);
or U20249 (N_20249,N_15724,N_15518);
nand U20250 (N_20250,N_19521,N_16899);
xnor U20251 (N_20251,N_19742,N_15184);
or U20252 (N_20252,N_18782,N_15316);
nand U20253 (N_20253,N_15889,N_15114);
nand U20254 (N_20254,N_17044,N_15642);
nand U20255 (N_20255,N_16714,N_18964);
and U20256 (N_20256,N_16898,N_19158);
xor U20257 (N_20257,N_15063,N_15067);
and U20258 (N_20258,N_15009,N_19414);
and U20259 (N_20259,N_15438,N_19025);
xnor U20260 (N_20260,N_17424,N_16538);
or U20261 (N_20261,N_19244,N_18748);
nand U20262 (N_20262,N_19093,N_16275);
or U20263 (N_20263,N_17341,N_17703);
or U20264 (N_20264,N_17557,N_15910);
nor U20265 (N_20265,N_17736,N_17806);
or U20266 (N_20266,N_15113,N_18872);
nand U20267 (N_20267,N_19402,N_15311);
nand U20268 (N_20268,N_17018,N_16459);
xnor U20269 (N_20269,N_16491,N_19866);
xor U20270 (N_20270,N_15287,N_19090);
or U20271 (N_20271,N_16051,N_17011);
xnor U20272 (N_20272,N_17377,N_18357);
or U20273 (N_20273,N_19852,N_16372);
and U20274 (N_20274,N_17970,N_18826);
xor U20275 (N_20275,N_17565,N_16940);
and U20276 (N_20276,N_16113,N_19453);
and U20277 (N_20277,N_15024,N_16620);
nor U20278 (N_20278,N_18497,N_17287);
and U20279 (N_20279,N_16438,N_18835);
or U20280 (N_20280,N_19682,N_19348);
or U20281 (N_20281,N_19313,N_19260);
nor U20282 (N_20282,N_18406,N_15811);
nand U20283 (N_20283,N_17388,N_18279);
nand U20284 (N_20284,N_18729,N_19591);
or U20285 (N_20285,N_15906,N_16291);
or U20286 (N_20286,N_16888,N_19118);
and U20287 (N_20287,N_17183,N_15607);
xor U20288 (N_20288,N_16640,N_15116);
xnor U20289 (N_20289,N_16827,N_17216);
and U20290 (N_20290,N_16567,N_15894);
and U20291 (N_20291,N_19325,N_15871);
nor U20292 (N_20292,N_17188,N_18353);
nand U20293 (N_20293,N_16831,N_17288);
xnor U20294 (N_20294,N_15172,N_16371);
and U20295 (N_20295,N_18156,N_17318);
nand U20296 (N_20296,N_19618,N_16585);
xnor U20297 (N_20297,N_17876,N_18247);
and U20298 (N_20298,N_16783,N_19854);
nor U20299 (N_20299,N_18395,N_18007);
and U20300 (N_20300,N_15405,N_18683);
xor U20301 (N_20301,N_18355,N_16651);
and U20302 (N_20302,N_18164,N_18151);
xnor U20303 (N_20303,N_17741,N_15254);
or U20304 (N_20304,N_15940,N_16376);
nand U20305 (N_20305,N_19928,N_16851);
or U20306 (N_20306,N_16440,N_17845);
xor U20307 (N_20307,N_16743,N_18753);
or U20308 (N_20308,N_15727,N_17793);
nor U20309 (N_20309,N_15748,N_16093);
xnor U20310 (N_20310,N_18898,N_16964);
nand U20311 (N_20311,N_17800,N_15592);
xnor U20312 (N_20312,N_19876,N_16064);
or U20313 (N_20313,N_16314,N_15057);
or U20314 (N_20314,N_18859,N_17154);
xor U20315 (N_20315,N_16812,N_17029);
or U20316 (N_20316,N_17783,N_18146);
or U20317 (N_20317,N_18376,N_16753);
and U20318 (N_20318,N_19557,N_19007);
or U20319 (N_20319,N_16424,N_17718);
and U20320 (N_20320,N_15633,N_19788);
nand U20321 (N_20321,N_19564,N_18197);
nand U20322 (N_20322,N_17853,N_16466);
xor U20323 (N_20323,N_19619,N_19199);
and U20324 (N_20324,N_17408,N_17271);
xor U20325 (N_20325,N_19699,N_15740);
xor U20326 (N_20326,N_16624,N_19142);
and U20327 (N_20327,N_19384,N_15170);
xnor U20328 (N_20328,N_18559,N_19144);
or U20329 (N_20329,N_16847,N_17969);
nor U20330 (N_20330,N_16340,N_18351);
or U20331 (N_20331,N_18422,N_15706);
and U20332 (N_20332,N_17340,N_19478);
nand U20333 (N_20333,N_18590,N_17207);
nor U20334 (N_20334,N_17948,N_19358);
nor U20335 (N_20335,N_15363,N_16297);
and U20336 (N_20336,N_15680,N_19713);
nand U20337 (N_20337,N_17458,N_16180);
xnor U20338 (N_20338,N_18747,N_15261);
nor U20339 (N_20339,N_17680,N_17767);
xnor U20340 (N_20340,N_19024,N_16845);
nor U20341 (N_20341,N_18597,N_17100);
xor U20342 (N_20342,N_18349,N_18897);
xor U20343 (N_20343,N_16800,N_16811);
or U20344 (N_20344,N_15503,N_16455);
or U20345 (N_20345,N_16678,N_19306);
xnor U20346 (N_20346,N_16499,N_18308);
xor U20347 (N_20347,N_16046,N_18464);
and U20348 (N_20348,N_18424,N_15088);
nor U20349 (N_20349,N_15976,N_19373);
nor U20350 (N_20350,N_15541,N_18973);
or U20351 (N_20351,N_17272,N_18893);
and U20352 (N_20352,N_15034,N_17448);
nand U20353 (N_20353,N_17418,N_16356);
nand U20354 (N_20354,N_16658,N_17517);
nor U20355 (N_20355,N_15183,N_18065);
or U20356 (N_20356,N_15621,N_17589);
nand U20357 (N_20357,N_18285,N_16479);
nand U20358 (N_20358,N_16184,N_18902);
xnor U20359 (N_20359,N_19182,N_19097);
and U20360 (N_20360,N_15844,N_19930);
and U20361 (N_20361,N_18906,N_15078);
and U20362 (N_20362,N_15578,N_17177);
and U20363 (N_20363,N_17603,N_19933);
and U20364 (N_20364,N_17593,N_19874);
or U20365 (N_20365,N_19562,N_16059);
nor U20366 (N_20366,N_16032,N_18054);
xor U20367 (N_20367,N_18104,N_16871);
nand U20368 (N_20368,N_16437,N_18767);
nand U20369 (N_20369,N_18137,N_17903);
or U20370 (N_20370,N_18298,N_18699);
nand U20371 (N_20371,N_18023,N_19639);
xor U20372 (N_20372,N_17145,N_15128);
nand U20373 (N_20373,N_19273,N_18294);
xor U20374 (N_20374,N_15373,N_19830);
nor U20375 (N_20375,N_18220,N_17337);
and U20376 (N_20376,N_17769,N_18189);
xor U20377 (N_20377,N_16629,N_15465);
nand U20378 (N_20378,N_15006,N_19466);
nand U20379 (N_20379,N_17815,N_15552);
nand U20380 (N_20380,N_15998,N_16842);
and U20381 (N_20381,N_16510,N_15949);
nand U20382 (N_20382,N_15107,N_15523);
xor U20383 (N_20383,N_15084,N_17255);
or U20384 (N_20384,N_18572,N_15505);
and U20385 (N_20385,N_19311,N_16417);
xor U20386 (N_20386,N_15228,N_17515);
nor U20387 (N_20387,N_15175,N_19341);
and U20388 (N_20388,N_16578,N_15753);
xnor U20389 (N_20389,N_16637,N_18141);
nor U20390 (N_20390,N_19772,N_16363);
nor U20391 (N_20391,N_16511,N_19708);
nor U20392 (N_20392,N_19420,N_18654);
nand U20393 (N_20393,N_19081,N_18352);
or U20394 (N_20394,N_17038,N_15730);
or U20395 (N_20395,N_16281,N_18943);
or U20396 (N_20396,N_19823,N_15721);
xor U20397 (N_20397,N_19431,N_16149);
and U20398 (N_20398,N_16112,N_15801);
and U20399 (N_20399,N_15595,N_16219);
nand U20400 (N_20400,N_17596,N_19732);
and U20401 (N_20401,N_19240,N_18981);
nor U20402 (N_20402,N_15927,N_18034);
or U20403 (N_20403,N_17066,N_16215);
or U20404 (N_20404,N_18495,N_16090);
and U20405 (N_20405,N_19630,N_16946);
nand U20406 (N_20406,N_19608,N_18739);
and U20407 (N_20407,N_18006,N_15046);
nand U20408 (N_20408,N_17752,N_15771);
xnor U20409 (N_20409,N_16191,N_16844);
and U20410 (N_20410,N_18134,N_17121);
nand U20411 (N_20411,N_15979,N_18466);
or U20412 (N_20412,N_17059,N_19644);
nor U20413 (N_20413,N_18712,N_15269);
nor U20414 (N_20414,N_19267,N_19976);
nand U20415 (N_20415,N_18233,N_18591);
and U20416 (N_20416,N_15897,N_18304);
nand U20417 (N_20417,N_18136,N_16397);
nand U20418 (N_20418,N_15247,N_19006);
and U20419 (N_20419,N_18312,N_17818);
and U20420 (N_20420,N_19038,N_17861);
nand U20421 (N_20421,N_15271,N_19360);
nand U20422 (N_20422,N_16932,N_19215);
and U20423 (N_20423,N_18758,N_18154);
xor U20424 (N_20424,N_19491,N_17601);
and U20425 (N_20425,N_19060,N_19867);
or U20426 (N_20426,N_19065,N_16156);
nand U20427 (N_20427,N_18802,N_16862);
or U20428 (N_20428,N_15029,N_19841);
xnor U20429 (N_20429,N_17090,N_16694);
or U20430 (N_20430,N_17362,N_16211);
nand U20431 (N_20431,N_17292,N_16120);
nand U20432 (N_20432,N_15540,N_19174);
or U20433 (N_20433,N_18208,N_19821);
and U20434 (N_20434,N_17844,N_17966);
or U20435 (N_20435,N_18599,N_18619);
xor U20436 (N_20436,N_15611,N_15717);
or U20437 (N_20437,N_15939,N_16865);
nand U20438 (N_20438,N_15507,N_19050);
nand U20439 (N_20439,N_16494,N_15484);
xnor U20440 (N_20440,N_19758,N_18343);
and U20441 (N_20441,N_16734,N_17582);
and U20442 (N_20442,N_15491,N_16342);
xor U20443 (N_20443,N_15276,N_17817);
xor U20444 (N_20444,N_15054,N_19096);
nor U20445 (N_20445,N_17397,N_19460);
and U20446 (N_20446,N_16664,N_17658);
and U20447 (N_20447,N_15676,N_15648);
nor U20448 (N_20448,N_15797,N_15869);
nand U20449 (N_20449,N_19689,N_17249);
xor U20450 (N_20450,N_16170,N_16029);
or U20451 (N_20451,N_16361,N_19763);
and U20452 (N_20452,N_19181,N_16174);
or U20453 (N_20453,N_16469,N_17170);
and U20454 (N_20454,N_18926,N_16715);
xor U20455 (N_20455,N_17655,N_16911);
and U20456 (N_20456,N_19221,N_18510);
nor U20457 (N_20457,N_15195,N_17636);
or U20458 (N_20458,N_16153,N_18133);
and U20459 (N_20459,N_19297,N_17089);
nor U20460 (N_20460,N_17553,N_16049);
or U20461 (N_20461,N_19801,N_15692);
and U20462 (N_20462,N_16548,N_17419);
xnor U20463 (N_20463,N_19069,N_16235);
nand U20464 (N_20464,N_15997,N_16303);
xor U20465 (N_20465,N_18168,N_17864);
or U20466 (N_20466,N_17671,N_19354);
nor U20467 (N_20467,N_18535,N_16960);
nor U20468 (N_20468,N_15212,N_17777);
nand U20469 (N_20469,N_17704,N_16636);
and U20470 (N_20470,N_19988,N_16134);
xor U20471 (N_20471,N_15273,N_18330);
and U20472 (N_20472,N_17708,N_15908);
and U20473 (N_20473,N_16422,N_19761);
nand U20474 (N_20474,N_17124,N_16105);
nor U20475 (N_20475,N_17771,N_18152);
xor U20476 (N_20476,N_17949,N_18016);
nor U20477 (N_20477,N_15710,N_17561);
nor U20478 (N_20478,N_16735,N_19095);
nor U20479 (N_20479,N_18120,N_17298);
and U20480 (N_20480,N_15565,N_17014);
xor U20481 (N_20481,N_17236,N_16700);
nand U20482 (N_20482,N_16824,N_17305);
and U20483 (N_20483,N_17315,N_15101);
nor U20484 (N_20484,N_19776,N_16638);
and U20485 (N_20485,N_16193,N_19587);
nor U20486 (N_20486,N_18010,N_15412);
nand U20487 (N_20487,N_17841,N_15358);
and U20488 (N_20488,N_19511,N_19155);
xnor U20489 (N_20489,N_19100,N_18819);
nand U20490 (N_20490,N_16254,N_15857);
or U20491 (N_20491,N_16897,N_15151);
or U20492 (N_20492,N_17878,N_17939);
nor U20493 (N_20493,N_18471,N_19434);
nand U20494 (N_20494,N_17076,N_15506);
and U20495 (N_20495,N_19499,N_17607);
nor U20496 (N_20496,N_16849,N_18937);
and U20497 (N_20497,N_19580,N_19035);
xnor U20498 (N_20498,N_16805,N_18128);
or U20499 (N_20499,N_19248,N_15384);
nand U20500 (N_20500,N_18640,N_18504);
or U20501 (N_20501,N_16308,N_17184);
nor U20502 (N_20502,N_16265,N_15495);
nor U20503 (N_20503,N_17118,N_18655);
xnor U20504 (N_20504,N_15434,N_18992);
or U20505 (N_20505,N_16534,N_19560);
and U20506 (N_20506,N_18255,N_18011);
xor U20507 (N_20507,N_19869,N_15489);
nor U20508 (N_20508,N_17523,N_19799);
or U20509 (N_20509,N_15688,N_17820);
and U20510 (N_20510,N_17158,N_17041);
nor U20511 (N_20511,N_19883,N_15926);
xor U20512 (N_20512,N_18083,N_19681);
xor U20513 (N_20513,N_15414,N_16206);
nand U20514 (N_20514,N_19949,N_19711);
nor U20515 (N_20515,N_15350,N_16606);
or U20516 (N_20516,N_17716,N_16568);
nand U20517 (N_20517,N_19904,N_17025);
nor U20518 (N_20518,N_19623,N_17862);
or U20519 (N_20519,N_19952,N_16222);
nand U20520 (N_20520,N_19858,N_19780);
and U20521 (N_20521,N_15085,N_18737);
xor U20522 (N_20522,N_15288,N_19686);
or U20523 (N_20523,N_17347,N_15360);
or U20524 (N_20524,N_17128,N_15509);
nor U20525 (N_20525,N_17135,N_16079);
xor U20526 (N_20526,N_18908,N_18374);
and U20527 (N_20527,N_17987,N_19284);
or U20528 (N_20528,N_19190,N_17050);
or U20529 (N_20529,N_19881,N_16592);
or U20530 (N_20530,N_19575,N_17737);
nand U20531 (N_20531,N_19518,N_19355);
nand U20532 (N_20532,N_19073,N_17281);
or U20533 (N_20533,N_16137,N_17846);
and U20534 (N_20534,N_16978,N_19146);
and U20535 (N_20535,N_18667,N_16116);
nor U20536 (N_20536,N_17387,N_15812);
or U20537 (N_20537,N_19405,N_16172);
nor U20538 (N_20538,N_19500,N_18576);
nand U20539 (N_20539,N_19394,N_18676);
or U20540 (N_20540,N_16118,N_17417);
and U20541 (N_20541,N_17087,N_15780);
xnor U20542 (N_20542,N_18024,N_18595);
xnor U20543 (N_20543,N_19307,N_19981);
or U20544 (N_20544,N_19489,N_15517);
or U20545 (N_20545,N_15326,N_19493);
xnor U20546 (N_20546,N_17733,N_16873);
or U20547 (N_20547,N_16902,N_19561);
nand U20548 (N_20548,N_16956,N_18302);
or U20549 (N_20549,N_18125,N_18423);
or U20550 (N_20550,N_15313,N_15312);
or U20551 (N_20551,N_18307,N_15751);
xor U20552 (N_20552,N_16389,N_18046);
nand U20553 (N_20553,N_18621,N_18776);
nor U20554 (N_20554,N_16976,N_18852);
nor U20555 (N_20555,N_18494,N_17951);
and U20556 (N_20556,N_15455,N_15833);
and U20557 (N_20557,N_17389,N_18492);
xnor U20558 (N_20558,N_19277,N_17791);
and U20559 (N_20559,N_18093,N_15354);
xnor U20560 (N_20560,N_18730,N_19167);
or U20561 (N_20561,N_19934,N_17280);
or U20562 (N_20562,N_18070,N_18169);
and U20563 (N_20563,N_16123,N_19335);
and U20564 (N_20564,N_18099,N_15615);
nand U20565 (N_20565,N_16159,N_18567);
or U20566 (N_20566,N_16834,N_17760);
or U20567 (N_20567,N_16826,N_16891);
and U20568 (N_20568,N_15792,N_17375);
nor U20569 (N_20569,N_16233,N_18420);
nand U20570 (N_20570,N_18324,N_19701);
nor U20571 (N_20571,N_16311,N_15514);
or U20572 (N_20572,N_15338,N_19051);
xor U20573 (N_20573,N_17574,N_16178);
or U20574 (N_20574,N_17509,N_19129);
or U20575 (N_20575,N_19265,N_17865);
xor U20576 (N_20576,N_16068,N_18372);
nor U20577 (N_20577,N_19400,N_19254);
or U20578 (N_20578,N_19913,N_17530);
nor U20579 (N_20579,N_16875,N_16903);
xor U20580 (N_20580,N_18386,N_16141);
xnor U20581 (N_20581,N_18606,N_18291);
nand U20582 (N_20582,N_16670,N_15716);
nor U20583 (N_20583,N_15055,N_18361);
nand U20584 (N_20584,N_18587,N_17977);
nand U20585 (N_20585,N_17773,N_19924);
xor U20586 (N_20586,N_16108,N_17711);
or U20587 (N_20587,N_17239,N_15922);
nor U20588 (N_20588,N_18309,N_15905);
xnor U20589 (N_20589,N_16053,N_15018);
xnor U20590 (N_20590,N_17807,N_17355);
or U20591 (N_20591,N_15817,N_15988);
xnor U20592 (N_20592,N_18254,N_19538);
or U20593 (N_20593,N_18664,N_17562);
nand U20594 (N_20594,N_18098,N_18622);
nor U20595 (N_20595,N_19889,N_18717);
nand U20596 (N_20596,N_15482,N_15488);
or U20597 (N_20597,N_15867,N_16704);
and U20598 (N_20598,N_17051,N_17631);
nor U20599 (N_20599,N_18284,N_16017);
and U20600 (N_20600,N_17908,N_16450);
nand U20601 (N_20601,N_15239,N_16742);
nor U20602 (N_20602,N_16489,N_18222);
nand U20603 (N_20603,N_17045,N_17492);
nand U20604 (N_20604,N_16011,N_15733);
nor U20605 (N_20605,N_15934,N_18397);
and U20606 (N_20606,N_18659,N_15265);
nand U20607 (N_20607,N_19653,N_18903);
nor U20608 (N_20608,N_18101,N_17489);
nand U20609 (N_20609,N_15962,N_16661);
or U20610 (N_20610,N_19448,N_16341);
or U20611 (N_20611,N_17317,N_15222);
nor U20612 (N_20612,N_15725,N_16791);
and U20613 (N_20613,N_15546,N_17712);
or U20614 (N_20614,N_17449,N_17663);
nand U20615 (N_20615,N_17300,N_16951);
nand U20616 (N_20616,N_17393,N_15701);
and U20617 (N_20617,N_16673,N_19863);
and U20618 (N_20618,N_15032,N_18738);
nor U20619 (N_20619,N_18658,N_15215);
and U20620 (N_20620,N_17136,N_17436);
nand U20621 (N_20621,N_18639,N_17008);
nor U20622 (N_20622,N_18235,N_17229);
and U20623 (N_20623,N_16449,N_17178);
nand U20624 (N_20624,N_17221,N_19894);
xor U20625 (N_20625,N_18704,N_17193);
nand U20626 (N_20626,N_17247,N_15399);
or U20627 (N_20627,N_18695,N_16892);
nor U20628 (N_20628,N_15293,N_18412);
xor U20629 (N_20629,N_17304,N_15712);
and U20630 (N_20630,N_15573,N_15383);
nand U20631 (N_20631,N_15071,N_15755);
xnor U20632 (N_20632,N_16196,N_19103);
nand U20633 (N_20633,N_19015,N_15421);
xnor U20634 (N_20634,N_19932,N_16201);
xor U20635 (N_20635,N_15446,N_18117);
and U20636 (N_20636,N_16048,N_19495);
xnor U20637 (N_20637,N_17911,N_16569);
or U20638 (N_20638,N_18751,N_15848);
or U20639 (N_20639,N_16119,N_18828);
or U20640 (N_20640,N_15367,N_16488);
and U20641 (N_20641,N_15525,N_17469);
xor U20642 (N_20642,N_19266,N_17117);
or U20643 (N_20643,N_18446,N_16436);
nand U20644 (N_20644,N_16705,N_15918);
xor U20645 (N_20645,N_15917,N_18956);
xnor U20646 (N_20646,N_16597,N_19600);
or U20647 (N_20647,N_15365,N_17754);
nand U20648 (N_20648,N_18020,N_15890);
nand U20649 (N_20649,N_15377,N_18398);
nor U20650 (N_20650,N_15987,N_17284);
and U20651 (N_20651,N_19520,N_15638);
xnor U20652 (N_20652,N_19049,N_16106);
and U20653 (N_20653,N_18339,N_16104);
or U20654 (N_20654,N_18295,N_15789);
nand U20655 (N_20655,N_19197,N_18493);
or U20656 (N_20656,N_18187,N_16840);
nor U20657 (N_20657,N_15798,N_18761);
and U20658 (N_20658,N_19259,N_18715);
xnor U20659 (N_20659,N_19000,N_19391);
nor U20660 (N_20660,N_15353,N_15073);
xnor U20661 (N_20661,N_19465,N_15931);
nand U20662 (N_20662,N_17204,N_18498);
xnor U20663 (N_20663,N_19421,N_15513);
xor U20664 (N_20664,N_18673,N_16486);
nor U20665 (N_20665,N_19547,N_17520);
xor U20666 (N_20666,N_19528,N_15060);
nor U20667 (N_20667,N_16313,N_16035);
nand U20668 (N_20668,N_15895,N_19346);
or U20669 (N_20669,N_17085,N_16262);
and U20670 (N_20670,N_17770,N_15723);
xor U20671 (N_20671,N_18925,N_17222);
or U20672 (N_20672,N_17446,N_15374);
nand U20673 (N_20673,N_19396,N_15548);
and U20674 (N_20674,N_17866,N_17457);
xnor U20675 (N_20675,N_18028,N_17617);
or U20676 (N_20676,N_18914,N_19813);
xor U20677 (N_20677,N_19722,N_17279);
or U20678 (N_20678,N_18705,N_19352);
and U20679 (N_20679,N_18569,N_16057);
nor U20680 (N_20680,N_16335,N_15442);
nand U20681 (N_20681,N_19786,N_19962);
xnor U20682 (N_20682,N_18733,N_16961);
nor U20683 (N_20683,N_15056,N_19359);
nor U20684 (N_20684,N_19995,N_18186);
nor U20685 (N_20685,N_18528,N_16695);
and U20686 (N_20686,N_18728,N_18890);
nor U20687 (N_20687,N_18548,N_15477);
nor U20688 (N_20688,N_15225,N_15661);
xnor U20689 (N_20689,N_19846,N_17999);
xor U20690 (N_20690,N_18100,N_16456);
and U20691 (N_20691,N_17167,N_18815);
nor U20692 (N_20692,N_18316,N_15855);
and U20693 (N_20693,N_19201,N_15767);
or U20694 (N_20694,N_19628,N_16870);
xor U20695 (N_20695,N_15913,N_15129);
and U20696 (N_20696,N_18886,N_19973);
nand U20697 (N_20697,N_19956,N_16273);
and U20698 (N_20698,N_16240,N_17597);
or U20699 (N_20699,N_16452,N_18297);
xor U20700 (N_20700,N_19900,N_16740);
nor U20701 (N_20701,N_15210,N_16589);
or U20702 (N_20702,N_15686,N_16416);
nand U20703 (N_20703,N_16545,N_19919);
and U20704 (N_20704,N_19378,N_17975);
nor U20705 (N_20705,N_15985,N_18399);
or U20706 (N_20706,N_18268,N_19896);
or U20707 (N_20707,N_19730,N_18626);
xor U20708 (N_20708,N_16493,N_17723);
xnor U20709 (N_20709,N_16292,N_16854);
nand U20710 (N_20710,N_18834,N_18527);
and U20711 (N_20711,N_16647,N_17438);
xnor U20712 (N_20712,N_18461,N_16249);
xnor U20713 (N_20713,N_18318,N_15560);
or U20714 (N_20714,N_16521,N_17782);
and U20715 (N_20715,N_19814,N_15900);
nand U20716 (N_20716,N_15834,N_18063);
nand U20717 (N_20717,N_15164,N_19832);
nand U20718 (N_20718,N_18391,N_16365);
xor U20719 (N_20719,N_16823,N_15389);
nand U20720 (N_20720,N_15847,N_15632);
nor U20721 (N_20721,N_15764,N_17366);
nor U20722 (N_20722,N_18696,N_17926);
and U20723 (N_20723,N_18450,N_15327);
or U20724 (N_20724,N_16642,N_15703);
xnor U20725 (N_20725,N_15836,N_15015);
nand U20726 (N_20726,N_17581,N_15372);
nand U20727 (N_20727,N_17302,N_16312);
nand U20728 (N_20728,N_18127,N_15850);
nand U20729 (N_20729,N_16143,N_18509);
nor U20730 (N_20730,N_15066,N_16217);
nand U20731 (N_20731,N_19320,N_17599);
nor U20732 (N_20732,N_17151,N_18322);
nand U20733 (N_20733,N_16081,N_18262);
xor U20734 (N_20734,N_19192,N_17022);
and U20735 (N_20735,N_17463,N_15270);
and U20736 (N_20736,N_15022,N_18700);
and U20737 (N_20737,N_18867,N_18411);
nand U20738 (N_20738,N_15961,N_16930);
nand U20739 (N_20739,N_17023,N_17972);
nand U20740 (N_20740,N_17619,N_16481);
nand U20741 (N_20741,N_15675,N_18161);
and U20742 (N_20742,N_19298,N_18680);
or U20743 (N_20743,N_19635,N_17394);
and U20744 (N_20744,N_18427,N_18797);
and U20745 (N_20745,N_19020,N_18641);
xnor U20746 (N_20746,N_18581,N_19300);
xor U20747 (N_20747,N_16445,N_18832);
nand U20748 (N_20748,N_19974,N_19198);
nand U20749 (N_20749,N_15761,N_16070);
or U20750 (N_20750,N_17486,N_19967);
and U20751 (N_20751,N_17798,N_18336);
xor U20752 (N_20752,N_18150,N_19583);
nor U20753 (N_20753,N_19517,N_19589);
nand U20754 (N_20754,N_19892,N_19068);
nand U20755 (N_20755,N_15213,N_15822);
nand U20756 (N_20756,N_15954,N_15569);
and U20757 (N_20757,N_17412,N_19023);
or U20758 (N_20758,N_15019,N_17490);
and U20759 (N_20759,N_19675,N_15424);
xor U20760 (N_20760,N_16770,N_17369);
or U20761 (N_20761,N_19977,N_16182);
xor U20762 (N_20762,N_15672,N_17161);
nand U20763 (N_20763,N_18012,N_17299);
nor U20764 (N_20764,N_17209,N_19878);
nor U20765 (N_20765,N_19897,N_19774);
nor U20766 (N_20766,N_19535,N_17953);
and U20767 (N_20767,N_17095,N_18190);
or U20768 (N_20768,N_16852,N_17838);
nand U20769 (N_20769,N_19855,N_16974);
nand U20770 (N_20770,N_18384,N_19274);
or U20771 (N_20771,N_19778,N_19698);
or U20772 (N_20772,N_16274,N_17738);
and U20773 (N_20773,N_16429,N_15331);
nand U20774 (N_20774,N_16853,N_19544);
or U20775 (N_20775,N_19275,N_16776);
or U20776 (N_20776,N_16878,N_15736);
or U20777 (N_20777,N_15694,N_19848);
nor U20778 (N_20778,N_17102,N_19409);
or U20779 (N_20779,N_17048,N_18175);
nand U20780 (N_20780,N_17350,N_16148);
nand U20781 (N_20781,N_17612,N_17743);
and U20782 (N_20782,N_16657,N_17348);
xor U20783 (N_20783,N_18800,N_18013);
nand U20784 (N_20784,N_15181,N_16763);
xor U20785 (N_20785,N_15787,N_16848);
xnor U20786 (N_20786,N_18919,N_16458);
and U20787 (N_20787,N_16204,N_15371);
xor U20788 (N_20788,N_18521,N_19503);
and U20789 (N_20789,N_15013,N_17875);
xnor U20790 (N_20790,N_19236,N_15325);
or U20791 (N_20791,N_15898,N_15841);
nand U20792 (N_20792,N_15854,N_16405);
xnor U20793 (N_20793,N_18511,N_15588);
nand U20794 (N_20794,N_18417,N_15294);
nand U20795 (N_20795,N_15148,N_15709);
nor U20796 (N_20796,N_15023,N_16485);
and U20797 (N_20797,N_17831,N_19596);
xnor U20798 (N_20798,N_17874,N_17465);
xor U20799 (N_20799,N_15426,N_18212);
xor U20800 (N_20800,N_18415,N_15923);
or U20801 (N_20801,N_16316,N_16351);
and U20802 (N_20802,N_17328,N_15253);
xnor U20803 (N_20803,N_18138,N_16781);
nand U20804 (N_20804,N_15310,N_19494);
or U20805 (N_20805,N_19411,N_15681);
xor U20806 (N_20806,N_17830,N_18091);
xnor U20807 (N_20807,N_19754,N_17453);
xnor U20808 (N_20808,N_15511,N_18375);
xnor U20809 (N_20809,N_18240,N_15763);
nor U20810 (N_20810,N_17495,N_18661);
xnor U20811 (N_20811,N_16711,N_15104);
nor U20812 (N_20812,N_19571,N_16427);
or U20813 (N_20813,N_17191,N_16650);
and U20814 (N_20814,N_18299,N_19439);
or U20815 (N_20815,N_18720,N_18447);
xor U20816 (N_20816,N_17905,N_16772);
nand U20817 (N_20817,N_17719,N_17171);
and U20818 (N_20818,N_16278,N_17740);
or U20819 (N_20819,N_17308,N_16272);
nand U20820 (N_20820,N_19101,N_18843);
and U20821 (N_20821,N_18062,N_15757);
xnor U20822 (N_20822,N_16364,N_16025);
nor U20823 (N_20823,N_17502,N_18039);
and U20824 (N_20824,N_18040,N_15396);
xor U20825 (N_20825,N_19012,N_18594);
nand U20826 (N_20826,N_18421,N_16085);
or U20827 (N_20827,N_16434,N_18770);
nand U20828 (N_20828,N_16229,N_16754);
or U20829 (N_20829,N_19663,N_16329);
xnor U20830 (N_20830,N_18122,N_17992);
nand U20831 (N_20831,N_18552,N_18965);
xnor U20832 (N_20832,N_15086,N_19251);
nor U20833 (N_20833,N_15357,N_15047);
xor U20834 (N_20834,N_19803,N_18644);
nand U20835 (N_20835,N_19137,N_18778);
xnor U20836 (N_20836,N_15427,N_16478);
and U20837 (N_20837,N_15671,N_19704);
nand U20838 (N_20838,N_18652,N_16198);
xnor U20839 (N_20839,N_19902,N_15231);
xor U20840 (N_20840,N_18088,N_16603);
and U20841 (N_20841,N_17654,N_18064);
and U20842 (N_20842,N_19921,N_16395);
nand U20843 (N_20843,N_16816,N_19526);
and U20844 (N_20844,N_16242,N_15816);
xnor U20845 (N_20845,N_19187,N_19660);
nor U20846 (N_20846,N_18648,N_15286);
nand U20847 (N_20847,N_15037,N_18097);
nand U20848 (N_20848,N_18841,N_15925);
or U20849 (N_20849,N_16981,N_19607);
or U20850 (N_20850,N_16841,N_17415);
nand U20851 (N_20851,N_16933,N_16212);
nor U20852 (N_20852,N_17033,N_17710);
xnor U20853 (N_20853,N_16767,N_18057);
nor U20854 (N_20854,N_19134,N_16267);
or U20855 (N_20855,N_15719,N_16687);
and U20856 (N_20856,N_19843,N_17555);
or U20857 (N_20857,N_17456,N_19258);
xor U20858 (N_20858,N_18075,N_18469);
and U20859 (N_20859,N_15456,N_17923);
xnor U20860 (N_20860,N_16359,N_15572);
nor U20861 (N_20861,N_16803,N_15447);
nor U20862 (N_20862,N_18242,N_15877);
or U20863 (N_20863,N_17244,N_19374);
nor U20864 (N_20864,N_18181,N_19039);
and U20865 (N_20865,N_19656,N_15644);
xor U20866 (N_20866,N_17586,N_15304);
and U20867 (N_20867,N_19614,N_15637);
nor U20868 (N_20868,N_19161,N_19545);
nor U20869 (N_20869,N_19558,N_16307);
or U20870 (N_20870,N_16175,N_16980);
xor U20871 (N_20871,N_17314,N_15448);
nor U20872 (N_20872,N_16346,N_17976);
nand U20873 (N_20873,N_16924,N_16015);
nor U20874 (N_20874,N_16163,N_17722);
xnor U20875 (N_20875,N_15915,N_19309);
nor U20876 (N_20876,N_16378,N_19611);
and U20877 (N_20877,N_17238,N_18258);
or U20878 (N_20878,N_16423,N_16598);
nor U20879 (N_20879,N_15219,N_18549);
nor U20880 (N_20880,N_15593,N_15419);
nor U20881 (N_20881,N_18604,N_15781);
nand U20882 (N_20882,N_17079,N_18025);
xnor U20883 (N_20883,N_16628,N_18001);
nand U20884 (N_20884,N_17967,N_19610);
and U20885 (N_20885,N_19898,N_16621);
nand U20886 (N_20886,N_16028,N_18385);
nor U20887 (N_20887,N_18887,N_16001);
nor U20888 (N_20888,N_17613,N_16320);
nor U20889 (N_20889,N_18979,N_16863);
nor U20890 (N_20890,N_19048,N_19567);
xnor U20891 (N_20891,N_16867,N_18930);
nand U20892 (N_20892,N_15403,N_18917);
nand U20893 (N_20893,N_19249,N_15005);
and U20894 (N_20894,N_19971,N_19332);
and U20895 (N_20895,N_19176,N_19188);
and U20896 (N_20896,N_15805,N_18967);
nand U20897 (N_20897,N_18433,N_17906);
nand U20898 (N_20898,N_16531,N_17243);
or U20899 (N_20899,N_17667,N_17194);
and U20900 (N_20900,N_16995,N_19271);
nor U20901 (N_20901,N_19148,N_17405);
and U20902 (N_20902,N_16076,N_15130);
and U20903 (N_20903,N_15045,N_16468);
or U20904 (N_20904,N_15027,N_16626);
or U20905 (N_20905,N_18871,N_16214);
or U20906 (N_20906,N_17852,N_16909);
or U20907 (N_20907,N_19152,N_15110);
and U20908 (N_20908,N_19207,N_17651);
nor U20909 (N_20909,N_15266,N_19357);
and U20910 (N_20910,N_18716,N_16707);
nor U20911 (N_20911,N_15970,N_16333);
nand U20912 (N_20912,N_15339,N_16525);
and U20913 (N_20913,N_15285,N_16912);
and U20914 (N_20914,N_17150,N_15221);
nand U20915 (N_20915,N_17529,N_15189);
nor U20916 (N_20916,N_19685,N_16533);
xnor U20917 (N_20917,N_18363,N_15278);
and U20918 (N_20918,N_17524,N_19490);
xnor U20919 (N_20919,N_18585,N_19741);
xor U20920 (N_20920,N_15217,N_19157);
xnor U20921 (N_20921,N_19935,N_19404);
nor U20922 (N_20922,N_17879,N_15631);
nand U20923 (N_20923,N_17323,N_16828);
xnor U20924 (N_20924,N_16896,N_15870);
or U20925 (N_20925,N_15142,N_19586);
and U20926 (N_20926,N_16052,N_19668);
nand U20927 (N_20927,N_19584,N_16952);
nand U20928 (N_20928,N_15702,N_15698);
xnor U20929 (N_20929,N_16590,N_18884);
nor U20930 (N_20930,N_15440,N_15444);
xnor U20931 (N_20931,N_19552,N_17122);
nand U20932 (N_20932,N_18132,N_18681);
and U20933 (N_20933,N_16250,N_19407);
nor U20934 (N_20934,N_18123,N_17310);
nor U20935 (N_20935,N_16248,N_18947);
nor U20936 (N_20936,N_19756,N_17539);
or U20937 (N_20937,N_17694,N_16126);
nand U20938 (N_20938,N_16073,N_16439);
nand U20939 (N_20939,N_15238,N_16165);
xor U20940 (N_20940,N_19927,N_15307);
nor U20941 (N_20941,N_18991,N_17568);
nor U20942 (N_20942,N_17823,N_16031);
nand U20943 (N_20943,N_17790,N_18409);
or U20944 (N_20944,N_16114,N_18830);
nor U20945 (N_20945,N_15705,N_15342);
or U20946 (N_20946,N_19716,N_19498);
nor U20947 (N_20947,N_18080,N_16693);
xnor U20948 (N_20948,N_19186,N_18891);
and U20949 (N_20949,N_16535,N_18455);
and U20950 (N_20950,N_17445,N_15971);
nand U20951 (N_20951,N_18870,N_18183);
and U20952 (N_20952,N_15144,N_16771);
nand U20953 (N_20953,N_15508,N_18766);
or U20954 (N_20954,N_19353,N_16710);
nor U20955 (N_20955,N_19573,N_18503);
nand U20956 (N_20956,N_18880,N_18044);
and U20957 (N_20957,N_19291,N_18310);
nor U20958 (N_20958,N_19269,N_18082);
nor U20959 (N_20959,N_17935,N_15937);
xnor U20960 (N_20960,N_17423,N_17664);
nand U20961 (N_20961,N_17669,N_17877);
and U20962 (N_20962,N_19323,N_17578);
or U20963 (N_20963,N_15308,N_19102);
nand U20964 (N_20964,N_18714,N_18955);
and U20965 (N_20965,N_19940,N_19113);
and U20966 (N_20966,N_16327,N_18008);
nand U20967 (N_20967,N_18631,N_17527);
or U20968 (N_20968,N_18816,N_16375);
xor U20969 (N_20969,N_16302,N_17914);
xor U20970 (N_20970,N_15300,N_19246);
nand U20971 (N_20971,N_18798,N_19418);
xnor U20972 (N_20972,N_16484,N_15975);
nand U20973 (N_20973,N_17162,N_16331);
xnor U20974 (N_20974,N_15000,N_19302);
or U20975 (N_20975,N_15933,N_19262);
nor U20976 (N_20976,N_17891,N_18568);
and U20977 (N_20977,N_18875,N_15492);
or U20978 (N_20978,N_18451,N_18829);
xor U20979 (N_20979,N_18671,N_17056);
xnor U20980 (N_20980,N_16874,N_18114);
xor U20981 (N_20981,N_19860,N_15443);
or U20982 (N_20982,N_15146,N_15628);
nand U20983 (N_20983,N_15745,N_18219);
nor U20984 (N_20984,N_19413,N_19462);
nor U20985 (N_20985,N_18325,N_17226);
nand U20986 (N_20986,N_15963,N_16122);
nor U20987 (N_20987,N_15813,N_17624);
nor U20988 (N_20988,N_19243,N_15912);
and U20989 (N_20989,N_19053,N_17788);
nor U20990 (N_20990,N_15245,N_18223);
nand U20991 (N_20991,N_19324,N_19170);
nor U20992 (N_20992,N_18530,N_15827);
and U20993 (N_20993,N_16360,N_16464);
nand U20994 (N_20994,N_18159,N_16200);
and U20995 (N_20995,N_17873,N_18272);
or U20996 (N_20996,N_17980,N_19632);
xnor U20997 (N_20997,N_19750,N_18236);
nor U20998 (N_20998,N_15177,N_15214);
nand U20999 (N_20999,N_16132,N_18702);
xnor U21000 (N_21000,N_17887,N_19617);
nand U21001 (N_21001,N_18777,N_18774);
or U21002 (N_21002,N_17705,N_17364);
and U21003 (N_21003,N_19957,N_17630);
and U21004 (N_21004,N_19795,N_19109);
nand U21005 (N_21005,N_18781,N_18532);
nor U21006 (N_21006,N_16793,N_17643);
or U21007 (N_21007,N_17251,N_19539);
and U21008 (N_21008,N_19121,N_17507);
and U21009 (N_21009,N_19083,N_18687);
xor U21010 (N_21010,N_18031,N_18584);
nand U21011 (N_21011,N_17109,N_19938);
or U21012 (N_21012,N_19415,N_19270);
xnor U21013 (N_21013,N_17871,N_16339);
xnor U21014 (N_21014,N_19293,N_15814);
and U21015 (N_21015,N_17978,N_16953);
nand U21016 (N_21016,N_16859,N_18201);
nor U21017 (N_21017,N_17536,N_15485);
and U21018 (N_21018,N_18095,N_19764);
xnor U21019 (N_21019,N_18056,N_19885);
or U21020 (N_21020,N_15314,N_18499);
and U21021 (N_21021,N_15697,N_19042);
and U21022 (N_21022,N_15916,N_17796);
xnor U21023 (N_21023,N_19027,N_19242);
nand U21024 (N_21024,N_19076,N_17729);
nand U21025 (N_21025,N_19914,N_19141);
and U21026 (N_21026,N_18940,N_16023);
and U21027 (N_21027,N_19471,N_18005);
nor U21028 (N_21028,N_18090,N_19047);
xnor U21029 (N_21029,N_17197,N_16410);
or U21030 (N_21030,N_18844,N_15268);
xor U21031 (N_21031,N_18986,N_15864);
or U21032 (N_21032,N_15617,N_17296);
nor U21033 (N_21033,N_16987,N_15668);
nor U21034 (N_21034,N_19753,N_17768);
nand U21035 (N_21035,N_17482,N_19676);
xnor U21036 (N_21036,N_17464,N_17180);
and U21037 (N_21037,N_15823,N_16906);
and U21038 (N_21038,N_15275,N_17735);
nor U21039 (N_21039,N_19524,N_17276);
and U21040 (N_21040,N_15785,N_15829);
nand U21041 (N_21041,N_17441,N_15227);
and U21042 (N_21042,N_15337,N_19757);
or U21043 (N_21043,N_18883,N_19112);
and U21044 (N_21044,N_15206,N_16723);
xor U21045 (N_21045,N_17513,N_17913);
and U21046 (N_21046,N_17210,N_17073);
or U21047 (N_21047,N_18079,N_18837);
or U21048 (N_21048,N_18293,N_19707);
and U21049 (N_21049,N_19063,N_19719);
and U21050 (N_21050,N_17274,N_19723);
and U21051 (N_21051,N_15674,N_16872);
nand U21052 (N_21052,N_17665,N_18109);
and U21053 (N_21053,N_17069,N_15160);
and U21054 (N_21054,N_17551,N_17531);
and U21055 (N_21055,N_17550,N_15040);
xnor U21056 (N_21056,N_17986,N_16690);
nor U21057 (N_21057,N_15953,N_18266);
or U21058 (N_21058,N_19944,N_19406);
nand U21059 (N_21059,N_18684,N_16608);
xnor U21060 (N_21060,N_18868,N_19314);
and U21061 (N_21061,N_18990,N_19991);
xnor U21062 (N_21062,N_19264,N_19172);
nor U21063 (N_21063,N_16210,N_16571);
xor U21064 (N_21064,N_17993,N_16943);
or U21065 (N_21065,N_16004,N_17587);
and U21066 (N_21066,N_19094,N_15252);
nand U21067 (N_21067,N_16008,N_15356);
and U21068 (N_21068,N_17932,N_19301);
nor U21069 (N_21069,N_17067,N_17896);
and U21070 (N_21070,N_15786,N_15531);
xor U21071 (N_21071,N_19895,N_16392);
or U21072 (N_21072,N_18666,N_16893);
xor U21073 (N_21073,N_16409,N_16084);
and U21074 (N_21074,N_17947,N_19205);
nor U21075 (N_21075,N_15159,N_17344);
or U21076 (N_21076,N_19784,N_18786);
xnor U21077 (N_21077,N_18444,N_16054);
and U21078 (N_21078,N_17511,N_17003);
xor U21079 (N_21079,N_18813,N_17605);
nand U21080 (N_21080,N_17885,N_18995);
nor U21081 (N_21081,N_16692,N_16373);
xor U21082 (N_21082,N_17840,N_17559);
nand U21083 (N_21083,N_15766,N_18688);
and U21084 (N_21084,N_19371,N_17042);
and U21085 (N_21085,N_17320,N_19387);
nor U21086 (N_21086,N_17357,N_15995);
nor U21087 (N_21087,N_15599,N_17488);
and U21088 (N_21088,N_16497,N_19283);
nand U21089 (N_21089,N_17922,N_18047);
nor U21090 (N_21090,N_15179,N_16973);
xor U21091 (N_21091,N_18789,N_17039);
or U21092 (N_21092,N_17413,N_17057);
nand U21093 (N_21093,N_17990,N_15775);
nor U21094 (N_21094,N_19227,N_17504);
nor U21095 (N_21095,N_15739,N_19868);
or U21096 (N_21096,N_15117,N_16610);
xnor U21097 (N_21097,N_17219,N_19829);
or U21098 (N_21098,N_19720,N_19910);
nor U21099 (N_21099,N_17105,N_18978);
nor U21100 (N_21100,N_17604,N_17563);
or U21101 (N_21101,N_18953,N_18862);
and U21102 (N_21102,N_15659,N_18693);
or U21103 (N_21103,N_19905,N_16387);
and U21104 (N_21104,N_19840,N_16207);
xnor U21105 (N_21105,N_16192,N_18380);
nor U21106 (N_21106,N_18346,N_16986);
and U21107 (N_21107,N_15295,N_15036);
and U21108 (N_21108,N_17832,N_15807);
xor U21109 (N_21109,N_15550,N_18094);
xor U21110 (N_21110,N_19473,N_16415);
nor U21111 (N_21111,N_18538,N_15519);
xor U21112 (N_21112,N_18488,N_18582);
nor U21113 (N_21113,N_15242,N_15802);
and U21114 (N_21114,N_18592,N_17784);
xor U21115 (N_21115,N_18885,N_18259);
nor U21116 (N_21116,N_18281,N_18033);
xor U21117 (N_21117,N_17112,N_18145);
and U21118 (N_21118,N_18757,N_19333);
xnor U21119 (N_21119,N_17657,N_19978);
nor U21120 (N_21120,N_17728,N_16306);
nor U21121 (N_21121,N_19286,N_15758);
or U21122 (N_21122,N_17696,N_17762);
or U21123 (N_21123,N_16547,N_15115);
nand U21124 (N_21124,N_17371,N_17131);
xnor U21125 (N_21125,N_19484,N_15576);
or U21126 (N_21126,N_19014,N_18944);
xor U21127 (N_21127,N_16938,N_15542);
or U21128 (N_21128,N_19037,N_19960);
and U21129 (N_21129,N_17538,N_17532);
nor U21130 (N_21130,N_16399,N_17358);
nand U21131 (N_21131,N_16722,N_18256);
xor U21132 (N_21132,N_18045,N_19110);
nand U21133 (N_21133,N_17402,N_19798);
nor U21134 (N_21134,N_19496,N_18542);
or U21135 (N_21135,N_16218,N_17206);
or U21136 (N_21136,N_16913,N_15409);
and U21137 (N_21137,N_16477,N_18634);
xor U21138 (N_21138,N_18746,N_17277);
and U21139 (N_21139,N_15035,N_15096);
or U21140 (N_21140,N_19838,N_17478);
nor U21141 (N_21141,N_17600,N_18575);
xor U21142 (N_21142,N_17755,N_18647);
nand U21143 (N_21143,N_16950,N_19721);
nor U21144 (N_21144,N_18787,N_15959);
or U21145 (N_21145,N_17411,N_15587);
nor U21146 (N_21146,N_17385,N_18119);
xnor U21147 (N_21147,N_19546,N_16739);
nand U21148 (N_21148,N_17761,N_18920);
xnor U21149 (N_21149,N_17648,N_18775);
or U21150 (N_21150,N_18858,N_18709);
xnor U21151 (N_21151,N_16785,N_16540);
nand U21152 (N_21152,N_18403,N_19485);
nand U21153 (N_21153,N_15173,N_18642);
nor U21154 (N_21154,N_16718,N_15203);
nand U21155 (N_21155,N_17262,N_16656);
and U21156 (N_21156,N_18241,N_18207);
or U21157 (N_21157,N_19483,N_19177);
nand U21158 (N_21158,N_19107,N_16573);
nor U21159 (N_21159,N_19362,N_16408);
and U21160 (N_21160,N_18579,N_17200);
xnor U21161 (N_21161,N_19775,N_15691);
nor U21162 (N_21162,N_18218,N_15951);
xnor U21163 (N_21163,N_18416,N_16448);
and U21164 (N_21164,N_15554,N_18999);
nand U21165 (N_21165,N_17324,N_17378);
or U21166 (N_21166,N_16092,N_15656);
xnor U21167 (N_21167,N_18052,N_16790);
xor U21168 (N_21168,N_19577,N_19505);
and U21169 (N_21169,N_19143,N_18265);
or U21170 (N_21170,N_17468,N_16041);
nand U21171 (N_21171,N_19222,N_19739);
and U21172 (N_21172,N_18449,N_17781);
or U21173 (N_21173,N_16584,N_16904);
nor U21174 (N_21174,N_18038,N_18792);
xor U21175 (N_21175,N_18993,N_19393);
nand U21176 (N_21176,N_18396,N_19138);
nand U21177 (N_21177,N_16418,N_16345);
xnor U21178 (N_21178,N_16433,N_18502);
xor U21179 (N_21179,N_15058,N_17684);
xnor U21180 (N_21180,N_16945,N_17342);
nand U21181 (N_21181,N_17525,N_18545);
and U21182 (N_21182,N_15026,N_15123);
and U21183 (N_21183,N_19180,N_16037);
xor U21184 (N_21184,N_19257,N_19555);
xnor U21185 (N_21185,N_15892,N_18846);
or U21186 (N_21186,N_15197,N_18525);
and U21187 (N_21187,N_19650,N_17283);
xor U21188 (N_21188,N_16556,N_15306);
nand U21189 (N_21189,N_19982,N_17179);
or U21190 (N_21190,N_17237,N_15355);
or U21191 (N_21191,N_16147,N_18998);
nand U21192 (N_21192,N_19228,N_19975);
nor U21193 (N_21193,N_18899,N_15974);
and U21194 (N_21194,N_19570,N_17751);
and U21195 (N_21195,N_18377,N_15903);
xnor U21196 (N_21196,N_19388,N_18476);
nand U21197 (N_21197,N_15153,N_15343);
and U21198 (N_21198,N_18633,N_15772);
nand U21199 (N_21199,N_16216,N_15768);
nand U21200 (N_21200,N_15191,N_18617);
xnor U21201 (N_21201,N_15154,N_15794);
nor U21202 (N_21202,N_17032,N_18711);
or U21203 (N_21203,N_18103,N_17944);
and U21204 (N_21204,N_17715,N_19044);
or U21205 (N_21205,N_18607,N_16012);
nor U21206 (N_21206,N_15432,N_16679);
xor U21207 (N_21207,N_17946,N_18303);
xnor U21208 (N_21208,N_16625,N_15220);
or U21209 (N_21209,N_19983,N_17242);
xor U21210 (N_21210,N_16304,N_16190);
nand U21211 (N_21211,N_17545,N_18050);
and U21212 (N_21212,N_15483,N_19245);
and U21213 (N_21213,N_16349,N_16140);
nor U21214 (N_21214,N_19694,N_19319);
and U21215 (N_21215,N_15319,N_15297);
or U21216 (N_21216,N_18818,N_16223);
nor U21217 (N_21217,N_16542,N_19011);
or U21218 (N_21218,N_17140,N_16864);
and U21219 (N_21219,N_15274,N_17061);
xor U21220 (N_21220,N_17138,N_17548);
nor U21221 (N_21221,N_19912,N_17091);
and U21222 (N_21222,N_18229,N_15425);
nand U21223 (N_21223,N_16970,N_18017);
xor U21224 (N_21224,N_18723,N_16269);
xnor U21225 (N_21225,N_16998,N_17129);
nor U21226 (N_21226,N_16821,N_15257);
nor U21227 (N_21227,N_19416,N_15711);
xor U21228 (N_21228,N_18173,N_19907);
xor U21229 (N_21229,N_18794,N_16736);
and U21230 (N_21230,N_17794,N_19202);
xor U21231 (N_21231,N_17460,N_18596);
xnor U21232 (N_21232,N_15404,N_15879);
nor U21233 (N_21233,N_17795,N_16065);
nor U21234 (N_21234,N_17496,N_17732);
or U21235 (N_21235,N_15643,N_17398);
or U21236 (N_21236,N_18866,N_18215);
or U21237 (N_21237,N_18645,N_16321);
nor U21238 (N_21238,N_15002,N_17505);
nor U21239 (N_21239,N_18086,N_17195);
nor U21240 (N_21240,N_15012,N_15199);
or U21241 (N_21241,N_18779,N_19968);
and U21242 (N_21242,N_17498,N_17598);
nor U21243 (N_21243,N_18320,N_18192);
nor U21244 (N_21244,N_15323,N_15654);
and U21245 (N_21245,N_17433,N_17019);
nand U21246 (N_21246,N_16721,N_16600);
nor U21247 (N_21247,N_15229,N_15695);
nor U21248 (N_21248,N_17166,N_15341);
xor U21249 (N_21249,N_19779,N_16645);
or U21250 (N_21250,N_19464,N_15613);
nor U21251 (N_21251,N_19289,N_15298);
or U21252 (N_21252,N_15391,N_17742);
nor U21253 (N_21253,N_17261,N_15563);
nand U21254 (N_21254,N_16725,N_19929);
or U21255 (N_21255,N_18166,N_15468);
nand U21256 (N_21256,N_16741,N_18110);
nand U21257 (N_21257,N_16588,N_16367);
xor U21258 (N_21258,N_18515,N_18179);
nor U21259 (N_21259,N_18041,N_18615);
nand U21260 (N_21260,N_18573,N_15291);
nor U21261 (N_21261,N_16447,N_19568);
nor U21262 (N_21262,N_16435,N_16993);
nand U21263 (N_21263,N_19691,N_16189);
nand U21264 (N_21264,N_16775,N_16560);
nor U21265 (N_21265,N_16205,N_17528);
nand U21266 (N_21266,N_15478,N_17231);
nor U21267 (N_21267,N_17758,N_15967);
or U21268 (N_21268,N_16465,N_16301);
and U21269 (N_21269,N_17331,N_17052);
nand U21270 (N_21270,N_18053,N_15579);
and U21271 (N_21271,N_19064,N_19705);
nor U21272 (N_21272,N_17668,N_19334);
nor U21273 (N_21273,N_19130,N_17142);
xor U21274 (N_21274,N_16130,N_19537);
nand U21275 (N_21275,N_17514,N_19807);
nor U21276 (N_21276,N_18513,N_18129);
xor U21277 (N_21277,N_17186,N_16747);
xnor U21278 (N_21278,N_17241,N_17602);
or U21279 (N_21279,N_17868,N_19120);
xnor U21280 (N_21280,N_18490,N_15935);
nor U21281 (N_21281,N_15911,N_19569);
xor U21282 (N_21282,N_15896,N_16413);
nor U21283 (N_21283,N_17902,N_15461);
and U21284 (N_21284,N_17148,N_15843);
or U21285 (N_21285,N_18945,N_17064);
or U21286 (N_21286,N_17146,N_17016);
or U21287 (N_21287,N_17855,N_15076);
xor U21288 (N_21288,N_15445,N_16602);
nand U21289 (N_21289,N_18609,N_18102);
nor U21290 (N_21290,N_16646,N_16483);
nor U21291 (N_21291,N_19031,N_16744);
nor U21292 (N_21292,N_19136,N_17230);
or U21293 (N_21293,N_16939,N_16033);
or U21294 (N_21294,N_18342,N_19749);
xnor U21295 (N_21295,N_18379,N_18785);
nor U21296 (N_21296,N_16609,N_17666);
nor U21297 (N_21297,N_18686,N_16696);
xor U21298 (N_21298,N_19218,N_17169);
xnor U21299 (N_21299,N_17681,N_15920);
nor U21300 (N_21300,N_19965,N_16730);
nor U21301 (N_21301,N_15500,N_15402);
nand U21302 (N_21302,N_16136,N_18389);
nand U21303 (N_21303,N_15335,N_15011);
or U21304 (N_21304,N_16716,N_19454);
xor U21305 (N_21305,N_19295,N_19941);
or U21306 (N_21306,N_18994,N_19594);
or U21307 (N_21307,N_16045,N_18649);
nand U21308 (N_21308,N_19239,N_19534);
nor U21309 (N_21309,N_16563,N_17144);
xnor U21310 (N_21310,N_15760,N_18989);
nand U21311 (N_21311,N_17322,N_15423);
and U21312 (N_21312,N_16503,N_17335);
nor U21313 (N_21313,N_19744,N_19828);
and U21314 (N_21314,N_17828,N_16348);
xnor U21315 (N_21315,N_16523,N_15368);
and U21316 (N_21316,N_16884,N_19550);
nand U21317 (N_21317,N_16111,N_19481);
nor U21318 (N_21318,N_16882,N_15473);
and U21319 (N_21319,N_18851,N_15224);
xnor U21320 (N_21320,N_15119,N_17407);
nand U21321 (N_21321,N_16765,N_15535);
or U21322 (N_21322,N_16779,N_16362);
or U21323 (N_21323,N_18701,N_15684);
nand U21324 (N_21324,N_16923,N_17646);
xor U21325 (N_21325,N_17899,N_19715);
or U21326 (N_21326,N_15603,N_18474);
or U21327 (N_21327,N_19999,N_18367);
and U21328 (N_21328,N_17172,N_16003);
or U21329 (N_21329,N_18603,N_18561);
or U21330 (N_21330,N_16764,N_18765);
nand U21331 (N_21331,N_16583,N_16398);
and U21332 (N_21332,N_15004,N_16616);
xnor U21333 (N_21333,N_18443,N_15369);
nand U21334 (N_21334,N_15577,N_15038);
nor U21335 (N_21335,N_16230,N_19961);
xor U21336 (N_21336,N_19165,N_18522);
nor U21337 (N_21337,N_19131,N_16453);
nand U21338 (N_21338,N_17113,N_15575);
xnor U21339 (N_21339,N_18206,N_19377);
and U21340 (N_21340,N_19084,N_18315);
nor U21341 (N_21341,N_19115,N_15469);
and U21342 (N_21342,N_18243,N_16731);
nand U21343 (N_21343,N_18555,N_17629);
nor U21344 (N_21344,N_18162,N_18113);
nor U21345 (N_21345,N_15052,N_18140);
or U21346 (N_21346,N_17269,N_19455);
or U21347 (N_21347,N_18896,N_18188);
xnor U21348 (N_21348,N_15264,N_15301);
or U21349 (N_21349,N_17685,N_16183);
and U21350 (N_21350,N_17383,N_19733);
nor U21351 (N_21351,N_17543,N_19735);
and U21352 (N_21352,N_17912,N_17610);
and U21353 (N_21353,N_19792,N_19959);
nor U21354 (N_21354,N_19890,N_18035);
nand U21355 (N_21355,N_16078,N_18710);
and U21356 (N_21356,N_15570,N_18675);
and U21357 (N_21357,N_15553,N_19887);
or U21358 (N_21358,N_16559,N_15394);
xnor U21359 (N_21359,N_18935,N_16890);
and U21360 (N_21360,N_15457,N_19474);
nor U21361 (N_21361,N_15283,N_17904);
and U21362 (N_21362,N_16251,N_18366);
and U21363 (N_21363,N_16879,N_15928);
nor U21364 (N_21364,N_19451,N_18276);
nand U21365 (N_21365,N_17890,N_19472);
and U21366 (N_21366,N_18067,N_15050);
nand U21367 (N_21367,N_18921,N_16290);
nand U21368 (N_21368,N_19041,N_15682);
and U21369 (N_21369,N_18938,N_17995);
xnor U21370 (N_21370,N_18741,N_15502);
nand U21371 (N_21371,N_16347,N_16187);
and U21372 (N_21372,N_18939,N_17535);
and U21373 (N_21373,N_17653,N_18009);
and U21374 (N_21374,N_18546,N_18252);
xnor U21375 (N_21375,N_16796,N_15699);
nand U21376 (N_21376,N_15364,N_15014);
nor U21377 (N_21377,N_15498,N_18996);
and U21378 (N_21378,N_16977,N_17725);
or U21379 (N_21379,N_15752,N_18682);
nand U21380 (N_21380,N_15126,N_15747);
and U21381 (N_21381,N_18752,N_19606);
xnor U21382 (N_21382,N_16965,N_18783);
and U21383 (N_21383,N_19636,N_16107);
and U21384 (N_21384,N_16271,N_19299);
and U21385 (N_21385,N_17111,N_17133);
nor U21386 (N_21386,N_15990,N_18390);
or U21387 (N_21387,N_16577,N_18796);
xor U21388 (N_21388,N_17430,N_18288);
or U21389 (N_21389,N_17429,N_15324);
nor U21390 (N_21390,N_18698,N_16145);
and U21391 (N_21391,N_19670,N_15729);
xnor U21392 (N_21392,N_17888,N_19164);
nand U21393 (N_21393,N_18030,N_19376);
nor U21394 (N_21394,N_19317,N_16789);
and U21395 (N_21395,N_16532,N_18124);
and U21396 (N_21396,N_19125,N_15660);
nor U21397 (N_21397,N_19717,N_15832);
nand U21398 (N_21398,N_16618,N_15137);
xor U21399 (N_21399,N_17275,N_15102);
nor U21400 (N_21400,N_15561,N_16755);
nand U21401 (N_21401,N_15818,N_15968);
xnor U21402 (N_21402,N_16719,N_18637);
xnor U21403 (N_21403,N_18270,N_19585);
or U21404 (N_21404,N_19990,N_17907);
or U21405 (N_21405,N_18074,N_19261);
or U21406 (N_21406,N_17886,N_16009);
or U21407 (N_21407,N_16901,N_18227);
xnor U21408 (N_21408,N_17941,N_18962);
nor U21409 (N_21409,N_15714,N_15240);
xor U21410 (N_21410,N_18356,N_19089);
nand U21411 (N_21411,N_17381,N_17623);
nand U21412 (N_21412,N_18430,N_15125);
or U21413 (N_21413,N_18139,N_17384);
nand U21414 (N_21414,N_19817,N_15176);
xor U21415 (N_21415,N_19058,N_19347);
xnor U21416 (N_21416,N_18373,N_16813);
or U21417 (N_21417,N_15831,N_17115);
or U21418 (N_21418,N_18685,N_16512);
xor U21419 (N_21419,N_15408,N_19816);
and U21420 (N_21420,N_18558,N_18048);
nand U21421 (N_21421,N_18337,N_17068);
nor U21422 (N_21422,N_15462,N_17440);
and U21423 (N_21423,N_19034,N_18087);
or U21424 (N_21424,N_15081,N_18946);
nand U21425 (N_21425,N_18332,N_15260);
nand U21426 (N_21426,N_19994,N_18734);
or U21427 (N_21427,N_16989,N_17727);
and U21428 (N_21428,N_18408,N_16644);
nand U21429 (N_21429,N_19424,N_19223);
nand U21430 (N_21430,N_18918,N_16727);
or U21431 (N_21431,N_17031,N_17576);
or U21432 (N_21432,N_19200,N_15948);
and U21433 (N_21433,N_15919,N_18199);
or U21434 (N_21434,N_17826,N_15042);
or U21435 (N_21435,N_19680,N_19734);
nor U21436 (N_21436,N_18060,N_16895);
nor U21437 (N_21437,N_16680,N_15872);
and U21438 (N_21438,N_16283,N_17965);
or U21439 (N_21439,N_16506,N_17053);
and U21440 (N_21440,N_17649,N_15647);
xnor U21441 (N_21441,N_19687,N_19287);
xor U21442 (N_21442,N_16225,N_16801);
or U21443 (N_21443,N_18894,N_17915);
nand U21444 (N_21444,N_19693,N_15079);
or U21445 (N_21445,N_18539,N_16036);
or U21446 (N_21446,N_17508,N_19969);
nor U21447 (N_21447,N_18529,N_17155);
nor U21448 (N_21448,N_17931,N_19008);
or U21449 (N_21449,N_19013,N_16377);
nor U21450 (N_21450,N_19501,N_17988);
or U21451 (N_21451,N_19859,N_19036);
nor U21452 (N_21452,N_17590,N_17246);
nand U21453 (N_21453,N_15734,N_15604);
or U21454 (N_21454,N_15201,N_17801);
xnor U21455 (N_21455,N_18482,N_17618);
or U21456 (N_21456,N_16305,N_17652);
and U21457 (N_21457,N_19616,N_15433);
xnor U21458 (N_21458,N_18578,N_19697);
xnor U21459 (N_21459,N_15420,N_19316);
xnor U21460 (N_21460,N_16572,N_16234);
nand U21461 (N_21461,N_15689,N_19203);
and U21462 (N_21462,N_19067,N_16883);
nand U21463 (N_21463,N_16566,N_17808);
or U21464 (N_21464,N_16060,N_18042);
nor U21465 (N_21465,N_17006,N_18345);
and U21466 (N_21466,N_17621,N_17804);
xnor U21467 (N_21467,N_19911,N_15544);
or U21468 (N_21468,N_15840,N_19942);
nand U21469 (N_21469,N_17130,N_19055);
nor U21470 (N_21470,N_18327,N_15649);
nor U21471 (N_21471,N_17937,N_17107);
or U21472 (N_21472,N_18836,N_18674);
xor U21473 (N_21473,N_19061,N_18211);
nor U21474 (N_21474,N_17493,N_17916);
or U21475 (N_21475,N_17034,N_18185);
and U21476 (N_21476,N_17676,N_18780);
nor U21477 (N_21477,N_15978,N_17106);
or U21478 (N_21478,N_19432,N_15400);
nand U21479 (N_21479,N_19375,N_19954);
and U21480 (N_21480,N_16125,N_17991);
or U21481 (N_21481,N_17744,N_17459);
nor U21482 (N_21482,N_18092,N_18148);
or U21483 (N_21483,N_19955,N_18949);
xnor U21484 (N_21484,N_16498,N_17228);
or U21485 (N_21485,N_17084,N_19622);
xnor U21486 (N_21486,N_19836,N_19370);
or U21487 (N_21487,N_16296,N_19649);
nor U21488 (N_21488,N_17699,N_16492);
xor U21489 (N_21489,N_17259,N_15586);
and U21490 (N_21490,N_19541,N_16194);
nor U21491 (N_21491,N_18853,N_15345);
nor U21492 (N_21492,N_15127,N_15873);
or U21493 (N_21493,N_16522,N_16635);
nand U21494 (N_21494,N_17072,N_15370);
or U21495 (N_21495,N_15281,N_18650);
and U21496 (N_21496,N_18669,N_19879);
and U21497 (N_21497,N_15112,N_18205);
and U21498 (N_21498,N_16653,N_18032);
xor U21499 (N_21499,N_19908,N_17766);
xnor U21500 (N_21500,N_19642,N_16894);
xnor U21501 (N_21501,N_16726,N_19529);
nand U21502 (N_21502,N_15982,N_15590);
nand U21503 (N_21503,N_17147,N_19939);
xor U21504 (N_21504,N_17637,N_17139);
xnor U21505 (N_21505,N_17470,N_17074);
and U21506 (N_21506,N_15362,N_16062);
or U21507 (N_21507,N_19872,N_15043);
or U21508 (N_21508,N_18200,N_18251);
nand U21509 (N_21509,N_16667,N_19777);
nand U21510 (N_21510,N_15411,N_15321);
nand U21511 (N_21511,N_18577,N_19059);
or U21512 (N_21512,N_17028,N_16910);
nor U21513 (N_21513,N_15208,N_18948);
xor U21514 (N_21514,N_15198,N_16876);
nand U21515 (N_21515,N_15236,N_16593);
nor U21516 (N_21516,N_18261,N_19140);
or U21517 (N_21517,N_15382,N_15437);
and U21518 (N_21518,N_18081,N_15431);
and U21519 (N_21519,N_17125,N_18627);
nor U21520 (N_21520,N_18465,N_16169);
or U21521 (N_21521,N_16920,N_19985);
nand U21522 (N_21522,N_16838,N_19522);
xnor U21523 (N_21523,N_16411,N_16666);
and U21524 (N_21524,N_19389,N_18453);
xnor U21525 (N_21525,N_19308,N_18043);
nor U21526 (N_21526,N_15235,N_15779);
and U21527 (N_21527,N_18516,N_18404);
nand U21528 (N_21528,N_16171,N_15690);
nor U21529 (N_21529,N_19175,N_15376);
nor U21530 (N_21530,N_18613,N_18483);
xnor U21531 (N_21531,N_19762,N_15292);
nand U21532 (N_21532,N_18600,N_18003);
and U21533 (N_21533,N_15769,N_18002);
or U21534 (N_21534,N_18588,N_19369);
or U21535 (N_21535,N_17642,N_19790);
and U21536 (N_21536,N_17165,N_18901);
xnor U21537 (N_21537,N_17484,N_18029);
or U21538 (N_21538,N_19519,N_19183);
nand U21539 (N_21539,N_15655,N_19818);
and U21540 (N_21540,N_17054,N_18611);
and U21541 (N_21541,N_19410,N_18280);
and U21542 (N_21542,N_19950,N_17159);
nand U21543 (N_21543,N_16097,N_19303);
xnor U21544 (N_21544,N_15859,N_19382);
nand U21545 (N_21545,N_18743,N_16115);
nor U21546 (N_21546,N_18232,N_16338);
and U21547 (N_21547,N_19783,N_19871);
or U21548 (N_21548,N_16310,N_15773);
and U21549 (N_21549,N_17952,N_15532);
or U21550 (N_21550,N_19951,N_15352);
nor U21551 (N_21551,N_15515,N_15641);
nand U21552 (N_21552,N_18202,N_15858);
or U21553 (N_21553,N_17103,N_16421);
and U21554 (N_21554,N_15289,N_15977);
nor U21555 (N_21555,N_19056,N_19506);
nand U21556 (N_21556,N_17848,N_15474);
nand U21557 (N_21557,N_17395,N_18305);
or U21558 (N_21558,N_17327,N_16382);
nand U21559 (N_21559,N_18459,N_19086);
or U21560 (N_21560,N_19820,N_17566);
xnor U21561 (N_21561,N_16055,N_15547);
nor U21562 (N_21562,N_15359,N_16990);
or U21563 (N_21563,N_18526,N_19104);
and U21564 (N_21564,N_16587,N_16886);
nor U21565 (N_21565,N_18657,N_16475);
and U21566 (N_21566,N_18651,N_19071);
or U21567 (N_21567,N_18825,N_15882);
nand U21568 (N_21568,N_19475,N_16712);
nand U21569 (N_21569,N_18740,N_19294);
or U21570 (N_21570,N_19679,N_16881);
or U21571 (N_21571,N_16619,N_18904);
xor U21572 (N_21572,N_18950,N_17116);
or U21573 (N_21573,N_18049,N_17985);
and U21574 (N_21574,N_16623,N_15330);
nand U21575 (N_21575,N_15512,N_16561);
nor U21576 (N_21576,N_17822,N_16030);
or U21577 (N_21577,N_15120,N_15893);
or U21578 (N_21578,N_17143,N_17881);
nor U21579 (N_21579,N_17934,N_16394);
xnor U21580 (N_21580,N_18801,N_17584);
nand U21581 (N_21581,N_19178,N_15909);
or U21582 (N_21582,N_15262,N_18437);
xnor U21583 (N_21583,N_18221,N_19343);
and U21584 (N_21584,N_19948,N_17811);
and U21585 (N_21585,N_17734,N_19070);
or U21586 (N_21586,N_16677,N_16684);
xnor U21587 (N_21587,N_16038,N_18821);
and U21588 (N_21588,N_17232,N_16786);
and U21589 (N_21589,N_16063,N_19565);
nor U21590 (N_21590,N_19553,N_19945);
and U21591 (N_21591,N_19193,N_18419);
nor U21592 (N_21592,N_16266,N_17724);
xor U21593 (N_21593,N_18756,N_19017);
and U21594 (N_21594,N_18066,N_19087);
and U21595 (N_21595,N_16850,N_15028);
nor U21596 (N_21596,N_19793,N_18888);
nor U21597 (N_21597,N_19549,N_19666);
xor U21598 (N_21598,N_19979,N_18418);
xnor U21599 (N_21599,N_19696,N_15001);
and U21600 (N_21600,N_16109,N_19781);
xor U21601 (N_21601,N_16018,N_17036);
or U21602 (N_21602,N_19390,N_18580);
or U21603 (N_21603,N_19964,N_16089);
xnor U21604 (N_21604,N_17747,N_19422);
or U21605 (N_21605,N_18245,N_15564);
xnor U21606 (N_21606,N_19150,N_19692);
xnor U21607 (N_21607,N_19123,N_15401);
nor U21608 (N_21608,N_17035,N_16580);
and U21609 (N_21609,N_18085,N_17936);
xnor U21610 (N_21610,N_15133,N_15407);
or U21611 (N_21611,N_16146,N_15666);
or U21612 (N_21612,N_16549,N_17573);
xnor U21613 (N_21613,N_19166,N_15080);
or U21614 (N_21614,N_15143,N_15099);
and U21615 (N_21615,N_19809,N_19398);
xnor U21616 (N_21616,N_19437,N_19808);
and U21617 (N_21617,N_18401,N_17628);
xnor U21618 (N_21618,N_17805,N_16164);
xnor U21619 (N_21619,N_17475,N_16737);
or U21620 (N_21620,N_17382,N_16988);
nand U21621 (N_21621,N_17625,N_18543);
nor U21622 (N_21622,N_19226,N_16002);
xnor U21623 (N_21623,N_15087,N_19213);
or U21624 (N_21624,N_16355,N_19477);
nor U21625 (N_21625,N_17940,N_17661);
and U21626 (N_21626,N_15665,N_17837);
or U21627 (N_21627,N_19349,N_16121);
and U21628 (N_21628,N_19737,N_17163);
nand U21629 (N_21629,N_15017,N_15770);
xor U21630 (N_21630,N_17647,N_16907);
and U21631 (N_21631,N_15460,N_19470);
and U21632 (N_21632,N_18089,N_17785);
xor U21633 (N_21633,N_19173,N_16246);
and U21634 (N_21634,N_17349,N_18480);
nand U21635 (N_21635,N_15743,N_17809);
nand U21636 (N_21636,N_18598,N_18506);
nor U21637 (N_21637,N_18849,N_17434);
or U21638 (N_21638,N_19345,N_17007);
or U21639 (N_21639,N_15385,N_15852);
nor U21640 (N_21640,N_17851,N_16277);
or U21641 (N_21641,N_17367,N_16622);
xor U21642 (N_21642,N_15778,N_16810);
xor U21643 (N_21643,N_17160,N_16067);
or U21644 (N_21644,N_17345,N_15493);
xnor U21645 (N_21645,N_17825,N_16403);
nand U21646 (N_21646,N_19381,N_18514);
nor U21647 (N_21647,N_19923,N_16391);
nand U21648 (N_21648,N_18560,N_19111);
or U21649 (N_21649,N_17152,N_17294);
nand U21650 (N_21650,N_17190,N_17212);
nand U21651 (N_21651,N_16856,N_19864);
or U21652 (N_21652,N_17677,N_19153);
xnor U21653 (N_21653,N_15340,N_18452);
nor U21654 (N_21654,N_18623,N_19225);
and U21655 (N_21655,N_18472,N_15946);
or U21656 (N_21656,N_16019,N_16815);
nor U21657 (N_21657,N_16352,N_15804);
xor U21658 (N_21658,N_19280,N_16639);
nor U21659 (N_21659,N_15302,N_16402);
xor U21660 (N_21660,N_16168,N_18536);
nand U21661 (N_21661,N_16047,N_16247);
or U21662 (N_21662,N_15986,N_18371);
and U21663 (N_21663,N_16968,N_17201);
xor U21664 (N_21664,N_15623,N_19738);
xnor U21665 (N_21665,N_19459,N_15625);
or U21666 (N_21666,N_19998,N_19826);
and U21667 (N_21667,N_16077,N_15272);
and U21668 (N_21668,N_18246,N_19925);
nor U21669 (N_21669,N_16724,N_19321);
and U21670 (N_21670,N_16576,N_18144);
nand U21671 (N_21671,N_18180,N_17365);
nor U21672 (N_21672,N_19497,N_19767);
and U21673 (N_21673,N_15790,N_17472);
and U21674 (N_21674,N_18719,N_15700);
or U21675 (N_21675,N_18204,N_18428);
nand U21676 (N_21676,N_18153,N_16931);
nand U21677 (N_21677,N_16069,N_18583);
xor U21678 (N_21678,N_18381,N_19984);
xor U21679 (N_21679,N_18807,N_17156);
or U21680 (N_21680,N_19162,N_16080);
nand U21681 (N_21681,N_15914,N_16228);
nor U21682 (N_21682,N_19220,N_16665);
and U21683 (N_21683,N_16135,N_19943);
and U21684 (N_21684,N_17547,N_16293);
nand U21685 (N_21685,N_16738,N_16985);
nand U21686 (N_21686,N_19770,N_19822);
nor U21687 (N_21687,N_19922,N_18565);
nand U21688 (N_21688,N_17707,N_16152);
xor U21689 (N_21689,N_17942,N_15156);
xor U21690 (N_21690,N_15390,N_18706);
nand U21691 (N_21691,N_18068,N_17585);
nor U21692 (N_21692,N_18929,N_15481);
nand U21693 (N_21693,N_15479,N_17001);
and U21694 (N_21694,N_15259,N_17775);
or U21695 (N_21695,N_15347,N_17083);
or U21696 (N_21696,N_19850,N_17267);
xnor U21697 (N_21697,N_15732,N_17753);
xor U21698 (N_21698,N_16386,N_15984);
or U21699 (N_21699,N_17608,N_19009);
and U21700 (N_21700,N_15942,N_15074);
or U21701 (N_21701,N_18334,N_19601);
xor U21702 (N_21702,N_17182,N_16103);
or U21703 (N_21703,N_18931,N_19458);
and U21704 (N_21704,N_18788,N_15728);
xnor U21705 (N_21705,N_19893,N_15958);
nand U21706 (N_21706,N_17750,N_19212);
or U21707 (N_21707,N_16467,N_18547);
or U21708 (N_21708,N_17945,N_16100);
or U21709 (N_21709,N_15720,N_15098);
nor U21710 (N_21710,N_18454,N_16885);
nand U21711 (N_21711,N_17688,N_18387);
nor U21712 (N_21712,N_17963,N_17497);
nor U21713 (N_21713,N_18456,N_19527);
nand U21714 (N_21714,N_17258,N_17984);
and U21715 (N_21715,N_17396,N_19703);
xor U21716 (N_21716,N_18331,N_16276);
nand U21717 (N_21717,N_17894,N_15650);
or U21718 (N_21718,N_19851,N_15169);
and U21719 (N_21719,N_19581,N_19683);
xor U21720 (N_21720,N_19326,N_18360);
xnor U21721 (N_21721,N_15993,N_16366);
nor U21722 (N_21722,N_15759,N_19819);
or U21723 (N_21723,N_15726,N_18413);
or U21724 (N_21724,N_18718,N_16565);
and U21725 (N_21725,N_16809,N_18571);
nand U21726 (N_21726,N_16236,N_16607);
or U21727 (N_21727,N_16474,N_17634);
xor U21728 (N_21728,N_17659,N_16287);
xnor U21729 (N_21729,N_16158,N_16905);
nand U21730 (N_21730,N_16098,N_18432);
and U21731 (N_21731,N_18228,N_15422);
xor U21732 (N_21732,N_15174,N_17627);
nand U21733 (N_21733,N_16927,N_19278);
and U21734 (N_21734,N_15279,N_19135);
nor U21735 (N_21735,N_18329,N_17004);
xnor U21736 (N_21736,N_15348,N_16022);
nand U21737 (N_21737,N_18881,N_18463);
nand U21738 (N_21738,N_19710,N_18004);
or U21739 (N_21739,N_17392,N_15334);
xor U21740 (N_21740,N_15318,N_18301);
xor U21741 (N_21741,N_16564,N_19847);
and U21742 (N_21742,N_17339,N_16676);
and U21743 (N_21743,N_15783,N_15161);
or U21744 (N_21744,N_19811,N_16756);
and U21745 (N_21745,N_16659,N_16203);
and U21746 (N_21746,N_18203,N_15584);
xnor U21747 (N_21747,N_18425,N_18541);
nand U21748 (N_21748,N_15536,N_17910);
nor U21749 (N_21749,N_18486,N_17726);
nand U21750 (N_21750,N_15744,N_18632);
nor U21751 (N_21751,N_15132,N_17312);
and U21752 (N_21752,N_16900,N_18635);
nand U21753 (N_21753,N_19888,N_16992);
xnor U21754 (N_21754,N_19667,N_16257);
or U21755 (N_21755,N_19987,N_16935);
or U21756 (N_21756,N_15742,N_17466);
and U21757 (N_21757,N_19620,N_19399);
xor U21758 (N_21758,N_17928,N_16117);
nor U21759 (N_21759,N_19018,N_19740);
xnor U21760 (N_21760,N_18562,N_18116);
xor U21761 (N_21761,N_15667,N_18198);
and U21762 (N_21762,N_16757,N_19671);
xnor U21763 (N_21763,N_18257,N_16016);
xnor U21764 (N_21764,N_18958,N_19206);
xor U21765 (N_21765,N_19452,N_15596);
and U21766 (N_21766,N_16529,N_15989);
nand U21767 (N_21767,N_18566,N_17391);
xor U21768 (N_21768,N_18895,N_17778);
nor U21769 (N_21769,N_17549,N_15309);
xor U21770 (N_21770,N_15640,N_16877);
nand U21771 (N_21771,N_18344,N_17883);
nor U21772 (N_21772,N_16701,N_17409);
nand U21773 (N_21773,N_19365,N_16683);
xor U21774 (N_21774,N_18037,N_15856);
or U21775 (N_21775,N_15863,N_19417);
or U21776 (N_21776,N_19005,N_15639);
and U21777 (N_21777,N_15851,N_17534);
xnor U21778 (N_21778,N_15880,N_15162);
and U21779 (N_21779,N_17656,N_18149);
nor U21780 (N_21780,N_17175,N_16381);
xor U21781 (N_21781,N_15476,N_18182);
nor U21782 (N_21782,N_19794,N_17400);
xor U21783 (N_21783,N_17506,N_18735);
nand U21784 (N_21784,N_16866,N_17483);
and U21785 (N_21785,N_18370,N_19891);
nand U21786 (N_21786,N_19456,N_18806);
xnor U21787 (N_21787,N_16915,N_15627);
or U21788 (N_21788,N_17295,N_18915);
or U21789 (N_21789,N_18226,N_19980);
nor U21790 (N_21790,N_15602,N_17013);
nand U21791 (N_21791,N_19920,N_17983);
xnor U21792 (N_21792,N_19873,N_19114);
nor U21793 (N_21793,N_16404,N_18475);
xnor U21794 (N_21794,N_18407,N_18115);
xor U21795 (N_21795,N_18313,N_16328);
nand U21796 (N_21796,N_17127,N_15077);
nand U21797 (N_21797,N_16515,N_18118);
nand U21798 (N_21798,N_16471,N_15996);
or U21799 (N_21799,N_19476,N_15051);
xor U21800 (N_21800,N_19281,N_18975);
xnor U21801 (N_21801,N_15200,N_16020);
nor U21802 (N_21802,N_19385,N_18365);
xor U21803 (N_21803,N_16319,N_16202);
nor U21804 (N_21804,N_16374,N_19706);
nand U21805 (N_21805,N_18879,N_16562);
and U21806 (N_21806,N_19208,N_17919);
and U21807 (N_21807,N_17858,N_17889);
and U21808 (N_21808,N_18759,N_16091);
nor U21809 (N_21809,N_18922,N_17971);
or U21810 (N_21810,N_18980,N_19634);
nor U21811 (N_21811,N_15956,N_18823);
nor U21812 (N_21812,N_16441,N_19364);
nor U21813 (N_21813,N_18564,N_15333);
or U21814 (N_21814,N_17361,N_15583);
xor U21815 (N_21815,N_17442,N_17319);
and U21816 (N_21816,N_17253,N_18269);
xnor U21817 (N_21817,N_15835,N_19419);
nor U21818 (N_21818,N_15608,N_17002);
xnor U21819 (N_21819,N_16554,N_19684);
nand U21820 (N_21820,N_18934,N_16808);
nand U21821 (N_21821,N_18773,N_17435);
xor U21822 (N_21822,N_19216,N_16139);
nand U21823 (N_21823,N_16581,N_15952);
and U21824 (N_21824,N_19966,N_15600);
xnor U21825 (N_21825,N_15620,N_19646);
nand U21826 (N_21826,N_18071,N_16750);
nor U21827 (N_21827,N_19621,N_16280);
or U21828 (N_21828,N_19880,N_15083);
and U21829 (N_21829,N_16887,N_16299);
xnor U21830 (N_21830,N_16936,N_15185);
xor U21831 (N_21831,N_15846,N_19310);
and U21832 (N_21832,N_15653,N_19709);
xor U21833 (N_21833,N_16963,N_19159);
nor U21834 (N_21834,N_19440,N_18410);
nand U21835 (N_21835,N_15670,N_15866);
and U21836 (N_21836,N_17954,N_16825);
nand U21837 (N_21837,N_19886,N_18625);
nor U21838 (N_21838,N_19536,N_16596);
or U21839 (N_21839,N_17964,N_19339);
nor U21840 (N_21840,N_16058,N_19080);
and U21841 (N_21841,N_16087,N_17043);
nand U21842 (N_21842,N_18392,N_17786);
nor U21843 (N_21843,N_18764,N_15441);
and U21844 (N_21844,N_19255,N_16221);
nor U21845 (N_21845,N_16094,N_19862);
and U21846 (N_21846,N_16997,N_15957);
and U21847 (N_21847,N_17329,N_15696);
nor U21848 (N_21848,N_15108,N_18745);
nand U21849 (N_21849,N_19825,N_17650);
nor U21850 (N_21850,N_18267,N_15436);
xor U21851 (N_21851,N_16720,N_17779);
or U21852 (N_21852,N_19322,N_19678);
or U21853 (N_21853,N_15451,N_15158);
and U21854 (N_21854,N_18909,N_17223);
and U21855 (N_21855,N_18593,N_15530);
or U21856 (N_21856,N_17765,N_15139);
nor U21857 (N_21857,N_17746,N_19677);
xor U21858 (N_21858,N_19530,N_17346);
nand U21859 (N_21859,N_17060,N_16713);
or U21860 (N_21860,N_17720,N_16101);
nand U21861 (N_21861,N_19947,N_15190);
xor U21862 (N_21862,N_17307,N_16655);
xor U21863 (N_21863,N_18311,N_16142);
xor U21864 (N_21864,N_19256,N_18882);
or U21865 (N_21865,N_18952,N_19214);
nor U21866 (N_21866,N_19233,N_16279);
and U21867 (N_21867,N_17897,N_16788);
and U21868 (N_21868,N_16914,N_16369);
and U21869 (N_21869,N_18605,N_15821);
and U21870 (N_21870,N_15003,N_16728);
nor U21871 (N_21871,N_16686,N_15233);
and U21872 (N_21872,N_15344,N_16509);
or U21873 (N_21873,N_19599,N_19771);
xor U21874 (N_21874,N_17522,N_19504);
xor U21875 (N_21875,N_15263,N_18557);
nor U21876 (N_21876,N_15594,N_17501);
nor U21877 (N_21877,N_16072,N_17189);
or U21878 (N_21878,N_16325,N_16928);
nand U21879 (N_21879,N_16197,N_17141);
xnor U21880 (N_21880,N_17462,N_18928);
and U21881 (N_21881,N_16752,N_17635);
nand U21882 (N_21882,N_15991,N_15980);
nor U21883 (N_21883,N_17594,N_19441);
nor U21884 (N_21884,N_19782,N_18414);
nand U21885 (N_21885,N_18326,N_17749);
nand U21886 (N_21886,N_15677,N_15157);
nor U21887 (N_21887,N_19837,N_19427);
nand U21888 (N_21888,N_18856,N_17088);
and U21889 (N_21889,N_16426,N_19429);
nor U21890 (N_21890,N_16444,N_15393);
or U21891 (N_21891,N_19285,N_15072);
nor U21892 (N_21892,N_16934,N_19372);
nor U21893 (N_21893,N_18263,N_16326);
nand U21894 (N_21894,N_18988,N_17257);
or U21895 (N_21895,N_17426,N_15093);
or U21896 (N_21896,N_16268,N_17968);
and U21897 (N_21897,N_18167,N_17420);
and U21898 (N_21898,N_17633,N_19461);
nand U21899 (N_21899,N_19631,N_19637);
or U21900 (N_21900,N_15486,N_17099);
xor U21901 (N_21901,N_17227,N_18653);
xnor U21902 (N_21902,N_16698,N_19361);
or U21903 (N_21903,N_16401,N_15065);
or U21904 (N_21904,N_19211,N_16432);
nor U21905 (N_21905,N_16769,N_16732);
nand U21906 (N_21906,N_15388,N_16237);
and U21907 (N_21907,N_19755,N_19082);
or U21908 (N_21908,N_15192,N_19856);
nor U21909 (N_21909,N_16528,N_17040);
xor U21910 (N_21910,N_17686,N_17476);
nand U21911 (N_21911,N_17234,N_18869);
nor U21912 (N_21912,N_15332,N_19796);
nor U21913 (N_21913,N_15837,N_15487);
or U21914 (N_21914,N_15784,N_18570);
nor U21915 (N_21915,N_19532,N_17096);
nor U21916 (N_21916,N_19831,N_17214);
or U21917 (N_21917,N_17422,N_19189);
nor U21918 (N_21918,N_17245,N_17380);
or U21919 (N_21919,N_15237,N_16615);
nand U21920 (N_21920,N_16014,N_16806);
or U21921 (N_21921,N_16550,N_16918);
xor U21922 (N_21922,N_19288,N_18084);
xnor U21923 (N_21923,N_19662,N_19543);
nor U21924 (N_21924,N_16818,N_16430);
nor U21925 (N_21925,N_18260,N_15387);
nor U21926 (N_21926,N_19833,N_15994);
nor U21927 (N_21927,N_15317,N_18178);
or U21928 (N_21928,N_15960,N_18496);
and U21929 (N_21929,N_17893,N_18854);
nand U21930 (N_21930,N_19030,N_17264);
and U21931 (N_21931,N_17872,N_19457);
and U21932 (N_21932,N_15545,N_15234);
or U21933 (N_21933,N_15999,N_17519);
nand U21934 (N_21934,N_19074,N_15585);
or U21935 (N_21935,N_16702,N_19688);
nor U21936 (N_21936,N_15091,N_18984);
nor U21937 (N_21937,N_17009,N_15806);
nor U21938 (N_21938,N_19835,N_17467);
xor U21939 (N_21939,N_19672,N_19184);
nand U21940 (N_21940,N_17626,N_18467);
and U21941 (N_21941,N_17892,N_19633);
and U21942 (N_21942,N_15379,N_15616);
xnor U21943 (N_21943,N_16157,N_19884);
xor U21944 (N_21944,N_18620,N_17406);
or U21945 (N_21945,N_18484,N_16160);
nand U21946 (N_21946,N_16922,N_18078);
nor U21947 (N_21947,N_16835,N_15795);
nand U21948 (N_21948,N_19029,N_17706);
xor U21949 (N_21949,N_15049,N_15329);
nand U21950 (N_21950,N_15652,N_17575);
nand U21951 (N_21951,N_15510,N_16762);
xnor U21952 (N_21952,N_15282,N_17491);
or U21953 (N_21953,N_19865,N_15782);
and U21954 (N_21954,N_16634,N_19279);
xor U21955 (N_21955,N_16446,N_19119);
nor U21956 (N_21956,N_17836,N_15534);
nand U21957 (N_21957,N_16336,N_16102);
xnor U21958 (N_21958,N_19963,N_19725);
xnor U21959 (N_21959,N_17884,N_16613);
or U21960 (N_21960,N_18554,N_17403);
or U21961 (N_21961,N_18969,N_19290);
or U21962 (N_21962,N_16627,N_17203);
nand U21963 (N_21963,N_19237,N_17595);
and U21964 (N_21964,N_15466,N_19296);
xor U21965 (N_21965,N_17437,N_18364);
xnor U21966 (N_21966,N_17839,N_15558);
xnor U21967 (N_21967,N_15875,N_16749);
xor U21968 (N_21968,N_16517,N_18643);
xor U21969 (N_21969,N_19647,N_15459);
nor U21970 (N_21970,N_19787,N_17046);
or U21971 (N_21971,N_19605,N_18878);
nand U21972 (N_21972,N_18861,N_17114);
xnor U21973 (N_21973,N_19075,N_16846);
or U21974 (N_21974,N_19331,N_17556);
nor U21975 (N_21975,N_16393,N_15328);
nand U21976 (N_21976,N_15947,N_15475);
xnor U21977 (N_21977,N_19915,N_16648);
and U21978 (N_21978,N_17082,N_15707);
or U21979 (N_21979,N_16689,N_15211);
and U21980 (N_21980,N_17973,N_18707);
xor U21981 (N_21981,N_15204,N_17037);
nor U21982 (N_21982,N_15606,N_16379);
nand U21983 (N_21983,N_16508,N_18278);
and U21984 (N_21984,N_17240,N_15800);
and U21985 (N_21985,N_18968,N_17829);
nor U21986 (N_21986,N_17370,N_18388);
nor U21987 (N_21987,N_18754,N_18174);
or U21988 (N_21988,N_17286,N_15516);
and U21989 (N_21989,N_19815,N_19906);
or U21990 (N_21990,N_16501,N_15746);
nand U21991 (N_21991,N_19426,N_19953);
nand U21992 (N_21992,N_17110,N_19751);
and U21993 (N_21993,N_15955,N_19502);
nand U21994 (N_21994,N_17431,N_17285);
nor U21995 (N_21995,N_18216,N_17047);
xor U21996 (N_21996,N_15008,N_18703);
nand U21997 (N_21997,N_17356,N_18500);
xnor U21998 (N_21998,N_16129,N_17473);
and U21999 (N_21999,N_19849,N_17812);
nand U22000 (N_22000,N_15738,N_16530);
xor U22001 (N_22001,N_18176,N_16209);
and U22002 (N_22002,N_19468,N_18121);
xor U22003 (N_22003,N_16461,N_17185);
nand U22004 (N_22004,N_16746,N_16099);
and U22005 (N_22005,N_19946,N_16921);
nor U22006 (N_22006,N_15435,N_19217);
or U22007 (N_22007,N_17235,N_17780);
or U22008 (N_22008,N_16128,N_15194);
nor U22009 (N_22009,N_16937,N_18328);
and U22010 (N_22010,N_18865,N_17757);
xor U22011 (N_22011,N_19627,N_16586);
nor U22012 (N_22012,N_15499,N_15430);
or U22013 (N_22013,N_17701,N_17639);
nand U22014 (N_22014,N_16761,N_16245);
nor U22015 (N_22015,N_18892,N_15539);
and U22016 (N_22016,N_19812,N_19124);
or U22017 (N_22017,N_16357,N_15196);
xor U22018 (N_22018,N_17933,N_18708);
nand U22019 (N_22019,N_17250,N_19235);
xor U22020 (N_22020,N_15216,N_18970);
xnor U22021 (N_22021,N_15020,N_19132);
nor U22022 (N_22022,N_17454,N_18170);
nor U22023 (N_22023,N_15529,N_17024);
nand U22024 (N_22024,N_18563,N_16252);
nor U22025 (N_22025,N_15567,N_17842);
nor U22026 (N_22026,N_17675,N_16270);
nand U22027 (N_22027,N_19392,N_16244);
or U22028 (N_22028,N_19673,N_18022);
or U22029 (N_22029,N_16294,N_16502);
and U22030 (N_22030,N_19724,N_15082);
xor U22031 (N_22031,N_15750,N_19467);
xnor U22032 (N_22032,N_18239,N_17925);
or U22033 (N_22033,N_16996,N_15209);
or U22034 (N_22034,N_17097,N_17847);
nor U22035 (N_22035,N_15522,N_16691);
nor U22036 (N_22036,N_15416,N_16161);
nand U22037 (N_22037,N_16282,N_15105);
xor U22038 (N_22038,N_16829,N_19116);
nand U22039 (N_22039,N_19282,N_15118);
xnor U22040 (N_22040,N_17787,N_16284);
nor U22041 (N_22041,N_15718,N_15826);
xnor U22042 (N_22042,N_18434,N_16778);
nor U22043 (N_22043,N_18663,N_17533);
xor U22044 (N_22044,N_18314,N_18725);
nand U22045 (N_22045,N_15526,N_15464);
nor U22046 (N_22046,N_16144,N_17774);
and U22047 (N_22047,N_15147,N_15673);
nor U22048 (N_22048,N_16074,N_17673);
xnor U22049 (N_22049,N_17799,N_15885);
nor U22050 (N_22050,N_16662,N_18997);
nand U22051 (N_22051,N_18983,N_15731);
nand U22052 (N_22052,N_18972,N_18026);
nand U22053 (N_22053,N_17093,N_18721);
nor U22054 (N_22054,N_19122,N_16256);
xor U22055 (N_22055,N_16729,N_18209);
or U22056 (N_22056,N_18963,N_15568);
nor U22057 (N_22057,N_15453,N_17819);
and U22058 (N_22058,N_15930,N_19844);
nand U22059 (N_22059,N_19318,N_18460);
and U22060 (N_22060,N_18055,N_17772);
and U22061 (N_22061,N_18762,N_15277);
or U22062 (N_22062,N_18692,N_17880);
nand U22063 (N_22063,N_15280,N_16487);
or U22064 (N_22064,N_18108,N_16955);
nor U22065 (N_22065,N_16095,N_18831);
nor U22066 (N_22066,N_15715,N_17108);
nand U22067 (N_22067,N_19435,N_19238);
nand U22068 (N_22068,N_16555,N_18264);
or U22069 (N_22069,N_19128,N_16066);
and U22070 (N_22070,N_15664,N_15865);
xnor U22071 (N_22071,N_16472,N_15791);
nor U22072 (N_22072,N_15679,N_17474);
nor U22073 (N_22073,N_17516,N_15708);
or U22074 (N_22074,N_19401,N_15992);
and U22075 (N_22075,N_15218,N_18193);
xnor U22076 (N_22076,N_19033,N_17512);
nor U22077 (N_22077,N_19875,N_15774);
nor U22078 (N_22078,N_18512,N_15533);
nand U22079 (N_22079,N_15267,N_15551);
and U22080 (N_22080,N_16383,N_16669);
xor U22081 (N_22081,N_17898,N_19609);
or U22082 (N_22082,N_18694,N_17882);
nor U22083 (N_22083,N_16595,N_15634);
nor U22084 (N_22084,N_16855,N_15062);
nor U22085 (N_22085,N_15722,N_17834);
or U22086 (N_22086,N_19463,N_15610);
xor U22087 (N_22087,N_16507,N_17123);
xor U22088 (N_22088,N_19804,N_15612);
nand U22089 (N_22089,N_17856,N_19010);
and U22090 (N_22090,N_17849,N_16005);
or U22091 (N_22091,N_15171,N_15497);
or U22092 (N_22092,N_17104,N_16807);
nor U22093 (N_22093,N_16286,N_16617);
nor U22094 (N_22094,N_16967,N_19163);
nor U22095 (N_22095,N_17015,N_16500);
or U22096 (N_22096,N_19229,N_16969);
nand U22097 (N_22097,N_17544,N_18319);
xnor U22098 (N_22098,N_17368,N_16185);
xnor U22099 (N_22099,N_18287,N_17692);
or U22100 (N_22100,N_15874,N_17098);
xnor U22101 (N_22101,N_16213,N_15395);
or U22102 (N_22102,N_15669,N_16632);
nor U22103 (N_22103,N_17181,N_18491);
xor U22104 (N_22104,N_18822,N_15315);
xnor U22105 (N_22105,N_17309,N_19516);
nor U22106 (N_22106,N_16176,N_18341);
or U22107 (N_22107,N_17334,N_15825);
nor U22108 (N_22108,N_15887,N_15463);
nor U22109 (N_22109,N_19592,N_17027);
nand U22110 (N_22110,N_17198,N_15899);
and U22111 (N_22111,N_19021,N_18429);
nand U22112 (N_22112,N_19329,N_16703);
nor U22113 (N_22113,N_15796,N_15810);
or U22114 (N_22114,N_17518,N_19877);
xnor U22115 (N_22115,N_19330,N_18959);
and U22116 (N_22116,N_18839,N_15815);
nor U22117 (N_22117,N_17591,N_15574);
or U22118 (N_22118,N_17644,N_19127);
xnor U22119 (N_22119,N_16941,N_18348);
nand U22120 (N_22120,N_17192,N_19731);
xnor U22121 (N_22121,N_19515,N_15878);
nor U22122 (N_22122,N_18439,N_17268);
and U22123 (N_22123,N_17000,N_17444);
nor U22124 (N_22124,N_16177,N_15756);
nor U22125 (N_22125,N_16558,N_17510);
nor U22126 (N_22126,N_19430,N_17077);
nand U22127 (N_22127,N_16226,N_15163);
nor U22128 (N_22128,N_16027,N_17461);
nor U22129 (N_22129,N_19579,N_15704);
nor U22130 (N_22130,N_19613,N_17792);
nor U22131 (N_22131,N_16979,N_15244);
xor U22132 (N_22132,N_18271,N_17410);
nand U22133 (N_22133,N_15031,N_18277);
xor U22134 (N_22134,N_15687,N_18210);
and U22135 (N_22135,N_16344,N_16697);
or U22136 (N_22136,N_18518,N_19486);
nand U22137 (N_22137,N_15256,N_17982);
and U22138 (N_22138,N_16957,N_19232);
or U22139 (N_22139,N_18755,N_16075);
or U22140 (N_22140,N_16822,N_17005);
xor U22141 (N_22141,N_16916,N_19615);
or U22142 (N_22142,N_19327,N_17979);
nand U22143 (N_22143,N_19085,N_19253);
nand U22144 (N_22144,N_18916,N_18487);
and U22145 (N_22145,N_19054,N_19661);
nor U22146 (N_22146,N_19185,N_15943);
xnor U22147 (N_22147,N_15075,N_17580);
nor U22148 (N_22148,N_16155,N_15737);
nor U22149 (N_22149,N_16420,N_15972);
xor U22150 (N_22150,N_15186,N_16463);
and U22151 (N_22151,N_19072,N_16368);
or U22152 (N_22152,N_17325,N_18927);
nor U22153 (N_22153,N_19937,N_16044);
xor U22154 (N_22154,N_15223,N_17196);
and U22155 (N_22155,N_15124,N_18369);
nand U22156 (N_22156,N_19350,N_17401);
nand U22157 (N_22157,N_15820,N_19224);
nand U22158 (N_22158,N_15094,N_19443);
nand U22159 (N_22159,N_19315,N_19403);
nand U22160 (N_22160,N_17202,N_19972);
or U22161 (N_22161,N_19156,N_18954);
or U22162 (N_22162,N_15929,N_18214);
xnor U22163 (N_22163,N_15965,N_16889);
nor U22164 (N_22164,N_18608,N_15685);
and U22165 (N_22165,N_18833,N_17756);
and U22166 (N_22166,N_19469,N_18672);
nor U22167 (N_22167,N_19449,N_18230);
and U22168 (N_22168,N_15983,N_15452);
xnor U22169 (N_22169,N_15973,N_15528);
and U22170 (N_22170,N_18508,N_17199);
or U22171 (N_22171,N_18231,N_18237);
nor U22172 (N_22172,N_18713,N_18157);
nand U22173 (N_22173,N_19659,N_16406);
nand U22174 (N_22174,N_18842,N_19917);
nand U22175 (N_22175,N_18106,N_19019);
or U22176 (N_22176,N_16384,N_15296);
and U22177 (N_22177,N_17427,N_19368);
xnor U22178 (N_22178,N_16124,N_17297);
or U22179 (N_22179,N_17567,N_19151);
and U22180 (N_22180,N_18556,N_18073);
or U22181 (N_22181,N_16774,N_18817);
or U22182 (N_22182,N_17278,N_16460);
nor U22183 (N_22183,N_18394,N_19909);
nand U22184 (N_22184,N_16082,N_18015);
nor U22185 (N_22185,N_18458,N_17901);
or U22186 (N_22186,N_16166,N_15597);
nor U22187 (N_22187,N_17081,N_18184);
nor U22188 (N_22188,N_18850,N_18335);
nor U22189 (N_22189,N_17332,N_15944);
xnor U22190 (N_22190,N_16631,N_17869);
xnor U22191 (N_22191,N_15168,N_19641);
and U22192 (N_22192,N_15166,N_19066);
or U22193 (N_22193,N_18574,N_18913);
or U22194 (N_22194,N_19091,N_19624);
nand U22195 (N_22195,N_19714,N_15496);
nor U22196 (N_22196,N_19996,N_15021);
or U22197 (N_22197,N_19548,N_15202);
and U22198 (N_22198,N_15150,N_17989);
or U22199 (N_22199,N_16151,N_17615);
nor U22200 (N_22200,N_17570,N_18479);
or U22201 (N_22201,N_17316,N_16599);
xnor U22202 (N_22202,N_18196,N_17390);
xnor U22203 (N_22203,N_16167,N_18848);
xnor U22204 (N_22204,N_19509,N_15619);
nand U22205 (N_22205,N_17670,N_16733);
xnor U22206 (N_22206,N_15178,N_15089);
nand U22207 (N_22207,N_18171,N_15248);
nor U22208 (N_22208,N_15571,N_15386);
xnor U22209 (N_22209,N_17961,N_18907);
and U22210 (N_22210,N_15070,N_19179);
or U22211 (N_22211,N_15290,N_17386);
nor U22212 (N_22212,N_17149,N_19640);
and U22213 (N_22213,N_19032,N_18289);
xnor U22214 (N_22214,N_19638,N_15167);
or U22215 (N_22215,N_15250,N_19305);
nor U22216 (N_22216,N_17455,N_19789);
xnor U22217 (N_22217,N_17918,N_16929);
xor U22218 (N_22218,N_17674,N_18553);
and U22219 (N_22219,N_19002,N_15601);
or U22220 (N_22220,N_15258,N_17363);
and U22221 (N_22221,N_15861,N_18855);
xor U22222 (N_22222,N_16056,N_19210);
and U22223 (N_22223,N_16820,N_15064);
xnor U22224 (N_22224,N_16013,N_16096);
xnor U22225 (N_22225,N_15048,N_19531);
or U22226 (N_22226,N_18359,N_15966);
xor U22227 (N_22227,N_17693,N_16794);
and U22228 (N_22228,N_17929,N_18292);
or U22229 (N_22229,N_16026,N_18668);
xor U22230 (N_22230,N_19380,N_16186);
xor U22231 (N_22231,N_18810,N_19149);
nand U22232 (N_22232,N_18194,N_16858);
and U22233 (N_22233,N_16672,N_16315);
or U22234 (N_22234,N_15095,N_18814);
or U22235 (N_22235,N_15678,N_17451);
or U22236 (N_22236,N_16959,N_16238);
xor U22237 (N_22237,N_19338,N_17336);
nor U22238 (N_22238,N_19191,N_19612);
and U22239 (N_22239,N_17974,N_19747);
xnor U22240 (N_22240,N_15187,N_15366);
or U22241 (N_22241,N_19052,N_18768);
nor U22242 (N_22242,N_17700,N_16110);
nand U22243 (N_22243,N_19016,N_16641);
and U22244 (N_22244,N_18982,N_15693);
nor U22245 (N_22245,N_19582,N_18900);
xnor U22246 (N_22246,N_15111,N_17917);
and U22247 (N_22247,N_17092,N_18501);
xnor U22248 (N_22248,N_19004,N_15549);
nor U22249 (N_22249,N_16706,N_19903);
xor U22250 (N_22250,N_16476,N_17863);
and U22251 (N_22251,N_16496,N_17260);
and U22252 (N_22252,N_17055,N_15044);
xor U22253 (N_22253,N_17480,N_18520);
and U22254 (N_22254,N_16231,N_17682);
or U22255 (N_22255,N_18021,N_15068);
and U22256 (N_22256,N_16414,N_19098);
nor U22257 (N_22257,N_19196,N_17763);
or U22258 (N_22258,N_15849,N_17959);
nor U22259 (N_22259,N_19077,N_16323);
nor U22260 (N_22260,N_16652,N_15467);
or U22261 (N_22261,N_18244,N_16232);
nand U22262 (N_22262,N_18224,N_15284);
nand U22263 (N_22263,N_17759,N_19746);
and U22264 (N_22264,N_19690,N_19572);
or U22265 (N_22265,N_19629,N_18165);
or U22266 (N_22266,N_16370,N_17352);
or U22267 (N_22267,N_18018,N_19383);
xnor U22268 (N_22268,N_16982,N_18874);
or U22269 (N_22269,N_17920,N_16179);
xnor U22270 (N_22270,N_16949,N_17049);
or U22271 (N_22271,N_18505,N_15149);
nor U22272 (N_22272,N_18470,N_18824);
nor U22273 (N_22273,N_19556,N_19773);
nand U22274 (N_22274,N_17731,N_18477);
nor U22275 (N_22275,N_18191,N_15061);
nor U22276 (N_22276,N_16984,N_18656);
nor U22277 (N_22277,N_15543,N_19559);
and U22278 (N_22278,N_17638,N_18772);
nor U22279 (N_22279,N_17439,N_16400);
nand U22280 (N_22280,N_16490,N_19351);
or U22281 (N_22281,N_17571,N_16688);
and U22282 (N_22282,N_17134,N_16758);
nand U22283 (N_22283,N_19507,N_19542);
and U22284 (N_22284,N_18096,N_18827);
and U22285 (N_22285,N_17137,N_18468);
nor U22286 (N_22286,N_18248,N_18440);
nand U22287 (N_22287,N_17303,N_15398);
nand U22288 (N_22288,N_17479,N_19045);
xnor U22289 (N_22289,N_17546,N_15122);
and U22290 (N_22290,N_17632,N_15830);
xnor U22291 (N_22291,N_16298,N_17471);
nor U22292 (N_22292,N_17012,N_16682);
nand U22293 (N_22293,N_17248,N_15454);
xor U22294 (N_22294,N_18077,N_19992);
and U22295 (N_22295,N_17306,N_16880);
nor U22296 (N_22296,N_16594,N_15097);
nor U22297 (N_22297,N_18534,N_17640);
nor U22298 (N_22298,N_16388,N_19336);
and U22299 (N_22299,N_19342,N_17833);
xnor U22300 (N_22300,N_19480,N_17691);
or U22301 (N_22301,N_16551,N_19785);
nand U22302 (N_22302,N_18441,N_17997);
and U22303 (N_22303,N_19126,N_16419);
or U22304 (N_22304,N_17333,N_19438);
and U22305 (N_22305,N_17270,N_18976);
or U22306 (N_22306,N_16264,N_16520);
and U22307 (N_22307,N_19645,N_17960);
and U22308 (N_22308,N_18238,N_19482);
xor U22309 (N_22309,N_15860,N_15322);
nand U22310 (N_22310,N_17827,N_15626);
and U22311 (N_22311,N_17481,N_15537);
or U22312 (N_22312,N_17126,N_19194);
or U22313 (N_22313,N_16088,N_15876);
nand U22314 (N_22314,N_16708,N_16975);
and U22315 (N_22315,N_18340,N_16505);
xor U22316 (N_22316,N_16574,N_18489);
and U22317 (N_22317,N_16649,N_18932);
nor U22318 (N_22318,N_16412,N_15092);
xnor U22319 (N_22319,N_16780,N_18877);
nand U22320 (N_22320,N_18638,N_17687);
or U22321 (N_22321,N_16473,N_19993);
nand U22322 (N_22322,N_16288,N_19727);
nor U22323 (N_22323,N_17291,N_16699);
nor U22324 (N_22324,N_16330,N_18382);
or U22325 (N_22325,N_18987,N_16717);
and U22326 (N_22326,N_15375,N_15589);
nand U22327 (N_22327,N_18820,N_19597);
or U22328 (N_22328,N_16255,N_18551);
and U22329 (N_22329,N_19916,N_19765);
or U22330 (N_22330,N_19970,N_16086);
nand U22331 (N_22331,N_18618,N_16050);
and U22332 (N_22332,N_16958,N_19363);
nor U22333 (N_22333,N_18936,N_16173);
nor U22334 (N_22334,N_17698,N_18321);
and U22335 (N_22335,N_16908,N_15381);
nor U22336 (N_22336,N_17614,N_18791);
and U22337 (N_22337,N_15351,N_16071);
and U22338 (N_22338,N_17376,N_15853);
xor U22339 (N_22339,N_15490,N_19312);
and U22340 (N_22340,N_18217,N_19797);
nand U22341 (N_22341,N_19845,N_18660);
xnor U22342 (N_22342,N_15439,N_19276);
xor U22343 (N_22343,N_18544,N_17101);
nand U22344 (N_22344,N_16643,N_18691);
xor U22345 (N_22345,N_15819,N_15059);
xnor U22346 (N_22346,N_19800,N_15152);
nor U22347 (N_22347,N_17588,N_16954);
nor U22348 (N_22348,N_18961,N_19169);
xnor U22349 (N_22349,N_17813,N_19752);
nand U22350 (N_22350,N_19654,N_18027);
xnor U22351 (N_22351,N_16350,N_17485);
and U22352 (N_22352,N_17168,N_19436);
nand U22353 (N_22353,N_17164,N_19657);
nand U22354 (N_22354,N_18172,N_17289);
or U22355 (N_22355,N_16131,N_19658);
nand U22356 (N_22356,N_17273,N_17721);
or U22357 (N_22357,N_18889,N_16782);
or U22358 (N_22358,N_15207,N_18234);
and U22359 (N_22359,N_16601,N_18763);
nand U22360 (N_22360,N_17450,N_15557);
or U22361 (N_22361,N_15131,N_15788);
and U22362 (N_22362,N_15749,N_19712);
and U22363 (N_22363,N_15429,N_15636);
or U22364 (N_22364,N_18795,N_15069);
xor U22365 (N_22365,N_15141,N_19088);
nand U22366 (N_22366,N_16150,N_19729);
and U22367 (N_22367,N_18058,N_15793);
xnor U22368 (N_22368,N_18393,N_19028);
or U22369 (N_22369,N_18749,N_17660);
nand U22370 (N_22370,N_18863,N_18805);
nor U22371 (N_22371,N_16839,N_17233);
or U22372 (N_22372,N_19263,N_19899);
or U22373 (N_22373,N_16539,N_18924);
or U22374 (N_22374,N_19986,N_19001);
nand U22375 (N_22375,N_15591,N_19810);
and U22376 (N_22376,N_19695,N_16006);
or U22377 (N_22377,N_17404,N_17835);
or U22378 (N_22378,N_17252,N_16709);
xnor U22379 (N_22379,N_16537,N_15109);
and U22380 (N_22380,N_18840,N_18923);
or U22381 (N_22381,N_16127,N_16671);
nor U22382 (N_22382,N_17996,N_17998);
or U22383 (N_22383,N_19367,N_17843);
nor U22384 (N_22384,N_19664,N_17215);
or U22385 (N_22385,N_19514,N_16358);
xnor U22386 (N_22386,N_16289,N_15140);
or U22387 (N_22387,N_19117,N_19340);
and U22388 (N_22388,N_16768,N_17854);
nor U22389 (N_22389,N_16544,N_15449);
or U22390 (N_22390,N_16536,N_16582);
nand U22391 (N_22391,N_16181,N_18354);
nor U22392 (N_22392,N_19643,N_17416);
or U22393 (N_22393,N_17540,N_17577);
and U22394 (N_22394,N_15030,N_18347);
and U22395 (N_22395,N_16857,N_16007);
nor U22396 (N_22396,N_17713,N_16748);
nor U22397 (N_22397,N_19133,N_16482);
nand U22398 (N_22398,N_17173,N_15799);
or U22399 (N_22399,N_19386,N_17293);
xnor U22400 (N_22400,N_16451,N_17620);
and U22401 (N_22401,N_18808,N_16630);
nand U22402 (N_22402,N_18744,N_15136);
nand U22403 (N_22403,N_18296,N_17662);
and U22404 (N_22404,N_15010,N_17343);
nand U22405 (N_22405,N_16188,N_17500);
nor U22406 (N_22406,N_18457,N_17764);
nand U22407 (N_22407,N_18135,N_16795);
or U22408 (N_22408,N_19026,N_18462);
xor U22409 (N_22409,N_17030,N_19425);
or U22410 (N_22410,N_18933,N_18517);
or U22411 (N_22411,N_15629,N_17730);
and U22412 (N_22412,N_17521,N_16804);
nand U22413 (N_22413,N_16042,N_17690);
nor U22414 (N_22414,N_19578,N_15103);
xor U22415 (N_22415,N_18960,N_19234);
and U22416 (N_22416,N_17425,N_17265);
and U22417 (N_22417,N_17205,N_16021);
or U22418 (N_22418,N_19736,N_17266);
and U22419 (N_22419,N_15299,N_16991);
nand U22420 (N_22420,N_17955,N_16454);
and U22421 (N_22421,N_16604,N_19525);
nand U22422 (N_22422,N_15378,N_19043);
nor U22423 (N_22423,N_18283,N_18436);
and U22424 (N_22424,N_16133,N_16972);
nand U22425 (N_22425,N_16681,N_17678);
xnor U22426 (N_22426,N_19397,N_19853);
nor U22427 (N_22427,N_17063,N_15883);
nor U22428 (N_22428,N_16239,N_17353);
nor U22429 (N_22429,N_16917,N_18036);
nand U22430 (N_22430,N_16285,N_18769);
nor U22431 (N_22431,N_19106,N_16524);
or U22432 (N_22432,N_17709,N_16760);
or U22433 (N_22433,N_15397,N_17609);
nor U22434 (N_22434,N_19062,N_16948);
or U22435 (N_22435,N_15380,N_15428);
nand U22436 (N_22436,N_19791,N_18249);
nor U22437 (N_22437,N_15614,N_19160);
nand U22438 (N_22438,N_17683,N_15053);
nand U22439 (N_22439,N_17748,N_18905);
or U22440 (N_22440,N_18624,N_17797);
or U22441 (N_22441,N_15868,N_15803);
xnor U22442 (N_22442,N_19824,N_19760);
or U22443 (N_22443,N_17132,N_19718);
or U22444 (N_22444,N_19241,N_17071);
nand U22445 (N_22445,N_18402,N_17080);
nand U22446 (N_22446,N_18400,N_19252);
nand U22447 (N_22447,N_16154,N_18383);
or U22448 (N_22448,N_17399,N_15241);
xnor U22449 (N_22449,N_15762,N_18793);
and U22450 (N_22450,N_18076,N_18000);
or U22451 (N_22451,N_19099,N_15921);
and U22452 (N_22452,N_16462,N_19554);
nand U22453 (N_22453,N_18306,N_16457);
or U22454 (N_22454,N_19745,N_16832);
xnor U22455 (N_22455,N_16263,N_16660);
xor U22456 (N_22456,N_19743,N_19145);
and U22457 (N_22457,N_19092,N_18519);
and U22458 (N_22458,N_18290,N_15777);
nand U22459 (N_22459,N_16787,N_16919);
nor U22460 (N_22460,N_17860,N_17579);
or U22461 (N_22461,N_19598,N_17256);
xnor U22462 (N_22462,N_19626,N_15559);
nand U22463 (N_22463,N_19563,N_17224);
nor U22464 (N_22464,N_16261,N_18533);
xnor U22465 (N_22465,N_16830,N_18481);
or U22466 (N_22466,N_18799,N_16227);
or U22467 (N_22467,N_18722,N_16220);
or U22468 (N_22468,N_17537,N_18612);
xor U22469 (N_22469,N_17900,N_18857);
or U22470 (N_22470,N_16966,N_17909);
nand U22471 (N_22471,N_19209,N_16208);
and U22472 (N_22472,N_16162,N_19219);
or U22473 (N_22473,N_16663,N_17477);
or U22474 (N_22474,N_15361,N_16861);
nand U22475 (N_22475,N_15635,N_19901);
nor U22476 (N_22476,N_19423,N_15713);
or U22477 (N_22477,N_19834,N_17802);
nand U22478 (N_22478,N_15188,N_16516);
nand U22479 (N_22479,N_18601,N_17867);
and U22480 (N_22480,N_15349,N_18368);
and U22481 (N_22481,N_17010,N_16243);
and U22482 (N_22482,N_18811,N_15521);
nand U22483 (N_22483,N_18072,N_19590);
or U22484 (N_22484,N_18338,N_15121);
and U22485 (N_22485,N_16034,N_17218);
nor U22486 (N_22486,N_16334,N_17414);
and U22487 (N_22487,N_19566,N_15415);
and U22488 (N_22488,N_17062,N_17924);
or U22489 (N_22489,N_18636,N_15605);
and U22490 (N_22490,N_15886,N_16480);
or U22491 (N_22491,N_15651,N_16541);
and U22492 (N_22492,N_19574,N_15205);
and U22493 (N_22493,N_19604,N_19022);
xor U22494 (N_22494,N_18742,N_18614);
nor U22495 (N_22495,N_16798,N_16332);
or U22496 (N_22496,N_18069,N_16685);
nand U22497 (N_22497,N_19669,N_17679);
and U22498 (N_22498,N_16354,N_19231);
or U22499 (N_22499,N_16258,N_17213);
xor U22500 (N_22500,N_17416,N_17900);
nor U22501 (N_22501,N_19692,N_17337);
xor U22502 (N_22502,N_15931,N_16954);
nor U22503 (N_22503,N_16587,N_19006);
xnor U22504 (N_22504,N_19850,N_16351);
nand U22505 (N_22505,N_18959,N_17663);
and U22506 (N_22506,N_15856,N_16810);
and U22507 (N_22507,N_17693,N_19316);
xor U22508 (N_22508,N_17026,N_19397);
nor U22509 (N_22509,N_17645,N_15133);
xor U22510 (N_22510,N_17387,N_17989);
and U22511 (N_22511,N_19514,N_17627);
and U22512 (N_22512,N_15221,N_16224);
nand U22513 (N_22513,N_17330,N_19312);
xor U22514 (N_22514,N_18242,N_18876);
nand U22515 (N_22515,N_15394,N_17520);
nand U22516 (N_22516,N_15015,N_18306);
and U22517 (N_22517,N_16913,N_19261);
and U22518 (N_22518,N_18547,N_18553);
nor U22519 (N_22519,N_16969,N_19955);
nor U22520 (N_22520,N_19028,N_19577);
nand U22521 (N_22521,N_16847,N_16381);
xor U22522 (N_22522,N_18072,N_18603);
xnor U22523 (N_22523,N_17919,N_16772);
nor U22524 (N_22524,N_15217,N_17402);
xnor U22525 (N_22525,N_16558,N_15405);
nand U22526 (N_22526,N_16949,N_17879);
nand U22527 (N_22527,N_17175,N_15789);
or U22528 (N_22528,N_16413,N_18676);
or U22529 (N_22529,N_15585,N_18934);
nand U22530 (N_22530,N_15623,N_15826);
and U22531 (N_22531,N_18325,N_19816);
and U22532 (N_22532,N_15752,N_19022);
and U22533 (N_22533,N_17636,N_17523);
nand U22534 (N_22534,N_19914,N_17904);
xor U22535 (N_22535,N_16202,N_19163);
nand U22536 (N_22536,N_17213,N_19292);
and U22537 (N_22537,N_19129,N_15755);
nor U22538 (N_22538,N_15183,N_18465);
nor U22539 (N_22539,N_16029,N_18383);
nor U22540 (N_22540,N_15965,N_19200);
nand U22541 (N_22541,N_17782,N_15671);
and U22542 (N_22542,N_18046,N_18025);
or U22543 (N_22543,N_16370,N_16606);
or U22544 (N_22544,N_15272,N_18250);
and U22545 (N_22545,N_16413,N_16748);
nor U22546 (N_22546,N_18483,N_19763);
xor U22547 (N_22547,N_15921,N_19557);
xor U22548 (N_22548,N_16985,N_16997);
and U22549 (N_22549,N_17981,N_19370);
nand U22550 (N_22550,N_16852,N_18135);
and U22551 (N_22551,N_17050,N_16064);
or U22552 (N_22552,N_19712,N_17517);
nand U22553 (N_22553,N_19815,N_19912);
xor U22554 (N_22554,N_16027,N_16592);
and U22555 (N_22555,N_17657,N_19138);
nor U22556 (N_22556,N_15815,N_19261);
and U22557 (N_22557,N_18342,N_17090);
nand U22558 (N_22558,N_19395,N_16150);
nand U22559 (N_22559,N_17203,N_15100);
nand U22560 (N_22560,N_18187,N_19397);
nand U22561 (N_22561,N_18957,N_17474);
nand U22562 (N_22562,N_19559,N_17428);
nor U22563 (N_22563,N_18811,N_18946);
xnor U22564 (N_22564,N_15927,N_16486);
and U22565 (N_22565,N_17494,N_16190);
and U22566 (N_22566,N_16014,N_17449);
nor U22567 (N_22567,N_18453,N_18621);
and U22568 (N_22568,N_19281,N_18908);
or U22569 (N_22569,N_16505,N_18745);
or U22570 (N_22570,N_19074,N_18094);
xor U22571 (N_22571,N_17860,N_15812);
or U22572 (N_22572,N_15301,N_19853);
nor U22573 (N_22573,N_18525,N_18825);
and U22574 (N_22574,N_19457,N_15619);
nor U22575 (N_22575,N_18029,N_15397);
and U22576 (N_22576,N_17149,N_17575);
nor U22577 (N_22577,N_18764,N_16366);
nor U22578 (N_22578,N_15889,N_15459);
and U22579 (N_22579,N_19999,N_18588);
or U22580 (N_22580,N_19217,N_16171);
and U22581 (N_22581,N_16887,N_19723);
nor U22582 (N_22582,N_17819,N_15188);
nor U22583 (N_22583,N_17346,N_17334);
or U22584 (N_22584,N_16180,N_18581);
xor U22585 (N_22585,N_17634,N_17940);
nand U22586 (N_22586,N_17053,N_18399);
nand U22587 (N_22587,N_15065,N_16662);
nor U22588 (N_22588,N_18392,N_16929);
nand U22589 (N_22589,N_16272,N_18097);
and U22590 (N_22590,N_15701,N_16936);
nor U22591 (N_22591,N_19919,N_17392);
and U22592 (N_22592,N_18911,N_17879);
or U22593 (N_22593,N_16181,N_18101);
and U22594 (N_22594,N_17740,N_15033);
and U22595 (N_22595,N_16318,N_19275);
nand U22596 (N_22596,N_17153,N_19886);
nor U22597 (N_22597,N_19720,N_15643);
nand U22598 (N_22598,N_17088,N_17592);
nand U22599 (N_22599,N_15346,N_15073);
nand U22600 (N_22600,N_19646,N_15801);
and U22601 (N_22601,N_16645,N_19691);
xor U22602 (N_22602,N_16540,N_18359);
nand U22603 (N_22603,N_17462,N_17971);
or U22604 (N_22604,N_19133,N_17208);
nand U22605 (N_22605,N_18351,N_16474);
and U22606 (N_22606,N_18762,N_18022);
and U22607 (N_22607,N_17422,N_19948);
and U22608 (N_22608,N_16839,N_15286);
and U22609 (N_22609,N_18182,N_16354);
and U22610 (N_22610,N_18275,N_17332);
and U22611 (N_22611,N_19940,N_15199);
xnor U22612 (N_22612,N_19341,N_15755);
and U22613 (N_22613,N_18376,N_19778);
xnor U22614 (N_22614,N_15799,N_15069);
nand U22615 (N_22615,N_15679,N_15105);
nor U22616 (N_22616,N_16228,N_17520);
nand U22617 (N_22617,N_15639,N_18481);
and U22618 (N_22618,N_16990,N_18873);
nand U22619 (N_22619,N_15737,N_18914);
and U22620 (N_22620,N_15665,N_15207);
and U22621 (N_22621,N_19962,N_16145);
nand U22622 (N_22622,N_16307,N_16062);
nor U22623 (N_22623,N_19696,N_19718);
xnor U22624 (N_22624,N_17320,N_15636);
or U22625 (N_22625,N_16300,N_15118);
nand U22626 (N_22626,N_16488,N_16704);
xnor U22627 (N_22627,N_15714,N_17853);
xor U22628 (N_22628,N_15317,N_16001);
xor U22629 (N_22629,N_18847,N_16802);
nor U22630 (N_22630,N_18805,N_19423);
or U22631 (N_22631,N_17361,N_15931);
xnor U22632 (N_22632,N_18658,N_16449);
nor U22633 (N_22633,N_16214,N_19065);
xor U22634 (N_22634,N_19005,N_18541);
nor U22635 (N_22635,N_17422,N_18855);
nor U22636 (N_22636,N_15960,N_15554);
or U22637 (N_22637,N_15239,N_16426);
nor U22638 (N_22638,N_16200,N_19968);
xnor U22639 (N_22639,N_15969,N_15127);
and U22640 (N_22640,N_17651,N_15929);
nor U22641 (N_22641,N_15571,N_16005);
nor U22642 (N_22642,N_16406,N_15761);
and U22643 (N_22643,N_15146,N_19741);
and U22644 (N_22644,N_18166,N_15442);
xor U22645 (N_22645,N_18909,N_17257);
xnor U22646 (N_22646,N_17361,N_19156);
or U22647 (N_22647,N_15204,N_16528);
nand U22648 (N_22648,N_16727,N_19326);
or U22649 (N_22649,N_19264,N_16637);
nor U22650 (N_22650,N_15678,N_15114);
and U22651 (N_22651,N_17325,N_18750);
and U22652 (N_22652,N_19952,N_19226);
nor U22653 (N_22653,N_19338,N_15027);
or U22654 (N_22654,N_17099,N_16257);
nor U22655 (N_22655,N_15112,N_15332);
nand U22656 (N_22656,N_17937,N_17585);
xor U22657 (N_22657,N_15972,N_16922);
nand U22658 (N_22658,N_16800,N_15136);
or U22659 (N_22659,N_19499,N_19163);
and U22660 (N_22660,N_19269,N_16332);
or U22661 (N_22661,N_18249,N_15600);
or U22662 (N_22662,N_19027,N_16519);
and U22663 (N_22663,N_19249,N_19992);
nand U22664 (N_22664,N_16355,N_17198);
or U22665 (N_22665,N_18806,N_17090);
nor U22666 (N_22666,N_17591,N_17721);
or U22667 (N_22667,N_16768,N_19144);
xor U22668 (N_22668,N_15310,N_17886);
and U22669 (N_22669,N_15411,N_15232);
or U22670 (N_22670,N_17302,N_17309);
nand U22671 (N_22671,N_17696,N_17006);
and U22672 (N_22672,N_17314,N_19041);
or U22673 (N_22673,N_16377,N_16119);
or U22674 (N_22674,N_18372,N_19094);
or U22675 (N_22675,N_18367,N_15421);
and U22676 (N_22676,N_19100,N_18707);
or U22677 (N_22677,N_17984,N_18074);
nand U22678 (N_22678,N_17907,N_16032);
nor U22679 (N_22679,N_18979,N_15915);
xnor U22680 (N_22680,N_16551,N_19665);
and U22681 (N_22681,N_19342,N_17991);
nor U22682 (N_22682,N_19661,N_18751);
and U22683 (N_22683,N_18781,N_19666);
xor U22684 (N_22684,N_17675,N_16944);
nand U22685 (N_22685,N_16489,N_18192);
xnor U22686 (N_22686,N_18003,N_18194);
nor U22687 (N_22687,N_17172,N_16326);
xnor U22688 (N_22688,N_17227,N_15518);
and U22689 (N_22689,N_15607,N_18497);
and U22690 (N_22690,N_18626,N_18910);
or U22691 (N_22691,N_17118,N_19739);
nand U22692 (N_22692,N_18454,N_18251);
nor U22693 (N_22693,N_15972,N_15031);
nor U22694 (N_22694,N_15311,N_15791);
xnor U22695 (N_22695,N_16023,N_17257);
nand U22696 (N_22696,N_15085,N_16470);
nand U22697 (N_22697,N_17901,N_18676);
xnor U22698 (N_22698,N_17683,N_17681);
nor U22699 (N_22699,N_18170,N_17017);
xnor U22700 (N_22700,N_17579,N_19299);
nor U22701 (N_22701,N_18553,N_16598);
and U22702 (N_22702,N_18051,N_16590);
xor U22703 (N_22703,N_19835,N_15195);
nor U22704 (N_22704,N_18839,N_19287);
or U22705 (N_22705,N_17211,N_15845);
and U22706 (N_22706,N_15626,N_17308);
and U22707 (N_22707,N_17170,N_19502);
or U22708 (N_22708,N_18957,N_15550);
nand U22709 (N_22709,N_19531,N_19582);
and U22710 (N_22710,N_16627,N_16348);
nor U22711 (N_22711,N_16772,N_17327);
nor U22712 (N_22712,N_15457,N_16867);
nor U22713 (N_22713,N_18687,N_18702);
xnor U22714 (N_22714,N_16714,N_17656);
nand U22715 (N_22715,N_17284,N_16168);
nand U22716 (N_22716,N_16342,N_19672);
nor U22717 (N_22717,N_18345,N_19513);
or U22718 (N_22718,N_16061,N_18667);
nand U22719 (N_22719,N_16390,N_17853);
and U22720 (N_22720,N_16329,N_17357);
nor U22721 (N_22721,N_15022,N_17357);
and U22722 (N_22722,N_17499,N_16753);
and U22723 (N_22723,N_15723,N_18636);
nand U22724 (N_22724,N_19281,N_16982);
or U22725 (N_22725,N_17189,N_18780);
and U22726 (N_22726,N_16833,N_15442);
nand U22727 (N_22727,N_18858,N_17976);
xor U22728 (N_22728,N_15686,N_15867);
or U22729 (N_22729,N_15923,N_16455);
nand U22730 (N_22730,N_15908,N_17546);
or U22731 (N_22731,N_18737,N_16319);
nor U22732 (N_22732,N_18097,N_15684);
and U22733 (N_22733,N_18805,N_19592);
nor U22734 (N_22734,N_16479,N_17981);
or U22735 (N_22735,N_17898,N_15414);
xor U22736 (N_22736,N_19355,N_15551);
xnor U22737 (N_22737,N_17759,N_16176);
xnor U22738 (N_22738,N_16484,N_15381);
xnor U22739 (N_22739,N_15758,N_19205);
xor U22740 (N_22740,N_19984,N_15241);
nand U22741 (N_22741,N_19202,N_19249);
and U22742 (N_22742,N_16375,N_15238);
and U22743 (N_22743,N_17155,N_17978);
xor U22744 (N_22744,N_16165,N_15071);
xor U22745 (N_22745,N_17630,N_17066);
and U22746 (N_22746,N_15452,N_17589);
or U22747 (N_22747,N_15991,N_16818);
nand U22748 (N_22748,N_16919,N_19982);
or U22749 (N_22749,N_15744,N_16200);
or U22750 (N_22750,N_16467,N_16536);
and U22751 (N_22751,N_19736,N_19328);
xnor U22752 (N_22752,N_18451,N_16341);
and U22753 (N_22753,N_19729,N_19565);
or U22754 (N_22754,N_16475,N_18998);
nor U22755 (N_22755,N_19496,N_17402);
xnor U22756 (N_22756,N_18487,N_18052);
xor U22757 (N_22757,N_15693,N_17215);
nor U22758 (N_22758,N_17709,N_19066);
or U22759 (N_22759,N_18185,N_18058);
or U22760 (N_22760,N_19050,N_17908);
xor U22761 (N_22761,N_16205,N_18764);
nand U22762 (N_22762,N_18124,N_17709);
and U22763 (N_22763,N_18710,N_19603);
or U22764 (N_22764,N_15766,N_17065);
and U22765 (N_22765,N_17655,N_16327);
nand U22766 (N_22766,N_16714,N_15907);
xor U22767 (N_22767,N_17522,N_18962);
or U22768 (N_22768,N_16565,N_19846);
and U22769 (N_22769,N_17678,N_18550);
nand U22770 (N_22770,N_19578,N_16870);
and U22771 (N_22771,N_16996,N_15307);
nand U22772 (N_22772,N_17211,N_18071);
and U22773 (N_22773,N_19835,N_19834);
xor U22774 (N_22774,N_19323,N_19124);
xnor U22775 (N_22775,N_15973,N_19444);
and U22776 (N_22776,N_15753,N_18067);
nor U22777 (N_22777,N_15099,N_15008);
or U22778 (N_22778,N_15347,N_18569);
nand U22779 (N_22779,N_18768,N_18795);
xnor U22780 (N_22780,N_19224,N_17583);
xnor U22781 (N_22781,N_16201,N_17571);
nand U22782 (N_22782,N_15311,N_18534);
xnor U22783 (N_22783,N_17840,N_16219);
xnor U22784 (N_22784,N_16667,N_17195);
xor U22785 (N_22785,N_18044,N_18380);
xnor U22786 (N_22786,N_17204,N_19343);
and U22787 (N_22787,N_16413,N_16585);
nand U22788 (N_22788,N_18344,N_16524);
or U22789 (N_22789,N_19219,N_19845);
and U22790 (N_22790,N_16855,N_16040);
nor U22791 (N_22791,N_15784,N_18690);
nand U22792 (N_22792,N_16422,N_19879);
nor U22793 (N_22793,N_19180,N_19604);
and U22794 (N_22794,N_16950,N_18060);
nand U22795 (N_22795,N_17332,N_18641);
nor U22796 (N_22796,N_18834,N_15590);
xnor U22797 (N_22797,N_17731,N_19930);
and U22798 (N_22798,N_18907,N_18955);
nand U22799 (N_22799,N_16942,N_17816);
or U22800 (N_22800,N_19192,N_18597);
or U22801 (N_22801,N_18794,N_15497);
or U22802 (N_22802,N_19756,N_16644);
xnor U22803 (N_22803,N_17287,N_18544);
or U22804 (N_22804,N_16611,N_17768);
nor U22805 (N_22805,N_17475,N_19287);
xor U22806 (N_22806,N_18427,N_17448);
xor U22807 (N_22807,N_15390,N_18598);
or U22808 (N_22808,N_19384,N_19645);
nand U22809 (N_22809,N_16128,N_18504);
nor U22810 (N_22810,N_18691,N_15579);
and U22811 (N_22811,N_18394,N_17297);
and U22812 (N_22812,N_16850,N_19827);
and U22813 (N_22813,N_16036,N_19222);
or U22814 (N_22814,N_17831,N_16809);
xor U22815 (N_22815,N_18641,N_16135);
xnor U22816 (N_22816,N_18601,N_15861);
nand U22817 (N_22817,N_18280,N_19826);
nor U22818 (N_22818,N_16059,N_17796);
xor U22819 (N_22819,N_18190,N_17446);
nor U22820 (N_22820,N_18811,N_15199);
or U22821 (N_22821,N_19256,N_17997);
or U22822 (N_22822,N_17166,N_15138);
nand U22823 (N_22823,N_16864,N_19397);
nor U22824 (N_22824,N_19586,N_15009);
or U22825 (N_22825,N_17696,N_18725);
nand U22826 (N_22826,N_17637,N_18390);
and U22827 (N_22827,N_17797,N_19180);
xnor U22828 (N_22828,N_15224,N_16711);
xnor U22829 (N_22829,N_18359,N_15063);
xor U22830 (N_22830,N_19901,N_17151);
nand U22831 (N_22831,N_17084,N_17678);
xor U22832 (N_22832,N_19600,N_19278);
and U22833 (N_22833,N_17391,N_17482);
nor U22834 (N_22834,N_19997,N_19062);
nor U22835 (N_22835,N_16865,N_19710);
nand U22836 (N_22836,N_19535,N_15038);
or U22837 (N_22837,N_18598,N_18763);
nand U22838 (N_22838,N_15048,N_18644);
nor U22839 (N_22839,N_16297,N_15289);
nand U22840 (N_22840,N_18692,N_15848);
nand U22841 (N_22841,N_19757,N_18630);
and U22842 (N_22842,N_19499,N_17932);
nand U22843 (N_22843,N_18482,N_16422);
nor U22844 (N_22844,N_15103,N_15593);
nand U22845 (N_22845,N_16832,N_18492);
or U22846 (N_22846,N_15973,N_18136);
nor U22847 (N_22847,N_18578,N_16568);
nor U22848 (N_22848,N_19925,N_17539);
or U22849 (N_22849,N_18742,N_18892);
and U22850 (N_22850,N_19752,N_19817);
nand U22851 (N_22851,N_17490,N_19932);
nand U22852 (N_22852,N_16474,N_19909);
and U22853 (N_22853,N_19470,N_16249);
or U22854 (N_22854,N_17585,N_18704);
nand U22855 (N_22855,N_17741,N_15214);
xor U22856 (N_22856,N_19152,N_19245);
xnor U22857 (N_22857,N_19115,N_18682);
and U22858 (N_22858,N_15668,N_18559);
or U22859 (N_22859,N_19704,N_17157);
or U22860 (N_22860,N_16081,N_15602);
nand U22861 (N_22861,N_17715,N_19287);
or U22862 (N_22862,N_16354,N_16976);
xor U22863 (N_22863,N_19270,N_17419);
or U22864 (N_22864,N_18251,N_19114);
and U22865 (N_22865,N_16061,N_18063);
nand U22866 (N_22866,N_16294,N_15270);
nor U22867 (N_22867,N_18028,N_17266);
xor U22868 (N_22868,N_18024,N_16053);
and U22869 (N_22869,N_15304,N_15776);
and U22870 (N_22870,N_17738,N_17105);
nor U22871 (N_22871,N_17740,N_16448);
and U22872 (N_22872,N_18090,N_16665);
nand U22873 (N_22873,N_19927,N_16948);
xor U22874 (N_22874,N_15928,N_19595);
nand U22875 (N_22875,N_19130,N_17289);
nand U22876 (N_22876,N_19873,N_19895);
nand U22877 (N_22877,N_16740,N_18820);
and U22878 (N_22878,N_17571,N_19751);
or U22879 (N_22879,N_19702,N_15277);
xor U22880 (N_22880,N_18076,N_18094);
nand U22881 (N_22881,N_19091,N_18799);
nand U22882 (N_22882,N_15649,N_15070);
nand U22883 (N_22883,N_16329,N_15945);
nand U22884 (N_22884,N_15015,N_19124);
or U22885 (N_22885,N_19809,N_18781);
xnor U22886 (N_22886,N_16877,N_16543);
nor U22887 (N_22887,N_17376,N_16405);
nor U22888 (N_22888,N_17885,N_19252);
xnor U22889 (N_22889,N_18474,N_17988);
xor U22890 (N_22890,N_18581,N_15764);
or U22891 (N_22891,N_19309,N_19269);
or U22892 (N_22892,N_17108,N_17038);
and U22893 (N_22893,N_17263,N_17503);
or U22894 (N_22894,N_15004,N_19897);
and U22895 (N_22895,N_19695,N_18994);
xnor U22896 (N_22896,N_16280,N_16564);
xnor U22897 (N_22897,N_16719,N_19022);
and U22898 (N_22898,N_17863,N_19817);
xnor U22899 (N_22899,N_18920,N_17804);
xnor U22900 (N_22900,N_16859,N_18464);
or U22901 (N_22901,N_19693,N_19991);
nor U22902 (N_22902,N_16713,N_18874);
and U22903 (N_22903,N_15063,N_17890);
nor U22904 (N_22904,N_19630,N_17677);
or U22905 (N_22905,N_15856,N_19020);
xor U22906 (N_22906,N_16393,N_19258);
nand U22907 (N_22907,N_15033,N_16315);
nor U22908 (N_22908,N_15205,N_19040);
and U22909 (N_22909,N_18151,N_16313);
or U22910 (N_22910,N_17317,N_18306);
nor U22911 (N_22911,N_15740,N_16358);
and U22912 (N_22912,N_15175,N_17989);
xnor U22913 (N_22913,N_17332,N_17412);
nor U22914 (N_22914,N_15521,N_18774);
xnor U22915 (N_22915,N_17536,N_19870);
xor U22916 (N_22916,N_17732,N_15667);
nand U22917 (N_22917,N_17123,N_18332);
and U22918 (N_22918,N_16107,N_18954);
and U22919 (N_22919,N_17589,N_15514);
and U22920 (N_22920,N_15524,N_17503);
or U22921 (N_22921,N_16208,N_19472);
nand U22922 (N_22922,N_16590,N_18157);
nand U22923 (N_22923,N_19024,N_19250);
xor U22924 (N_22924,N_16113,N_16862);
nor U22925 (N_22925,N_16864,N_15273);
and U22926 (N_22926,N_15622,N_16728);
nand U22927 (N_22927,N_15999,N_15543);
nand U22928 (N_22928,N_15412,N_19064);
nand U22929 (N_22929,N_15641,N_18784);
nor U22930 (N_22930,N_18353,N_16619);
and U22931 (N_22931,N_16538,N_17093);
nand U22932 (N_22932,N_19877,N_18268);
nor U22933 (N_22933,N_19729,N_15166);
xnor U22934 (N_22934,N_17958,N_19835);
xor U22935 (N_22935,N_17469,N_16300);
and U22936 (N_22936,N_19668,N_15103);
or U22937 (N_22937,N_16336,N_18344);
and U22938 (N_22938,N_16074,N_15403);
nor U22939 (N_22939,N_16471,N_16422);
nor U22940 (N_22940,N_18855,N_16513);
nand U22941 (N_22941,N_19943,N_15459);
xor U22942 (N_22942,N_18662,N_18293);
nor U22943 (N_22943,N_17954,N_19392);
nor U22944 (N_22944,N_19205,N_19133);
or U22945 (N_22945,N_17642,N_17522);
xor U22946 (N_22946,N_18473,N_16195);
or U22947 (N_22947,N_19579,N_19575);
nor U22948 (N_22948,N_18331,N_16991);
xnor U22949 (N_22949,N_16758,N_15623);
and U22950 (N_22950,N_16405,N_15678);
and U22951 (N_22951,N_16118,N_16300);
xor U22952 (N_22952,N_19282,N_15500);
nand U22953 (N_22953,N_16332,N_16710);
and U22954 (N_22954,N_17390,N_15013);
or U22955 (N_22955,N_18415,N_15902);
nor U22956 (N_22956,N_16776,N_17466);
nor U22957 (N_22957,N_15979,N_16580);
and U22958 (N_22958,N_18289,N_17035);
nand U22959 (N_22959,N_16766,N_16339);
nor U22960 (N_22960,N_19869,N_15024);
and U22961 (N_22961,N_17452,N_16240);
xnor U22962 (N_22962,N_17032,N_15581);
nand U22963 (N_22963,N_15937,N_15697);
xor U22964 (N_22964,N_17924,N_16967);
nand U22965 (N_22965,N_19954,N_19596);
nand U22966 (N_22966,N_18528,N_17139);
nor U22967 (N_22967,N_17583,N_19575);
nor U22968 (N_22968,N_18688,N_18338);
nor U22969 (N_22969,N_18767,N_18106);
or U22970 (N_22970,N_18513,N_18796);
nor U22971 (N_22971,N_19629,N_17782);
nand U22972 (N_22972,N_17860,N_16060);
and U22973 (N_22973,N_15502,N_15001);
and U22974 (N_22974,N_16611,N_18042);
and U22975 (N_22975,N_16380,N_15601);
or U22976 (N_22976,N_19258,N_17386);
xor U22977 (N_22977,N_15434,N_18561);
nor U22978 (N_22978,N_16534,N_18534);
nor U22979 (N_22979,N_15868,N_15248);
or U22980 (N_22980,N_15667,N_15999);
nand U22981 (N_22981,N_15037,N_15772);
nand U22982 (N_22982,N_18619,N_18052);
and U22983 (N_22983,N_16611,N_15960);
or U22984 (N_22984,N_16425,N_17198);
nor U22985 (N_22985,N_15353,N_16685);
xnor U22986 (N_22986,N_17778,N_16668);
nor U22987 (N_22987,N_16167,N_16541);
and U22988 (N_22988,N_19331,N_16856);
nor U22989 (N_22989,N_15605,N_19157);
xor U22990 (N_22990,N_17827,N_19955);
nor U22991 (N_22991,N_15869,N_15527);
nand U22992 (N_22992,N_19891,N_16936);
or U22993 (N_22993,N_16021,N_19890);
or U22994 (N_22994,N_16240,N_17939);
nor U22995 (N_22995,N_15068,N_17001);
and U22996 (N_22996,N_19850,N_16483);
nand U22997 (N_22997,N_16800,N_19418);
or U22998 (N_22998,N_18622,N_15150);
nand U22999 (N_22999,N_16622,N_17703);
or U23000 (N_23000,N_18304,N_19976);
xnor U23001 (N_23001,N_17254,N_17381);
or U23002 (N_23002,N_15460,N_18199);
or U23003 (N_23003,N_15070,N_17991);
nand U23004 (N_23004,N_18436,N_17344);
nor U23005 (N_23005,N_18609,N_17016);
nor U23006 (N_23006,N_18794,N_19574);
nand U23007 (N_23007,N_15970,N_19777);
or U23008 (N_23008,N_16103,N_16968);
nor U23009 (N_23009,N_15624,N_16803);
nand U23010 (N_23010,N_19755,N_18635);
nor U23011 (N_23011,N_19819,N_19725);
and U23012 (N_23012,N_18431,N_15851);
and U23013 (N_23013,N_19160,N_16710);
and U23014 (N_23014,N_15828,N_15110);
nor U23015 (N_23015,N_18022,N_18262);
nor U23016 (N_23016,N_17521,N_16838);
and U23017 (N_23017,N_19655,N_16835);
or U23018 (N_23018,N_17856,N_16650);
and U23019 (N_23019,N_16907,N_17632);
nand U23020 (N_23020,N_17891,N_18144);
nand U23021 (N_23021,N_15615,N_16327);
and U23022 (N_23022,N_18560,N_19006);
nand U23023 (N_23023,N_15703,N_16204);
xnor U23024 (N_23024,N_19276,N_15045);
or U23025 (N_23025,N_16762,N_19892);
nor U23026 (N_23026,N_19538,N_16837);
nand U23027 (N_23027,N_15490,N_17814);
and U23028 (N_23028,N_19787,N_17623);
xor U23029 (N_23029,N_18706,N_18728);
nand U23030 (N_23030,N_17545,N_17060);
xnor U23031 (N_23031,N_18296,N_18530);
and U23032 (N_23032,N_15586,N_18194);
xnor U23033 (N_23033,N_16132,N_16702);
and U23034 (N_23034,N_17682,N_19321);
xor U23035 (N_23035,N_15601,N_17366);
or U23036 (N_23036,N_19129,N_17965);
or U23037 (N_23037,N_18988,N_15232);
xnor U23038 (N_23038,N_18548,N_16627);
xnor U23039 (N_23039,N_17838,N_19098);
and U23040 (N_23040,N_17281,N_19865);
and U23041 (N_23041,N_19264,N_17612);
and U23042 (N_23042,N_16682,N_19339);
and U23043 (N_23043,N_16083,N_17765);
or U23044 (N_23044,N_16753,N_17439);
or U23045 (N_23045,N_18046,N_15720);
or U23046 (N_23046,N_16342,N_15994);
nand U23047 (N_23047,N_17968,N_15156);
xnor U23048 (N_23048,N_18938,N_18396);
or U23049 (N_23049,N_19363,N_15711);
nand U23050 (N_23050,N_16542,N_18984);
nor U23051 (N_23051,N_15067,N_15475);
nor U23052 (N_23052,N_15177,N_16529);
nand U23053 (N_23053,N_15895,N_17173);
and U23054 (N_23054,N_17542,N_15745);
and U23055 (N_23055,N_15534,N_16339);
xor U23056 (N_23056,N_16508,N_16493);
nor U23057 (N_23057,N_17788,N_17891);
or U23058 (N_23058,N_19242,N_18433);
xnor U23059 (N_23059,N_17695,N_18737);
and U23060 (N_23060,N_18758,N_15423);
and U23061 (N_23061,N_17573,N_18294);
nor U23062 (N_23062,N_19483,N_17210);
nor U23063 (N_23063,N_18686,N_15952);
nand U23064 (N_23064,N_16480,N_17909);
xnor U23065 (N_23065,N_18972,N_16434);
nand U23066 (N_23066,N_18732,N_17664);
or U23067 (N_23067,N_16849,N_19257);
nor U23068 (N_23068,N_19987,N_19180);
xor U23069 (N_23069,N_18826,N_19448);
nor U23070 (N_23070,N_19486,N_15349);
and U23071 (N_23071,N_16542,N_19938);
and U23072 (N_23072,N_17939,N_17800);
nor U23073 (N_23073,N_16536,N_18752);
nor U23074 (N_23074,N_15493,N_19045);
or U23075 (N_23075,N_16635,N_18820);
and U23076 (N_23076,N_18940,N_15484);
nor U23077 (N_23077,N_18249,N_15296);
xor U23078 (N_23078,N_18170,N_17712);
xor U23079 (N_23079,N_17773,N_15497);
nor U23080 (N_23080,N_18721,N_15190);
nor U23081 (N_23081,N_17841,N_16339);
or U23082 (N_23082,N_16509,N_17481);
and U23083 (N_23083,N_19889,N_16976);
or U23084 (N_23084,N_15773,N_17328);
or U23085 (N_23085,N_17258,N_17817);
nor U23086 (N_23086,N_15626,N_17156);
and U23087 (N_23087,N_17039,N_15988);
nand U23088 (N_23088,N_18901,N_17249);
nand U23089 (N_23089,N_15824,N_15622);
xnor U23090 (N_23090,N_16329,N_19169);
xnor U23091 (N_23091,N_19071,N_19067);
nor U23092 (N_23092,N_18857,N_17684);
nand U23093 (N_23093,N_19515,N_16699);
nor U23094 (N_23094,N_18671,N_19012);
and U23095 (N_23095,N_17144,N_17931);
nand U23096 (N_23096,N_17733,N_17067);
nor U23097 (N_23097,N_17322,N_19911);
and U23098 (N_23098,N_16061,N_17202);
nor U23099 (N_23099,N_16614,N_16154);
or U23100 (N_23100,N_15037,N_15949);
nand U23101 (N_23101,N_17839,N_19395);
and U23102 (N_23102,N_19817,N_15590);
and U23103 (N_23103,N_19720,N_15814);
nand U23104 (N_23104,N_17129,N_17862);
nor U23105 (N_23105,N_19066,N_19302);
or U23106 (N_23106,N_15037,N_16420);
nand U23107 (N_23107,N_19810,N_18180);
nor U23108 (N_23108,N_16079,N_17363);
nand U23109 (N_23109,N_16213,N_15700);
and U23110 (N_23110,N_18894,N_16691);
and U23111 (N_23111,N_19288,N_19180);
and U23112 (N_23112,N_15849,N_18327);
xor U23113 (N_23113,N_15590,N_16241);
or U23114 (N_23114,N_19979,N_18803);
xnor U23115 (N_23115,N_15961,N_15000);
xnor U23116 (N_23116,N_16431,N_19589);
nand U23117 (N_23117,N_17330,N_18089);
or U23118 (N_23118,N_18097,N_18361);
xnor U23119 (N_23119,N_18880,N_16463);
xor U23120 (N_23120,N_16271,N_17456);
nor U23121 (N_23121,N_16676,N_15966);
nor U23122 (N_23122,N_17410,N_15449);
or U23123 (N_23123,N_19307,N_17114);
xor U23124 (N_23124,N_15579,N_16038);
xor U23125 (N_23125,N_15479,N_16927);
nor U23126 (N_23126,N_16454,N_19670);
nand U23127 (N_23127,N_15248,N_19877);
xnor U23128 (N_23128,N_17639,N_19248);
or U23129 (N_23129,N_15556,N_15240);
nand U23130 (N_23130,N_19085,N_15302);
or U23131 (N_23131,N_19414,N_16853);
and U23132 (N_23132,N_16573,N_18785);
nand U23133 (N_23133,N_15959,N_16024);
or U23134 (N_23134,N_19992,N_18087);
xnor U23135 (N_23135,N_15792,N_18889);
nand U23136 (N_23136,N_15113,N_19189);
nor U23137 (N_23137,N_17246,N_17192);
and U23138 (N_23138,N_18585,N_19657);
nand U23139 (N_23139,N_16576,N_15634);
and U23140 (N_23140,N_15706,N_16290);
or U23141 (N_23141,N_19317,N_18939);
nor U23142 (N_23142,N_17805,N_18978);
nor U23143 (N_23143,N_18236,N_17663);
nor U23144 (N_23144,N_19351,N_15861);
xnor U23145 (N_23145,N_17981,N_15856);
xor U23146 (N_23146,N_19599,N_17247);
xor U23147 (N_23147,N_18156,N_15222);
and U23148 (N_23148,N_18173,N_17408);
xor U23149 (N_23149,N_17562,N_17666);
nand U23150 (N_23150,N_17505,N_15017);
nor U23151 (N_23151,N_17703,N_15715);
or U23152 (N_23152,N_15994,N_15769);
xor U23153 (N_23153,N_16727,N_18321);
xnor U23154 (N_23154,N_15760,N_15097);
or U23155 (N_23155,N_15159,N_16584);
and U23156 (N_23156,N_19907,N_17737);
nand U23157 (N_23157,N_19693,N_17108);
xor U23158 (N_23158,N_17989,N_19169);
xor U23159 (N_23159,N_19839,N_15081);
nor U23160 (N_23160,N_15007,N_15582);
xor U23161 (N_23161,N_17533,N_18818);
nand U23162 (N_23162,N_17021,N_16761);
or U23163 (N_23163,N_15344,N_16567);
xor U23164 (N_23164,N_19267,N_17642);
or U23165 (N_23165,N_16768,N_19817);
and U23166 (N_23166,N_18136,N_19712);
or U23167 (N_23167,N_19912,N_17384);
xnor U23168 (N_23168,N_19444,N_16209);
nand U23169 (N_23169,N_19216,N_19726);
xor U23170 (N_23170,N_15879,N_16722);
xnor U23171 (N_23171,N_18270,N_15586);
nor U23172 (N_23172,N_16676,N_17506);
xnor U23173 (N_23173,N_19600,N_17750);
nor U23174 (N_23174,N_17764,N_18949);
nand U23175 (N_23175,N_18272,N_18489);
and U23176 (N_23176,N_16610,N_17125);
and U23177 (N_23177,N_16634,N_15532);
xor U23178 (N_23178,N_18818,N_16787);
or U23179 (N_23179,N_19076,N_15966);
xnor U23180 (N_23180,N_15803,N_15638);
nor U23181 (N_23181,N_19503,N_19471);
and U23182 (N_23182,N_19100,N_18734);
xor U23183 (N_23183,N_19798,N_17293);
nor U23184 (N_23184,N_18183,N_18948);
xnor U23185 (N_23185,N_17257,N_18245);
and U23186 (N_23186,N_17567,N_16889);
xor U23187 (N_23187,N_17324,N_17489);
xnor U23188 (N_23188,N_15965,N_16821);
xor U23189 (N_23189,N_17642,N_15911);
or U23190 (N_23190,N_15079,N_16014);
nand U23191 (N_23191,N_16084,N_15896);
and U23192 (N_23192,N_18881,N_16814);
and U23193 (N_23193,N_16161,N_15398);
xor U23194 (N_23194,N_17431,N_19868);
or U23195 (N_23195,N_16015,N_17413);
nor U23196 (N_23196,N_17461,N_15164);
and U23197 (N_23197,N_19883,N_16054);
or U23198 (N_23198,N_15587,N_15409);
and U23199 (N_23199,N_15580,N_15293);
or U23200 (N_23200,N_15496,N_17576);
or U23201 (N_23201,N_17656,N_18792);
and U23202 (N_23202,N_17870,N_17652);
nor U23203 (N_23203,N_16433,N_17072);
nand U23204 (N_23204,N_18707,N_15265);
nand U23205 (N_23205,N_16301,N_15157);
xnor U23206 (N_23206,N_18800,N_15514);
nand U23207 (N_23207,N_15381,N_18894);
nor U23208 (N_23208,N_17957,N_17696);
nor U23209 (N_23209,N_17838,N_18129);
nor U23210 (N_23210,N_17981,N_17903);
and U23211 (N_23211,N_17982,N_16962);
nand U23212 (N_23212,N_19339,N_15999);
and U23213 (N_23213,N_15461,N_17635);
or U23214 (N_23214,N_17592,N_16677);
and U23215 (N_23215,N_17113,N_18117);
nor U23216 (N_23216,N_17667,N_19941);
and U23217 (N_23217,N_15328,N_16501);
nand U23218 (N_23218,N_15283,N_15590);
and U23219 (N_23219,N_18259,N_19829);
nand U23220 (N_23220,N_19239,N_18138);
or U23221 (N_23221,N_17233,N_15870);
nor U23222 (N_23222,N_19515,N_18084);
nor U23223 (N_23223,N_17434,N_17195);
nor U23224 (N_23224,N_16076,N_17710);
xor U23225 (N_23225,N_15968,N_16499);
or U23226 (N_23226,N_18992,N_16413);
nand U23227 (N_23227,N_15856,N_17175);
nor U23228 (N_23228,N_17937,N_18190);
nand U23229 (N_23229,N_16889,N_18114);
xor U23230 (N_23230,N_18417,N_17256);
nor U23231 (N_23231,N_18816,N_17067);
and U23232 (N_23232,N_19109,N_15041);
nor U23233 (N_23233,N_16289,N_19171);
or U23234 (N_23234,N_18993,N_19021);
nand U23235 (N_23235,N_16039,N_19522);
nor U23236 (N_23236,N_18785,N_15133);
nor U23237 (N_23237,N_15608,N_18111);
nand U23238 (N_23238,N_18572,N_15295);
nor U23239 (N_23239,N_16377,N_17682);
xnor U23240 (N_23240,N_16721,N_18202);
and U23241 (N_23241,N_15732,N_17246);
or U23242 (N_23242,N_16981,N_17634);
or U23243 (N_23243,N_16128,N_18874);
xor U23244 (N_23244,N_18618,N_18446);
nand U23245 (N_23245,N_17587,N_16714);
nand U23246 (N_23246,N_18822,N_16167);
nand U23247 (N_23247,N_19171,N_15127);
or U23248 (N_23248,N_19930,N_15885);
or U23249 (N_23249,N_19713,N_19842);
and U23250 (N_23250,N_17517,N_19328);
xnor U23251 (N_23251,N_17079,N_19081);
or U23252 (N_23252,N_19642,N_17492);
nor U23253 (N_23253,N_19452,N_18189);
nor U23254 (N_23254,N_16784,N_19593);
and U23255 (N_23255,N_17944,N_15983);
or U23256 (N_23256,N_16563,N_17705);
xor U23257 (N_23257,N_16270,N_19853);
and U23258 (N_23258,N_18349,N_15063);
nor U23259 (N_23259,N_19205,N_18141);
xor U23260 (N_23260,N_16457,N_19293);
nand U23261 (N_23261,N_19110,N_17412);
xor U23262 (N_23262,N_15663,N_17287);
nand U23263 (N_23263,N_17486,N_17000);
nor U23264 (N_23264,N_18266,N_19474);
nor U23265 (N_23265,N_19334,N_19234);
xnor U23266 (N_23266,N_18925,N_15269);
or U23267 (N_23267,N_15791,N_18343);
nand U23268 (N_23268,N_19266,N_19217);
xnor U23269 (N_23269,N_17454,N_16063);
or U23270 (N_23270,N_17176,N_15746);
nand U23271 (N_23271,N_18174,N_18785);
and U23272 (N_23272,N_19963,N_16322);
xnor U23273 (N_23273,N_15656,N_16130);
nor U23274 (N_23274,N_15957,N_18489);
or U23275 (N_23275,N_17085,N_19390);
nor U23276 (N_23276,N_19847,N_15590);
nor U23277 (N_23277,N_19533,N_15116);
xor U23278 (N_23278,N_17633,N_15326);
and U23279 (N_23279,N_18936,N_15022);
or U23280 (N_23280,N_19128,N_18900);
or U23281 (N_23281,N_16613,N_19282);
or U23282 (N_23282,N_18351,N_15668);
or U23283 (N_23283,N_18370,N_15499);
and U23284 (N_23284,N_18234,N_18065);
nor U23285 (N_23285,N_19823,N_17659);
xor U23286 (N_23286,N_16543,N_18095);
and U23287 (N_23287,N_15498,N_16543);
xnor U23288 (N_23288,N_15533,N_15115);
xnor U23289 (N_23289,N_16977,N_19734);
and U23290 (N_23290,N_16258,N_16851);
nor U23291 (N_23291,N_19205,N_17871);
nand U23292 (N_23292,N_18226,N_17998);
nor U23293 (N_23293,N_15116,N_15020);
or U23294 (N_23294,N_19647,N_19353);
nand U23295 (N_23295,N_16982,N_18679);
nand U23296 (N_23296,N_18283,N_17067);
or U23297 (N_23297,N_16467,N_19899);
xnor U23298 (N_23298,N_18118,N_17937);
or U23299 (N_23299,N_16856,N_18194);
and U23300 (N_23300,N_19208,N_19701);
nor U23301 (N_23301,N_19175,N_15069);
or U23302 (N_23302,N_19147,N_16405);
or U23303 (N_23303,N_17661,N_15497);
xnor U23304 (N_23304,N_18058,N_17759);
nand U23305 (N_23305,N_17103,N_15521);
xnor U23306 (N_23306,N_17454,N_18608);
nor U23307 (N_23307,N_17163,N_15461);
and U23308 (N_23308,N_19326,N_19227);
xor U23309 (N_23309,N_19232,N_18112);
and U23310 (N_23310,N_18694,N_17697);
and U23311 (N_23311,N_15690,N_17443);
or U23312 (N_23312,N_18053,N_17415);
nand U23313 (N_23313,N_19274,N_15923);
xnor U23314 (N_23314,N_16986,N_18626);
nand U23315 (N_23315,N_16688,N_16289);
xor U23316 (N_23316,N_17826,N_16485);
or U23317 (N_23317,N_17163,N_19709);
nor U23318 (N_23318,N_18220,N_15996);
and U23319 (N_23319,N_16205,N_15735);
nor U23320 (N_23320,N_17003,N_16712);
nand U23321 (N_23321,N_19783,N_17557);
or U23322 (N_23322,N_17399,N_16419);
xnor U23323 (N_23323,N_15009,N_16198);
xor U23324 (N_23324,N_17861,N_19676);
xor U23325 (N_23325,N_16450,N_19925);
or U23326 (N_23326,N_15836,N_15075);
nand U23327 (N_23327,N_19083,N_15901);
nor U23328 (N_23328,N_15231,N_18391);
nor U23329 (N_23329,N_19801,N_15203);
nand U23330 (N_23330,N_16172,N_15978);
nand U23331 (N_23331,N_19565,N_18267);
nand U23332 (N_23332,N_18827,N_19871);
or U23333 (N_23333,N_17893,N_19224);
nor U23334 (N_23334,N_16933,N_16926);
nor U23335 (N_23335,N_15147,N_17741);
xor U23336 (N_23336,N_18399,N_15431);
and U23337 (N_23337,N_19648,N_19822);
and U23338 (N_23338,N_18967,N_16734);
and U23339 (N_23339,N_18064,N_17134);
nor U23340 (N_23340,N_17462,N_15815);
xnor U23341 (N_23341,N_16887,N_15614);
and U23342 (N_23342,N_19503,N_16415);
and U23343 (N_23343,N_19043,N_15838);
xor U23344 (N_23344,N_15227,N_18933);
and U23345 (N_23345,N_15745,N_18703);
xor U23346 (N_23346,N_19921,N_16338);
nor U23347 (N_23347,N_19725,N_19321);
nand U23348 (N_23348,N_15697,N_18802);
or U23349 (N_23349,N_17537,N_16435);
or U23350 (N_23350,N_16092,N_19767);
or U23351 (N_23351,N_15761,N_15887);
and U23352 (N_23352,N_16383,N_18613);
nor U23353 (N_23353,N_19667,N_18385);
nand U23354 (N_23354,N_15941,N_16533);
or U23355 (N_23355,N_16786,N_17633);
and U23356 (N_23356,N_16469,N_19624);
nand U23357 (N_23357,N_18042,N_15855);
xor U23358 (N_23358,N_17295,N_17373);
nor U23359 (N_23359,N_15128,N_19186);
nand U23360 (N_23360,N_16981,N_19324);
nor U23361 (N_23361,N_19081,N_17666);
xnor U23362 (N_23362,N_19824,N_16957);
nor U23363 (N_23363,N_17027,N_19005);
nand U23364 (N_23364,N_17834,N_19563);
or U23365 (N_23365,N_19938,N_18067);
and U23366 (N_23366,N_15770,N_15549);
nand U23367 (N_23367,N_16041,N_17658);
nor U23368 (N_23368,N_18798,N_18970);
xor U23369 (N_23369,N_19738,N_19758);
nand U23370 (N_23370,N_17949,N_18518);
xor U23371 (N_23371,N_18285,N_15942);
and U23372 (N_23372,N_19366,N_17357);
nor U23373 (N_23373,N_15022,N_16225);
or U23374 (N_23374,N_19498,N_17584);
nand U23375 (N_23375,N_18119,N_18946);
nor U23376 (N_23376,N_16241,N_15470);
nand U23377 (N_23377,N_18579,N_15293);
xnor U23378 (N_23378,N_17921,N_18301);
nand U23379 (N_23379,N_18168,N_15646);
and U23380 (N_23380,N_18447,N_19745);
nor U23381 (N_23381,N_19771,N_18333);
xnor U23382 (N_23382,N_18107,N_19568);
xor U23383 (N_23383,N_17905,N_19906);
and U23384 (N_23384,N_18640,N_17651);
nor U23385 (N_23385,N_16972,N_15349);
xor U23386 (N_23386,N_17006,N_19840);
nor U23387 (N_23387,N_19819,N_16016);
and U23388 (N_23388,N_15617,N_15869);
nand U23389 (N_23389,N_19973,N_17867);
nor U23390 (N_23390,N_16037,N_18313);
or U23391 (N_23391,N_19483,N_19797);
or U23392 (N_23392,N_18660,N_19631);
nor U23393 (N_23393,N_15061,N_16264);
or U23394 (N_23394,N_17726,N_17708);
or U23395 (N_23395,N_16333,N_16597);
or U23396 (N_23396,N_16353,N_15176);
and U23397 (N_23397,N_17163,N_16173);
nand U23398 (N_23398,N_16100,N_18026);
and U23399 (N_23399,N_16377,N_18965);
or U23400 (N_23400,N_18060,N_19785);
nand U23401 (N_23401,N_19457,N_18361);
or U23402 (N_23402,N_16643,N_17395);
or U23403 (N_23403,N_18230,N_18408);
nor U23404 (N_23404,N_16782,N_18174);
nor U23405 (N_23405,N_19710,N_19043);
or U23406 (N_23406,N_15053,N_18399);
and U23407 (N_23407,N_18186,N_19890);
nand U23408 (N_23408,N_16558,N_19254);
xnor U23409 (N_23409,N_17576,N_16389);
nor U23410 (N_23410,N_18553,N_17548);
xor U23411 (N_23411,N_18139,N_17845);
and U23412 (N_23412,N_15537,N_17926);
xnor U23413 (N_23413,N_16292,N_16682);
nor U23414 (N_23414,N_19592,N_16770);
nand U23415 (N_23415,N_19036,N_16876);
xor U23416 (N_23416,N_18271,N_16258);
or U23417 (N_23417,N_16522,N_19157);
nor U23418 (N_23418,N_16905,N_15436);
and U23419 (N_23419,N_18069,N_15393);
nand U23420 (N_23420,N_15124,N_18279);
and U23421 (N_23421,N_19978,N_19487);
or U23422 (N_23422,N_15432,N_16170);
nor U23423 (N_23423,N_15142,N_17959);
or U23424 (N_23424,N_16565,N_19241);
xor U23425 (N_23425,N_15911,N_17853);
xnor U23426 (N_23426,N_19558,N_19169);
xor U23427 (N_23427,N_19620,N_16127);
and U23428 (N_23428,N_16990,N_18670);
nor U23429 (N_23429,N_15635,N_19086);
nand U23430 (N_23430,N_15067,N_15808);
xnor U23431 (N_23431,N_16953,N_16739);
xnor U23432 (N_23432,N_15138,N_18085);
nand U23433 (N_23433,N_16974,N_17979);
nand U23434 (N_23434,N_15580,N_19719);
or U23435 (N_23435,N_19963,N_16105);
nand U23436 (N_23436,N_15963,N_18183);
xnor U23437 (N_23437,N_18275,N_15099);
and U23438 (N_23438,N_16743,N_18704);
nand U23439 (N_23439,N_15571,N_18224);
nor U23440 (N_23440,N_18236,N_18807);
and U23441 (N_23441,N_19599,N_17317);
xnor U23442 (N_23442,N_16330,N_16282);
and U23443 (N_23443,N_18713,N_17868);
nor U23444 (N_23444,N_17121,N_19504);
nand U23445 (N_23445,N_15515,N_15304);
or U23446 (N_23446,N_17225,N_17541);
nand U23447 (N_23447,N_15441,N_18334);
nor U23448 (N_23448,N_17212,N_16230);
and U23449 (N_23449,N_18667,N_18502);
or U23450 (N_23450,N_17593,N_17873);
and U23451 (N_23451,N_16627,N_17827);
nand U23452 (N_23452,N_18781,N_16780);
nand U23453 (N_23453,N_16129,N_15860);
or U23454 (N_23454,N_17612,N_16020);
nor U23455 (N_23455,N_18523,N_18236);
or U23456 (N_23456,N_16560,N_18965);
or U23457 (N_23457,N_16530,N_15229);
or U23458 (N_23458,N_15347,N_16810);
nand U23459 (N_23459,N_17615,N_15591);
nor U23460 (N_23460,N_19048,N_17200);
and U23461 (N_23461,N_19954,N_19536);
nand U23462 (N_23462,N_18401,N_17047);
and U23463 (N_23463,N_18436,N_15647);
or U23464 (N_23464,N_15713,N_18136);
and U23465 (N_23465,N_16524,N_17202);
xor U23466 (N_23466,N_18056,N_18305);
and U23467 (N_23467,N_19808,N_18329);
xnor U23468 (N_23468,N_15537,N_18401);
and U23469 (N_23469,N_17525,N_15008);
nand U23470 (N_23470,N_19777,N_15850);
or U23471 (N_23471,N_15463,N_16146);
nor U23472 (N_23472,N_17254,N_19734);
and U23473 (N_23473,N_18126,N_19548);
and U23474 (N_23474,N_15993,N_15084);
or U23475 (N_23475,N_19088,N_16781);
and U23476 (N_23476,N_19399,N_16377);
or U23477 (N_23477,N_17245,N_16477);
nor U23478 (N_23478,N_17559,N_19838);
and U23479 (N_23479,N_18301,N_15524);
nand U23480 (N_23480,N_17188,N_17701);
nand U23481 (N_23481,N_16221,N_15577);
and U23482 (N_23482,N_15145,N_15267);
or U23483 (N_23483,N_15327,N_15662);
and U23484 (N_23484,N_16229,N_18780);
nand U23485 (N_23485,N_17293,N_17099);
nand U23486 (N_23486,N_16876,N_17707);
xnor U23487 (N_23487,N_16623,N_15661);
nand U23488 (N_23488,N_18212,N_17510);
nand U23489 (N_23489,N_17599,N_17019);
nand U23490 (N_23490,N_18735,N_16037);
nand U23491 (N_23491,N_18920,N_18636);
and U23492 (N_23492,N_19554,N_16803);
nand U23493 (N_23493,N_17513,N_15230);
nand U23494 (N_23494,N_18157,N_17143);
and U23495 (N_23495,N_16338,N_16235);
nand U23496 (N_23496,N_16545,N_17207);
xnor U23497 (N_23497,N_17936,N_18430);
nand U23498 (N_23498,N_19152,N_17130);
xor U23499 (N_23499,N_18499,N_15014);
and U23500 (N_23500,N_16632,N_18236);
nor U23501 (N_23501,N_15610,N_18502);
nor U23502 (N_23502,N_19081,N_18425);
nor U23503 (N_23503,N_19954,N_19795);
or U23504 (N_23504,N_16504,N_15204);
nor U23505 (N_23505,N_17021,N_16486);
or U23506 (N_23506,N_18482,N_17223);
xor U23507 (N_23507,N_18235,N_19174);
or U23508 (N_23508,N_16393,N_15618);
or U23509 (N_23509,N_17317,N_19638);
nand U23510 (N_23510,N_16654,N_15761);
or U23511 (N_23511,N_16304,N_16912);
nand U23512 (N_23512,N_15324,N_18907);
xnor U23513 (N_23513,N_16339,N_15923);
nor U23514 (N_23514,N_19194,N_17414);
nor U23515 (N_23515,N_15999,N_17018);
or U23516 (N_23516,N_18960,N_15364);
and U23517 (N_23517,N_17776,N_19211);
nand U23518 (N_23518,N_16280,N_17142);
and U23519 (N_23519,N_16741,N_18005);
and U23520 (N_23520,N_15037,N_16604);
nor U23521 (N_23521,N_17096,N_16565);
nor U23522 (N_23522,N_17985,N_19990);
or U23523 (N_23523,N_17609,N_18946);
nand U23524 (N_23524,N_16878,N_17066);
nor U23525 (N_23525,N_16097,N_17531);
nor U23526 (N_23526,N_15048,N_17838);
and U23527 (N_23527,N_16502,N_16429);
nand U23528 (N_23528,N_17374,N_19838);
nor U23529 (N_23529,N_16740,N_16886);
xnor U23530 (N_23530,N_15220,N_18733);
and U23531 (N_23531,N_18286,N_18671);
nand U23532 (N_23532,N_18363,N_18548);
xor U23533 (N_23533,N_18982,N_16435);
nor U23534 (N_23534,N_17081,N_17094);
xnor U23535 (N_23535,N_19350,N_16677);
or U23536 (N_23536,N_18065,N_18288);
xnor U23537 (N_23537,N_16752,N_18022);
xnor U23538 (N_23538,N_16403,N_18173);
or U23539 (N_23539,N_17222,N_17700);
nor U23540 (N_23540,N_16712,N_18910);
nor U23541 (N_23541,N_18045,N_17171);
nand U23542 (N_23542,N_16990,N_16961);
xnor U23543 (N_23543,N_17775,N_18957);
nand U23544 (N_23544,N_17154,N_19727);
nand U23545 (N_23545,N_15276,N_16285);
nand U23546 (N_23546,N_19606,N_16764);
xnor U23547 (N_23547,N_18499,N_16476);
nand U23548 (N_23548,N_17026,N_18403);
nor U23549 (N_23549,N_15812,N_15211);
nor U23550 (N_23550,N_18011,N_17624);
xor U23551 (N_23551,N_19830,N_15845);
and U23552 (N_23552,N_18201,N_18132);
and U23553 (N_23553,N_17977,N_17615);
or U23554 (N_23554,N_16971,N_16882);
and U23555 (N_23555,N_17640,N_17121);
or U23556 (N_23556,N_16027,N_17797);
nor U23557 (N_23557,N_16912,N_17892);
nor U23558 (N_23558,N_16605,N_19253);
or U23559 (N_23559,N_17893,N_16724);
or U23560 (N_23560,N_17881,N_18123);
nor U23561 (N_23561,N_19632,N_18387);
and U23562 (N_23562,N_19283,N_15735);
and U23563 (N_23563,N_16676,N_17725);
xor U23564 (N_23564,N_17682,N_16827);
nor U23565 (N_23565,N_16344,N_19556);
xor U23566 (N_23566,N_19299,N_17267);
nand U23567 (N_23567,N_16366,N_17232);
nor U23568 (N_23568,N_15601,N_15174);
nand U23569 (N_23569,N_16772,N_19734);
and U23570 (N_23570,N_18593,N_17985);
and U23571 (N_23571,N_17921,N_15817);
nor U23572 (N_23572,N_19720,N_19161);
xor U23573 (N_23573,N_15787,N_15463);
xnor U23574 (N_23574,N_19434,N_17122);
or U23575 (N_23575,N_17802,N_16931);
and U23576 (N_23576,N_15135,N_15629);
or U23577 (N_23577,N_16631,N_19707);
nand U23578 (N_23578,N_19004,N_18108);
nand U23579 (N_23579,N_16101,N_16247);
nand U23580 (N_23580,N_15563,N_15405);
xnor U23581 (N_23581,N_16683,N_18769);
xor U23582 (N_23582,N_17457,N_19617);
xor U23583 (N_23583,N_15588,N_17956);
and U23584 (N_23584,N_18784,N_17777);
nand U23585 (N_23585,N_16999,N_18787);
nor U23586 (N_23586,N_18176,N_18865);
or U23587 (N_23587,N_16396,N_18986);
and U23588 (N_23588,N_17501,N_15413);
nor U23589 (N_23589,N_16084,N_18398);
nand U23590 (N_23590,N_17888,N_18117);
or U23591 (N_23591,N_18051,N_18814);
and U23592 (N_23592,N_17353,N_19302);
nor U23593 (N_23593,N_18673,N_19256);
nor U23594 (N_23594,N_19156,N_17106);
and U23595 (N_23595,N_19758,N_16447);
nand U23596 (N_23596,N_19325,N_19040);
nor U23597 (N_23597,N_19402,N_16476);
or U23598 (N_23598,N_16258,N_19273);
xor U23599 (N_23599,N_19698,N_15268);
or U23600 (N_23600,N_15251,N_19247);
or U23601 (N_23601,N_17243,N_18593);
and U23602 (N_23602,N_19434,N_19309);
nand U23603 (N_23603,N_18586,N_16780);
nand U23604 (N_23604,N_17118,N_15795);
nor U23605 (N_23605,N_15772,N_17331);
nor U23606 (N_23606,N_18332,N_16564);
and U23607 (N_23607,N_18124,N_19370);
nor U23608 (N_23608,N_18664,N_16308);
xnor U23609 (N_23609,N_16631,N_15794);
nor U23610 (N_23610,N_17910,N_15557);
and U23611 (N_23611,N_17399,N_15392);
and U23612 (N_23612,N_17983,N_19829);
xor U23613 (N_23613,N_17561,N_18003);
and U23614 (N_23614,N_19944,N_18401);
nand U23615 (N_23615,N_17448,N_17059);
and U23616 (N_23616,N_15047,N_18255);
xor U23617 (N_23617,N_15517,N_15999);
nor U23618 (N_23618,N_16477,N_19160);
xor U23619 (N_23619,N_17569,N_16793);
and U23620 (N_23620,N_19711,N_16532);
nor U23621 (N_23621,N_19995,N_15123);
and U23622 (N_23622,N_17046,N_19646);
and U23623 (N_23623,N_17199,N_19539);
or U23624 (N_23624,N_19596,N_15342);
xnor U23625 (N_23625,N_15973,N_17053);
and U23626 (N_23626,N_15542,N_16443);
or U23627 (N_23627,N_19619,N_19604);
or U23628 (N_23628,N_16535,N_18729);
or U23629 (N_23629,N_16798,N_16202);
nand U23630 (N_23630,N_18783,N_15241);
nand U23631 (N_23631,N_17473,N_15683);
nor U23632 (N_23632,N_18653,N_18547);
nor U23633 (N_23633,N_19944,N_15307);
xor U23634 (N_23634,N_17474,N_18063);
nand U23635 (N_23635,N_16295,N_17994);
or U23636 (N_23636,N_17240,N_17948);
or U23637 (N_23637,N_17499,N_16278);
xor U23638 (N_23638,N_17840,N_19117);
xnor U23639 (N_23639,N_16252,N_16014);
nor U23640 (N_23640,N_18424,N_16921);
and U23641 (N_23641,N_19782,N_18844);
nor U23642 (N_23642,N_19298,N_18197);
or U23643 (N_23643,N_17825,N_15296);
nor U23644 (N_23644,N_19790,N_19721);
or U23645 (N_23645,N_17686,N_19322);
nor U23646 (N_23646,N_18202,N_18083);
nand U23647 (N_23647,N_18720,N_19720);
and U23648 (N_23648,N_15861,N_16838);
nor U23649 (N_23649,N_17497,N_18745);
nand U23650 (N_23650,N_15091,N_17812);
nor U23651 (N_23651,N_15909,N_17081);
and U23652 (N_23652,N_16601,N_16576);
and U23653 (N_23653,N_16977,N_19711);
and U23654 (N_23654,N_18872,N_19556);
and U23655 (N_23655,N_15738,N_19327);
nand U23656 (N_23656,N_15755,N_16363);
nor U23657 (N_23657,N_15549,N_15740);
and U23658 (N_23658,N_15649,N_16987);
and U23659 (N_23659,N_17843,N_15729);
and U23660 (N_23660,N_19867,N_17656);
and U23661 (N_23661,N_18302,N_17414);
and U23662 (N_23662,N_18668,N_18566);
nand U23663 (N_23663,N_16348,N_17628);
and U23664 (N_23664,N_19754,N_16081);
xor U23665 (N_23665,N_15315,N_16778);
nand U23666 (N_23666,N_19394,N_19056);
xnor U23667 (N_23667,N_18959,N_17245);
nor U23668 (N_23668,N_18231,N_15304);
xor U23669 (N_23669,N_16002,N_17038);
xor U23670 (N_23670,N_18907,N_19260);
nand U23671 (N_23671,N_17916,N_19227);
nor U23672 (N_23672,N_15710,N_19067);
and U23673 (N_23673,N_18765,N_18199);
xnor U23674 (N_23674,N_18995,N_19150);
xnor U23675 (N_23675,N_18737,N_16474);
or U23676 (N_23676,N_16525,N_15194);
nor U23677 (N_23677,N_16266,N_19152);
nor U23678 (N_23678,N_17305,N_18195);
xor U23679 (N_23679,N_18217,N_16170);
and U23680 (N_23680,N_16993,N_15086);
nand U23681 (N_23681,N_18997,N_17334);
xor U23682 (N_23682,N_15467,N_18806);
xnor U23683 (N_23683,N_17810,N_17214);
nor U23684 (N_23684,N_19996,N_17613);
nand U23685 (N_23685,N_18857,N_17167);
nor U23686 (N_23686,N_15647,N_17782);
nor U23687 (N_23687,N_15085,N_15076);
nor U23688 (N_23688,N_18188,N_17159);
xnor U23689 (N_23689,N_17944,N_15616);
xor U23690 (N_23690,N_18901,N_15155);
and U23691 (N_23691,N_15424,N_19220);
nor U23692 (N_23692,N_18237,N_17600);
and U23693 (N_23693,N_17860,N_19977);
xor U23694 (N_23694,N_16950,N_18601);
or U23695 (N_23695,N_15985,N_17650);
nand U23696 (N_23696,N_15581,N_18199);
xor U23697 (N_23697,N_16178,N_16632);
xor U23698 (N_23698,N_15685,N_17757);
or U23699 (N_23699,N_18062,N_15426);
or U23700 (N_23700,N_16317,N_17425);
nor U23701 (N_23701,N_15647,N_15454);
and U23702 (N_23702,N_17582,N_16487);
and U23703 (N_23703,N_18567,N_17597);
and U23704 (N_23704,N_19569,N_17381);
and U23705 (N_23705,N_15609,N_19009);
or U23706 (N_23706,N_19334,N_19065);
nand U23707 (N_23707,N_17296,N_16522);
and U23708 (N_23708,N_19177,N_18477);
or U23709 (N_23709,N_17022,N_17835);
or U23710 (N_23710,N_17436,N_15394);
nor U23711 (N_23711,N_18908,N_16848);
or U23712 (N_23712,N_15068,N_18839);
nor U23713 (N_23713,N_16171,N_16749);
xor U23714 (N_23714,N_17208,N_19634);
nor U23715 (N_23715,N_17091,N_19875);
xor U23716 (N_23716,N_17614,N_19772);
xor U23717 (N_23717,N_18909,N_16432);
or U23718 (N_23718,N_19924,N_15477);
xnor U23719 (N_23719,N_17093,N_17980);
nor U23720 (N_23720,N_15155,N_18777);
and U23721 (N_23721,N_15367,N_17150);
nor U23722 (N_23722,N_18715,N_17991);
or U23723 (N_23723,N_15628,N_15617);
and U23724 (N_23724,N_18786,N_18904);
or U23725 (N_23725,N_18229,N_17507);
and U23726 (N_23726,N_19434,N_16794);
xor U23727 (N_23727,N_17894,N_19758);
or U23728 (N_23728,N_18795,N_15575);
and U23729 (N_23729,N_18273,N_18457);
nor U23730 (N_23730,N_18947,N_15354);
or U23731 (N_23731,N_17832,N_16371);
nand U23732 (N_23732,N_15287,N_16076);
and U23733 (N_23733,N_17291,N_15770);
xnor U23734 (N_23734,N_16286,N_16831);
xnor U23735 (N_23735,N_18698,N_15353);
xnor U23736 (N_23736,N_15269,N_18902);
nor U23737 (N_23737,N_15709,N_18271);
nor U23738 (N_23738,N_19703,N_17278);
nor U23739 (N_23739,N_18031,N_19234);
nor U23740 (N_23740,N_18976,N_17527);
nor U23741 (N_23741,N_17760,N_17094);
or U23742 (N_23742,N_19943,N_19883);
and U23743 (N_23743,N_15127,N_16634);
nand U23744 (N_23744,N_17037,N_19312);
nand U23745 (N_23745,N_19607,N_16844);
and U23746 (N_23746,N_16718,N_17004);
or U23747 (N_23747,N_19862,N_16263);
or U23748 (N_23748,N_19130,N_15716);
and U23749 (N_23749,N_19589,N_16811);
or U23750 (N_23750,N_16214,N_19734);
or U23751 (N_23751,N_18922,N_19232);
xor U23752 (N_23752,N_17053,N_17751);
or U23753 (N_23753,N_17263,N_15686);
nand U23754 (N_23754,N_16984,N_16435);
or U23755 (N_23755,N_16942,N_15886);
nand U23756 (N_23756,N_17376,N_18988);
and U23757 (N_23757,N_18593,N_16911);
or U23758 (N_23758,N_16246,N_16034);
nor U23759 (N_23759,N_18048,N_17804);
nand U23760 (N_23760,N_16572,N_15513);
and U23761 (N_23761,N_18823,N_19301);
nor U23762 (N_23762,N_15269,N_17367);
or U23763 (N_23763,N_15320,N_16915);
xnor U23764 (N_23764,N_16280,N_18114);
or U23765 (N_23765,N_16909,N_18945);
or U23766 (N_23766,N_15688,N_19210);
or U23767 (N_23767,N_17566,N_16675);
nand U23768 (N_23768,N_15230,N_15526);
and U23769 (N_23769,N_15039,N_18830);
or U23770 (N_23770,N_18631,N_16146);
nand U23771 (N_23771,N_17799,N_19478);
and U23772 (N_23772,N_19048,N_19167);
nor U23773 (N_23773,N_15152,N_16780);
nor U23774 (N_23774,N_19532,N_19713);
nand U23775 (N_23775,N_19243,N_18325);
nor U23776 (N_23776,N_16249,N_18163);
nor U23777 (N_23777,N_15986,N_17682);
or U23778 (N_23778,N_19696,N_19159);
nand U23779 (N_23779,N_15270,N_15240);
nor U23780 (N_23780,N_19511,N_19832);
nor U23781 (N_23781,N_17001,N_17733);
nand U23782 (N_23782,N_19316,N_16270);
nand U23783 (N_23783,N_15222,N_16076);
nor U23784 (N_23784,N_15351,N_15679);
or U23785 (N_23785,N_17744,N_16190);
xnor U23786 (N_23786,N_17881,N_18872);
nand U23787 (N_23787,N_19218,N_15102);
nor U23788 (N_23788,N_18381,N_17926);
or U23789 (N_23789,N_18895,N_17066);
nand U23790 (N_23790,N_17691,N_19461);
or U23791 (N_23791,N_15183,N_16104);
xnor U23792 (N_23792,N_19294,N_18322);
nand U23793 (N_23793,N_16565,N_15680);
and U23794 (N_23794,N_19702,N_18285);
nor U23795 (N_23795,N_15241,N_18289);
and U23796 (N_23796,N_15493,N_15324);
nor U23797 (N_23797,N_17541,N_18502);
xor U23798 (N_23798,N_15215,N_16418);
nor U23799 (N_23799,N_16851,N_15935);
xor U23800 (N_23800,N_17467,N_17684);
or U23801 (N_23801,N_17504,N_15095);
or U23802 (N_23802,N_18346,N_19802);
nor U23803 (N_23803,N_15015,N_18397);
nand U23804 (N_23804,N_18022,N_17749);
nor U23805 (N_23805,N_16112,N_18131);
xnor U23806 (N_23806,N_16232,N_17434);
xor U23807 (N_23807,N_16681,N_19774);
and U23808 (N_23808,N_18636,N_15107);
xor U23809 (N_23809,N_18312,N_17243);
xnor U23810 (N_23810,N_19664,N_17617);
xor U23811 (N_23811,N_19406,N_17833);
nor U23812 (N_23812,N_19115,N_18057);
nand U23813 (N_23813,N_19848,N_15205);
and U23814 (N_23814,N_16631,N_17189);
and U23815 (N_23815,N_16279,N_16393);
nor U23816 (N_23816,N_18748,N_19026);
nor U23817 (N_23817,N_15547,N_17099);
and U23818 (N_23818,N_18062,N_18535);
nor U23819 (N_23819,N_18581,N_17535);
nor U23820 (N_23820,N_16641,N_16232);
and U23821 (N_23821,N_15153,N_19659);
or U23822 (N_23822,N_16614,N_16975);
or U23823 (N_23823,N_17763,N_19997);
xnor U23824 (N_23824,N_15681,N_19390);
or U23825 (N_23825,N_17775,N_19751);
xnor U23826 (N_23826,N_17849,N_16935);
xor U23827 (N_23827,N_18597,N_17892);
xnor U23828 (N_23828,N_17488,N_19335);
nor U23829 (N_23829,N_18395,N_17081);
nor U23830 (N_23830,N_16857,N_15939);
nor U23831 (N_23831,N_19725,N_16839);
nand U23832 (N_23832,N_16160,N_17882);
and U23833 (N_23833,N_15541,N_16303);
or U23834 (N_23834,N_15835,N_16502);
nand U23835 (N_23835,N_15108,N_18918);
or U23836 (N_23836,N_18405,N_15718);
and U23837 (N_23837,N_18503,N_16480);
and U23838 (N_23838,N_18198,N_16816);
or U23839 (N_23839,N_17285,N_18006);
nor U23840 (N_23840,N_19971,N_18319);
and U23841 (N_23841,N_16540,N_19553);
nor U23842 (N_23842,N_19946,N_16481);
or U23843 (N_23843,N_18079,N_19592);
nor U23844 (N_23844,N_15423,N_18792);
nor U23845 (N_23845,N_16280,N_18013);
nand U23846 (N_23846,N_18475,N_19661);
nor U23847 (N_23847,N_16843,N_18458);
and U23848 (N_23848,N_18753,N_17428);
nor U23849 (N_23849,N_18349,N_18226);
xnor U23850 (N_23850,N_16147,N_18600);
and U23851 (N_23851,N_16332,N_16404);
and U23852 (N_23852,N_15427,N_15495);
xor U23853 (N_23853,N_17670,N_16938);
or U23854 (N_23854,N_19954,N_19397);
xor U23855 (N_23855,N_17328,N_19745);
xor U23856 (N_23856,N_17767,N_18693);
nand U23857 (N_23857,N_18367,N_19520);
nand U23858 (N_23858,N_16337,N_19323);
xor U23859 (N_23859,N_15548,N_19942);
nor U23860 (N_23860,N_18261,N_18320);
or U23861 (N_23861,N_15671,N_19272);
nand U23862 (N_23862,N_15671,N_17976);
xor U23863 (N_23863,N_19832,N_15004);
or U23864 (N_23864,N_16090,N_18119);
nor U23865 (N_23865,N_17878,N_16827);
or U23866 (N_23866,N_16619,N_16584);
nand U23867 (N_23867,N_17344,N_18183);
or U23868 (N_23868,N_17724,N_17854);
or U23869 (N_23869,N_17911,N_17517);
xnor U23870 (N_23870,N_15041,N_18525);
or U23871 (N_23871,N_15023,N_19825);
xor U23872 (N_23872,N_17967,N_19448);
or U23873 (N_23873,N_15977,N_18128);
or U23874 (N_23874,N_16321,N_16981);
nor U23875 (N_23875,N_18673,N_16295);
and U23876 (N_23876,N_16838,N_16722);
nor U23877 (N_23877,N_15937,N_19712);
xnor U23878 (N_23878,N_15230,N_18596);
or U23879 (N_23879,N_19065,N_16417);
nand U23880 (N_23880,N_17137,N_17497);
xnor U23881 (N_23881,N_17267,N_17573);
nor U23882 (N_23882,N_15686,N_18856);
xor U23883 (N_23883,N_17957,N_19347);
or U23884 (N_23884,N_15885,N_17056);
and U23885 (N_23885,N_17305,N_15761);
nor U23886 (N_23886,N_17766,N_19104);
or U23887 (N_23887,N_19533,N_18017);
and U23888 (N_23888,N_17886,N_18383);
or U23889 (N_23889,N_15672,N_17654);
xor U23890 (N_23890,N_19612,N_19769);
nor U23891 (N_23891,N_16690,N_18432);
or U23892 (N_23892,N_16042,N_18262);
nand U23893 (N_23893,N_19460,N_15381);
xor U23894 (N_23894,N_16371,N_17010);
nand U23895 (N_23895,N_17510,N_17486);
or U23896 (N_23896,N_19248,N_15417);
nand U23897 (N_23897,N_17941,N_16890);
or U23898 (N_23898,N_16601,N_16843);
and U23899 (N_23899,N_17927,N_19688);
or U23900 (N_23900,N_19839,N_15174);
nand U23901 (N_23901,N_18669,N_18535);
and U23902 (N_23902,N_19038,N_18207);
nand U23903 (N_23903,N_19324,N_17331);
and U23904 (N_23904,N_18472,N_18240);
nor U23905 (N_23905,N_18868,N_18501);
or U23906 (N_23906,N_16320,N_18783);
and U23907 (N_23907,N_19044,N_15654);
nand U23908 (N_23908,N_17762,N_19509);
and U23909 (N_23909,N_19454,N_16475);
nand U23910 (N_23910,N_15638,N_15065);
nand U23911 (N_23911,N_16696,N_19416);
and U23912 (N_23912,N_16379,N_18767);
nand U23913 (N_23913,N_15664,N_15941);
and U23914 (N_23914,N_19350,N_19197);
nor U23915 (N_23915,N_15511,N_18802);
nand U23916 (N_23916,N_17454,N_15461);
nor U23917 (N_23917,N_19474,N_19483);
and U23918 (N_23918,N_16872,N_16223);
xor U23919 (N_23919,N_17201,N_15811);
xnor U23920 (N_23920,N_15628,N_15155);
nor U23921 (N_23921,N_19266,N_15248);
xnor U23922 (N_23922,N_17572,N_19624);
xnor U23923 (N_23923,N_18325,N_19611);
and U23924 (N_23924,N_18424,N_18144);
and U23925 (N_23925,N_16224,N_19845);
nor U23926 (N_23926,N_19834,N_15239);
nand U23927 (N_23927,N_17709,N_16608);
and U23928 (N_23928,N_19131,N_16017);
nand U23929 (N_23929,N_19027,N_16696);
xor U23930 (N_23930,N_17176,N_18350);
and U23931 (N_23931,N_19438,N_18476);
nor U23932 (N_23932,N_19073,N_15246);
nor U23933 (N_23933,N_15004,N_15811);
nor U23934 (N_23934,N_18906,N_19775);
nor U23935 (N_23935,N_18006,N_19055);
nor U23936 (N_23936,N_16832,N_19479);
xnor U23937 (N_23937,N_17767,N_18193);
nand U23938 (N_23938,N_16761,N_19457);
nand U23939 (N_23939,N_18187,N_15915);
nor U23940 (N_23940,N_18444,N_18996);
or U23941 (N_23941,N_18184,N_15928);
xor U23942 (N_23942,N_16410,N_18248);
nor U23943 (N_23943,N_19891,N_18802);
xor U23944 (N_23944,N_17153,N_18232);
xnor U23945 (N_23945,N_15099,N_17707);
or U23946 (N_23946,N_15059,N_16769);
nor U23947 (N_23947,N_16915,N_18850);
or U23948 (N_23948,N_16342,N_19683);
and U23949 (N_23949,N_15894,N_15834);
nor U23950 (N_23950,N_15083,N_16725);
and U23951 (N_23951,N_19729,N_17213);
and U23952 (N_23952,N_19480,N_18812);
and U23953 (N_23953,N_15472,N_15215);
and U23954 (N_23954,N_16601,N_15913);
xor U23955 (N_23955,N_15724,N_16557);
nor U23956 (N_23956,N_17863,N_15482);
nor U23957 (N_23957,N_18556,N_15572);
or U23958 (N_23958,N_16512,N_17672);
nand U23959 (N_23959,N_18634,N_19235);
nand U23960 (N_23960,N_17181,N_19489);
xor U23961 (N_23961,N_18039,N_19589);
xnor U23962 (N_23962,N_16945,N_15516);
xor U23963 (N_23963,N_16794,N_18423);
nor U23964 (N_23964,N_18102,N_19178);
and U23965 (N_23965,N_19363,N_16714);
or U23966 (N_23966,N_19430,N_17043);
nand U23967 (N_23967,N_15641,N_19986);
nand U23968 (N_23968,N_15698,N_16160);
or U23969 (N_23969,N_17387,N_19231);
xor U23970 (N_23970,N_15503,N_16899);
or U23971 (N_23971,N_17510,N_17687);
nand U23972 (N_23972,N_19448,N_19701);
xnor U23973 (N_23973,N_18570,N_16609);
or U23974 (N_23974,N_17037,N_15405);
and U23975 (N_23975,N_15572,N_17629);
nand U23976 (N_23976,N_19412,N_16618);
nand U23977 (N_23977,N_17705,N_17052);
xnor U23978 (N_23978,N_18753,N_18909);
nor U23979 (N_23979,N_16339,N_15426);
or U23980 (N_23980,N_19037,N_18356);
xnor U23981 (N_23981,N_15719,N_17905);
or U23982 (N_23982,N_16250,N_17873);
xnor U23983 (N_23983,N_16619,N_16359);
and U23984 (N_23984,N_15859,N_18914);
and U23985 (N_23985,N_17065,N_17512);
nand U23986 (N_23986,N_16388,N_15969);
or U23987 (N_23987,N_16857,N_17961);
nor U23988 (N_23988,N_16648,N_16870);
or U23989 (N_23989,N_19327,N_17884);
and U23990 (N_23990,N_15995,N_15016);
or U23991 (N_23991,N_17717,N_19199);
nor U23992 (N_23992,N_19781,N_16075);
or U23993 (N_23993,N_19697,N_15057);
xor U23994 (N_23994,N_16149,N_17990);
or U23995 (N_23995,N_15549,N_16681);
and U23996 (N_23996,N_15863,N_16526);
or U23997 (N_23997,N_16637,N_15888);
xor U23998 (N_23998,N_19689,N_16668);
nor U23999 (N_23999,N_15054,N_16195);
nor U24000 (N_24000,N_15087,N_18896);
nand U24001 (N_24001,N_19933,N_19155);
or U24002 (N_24002,N_16518,N_18639);
or U24003 (N_24003,N_15002,N_15108);
or U24004 (N_24004,N_15896,N_19648);
and U24005 (N_24005,N_18889,N_17809);
and U24006 (N_24006,N_17601,N_17614);
nor U24007 (N_24007,N_16866,N_16550);
or U24008 (N_24008,N_18722,N_19105);
and U24009 (N_24009,N_16947,N_19490);
and U24010 (N_24010,N_18122,N_16801);
nor U24011 (N_24011,N_19023,N_17196);
nand U24012 (N_24012,N_19853,N_17354);
or U24013 (N_24013,N_18337,N_18792);
xnor U24014 (N_24014,N_19654,N_15793);
xnor U24015 (N_24015,N_15262,N_19542);
xnor U24016 (N_24016,N_15490,N_18074);
nor U24017 (N_24017,N_16568,N_15880);
xnor U24018 (N_24018,N_18388,N_17002);
nor U24019 (N_24019,N_15940,N_17603);
nand U24020 (N_24020,N_15197,N_17510);
and U24021 (N_24021,N_18450,N_19048);
or U24022 (N_24022,N_17300,N_18240);
nor U24023 (N_24023,N_16962,N_17787);
nor U24024 (N_24024,N_18419,N_16617);
or U24025 (N_24025,N_16746,N_19935);
nor U24026 (N_24026,N_18322,N_15284);
or U24027 (N_24027,N_19482,N_17012);
xnor U24028 (N_24028,N_15961,N_15292);
or U24029 (N_24029,N_15939,N_16799);
and U24030 (N_24030,N_17619,N_19495);
nor U24031 (N_24031,N_16725,N_18938);
xor U24032 (N_24032,N_19593,N_19036);
nand U24033 (N_24033,N_17373,N_16549);
and U24034 (N_24034,N_16693,N_16516);
nor U24035 (N_24035,N_17401,N_18718);
nand U24036 (N_24036,N_15798,N_17089);
nor U24037 (N_24037,N_17005,N_17635);
and U24038 (N_24038,N_19826,N_16633);
or U24039 (N_24039,N_19273,N_19916);
and U24040 (N_24040,N_16856,N_17843);
nand U24041 (N_24041,N_16147,N_19140);
nor U24042 (N_24042,N_15761,N_15502);
nand U24043 (N_24043,N_16649,N_15153);
nand U24044 (N_24044,N_16255,N_17973);
xor U24045 (N_24045,N_18130,N_17535);
and U24046 (N_24046,N_18324,N_18247);
nand U24047 (N_24047,N_16322,N_18490);
nor U24048 (N_24048,N_16135,N_18649);
xnor U24049 (N_24049,N_15304,N_16730);
or U24050 (N_24050,N_17891,N_15400);
or U24051 (N_24051,N_15696,N_18293);
nor U24052 (N_24052,N_16179,N_15062);
nand U24053 (N_24053,N_18531,N_15220);
nor U24054 (N_24054,N_17968,N_16490);
nor U24055 (N_24055,N_17595,N_15113);
or U24056 (N_24056,N_19014,N_16230);
nand U24057 (N_24057,N_16644,N_18026);
xor U24058 (N_24058,N_15030,N_16771);
nor U24059 (N_24059,N_15018,N_18582);
xor U24060 (N_24060,N_16536,N_15214);
nor U24061 (N_24061,N_19957,N_19141);
and U24062 (N_24062,N_17573,N_19588);
nand U24063 (N_24063,N_16348,N_18992);
nor U24064 (N_24064,N_17347,N_19226);
nor U24065 (N_24065,N_19138,N_18512);
nand U24066 (N_24066,N_19612,N_18255);
nand U24067 (N_24067,N_18422,N_18080);
or U24068 (N_24068,N_16230,N_17812);
nand U24069 (N_24069,N_17671,N_15197);
nand U24070 (N_24070,N_15538,N_15094);
xnor U24071 (N_24071,N_17453,N_19529);
nor U24072 (N_24072,N_19187,N_17133);
nand U24073 (N_24073,N_15893,N_17464);
and U24074 (N_24074,N_16706,N_16955);
and U24075 (N_24075,N_16441,N_19204);
xor U24076 (N_24076,N_19707,N_15134);
or U24077 (N_24077,N_16526,N_19570);
nand U24078 (N_24078,N_16062,N_18018);
nor U24079 (N_24079,N_19070,N_18170);
and U24080 (N_24080,N_15871,N_17163);
nand U24081 (N_24081,N_19312,N_17636);
nor U24082 (N_24082,N_18036,N_19101);
nand U24083 (N_24083,N_16889,N_15737);
xnor U24084 (N_24084,N_17018,N_19977);
and U24085 (N_24085,N_17270,N_15326);
or U24086 (N_24086,N_18744,N_17708);
or U24087 (N_24087,N_16822,N_18236);
and U24088 (N_24088,N_19366,N_18410);
or U24089 (N_24089,N_18360,N_18181);
and U24090 (N_24090,N_18737,N_19418);
xnor U24091 (N_24091,N_17896,N_15164);
and U24092 (N_24092,N_19993,N_19588);
nand U24093 (N_24093,N_17039,N_19179);
and U24094 (N_24094,N_16590,N_16026);
nand U24095 (N_24095,N_17303,N_17022);
or U24096 (N_24096,N_17723,N_19662);
and U24097 (N_24097,N_17212,N_19808);
xor U24098 (N_24098,N_16044,N_18181);
nand U24099 (N_24099,N_17845,N_16537);
nor U24100 (N_24100,N_17595,N_16117);
nand U24101 (N_24101,N_15889,N_15017);
nor U24102 (N_24102,N_15455,N_18335);
xnor U24103 (N_24103,N_18862,N_18519);
or U24104 (N_24104,N_15539,N_16595);
xor U24105 (N_24105,N_15739,N_18014);
nand U24106 (N_24106,N_17413,N_15631);
nand U24107 (N_24107,N_16290,N_16503);
nand U24108 (N_24108,N_16989,N_15949);
or U24109 (N_24109,N_18877,N_15389);
and U24110 (N_24110,N_19646,N_15090);
and U24111 (N_24111,N_18923,N_15292);
nand U24112 (N_24112,N_15750,N_19478);
xor U24113 (N_24113,N_18257,N_18803);
nor U24114 (N_24114,N_18128,N_15076);
or U24115 (N_24115,N_19430,N_18981);
xnor U24116 (N_24116,N_15632,N_16564);
and U24117 (N_24117,N_17028,N_15175);
and U24118 (N_24118,N_19487,N_17160);
or U24119 (N_24119,N_16207,N_17350);
and U24120 (N_24120,N_15870,N_19672);
nand U24121 (N_24121,N_16995,N_19452);
or U24122 (N_24122,N_19964,N_15452);
and U24123 (N_24123,N_15248,N_15875);
and U24124 (N_24124,N_16861,N_16791);
nor U24125 (N_24125,N_16845,N_16657);
nor U24126 (N_24126,N_18221,N_18397);
or U24127 (N_24127,N_16151,N_18788);
nor U24128 (N_24128,N_17652,N_17011);
and U24129 (N_24129,N_18345,N_19732);
nor U24130 (N_24130,N_15257,N_16715);
nor U24131 (N_24131,N_19572,N_17500);
nor U24132 (N_24132,N_19585,N_18104);
or U24133 (N_24133,N_16887,N_15850);
xnor U24134 (N_24134,N_18594,N_19229);
or U24135 (N_24135,N_16774,N_18121);
nor U24136 (N_24136,N_17589,N_18065);
or U24137 (N_24137,N_17488,N_17358);
nor U24138 (N_24138,N_16121,N_19335);
and U24139 (N_24139,N_19119,N_18336);
and U24140 (N_24140,N_15726,N_16416);
or U24141 (N_24141,N_15946,N_16324);
and U24142 (N_24142,N_18182,N_18498);
and U24143 (N_24143,N_17922,N_15638);
nor U24144 (N_24144,N_18785,N_17624);
and U24145 (N_24145,N_15237,N_17155);
nor U24146 (N_24146,N_16054,N_16228);
nor U24147 (N_24147,N_17743,N_15005);
nor U24148 (N_24148,N_19214,N_19123);
and U24149 (N_24149,N_15564,N_15914);
nor U24150 (N_24150,N_16338,N_19094);
xor U24151 (N_24151,N_19905,N_18999);
xor U24152 (N_24152,N_16095,N_16287);
or U24153 (N_24153,N_19755,N_15710);
xnor U24154 (N_24154,N_16831,N_17403);
nor U24155 (N_24155,N_19892,N_16148);
and U24156 (N_24156,N_17243,N_18985);
nand U24157 (N_24157,N_16757,N_16342);
nand U24158 (N_24158,N_17102,N_18705);
and U24159 (N_24159,N_18870,N_19569);
xor U24160 (N_24160,N_16838,N_16035);
nand U24161 (N_24161,N_19402,N_15431);
and U24162 (N_24162,N_15426,N_17120);
nor U24163 (N_24163,N_17792,N_16513);
nor U24164 (N_24164,N_15509,N_18620);
or U24165 (N_24165,N_18109,N_19395);
or U24166 (N_24166,N_18083,N_15759);
xor U24167 (N_24167,N_17077,N_15348);
xnor U24168 (N_24168,N_19343,N_17767);
and U24169 (N_24169,N_16386,N_17701);
xnor U24170 (N_24170,N_19552,N_16581);
and U24171 (N_24171,N_17791,N_15092);
xor U24172 (N_24172,N_16625,N_17552);
nor U24173 (N_24173,N_15169,N_17780);
nor U24174 (N_24174,N_18130,N_18977);
or U24175 (N_24175,N_15834,N_16268);
nor U24176 (N_24176,N_19450,N_17787);
or U24177 (N_24177,N_17014,N_18225);
nand U24178 (N_24178,N_15576,N_15641);
and U24179 (N_24179,N_19044,N_18367);
nand U24180 (N_24180,N_15410,N_18553);
or U24181 (N_24181,N_19278,N_16189);
or U24182 (N_24182,N_16263,N_17740);
xnor U24183 (N_24183,N_19978,N_18671);
or U24184 (N_24184,N_16141,N_19530);
nor U24185 (N_24185,N_19543,N_17094);
and U24186 (N_24186,N_15352,N_18359);
xor U24187 (N_24187,N_17122,N_16957);
nand U24188 (N_24188,N_15044,N_15417);
nand U24189 (N_24189,N_17849,N_17177);
xnor U24190 (N_24190,N_17558,N_16942);
nand U24191 (N_24191,N_15256,N_15803);
nor U24192 (N_24192,N_18877,N_18736);
and U24193 (N_24193,N_17316,N_18551);
xnor U24194 (N_24194,N_17885,N_19333);
nand U24195 (N_24195,N_19351,N_19234);
nand U24196 (N_24196,N_18182,N_15240);
nand U24197 (N_24197,N_15943,N_19516);
nand U24198 (N_24198,N_18927,N_19770);
xnor U24199 (N_24199,N_19255,N_17029);
or U24200 (N_24200,N_15053,N_17787);
or U24201 (N_24201,N_15844,N_17899);
and U24202 (N_24202,N_16870,N_16160);
nand U24203 (N_24203,N_19020,N_19211);
xor U24204 (N_24204,N_19041,N_16083);
or U24205 (N_24205,N_15058,N_17569);
nor U24206 (N_24206,N_18783,N_18433);
nor U24207 (N_24207,N_17938,N_16643);
nor U24208 (N_24208,N_15686,N_15026);
xnor U24209 (N_24209,N_16749,N_15413);
nor U24210 (N_24210,N_18668,N_17977);
nor U24211 (N_24211,N_16495,N_15084);
or U24212 (N_24212,N_17487,N_16766);
xnor U24213 (N_24213,N_18433,N_16152);
or U24214 (N_24214,N_15471,N_17929);
and U24215 (N_24215,N_17933,N_19327);
or U24216 (N_24216,N_16842,N_17970);
or U24217 (N_24217,N_19078,N_18956);
or U24218 (N_24218,N_17720,N_16448);
xor U24219 (N_24219,N_18347,N_18779);
or U24220 (N_24220,N_17358,N_18663);
nand U24221 (N_24221,N_16129,N_18235);
and U24222 (N_24222,N_18246,N_16518);
or U24223 (N_24223,N_15232,N_19142);
xor U24224 (N_24224,N_15865,N_16494);
or U24225 (N_24225,N_18859,N_17324);
xor U24226 (N_24226,N_19240,N_16924);
and U24227 (N_24227,N_19320,N_19815);
and U24228 (N_24228,N_18339,N_18440);
nor U24229 (N_24229,N_17725,N_17416);
nor U24230 (N_24230,N_19285,N_19204);
nor U24231 (N_24231,N_18192,N_17446);
nor U24232 (N_24232,N_17630,N_18483);
xor U24233 (N_24233,N_19133,N_17401);
xnor U24234 (N_24234,N_18169,N_19892);
nand U24235 (N_24235,N_16980,N_18140);
and U24236 (N_24236,N_19045,N_18532);
nor U24237 (N_24237,N_19549,N_16708);
xor U24238 (N_24238,N_15983,N_16614);
nand U24239 (N_24239,N_17845,N_19805);
nor U24240 (N_24240,N_18512,N_17751);
xor U24241 (N_24241,N_16372,N_18330);
nor U24242 (N_24242,N_18352,N_16213);
nor U24243 (N_24243,N_18798,N_16520);
nor U24244 (N_24244,N_15884,N_17489);
nor U24245 (N_24245,N_19228,N_19598);
nand U24246 (N_24246,N_16988,N_17033);
or U24247 (N_24247,N_16687,N_16895);
and U24248 (N_24248,N_17695,N_16988);
nand U24249 (N_24249,N_16765,N_18473);
nor U24250 (N_24250,N_19545,N_18247);
nor U24251 (N_24251,N_16725,N_15034);
or U24252 (N_24252,N_17807,N_15906);
xor U24253 (N_24253,N_18853,N_15987);
xor U24254 (N_24254,N_15144,N_15779);
or U24255 (N_24255,N_16236,N_17157);
nor U24256 (N_24256,N_19356,N_19432);
or U24257 (N_24257,N_16668,N_16892);
nor U24258 (N_24258,N_15863,N_15735);
nand U24259 (N_24259,N_17609,N_18047);
nor U24260 (N_24260,N_17849,N_19341);
nor U24261 (N_24261,N_15523,N_18957);
or U24262 (N_24262,N_16816,N_18789);
nor U24263 (N_24263,N_15021,N_16986);
xnor U24264 (N_24264,N_19856,N_19750);
nand U24265 (N_24265,N_16505,N_17069);
nor U24266 (N_24266,N_18825,N_17468);
xnor U24267 (N_24267,N_16894,N_16856);
or U24268 (N_24268,N_18979,N_19591);
xnor U24269 (N_24269,N_15483,N_16552);
or U24270 (N_24270,N_17070,N_16369);
nand U24271 (N_24271,N_15173,N_17586);
or U24272 (N_24272,N_18330,N_16865);
nand U24273 (N_24273,N_19811,N_18066);
nand U24274 (N_24274,N_16616,N_15536);
and U24275 (N_24275,N_18669,N_17156);
nand U24276 (N_24276,N_17116,N_16549);
and U24277 (N_24277,N_16097,N_16150);
xor U24278 (N_24278,N_17408,N_19106);
and U24279 (N_24279,N_16009,N_17036);
xnor U24280 (N_24280,N_15220,N_17821);
or U24281 (N_24281,N_18732,N_18549);
nor U24282 (N_24282,N_17241,N_19441);
and U24283 (N_24283,N_15011,N_19086);
xor U24284 (N_24284,N_15779,N_16015);
xor U24285 (N_24285,N_18793,N_16023);
xnor U24286 (N_24286,N_19392,N_17449);
or U24287 (N_24287,N_16222,N_18563);
nand U24288 (N_24288,N_17824,N_17029);
or U24289 (N_24289,N_19952,N_19482);
and U24290 (N_24290,N_16943,N_16681);
nand U24291 (N_24291,N_17893,N_19941);
nor U24292 (N_24292,N_17207,N_15065);
xnor U24293 (N_24293,N_16797,N_19979);
nor U24294 (N_24294,N_15299,N_18971);
nand U24295 (N_24295,N_18525,N_16517);
xnor U24296 (N_24296,N_19304,N_16506);
nand U24297 (N_24297,N_15544,N_19699);
xor U24298 (N_24298,N_17086,N_16487);
and U24299 (N_24299,N_18068,N_15133);
xor U24300 (N_24300,N_18383,N_17917);
nand U24301 (N_24301,N_18962,N_16364);
or U24302 (N_24302,N_16410,N_15011);
and U24303 (N_24303,N_16422,N_18079);
nor U24304 (N_24304,N_18088,N_17224);
or U24305 (N_24305,N_16691,N_19556);
and U24306 (N_24306,N_15227,N_18298);
nor U24307 (N_24307,N_16630,N_16690);
nand U24308 (N_24308,N_18574,N_16502);
nor U24309 (N_24309,N_15022,N_19239);
nor U24310 (N_24310,N_18980,N_18220);
nand U24311 (N_24311,N_16491,N_15294);
nand U24312 (N_24312,N_17474,N_18814);
or U24313 (N_24313,N_18588,N_18824);
xor U24314 (N_24314,N_18650,N_15377);
nor U24315 (N_24315,N_16470,N_17024);
nand U24316 (N_24316,N_16224,N_17150);
xnor U24317 (N_24317,N_16445,N_16978);
and U24318 (N_24318,N_16039,N_18065);
or U24319 (N_24319,N_16336,N_19410);
and U24320 (N_24320,N_15361,N_18857);
nand U24321 (N_24321,N_19040,N_16715);
nand U24322 (N_24322,N_16426,N_17056);
xor U24323 (N_24323,N_18604,N_15556);
nand U24324 (N_24324,N_15599,N_18126);
nand U24325 (N_24325,N_16580,N_18112);
or U24326 (N_24326,N_19777,N_15805);
xor U24327 (N_24327,N_16824,N_17109);
xor U24328 (N_24328,N_17850,N_19353);
nand U24329 (N_24329,N_15178,N_16472);
xnor U24330 (N_24330,N_18740,N_19851);
and U24331 (N_24331,N_18012,N_19391);
nor U24332 (N_24332,N_15303,N_15654);
xnor U24333 (N_24333,N_16421,N_15431);
nor U24334 (N_24334,N_15458,N_18374);
or U24335 (N_24335,N_19526,N_18476);
nand U24336 (N_24336,N_16183,N_15966);
nor U24337 (N_24337,N_18440,N_15086);
nor U24338 (N_24338,N_18842,N_18983);
nor U24339 (N_24339,N_18219,N_18064);
xor U24340 (N_24340,N_16260,N_17402);
nand U24341 (N_24341,N_17329,N_16980);
xor U24342 (N_24342,N_18083,N_18898);
nand U24343 (N_24343,N_15076,N_19750);
and U24344 (N_24344,N_19432,N_16650);
or U24345 (N_24345,N_18035,N_16595);
or U24346 (N_24346,N_15212,N_17776);
nor U24347 (N_24347,N_15464,N_17674);
or U24348 (N_24348,N_19393,N_19982);
xnor U24349 (N_24349,N_19959,N_18389);
or U24350 (N_24350,N_19946,N_19249);
and U24351 (N_24351,N_18265,N_16709);
nand U24352 (N_24352,N_15509,N_17585);
and U24353 (N_24353,N_16432,N_18828);
nand U24354 (N_24354,N_15885,N_15921);
nand U24355 (N_24355,N_16848,N_15939);
nand U24356 (N_24356,N_17760,N_18255);
nor U24357 (N_24357,N_17500,N_16045);
nand U24358 (N_24358,N_19706,N_15121);
and U24359 (N_24359,N_17878,N_18867);
and U24360 (N_24360,N_17668,N_15432);
nor U24361 (N_24361,N_19043,N_19757);
or U24362 (N_24362,N_17203,N_15023);
nand U24363 (N_24363,N_19548,N_17843);
or U24364 (N_24364,N_17738,N_19760);
xor U24365 (N_24365,N_16413,N_18437);
or U24366 (N_24366,N_16727,N_19863);
nor U24367 (N_24367,N_19440,N_16290);
and U24368 (N_24368,N_18825,N_17783);
nand U24369 (N_24369,N_15981,N_16293);
nor U24370 (N_24370,N_15371,N_15863);
nor U24371 (N_24371,N_18852,N_15945);
or U24372 (N_24372,N_18986,N_16648);
xor U24373 (N_24373,N_18134,N_17111);
and U24374 (N_24374,N_18913,N_18859);
xnor U24375 (N_24375,N_16513,N_17145);
and U24376 (N_24376,N_15410,N_19273);
and U24377 (N_24377,N_19638,N_18627);
and U24378 (N_24378,N_18114,N_15084);
or U24379 (N_24379,N_18683,N_17976);
nor U24380 (N_24380,N_16441,N_18188);
or U24381 (N_24381,N_15965,N_19090);
nor U24382 (N_24382,N_16527,N_18807);
xor U24383 (N_24383,N_17430,N_16441);
and U24384 (N_24384,N_16477,N_15696);
xnor U24385 (N_24385,N_19055,N_16666);
or U24386 (N_24386,N_18071,N_16771);
xor U24387 (N_24387,N_18567,N_17607);
and U24388 (N_24388,N_19101,N_18695);
nor U24389 (N_24389,N_18358,N_16504);
or U24390 (N_24390,N_18437,N_16190);
nor U24391 (N_24391,N_19271,N_17785);
or U24392 (N_24392,N_16507,N_16794);
nor U24393 (N_24393,N_17328,N_18955);
nand U24394 (N_24394,N_16884,N_15204);
nor U24395 (N_24395,N_19748,N_19690);
nand U24396 (N_24396,N_19825,N_17192);
xor U24397 (N_24397,N_18527,N_18023);
nor U24398 (N_24398,N_18569,N_19043);
xnor U24399 (N_24399,N_15254,N_19777);
nor U24400 (N_24400,N_15815,N_17178);
nor U24401 (N_24401,N_17246,N_16422);
or U24402 (N_24402,N_15756,N_15064);
nor U24403 (N_24403,N_18692,N_15334);
xnor U24404 (N_24404,N_19709,N_16662);
nand U24405 (N_24405,N_18984,N_16997);
nor U24406 (N_24406,N_19397,N_15196);
nand U24407 (N_24407,N_15219,N_16164);
or U24408 (N_24408,N_15710,N_19138);
and U24409 (N_24409,N_19917,N_15976);
xnor U24410 (N_24410,N_15343,N_16345);
or U24411 (N_24411,N_18014,N_19173);
nor U24412 (N_24412,N_19857,N_19391);
and U24413 (N_24413,N_19093,N_15248);
or U24414 (N_24414,N_17184,N_19091);
nand U24415 (N_24415,N_18094,N_18595);
and U24416 (N_24416,N_17860,N_18372);
and U24417 (N_24417,N_17358,N_17471);
or U24418 (N_24418,N_17904,N_15455);
or U24419 (N_24419,N_19361,N_15489);
and U24420 (N_24420,N_16362,N_16373);
and U24421 (N_24421,N_15952,N_15236);
xnor U24422 (N_24422,N_18066,N_15642);
xor U24423 (N_24423,N_17113,N_15797);
and U24424 (N_24424,N_16566,N_15059);
nor U24425 (N_24425,N_16380,N_17753);
nand U24426 (N_24426,N_15738,N_17943);
and U24427 (N_24427,N_15287,N_17842);
and U24428 (N_24428,N_17967,N_18324);
or U24429 (N_24429,N_17430,N_17592);
nor U24430 (N_24430,N_15794,N_17192);
or U24431 (N_24431,N_15468,N_17208);
xor U24432 (N_24432,N_17709,N_19062);
or U24433 (N_24433,N_18134,N_18390);
and U24434 (N_24434,N_19628,N_18645);
xor U24435 (N_24435,N_19616,N_15586);
nand U24436 (N_24436,N_17332,N_17688);
nor U24437 (N_24437,N_18558,N_17973);
or U24438 (N_24438,N_15841,N_18306);
nor U24439 (N_24439,N_16972,N_18596);
or U24440 (N_24440,N_18577,N_17009);
nand U24441 (N_24441,N_19535,N_18101);
and U24442 (N_24442,N_17085,N_19448);
nand U24443 (N_24443,N_15535,N_19325);
and U24444 (N_24444,N_15668,N_17060);
nor U24445 (N_24445,N_19542,N_18120);
xor U24446 (N_24446,N_17421,N_16155);
nand U24447 (N_24447,N_19076,N_16242);
nand U24448 (N_24448,N_16884,N_19193);
nor U24449 (N_24449,N_15508,N_17817);
and U24450 (N_24450,N_18086,N_18107);
nor U24451 (N_24451,N_16487,N_16497);
xnor U24452 (N_24452,N_18736,N_18978);
xor U24453 (N_24453,N_19534,N_19673);
nor U24454 (N_24454,N_15245,N_15771);
xnor U24455 (N_24455,N_19296,N_19702);
xor U24456 (N_24456,N_19079,N_18122);
nor U24457 (N_24457,N_16789,N_15382);
or U24458 (N_24458,N_15188,N_17778);
nor U24459 (N_24459,N_19571,N_19501);
and U24460 (N_24460,N_17640,N_18150);
and U24461 (N_24461,N_17704,N_17162);
nor U24462 (N_24462,N_15407,N_18292);
nand U24463 (N_24463,N_16112,N_16284);
nand U24464 (N_24464,N_17821,N_15763);
nor U24465 (N_24465,N_18435,N_19485);
or U24466 (N_24466,N_16887,N_19895);
and U24467 (N_24467,N_17449,N_19856);
nand U24468 (N_24468,N_15884,N_15702);
nor U24469 (N_24469,N_18593,N_15242);
nor U24470 (N_24470,N_17931,N_16091);
xor U24471 (N_24471,N_15026,N_16894);
or U24472 (N_24472,N_17451,N_15700);
and U24473 (N_24473,N_17300,N_19831);
or U24474 (N_24474,N_18282,N_19841);
and U24475 (N_24475,N_16039,N_18390);
nand U24476 (N_24476,N_19470,N_15040);
nor U24477 (N_24477,N_17722,N_16294);
nand U24478 (N_24478,N_18622,N_18841);
nor U24479 (N_24479,N_19867,N_16305);
and U24480 (N_24480,N_18035,N_17277);
or U24481 (N_24481,N_19008,N_16105);
and U24482 (N_24482,N_19975,N_16992);
nor U24483 (N_24483,N_19144,N_17027);
and U24484 (N_24484,N_15718,N_18933);
nand U24485 (N_24485,N_18591,N_18308);
nand U24486 (N_24486,N_19795,N_18112);
xor U24487 (N_24487,N_18550,N_16832);
and U24488 (N_24488,N_19270,N_16989);
or U24489 (N_24489,N_16719,N_18824);
nand U24490 (N_24490,N_17387,N_19783);
nand U24491 (N_24491,N_19551,N_17370);
nor U24492 (N_24492,N_18140,N_15599);
or U24493 (N_24493,N_17691,N_17339);
nor U24494 (N_24494,N_16838,N_16227);
and U24495 (N_24495,N_18562,N_17083);
nand U24496 (N_24496,N_15439,N_18966);
xor U24497 (N_24497,N_16505,N_18335);
or U24498 (N_24498,N_17747,N_16358);
or U24499 (N_24499,N_19697,N_19903);
and U24500 (N_24500,N_16056,N_17084);
and U24501 (N_24501,N_18496,N_19059);
nor U24502 (N_24502,N_16131,N_18646);
nor U24503 (N_24503,N_15471,N_18484);
nand U24504 (N_24504,N_15581,N_17173);
or U24505 (N_24505,N_19576,N_16037);
xor U24506 (N_24506,N_15104,N_16504);
nand U24507 (N_24507,N_17873,N_17273);
and U24508 (N_24508,N_15775,N_18182);
and U24509 (N_24509,N_19196,N_17041);
or U24510 (N_24510,N_18435,N_17746);
and U24511 (N_24511,N_17645,N_15347);
nand U24512 (N_24512,N_19671,N_18481);
xor U24513 (N_24513,N_18059,N_19829);
xnor U24514 (N_24514,N_15844,N_15703);
nand U24515 (N_24515,N_16277,N_17950);
or U24516 (N_24516,N_16686,N_15677);
xnor U24517 (N_24517,N_19290,N_19514);
and U24518 (N_24518,N_16942,N_16101);
and U24519 (N_24519,N_18567,N_17915);
and U24520 (N_24520,N_15088,N_16986);
and U24521 (N_24521,N_19859,N_17032);
or U24522 (N_24522,N_15878,N_19176);
or U24523 (N_24523,N_15940,N_18094);
nand U24524 (N_24524,N_19202,N_15085);
nor U24525 (N_24525,N_15213,N_15207);
nand U24526 (N_24526,N_18539,N_16564);
nor U24527 (N_24527,N_19439,N_16827);
and U24528 (N_24528,N_17315,N_19984);
and U24529 (N_24529,N_16628,N_19936);
and U24530 (N_24530,N_17346,N_16684);
or U24531 (N_24531,N_16090,N_18101);
xor U24532 (N_24532,N_16597,N_16353);
and U24533 (N_24533,N_18030,N_18590);
nand U24534 (N_24534,N_16831,N_19688);
xor U24535 (N_24535,N_16484,N_18333);
nand U24536 (N_24536,N_18591,N_19030);
xor U24537 (N_24537,N_16276,N_18362);
xnor U24538 (N_24538,N_19950,N_15899);
or U24539 (N_24539,N_16204,N_15336);
nand U24540 (N_24540,N_18169,N_17917);
nor U24541 (N_24541,N_18098,N_18006);
nand U24542 (N_24542,N_17214,N_15503);
nand U24543 (N_24543,N_17002,N_17816);
nor U24544 (N_24544,N_17001,N_18810);
or U24545 (N_24545,N_15303,N_16189);
xor U24546 (N_24546,N_17806,N_15017);
or U24547 (N_24547,N_17556,N_15715);
nand U24548 (N_24548,N_15447,N_15266);
nor U24549 (N_24549,N_18756,N_19365);
nor U24550 (N_24550,N_16822,N_15062);
or U24551 (N_24551,N_17996,N_18131);
nor U24552 (N_24552,N_15089,N_16964);
or U24553 (N_24553,N_19400,N_18211);
nand U24554 (N_24554,N_16118,N_18132);
nand U24555 (N_24555,N_16844,N_16626);
or U24556 (N_24556,N_19932,N_16346);
or U24557 (N_24557,N_16061,N_15514);
and U24558 (N_24558,N_15105,N_18914);
nand U24559 (N_24559,N_16480,N_16965);
xor U24560 (N_24560,N_15563,N_16595);
nor U24561 (N_24561,N_19908,N_16822);
nor U24562 (N_24562,N_19614,N_17469);
nor U24563 (N_24563,N_17563,N_15552);
and U24564 (N_24564,N_18542,N_19787);
or U24565 (N_24565,N_18997,N_19545);
nor U24566 (N_24566,N_18763,N_17984);
xor U24567 (N_24567,N_19509,N_16540);
xor U24568 (N_24568,N_17885,N_17218);
xor U24569 (N_24569,N_19601,N_19179);
or U24570 (N_24570,N_17137,N_16372);
nand U24571 (N_24571,N_17215,N_15050);
nor U24572 (N_24572,N_19985,N_17982);
nor U24573 (N_24573,N_17102,N_17818);
nor U24574 (N_24574,N_16740,N_17389);
xnor U24575 (N_24575,N_16664,N_17512);
nand U24576 (N_24576,N_17099,N_16446);
or U24577 (N_24577,N_18951,N_18858);
nor U24578 (N_24578,N_18260,N_16631);
xnor U24579 (N_24579,N_16525,N_16980);
nor U24580 (N_24580,N_18564,N_17204);
nand U24581 (N_24581,N_16652,N_19618);
and U24582 (N_24582,N_18151,N_16034);
xor U24583 (N_24583,N_19561,N_16830);
nand U24584 (N_24584,N_16495,N_17568);
nor U24585 (N_24585,N_15047,N_15799);
xnor U24586 (N_24586,N_19198,N_15618);
or U24587 (N_24587,N_17637,N_18542);
and U24588 (N_24588,N_15537,N_19780);
nor U24589 (N_24589,N_18847,N_16126);
nand U24590 (N_24590,N_19584,N_18945);
or U24591 (N_24591,N_15458,N_16791);
xor U24592 (N_24592,N_18585,N_17249);
or U24593 (N_24593,N_15708,N_18894);
nand U24594 (N_24594,N_19994,N_18427);
xor U24595 (N_24595,N_16264,N_19759);
and U24596 (N_24596,N_18229,N_19804);
or U24597 (N_24597,N_18413,N_19659);
xor U24598 (N_24598,N_17708,N_16758);
and U24599 (N_24599,N_16379,N_17785);
xor U24600 (N_24600,N_17413,N_18694);
xnor U24601 (N_24601,N_18070,N_16454);
and U24602 (N_24602,N_15692,N_15092);
and U24603 (N_24603,N_16668,N_18296);
nand U24604 (N_24604,N_15597,N_17784);
and U24605 (N_24605,N_17813,N_19522);
xor U24606 (N_24606,N_18314,N_18751);
nor U24607 (N_24607,N_15772,N_18196);
nand U24608 (N_24608,N_16151,N_16591);
nand U24609 (N_24609,N_18262,N_18833);
xor U24610 (N_24610,N_19867,N_17930);
and U24611 (N_24611,N_16371,N_18923);
nor U24612 (N_24612,N_16839,N_17510);
xnor U24613 (N_24613,N_18221,N_18808);
nand U24614 (N_24614,N_15358,N_16399);
xor U24615 (N_24615,N_15625,N_19847);
or U24616 (N_24616,N_17338,N_15604);
nand U24617 (N_24617,N_17080,N_16421);
nand U24618 (N_24618,N_15972,N_15355);
xnor U24619 (N_24619,N_19288,N_18314);
nand U24620 (N_24620,N_16577,N_18109);
nor U24621 (N_24621,N_16201,N_19054);
or U24622 (N_24622,N_15979,N_17560);
nor U24623 (N_24623,N_19200,N_18191);
and U24624 (N_24624,N_17457,N_19522);
xnor U24625 (N_24625,N_19535,N_16606);
xor U24626 (N_24626,N_19868,N_15985);
xor U24627 (N_24627,N_15845,N_19541);
nor U24628 (N_24628,N_15526,N_18452);
or U24629 (N_24629,N_16452,N_18572);
or U24630 (N_24630,N_19408,N_17375);
and U24631 (N_24631,N_15690,N_16183);
xnor U24632 (N_24632,N_15990,N_17014);
nand U24633 (N_24633,N_19014,N_16793);
xnor U24634 (N_24634,N_15711,N_18404);
and U24635 (N_24635,N_18727,N_18855);
nor U24636 (N_24636,N_16988,N_18807);
xnor U24637 (N_24637,N_18227,N_18154);
nor U24638 (N_24638,N_16151,N_18646);
or U24639 (N_24639,N_15605,N_19139);
and U24640 (N_24640,N_19282,N_19400);
nor U24641 (N_24641,N_15604,N_17248);
nor U24642 (N_24642,N_15324,N_18956);
or U24643 (N_24643,N_17863,N_18360);
nand U24644 (N_24644,N_16278,N_15734);
or U24645 (N_24645,N_15007,N_17280);
nand U24646 (N_24646,N_18381,N_17935);
or U24647 (N_24647,N_17426,N_16399);
xnor U24648 (N_24648,N_18739,N_15017);
or U24649 (N_24649,N_19151,N_19778);
xor U24650 (N_24650,N_16941,N_15309);
xnor U24651 (N_24651,N_19343,N_17308);
nor U24652 (N_24652,N_19024,N_17276);
nor U24653 (N_24653,N_19526,N_15686);
and U24654 (N_24654,N_17268,N_16979);
xor U24655 (N_24655,N_15292,N_18588);
and U24656 (N_24656,N_18515,N_16476);
nand U24657 (N_24657,N_19267,N_16406);
and U24658 (N_24658,N_17022,N_18137);
xnor U24659 (N_24659,N_17587,N_15580);
and U24660 (N_24660,N_16569,N_17062);
or U24661 (N_24661,N_18561,N_18398);
and U24662 (N_24662,N_16794,N_17510);
xnor U24663 (N_24663,N_16013,N_15778);
nor U24664 (N_24664,N_18636,N_17480);
nand U24665 (N_24665,N_17361,N_18678);
nand U24666 (N_24666,N_17188,N_17251);
or U24667 (N_24667,N_16589,N_15867);
or U24668 (N_24668,N_16861,N_17316);
xnor U24669 (N_24669,N_15951,N_18934);
or U24670 (N_24670,N_16460,N_19157);
nand U24671 (N_24671,N_17760,N_17731);
or U24672 (N_24672,N_18741,N_19029);
nor U24673 (N_24673,N_18127,N_17819);
or U24674 (N_24674,N_18596,N_16223);
or U24675 (N_24675,N_19293,N_19630);
nand U24676 (N_24676,N_17994,N_15702);
nand U24677 (N_24677,N_16890,N_18568);
xnor U24678 (N_24678,N_19587,N_16878);
and U24679 (N_24679,N_16589,N_18716);
or U24680 (N_24680,N_19850,N_18711);
xor U24681 (N_24681,N_19849,N_17575);
nor U24682 (N_24682,N_16855,N_17365);
nand U24683 (N_24683,N_15378,N_19261);
or U24684 (N_24684,N_16144,N_15575);
or U24685 (N_24685,N_18130,N_17831);
xor U24686 (N_24686,N_19570,N_17194);
nand U24687 (N_24687,N_18121,N_18506);
and U24688 (N_24688,N_16065,N_15263);
nand U24689 (N_24689,N_17781,N_18681);
nand U24690 (N_24690,N_15994,N_16707);
nand U24691 (N_24691,N_18558,N_16759);
or U24692 (N_24692,N_19163,N_17625);
and U24693 (N_24693,N_18460,N_16592);
xnor U24694 (N_24694,N_15687,N_16786);
nor U24695 (N_24695,N_18649,N_16450);
nand U24696 (N_24696,N_19281,N_19644);
and U24697 (N_24697,N_16370,N_19858);
xnor U24698 (N_24698,N_17370,N_17627);
and U24699 (N_24699,N_18939,N_15930);
xor U24700 (N_24700,N_16834,N_16770);
or U24701 (N_24701,N_19283,N_19017);
xor U24702 (N_24702,N_17363,N_18374);
nor U24703 (N_24703,N_18456,N_17273);
xor U24704 (N_24704,N_17214,N_18016);
xnor U24705 (N_24705,N_16779,N_17089);
and U24706 (N_24706,N_17717,N_18198);
and U24707 (N_24707,N_17076,N_19513);
or U24708 (N_24708,N_15038,N_16297);
or U24709 (N_24709,N_16692,N_17884);
nand U24710 (N_24710,N_17757,N_17966);
nand U24711 (N_24711,N_18911,N_18345);
or U24712 (N_24712,N_18462,N_19198);
nor U24713 (N_24713,N_16338,N_17913);
and U24714 (N_24714,N_19646,N_19096);
xnor U24715 (N_24715,N_15910,N_18445);
xor U24716 (N_24716,N_19208,N_16007);
nor U24717 (N_24717,N_18946,N_16103);
and U24718 (N_24718,N_17951,N_18606);
xor U24719 (N_24719,N_19487,N_16238);
or U24720 (N_24720,N_19334,N_16126);
xor U24721 (N_24721,N_15886,N_16372);
nand U24722 (N_24722,N_15071,N_18503);
nor U24723 (N_24723,N_17839,N_19905);
or U24724 (N_24724,N_15055,N_16029);
nand U24725 (N_24725,N_19230,N_15422);
xnor U24726 (N_24726,N_15772,N_16634);
xor U24727 (N_24727,N_15318,N_17283);
nand U24728 (N_24728,N_19713,N_16283);
xnor U24729 (N_24729,N_19864,N_16093);
nor U24730 (N_24730,N_18269,N_17599);
nor U24731 (N_24731,N_15663,N_17942);
or U24732 (N_24732,N_15599,N_19756);
nor U24733 (N_24733,N_16694,N_19721);
xor U24734 (N_24734,N_16900,N_17034);
and U24735 (N_24735,N_18387,N_16890);
or U24736 (N_24736,N_19629,N_16950);
nand U24737 (N_24737,N_17098,N_18795);
xor U24738 (N_24738,N_15608,N_18188);
nand U24739 (N_24739,N_19859,N_17832);
or U24740 (N_24740,N_17465,N_17525);
xor U24741 (N_24741,N_15428,N_15744);
nor U24742 (N_24742,N_19951,N_17740);
nand U24743 (N_24743,N_17344,N_18403);
xnor U24744 (N_24744,N_16484,N_17215);
nand U24745 (N_24745,N_16058,N_18598);
and U24746 (N_24746,N_18657,N_18865);
nand U24747 (N_24747,N_18269,N_15474);
nand U24748 (N_24748,N_16962,N_16719);
nor U24749 (N_24749,N_18769,N_15981);
or U24750 (N_24750,N_18241,N_17628);
nor U24751 (N_24751,N_16301,N_19120);
and U24752 (N_24752,N_18041,N_17630);
and U24753 (N_24753,N_19036,N_18175);
nand U24754 (N_24754,N_19774,N_19747);
nand U24755 (N_24755,N_17531,N_17610);
xor U24756 (N_24756,N_19530,N_18410);
nand U24757 (N_24757,N_15892,N_19647);
nand U24758 (N_24758,N_19035,N_17174);
or U24759 (N_24759,N_15324,N_19372);
xor U24760 (N_24760,N_19380,N_19655);
xor U24761 (N_24761,N_18410,N_17769);
nor U24762 (N_24762,N_16747,N_18858);
and U24763 (N_24763,N_19516,N_15293);
nand U24764 (N_24764,N_18755,N_18092);
xnor U24765 (N_24765,N_17631,N_18455);
nor U24766 (N_24766,N_18889,N_18382);
or U24767 (N_24767,N_15343,N_17312);
xnor U24768 (N_24768,N_17395,N_17695);
and U24769 (N_24769,N_17407,N_16421);
or U24770 (N_24770,N_16692,N_18317);
and U24771 (N_24771,N_18811,N_19742);
nand U24772 (N_24772,N_19049,N_16349);
xor U24773 (N_24773,N_15741,N_15593);
xnor U24774 (N_24774,N_19767,N_16424);
nor U24775 (N_24775,N_19459,N_17902);
nand U24776 (N_24776,N_19856,N_17611);
nor U24777 (N_24777,N_18049,N_17327);
nand U24778 (N_24778,N_15061,N_17187);
and U24779 (N_24779,N_18328,N_19733);
nand U24780 (N_24780,N_18650,N_18265);
xnor U24781 (N_24781,N_18308,N_18642);
and U24782 (N_24782,N_15083,N_18897);
nand U24783 (N_24783,N_18837,N_18322);
and U24784 (N_24784,N_15373,N_15699);
nor U24785 (N_24785,N_19551,N_15441);
nor U24786 (N_24786,N_17409,N_15132);
and U24787 (N_24787,N_18337,N_17040);
nand U24788 (N_24788,N_17144,N_17581);
xor U24789 (N_24789,N_19023,N_19161);
and U24790 (N_24790,N_19321,N_15501);
nand U24791 (N_24791,N_18127,N_18554);
xnor U24792 (N_24792,N_19482,N_18962);
nand U24793 (N_24793,N_15922,N_15649);
and U24794 (N_24794,N_15010,N_17789);
nor U24795 (N_24795,N_17651,N_16201);
or U24796 (N_24796,N_19519,N_15582);
nor U24797 (N_24797,N_19662,N_17359);
nor U24798 (N_24798,N_16885,N_16900);
nor U24799 (N_24799,N_19961,N_17997);
nor U24800 (N_24800,N_16107,N_17619);
nand U24801 (N_24801,N_16362,N_15638);
nor U24802 (N_24802,N_17417,N_17089);
and U24803 (N_24803,N_15148,N_18941);
xor U24804 (N_24804,N_16357,N_19568);
xor U24805 (N_24805,N_18129,N_18308);
or U24806 (N_24806,N_18748,N_16729);
nand U24807 (N_24807,N_19654,N_16000);
and U24808 (N_24808,N_17620,N_15745);
xor U24809 (N_24809,N_18218,N_15684);
and U24810 (N_24810,N_17485,N_16569);
nand U24811 (N_24811,N_19582,N_17819);
and U24812 (N_24812,N_16102,N_17138);
or U24813 (N_24813,N_18561,N_16286);
nor U24814 (N_24814,N_18203,N_16640);
nor U24815 (N_24815,N_16218,N_19659);
or U24816 (N_24816,N_16316,N_16081);
nand U24817 (N_24817,N_19863,N_15653);
and U24818 (N_24818,N_18765,N_16153);
and U24819 (N_24819,N_17025,N_18863);
nand U24820 (N_24820,N_15834,N_17135);
xor U24821 (N_24821,N_17731,N_19635);
and U24822 (N_24822,N_17124,N_15916);
nor U24823 (N_24823,N_18693,N_16749);
xor U24824 (N_24824,N_15061,N_16977);
nand U24825 (N_24825,N_19937,N_18512);
or U24826 (N_24826,N_18053,N_16767);
nand U24827 (N_24827,N_18891,N_19292);
nand U24828 (N_24828,N_16828,N_18476);
nor U24829 (N_24829,N_17015,N_17503);
or U24830 (N_24830,N_16183,N_15557);
xnor U24831 (N_24831,N_16843,N_19162);
nor U24832 (N_24832,N_19882,N_18751);
or U24833 (N_24833,N_16180,N_16232);
nor U24834 (N_24834,N_17875,N_18300);
nor U24835 (N_24835,N_18257,N_16173);
nor U24836 (N_24836,N_16638,N_16808);
nand U24837 (N_24837,N_17328,N_15772);
and U24838 (N_24838,N_17149,N_16748);
nor U24839 (N_24839,N_16362,N_15450);
and U24840 (N_24840,N_15558,N_16537);
and U24841 (N_24841,N_18839,N_17457);
nor U24842 (N_24842,N_18416,N_19511);
and U24843 (N_24843,N_15874,N_17738);
or U24844 (N_24844,N_16201,N_15141);
or U24845 (N_24845,N_16462,N_17257);
nor U24846 (N_24846,N_18795,N_16510);
and U24847 (N_24847,N_15580,N_18598);
or U24848 (N_24848,N_16998,N_15894);
nand U24849 (N_24849,N_15343,N_17622);
or U24850 (N_24850,N_15129,N_15744);
nand U24851 (N_24851,N_17200,N_16871);
nor U24852 (N_24852,N_19494,N_17512);
and U24853 (N_24853,N_19234,N_16727);
and U24854 (N_24854,N_19649,N_19803);
nor U24855 (N_24855,N_16255,N_17307);
and U24856 (N_24856,N_17994,N_16293);
xnor U24857 (N_24857,N_18826,N_19391);
nor U24858 (N_24858,N_18243,N_17015);
nor U24859 (N_24859,N_19208,N_17516);
nand U24860 (N_24860,N_19325,N_16269);
nor U24861 (N_24861,N_19745,N_17340);
xor U24862 (N_24862,N_19866,N_15086);
or U24863 (N_24863,N_19037,N_15407);
nor U24864 (N_24864,N_16518,N_19520);
nand U24865 (N_24865,N_18998,N_16775);
or U24866 (N_24866,N_19604,N_19023);
nor U24867 (N_24867,N_16769,N_16835);
xnor U24868 (N_24868,N_16890,N_16373);
and U24869 (N_24869,N_17266,N_16092);
xnor U24870 (N_24870,N_18354,N_18770);
and U24871 (N_24871,N_17338,N_19298);
nand U24872 (N_24872,N_17143,N_16537);
nand U24873 (N_24873,N_18501,N_17070);
xnor U24874 (N_24874,N_17983,N_19763);
nor U24875 (N_24875,N_19450,N_17730);
nor U24876 (N_24876,N_17146,N_17110);
nand U24877 (N_24877,N_17264,N_19412);
nor U24878 (N_24878,N_15533,N_17011);
and U24879 (N_24879,N_18352,N_15835);
or U24880 (N_24880,N_15051,N_15957);
nand U24881 (N_24881,N_15255,N_15562);
nor U24882 (N_24882,N_15745,N_19687);
and U24883 (N_24883,N_18231,N_19610);
nand U24884 (N_24884,N_19340,N_17994);
xnor U24885 (N_24885,N_15303,N_16975);
nand U24886 (N_24886,N_17448,N_16925);
nand U24887 (N_24887,N_16918,N_17927);
nor U24888 (N_24888,N_15456,N_18822);
or U24889 (N_24889,N_17821,N_18550);
or U24890 (N_24890,N_17260,N_17632);
xor U24891 (N_24891,N_15753,N_15687);
or U24892 (N_24892,N_17395,N_15557);
xnor U24893 (N_24893,N_16067,N_15347);
nand U24894 (N_24894,N_16904,N_19836);
nand U24895 (N_24895,N_17161,N_19812);
nand U24896 (N_24896,N_19486,N_16779);
xnor U24897 (N_24897,N_17538,N_16800);
and U24898 (N_24898,N_19813,N_16974);
and U24899 (N_24899,N_18976,N_17491);
nand U24900 (N_24900,N_15576,N_15931);
nand U24901 (N_24901,N_15534,N_16909);
nand U24902 (N_24902,N_16043,N_19742);
nand U24903 (N_24903,N_18212,N_15495);
nand U24904 (N_24904,N_17753,N_15345);
or U24905 (N_24905,N_15619,N_17905);
xor U24906 (N_24906,N_17284,N_19515);
or U24907 (N_24907,N_15725,N_18918);
xor U24908 (N_24908,N_15499,N_17412);
and U24909 (N_24909,N_16982,N_15810);
nor U24910 (N_24910,N_15590,N_19057);
nor U24911 (N_24911,N_19048,N_17683);
and U24912 (N_24912,N_19458,N_15121);
and U24913 (N_24913,N_19321,N_16964);
nor U24914 (N_24914,N_15651,N_17069);
xnor U24915 (N_24915,N_15032,N_16421);
or U24916 (N_24916,N_16214,N_18994);
nor U24917 (N_24917,N_16399,N_17349);
nor U24918 (N_24918,N_17882,N_15895);
xnor U24919 (N_24919,N_19867,N_15961);
or U24920 (N_24920,N_18856,N_17231);
nand U24921 (N_24921,N_19398,N_17402);
and U24922 (N_24922,N_17167,N_18630);
xnor U24923 (N_24923,N_15295,N_17351);
or U24924 (N_24924,N_15971,N_19056);
nor U24925 (N_24925,N_19336,N_19091);
nand U24926 (N_24926,N_15583,N_18087);
xnor U24927 (N_24927,N_15294,N_19678);
nand U24928 (N_24928,N_16375,N_16055);
xor U24929 (N_24929,N_16368,N_18025);
and U24930 (N_24930,N_16369,N_19954);
and U24931 (N_24931,N_19119,N_15265);
or U24932 (N_24932,N_16874,N_18814);
xnor U24933 (N_24933,N_19414,N_18143);
nand U24934 (N_24934,N_15164,N_19534);
nor U24935 (N_24935,N_15465,N_15034);
xnor U24936 (N_24936,N_15599,N_18886);
xor U24937 (N_24937,N_15957,N_18733);
or U24938 (N_24938,N_16052,N_15964);
xor U24939 (N_24939,N_18019,N_15224);
xor U24940 (N_24940,N_16243,N_18395);
or U24941 (N_24941,N_19879,N_16972);
nand U24942 (N_24942,N_15534,N_15844);
or U24943 (N_24943,N_16276,N_19462);
nand U24944 (N_24944,N_16762,N_16431);
or U24945 (N_24945,N_16557,N_15525);
or U24946 (N_24946,N_18420,N_17680);
or U24947 (N_24947,N_15495,N_19741);
nand U24948 (N_24948,N_15435,N_16978);
or U24949 (N_24949,N_15862,N_19880);
xnor U24950 (N_24950,N_15316,N_18375);
or U24951 (N_24951,N_15064,N_16654);
nor U24952 (N_24952,N_19945,N_16581);
nand U24953 (N_24953,N_19104,N_17172);
nand U24954 (N_24954,N_17651,N_17986);
nand U24955 (N_24955,N_18956,N_19277);
and U24956 (N_24956,N_15284,N_19011);
nor U24957 (N_24957,N_16216,N_19618);
nand U24958 (N_24958,N_17641,N_18591);
xor U24959 (N_24959,N_17548,N_16304);
nand U24960 (N_24960,N_18084,N_17564);
xor U24961 (N_24961,N_16626,N_18857);
nand U24962 (N_24962,N_17616,N_16824);
or U24963 (N_24963,N_19085,N_16721);
nor U24964 (N_24964,N_18269,N_19898);
nor U24965 (N_24965,N_16356,N_15421);
or U24966 (N_24966,N_16753,N_15339);
nor U24967 (N_24967,N_15647,N_19708);
or U24968 (N_24968,N_19322,N_19207);
or U24969 (N_24969,N_15947,N_15452);
and U24970 (N_24970,N_18809,N_19477);
xnor U24971 (N_24971,N_16553,N_19867);
or U24972 (N_24972,N_18834,N_15863);
or U24973 (N_24973,N_16028,N_15851);
or U24974 (N_24974,N_15841,N_18730);
xnor U24975 (N_24975,N_18579,N_15831);
and U24976 (N_24976,N_19683,N_18931);
xnor U24977 (N_24977,N_18189,N_18233);
or U24978 (N_24978,N_15539,N_17613);
or U24979 (N_24979,N_16495,N_18713);
nand U24980 (N_24980,N_17527,N_16802);
nor U24981 (N_24981,N_18836,N_17552);
xor U24982 (N_24982,N_19265,N_16848);
and U24983 (N_24983,N_18416,N_18498);
nand U24984 (N_24984,N_15528,N_15410);
xnor U24985 (N_24985,N_17605,N_18783);
nor U24986 (N_24986,N_19452,N_15677);
nor U24987 (N_24987,N_15074,N_19091);
nand U24988 (N_24988,N_18388,N_15502);
xor U24989 (N_24989,N_15573,N_15945);
nor U24990 (N_24990,N_17086,N_17401);
and U24991 (N_24991,N_19283,N_16429);
nand U24992 (N_24992,N_15505,N_16924);
nand U24993 (N_24993,N_18148,N_17127);
nand U24994 (N_24994,N_15268,N_15078);
nor U24995 (N_24995,N_18206,N_16088);
nand U24996 (N_24996,N_18845,N_19640);
nand U24997 (N_24997,N_15240,N_17955);
nand U24998 (N_24998,N_19230,N_17963);
and U24999 (N_24999,N_15153,N_15180);
nand UO_0 (O_0,N_22401,N_22693);
nor UO_1 (O_1,N_20147,N_24249);
or UO_2 (O_2,N_22407,N_20287);
or UO_3 (O_3,N_20776,N_23961);
nand UO_4 (O_4,N_22737,N_23695);
nand UO_5 (O_5,N_24472,N_21136);
nand UO_6 (O_6,N_24256,N_23095);
xnor UO_7 (O_7,N_24713,N_24737);
nor UO_8 (O_8,N_20394,N_23399);
nor UO_9 (O_9,N_23139,N_20915);
and UO_10 (O_10,N_22250,N_20340);
nand UO_11 (O_11,N_21260,N_20241);
nor UO_12 (O_12,N_22756,N_22220);
nand UO_13 (O_13,N_24418,N_24977);
nor UO_14 (O_14,N_21480,N_24185);
or UO_15 (O_15,N_20438,N_22070);
xnor UO_16 (O_16,N_22248,N_22919);
nand UO_17 (O_17,N_24123,N_20286);
xnor UO_18 (O_18,N_23799,N_21975);
nand UO_19 (O_19,N_23047,N_20977);
and UO_20 (O_20,N_24706,N_20827);
xor UO_21 (O_21,N_23432,N_22568);
or UO_22 (O_22,N_23062,N_22009);
and UO_23 (O_23,N_23573,N_22062);
nand UO_24 (O_24,N_20755,N_21861);
nor UO_25 (O_25,N_21345,N_23759);
xnor UO_26 (O_26,N_23328,N_23031);
nand UO_27 (O_27,N_22569,N_23692);
or UO_28 (O_28,N_20550,N_22365);
xnor UO_29 (O_29,N_21563,N_24881);
nand UO_30 (O_30,N_22322,N_24117);
and UO_31 (O_31,N_22409,N_22246);
xor UO_32 (O_32,N_24612,N_20597);
nor UO_33 (O_33,N_21380,N_20732);
nor UO_34 (O_34,N_21920,N_20861);
nor UO_35 (O_35,N_24459,N_21342);
xnor UO_36 (O_36,N_22271,N_20926);
and UO_37 (O_37,N_24153,N_24658);
xnor UO_38 (O_38,N_23669,N_23473);
nand UO_39 (O_39,N_23216,N_20001);
and UO_40 (O_40,N_22895,N_24986);
nand UO_41 (O_41,N_20969,N_23323);
xor UO_42 (O_42,N_20354,N_22635);
or UO_43 (O_43,N_23133,N_24481);
nand UO_44 (O_44,N_21019,N_23896);
or UO_45 (O_45,N_23395,N_21190);
nor UO_46 (O_46,N_20015,N_22889);
xor UO_47 (O_47,N_23276,N_21372);
and UO_48 (O_48,N_21403,N_22770);
xnor UO_49 (O_49,N_23373,N_21831);
nand UO_50 (O_50,N_20335,N_20898);
and UO_51 (O_51,N_21173,N_20822);
or UO_52 (O_52,N_23726,N_24885);
and UO_53 (O_53,N_24622,N_23618);
nor UO_54 (O_54,N_20355,N_23859);
nand UO_55 (O_55,N_23540,N_22544);
nand UO_56 (O_56,N_21691,N_21411);
xnor UO_57 (O_57,N_24944,N_23097);
and UO_58 (O_58,N_23592,N_23601);
xnor UO_59 (O_59,N_20906,N_21484);
nand UO_60 (O_60,N_21401,N_20874);
nor UO_61 (O_61,N_20965,N_22091);
nor UO_62 (O_62,N_21589,N_23583);
xnor UO_63 (O_63,N_22597,N_24184);
or UO_64 (O_64,N_21616,N_21745);
or UO_65 (O_65,N_20745,N_21517);
nand UO_66 (O_66,N_23390,N_23083);
nor UO_67 (O_67,N_22079,N_24815);
xnor UO_68 (O_68,N_22816,N_20256);
nor UO_69 (O_69,N_20139,N_24801);
nor UO_70 (O_70,N_20700,N_22982);
or UO_71 (O_71,N_24639,N_22236);
or UO_72 (O_72,N_21984,N_24397);
xor UO_73 (O_73,N_24679,N_22117);
or UO_74 (O_74,N_23679,N_20677);
nand UO_75 (O_75,N_21926,N_21894);
or UO_76 (O_76,N_23496,N_20150);
xor UO_77 (O_77,N_24112,N_24542);
xnor UO_78 (O_78,N_23306,N_22383);
xnor UO_79 (O_79,N_24191,N_24571);
or UO_80 (O_80,N_21117,N_21991);
or UO_81 (O_81,N_21358,N_21573);
or UO_82 (O_82,N_23534,N_24322);
nand UO_83 (O_83,N_23078,N_23713);
and UO_84 (O_84,N_20653,N_20123);
nand UO_85 (O_85,N_21317,N_20538);
xor UO_86 (O_86,N_23720,N_22791);
xor UO_87 (O_87,N_23998,N_21077);
and UO_88 (O_88,N_21516,N_20586);
or UO_89 (O_89,N_24309,N_23696);
xnor UO_90 (O_90,N_23449,N_20231);
nor UO_91 (O_91,N_20531,N_23146);
xnor UO_92 (O_92,N_21385,N_22461);
nor UO_93 (O_93,N_24467,N_23264);
or UO_94 (O_94,N_24029,N_23034);
xor UO_95 (O_95,N_22880,N_23552);
xnor UO_96 (O_96,N_20879,N_21614);
or UO_97 (O_97,N_23587,N_22538);
nor UO_98 (O_98,N_20963,N_20307);
and UO_99 (O_99,N_21112,N_20656);
xnor UO_100 (O_100,N_22267,N_22374);
and UO_101 (O_101,N_24246,N_23558);
nor UO_102 (O_102,N_22292,N_23008);
nor UO_103 (O_103,N_23671,N_23162);
or UO_104 (O_104,N_21125,N_24124);
nand UO_105 (O_105,N_22549,N_20048);
nor UO_106 (O_106,N_20130,N_24167);
or UO_107 (O_107,N_24279,N_20589);
xor UO_108 (O_108,N_23050,N_21650);
nand UO_109 (O_109,N_23820,N_22204);
and UO_110 (O_110,N_24891,N_20444);
nor UO_111 (O_111,N_22350,N_20659);
and UO_112 (O_112,N_21980,N_22475);
xnor UO_113 (O_113,N_23093,N_20931);
or UO_114 (O_114,N_20456,N_21545);
nand UO_115 (O_115,N_24704,N_24857);
nand UO_116 (O_116,N_21459,N_23379);
or UO_117 (O_117,N_20398,N_21715);
xor UO_118 (O_118,N_23983,N_22100);
and UO_119 (O_119,N_20506,N_20290);
and UO_120 (O_120,N_24513,N_23885);
or UO_121 (O_121,N_21554,N_20573);
nor UO_122 (O_122,N_20640,N_24060);
and UO_123 (O_123,N_22726,N_20493);
nor UO_124 (O_124,N_22139,N_24516);
xnor UO_125 (O_125,N_21449,N_23658);
or UO_126 (O_126,N_23833,N_21905);
or UO_127 (O_127,N_21096,N_21668);
or UO_128 (O_128,N_23974,N_20433);
and UO_129 (O_129,N_24861,N_24305);
xnor UO_130 (O_130,N_24973,N_24331);
nor UO_131 (O_131,N_22180,N_20187);
xnor UO_132 (O_132,N_23284,N_24217);
nand UO_133 (O_133,N_21731,N_23459);
nand UO_134 (O_134,N_21594,N_20577);
xnor UO_135 (O_135,N_24365,N_20804);
and UO_136 (O_136,N_21126,N_24209);
and UO_137 (O_137,N_22329,N_22964);
nand UO_138 (O_138,N_23074,N_24386);
xnor UO_139 (O_139,N_21597,N_23442);
and UO_140 (O_140,N_20948,N_23843);
nand UO_141 (O_141,N_24049,N_21038);
nor UO_142 (O_142,N_23653,N_21965);
and UO_143 (O_143,N_24489,N_24818);
xor UO_144 (O_144,N_20803,N_24719);
nand UO_145 (O_145,N_21321,N_23220);
xnor UO_146 (O_146,N_21999,N_24338);
and UO_147 (O_147,N_20556,N_21607);
nand UO_148 (O_148,N_22662,N_23588);
xnor UO_149 (O_149,N_20191,N_22525);
and UO_150 (O_150,N_24308,N_23982);
nand UO_151 (O_151,N_20784,N_22928);
xnor UO_152 (O_152,N_23438,N_22338);
or UO_153 (O_153,N_22053,N_23538);
xnor UO_154 (O_154,N_20013,N_22358);
nor UO_155 (O_155,N_23755,N_20571);
nor UO_156 (O_156,N_22438,N_20964);
or UO_157 (O_157,N_23064,N_22870);
nand UO_158 (O_158,N_20294,N_20759);
or UO_159 (O_159,N_24919,N_22171);
xnor UO_160 (O_160,N_20664,N_20734);
nor UO_161 (O_161,N_22650,N_22565);
and UO_162 (O_162,N_23965,N_21259);
nand UO_163 (O_163,N_22952,N_23141);
or UO_164 (O_164,N_20389,N_22611);
or UO_165 (O_165,N_20821,N_23925);
or UO_166 (O_166,N_21885,N_21893);
or UO_167 (O_167,N_21955,N_21307);
or UO_168 (O_168,N_22670,N_24884);
and UO_169 (O_169,N_22683,N_23582);
xnor UO_170 (O_170,N_20315,N_22480);
nand UO_171 (O_171,N_22205,N_20809);
nor UO_172 (O_172,N_23711,N_21870);
or UO_173 (O_173,N_23299,N_21237);
or UO_174 (O_174,N_22760,N_24187);
and UO_175 (O_175,N_23037,N_21532);
xnor UO_176 (O_176,N_22778,N_23955);
nand UO_177 (O_177,N_22231,N_24194);
nand UO_178 (O_178,N_23196,N_20660);
or UO_179 (O_179,N_24160,N_20635);
nor UO_180 (O_180,N_22467,N_24414);
or UO_181 (O_181,N_23836,N_24183);
nor UO_182 (O_182,N_21697,N_22768);
xnor UO_183 (O_183,N_21462,N_23949);
nand UO_184 (O_184,N_24528,N_23142);
and UO_185 (O_185,N_20682,N_20100);
xor UO_186 (O_186,N_23163,N_23404);
or UO_187 (O_187,N_21109,N_21193);
xnor UO_188 (O_188,N_24747,N_24053);
and UO_189 (O_189,N_20249,N_23173);
and UO_190 (O_190,N_22418,N_22061);
and UO_191 (O_191,N_22025,N_24450);
or UO_192 (O_192,N_20369,N_21337);
and UO_193 (O_193,N_23458,N_20869);
nor UO_194 (O_194,N_22107,N_20904);
xor UO_195 (O_195,N_20667,N_21579);
and UO_196 (O_196,N_21371,N_24054);
nand UO_197 (O_197,N_24549,N_22226);
nor UO_198 (O_198,N_20950,N_20328);
xnor UO_199 (O_199,N_21147,N_21601);
xnor UO_200 (O_200,N_23756,N_23474);
nand UO_201 (O_201,N_24255,N_20630);
and UO_202 (O_202,N_22798,N_23224);
nor UO_203 (O_203,N_21339,N_20975);
nor UO_204 (O_204,N_22188,N_20972);
nand UO_205 (O_205,N_21394,N_23780);
nor UO_206 (O_206,N_22599,N_24650);
or UO_207 (O_207,N_23007,N_22189);
xor UO_208 (O_208,N_21246,N_24948);
and UO_209 (O_209,N_24225,N_20595);
or UO_210 (O_210,N_23167,N_23161);
xor UO_211 (O_211,N_24289,N_22651);
nand UO_212 (O_212,N_22851,N_20634);
xor UO_213 (O_213,N_21369,N_21033);
nand UO_214 (O_214,N_23884,N_20508);
and UO_215 (O_215,N_23563,N_20554);
or UO_216 (O_216,N_21994,N_23543);
xor UO_217 (O_217,N_22970,N_21872);
nand UO_218 (O_218,N_20185,N_20450);
xnor UO_219 (O_219,N_24473,N_24692);
nor UO_220 (O_220,N_23227,N_21859);
xnor UO_221 (O_221,N_20830,N_23514);
xor UO_222 (O_222,N_24905,N_23553);
nand UO_223 (O_223,N_21599,N_21795);
nand UO_224 (O_224,N_24080,N_21226);
xor UO_225 (O_225,N_22160,N_23740);
or UO_226 (O_226,N_23017,N_21303);
or UO_227 (O_227,N_20889,N_23959);
or UO_228 (O_228,N_23169,N_20757);
xor UO_229 (O_229,N_21029,N_24617);
nand UO_230 (O_230,N_23024,N_20725);
xor UO_231 (O_231,N_20441,N_23441);
or UO_232 (O_232,N_24941,N_22933);
nand UO_233 (O_233,N_22479,N_23634);
nor UO_234 (O_234,N_22658,N_21299);
xor UO_235 (O_235,N_23877,N_23656);
or UO_236 (O_236,N_22999,N_20498);
nor UO_237 (O_237,N_20912,N_22716);
xnor UO_238 (O_238,N_24630,N_20982);
xor UO_239 (O_239,N_23347,N_24302);
or UO_240 (O_240,N_23565,N_21432);
nor UO_241 (O_241,N_22747,N_20302);
xor UO_242 (O_242,N_21510,N_21967);
nor UO_243 (O_243,N_23758,N_21521);
nand UO_244 (O_244,N_21842,N_21276);
or UO_245 (O_245,N_24429,N_21210);
nor UO_246 (O_246,N_24792,N_23924);
and UO_247 (O_247,N_24079,N_23997);
nand UO_248 (O_248,N_22486,N_24264);
and UO_249 (O_249,N_20579,N_20618);
and UO_250 (O_250,N_21824,N_23409);
xnor UO_251 (O_251,N_21085,N_24506);
or UO_252 (O_252,N_24889,N_24886);
nor UO_253 (O_253,N_21910,N_23411);
xnor UO_254 (O_254,N_21215,N_23421);
or UO_255 (O_255,N_21940,N_21290);
or UO_256 (O_256,N_21914,N_22618);
nor UO_257 (O_257,N_23928,N_24099);
or UO_258 (O_258,N_24929,N_23235);
xnor UO_259 (O_259,N_23886,N_21111);
xnor UO_260 (O_260,N_21923,N_24257);
or UO_261 (O_261,N_23913,N_21067);
nand UO_262 (O_262,N_20712,N_21558);
or UO_263 (O_263,N_24376,N_24015);
and UO_264 (O_264,N_20269,N_20258);
nor UO_265 (O_265,N_24782,N_22375);
and UO_266 (O_266,N_22595,N_20133);
nand UO_267 (O_267,N_21797,N_23419);
nor UO_268 (O_268,N_24030,N_24286);
nand UO_269 (O_269,N_21266,N_22540);
xnor UO_270 (O_270,N_21674,N_22020);
or UO_271 (O_271,N_24446,N_24457);
or UO_272 (O_272,N_20815,N_22482);
xor UO_273 (O_273,N_23422,N_20704);
or UO_274 (O_274,N_21622,N_24841);
or UO_275 (O_275,N_23505,N_22224);
and UO_276 (O_276,N_24608,N_22998);
nand UO_277 (O_277,N_20312,N_24972);
nor UO_278 (O_278,N_24424,N_20181);
nand UO_279 (O_279,N_23665,N_21387);
nor UO_280 (O_280,N_24780,N_20467);
nor UO_281 (O_281,N_20756,N_22377);
or UO_282 (O_282,N_22724,N_24508);
or UO_283 (O_283,N_20747,N_23721);
nor UO_284 (O_284,N_21743,N_20386);
and UO_285 (O_285,N_24064,N_22311);
nor UO_286 (O_286,N_22974,N_20214);
nor UO_287 (O_287,N_22628,N_24922);
and UO_288 (O_288,N_23475,N_21243);
or UO_289 (O_289,N_22811,N_23072);
or UO_290 (O_290,N_20316,N_24867);
xor UO_291 (O_291,N_20113,N_23628);
xnor UO_292 (O_292,N_21057,N_24911);
xnor UO_293 (O_293,N_22578,N_23944);
nor UO_294 (O_294,N_24765,N_22588);
xnor UO_295 (O_295,N_21638,N_23545);
or UO_296 (O_296,N_20616,N_20853);
nand UO_297 (O_297,N_20410,N_21784);
xor UO_298 (O_298,N_23868,N_24059);
nor UO_299 (O_299,N_23283,N_23106);
nand UO_300 (O_300,N_22874,N_24487);
or UO_301 (O_301,N_24565,N_20141);
nand UO_302 (O_302,N_21165,N_21672);
nand UO_303 (O_303,N_21884,N_21935);
and UO_304 (O_304,N_24477,N_23427);
xnor UO_305 (O_305,N_22641,N_21927);
or UO_306 (O_306,N_22228,N_20714);
xnor UO_307 (O_307,N_24748,N_20097);
nand UO_308 (O_308,N_24699,N_24169);
nand UO_309 (O_309,N_24816,N_21922);
xor UO_310 (O_310,N_20032,N_20933);
nand UO_311 (O_311,N_21906,N_22687);
nand UO_312 (O_312,N_23844,N_22531);
and UO_313 (O_313,N_23567,N_23662);
nor UO_314 (O_314,N_24652,N_21204);
xnor UO_315 (O_315,N_21479,N_20727);
or UO_316 (O_316,N_23281,N_22111);
and UO_317 (O_317,N_20158,N_21061);
and UO_318 (O_318,N_23433,N_24018);
nor UO_319 (O_319,N_20031,N_20080);
xor UO_320 (O_320,N_21698,N_21883);
xnor UO_321 (O_321,N_20517,N_20276);
nand UO_322 (O_322,N_24090,N_20136);
and UO_323 (O_323,N_20205,N_24956);
or UO_324 (O_324,N_23785,N_21491);
xor UO_325 (O_325,N_23909,N_24382);
xor UO_326 (O_326,N_24970,N_23800);
or UO_327 (O_327,N_21045,N_24654);
nand UO_328 (O_328,N_21168,N_22715);
nand UO_329 (O_329,N_21113,N_23055);
nand UO_330 (O_330,N_22256,N_22398);
or UO_331 (O_331,N_24702,N_24304);
xor UO_332 (O_332,N_22696,N_24644);
or UO_333 (O_333,N_20826,N_22539);
and UO_334 (O_334,N_24683,N_22326);
nor UO_335 (O_335,N_21714,N_23643);
nand UO_336 (O_336,N_23352,N_24356);
nor UO_337 (O_337,N_20689,N_23479);
xnor UO_338 (O_338,N_23091,N_21669);
or UO_339 (O_339,N_22487,N_21468);
nor UO_340 (O_340,N_22201,N_21115);
or UO_341 (O_341,N_22470,N_20344);
or UO_342 (O_342,N_23969,N_23701);
and UO_343 (O_343,N_20235,N_20884);
nor UO_344 (O_344,N_23585,N_20768);
nand UO_345 (O_345,N_23994,N_22782);
nor UO_346 (O_346,N_22163,N_21461);
nand UO_347 (O_347,N_22572,N_23971);
nor UO_348 (O_348,N_24326,N_24423);
nor UO_349 (O_349,N_23314,N_23619);
nand UO_350 (O_350,N_24842,N_21262);
and UO_351 (O_351,N_22986,N_21708);
and UO_352 (O_352,N_21586,N_23245);
nor UO_353 (O_353,N_21181,N_24701);
and UO_354 (O_354,N_22404,N_22632);
and UO_355 (O_355,N_22838,N_24484);
nand UO_356 (O_356,N_24828,N_21684);
and UO_357 (O_357,N_22527,N_23136);
or UO_358 (O_358,N_20695,N_24372);
xor UO_359 (O_359,N_22653,N_20499);
or UO_360 (O_360,N_24004,N_21993);
or UO_361 (O_361,N_21239,N_23883);
or UO_362 (O_362,N_21962,N_22303);
and UO_363 (O_363,N_23137,N_22232);
xor UO_364 (O_364,N_24375,N_21727);
nand UO_365 (O_365,N_21140,N_24456);
nor UO_366 (O_366,N_24733,N_20348);
xor UO_367 (O_367,N_20673,N_22242);
or UO_368 (O_368,N_22499,N_21124);
nand UO_369 (O_369,N_22314,N_24518);
xnor UO_370 (O_370,N_23388,N_23272);
or UO_371 (O_371,N_20829,N_21890);
nor UO_372 (O_372,N_24339,N_21982);
nor UO_373 (O_373,N_21690,N_22215);
nor UO_374 (O_374,N_22223,N_23155);
and UO_375 (O_375,N_22086,N_24129);
xor UO_376 (O_376,N_22315,N_20060);
nand UO_377 (O_377,N_23025,N_23026);
xnor UO_378 (O_378,N_21966,N_24735);
xor UO_379 (O_379,N_22177,N_24812);
nand UO_380 (O_380,N_20468,N_21087);
xnor UO_381 (O_381,N_22609,N_22825);
xor UO_382 (O_382,N_20958,N_21556);
or UO_383 (O_383,N_20449,N_20738);
nor UO_384 (O_384,N_23544,N_23180);
or UO_385 (O_385,N_23461,N_20116);
xnor UO_386 (O_386,N_23804,N_24352);
and UO_387 (O_387,N_20519,N_21222);
or UO_388 (O_388,N_20271,N_21064);
or UO_389 (O_389,N_20718,N_20036);
nor UO_390 (O_390,N_21329,N_22508);
or UO_391 (O_391,N_24177,N_23663);
xnor UO_392 (O_392,N_21309,N_21242);
nand UO_393 (O_393,N_20180,N_20708);
nand UO_394 (O_394,N_24433,N_24656);
nand UO_395 (O_395,N_22534,N_22925);
nand UO_396 (O_396,N_20417,N_21687);
xnor UO_397 (O_397,N_24496,N_20971);
and UO_398 (O_398,N_20140,N_20485);
and UO_399 (O_399,N_21815,N_21676);
nor UO_400 (O_400,N_23633,N_20529);
nand UO_401 (O_401,N_23077,N_22257);
nor UO_402 (O_402,N_21700,N_22755);
or UO_403 (O_403,N_23621,N_21465);
xor UO_404 (O_404,N_21902,N_22659);
and UO_405 (O_405,N_24537,N_24999);
or UO_406 (O_406,N_23152,N_21716);
and UO_407 (O_407,N_20367,N_21288);
xor UO_408 (O_408,N_24208,N_23867);
nand UO_409 (O_409,N_21364,N_20916);
nor UO_410 (O_410,N_23980,N_20119);
nand UO_411 (O_411,N_22930,N_20413);
and UO_412 (O_412,N_21245,N_22808);
nor UO_413 (O_413,N_22173,N_24510);
nor UO_414 (O_414,N_21350,N_21398);
or UO_415 (O_415,N_23853,N_23502);
nand UO_416 (O_416,N_24913,N_23691);
xor UO_417 (O_417,N_21696,N_22932);
and UO_418 (O_418,N_24779,N_20373);
nand UO_419 (O_419,N_20137,N_22875);
nor UO_420 (O_420,N_22510,N_22330);
nand UO_421 (O_421,N_20012,N_24743);
xnor UO_422 (O_422,N_21410,N_24141);
xnor UO_423 (O_423,N_24883,N_23297);
or UO_424 (O_424,N_23765,N_20284);
or UO_425 (O_425,N_22823,N_23204);
and UO_426 (O_426,N_20382,N_23996);
nor UO_427 (O_427,N_21882,N_24887);
and UO_428 (O_428,N_21283,N_23946);
or UO_429 (O_429,N_21527,N_21161);
xor UO_430 (O_430,N_21406,N_22502);
xnor UO_431 (O_431,N_21777,N_23401);
xnor UO_432 (O_432,N_22037,N_21051);
nor UO_433 (O_433,N_23899,N_24950);
nor UO_434 (O_434,N_21677,N_20855);
nor UO_435 (O_435,N_23747,N_21875);
or UO_436 (O_436,N_21666,N_21066);
and UO_437 (O_437,N_22151,N_20108);
nand UO_438 (O_438,N_24104,N_21811);
nand UO_439 (O_439,N_23851,N_24277);
nand UO_440 (O_440,N_22801,N_21808);
nand UO_441 (O_441,N_23798,N_24336);
and UO_442 (O_442,N_23525,N_23606);
and UO_443 (O_443,N_23864,N_24763);
xor UO_444 (O_444,N_21794,N_24354);
and UO_445 (O_445,N_21663,N_21813);
or UO_446 (O_446,N_22981,N_20466);
and UO_447 (O_447,N_24784,N_22985);
and UO_448 (O_448,N_20897,N_21759);
nand UO_449 (O_449,N_21344,N_22633);
nand UO_450 (O_450,N_22230,N_24628);
nor UO_451 (O_451,N_20801,N_21105);
xor UO_452 (O_452,N_22247,N_22497);
or UO_453 (O_453,N_24586,N_23999);
nor UO_454 (O_454,N_21804,N_20793);
nand UO_455 (O_455,N_20486,N_20018);
nand UO_456 (O_456,N_22844,N_20512);
nor UO_457 (O_457,N_20038,N_20358);
nor UO_458 (O_458,N_20201,N_23580);
xnor UO_459 (O_459,N_22213,N_23454);
and UO_460 (O_460,N_20285,N_21343);
xor UO_461 (O_461,N_21056,N_22217);
or UO_462 (O_462,N_22698,N_22800);
xnor UO_463 (O_463,N_21234,N_21623);
and UO_464 (O_464,N_23751,N_22353);
nor UO_465 (O_465,N_22742,N_24503);
nor UO_466 (O_466,N_23476,N_23214);
nor UO_467 (O_467,N_20423,N_20749);
or UO_468 (O_468,N_23767,N_21658);
nand UO_469 (O_469,N_23154,N_22666);
nor UO_470 (O_470,N_23042,N_24342);
nand UO_471 (O_471,N_22165,N_20127);
or UO_472 (O_472,N_23905,N_20935);
or UO_473 (O_473,N_21958,N_20525);
nor UO_474 (O_474,N_20135,N_20240);
and UO_475 (O_475,N_22123,N_24943);
and UO_476 (O_476,N_21835,N_24925);
nand UO_477 (O_477,N_24927,N_23117);
or UO_478 (O_478,N_24135,N_22523);
and UO_479 (O_479,N_20944,N_22402);
and UO_480 (O_480,N_21604,N_22594);
nand UO_481 (O_481,N_23362,N_24105);
xnor UO_482 (O_482,N_24495,N_24437);
nand UO_483 (O_483,N_23712,N_23862);
nor UO_484 (O_484,N_20802,N_23116);
xnor UO_485 (O_485,N_20816,N_24872);
or UO_486 (O_486,N_23102,N_24394);
nor UO_487 (O_487,N_24688,N_22119);
or UO_488 (O_488,N_21722,N_20516);
xnor UO_489 (O_489,N_24625,N_20733);
or UO_490 (O_490,N_24928,N_21968);
and UO_491 (O_491,N_20064,N_21720);
or UO_492 (O_492,N_21457,N_21544);
or UO_493 (O_493,N_23014,N_24421);
nor UO_494 (O_494,N_20028,N_20268);
nand UO_495 (O_495,N_22172,N_21617);
nor UO_496 (O_496,N_24198,N_20987);
xnor UO_497 (O_497,N_20938,N_23005);
nor UO_498 (O_498,N_22779,N_21944);
nand UO_499 (O_499,N_24300,N_22396);
nand UO_500 (O_500,N_21306,N_21102);
and UO_501 (O_501,N_20692,N_20457);
xnor UO_502 (O_502,N_20772,N_21379);
nand UO_503 (O_503,N_24100,N_20521);
or UO_504 (O_504,N_24752,N_23316);
or UO_505 (O_505,N_24581,N_24000);
or UO_506 (O_506,N_24468,N_21588);
nor UO_507 (O_507,N_23035,N_21609);
and UO_508 (O_508,N_21175,N_20115);
xor UO_509 (O_509,N_21528,N_21196);
nand UO_510 (O_510,N_23127,N_24161);
or UO_511 (O_511,N_21869,N_20992);
nor UO_512 (O_512,N_24061,N_22781);
and UO_513 (O_513,N_24512,N_23003);
and UO_514 (O_514,N_21378,N_21856);
or UO_515 (O_515,N_21695,N_21571);
nor UO_516 (O_516,N_21936,N_22552);
nand UO_517 (O_517,N_22045,N_21017);
nor UO_518 (O_518,N_23387,N_20887);
or UO_519 (O_519,N_24520,N_23624);
xnor UO_520 (O_520,N_20917,N_21657);
and UO_521 (O_521,N_20247,N_22416);
and UO_522 (O_522,N_24521,N_24708);
nand UO_523 (O_523,N_21421,N_20156);
nand UO_524 (O_524,N_21450,N_23194);
nand UO_525 (O_525,N_22916,N_24449);
nor UO_526 (O_526,N_24971,N_23082);
xnor UO_527 (O_527,N_21662,N_22968);
nand UO_528 (O_528,N_21500,N_21610);
and UO_529 (O_529,N_24830,N_22856);
or UO_530 (O_530,N_20561,N_21782);
nand UO_531 (O_531,N_23791,N_24539);
or UO_532 (O_532,N_20722,N_21208);
nor UO_533 (O_533,N_20099,N_24074);
and UO_534 (O_534,N_23285,N_23271);
and UO_535 (O_535,N_21997,N_20758);
and UO_536 (O_536,N_21624,N_24084);
nand UO_537 (O_537,N_24619,N_23940);
and UO_538 (O_538,N_23934,N_24103);
nand UO_539 (O_539,N_20957,N_20049);
nand UO_540 (O_540,N_23400,N_24332);
and UO_541 (O_541,N_24964,N_21478);
and UO_542 (O_542,N_22614,N_22717);
nor UO_543 (O_543,N_20228,N_24501);
nand UO_544 (O_544,N_22048,N_22042);
nand UO_545 (O_545,N_22701,N_23175);
and UO_546 (O_546,N_22988,N_24805);
xor UO_547 (O_547,N_20715,N_22557);
or UO_548 (O_548,N_23783,N_21786);
nand UO_549 (O_549,N_21048,N_22753);
or UO_550 (O_550,N_24091,N_22979);
nand UO_551 (O_551,N_23600,N_22674);
and UO_552 (O_552,N_22959,N_22512);
or UO_553 (O_553,N_23099,N_23894);
nor UO_554 (O_554,N_24254,N_22777);
nor UO_555 (O_555,N_24139,N_22385);
or UO_556 (O_556,N_22965,N_20911);
nor UO_557 (O_557,N_20845,N_22076);
nor UO_558 (O_558,N_23937,N_20598);
nand UO_559 (O_559,N_21717,N_20282);
xor UO_560 (O_560,N_21809,N_24963);
nand UO_561 (O_561,N_22553,N_21131);
or UO_562 (O_562,N_23488,N_21707);
xnor UO_563 (O_563,N_23208,N_21474);
nand UO_564 (O_564,N_20061,N_24204);
xnor UO_565 (O_565,N_20905,N_20668);
and UO_566 (O_566,N_22832,N_23207);
and UO_567 (O_567,N_20005,N_22921);
nand UO_568 (O_568,N_24725,N_24233);
xnor UO_569 (O_569,N_21171,N_24131);
or UO_570 (O_570,N_23687,N_23429);
nand UO_571 (O_571,N_22073,N_23318);
nand UO_572 (O_572,N_22810,N_20593);
or UO_573 (O_573,N_24535,N_23547);
xor UO_574 (O_574,N_23970,N_20500);
or UO_575 (O_575,N_24534,N_23818);
nor UO_576 (O_576,N_22229,N_24620);
xor UO_577 (O_577,N_23494,N_20709);
xor UO_578 (O_578,N_21186,N_21596);
or UO_579 (O_579,N_22312,N_23090);
or UO_580 (O_580,N_20277,N_23515);
and UO_581 (O_581,N_21355,N_22967);
and UO_582 (O_582,N_24632,N_24479);
nor UO_583 (O_583,N_20469,N_23673);
xnor UO_584 (O_584,N_22940,N_20305);
or UO_585 (O_585,N_22740,N_22563);
xnor UO_586 (O_586,N_24417,N_20289);
nor UO_587 (O_587,N_23892,N_20563);
xnor UO_588 (O_588,N_22547,N_20539);
nand UO_589 (O_589,N_22601,N_20763);
nor UO_590 (O_590,N_21939,N_20541);
or UO_591 (O_591,N_21157,N_22361);
and UO_592 (O_592,N_23604,N_20913);
or UO_593 (O_593,N_21858,N_23330);
and UO_594 (O_594,N_20318,N_23020);
nor UO_595 (O_595,N_21332,N_21408);
xnor UO_596 (O_596,N_24554,N_22132);
xnor UO_597 (O_597,N_22743,N_21789);
and UO_598 (O_598,N_23728,N_24968);
and UO_599 (O_599,N_21986,N_24324);
or UO_600 (O_600,N_21888,N_24012);
and UO_601 (O_601,N_24937,N_20775);
or UO_602 (O_602,N_21172,N_22710);
nor UO_603 (O_603,N_24034,N_24474);
and UO_604 (O_604,N_24299,N_23156);
nand UO_605 (O_605,N_23493,N_22663);
nor UO_606 (O_606,N_23251,N_24915);
and UO_607 (O_607,N_22174,N_24720);
or UO_608 (O_608,N_21489,N_23654);
and UO_609 (O_609,N_24594,N_23120);
nand UO_610 (O_610,N_21688,N_20762);
nor UO_611 (O_611,N_22016,N_20723);
and UO_612 (O_612,N_20057,N_21713);
or UO_613 (O_613,N_22018,N_23168);
and UO_614 (O_614,N_24036,N_21721);
or UO_615 (O_615,N_20617,N_20027);
nor UO_616 (O_616,N_24447,N_24301);
or UO_617 (O_617,N_20209,N_23891);
xnor UO_618 (O_618,N_22829,N_24207);
nand UO_619 (O_619,N_24073,N_22634);
xnor UO_620 (O_620,N_24651,N_23507);
xor UO_621 (O_621,N_24646,N_20296);
and UO_622 (O_622,N_20076,N_24712);
nor UO_623 (O_623,N_23040,N_24672);
nor UO_624 (O_624,N_23424,N_23732);
or UO_625 (O_625,N_20474,N_20980);
or UO_626 (O_626,N_23914,N_20443);
xor UO_627 (O_627,N_21134,N_23049);
nand UO_628 (O_628,N_20602,N_22676);
xor UO_629 (O_629,N_21961,N_20927);
or UO_630 (O_630,N_23470,N_24327);
and UO_631 (O_631,N_23298,N_21368);
nor UO_632 (O_632,N_23848,N_21852);
nand UO_633 (O_633,N_20691,N_23960);
xnor UO_634 (O_634,N_21354,N_23554);
nand UO_635 (O_635,N_20546,N_22606);
nor UO_636 (O_636,N_22947,N_21664);
xor UO_637 (O_637,N_23267,N_20159);
xnor UO_638 (O_638,N_22254,N_22277);
nor UO_639 (O_639,N_22884,N_20054);
xor UO_640 (O_640,N_21998,N_23815);
and UO_641 (O_641,N_22962,N_20458);
nand UO_642 (O_642,N_21107,N_20644);
or UO_643 (O_643,N_24961,N_23255);
nor UO_644 (O_644,N_23398,N_22616);
or UO_645 (O_645,N_20088,N_22176);
or UO_646 (O_646,N_24285,N_22529);
nand UO_647 (O_647,N_22944,N_21063);
nor UO_648 (O_648,N_23918,N_23484);
nor UO_649 (O_649,N_21564,N_23089);
nand UO_650 (O_650,N_21294,N_22038);
or UO_651 (O_651,N_20067,N_20199);
nor UO_652 (O_652,N_21311,N_23234);
and UO_653 (O_653,N_21145,N_24575);
nor UO_654 (O_654,N_24025,N_22170);
nor UO_655 (O_655,N_21143,N_20259);
nand UO_656 (O_656,N_22183,N_21860);
nor UO_657 (O_657,N_24452,N_20182);
nand UO_658 (O_658,N_21757,N_22146);
xnor UO_659 (O_659,N_21334,N_22922);
nand UO_660 (O_660,N_22685,N_21331);
and UO_661 (O_661,N_22835,N_24404);
or UO_662 (O_662,N_23407,N_20188);
and UO_663 (O_663,N_20729,N_20846);
and UO_664 (O_664,N_22927,N_22084);
or UO_665 (O_665,N_21689,N_22918);
nor UO_666 (O_666,N_21499,N_21308);
nand UO_667 (O_667,N_24111,N_24860);
and UO_668 (O_668,N_22975,N_23810);
xor UO_669 (O_669,N_22127,N_24715);
nand UO_670 (O_670,N_21542,N_20189);
xnor UO_671 (O_671,N_23113,N_23426);
or UO_672 (O_672,N_20837,N_22089);
and UO_673 (O_673,N_22708,N_24729);
nand UO_674 (O_674,N_20900,N_22270);
xnor UO_675 (O_675,N_24696,N_21818);
and UO_676 (O_676,N_20047,N_23164);
xnor UO_677 (O_677,N_23852,N_21091);
nand UO_678 (O_678,N_22423,N_23392);
nor UO_679 (O_679,N_20362,N_22491);
nand UO_680 (O_680,N_22010,N_21090);
nor UO_681 (O_681,N_22516,N_20233);
nor UO_682 (O_682,N_21762,N_24465);
and UO_683 (O_683,N_24838,N_22713);
or UO_684 (O_684,N_21300,N_21990);
nor UO_685 (O_685,N_20352,N_22963);
or UO_686 (O_686,N_24017,N_20033);
or UO_687 (O_687,N_23257,N_22524);
or UO_688 (O_688,N_20424,N_20937);
nand UO_689 (O_689,N_21728,N_23875);
and UO_690 (O_690,N_23250,N_21733);
nand UO_691 (O_691,N_21778,N_21506);
nor UO_692 (O_692,N_20878,N_23828);
and UO_693 (O_693,N_23698,N_24031);
nor UO_694 (O_694,N_23066,N_22030);
and UO_695 (O_695,N_22994,N_20582);
xor UO_696 (O_696,N_22046,N_24808);
nor UO_697 (O_697,N_20651,N_23492);
or UO_698 (O_698,N_22434,N_22343);
nand UO_699 (O_699,N_23676,N_22290);
xnor UO_700 (O_700,N_22677,N_21874);
and UO_701 (O_701,N_24798,N_23953);
nand UO_702 (O_702,N_24284,N_21803);
and UO_703 (O_703,N_23126,N_22993);
or UO_704 (O_704,N_20633,N_23598);
nand UO_705 (O_705,N_24493,N_24978);
or UO_706 (O_706,N_21429,N_22463);
or UO_707 (O_707,N_23976,N_20818);
xor UO_708 (O_708,N_24827,N_24543);
and UO_709 (O_709,N_20196,N_20210);
nand UO_710 (O_710,N_21278,N_21152);
nand UO_711 (O_711,N_20206,N_23978);
nor UO_712 (O_712,N_20697,N_20337);
nor UO_713 (O_713,N_21426,N_21791);
nand UO_714 (O_714,N_21483,N_22886);
and UO_715 (O_715,N_20491,N_20055);
and UO_716 (O_716,N_23988,N_21889);
nand UO_717 (O_717,N_20347,N_20451);
or UO_718 (O_718,N_23181,N_20171);
or UO_719 (O_719,N_23478,N_22181);
xor UO_720 (O_720,N_24127,N_24945);
nand UO_721 (O_721,N_21055,N_23324);
nor UO_722 (O_722,N_21865,N_22219);
or UO_723 (O_723,N_23769,N_23956);
or UO_724 (O_724,N_20224,N_24669);
nand UO_725 (O_725,N_23569,N_23575);
nand UO_726 (O_726,N_22441,N_20902);
or UO_727 (O_727,N_24781,N_22301);
and UO_728 (O_728,N_24399,N_23481);
nand UO_729 (O_729,N_20785,N_22624);
nand UO_730 (O_730,N_22905,N_20492);
nand UO_731 (O_731,N_24890,N_21730);
and UO_732 (O_732,N_20040,N_23443);
nand UO_733 (O_733,N_20408,N_20391);
nor UO_734 (O_734,N_20823,N_24388);
or UO_735 (O_735,N_22764,N_24871);
nand UO_736 (O_736,N_24755,N_20730);
nor UO_737 (O_737,N_21319,N_24580);
nor UO_738 (O_738,N_23648,N_23957);
or UO_739 (O_739,N_24789,N_23319);
or UO_740 (O_740,N_23221,N_22697);
and UO_741 (O_741,N_24239,N_20873);
nand UO_742 (O_742,N_22352,N_21705);
xnor UO_743 (O_743,N_21981,N_23358);
nand UO_744 (O_744,N_20342,N_23170);
xor UO_745 (O_745,N_23830,N_21189);
and UO_746 (O_746,N_23140,N_20392);
and UO_747 (O_747,N_20454,N_24635);
and UO_748 (O_748,N_21792,N_20773);
or UO_749 (O_749,N_22104,N_23733);
nor UO_750 (O_750,N_23218,N_23797);
nor UO_751 (O_751,N_20083,N_24316);
xnor UO_752 (O_752,N_20871,N_24016);
or UO_753 (O_753,N_21282,N_23813);
nand UO_754 (O_754,N_24577,N_24095);
xnor UO_755 (O_755,N_20649,N_23559);
nor UO_756 (O_756,N_20592,N_23512);
xor UO_757 (O_757,N_20612,N_22969);
and UO_758 (O_758,N_23773,N_21418);
or UO_759 (O_759,N_23109,N_21076);
and UO_760 (O_760,N_21009,N_20688);
and UO_761 (O_761,N_21392,N_22367);
or UO_762 (O_762,N_20888,N_22096);
or UO_763 (O_763,N_20094,N_22047);
xnor UO_764 (O_764,N_21877,N_21620);
nand UO_765 (O_765,N_23002,N_24089);
nand UO_766 (O_766,N_22272,N_20780);
nand UO_767 (O_767,N_22605,N_22415);
and UO_768 (O_768,N_24215,N_20711);
xor UO_769 (O_769,N_20003,N_24985);
nor UO_770 (O_770,N_20422,N_24303);
nor UO_771 (O_771,N_24063,N_24211);
nor UO_772 (O_772,N_23840,N_23531);
nor UO_773 (O_773,N_24389,N_20223);
and UO_774 (O_774,N_20783,N_23315);
and UO_775 (O_775,N_21082,N_22977);
xor UO_776 (O_776,N_22431,N_20166);
xor UO_777 (O_777,N_23103,N_24797);
nand UO_778 (O_778,N_21807,N_20588);
or UO_779 (O_779,N_21566,N_21146);
or UO_780 (O_780,N_21488,N_20145);
nand UO_781 (O_781,N_22853,N_20429);
or UO_782 (O_782,N_20161,N_22954);
and UO_783 (O_783,N_22112,N_21182);
nand UO_784 (O_784,N_21273,N_24923);
nand UO_785 (O_785,N_23880,N_20042);
nor UO_786 (O_786,N_22671,N_20681);
xnor UO_787 (O_787,N_24483,N_24834);
and UO_788 (O_788,N_20522,N_20148);
and UO_789 (O_789,N_24368,N_21099);
xor UO_790 (O_790,N_22258,N_24666);
nor UO_791 (O_791,N_23135,N_21648);
nand UO_792 (O_792,N_22306,N_22297);
and UO_793 (O_793,N_21220,N_20741);
xor UO_794 (O_794,N_23968,N_24693);
xor UO_795 (O_795,N_21219,N_23325);
xor UO_796 (O_796,N_24023,N_22603);
xor UO_797 (O_797,N_23594,N_21233);
and UO_798 (O_798,N_20198,N_24631);
and UO_799 (O_799,N_24924,N_20363);
nand UO_800 (O_800,N_24164,N_20056);
and UO_801 (O_801,N_21855,N_22850);
xnor UO_802 (O_802,N_20750,N_23744);
nor UO_803 (O_803,N_24058,N_20960);
and UO_804 (O_804,N_20832,N_20817);
xor UO_805 (O_805,N_24946,N_20596);
and UO_806 (O_806,N_23213,N_22668);
nand UO_807 (O_807,N_22804,N_23345);
nand UO_808 (O_808,N_21508,N_23205);
nor UO_809 (O_809,N_20868,N_24906);
nand UO_810 (O_810,N_20396,N_22198);
or UO_811 (O_811,N_21073,N_22942);
xor UO_812 (O_812,N_23586,N_20872);
nand UO_813 (O_813,N_22035,N_21149);
nor UO_814 (O_814,N_21569,N_22308);
xor UO_815 (O_815,N_21270,N_21008);
xor UO_816 (O_816,N_21568,N_22865);
nor UO_817 (O_817,N_21825,N_21428);
and UO_818 (O_818,N_23334,N_23823);
and UO_819 (O_819,N_23664,N_22911);
nand UO_820 (O_820,N_21636,N_21531);
nand UO_821 (O_821,N_22408,N_21327);
and UO_822 (O_822,N_20366,N_24297);
xor UO_823 (O_823,N_22291,N_20026);
nor UO_824 (O_824,N_23471,N_23620);
xor UO_825 (O_825,N_22759,N_22087);
and UO_826 (O_826,N_22868,N_20643);
nor UO_827 (O_827,N_20854,N_20626);
and UO_828 (O_828,N_23053,N_23353);
nand UO_829 (O_829,N_21627,N_22360);
xor UO_830 (O_830,N_24227,N_22950);
and UO_831 (O_831,N_22758,N_24334);
and UO_832 (O_832,N_23394,N_23987);
xnor UO_833 (O_833,N_24355,N_24572);
xnor UO_834 (O_834,N_22700,N_22514);
nor UO_835 (O_835,N_20796,N_23693);
or UO_836 (O_836,N_24603,N_24909);
xor UO_837 (O_837,N_22924,N_21886);
nand UO_838 (O_838,N_21774,N_23770);
nor UO_839 (O_839,N_23703,N_23489);
xnor UO_840 (O_840,N_21191,N_22462);
xor UO_841 (O_841,N_20483,N_22876);
or UO_842 (O_842,N_22108,N_21200);
nand UO_843 (O_843,N_21495,N_24329);
xnor UO_844 (O_844,N_24875,N_21375);
or UO_845 (O_845,N_24564,N_24851);
nand UO_846 (O_846,N_22004,N_23645);
xor UO_847 (O_847,N_20153,N_20791);
xor UO_848 (O_848,N_21423,N_24505);
nor UO_849 (O_849,N_21249,N_24547);
or UO_850 (O_850,N_22321,N_23903);
xnor UO_851 (O_851,N_20351,N_21509);
or UO_852 (O_852,N_24043,N_22476);
xor UO_853 (O_853,N_24197,N_23070);
or UO_854 (O_854,N_21640,N_21954);
or UO_855 (O_855,N_24601,N_22075);
xnor UO_856 (O_856,N_23329,N_21699);
and UO_857 (O_857,N_20254,N_24854);
or UO_858 (O_858,N_22560,N_24419);
nand UO_859 (O_859,N_24463,N_22520);
and UO_860 (O_860,N_24454,N_21054);
nor UO_861 (O_861,N_21490,N_20859);
nor UO_862 (O_862,N_21015,N_20440);
xnor UO_863 (O_863,N_20107,N_23351);
nor UO_864 (O_864,N_23051,N_24214);
nor UO_865 (O_865,N_20331,N_23437);
xnor UO_866 (O_866,N_21755,N_24333);
nor UO_867 (O_867,N_20895,N_20613);
nor UO_868 (O_868,N_22464,N_20842);
xnor UO_869 (O_869,N_22318,N_20283);
nand UO_870 (O_870,N_23660,N_22208);
or UO_871 (O_871,N_20581,N_22766);
and UO_872 (O_872,N_21211,N_24144);
nor UO_873 (O_873,N_21549,N_22394);
nand UO_874 (O_874,N_24445,N_21530);
or UO_875 (O_875,N_23599,N_23439);
or UO_876 (O_876,N_23869,N_21848);
xor UO_877 (O_877,N_24240,N_22664);
or UO_878 (O_878,N_21496,N_23355);
or UO_879 (O_879,N_23895,N_21199);
xnor UO_880 (O_880,N_23254,N_20666);
and UO_881 (O_881,N_22725,N_22427);
and UO_882 (O_882,N_23963,N_21652);
nor UO_883 (O_883,N_23209,N_21760);
nand UO_884 (O_884,N_22355,N_24205);
and UO_885 (O_885,N_22354,N_22333);
nand UO_886 (O_886,N_22902,N_23617);
and UO_887 (O_887,N_21843,N_23046);
and UO_888 (O_888,N_23199,N_24990);
nand UO_889 (O_889,N_21507,N_21866);
nor UO_890 (O_890,N_21641,N_23964);
and UO_891 (O_891,N_24163,N_20530);
nor UO_892 (O_892,N_24062,N_23898);
and UO_893 (O_893,N_24843,N_23177);
nand UO_894 (O_894,N_24330,N_23819);
xor UO_895 (O_895,N_23657,N_20420);
and UO_896 (O_896,N_23816,N_21252);
or UO_897 (O_897,N_24408,N_20232);
or UO_898 (O_898,N_22243,N_21002);
nand UO_899 (O_899,N_23950,N_24294);
nor UO_900 (O_900,N_24152,N_22493);
nand UO_901 (O_901,N_22718,N_20962);
or UO_902 (O_902,N_22364,N_21313);
nand UO_903 (O_903,N_23907,N_22197);
nor UO_904 (O_904,N_23707,N_24055);
xnor UO_905 (O_905,N_24556,N_21829);
and UO_906 (O_906,N_22709,N_22466);
or UO_907 (O_907,N_21178,N_22064);
nand UO_908 (O_908,N_24536,N_23768);
or UO_909 (O_909,N_20341,N_21963);
nand UO_910 (O_910,N_20631,N_23301);
xor UO_911 (O_911,N_23242,N_21526);
or UO_912 (O_912,N_24235,N_23241);
and UO_913 (O_913,N_23151,N_22941);
nand UO_914 (O_914,N_20765,N_20152);
and UO_915 (O_915,N_24926,N_22386);
or UO_916 (O_916,N_24606,N_21692);
and UO_917 (O_917,N_21585,N_24877);
xnor UO_918 (O_918,N_21000,N_23837);
and UO_919 (O_919,N_20792,N_24710);
xor UO_920 (O_920,N_22251,N_22342);
nor UO_921 (O_921,N_21557,N_20808);
and UO_922 (O_922,N_21039,N_21634);
nor UO_923 (O_923,N_24026,N_20555);
nor UO_924 (O_924,N_20686,N_20743);
nand UO_925 (O_925,N_23795,N_23724);
or UO_926 (O_926,N_22244,N_21943);
nand UO_927 (O_927,N_20143,N_24102);
xnor UO_928 (O_928,N_23933,N_24562);
and UO_929 (O_929,N_24588,N_21224);
nor UO_930 (O_930,N_21322,N_21214);
xnor UO_931 (O_931,N_22997,N_22972);
or UO_932 (O_932,N_23033,N_23317);
or UO_933 (O_933,N_23929,N_22069);
nor UO_934 (O_934,N_23165,N_24364);
nor UO_935 (O_935,N_22805,N_21241);
nor UO_936 (O_936,N_23735,N_20095);
and UO_937 (O_937,N_24994,N_23435);
nor UO_938 (O_938,N_23472,N_20407);
and UO_939 (O_939,N_21185,N_23566);
or UO_940 (O_940,N_24272,N_20266);
nor UO_941 (O_941,N_22307,N_23821);
xnor UO_942 (O_942,N_23348,N_24987);
xnor UO_943 (O_943,N_23535,N_20081);
xor UO_944 (O_944,N_22847,N_24200);
nor UO_945 (O_945,N_24846,N_24425);
or UO_946 (O_946,N_23548,N_23396);
nand UO_947 (O_947,N_21130,N_23028);
nand UO_948 (O_948,N_24659,N_24262);
nor UO_949 (O_949,N_21796,N_21864);
and UO_950 (O_950,N_20942,N_24947);
and UO_951 (O_951,N_20896,N_24271);
nor UO_952 (O_952,N_22000,N_22237);
or UO_953 (O_953,N_20954,N_21747);
xnor UO_954 (O_954,N_21711,N_22731);
nand UO_955 (O_955,N_24310,N_21042);
or UO_956 (O_956,N_24839,N_24967);
and UO_957 (O_957,N_22788,N_24068);
xnor UO_958 (O_958,N_22182,N_24629);
or UO_959 (O_959,N_23776,N_21424);
nor UO_960 (O_960,N_21376,N_21775);
or UO_961 (O_961,N_21862,N_20985);
and UO_962 (O_962,N_22212,N_23504);
and UO_963 (O_963,N_24874,N_23754);
or UO_964 (O_964,N_24653,N_21248);
nor UO_965 (O_965,N_21030,N_23371);
xor UO_966 (O_966,N_21289,N_23122);
nor UO_967 (O_967,N_22013,N_24904);
xor UO_968 (O_968,N_24661,N_23185);
and UO_969 (O_969,N_20487,N_22734);
xor UO_970 (O_970,N_22507,N_24989);
nor UO_971 (O_971,N_24448,N_22150);
nor UO_972 (O_972,N_22780,N_23562);
and UO_973 (O_973,N_20418,N_24979);
or UO_974 (O_974,N_20178,N_24823);
and UO_975 (O_975,N_21937,N_22796);
xor UO_976 (O_976,N_24933,N_22625);
or UO_977 (O_977,N_20576,N_24959);
or UO_978 (O_978,N_21916,N_21230);
xor UO_979 (O_979,N_20216,N_21771);
and UO_980 (O_980,N_24745,N_21352);
nor UO_981 (O_981,N_20447,N_23926);
and UO_982 (O_982,N_24689,N_22877);
xnor UO_983 (O_983,N_23382,N_21485);
and UO_984 (O_984,N_22754,N_21166);
and UO_985 (O_985,N_23992,N_20657);
or UO_986 (O_986,N_24274,N_24002);
and UO_987 (O_987,N_24178,N_21702);
nor UO_988 (O_988,N_22019,N_21522);
xor UO_989 (O_989,N_22335,N_22532);
and UO_990 (O_990,N_23832,N_22757);
and UO_991 (O_991,N_24787,N_24427);
nor UO_992 (O_992,N_24907,N_24252);
nor UO_993 (O_993,N_22773,N_20332);
nor UO_994 (O_994,N_20713,N_23709);
nand UO_995 (O_995,N_22723,N_21482);
xnor UO_996 (O_996,N_23684,N_22570);
nor UO_997 (O_997,N_20208,N_22961);
and UO_998 (O_998,N_21909,N_21381);
nand UO_999 (O_999,N_24440,N_21851);
xnor UO_1000 (O_1000,N_21118,N_23995);
nand UO_1001 (O_1001,N_23406,N_22346);
or UO_1002 (O_1002,N_24269,N_24517);
nor UO_1003 (O_1003,N_21693,N_23874);
nand UO_1004 (O_1004,N_21255,N_24362);
nor UO_1005 (O_1005,N_23609,N_20125);
nand UO_1006 (O_1006,N_21686,N_23666);
nand UO_1007 (O_1007,N_23872,N_24032);
nand UO_1008 (O_1008,N_20303,N_21027);
and UO_1009 (O_1009,N_22561,N_21719);
and UO_1010 (O_1010,N_23973,N_23184);
or UO_1011 (O_1011,N_23811,N_24804);
and UO_1012 (O_1012,N_22909,N_23876);
xnor UO_1013 (O_1013,N_22906,N_20298);
nand UO_1014 (O_1014,N_24640,N_22517);
or UO_1015 (O_1015,N_20672,N_23374);
xor UO_1016 (O_1016,N_20505,N_20946);
or UO_1017 (O_1017,N_22577,N_22161);
or UO_1018 (O_1018,N_22881,N_22783);
nor UO_1019 (O_1019,N_23736,N_21907);
nand UO_1020 (O_1020,N_24345,N_20922);
xnor UO_1021 (O_1021,N_24232,N_23850);
xnor UO_1022 (O_1022,N_23287,N_20952);
xor UO_1023 (O_1023,N_24958,N_23112);
and UO_1024 (O_1024,N_21216,N_20165);
nor UO_1025 (O_1025,N_21437,N_21584);
xor UO_1026 (O_1026,N_24101,N_22263);
and UO_1027 (O_1027,N_23863,N_22265);
nand UO_1028 (O_1028,N_24476,N_21979);
nand UO_1029 (O_1029,N_21271,N_21005);
nor UO_1030 (O_1030,N_22582,N_21974);
or UO_1031 (O_1031,N_21213,N_22054);
or UO_1032 (O_1032,N_24935,N_23201);
or UO_1033 (O_1033,N_24774,N_23774);
and UO_1034 (O_1034,N_24266,N_22320);
nand UO_1035 (O_1035,N_22492,N_20092);
xor UO_1036 (O_1036,N_21660,N_20735);
or UO_1037 (O_1037,N_21274,N_23290);
and UO_1038 (O_1038,N_20020,N_24248);
or UO_1039 (O_1039,N_21492,N_23865);
nand UO_1040 (O_1040,N_23430,N_22193);
nand UO_1041 (O_1041,N_21148,N_20676);
nor UO_1042 (O_1042,N_24613,N_22719);
or UO_1043 (O_1043,N_20812,N_22299);
and UO_1044 (O_1044,N_20155,N_22980);
nand UO_1045 (O_1045,N_20222,N_20737);
nor UO_1046 (O_1046,N_22813,N_23499);
or UO_1047 (O_1047,N_22645,N_21301);
and UO_1048 (O_1048,N_20543,N_20518);
nor UO_1049 (O_1049,N_24021,N_24174);
and UO_1050 (O_1050,N_21605,N_24835);
nor UO_1051 (O_1051,N_22675,N_23219);
xnor UO_1052 (O_1052,N_21919,N_21139);
or UO_1053 (O_1053,N_20242,N_22699);
nor UO_1054 (O_1054,N_20460,N_24107);
and UO_1055 (O_1055,N_24346,N_22382);
and UO_1056 (O_1056,N_23729,N_24976);
nor UO_1057 (O_1057,N_21456,N_20129);
or UO_1058 (O_1058,N_23841,N_24738);
or UO_1059 (O_1059,N_24146,N_24488);
and UO_1060 (O_1060,N_20645,N_22095);
and UO_1061 (O_1061,N_20532,N_20675);
and UO_1062 (O_1062,N_21359,N_22106);
or UO_1063 (O_1063,N_24218,N_20146);
nor UO_1064 (O_1064,N_20509,N_23561);
xnor UO_1065 (O_1065,N_24298,N_21912);
xor UO_1066 (O_1066,N_24134,N_24395);
and UO_1067 (O_1067,N_24621,N_24442);
nand UO_1068 (O_1068,N_23132,N_24502);
xnor UO_1069 (O_1069,N_22515,N_22362);
nand UO_1070 (O_1070,N_24186,N_21512);
xnor UO_1071 (O_1071,N_22124,N_21536);
and UO_1072 (O_1072,N_20253,N_22113);
and UO_1073 (O_1073,N_22003,N_20893);
or UO_1074 (O_1074,N_22319,N_23857);
nand UO_1075 (O_1075,N_22834,N_23247);
nor UO_1076 (O_1076,N_23589,N_24293);
xnor UO_1077 (O_1077,N_24311,N_24048);
nand UO_1078 (O_1078,N_22332,N_22971);
and UO_1079 (O_1079,N_21293,N_23942);
and UO_1080 (O_1080,N_24438,N_20046);
or UO_1081 (O_1081,N_21287,N_20239);
or UO_1082 (O_1082,N_24582,N_23423);
xnor UO_1083 (O_1083,N_20346,N_24156);
nor UO_1084 (O_1084,N_23009,N_21093);
xor UO_1085 (O_1085,N_22840,N_23870);
nand UO_1086 (O_1086,N_20377,N_23530);
nor UO_1087 (O_1087,N_24691,N_22295);
xor UO_1088 (O_1088,N_23350,N_21635);
and UO_1089 (O_1089,N_22456,N_21656);
nor UO_1090 (O_1090,N_22660,N_21973);
nor UO_1091 (O_1091,N_20270,N_20720);
or UO_1092 (O_1092,N_24751,N_22953);
and UO_1093 (O_1093,N_23742,N_20751);
nor UO_1094 (O_1094,N_20628,N_20840);
and UO_1095 (O_1095,N_20545,N_23456);
and UO_1096 (O_1096,N_22454,N_20862);
and UO_1097 (O_1097,N_23670,N_21911);
and UO_1098 (O_1098,N_22914,N_20497);
and UO_1099 (O_1099,N_22960,N_23506);
and UO_1100 (O_1100,N_23967,N_20197);
nor UO_1101 (O_1101,N_24544,N_20836);
xor UO_1102 (O_1102,N_22238,N_23993);
xor UO_1103 (O_1103,N_21156,N_23309);
nor UO_1104 (O_1104,N_21938,N_24460);
nand UO_1105 (O_1105,N_21853,N_21453);
xor UO_1106 (O_1106,N_20227,N_21734);
nor UO_1107 (O_1107,N_20558,N_21600);
or UO_1108 (O_1108,N_22935,N_23760);
and UO_1109 (O_1109,N_23668,N_22392);
and UO_1110 (O_1110,N_21983,N_23121);
or UO_1111 (O_1111,N_21917,N_21383);
and UO_1112 (O_1112,N_23303,N_20273);
xor UO_1113 (O_1113,N_23990,N_24273);
or UO_1114 (O_1114,N_21749,N_20104);
xor UO_1115 (O_1115,N_24773,N_22720);
or UO_1116 (O_1116,N_24515,N_20814);
or UO_1117 (O_1117,N_22519,N_23331);
and UO_1118 (O_1118,N_24003,N_24681);
and UO_1119 (O_1119,N_24932,N_22339);
or UO_1120 (O_1120,N_21575,N_24850);
and UO_1121 (O_1121,N_22647,N_21104);
and UO_1122 (O_1122,N_21988,N_20805);
and UO_1123 (O_1123,N_20607,N_24992);
nand UO_1124 (O_1124,N_20599,N_20448);
and UO_1125 (O_1125,N_22414,N_24428);
nand UO_1126 (O_1126,N_20760,N_22682);
xnor UO_1127 (O_1127,N_22128,N_24243);
xor UO_1128 (O_1128,N_23268,N_22439);
nor UO_1129 (O_1129,N_21631,N_22841);
nor UO_1130 (O_1130,N_23827,N_21333);
nor UO_1131 (O_1131,N_24391,N_24154);
nand UO_1132 (O_1132,N_24845,N_24788);
nand UO_1133 (O_1133,N_20257,N_22447);
xor UO_1134 (O_1134,N_21583,N_23847);
or UO_1135 (O_1135,N_20510,N_22430);
xor UO_1136 (O_1136,N_21957,N_23659);
or UO_1137 (O_1137,N_24991,N_23786);
nand UO_1138 (O_1138,N_20943,N_21577);
xnor UO_1139 (O_1139,N_22631,N_21250);
xor UO_1140 (O_1140,N_23500,N_20920);
or UO_1141 (O_1141,N_20109,N_24092);
nor UO_1142 (O_1142,N_21430,N_21633);
nand UO_1143 (O_1143,N_24697,N_23460);
xnor UO_1144 (O_1144,N_21314,N_23610);
or UO_1145 (O_1145,N_21934,N_22262);
and UO_1146 (O_1146,N_24358,N_20463);
and UO_1147 (O_1147,N_23100,N_24509);
and UO_1148 (O_1148,N_21467,N_22518);
and UO_1149 (O_1149,N_22289,N_23954);
nor UO_1150 (O_1150,N_23685,N_22023);
or UO_1151 (O_1151,N_22002,N_24918);
or UO_1152 (O_1152,N_20068,N_23834);
or UO_1153 (O_1153,N_23527,N_24567);
nand UO_1154 (O_1154,N_22819,N_20690);
xor UO_1155 (O_1155,N_23699,N_23270);
nand UO_1156 (O_1156,N_23887,N_22141);
and UO_1157 (O_1157,N_20687,N_24576);
nor UO_1158 (O_1158,N_23532,N_23904);
xor UO_1159 (O_1159,N_21225,N_20578);
xnor UO_1160 (O_1160,N_20203,N_23674);
and UO_1161 (O_1161,N_20655,N_23171);
nor UO_1162 (O_1162,N_20559,N_24097);
nor UO_1163 (O_1163,N_24848,N_23372);
nand UO_1164 (O_1164,N_21142,N_20833);
nand UO_1165 (O_1165,N_20748,N_23340);
or UO_1166 (O_1166,N_23436,N_24148);
nor UO_1167 (O_1167,N_21155,N_22012);
and UO_1168 (O_1168,N_24162,N_22892);
and UO_1169 (O_1169,N_22300,N_23838);
xor UO_1170 (O_1170,N_21320,N_20470);
nor UO_1171 (O_1171,N_20699,N_24749);
and UO_1172 (O_1172,N_21415,N_20537);
or UO_1173 (O_1173,N_21026,N_21494);
nand UO_1174 (O_1174,N_21565,N_24435);
and UO_1175 (O_1175,N_23595,N_23210);
xor UO_1176 (O_1176,N_22310,N_22888);
or UO_1177 (O_1177,N_21138,N_24219);
nor UO_1178 (O_1178,N_24276,N_22359);
nor UO_1179 (O_1179,N_20986,N_21952);
nor UO_1180 (O_1180,N_20976,N_23739);
nand UO_1181 (O_1181,N_20488,N_21928);
nor UO_1182 (O_1182,N_24511,N_21212);
or UO_1183 (O_1183,N_20215,N_22831);
or UO_1184 (O_1184,N_22689,N_20961);
xnor UO_1185 (O_1185,N_21046,N_21735);
or UO_1186 (O_1186,N_24902,N_24607);
xor UO_1187 (O_1187,N_20535,N_20901);
and UO_1188 (O_1188,N_24519,N_23753);
nand UO_1189 (O_1189,N_24552,N_22555);
nor UO_1190 (O_1190,N_22420,N_23762);
nor UO_1191 (O_1191,N_23338,N_22596);
or UO_1192 (O_1192,N_24760,N_21847);
and UO_1193 (O_1193,N_24698,N_22522);
nor UO_1194 (O_1194,N_21772,N_24878);
xor UO_1195 (O_1195,N_20511,N_21079);
nor UO_1196 (O_1196,N_21513,N_22714);
nor UO_1197 (O_1197,N_21469,N_21812);
or UO_1198 (O_1198,N_21275,N_21035);
xor UO_1199 (O_1199,N_21823,N_22695);
and UO_1200 (O_1200,N_22908,N_21953);
or UO_1201 (O_1201,N_22175,N_23749);
or UO_1202 (O_1202,N_23058,N_22294);
or UO_1203 (O_1203,N_21330,N_24551);
or UO_1204 (O_1204,N_24173,N_24315);
xor UO_1205 (O_1205,N_21891,N_21341);
nand UO_1206 (O_1206,N_23640,N_21887);
nand UO_1207 (O_1207,N_20121,N_21040);
and UO_1208 (O_1208,N_21581,N_24317);
and UO_1209 (O_1209,N_20016,N_23420);
nor UO_1210 (O_1210,N_22581,N_23866);
nor UO_1211 (O_1211,N_21049,N_21978);
and UO_1212 (O_1212,N_24125,N_22610);
or UO_1213 (O_1213,N_22050,N_23397);
xor UO_1214 (O_1214,N_20908,N_24727);
or UO_1215 (O_1215,N_22327,N_21519);
or UO_1216 (O_1216,N_24917,N_22060);
nor UO_1217 (O_1217,N_23854,N_20542);
nand UO_1218 (O_1218,N_21726,N_23796);
nor UO_1219 (O_1219,N_23104,N_22926);
or UO_1220 (O_1220,N_20311,N_23341);
and UO_1221 (O_1221,N_21433,N_24369);
and UO_1222 (O_1222,N_20017,N_22537);
and UO_1223 (O_1223,N_24687,N_22973);
or UO_1224 (O_1224,N_24759,N_24242);
nand UO_1225 (O_1225,N_20476,N_23831);
nor UO_1226 (O_1226,N_20037,N_23182);
and UO_1227 (O_1227,N_21628,N_21873);
nand UO_1228 (O_1228,N_23890,N_21386);
nand UO_1229 (O_1229,N_21618,N_20870);
and UO_1230 (O_1230,N_22218,N_24381);
nand UO_1231 (O_1231,N_20275,N_21625);
nand UO_1232 (O_1232,N_22621,N_21407);
nand UO_1233 (O_1233,N_23237,N_23487);
or UO_1234 (O_1234,N_23041,N_24514);
nand UO_1235 (O_1235,N_24811,N_22437);
nor UO_1236 (O_1236,N_20642,N_24341);
and UO_1237 (O_1237,N_24296,N_22820);
or UO_1238 (O_1238,N_20267,N_21505);
and UO_1239 (O_1239,N_23450,N_22252);
nor UO_1240 (O_1240,N_20009,N_23092);
or UO_1241 (O_1241,N_21037,N_24441);
or UO_1242 (O_1242,N_22646,N_23518);
or UO_1243 (O_1243,N_20813,N_22752);
nor UO_1244 (O_1244,N_22304,N_23706);
nor UO_1245 (O_1245,N_24952,N_24642);
nor UO_1246 (O_1246,N_24764,N_23731);
and UO_1247 (O_1247,N_23265,N_22546);
xor UO_1248 (O_1248,N_22485,N_21206);
xor UO_1249 (O_1249,N_22774,N_22334);
and UO_1250 (O_1250,N_21768,N_24013);
xnor UO_1251 (O_1251,N_21081,N_22842);
and UO_1252 (O_1252,N_24892,N_22590);
nand UO_1253 (O_1253,N_22748,N_20601);
nor UO_1254 (O_1254,N_22040,N_21158);
nor UO_1255 (O_1255,N_23680,N_22276);
nand UO_1256 (O_1256,N_24864,N_23482);
or UO_1257 (O_1257,N_24530,N_20219);
and UO_1258 (O_1258,N_21121,N_24758);
nand UO_1259 (O_1259,N_23636,N_24044);
nand UO_1260 (O_1260,N_22142,N_20051);
nor UO_1261 (O_1261,N_20374,N_21402);
xnor UO_1262 (O_1262,N_24007,N_20639);
or UO_1263 (O_1263,N_21561,N_24602);
and UO_1264 (O_1264,N_20572,N_20671);
nor UO_1265 (O_1265,N_23190,N_20144);
nor UO_1266 (O_1266,N_20039,N_22848);
xnor UO_1267 (O_1267,N_23497,N_20388);
and UO_1268 (O_1268,N_24335,N_23627);
and UO_1269 (O_1269,N_24393,N_23057);
nand UO_1270 (O_1270,N_20728,N_22883);
and UO_1271 (O_1271,N_22085,N_24726);
nor UO_1272 (O_1272,N_23788,N_20534);
nand UO_1273 (O_1273,N_20507,N_24379);
nand UO_1274 (O_1274,N_24407,N_24723);
or UO_1275 (O_1275,N_21232,N_23236);
or UO_1276 (O_1276,N_21267,N_24569);
xor UO_1277 (O_1277,N_20255,N_23787);
xnor UO_1278 (O_1278,N_21524,N_23935);
or UO_1279 (O_1279,N_20114,N_22481);
and UO_1280 (O_1280,N_22503,N_21572);
nand UO_1281 (O_1281,N_24110,N_21562);
and UO_1282 (O_1282,N_20564,N_20230);
nand UO_1283 (O_1283,N_23510,N_22872);
nand UO_1284 (O_1284,N_23738,N_21645);
and UO_1285 (O_1285,N_21785,N_21305);
xor UO_1286 (O_1286,N_20502,N_21897);
xor UO_1287 (O_1287,N_24385,N_24314);
nor UO_1288 (O_1288,N_20226,N_21022);
nor UO_1289 (O_1289,N_22937,N_20603);
nand UO_1290 (O_1290,N_24085,N_21892);
and UO_1291 (O_1291,N_21167,N_24290);
xnor UO_1292 (O_1292,N_21964,N_20445);
or UO_1293 (O_1293,N_21059,N_24390);
or UO_1294 (O_1294,N_24411,N_22575);
nor UO_1295 (O_1295,N_21097,N_21382);
or UO_1296 (O_1296,N_23183,N_21393);
nand UO_1297 (O_1297,N_24347,N_21116);
nand UO_1298 (O_1298,N_20568,N_24674);
and UO_1299 (O_1299,N_22286,N_23792);
and UO_1300 (O_1300,N_21655,N_22331);
and UO_1301 (O_1301,N_23431,N_22496);
or UO_1302 (O_1302,N_20998,N_24695);
xor UO_1303 (O_1303,N_20087,N_24563);
and UO_1304 (O_1304,N_23307,N_24548);
nand UO_1305 (O_1305,N_21518,N_22567);
nor UO_1306 (O_1306,N_23378,N_22899);
and UO_1307 (O_1307,N_20414,N_20605);
and UO_1308 (O_1308,N_20624,N_21481);
nor UO_1309 (O_1309,N_24880,N_23386);
and UO_1310 (O_1310,N_21170,N_21486);
and UO_1311 (O_1311,N_20652,N_21032);
nor UO_1312 (O_1312,N_20619,N_23263);
or UO_1313 (O_1313,N_24982,N_20295);
nand UO_1314 (O_1314,N_20234,N_23178);
and UO_1315 (O_1315,N_22452,N_21802);
or UO_1316 (O_1316,N_20264,N_21615);
and UO_1317 (O_1317,N_22395,N_22098);
or UO_1318 (O_1318,N_24461,N_22403);
xnor UO_1319 (O_1319,N_22152,N_22387);
xor UO_1320 (O_1320,N_23608,N_21235);
nor UO_1321 (O_1321,N_20322,N_23384);
and UO_1322 (O_1322,N_23932,N_24559);
xor UO_1323 (O_1323,N_21265,N_22885);
xor UO_1324 (O_1324,N_24993,N_21068);
nand UO_1325 (O_1325,N_22147,N_23919);
nor UO_1326 (O_1326,N_24680,N_20021);
nand UO_1327 (O_1327,N_22694,N_21710);
or UO_1328 (O_1328,N_21740,N_24130);
nand UO_1329 (O_1329,N_23511,N_20515);
or UO_1330 (O_1330,N_20310,N_24357);
xor UO_1331 (O_1331,N_21442,N_20705);
xor UO_1332 (O_1332,N_21463,N_24598);
and UO_1333 (O_1333,N_23931,N_21679);
or UO_1334 (O_1334,N_21409,N_23107);
or UO_1335 (O_1335,N_24157,N_22233);
and UO_1336 (O_1336,N_24673,N_24615);
and UO_1337 (O_1337,N_24469,N_21989);
and UO_1338 (O_1338,N_24809,N_23715);
or UO_1339 (O_1339,N_21296,N_20540);
and UO_1340 (O_1340,N_22041,N_21279);
and UO_1341 (O_1341,N_22574,N_24714);
and UO_1342 (O_1342,N_21154,N_21946);
xnor UO_1343 (O_1343,N_22043,N_22535);
xor UO_1344 (O_1344,N_24717,N_24067);
or UO_1345 (O_1345,N_24475,N_23782);
or UO_1346 (O_1346,N_23342,N_24761);
nor UO_1347 (O_1347,N_20560,N_21201);
nand UO_1348 (O_1348,N_24876,N_20406);
and UO_1349 (O_1349,N_22704,N_21800);
and UO_1350 (O_1350,N_21876,N_21598);
and UO_1351 (O_1351,N_20073,N_24772);
xnor UO_1352 (O_1352,N_22468,N_24897);
or UO_1353 (O_1353,N_21942,N_23778);
nor UO_1354 (O_1354,N_22795,N_22984);
nand UO_1355 (O_1355,N_24643,N_23446);
xnor UO_1356 (O_1356,N_23958,N_24595);
or UO_1357 (O_1357,N_23772,N_21630);
and UO_1358 (O_1358,N_21399,N_24405);
or UO_1359 (O_1359,N_20082,N_24126);
xnor UO_1360 (O_1360,N_21739,N_24353);
nor UO_1361 (O_1361,N_23223,N_24014);
nand UO_1362 (O_1362,N_23094,N_24868);
xor UO_1363 (O_1363,N_22637,N_24422);
xnor UO_1364 (O_1364,N_21151,N_22126);
xnor UO_1365 (O_1365,N_23808,N_24192);
nor UO_1366 (O_1366,N_22771,N_24106);
nor UO_1367 (O_1367,N_20280,N_20324);
xnor UO_1368 (O_1368,N_20638,N_22864);
or UO_1369 (O_1369,N_22736,N_20503);
nand UO_1370 (O_1370,N_22566,N_20035);
xnor UO_1371 (O_1371,N_20536,N_22684);
nand UO_1372 (O_1372,N_21817,N_23312);
or UO_1373 (O_1373,N_21925,N_21951);
and UO_1374 (O_1374,N_24722,N_23467);
and UO_1375 (O_1375,N_24579,N_20278);
and UO_1376 (O_1376,N_21084,N_22690);
nand UO_1377 (O_1377,N_20411,N_22587);
or UO_1378 (O_1378,N_21240,N_24416);
nand UO_1379 (O_1379,N_23807,N_20504);
or UO_1380 (O_1380,N_24894,N_20079);
nor UO_1381 (O_1381,N_20164,N_23688);
nor UO_1382 (O_1382,N_21763,N_21816);
nand UO_1383 (O_1383,N_24230,N_23075);
or UO_1384 (O_1384,N_22478,N_23781);
and UO_1385 (O_1385,N_22593,N_22051);
nand UO_1386 (O_1386,N_23149,N_22285);
nand UO_1387 (O_1387,N_22772,N_21353);
and UO_1388 (O_1388,N_23825,N_21941);
and UO_1389 (O_1389,N_20949,N_21041);
or UO_1390 (O_1390,N_23080,N_24458);
xnor UO_1391 (O_1391,N_21318,N_20719);
nor UO_1392 (O_1392,N_22122,N_24671);
xor UO_1393 (O_1393,N_23945,N_20885);
and UO_1394 (O_1394,N_20168,N_22417);
nand UO_1395 (O_1395,N_20434,N_20636);
xor UO_1396 (O_1396,N_22474,N_21231);
and UO_1397 (O_1397,N_24771,N_21972);
or UO_1398 (O_1398,N_20183,N_21236);
xor UO_1399 (O_1399,N_21736,N_20955);
nor UO_1400 (O_1400,N_24137,N_20841);
nor UO_1401 (O_1401,N_22259,N_23842);
nand UO_1402 (O_1402,N_21781,N_23158);
nand UO_1403 (O_1403,N_20513,N_21217);
nand UO_1404 (O_1404,N_23717,N_24538);
xor UO_1405 (O_1405,N_23466,N_24526);
nand UO_1406 (O_1406,N_21050,N_23650);
or UO_1407 (O_1407,N_24856,N_20779);
xor UO_1408 (O_1408,N_22900,N_23311);
xor UO_1409 (O_1409,N_21497,N_20608);
nor UO_1410 (O_1410,N_23068,N_21828);
nand UO_1411 (O_1411,N_23503,N_23521);
xor UO_1412 (O_1412,N_22833,N_23734);
xnor UO_1413 (O_1413,N_22732,N_23225);
and UO_1414 (O_1414,N_21052,N_22316);
nand UO_1415 (O_1415,N_21365,N_20265);
nand UO_1416 (O_1416,N_22008,N_23597);
nor UO_1417 (O_1417,N_21498,N_24490);
and UO_1418 (O_1418,N_23010,N_24193);
and UO_1419 (O_1419,N_23523,N_23989);
and UO_1420 (O_1420,N_24969,N_21932);
xnor UO_1421 (O_1421,N_21895,N_20637);
nor UO_1422 (O_1422,N_22116,N_24189);
or UO_1423 (O_1423,N_20292,N_24596);
xor UO_1424 (O_1424,N_24231,N_24155);
nor UO_1425 (O_1425,N_20849,N_23716);
and UO_1426 (O_1426,N_20353,N_24611);
nor UO_1427 (O_1427,N_23605,N_23153);
or UO_1428 (O_1428,N_24328,N_20721);
nor UO_1429 (O_1429,N_22279,N_20648);
or UO_1430 (O_1430,N_22857,N_23176);
nor UO_1431 (O_1431,N_23001,N_20356);
or UO_1432 (O_1432,N_20034,N_24035);
and UO_1433 (O_1433,N_20446,N_22602);
xor UO_1434 (O_1434,N_20065,N_21025);
or UO_1435 (O_1435,N_21592,N_22168);
or UO_1436 (O_1436,N_20799,N_20770);
or UO_1437 (O_1437,N_21879,N_24413);
nand UO_1438 (O_1438,N_24584,N_23202);
nor UO_1439 (O_1439,N_24793,N_21539);
nand UO_1440 (O_1440,N_24721,N_21464);
and UO_1441 (O_1441,N_20533,N_24360);
nand UO_1442 (O_1442,N_22245,N_20072);
and UO_1443 (O_1443,N_23232,N_22337);
xor UO_1444 (O_1444,N_23238,N_21637);
nand UO_1445 (O_1445,N_23361,N_22989);
and UO_1446 (O_1446,N_21431,N_23802);
nor UO_1447 (O_1447,N_24593,N_23230);
or UO_1448 (O_1448,N_20600,N_21291);
or UO_1449 (O_1449,N_23806,N_23611);
and UO_1450 (O_1450,N_21133,N_22227);
nand UO_1451 (O_1451,N_20400,N_24451);
nor UO_1452 (O_1452,N_22274,N_20402);
and UO_1453 (O_1453,N_23418,N_20929);
xor UO_1454 (O_1454,N_20662,N_23052);
and UO_1455 (O_1455,N_20754,N_21455);
or UO_1456 (O_1456,N_24253,N_23629);
or UO_1457 (O_1457,N_21119,N_24803);
nor UO_1458 (O_1458,N_21218,N_22380);
xor UO_1459 (O_1459,N_23118,N_21767);
and UO_1460 (O_1460,N_24321,N_22790);
and UO_1461 (O_1461,N_22136,N_23469);
nor UO_1462 (O_1462,N_22501,N_22199);
nor UO_1463 (O_1463,N_22155,N_20838);
nand UO_1464 (O_1464,N_23327,N_21839);
nand UO_1465 (O_1465,N_21227,N_20105);
nor UO_1466 (O_1466,N_22287,N_21060);
xnor UO_1467 (O_1467,N_24682,N_23809);
nand UO_1468 (O_1468,N_24280,N_24478);
nor UO_1469 (O_1469,N_22444,N_22852);
and UO_1470 (O_1470,N_22765,N_20200);
xor UO_1471 (O_1471,N_21987,N_22302);
nor UO_1472 (O_1472,N_20941,N_23322);
nand UO_1473 (O_1473,N_22987,N_23541);
xnor UO_1474 (O_1474,N_23613,N_22613);
xnor UO_1475 (O_1475,N_23952,N_21578);
xor UO_1476 (O_1476,N_20918,N_22240);
nand UO_1477 (O_1477,N_21286,N_23966);
or UO_1478 (O_1478,N_23901,N_21881);
xnor UO_1479 (O_1479,N_22078,N_23704);
xor UO_1480 (O_1480,N_24492,N_21351);
nor UO_1481 (O_1481,N_21315,N_20551);
or UO_1482 (O_1482,N_20663,N_24195);
nor UO_1483 (O_1483,N_23757,N_20956);
nand UO_1484 (O_1484,N_21183,N_20091);
nand UO_1485 (O_1485,N_22513,N_22494);
xnor UO_1486 (O_1486,N_20701,N_21435);
nor UO_1487 (O_1487,N_24662,N_23278);
and UO_1488 (O_1488,N_20058,N_22099);
or UO_1489 (O_1489,N_22639,N_23465);
xor UO_1490 (O_1490,N_22542,N_23148);
xnor UO_1491 (O_1491,N_20380,N_20212);
xnor UO_1492 (O_1492,N_22371,N_20131);
nor UO_1493 (O_1493,N_20075,N_23006);
nor UO_1494 (O_1494,N_23061,N_21515);
nor UO_1495 (O_1495,N_21591,N_22325);
nand UO_1496 (O_1496,N_20112,N_22592);
xnor UO_1497 (O_1497,N_22629,N_21703);
xor UO_1498 (O_1498,N_24966,N_20154);
nor UO_1499 (O_1499,N_21904,N_20174);
xnor UO_1500 (O_1500,N_21179,N_21551);
and UO_1501 (O_1501,N_24645,N_22739);
nand UO_1502 (O_1502,N_23310,N_24930);
nor UO_1503 (O_1503,N_23198,N_22548);
nor UO_1504 (O_1504,N_24524,N_22406);
and UO_1505 (O_1505,N_23124,N_23860);
nor UO_1506 (O_1506,N_23282,N_21247);
nor UO_1507 (O_1507,N_22110,N_20084);
nor UO_1508 (O_1508,N_20007,N_23641);
nand UO_1509 (O_1509,N_24196,N_21070);
or UO_1510 (O_1510,N_20365,N_22114);
xor UO_1511 (O_1511,N_23108,N_22551);
xnor UO_1512 (O_1512,N_22913,N_21108);
nand UO_1513 (O_1513,N_24638,N_22372);
and UO_1514 (O_1514,N_20610,N_24377);
xor UO_1515 (O_1515,N_22990,N_23639);
nor UO_1516 (O_1516,N_23632,N_22679);
nand UO_1517 (O_1517,N_20062,N_21264);
or UO_1518 (O_1518,N_22080,N_24046);
or UO_1519 (O_1519,N_24361,N_23908);
nor UO_1520 (O_1520,N_21284,N_24241);
and UO_1521 (O_1521,N_21770,N_24094);
and UO_1522 (O_1522,N_20694,N_24291);
nor UO_1523 (O_1523,N_22688,N_23723);
nor UO_1524 (O_1524,N_21924,N_24040);
and UO_1525 (O_1525,N_21670,N_22580);
nand UO_1526 (O_1526,N_20767,N_23930);
or UO_1527 (O_1527,N_20179,N_22495);
or UO_1528 (O_1528,N_23011,N_20195);
or UO_1529 (O_1529,N_21251,N_22455);
and UO_1530 (O_1530,N_22275,N_22445);
or UO_1531 (O_1531,N_21868,N_23022);
xnor UO_1532 (O_1532,N_22622,N_24020);
nor UO_1533 (O_1533,N_24664,N_24570);
and UO_1534 (O_1534,N_22049,N_22143);
nand UO_1535 (O_1535,N_24527,N_24343);
or UO_1536 (O_1536,N_20023,N_21349);
xnor UO_1537 (O_1537,N_22951,N_20824);
and UO_1538 (O_1538,N_20149,N_24363);
xor UO_1539 (O_1539,N_23529,N_24190);
and UO_1540 (O_1540,N_21425,N_21546);
or UO_1541 (O_1541,N_24083,N_23246);
or UO_1542 (O_1542,N_21501,N_21724);
nor UO_1543 (O_1543,N_23279,N_20421);
or UO_1544 (O_1544,N_23292,N_20250);
nand UO_1545 (O_1545,N_21673,N_24859);
and UO_1546 (O_1546,N_24229,N_20661);
nor UO_1547 (O_1547,N_20746,N_22097);
xor UO_1548 (O_1548,N_24523,N_23873);
nand UO_1549 (O_1549,N_21312,N_21995);
or UO_1550 (O_1550,N_24920,N_23391);
and UO_1551 (O_1551,N_20437,N_24319);
nand UO_1552 (O_1552,N_22839,N_23986);
or UO_1553 (O_1553,N_22750,N_21765);
nand UO_1554 (O_1554,N_23088,N_24730);
and UO_1555 (O_1555,N_20590,N_20225);
and UO_1556 (O_1556,N_22733,N_21412);
nor UO_1557 (O_1557,N_21397,N_22992);
nor UO_1558 (O_1558,N_22623,N_24149);
nor UO_1559 (O_1559,N_20866,N_23417);
and UO_1560 (O_1560,N_20050,N_23111);
or UO_1561 (O_1561,N_24132,N_24951);
or UO_1562 (O_1562,N_21799,N_20419);
and UO_1563 (O_1563,N_20811,N_20432);
nand UO_1564 (O_1564,N_21202,N_21335);
xor UO_1565 (O_1565,N_20877,N_24599);
and UO_1566 (O_1566,N_24281,N_21783);
nand UO_1567 (O_1567,N_21254,N_24283);
nor UO_1568 (O_1568,N_24997,N_23519);
xnor UO_1569 (O_1569,N_21205,N_22854);
nand UO_1570 (O_1570,N_21120,N_22638);
and UO_1571 (O_1571,N_20886,N_22059);
or UO_1572 (O_1572,N_23349,N_21849);
nor UO_1573 (O_1573,N_23551,N_23766);
nor UO_1574 (O_1574,N_22667,N_22995);
nand UO_1575 (O_1575,N_21310,N_24202);
nor UO_1576 (O_1576,N_21447,N_23858);
xnor UO_1577 (O_1577,N_23243,N_20415);
and UO_1578 (O_1578,N_22589,N_24228);
nand UO_1579 (O_1579,N_22034,N_23622);
nand UO_1580 (O_1580,N_22366,N_22363);
or UO_1581 (O_1581,N_24203,N_22802);
xnor UO_1582 (O_1582,N_20397,N_23150);
nand UO_1583 (O_1583,N_23745,N_24366);
xnor UO_1584 (O_1584,N_21074,N_23195);
xnor UO_1585 (O_1585,N_21188,N_22133);
or UO_1586 (O_1586,N_22185,N_23975);
and UO_1587 (O_1587,N_21098,N_20320);
or UO_1588 (O_1588,N_23147,N_23784);
xor UO_1589 (O_1589,N_24275,N_22144);
or UO_1590 (O_1590,N_21396,N_20101);
and UO_1591 (O_1591,N_23160,N_20740);
nor UO_1592 (O_1592,N_21820,N_22135);
or UO_1593 (O_1593,N_20580,N_20288);
and UO_1594 (O_1594,N_20778,N_21553);
xor UO_1595 (O_1595,N_21304,N_21261);
nand UO_1596 (O_1596,N_22118,N_22912);
xnor UO_1597 (O_1597,N_24806,N_24953);
and UO_1598 (O_1598,N_24777,N_20163);
and UO_1599 (O_1599,N_23333,N_24942);
nand UO_1600 (O_1600,N_22721,N_21024);
xnor UO_1601 (O_1601,N_21295,N_22433);
xnor UO_1602 (O_1602,N_21285,N_20379);
or UO_1603 (O_1603,N_23302,N_24348);
and UO_1604 (O_1604,N_24206,N_23032);
and UO_1605 (O_1605,N_22203,N_24711);
xnor UO_1606 (O_1606,N_24113,N_22393);
xor UO_1607 (O_1607,N_24724,N_20683);
xor UO_1608 (O_1608,N_24431,N_20330);
nand UO_1609 (O_1609,N_23289,N_23570);
xnor UO_1610 (O_1610,N_24056,N_23805);
or UO_1611 (O_1611,N_21141,N_22067);
nand UO_1612 (O_1612,N_21602,N_24337);
nor UO_1613 (O_1613,N_22915,N_20246);
nand UO_1614 (O_1614,N_24371,N_21058);
nor UO_1615 (O_1615,N_24140,N_24261);
nor UO_1616 (O_1616,N_24840,N_21162);
nor UO_1617 (O_1617,N_22471,N_22859);
nand UO_1618 (O_1618,N_22391,N_21475);
xnor UO_1619 (O_1619,N_21826,N_21582);
xor UO_1620 (O_1620,N_24858,N_24633);
or UO_1621 (O_1621,N_20345,N_23288);
xor UO_1622 (O_1622,N_24938,N_22006);
xnor UO_1623 (O_1623,N_20338,N_23746);
or UO_1624 (O_1624,N_21363,N_23697);
xor UO_1625 (O_1625,N_24076,N_20349);
xnor UO_1626 (O_1626,N_22812,N_22626);
nand UO_1627 (O_1627,N_23044,N_21177);
and UO_1628 (O_1628,N_20128,N_24041);
nand UO_1629 (O_1629,N_20482,N_24590);
or UO_1630 (O_1630,N_22536,N_21945);
and UO_1631 (O_1631,N_23977,N_20547);
and UO_1632 (O_1632,N_23452,N_24609);
nor UO_1633 (O_1633,N_23016,N_22955);
xor UO_1634 (O_1634,N_23979,N_21819);
and UO_1635 (O_1635,N_22686,N_23252);
and UO_1636 (O_1636,N_23073,N_24837);
or UO_1637 (O_1637,N_23200,N_21016);
nor UO_1638 (O_1638,N_21088,N_22897);
xor UO_1639 (O_1639,N_22821,N_22956);
xor UO_1640 (O_1640,N_24573,N_24120);
and UO_1641 (O_1641,N_24380,N_21012);
nor UO_1642 (O_1642,N_20574,N_23027);
or UO_1643 (O_1643,N_20843,N_20806);
or UO_1644 (O_1644,N_20455,N_20006);
xor UO_1645 (O_1645,N_22253,N_23803);
xor UO_1646 (O_1646,N_21164,N_24796);
nor UO_1647 (O_1647,N_22381,N_23364);
xor UO_1648 (O_1648,N_24180,N_22449);
nor UO_1649 (O_1649,N_22225,N_20192);
nor UO_1650 (O_1650,N_21704,N_22860);
xnor UO_1651 (O_1651,N_22767,N_22145);
or UO_1652 (O_1652,N_22945,N_20475);
or UO_1653 (O_1653,N_20333,N_21472);
nor UO_1654 (O_1654,N_22105,N_24766);
and UO_1655 (O_1655,N_23197,N_23389);
nand UO_1656 (O_1656,N_21718,N_20609);
xor UO_1657 (O_1657,N_24087,N_23212);
nand UO_1658 (O_1658,N_21737,N_20989);
nand UO_1659 (O_1659,N_23625,N_20970);
nand UO_1660 (O_1660,N_21787,N_24826);
xnor UO_1661 (O_1661,N_23939,N_20162);
xor UO_1662 (O_1662,N_24415,N_22039);
nor UO_1663 (O_1663,N_22887,N_20553);
xnor UO_1664 (O_1664,N_22661,N_24260);
xor UO_1665 (O_1665,N_24541,N_22604);
xor UO_1666 (O_1666,N_24081,N_24578);
nor UO_1667 (O_1667,N_22855,N_24011);
nand UO_1668 (O_1668,N_22421,N_23367);
nor UO_1669 (O_1669,N_20211,N_22027);
nor UO_1670 (O_1670,N_23249,N_24470);
nand UO_1671 (O_1671,N_23612,N_23416);
or UO_1672 (O_1672,N_20790,N_24147);
nor UO_1673 (O_1673,N_23871,N_21053);
nor UO_1674 (O_1674,N_20002,N_20625);
nand UO_1675 (O_1675,N_20473,N_21400);
or UO_1676 (O_1676,N_21880,N_20157);
and UO_1677 (O_1677,N_24047,N_24313);
or UO_1678 (O_1678,N_24678,N_23539);
or UO_1679 (O_1679,N_23635,N_22413);
nand UO_1680 (O_1680,N_20514,N_23546);
and UO_1681 (O_1681,N_21362,N_23524);
xor UO_1682 (O_1682,N_21357,N_22376);
xor UO_1683 (O_1683,N_23686,N_20968);
nand UO_1684 (O_1684,N_23266,N_21458);
nor UO_1685 (O_1685,N_20831,N_23794);
and UO_1686 (O_1686,N_23480,N_23761);
nor UO_1687 (O_1687,N_20399,N_24998);
nand UO_1688 (O_1688,N_21559,N_24010);
nand UO_1689 (O_1689,N_24546,N_24171);
nand UO_1690 (O_1690,N_23483,N_20177);
nor UO_1691 (O_1691,N_24122,N_23273);
xnor UO_1692 (O_1692,N_20279,N_21328);
xnor UO_1693 (O_1693,N_22093,N_23498);
xnor UO_1694 (O_1694,N_21976,N_22033);
nor UO_1695 (O_1695,N_23023,N_22741);
xor UO_1696 (O_1696,N_21129,N_23332);
xnor UO_1697 (O_1697,N_22378,N_22255);
or UO_1698 (O_1698,N_23428,N_24384);
or UO_1699 (O_1699,N_23369,N_21454);
nor UO_1700 (O_1700,N_21754,N_23801);
and UO_1701 (O_1701,N_24939,N_22827);
nand UO_1702 (O_1702,N_24934,N_21913);
xor UO_1703 (O_1703,N_24383,N_24444);
and UO_1704 (O_1704,N_24965,N_21047);
and UO_1705 (O_1705,N_21078,N_20606);
nor UO_1706 (O_1706,N_24075,N_23556);
nand UO_1707 (O_1707,N_24268,N_23536);
nand UO_1708 (O_1708,N_22867,N_22210);
or UO_1709 (O_1709,N_23719,N_20096);
or UO_1710 (O_1710,N_21419,N_20567);
xnor UO_1711 (O_1711,N_22598,N_23189);
or UO_1712 (O_1712,N_20702,N_22530);
or UO_1713 (O_1713,N_24182,N_24744);
xor UO_1714 (O_1714,N_24188,N_24984);
and UO_1715 (O_1715,N_20569,N_23065);
nor UO_1716 (O_1716,N_23593,N_22453);
nor UO_1717 (O_1717,N_24960,N_22541);
nand UO_1718 (O_1718,N_20393,N_22192);
nor UO_1719 (O_1719,N_24742,N_24648);
and UO_1720 (O_1720,N_20059,N_20835);
and UO_1721 (O_1721,N_21548,N_21845);
xnor UO_1722 (O_1722,N_22241,N_20194);
xor UO_1723 (O_1723,N_24170,N_24663);
and UO_1724 (O_1724,N_20442,N_22692);
nor UO_1725 (O_1725,N_23206,N_24216);
xor UO_1726 (O_1726,N_22169,N_24533);
nand UO_1727 (O_1727,N_22550,N_24732);
nand UO_1728 (O_1728,N_24166,N_24320);
and UO_1729 (O_1729,N_22159,N_24430);
xnor UO_1730 (O_1730,N_24288,N_23771);
nor UO_1731 (O_1731,N_21555,N_21732);
nor UO_1732 (O_1732,N_23972,N_24995);
or UO_1733 (O_1733,N_21443,N_24251);
xor UO_1734 (O_1734,N_21439,N_22134);
nand UO_1735 (O_1735,N_20951,N_20465);
nor UO_1736 (O_1736,N_22460,N_22861);
nand UO_1737 (O_1737,N_22976,N_20172);
nor UO_1738 (O_1738,N_20739,N_23056);
xnor UO_1739 (O_1739,N_20489,N_24525);
xnor UO_1740 (O_1740,N_20375,N_21346);
or UO_1741 (O_1741,N_22011,N_23129);
nor UO_1742 (O_1742,N_21198,N_23233);
and UO_1743 (O_1743,N_22058,N_20520);
nand UO_1744 (O_1744,N_21950,N_21003);
nor UO_1745 (O_1745,N_20899,N_20724);
nor UO_1746 (O_1746,N_21374,N_20008);
and UO_1747 (O_1747,N_20629,N_22388);
nand UO_1748 (O_1748,N_21473,N_22349);
or UO_1749 (O_1749,N_24434,N_23244);
nor UO_1750 (O_1750,N_22809,N_21706);
xor UO_1751 (O_1751,N_22472,N_24082);
or UO_1752 (O_1752,N_21651,N_23119);
or UO_1753 (O_1753,N_22504,N_20807);
nor UO_1754 (O_1754,N_23572,N_20771);
nor UO_1755 (O_1755,N_22345,N_23360);
or UO_1756 (O_1756,N_20176,N_21007);
and UO_1757 (O_1757,N_20368,N_21681);
and UO_1758 (O_1758,N_21741,N_22186);
nand UO_1759 (O_1759,N_21644,N_23637);
and UO_1760 (O_1760,N_23855,N_20360);
and UO_1761 (O_1761,N_21195,N_23631);
nor UO_1762 (O_1762,N_23248,N_22120);
xnor UO_1763 (O_1763,N_23258,N_22194);
xor UO_1764 (O_1764,N_24292,N_23579);
nor UO_1765 (O_1765,N_24940,N_21209);
nor UO_1766 (O_1766,N_20306,N_22178);
nand UO_1767 (O_1767,N_23649,N_21537);
nor UO_1768 (O_1768,N_22803,N_22130);
nand UO_1769 (O_1769,N_21028,N_23814);
nand UO_1770 (O_1770,N_22730,N_24052);
xor UO_1771 (O_1771,N_22211,N_21502);
and UO_1772 (O_1772,N_22411,N_24350);
nand UO_1773 (O_1773,N_21850,N_21761);
nor UO_1774 (O_1774,N_21764,N_24019);
and UO_1775 (O_1775,N_23921,N_24873);
or UO_1776 (O_1776,N_20856,N_20453);
and UO_1777 (O_1777,N_23985,N_20710);
or UO_1778 (O_1778,N_22369,N_22031);
nor UO_1779 (O_1779,N_23672,N_21176);
xnor UO_1780 (O_1780,N_22584,N_22879);
nand UO_1781 (O_1781,N_22869,N_24767);
xnor UO_1782 (O_1782,N_24627,N_21361);
xor UO_1783 (O_1783,N_20014,N_22007);
or UO_1784 (O_1784,N_20788,N_21221);
and UO_1785 (O_1785,N_22200,N_20000);
nand UO_1786 (O_1786,N_22029,N_23578);
nand UO_1787 (O_1787,N_20086,N_22904);
or UO_1788 (O_1788,N_23081,N_23667);
nor UO_1789 (O_1789,N_20327,N_21277);
nand UO_1790 (O_1790,N_22422,N_21857);
and UO_1791 (O_1791,N_21269,N_20069);
xor UO_1792 (O_1792,N_22815,N_20800);
nand UO_1793 (O_1793,N_22222,N_24676);
nor UO_1794 (O_1794,N_20071,N_23675);
nand UO_1795 (O_1795,N_22140,N_24550);
or UO_1796 (O_1796,N_22088,N_22336);
and UO_1797 (O_1797,N_20190,N_22822);
xnor UO_1798 (O_1798,N_24820,N_21095);
xor UO_1799 (O_1799,N_21062,N_22052);
nor UO_1800 (O_1800,N_20526,N_21533);
xor UO_1801 (O_1801,N_22917,N_21441);
and UO_1802 (O_1802,N_20990,N_23157);
xor UO_1803 (O_1803,N_24287,N_20387);
or UO_1804 (O_1804,N_21023,N_23591);
or UO_1805 (O_1805,N_22429,N_21159);
or UO_1806 (O_1806,N_20865,N_20024);
or UO_1807 (O_1807,N_22665,N_24402);
and UO_1808 (O_1808,N_20693,N_24159);
nand UO_1809 (O_1809,N_24553,N_21683);
xnor UO_1810 (O_1810,N_22483,N_20430);
xnor UO_1811 (O_1811,N_23366,N_22543);
and UO_1812 (O_1812,N_21069,N_20665);
nand UO_1813 (O_1813,N_22728,N_20834);
and UO_1814 (O_1814,N_22026,N_24705);
xnor UO_1815 (O_1815,N_24323,N_24086);
and UO_1816 (O_1816,N_21244,N_23644);
and UO_1817 (O_1817,N_24962,N_22863);
and UO_1818 (O_1818,N_24001,N_21114);
xor UO_1819 (O_1819,N_24529,N_24426);
nand UO_1820 (O_1820,N_23262,N_21629);
and UO_1821 (O_1821,N_22115,N_22866);
xor UO_1822 (O_1822,N_20848,N_22298);
xnor UO_1823 (O_1823,N_24312,N_22776);
or UO_1824 (O_1824,N_24179,N_23581);
or UO_1825 (O_1825,N_23296,N_20390);
xnor UO_1826 (O_1826,N_23239,N_24833);
nand UO_1827 (O_1827,N_21080,N_23623);
xnor UO_1828 (O_1828,N_21960,N_23114);
and UO_1829 (O_1829,N_20339,N_20428);
nand UO_1830 (O_1830,N_23501,N_23555);
xor UO_1831 (O_1831,N_23900,N_23689);
nor UO_1832 (O_1832,N_24351,N_24677);
xnor UO_1833 (O_1833,N_23123,N_20077);
nor UO_1834 (O_1834,N_24817,N_24263);
nand UO_1835 (O_1835,N_21918,N_24634);
and UO_1836 (O_1836,N_20696,N_24455);
nor UO_1837 (O_1837,N_20304,N_22949);
or UO_1838 (O_1838,N_21169,N_22153);
or UO_1839 (O_1839,N_22399,N_20435);
xnor UO_1840 (O_1840,N_23226,N_23951);
or UO_1841 (O_1841,N_24151,N_24540);
xor UO_1842 (O_1842,N_24374,N_22351);
nor UO_1843 (O_1843,N_22082,N_24500);
xnor UO_1844 (O_1844,N_21723,N_22068);
nor UO_1845 (O_1845,N_23376,N_23039);
or UO_1846 (O_1846,N_23304,N_21603);
nor UO_1847 (O_1847,N_22939,N_22191);
nand UO_1848 (O_1848,N_21947,N_22591);
nand UO_1849 (O_1849,N_20370,N_24707);
and UO_1850 (O_1850,N_24443,N_24718);
or UO_1851 (O_1851,N_23188,N_23642);
xnor UO_1852 (O_1852,N_20220,N_24409);
or UO_1853 (O_1853,N_23425,N_20291);
and UO_1854 (O_1854,N_24844,N_21325);
xnor UO_1855 (O_1855,N_22896,N_22703);
nand UO_1856 (O_1856,N_24954,N_21846);
nor UO_1857 (O_1857,N_23174,N_21470);
xnor UO_1858 (O_1858,N_21574,N_20207);
nand UO_1859 (O_1859,N_21956,N_21930);
or UO_1860 (O_1860,N_20481,N_20496);
xor UO_1861 (O_1861,N_22022,N_22469);
nor UO_1862 (O_1862,N_23115,N_21257);
or UO_1863 (O_1863,N_23375,N_21642);
xnor UO_1864 (O_1864,N_20263,N_20376);
or UO_1865 (O_1865,N_20301,N_22644);
xor UO_1866 (O_1866,N_22077,N_22615);
xor UO_1867 (O_1867,N_23574,N_22936);
nor UO_1868 (O_1868,N_23571,N_20425);
and UO_1869 (O_1869,N_21476,N_23260);
and UO_1870 (O_1870,N_20218,N_24802);
xor UO_1871 (O_1871,N_23087,N_23381);
or UO_1872 (O_1872,N_23211,N_20110);
and UO_1873 (O_1873,N_22583,N_22727);
or UO_1874 (O_1874,N_22340,N_24119);
or UO_1875 (O_1875,N_24295,N_21180);
or UO_1876 (O_1876,N_22235,N_22443);
xnor UO_1877 (O_1877,N_21611,N_22261);
or UO_1878 (O_1878,N_20798,N_20299);
nor UO_1879 (O_1879,N_22873,N_20934);
nor UO_1880 (O_1880,N_20193,N_23405);
nand UO_1881 (O_1881,N_21701,N_22092);
xnor UO_1882 (O_1882,N_24420,N_21647);
and UO_1883 (O_1883,N_24807,N_21302);
and UO_1884 (O_1884,N_21427,N_22370);
nor UO_1885 (O_1885,N_24400,N_23943);
and UO_1886 (O_1886,N_22702,N_22164);
xor UO_1887 (O_1887,N_20797,N_23614);
xnor UO_1888 (O_1888,N_24585,N_21128);
nor UO_1889 (O_1889,N_22789,N_20622);
nor UO_1890 (O_1890,N_20169,N_20229);
xnor UO_1891 (O_1891,N_20858,N_20764);
nand UO_1892 (O_1892,N_23652,N_22103);
xnor UO_1893 (O_1893,N_24143,N_22711);
and UO_1894 (O_1894,N_23084,N_24750);
nand UO_1895 (O_1895,N_23526,N_20565);
xnor UO_1896 (O_1896,N_21384,N_20204);
and UO_1897 (O_1897,N_23455,N_20308);
nand UO_1898 (O_1898,N_22400,N_20243);
or UO_1899 (O_1899,N_24378,N_21593);
nand UO_1900 (O_1900,N_21520,N_22797);
and UO_1901 (O_1901,N_24649,N_22729);
nor UO_1902 (O_1902,N_23708,N_22017);
or UO_1903 (O_1903,N_22554,N_22436);
and UO_1904 (O_1904,N_22526,N_20117);
or UO_1905 (O_1905,N_24829,N_22882);
or UO_1906 (O_1906,N_23004,N_21535);
nand UO_1907 (O_1907,N_20852,N_24983);
nor UO_1908 (O_1908,N_20726,N_24359);
nand UO_1909 (O_1909,N_24096,N_24223);
or UO_1910 (O_1910,N_21751,N_20789);
nor UO_1911 (O_1911,N_20966,N_23916);
or UO_1912 (O_1912,N_24037,N_20632);
nor UO_1913 (O_1913,N_23879,N_21160);
xnor UO_1914 (O_1914,N_21769,N_20160);
xor UO_1915 (O_1915,N_22983,N_23172);
or UO_1916 (O_1916,N_24158,N_21253);
nand UO_1917 (O_1917,N_22958,N_23647);
xnor UO_1918 (O_1918,N_24558,N_23560);
nand UO_1919 (O_1919,N_21694,N_21899);
or UO_1920 (O_1920,N_23743,N_24531);
xor UO_1921 (O_1921,N_20523,N_22562);
nand UO_1922 (O_1922,N_23191,N_21639);
nor UO_1923 (O_1923,N_20867,N_23603);
or UO_1924 (O_1924,N_24038,N_22405);
or UO_1925 (O_1925,N_23646,N_23101);
and UO_1926 (O_1926,N_23638,N_23775);
nor UO_1927 (O_1927,N_21832,N_21753);
and UO_1928 (O_1928,N_23910,N_24065);
or UO_1929 (O_1929,N_24914,N_23187);
and UO_1930 (O_1930,N_22576,N_22347);
or UO_1931 (O_1931,N_22620,N_22705);
nand UO_1932 (O_1932,N_22746,N_20439);
nand UO_1933 (O_1933,N_24949,N_24238);
and UO_1934 (O_1934,N_21440,N_21504);
xnor UO_1935 (O_1935,N_24432,N_23948);
and UO_1936 (O_1936,N_21675,N_22761);
and UO_1937 (O_1937,N_20731,N_21929);
nor UO_1938 (O_1938,N_22102,N_24497);
nor UO_1939 (O_1939,N_23677,N_21654);
nand UO_1940 (O_1940,N_24600,N_24024);
and UO_1941 (O_1941,N_22600,N_20262);
or UO_1942 (O_1942,N_20892,N_22806);
and UO_1943 (O_1943,N_24637,N_22268);
xnor UO_1944 (O_1944,N_20544,N_20472);
xor UO_1945 (O_1945,N_23520,N_20251);
nand UO_1946 (O_1946,N_21595,N_20883);
nand UO_1947 (O_1947,N_20383,N_23710);
nand UO_1948 (O_1948,N_23533,N_22745);
or UO_1949 (O_1949,N_20646,N_20404);
or UO_1950 (O_1950,N_24114,N_23343);
xnor UO_1951 (O_1951,N_24936,N_24236);
and UO_1952 (O_1952,N_23779,N_21422);
nor UO_1953 (O_1953,N_20782,N_24824);
xor UO_1954 (O_1954,N_22923,N_23856);
or UO_1955 (O_1955,N_24955,N_21014);
nor UO_1956 (O_1956,N_21298,N_21018);
nand UO_1957 (O_1957,N_23385,N_21044);
or UO_1958 (O_1958,N_22775,N_22934);
nand UO_1959 (O_1959,N_22652,N_23344);
nand UO_1960 (O_1960,N_23291,N_24597);
xnor UO_1961 (O_1961,N_23528,N_24852);
and UO_1962 (O_1962,N_20864,N_22032);
nand UO_1963 (O_1963,N_22807,N_23513);
xnor UO_1964 (O_1964,N_20910,N_24791);
or UO_1965 (O_1965,N_21466,N_22081);
nand UO_1966 (O_1966,N_20552,N_21272);
xnor UO_1967 (O_1967,N_23145,N_22505);
nand UO_1968 (O_1968,N_20999,N_22138);
or UO_1969 (O_1969,N_24757,N_23750);
nor UO_1970 (O_1970,N_23277,N_23067);
nand UO_1971 (O_1971,N_22066,N_23616);
nand UO_1972 (O_1972,N_20381,N_22063);
and UO_1973 (O_1973,N_20851,N_21834);
nand UO_1974 (O_1974,N_22216,N_22846);
xor UO_1975 (O_1975,N_22465,N_22195);
nand UO_1976 (O_1976,N_21089,N_20019);
nand UO_1977 (O_1977,N_20045,N_24033);
nand UO_1978 (O_1978,N_23468,N_21438);
nand UO_1979 (O_1979,N_20022,N_21110);
xnor UO_1980 (O_1980,N_20236,N_20736);
nor UO_1981 (O_1981,N_22707,N_23651);
or UO_1982 (O_1982,N_20378,N_23517);
nor UO_1983 (O_1983,N_21729,N_21460);
or UO_1984 (O_1984,N_21292,N_23030);
and UO_1985 (O_1985,N_23777,N_22074);
and UO_1986 (O_1986,N_20978,N_20974);
nand UO_1987 (O_1987,N_22903,N_23718);
nor UO_1988 (O_1988,N_24589,N_21921);
or UO_1989 (O_1989,N_23577,N_21560);
and UO_1990 (O_1990,N_22636,N_24557);
or UO_1991 (O_1991,N_21391,N_20118);
nor UO_1992 (O_1992,N_21931,N_23215);
xor UO_1993 (O_1993,N_20562,N_21348);
xnor UO_1994 (O_1994,N_24340,N_23462);
or UO_1995 (O_1995,N_23029,N_23286);
xnor UO_1996 (O_1996,N_21187,N_22202);
or UO_1997 (O_1997,N_20967,N_24410);
and UO_1998 (O_1998,N_24623,N_22368);
and UO_1999 (O_1999,N_21338,N_20819);
xor UO_2000 (O_2000,N_23509,N_24703);
nand UO_2001 (O_2001,N_20426,N_20074);
nor UO_2002 (O_2002,N_24555,N_24464);
or UO_2003 (O_2003,N_24957,N_20627);
or UO_2004 (O_2004,N_21071,N_21238);
nand UO_2005 (O_2005,N_24142,N_24684);
xor UO_2006 (O_2006,N_22269,N_24175);
nand UO_2007 (O_2007,N_20343,N_22898);
or UO_2008 (O_2008,N_24499,N_20364);
or UO_2009 (O_2009,N_21326,N_22751);
or UO_2010 (O_2010,N_22457,N_21336);
or UO_2011 (O_2011,N_23882,N_21959);
nor UO_2012 (O_2012,N_20490,N_20654);
xor UO_2013 (O_2013,N_22735,N_22784);
xor UO_2014 (O_2014,N_24898,N_24753);
xor UO_2015 (O_2015,N_20371,N_24716);
nor UO_2016 (O_2016,N_23445,N_22871);
xnor UO_2017 (O_2017,N_23363,N_24212);
xor UO_2018 (O_2018,N_20570,N_20134);
nor UO_2019 (O_2019,N_22657,N_20945);
and UO_2020 (O_2020,N_23681,N_20261);
and UO_2021 (O_2021,N_20549,N_20237);
or UO_2022 (O_2022,N_23826,N_20839);
nor UO_2023 (O_2023,N_20587,N_20173);
xnor UO_2024 (O_2024,N_20321,N_23457);
or UO_2025 (O_2025,N_21413,N_20761);
nand UO_2026 (O_2026,N_24668,N_23590);
nor UO_2027 (O_2027,N_24072,N_23410);
and UO_2028 (O_2028,N_23655,N_20925);
xor UO_2029 (O_2029,N_23368,N_24412);
and UO_2030 (O_2030,N_22293,N_20336);
nor UO_2031 (O_2031,N_21659,N_24237);
and UO_2032 (O_2032,N_22459,N_24847);
nor UO_2033 (O_2033,N_23063,N_22793);
or UO_2034 (O_2034,N_23448,N_23835);
xor UO_2035 (O_2035,N_24224,N_24306);
nor UO_2036 (O_2036,N_24482,N_24027);
nor UO_2037 (O_2037,N_21682,N_21001);
and UO_2038 (O_2038,N_22148,N_24121);
nand UO_2039 (O_2039,N_21547,N_20217);
nand UO_2040 (O_2040,N_22094,N_23346);
xnor UO_2041 (O_2041,N_24762,N_23313);
xnor UO_2042 (O_2042,N_20480,N_21671);
and UO_2043 (O_2043,N_22642,N_24882);
and UO_2044 (O_2044,N_21752,N_23308);
or UO_2045 (O_2045,N_23917,N_24396);
nor UO_2046 (O_2046,N_24821,N_23130);
or UO_2047 (O_2047,N_20658,N_21043);
or UO_2048 (O_2048,N_24138,N_22858);
or UO_2049 (O_2049,N_20314,N_22344);
and UO_2050 (O_2050,N_21949,N_23447);
nor UO_2051 (O_2051,N_20350,N_21612);
nand UO_2052 (O_2052,N_21436,N_22738);
and UO_2053 (O_2053,N_22442,N_23036);
xnor UO_2054 (O_2054,N_23789,N_22065);
or UO_2055 (O_2055,N_24172,N_21011);
xnor UO_2056 (O_2056,N_22744,N_23021);
nor UO_2057 (O_2057,N_20494,N_24115);
xor UO_2058 (O_2058,N_24618,N_21228);
nor UO_2059 (O_2059,N_20066,N_21036);
and UO_2060 (O_2060,N_23722,N_24247);
xor UO_2061 (O_2061,N_21871,N_22843);
nand UO_2062 (O_2062,N_23463,N_22196);
or UO_2063 (O_2063,N_23727,N_20409);
or UO_2064 (O_2064,N_22101,N_21590);
and UO_2065 (O_2065,N_23602,N_24768);
or UO_2066 (O_2066,N_23491,N_23845);
nand UO_2067 (O_2067,N_20459,N_24116);
nor UO_2068 (O_2068,N_22283,N_23143);
and UO_2069 (O_2069,N_20575,N_22640);
and UO_2070 (O_2070,N_22323,N_20594);
xor UO_2071 (O_2071,N_20997,N_21552);
and UO_2072 (O_2072,N_21827,N_21903);
xor UO_2073 (O_2073,N_20707,N_23336);
or UO_2074 (O_2074,N_22426,N_23128);
nor UO_2075 (O_2075,N_22691,N_24373);
nand UO_2076 (O_2076,N_24741,N_20501);
and UO_2077 (O_2077,N_23763,N_24731);
or UO_2078 (O_2078,N_20994,N_20548);
xor UO_2079 (O_2079,N_20053,N_20403);
nor UO_2080 (O_2080,N_23012,N_23846);
or UO_2081 (O_2081,N_22214,N_24008);
nand UO_2082 (O_2082,N_22511,N_20395);
nand UO_2083 (O_2083,N_21416,N_21203);
and UO_2084 (O_2084,N_20996,N_22826);
nand UO_2085 (O_2085,N_20881,N_22617);
and UO_2086 (O_2086,N_24786,N_20919);
xor UO_2087 (O_2087,N_23683,N_21678);
and UO_2088 (O_2088,N_24690,N_22458);
xor UO_2089 (O_2089,N_22792,N_24318);
and UO_2090 (O_2090,N_23380,N_20272);
nand UO_2091 (O_2091,N_24996,N_20787);
nor UO_2092 (O_2092,N_22167,N_24439);
and UO_2093 (O_2093,N_22528,N_23893);
nor UO_2094 (O_2094,N_23076,N_22894);
nor UO_2095 (O_2095,N_24498,N_22341);
nor UO_2096 (O_2096,N_20142,N_22500);
and UO_2097 (O_2097,N_20325,N_22055);
nor UO_2098 (O_2098,N_24888,N_24667);
and UO_2099 (O_2099,N_20070,N_21477);
or UO_2100 (O_2100,N_22607,N_21948);
and UO_2101 (O_2101,N_24436,N_20416);
nand UO_2102 (O_2102,N_24665,N_22288);
nor UO_2103 (O_2103,N_22948,N_21153);
xor UO_2104 (O_2104,N_23131,N_22966);
nand UO_2105 (O_2105,N_21773,N_24870);
or UO_2106 (O_2106,N_20167,N_24226);
and UO_2107 (O_2107,N_24814,N_21452);
nor UO_2108 (O_2108,N_21837,N_22938);
or UO_2109 (O_2109,N_24401,N_24005);
nor UO_2110 (O_2110,N_23071,N_22221);
xnor UO_2111 (O_2111,N_21543,N_23261);
or UO_2112 (O_2112,N_22849,N_20479);
nand UO_2113 (O_2113,N_22828,N_20939);
nor UO_2114 (O_2114,N_21632,N_23356);
and UO_2115 (O_2115,N_24785,N_20089);
or UO_2116 (O_2116,N_24825,N_23293);
or UO_2117 (O_2117,N_22627,N_23522);
and UO_2118 (O_2118,N_20527,N_24387);
xor UO_2119 (O_2119,N_22397,N_22957);
or UO_2120 (O_2120,N_21985,N_21744);
xnor UO_2121 (O_2121,N_22643,N_22762);
and UO_2122 (O_2122,N_24879,N_24344);
and UO_2123 (O_2123,N_20979,N_20124);
nand UO_2124 (O_2124,N_23839,N_23274);
or UO_2125 (O_2125,N_23000,N_24070);
nor UO_2126 (O_2126,N_24980,N_24783);
and UO_2127 (O_2127,N_23186,N_20030);
xor UO_2128 (O_2128,N_20983,N_22057);
xnor UO_2129 (O_2129,N_21031,N_22184);
or UO_2130 (O_2130,N_23516,N_23018);
and UO_2131 (O_2131,N_20106,N_23326);
and UO_2132 (O_2132,N_21969,N_20281);
xor UO_2133 (O_2133,N_23019,N_20932);
nor UO_2134 (O_2134,N_22280,N_21587);
or UO_2135 (O_2135,N_24118,N_21750);
nand UO_2136 (O_2136,N_20923,N_20585);
and UO_2137 (O_2137,N_22649,N_22190);
or UO_2138 (O_2138,N_23402,N_23626);
nor UO_2139 (O_2139,N_22448,N_24831);
or UO_2140 (O_2140,N_24244,N_23984);
xor UO_2141 (O_2141,N_22488,N_24921);
xor UO_2142 (O_2142,N_22357,N_20495);
and UO_2143 (O_2143,N_24813,N_24403);
and UO_2144 (O_2144,N_24893,N_24485);
and UO_2145 (O_2145,N_20317,N_24282);
or UO_2146 (O_2146,N_20959,N_24910);
and UO_2147 (O_2147,N_21821,N_24532);
and UO_2148 (O_2148,N_22313,N_22630);
and UO_2149 (O_2149,N_22044,N_21106);
nand UO_2150 (O_2150,N_23915,N_24916);
or UO_2151 (O_2151,N_20245,N_23812);
nand UO_2152 (O_2152,N_20820,N_21297);
nor UO_2153 (O_2153,N_22814,N_23295);
xnor UO_2154 (O_2154,N_21370,N_21367);
and UO_2155 (O_2155,N_21746,N_23069);
and UO_2156 (O_2156,N_24176,N_23941);
and UO_2157 (O_2157,N_22154,N_24213);
xnor UO_2158 (O_2158,N_23615,N_21444);
and UO_2159 (O_2159,N_23495,N_21992);
nor UO_2160 (O_2160,N_23045,N_22559);
xor UO_2161 (O_2161,N_23043,N_24795);
nor UO_2162 (O_2162,N_24641,N_22669);
or UO_2163 (O_2163,N_21448,N_23878);
and UO_2164 (O_2164,N_21580,N_21389);
nor UO_2165 (O_2165,N_24307,N_20611);
nor UO_2166 (O_2166,N_22410,N_20063);
nand UO_2167 (O_2167,N_24051,N_21709);
nor UO_2168 (O_2168,N_21281,N_20781);
nand UO_2169 (O_2169,N_24471,N_24370);
or UO_2170 (O_2170,N_20102,N_21838);
or UO_2171 (O_2171,N_20452,N_24507);
nor UO_2172 (O_2172,N_23166,N_24853);
nand UO_2173 (O_2173,N_22419,N_21830);
nor UO_2174 (O_2174,N_23339,N_22435);
or UO_2175 (O_2175,N_24700,N_21534);
xnor UO_2176 (O_2176,N_22996,N_23936);
nand UO_2177 (O_2177,N_23408,N_24168);
xnor UO_2178 (O_2178,N_21144,N_24566);
nor UO_2179 (O_2179,N_20981,N_20361);
and UO_2180 (O_2180,N_24616,N_23817);
or UO_2181 (O_2181,N_22014,N_24109);
xnor UO_2182 (O_2182,N_23824,N_24908);
and UO_2183 (O_2183,N_20484,N_23661);
or UO_2184 (O_2184,N_24150,N_23906);
xor UO_2185 (O_2185,N_22206,N_22878);
nor UO_2186 (O_2186,N_22207,N_24349);
nand UO_2187 (O_2187,N_20093,N_22425);
or UO_2188 (O_2188,N_20876,N_24258);
xor UO_2189 (O_2189,N_24675,N_21606);
xor UO_2190 (O_2190,N_21163,N_21779);
and UO_2191 (O_2191,N_23414,N_20025);
nand UO_2192 (O_2192,N_21135,N_23752);
nand UO_2193 (O_2193,N_20436,N_22678);
nor UO_2194 (O_2194,N_23911,N_21841);
and UO_2195 (O_2195,N_22506,N_23370);
xor UO_2196 (O_2196,N_21970,N_22234);
and UO_2197 (O_2197,N_24800,N_20995);
xor UO_2198 (O_2198,N_24866,N_20090);
and UO_2199 (O_2199,N_20471,N_23705);
xnor UO_2200 (O_2200,N_23748,N_24108);
or UO_2201 (O_2201,N_24739,N_24088);
or UO_2202 (O_2202,N_22787,N_20752);
xnor UO_2203 (O_2203,N_20478,N_23584);
or UO_2204 (O_2204,N_20405,N_23861);
xnor UO_2205 (O_2205,N_24819,N_20717);
xor UO_2206 (O_2206,N_24770,N_23508);
nor UO_2207 (O_2207,N_23048,N_21263);
or UO_2208 (O_2208,N_24900,N_22786);
and UO_2209 (O_2209,N_22749,N_22024);
nand UO_2210 (O_2210,N_23897,N_21086);
and UO_2211 (O_2211,N_20384,N_22157);
nor UO_2212 (O_2212,N_20175,N_23110);
nor UO_2213 (O_2213,N_21340,N_21223);
and UO_2214 (O_2214,N_21127,N_21738);
nand UO_2215 (O_2215,N_22585,N_21194);
xnor UO_2216 (O_2216,N_24583,N_21405);
nor UO_2217 (O_2217,N_24849,N_21420);
xor UO_2218 (O_2218,N_23159,N_20825);
or UO_2219 (O_2219,N_22028,N_22680);
nand UO_2220 (O_2220,N_20524,N_24078);
or UO_2221 (O_2221,N_21013,N_20528);
or UO_2222 (O_2222,N_20462,N_23793);
and UO_2223 (O_2223,N_20928,N_20650);
or UO_2224 (O_2224,N_22356,N_22260);
nor UO_2225 (O_2225,N_24636,N_24220);
xnor UO_2226 (O_2226,N_20716,N_22571);
and UO_2227 (O_2227,N_21541,N_23096);
nand UO_2228 (O_2228,N_22672,N_20875);
or UO_2229 (O_2229,N_23568,N_24865);
nor UO_2230 (O_2230,N_22619,N_21184);
or UO_2231 (O_2231,N_24210,N_24912);
nor UO_2232 (O_2232,N_21908,N_20810);
nor UO_2233 (O_2233,N_20769,N_21197);
or UO_2234 (O_2234,N_22837,N_23888);
nand UO_2235 (O_2235,N_22673,N_21643);
and UO_2236 (O_2236,N_24592,N_23453);
or UO_2237 (O_2237,N_21996,N_21900);
nor UO_2238 (O_2238,N_23737,N_23549);
or UO_2239 (O_2239,N_21020,N_22071);
or UO_2240 (O_2240,N_24655,N_22239);
nor UO_2241 (O_2241,N_20991,N_22450);
nor UO_2242 (O_2242,N_23902,N_20620);
xor UO_2243 (O_2243,N_21780,N_20274);
and UO_2244 (O_2244,N_22412,N_24234);
nor UO_2245 (O_2245,N_20753,N_21840);
and UO_2246 (O_2246,N_22328,N_24810);
nor UO_2247 (O_2247,N_22763,N_24128);
nor UO_2248 (O_2248,N_21373,N_24895);
or UO_2249 (O_2249,N_20670,N_24626);
nor UO_2250 (O_2250,N_22978,N_20930);
nand UO_2251 (O_2251,N_21006,N_23415);
or UO_2252 (O_2252,N_21417,N_21192);
xnor UO_2253 (O_2253,N_23269,N_24270);
nor UO_2254 (O_2254,N_21075,N_20794);
xnor UO_2255 (O_2255,N_20300,N_21094);
or UO_2256 (O_2256,N_22109,N_22890);
nand UO_2257 (O_2257,N_22907,N_22862);
nand UO_2258 (O_2258,N_24775,N_23059);
nor UO_2259 (O_2259,N_22943,N_23829);
nand UO_2260 (O_2260,N_24836,N_24181);
or UO_2261 (O_2261,N_24896,N_20372);
and UO_2262 (O_2262,N_20936,N_24392);
nor UO_2263 (O_2263,N_21388,N_22484);
nand UO_2264 (O_2264,N_21915,N_21898);
or UO_2265 (O_2265,N_22533,N_23550);
or UO_2266 (O_2266,N_20244,N_20614);
nor UO_2267 (O_2267,N_20786,N_23564);
nand UO_2268 (O_2268,N_23730,N_21404);
and UO_2269 (O_2269,N_24245,N_24746);
xnor UO_2270 (O_2270,N_23320,N_20238);
nor UO_2271 (O_2271,N_24009,N_23013);
xor UO_2272 (O_2272,N_21092,N_21538);
and UO_2273 (O_2273,N_22324,N_24250);
or UO_2274 (O_2274,N_22156,N_24855);
and UO_2275 (O_2275,N_22893,N_24863);
nand UO_2276 (O_2276,N_20621,N_24453);
and UO_2277 (O_2277,N_21137,N_20903);
and UO_2278 (O_2278,N_20427,N_20742);
and UO_2279 (O_2279,N_24325,N_21377);
and UO_2280 (O_2280,N_20120,N_22722);
xnor UO_2281 (O_2281,N_21788,N_21854);
or UO_2282 (O_2282,N_24165,N_24647);
xnor UO_2283 (O_2283,N_21776,N_22021);
and UO_2284 (O_2284,N_22273,N_21608);
xnor UO_2285 (O_2285,N_21790,N_21347);
xnor UO_2286 (O_2286,N_22910,N_23015);
or UO_2287 (O_2287,N_23229,N_22836);
and UO_2288 (O_2288,N_20857,N_22521);
nand UO_2289 (O_2289,N_23790,N_22166);
nor UO_2290 (O_2290,N_20615,N_20678);
and UO_2291 (O_2291,N_21613,N_23434);
xor UO_2292 (O_2292,N_20891,N_23927);
xor UO_2293 (O_2293,N_21395,N_23231);
and UO_2294 (O_2294,N_22432,N_22608);
nor UO_2295 (O_2295,N_22891,N_20461);
nand UO_2296 (O_2296,N_23393,N_20993);
or UO_2297 (O_2297,N_21977,N_20334);
xor UO_2298 (O_2298,N_20909,N_23294);
nand UO_2299 (O_2299,N_23359,N_22681);
or UO_2300 (O_2300,N_20052,N_21356);
nor UO_2301 (O_2301,N_23962,N_22785);
xnor UO_2302 (O_2302,N_23383,N_24709);
or UO_2303 (O_2303,N_20477,N_20359);
and UO_2304 (O_2304,N_21646,N_22769);
nand UO_2305 (O_2305,N_21174,N_24560);
and UO_2306 (O_2306,N_20921,N_23179);
or UO_2307 (O_2307,N_21836,N_21487);
nor UO_2308 (O_2308,N_21667,N_21072);
xnor UO_2309 (O_2309,N_20221,N_21742);
or UO_2310 (O_2310,N_20309,N_24832);
xor UO_2311 (O_2311,N_20774,N_20850);
and UO_2312 (O_2312,N_22131,N_20213);
or UO_2313 (O_2313,N_21685,N_22348);
or UO_2314 (O_2314,N_24728,N_22446);
or UO_2315 (O_2315,N_20679,N_22991);
xor UO_2316 (O_2316,N_21680,N_22799);
and UO_2317 (O_2317,N_22656,N_20844);
or UO_2318 (O_2318,N_21523,N_20085);
xnor UO_2319 (O_2319,N_24778,N_22296);
nor UO_2320 (O_2320,N_20641,N_22929);
nand UO_2321 (O_2321,N_23357,N_22056);
or UO_2322 (O_2322,N_21653,N_22794);
nor UO_2323 (O_2323,N_23144,N_20890);
xor UO_2324 (O_2324,N_24769,N_24974);
and UO_2325 (O_2325,N_20078,N_22901);
nand UO_2326 (O_2326,N_23444,N_20010);
nor UO_2327 (O_2327,N_24201,N_22477);
xor UO_2328 (O_2328,N_21471,N_24071);
nor UO_2329 (O_2329,N_23923,N_24901);
or UO_2330 (O_2330,N_24670,N_23256);
or UO_2331 (O_2331,N_20132,N_22473);
xnor UO_2332 (O_2332,N_21712,N_22384);
nor UO_2333 (O_2333,N_20293,N_22379);
nand UO_2334 (O_2334,N_24776,N_21100);
nor UO_2335 (O_2335,N_20604,N_20924);
nand UO_2336 (O_2336,N_21445,N_20744);
and UO_2337 (O_2337,N_22249,N_24734);
and UO_2338 (O_2338,N_21576,N_24822);
and UO_2339 (O_2339,N_21451,N_24466);
nor UO_2340 (O_2340,N_21649,N_21122);
and UO_2341 (O_2341,N_23403,N_24561);
nor UO_2342 (O_2342,N_22509,N_22015);
nand UO_2343 (O_2343,N_24799,N_22005);
xor UO_2344 (O_2344,N_22083,N_21229);
or UO_2345 (O_2345,N_23947,N_21390);
xnor UO_2346 (O_2346,N_20111,N_24398);
nand UO_2347 (O_2347,N_22490,N_24604);
xor UO_2348 (O_2348,N_20098,N_21323);
nand UO_2349 (O_2349,N_21806,N_24574);
nor UO_2350 (O_2350,N_21503,N_20863);
or UO_2351 (O_2351,N_24491,N_21525);
or UO_2352 (O_2352,N_22573,N_21434);
nand UO_2353 (O_2353,N_23054,N_24098);
or UO_2354 (O_2354,N_24614,N_24740);
nor UO_2355 (O_2355,N_21414,N_23881);
nand UO_2356 (O_2356,N_22072,N_24568);
nor UO_2357 (O_2357,N_21446,N_20248);
and UO_2358 (O_2358,N_21268,N_20947);
or UO_2359 (O_2359,N_21540,N_24522);
xnor UO_2360 (O_2360,N_24028,N_23412);
and UO_2361 (O_2361,N_20953,N_21621);
and UO_2362 (O_2362,N_22931,N_20777);
nor UO_2363 (O_2363,N_20795,N_22586);
nand UO_2364 (O_2364,N_23700,N_23938);
nor UO_2365 (O_2365,N_20680,N_23253);
nor UO_2366 (O_2366,N_23337,N_20685);
or UO_2367 (O_2367,N_23607,N_21901);
or UO_2368 (O_2368,N_21665,N_21766);
or UO_2369 (O_2369,N_22036,N_24039);
nand UO_2370 (O_2370,N_23490,N_22556);
xor UO_2371 (O_2371,N_22818,N_23630);
nor UO_2372 (O_2372,N_23451,N_22125);
or UO_2373 (O_2373,N_23682,N_20706);
nand UO_2374 (O_2374,N_23275,N_22266);
or UO_2375 (O_2375,N_20126,N_23079);
nand UO_2376 (O_2376,N_21933,N_20202);
and UO_2377 (O_2377,N_20847,N_20103);
nor UO_2378 (O_2378,N_21971,N_20323);
xnor UO_2379 (O_2379,N_21021,N_23354);
and UO_2380 (O_2380,N_20464,N_24975);
and UO_2381 (O_2381,N_22278,N_20412);
and UO_2382 (O_2382,N_23085,N_22824);
nor UO_2383 (O_2383,N_23764,N_20004);
and UO_2384 (O_2384,N_22179,N_21258);
and UO_2385 (O_2385,N_22654,N_23365);
and UO_2386 (O_2386,N_23217,N_20984);
nand UO_2387 (O_2387,N_21280,N_23060);
xor UO_2388 (O_2388,N_23125,N_24145);
or UO_2389 (O_2389,N_24133,N_20357);
nor UO_2390 (O_2390,N_20326,N_21661);
or UO_2391 (O_2391,N_24486,N_22845);
or UO_2392 (O_2392,N_24660,N_23486);
nor UO_2393 (O_2393,N_20623,N_22121);
and UO_2394 (O_2394,N_24794,N_24591);
and UO_2395 (O_2395,N_22390,N_24267);
and UO_2396 (O_2396,N_23694,N_24480);
nand UO_2397 (O_2397,N_24587,N_24050);
and UO_2398 (O_2398,N_24494,N_20669);
nor UO_2399 (O_2399,N_21801,N_20319);
and UO_2400 (O_2400,N_23193,N_20698);
or UO_2401 (O_2401,N_20138,N_20029);
and UO_2402 (O_2402,N_23912,N_22187);
nor UO_2403 (O_2403,N_21324,N_24259);
nand UO_2404 (O_2404,N_21878,N_20684);
xor UO_2405 (O_2405,N_24685,N_22317);
and UO_2406 (O_2406,N_22209,N_23889);
nand UO_2407 (O_2407,N_20583,N_23714);
and UO_2408 (O_2408,N_22564,N_23741);
xor UO_2409 (O_2409,N_23105,N_22558);
nor UO_2410 (O_2410,N_20988,N_24278);
xor UO_2411 (O_2411,N_20907,N_21756);
and UO_2412 (O_2412,N_21316,N_23240);
xor UO_2413 (O_2413,N_23477,N_21814);
nand UO_2414 (O_2414,N_21083,N_20122);
xor UO_2415 (O_2415,N_23228,N_21360);
xnor UO_2416 (O_2416,N_20940,N_23690);
xnor UO_2417 (O_2417,N_21514,N_21758);
nand UO_2418 (O_2418,N_23542,N_24136);
xnor UO_2419 (O_2419,N_24199,N_21867);
or UO_2420 (O_2420,N_23702,N_22129);
nor UO_2421 (O_2421,N_23086,N_20313);
nand UO_2422 (O_2422,N_21822,N_21103);
and UO_2423 (O_2423,N_23464,N_20151);
nor UO_2424 (O_2424,N_20329,N_23335);
or UO_2425 (O_2425,N_22090,N_23485);
nand UO_2426 (O_2426,N_22489,N_21570);
or UO_2427 (O_2427,N_24057,N_23192);
or UO_2428 (O_2428,N_21123,N_22946);
or UO_2429 (O_2429,N_22440,N_21493);
nand UO_2430 (O_2430,N_22817,N_23725);
nand UO_2431 (O_2431,N_22264,N_23920);
or UO_2432 (O_2432,N_22428,N_20894);
xor UO_2433 (O_2433,N_24504,N_20011);
nor UO_2434 (O_2434,N_20252,N_23822);
nor UO_2435 (O_2435,N_21065,N_20566);
xor UO_2436 (O_2436,N_21798,N_23596);
nand UO_2437 (O_2437,N_20186,N_22281);
or UO_2438 (O_2438,N_23440,N_24790);
xor UO_2439 (O_2439,N_22282,N_24694);
and UO_2440 (O_2440,N_21725,N_23377);
nand UO_2441 (O_2441,N_21511,N_20766);
nor UO_2442 (O_2442,N_21844,N_20557);
and UO_2443 (O_2443,N_23280,N_20170);
or UO_2444 (O_2444,N_21207,N_23922);
or UO_2445 (O_2445,N_24605,N_22712);
nand UO_2446 (O_2446,N_21132,N_24093);
xor UO_2447 (O_2447,N_20674,N_21101);
nor UO_2448 (O_2448,N_24903,N_23321);
xnor UO_2449 (O_2449,N_23203,N_21529);
nand UO_2450 (O_2450,N_23557,N_21833);
or UO_2451 (O_2451,N_23991,N_24006);
xnor UO_2452 (O_2452,N_22830,N_20882);
and UO_2453 (O_2453,N_24545,N_24610);
nor UO_2454 (O_2454,N_20401,N_20260);
xnor UO_2455 (O_2455,N_24899,N_23038);
nor UO_2456 (O_2456,N_22655,N_24367);
xor UO_2457 (O_2457,N_23259,N_21034);
xor UO_2458 (O_2458,N_22706,N_23537);
nor UO_2459 (O_2459,N_24988,N_22309);
and UO_2460 (O_2460,N_20043,N_24265);
xor UO_2461 (O_2461,N_24624,N_21810);
or UO_2462 (O_2462,N_22284,N_22137);
nand UO_2463 (O_2463,N_24686,N_22579);
xor UO_2464 (O_2464,N_20044,N_24657);
nor UO_2465 (O_2465,N_24045,N_24931);
and UO_2466 (O_2466,N_21626,N_20041);
and UO_2467 (O_2467,N_22389,N_24069);
xor UO_2468 (O_2468,N_21793,N_20297);
or UO_2469 (O_2469,N_21550,N_20385);
or UO_2470 (O_2470,N_24862,N_20880);
xnor UO_2471 (O_2471,N_23134,N_20914);
and UO_2472 (O_2472,N_20647,N_24754);
or UO_2473 (O_2473,N_23413,N_20591);
nand UO_2474 (O_2474,N_22001,N_24869);
nand UO_2475 (O_2475,N_24756,N_22498);
xor UO_2476 (O_2476,N_23305,N_24981);
nor UO_2477 (O_2477,N_24736,N_21863);
nand UO_2478 (O_2478,N_21150,N_21748);
nand UO_2479 (O_2479,N_22612,N_23222);
nor UO_2480 (O_2480,N_22305,N_22451);
nor UO_2481 (O_2481,N_23981,N_21896);
nand UO_2482 (O_2482,N_24462,N_23098);
nand UO_2483 (O_2483,N_22920,N_23678);
or UO_2484 (O_2484,N_23300,N_24022);
or UO_2485 (O_2485,N_24066,N_20703);
nor UO_2486 (O_2486,N_24222,N_20828);
or UO_2487 (O_2487,N_22158,N_20860);
nand UO_2488 (O_2488,N_22162,N_23138);
and UO_2489 (O_2489,N_21567,N_22424);
or UO_2490 (O_2490,N_24221,N_20431);
and UO_2491 (O_2491,N_22545,N_23849);
or UO_2492 (O_2492,N_21256,N_21805);
and UO_2493 (O_2493,N_21366,N_24042);
xnor UO_2494 (O_2494,N_22149,N_21004);
and UO_2495 (O_2495,N_23576,N_22373);
xnor UO_2496 (O_2496,N_24406,N_20184);
xnor UO_2497 (O_2497,N_21619,N_22648);
nor UO_2498 (O_2498,N_21010,N_24077);
or UO_2499 (O_2499,N_20584,N_20973);
xor UO_2500 (O_2500,N_21196,N_21423);
or UO_2501 (O_2501,N_20248,N_20225);
nand UO_2502 (O_2502,N_23060,N_20628);
and UO_2503 (O_2503,N_23321,N_20959);
nor UO_2504 (O_2504,N_24435,N_20142);
nand UO_2505 (O_2505,N_20921,N_22149);
or UO_2506 (O_2506,N_22171,N_21455);
nor UO_2507 (O_2507,N_23736,N_24278);
or UO_2508 (O_2508,N_22040,N_22886);
nor UO_2509 (O_2509,N_21650,N_23957);
xor UO_2510 (O_2510,N_24980,N_20580);
or UO_2511 (O_2511,N_20940,N_21360);
xor UO_2512 (O_2512,N_22796,N_22681);
nor UO_2513 (O_2513,N_23075,N_20127);
xnor UO_2514 (O_2514,N_21630,N_23769);
nor UO_2515 (O_2515,N_23571,N_20526);
nor UO_2516 (O_2516,N_23911,N_23999);
xor UO_2517 (O_2517,N_24819,N_22192);
or UO_2518 (O_2518,N_24466,N_20134);
nand UO_2519 (O_2519,N_20574,N_20957);
and UO_2520 (O_2520,N_24174,N_22698);
xnor UO_2521 (O_2521,N_22920,N_24032);
nor UO_2522 (O_2522,N_21549,N_23021);
nand UO_2523 (O_2523,N_22675,N_20391);
nor UO_2524 (O_2524,N_23984,N_22731);
xor UO_2525 (O_2525,N_22543,N_20864);
nand UO_2526 (O_2526,N_21094,N_20771);
xor UO_2527 (O_2527,N_20923,N_20969);
or UO_2528 (O_2528,N_24597,N_20463);
and UO_2529 (O_2529,N_22610,N_20459);
and UO_2530 (O_2530,N_22758,N_21635);
nor UO_2531 (O_2531,N_23376,N_21831);
and UO_2532 (O_2532,N_20091,N_23884);
nand UO_2533 (O_2533,N_24341,N_22938);
nor UO_2534 (O_2534,N_21237,N_22733);
and UO_2535 (O_2535,N_24679,N_21918);
xnor UO_2536 (O_2536,N_20084,N_21916);
or UO_2537 (O_2537,N_20245,N_21231);
nand UO_2538 (O_2538,N_22143,N_21206);
nor UO_2539 (O_2539,N_23957,N_22936);
nor UO_2540 (O_2540,N_20955,N_24298);
xnor UO_2541 (O_2541,N_23900,N_23516);
nor UO_2542 (O_2542,N_21396,N_24668);
xor UO_2543 (O_2543,N_22175,N_23573);
or UO_2544 (O_2544,N_21485,N_23204);
nand UO_2545 (O_2545,N_21045,N_24339);
and UO_2546 (O_2546,N_24924,N_21857);
and UO_2547 (O_2547,N_22785,N_21383);
and UO_2548 (O_2548,N_20008,N_20606);
and UO_2549 (O_2549,N_24931,N_21905);
xor UO_2550 (O_2550,N_21883,N_20244);
or UO_2551 (O_2551,N_22383,N_24874);
nor UO_2552 (O_2552,N_24397,N_23647);
and UO_2553 (O_2553,N_20408,N_23896);
nor UO_2554 (O_2554,N_20002,N_24589);
and UO_2555 (O_2555,N_23174,N_22036);
or UO_2556 (O_2556,N_20471,N_20418);
xnor UO_2557 (O_2557,N_21741,N_24905);
nor UO_2558 (O_2558,N_24962,N_20338);
or UO_2559 (O_2559,N_20999,N_21424);
xnor UO_2560 (O_2560,N_23576,N_24634);
nor UO_2561 (O_2561,N_21306,N_24757);
nor UO_2562 (O_2562,N_23960,N_22432);
and UO_2563 (O_2563,N_22567,N_22197);
and UO_2564 (O_2564,N_22995,N_21066);
nor UO_2565 (O_2565,N_24044,N_20013);
and UO_2566 (O_2566,N_23488,N_24710);
or UO_2567 (O_2567,N_24200,N_21641);
xor UO_2568 (O_2568,N_22534,N_24741);
and UO_2569 (O_2569,N_20899,N_24937);
nand UO_2570 (O_2570,N_22065,N_24743);
nor UO_2571 (O_2571,N_22284,N_23621);
xor UO_2572 (O_2572,N_22571,N_22954);
and UO_2573 (O_2573,N_20635,N_22014);
xnor UO_2574 (O_2574,N_20406,N_24359);
or UO_2575 (O_2575,N_20741,N_22408);
nand UO_2576 (O_2576,N_23585,N_23984);
or UO_2577 (O_2577,N_24535,N_24693);
or UO_2578 (O_2578,N_22596,N_24677);
and UO_2579 (O_2579,N_23467,N_24122);
nand UO_2580 (O_2580,N_24250,N_23844);
nand UO_2581 (O_2581,N_21226,N_22972);
and UO_2582 (O_2582,N_21925,N_21643);
nand UO_2583 (O_2583,N_22213,N_22459);
and UO_2584 (O_2584,N_21506,N_21741);
xnor UO_2585 (O_2585,N_22147,N_20560);
xnor UO_2586 (O_2586,N_20311,N_22044);
nand UO_2587 (O_2587,N_23913,N_21598);
and UO_2588 (O_2588,N_24057,N_21486);
nand UO_2589 (O_2589,N_24619,N_23372);
xnor UO_2590 (O_2590,N_20727,N_23383);
xnor UO_2591 (O_2591,N_20429,N_22955);
nor UO_2592 (O_2592,N_24638,N_21026);
xor UO_2593 (O_2593,N_24564,N_21217);
and UO_2594 (O_2594,N_23537,N_23733);
or UO_2595 (O_2595,N_20793,N_24532);
and UO_2596 (O_2596,N_23081,N_22436);
nor UO_2597 (O_2597,N_20316,N_22105);
nand UO_2598 (O_2598,N_21470,N_20400);
or UO_2599 (O_2599,N_21152,N_21268);
nand UO_2600 (O_2600,N_23444,N_20917);
or UO_2601 (O_2601,N_22803,N_20335);
nand UO_2602 (O_2602,N_24712,N_21384);
nor UO_2603 (O_2603,N_21690,N_24601);
or UO_2604 (O_2604,N_22000,N_24344);
nand UO_2605 (O_2605,N_20149,N_23263);
nand UO_2606 (O_2606,N_21456,N_22044);
nand UO_2607 (O_2607,N_23579,N_22083);
nand UO_2608 (O_2608,N_24378,N_20779);
nand UO_2609 (O_2609,N_20292,N_20055);
nand UO_2610 (O_2610,N_24771,N_21454);
nand UO_2611 (O_2611,N_21842,N_24600);
or UO_2612 (O_2612,N_20103,N_24112);
or UO_2613 (O_2613,N_20821,N_20960);
and UO_2614 (O_2614,N_22405,N_22137);
and UO_2615 (O_2615,N_21186,N_21702);
xor UO_2616 (O_2616,N_21314,N_21867);
and UO_2617 (O_2617,N_23581,N_21971);
or UO_2618 (O_2618,N_21840,N_22590);
and UO_2619 (O_2619,N_22814,N_21518);
and UO_2620 (O_2620,N_20767,N_21549);
nor UO_2621 (O_2621,N_20829,N_22262);
nand UO_2622 (O_2622,N_20883,N_24858);
nor UO_2623 (O_2623,N_22602,N_23017);
or UO_2624 (O_2624,N_23732,N_21674);
nor UO_2625 (O_2625,N_22725,N_23846);
or UO_2626 (O_2626,N_23243,N_22401);
or UO_2627 (O_2627,N_23447,N_24592);
nor UO_2628 (O_2628,N_22725,N_20649);
nor UO_2629 (O_2629,N_21059,N_24015);
and UO_2630 (O_2630,N_22215,N_23629);
xnor UO_2631 (O_2631,N_21385,N_21231);
nor UO_2632 (O_2632,N_23834,N_23334);
and UO_2633 (O_2633,N_20307,N_21610);
nor UO_2634 (O_2634,N_24485,N_22689);
xnor UO_2635 (O_2635,N_21853,N_23585);
or UO_2636 (O_2636,N_22723,N_24278);
xnor UO_2637 (O_2637,N_24886,N_23703);
xor UO_2638 (O_2638,N_23899,N_23064);
nor UO_2639 (O_2639,N_20865,N_20747);
nand UO_2640 (O_2640,N_22609,N_20959);
xnor UO_2641 (O_2641,N_21640,N_21961);
nor UO_2642 (O_2642,N_20254,N_22628);
nor UO_2643 (O_2643,N_24689,N_22595);
nor UO_2644 (O_2644,N_20577,N_24860);
nor UO_2645 (O_2645,N_22908,N_23267);
nand UO_2646 (O_2646,N_21051,N_20307);
nand UO_2647 (O_2647,N_21815,N_24699);
nand UO_2648 (O_2648,N_24368,N_24053);
xor UO_2649 (O_2649,N_21781,N_20002);
xnor UO_2650 (O_2650,N_23778,N_22150);
nand UO_2651 (O_2651,N_21341,N_23881);
xor UO_2652 (O_2652,N_24558,N_21997);
xor UO_2653 (O_2653,N_24001,N_23659);
nor UO_2654 (O_2654,N_24079,N_20451);
nor UO_2655 (O_2655,N_22541,N_20206);
nor UO_2656 (O_2656,N_23581,N_21973);
or UO_2657 (O_2657,N_22716,N_20693);
nor UO_2658 (O_2658,N_20186,N_20125);
and UO_2659 (O_2659,N_24116,N_23432);
nor UO_2660 (O_2660,N_24477,N_21689);
xnor UO_2661 (O_2661,N_22786,N_24288);
xor UO_2662 (O_2662,N_22141,N_20513);
or UO_2663 (O_2663,N_21646,N_23038);
or UO_2664 (O_2664,N_24498,N_21046);
nand UO_2665 (O_2665,N_21161,N_20776);
xnor UO_2666 (O_2666,N_23111,N_24083);
nand UO_2667 (O_2667,N_21026,N_22760);
nor UO_2668 (O_2668,N_20597,N_21072);
nor UO_2669 (O_2669,N_21573,N_20993);
or UO_2670 (O_2670,N_24169,N_20371);
nand UO_2671 (O_2671,N_21203,N_23078);
xnor UO_2672 (O_2672,N_24431,N_21088);
and UO_2673 (O_2673,N_24769,N_20417);
and UO_2674 (O_2674,N_23285,N_24131);
or UO_2675 (O_2675,N_24475,N_24744);
xor UO_2676 (O_2676,N_23597,N_23464);
and UO_2677 (O_2677,N_23418,N_22326);
nand UO_2678 (O_2678,N_20913,N_20125);
xnor UO_2679 (O_2679,N_21727,N_21291);
xnor UO_2680 (O_2680,N_22656,N_24969);
or UO_2681 (O_2681,N_23926,N_20901);
xnor UO_2682 (O_2682,N_21688,N_22706);
nor UO_2683 (O_2683,N_23271,N_21519);
nand UO_2684 (O_2684,N_24112,N_22204);
nor UO_2685 (O_2685,N_24252,N_23336);
and UO_2686 (O_2686,N_21224,N_23463);
nor UO_2687 (O_2687,N_24314,N_22618);
or UO_2688 (O_2688,N_22207,N_24782);
and UO_2689 (O_2689,N_23815,N_23986);
nand UO_2690 (O_2690,N_21795,N_23380);
and UO_2691 (O_2691,N_24300,N_22831);
and UO_2692 (O_2692,N_24815,N_21184);
and UO_2693 (O_2693,N_20185,N_21396);
nor UO_2694 (O_2694,N_20147,N_24478);
xor UO_2695 (O_2695,N_21429,N_20065);
or UO_2696 (O_2696,N_20150,N_20032);
or UO_2697 (O_2697,N_22282,N_24907);
and UO_2698 (O_2698,N_20521,N_23423);
or UO_2699 (O_2699,N_23331,N_20742);
and UO_2700 (O_2700,N_24495,N_24282);
xor UO_2701 (O_2701,N_22226,N_24442);
or UO_2702 (O_2702,N_23312,N_22230);
nor UO_2703 (O_2703,N_21089,N_22619);
or UO_2704 (O_2704,N_21762,N_21248);
and UO_2705 (O_2705,N_21809,N_21875);
nor UO_2706 (O_2706,N_23778,N_24169);
and UO_2707 (O_2707,N_21013,N_24084);
nor UO_2708 (O_2708,N_20245,N_22375);
and UO_2709 (O_2709,N_24797,N_24337);
xor UO_2710 (O_2710,N_24952,N_24681);
and UO_2711 (O_2711,N_23814,N_23122);
or UO_2712 (O_2712,N_24930,N_20717);
nor UO_2713 (O_2713,N_20993,N_21781);
nor UO_2714 (O_2714,N_21840,N_23860);
nor UO_2715 (O_2715,N_24868,N_22547);
nand UO_2716 (O_2716,N_24196,N_24623);
or UO_2717 (O_2717,N_24023,N_24075);
and UO_2718 (O_2718,N_20755,N_20058);
xnor UO_2719 (O_2719,N_20766,N_23039);
nor UO_2720 (O_2720,N_20700,N_24997);
nor UO_2721 (O_2721,N_23253,N_21645);
nor UO_2722 (O_2722,N_20548,N_24404);
xnor UO_2723 (O_2723,N_21099,N_24221);
or UO_2724 (O_2724,N_23739,N_23484);
xnor UO_2725 (O_2725,N_20849,N_24286);
nand UO_2726 (O_2726,N_24059,N_20624);
xnor UO_2727 (O_2727,N_22052,N_22610);
nand UO_2728 (O_2728,N_23625,N_22726);
and UO_2729 (O_2729,N_22904,N_22877);
or UO_2730 (O_2730,N_22744,N_22244);
and UO_2731 (O_2731,N_24753,N_21872);
xor UO_2732 (O_2732,N_22913,N_20000);
and UO_2733 (O_2733,N_20834,N_22951);
nor UO_2734 (O_2734,N_20665,N_22414);
or UO_2735 (O_2735,N_23703,N_20423);
nor UO_2736 (O_2736,N_20913,N_21744);
nor UO_2737 (O_2737,N_21933,N_22516);
nor UO_2738 (O_2738,N_20797,N_21501);
xnor UO_2739 (O_2739,N_21071,N_23450);
and UO_2740 (O_2740,N_20024,N_21042);
and UO_2741 (O_2741,N_24815,N_23256);
xor UO_2742 (O_2742,N_23462,N_20880);
nand UO_2743 (O_2743,N_24162,N_21561);
or UO_2744 (O_2744,N_21873,N_23515);
nor UO_2745 (O_2745,N_23759,N_24591);
xnor UO_2746 (O_2746,N_23718,N_23848);
or UO_2747 (O_2747,N_21079,N_24848);
xor UO_2748 (O_2748,N_23423,N_24578);
and UO_2749 (O_2749,N_22717,N_23175);
xnor UO_2750 (O_2750,N_20714,N_20688);
and UO_2751 (O_2751,N_21144,N_21084);
nand UO_2752 (O_2752,N_21908,N_20121);
xor UO_2753 (O_2753,N_23368,N_22231);
xnor UO_2754 (O_2754,N_24197,N_20527);
nor UO_2755 (O_2755,N_22373,N_20576);
xnor UO_2756 (O_2756,N_20255,N_24854);
nor UO_2757 (O_2757,N_23277,N_21678);
nor UO_2758 (O_2758,N_20068,N_23936);
and UO_2759 (O_2759,N_24194,N_21218);
and UO_2760 (O_2760,N_24545,N_20331);
nor UO_2761 (O_2761,N_24496,N_23558);
or UO_2762 (O_2762,N_20387,N_23901);
or UO_2763 (O_2763,N_22694,N_23994);
and UO_2764 (O_2764,N_20436,N_22169);
and UO_2765 (O_2765,N_24698,N_23749);
nor UO_2766 (O_2766,N_22334,N_21119);
xnor UO_2767 (O_2767,N_20042,N_20160);
xnor UO_2768 (O_2768,N_23653,N_20767);
and UO_2769 (O_2769,N_23568,N_21862);
xnor UO_2770 (O_2770,N_20147,N_22337);
nor UO_2771 (O_2771,N_23119,N_23026);
nand UO_2772 (O_2772,N_24590,N_23008);
or UO_2773 (O_2773,N_21606,N_20919);
and UO_2774 (O_2774,N_24782,N_21401);
nor UO_2775 (O_2775,N_24490,N_21590);
or UO_2776 (O_2776,N_24701,N_21689);
nor UO_2777 (O_2777,N_20097,N_24874);
and UO_2778 (O_2778,N_24575,N_21731);
or UO_2779 (O_2779,N_22583,N_22591);
nand UO_2780 (O_2780,N_21740,N_22512);
nor UO_2781 (O_2781,N_23685,N_21942);
xnor UO_2782 (O_2782,N_22444,N_23648);
nand UO_2783 (O_2783,N_21009,N_20534);
nand UO_2784 (O_2784,N_20982,N_21545);
nor UO_2785 (O_2785,N_21503,N_23475);
and UO_2786 (O_2786,N_23741,N_24977);
nor UO_2787 (O_2787,N_22684,N_21757);
or UO_2788 (O_2788,N_22251,N_22274);
nor UO_2789 (O_2789,N_22639,N_24078);
nand UO_2790 (O_2790,N_23878,N_22044);
xnor UO_2791 (O_2791,N_24962,N_21764);
xnor UO_2792 (O_2792,N_22795,N_20020);
and UO_2793 (O_2793,N_22631,N_20686);
xor UO_2794 (O_2794,N_23710,N_24496);
and UO_2795 (O_2795,N_21314,N_23129);
nand UO_2796 (O_2796,N_20573,N_21825);
and UO_2797 (O_2797,N_21286,N_21079);
and UO_2798 (O_2798,N_23510,N_24879);
xor UO_2799 (O_2799,N_23511,N_24172);
and UO_2800 (O_2800,N_24146,N_23917);
nor UO_2801 (O_2801,N_20828,N_23079);
nor UO_2802 (O_2802,N_20072,N_24918);
xnor UO_2803 (O_2803,N_20456,N_24665);
and UO_2804 (O_2804,N_24924,N_22206);
or UO_2805 (O_2805,N_21173,N_24322);
nand UO_2806 (O_2806,N_21773,N_24827);
nor UO_2807 (O_2807,N_22806,N_23662);
nand UO_2808 (O_2808,N_24110,N_21528);
nor UO_2809 (O_2809,N_20492,N_20026);
and UO_2810 (O_2810,N_21295,N_22399);
nand UO_2811 (O_2811,N_24248,N_24028);
and UO_2812 (O_2812,N_23510,N_20573);
and UO_2813 (O_2813,N_23555,N_22447);
and UO_2814 (O_2814,N_20615,N_20346);
nor UO_2815 (O_2815,N_20178,N_22402);
nand UO_2816 (O_2816,N_22302,N_21923);
or UO_2817 (O_2817,N_21165,N_23790);
nor UO_2818 (O_2818,N_23798,N_20272);
nor UO_2819 (O_2819,N_24419,N_22389);
nand UO_2820 (O_2820,N_24673,N_20654);
xor UO_2821 (O_2821,N_24763,N_24092);
and UO_2822 (O_2822,N_23240,N_22106);
nor UO_2823 (O_2823,N_20328,N_21838);
or UO_2824 (O_2824,N_21112,N_23005);
xnor UO_2825 (O_2825,N_21344,N_23262);
xor UO_2826 (O_2826,N_20704,N_22906);
nand UO_2827 (O_2827,N_20600,N_24328);
and UO_2828 (O_2828,N_20873,N_20454);
and UO_2829 (O_2829,N_21148,N_23651);
nor UO_2830 (O_2830,N_21422,N_22323);
xor UO_2831 (O_2831,N_24757,N_23936);
nand UO_2832 (O_2832,N_23776,N_24735);
nand UO_2833 (O_2833,N_24072,N_24427);
or UO_2834 (O_2834,N_20632,N_21000);
nor UO_2835 (O_2835,N_24991,N_21425);
xor UO_2836 (O_2836,N_21885,N_24447);
nor UO_2837 (O_2837,N_24281,N_24912);
and UO_2838 (O_2838,N_24239,N_22074);
xor UO_2839 (O_2839,N_20599,N_24589);
xnor UO_2840 (O_2840,N_20270,N_20696);
nand UO_2841 (O_2841,N_20777,N_23013);
nor UO_2842 (O_2842,N_20115,N_24153);
xnor UO_2843 (O_2843,N_21799,N_23867);
nor UO_2844 (O_2844,N_22285,N_22365);
nor UO_2845 (O_2845,N_22226,N_23735);
xnor UO_2846 (O_2846,N_23213,N_24198);
xnor UO_2847 (O_2847,N_21320,N_23687);
nor UO_2848 (O_2848,N_20119,N_20573);
xor UO_2849 (O_2849,N_24315,N_24593);
nor UO_2850 (O_2850,N_20787,N_23650);
xnor UO_2851 (O_2851,N_21967,N_20397);
xnor UO_2852 (O_2852,N_24285,N_20881);
xor UO_2853 (O_2853,N_24336,N_23487);
xor UO_2854 (O_2854,N_24581,N_20538);
or UO_2855 (O_2855,N_20389,N_22325);
nand UO_2856 (O_2856,N_22471,N_24608);
nor UO_2857 (O_2857,N_20330,N_24635);
nand UO_2858 (O_2858,N_22026,N_23399);
and UO_2859 (O_2859,N_20146,N_21054);
nand UO_2860 (O_2860,N_23240,N_21287);
xor UO_2861 (O_2861,N_22831,N_20519);
or UO_2862 (O_2862,N_24358,N_20600);
nand UO_2863 (O_2863,N_20873,N_20110);
and UO_2864 (O_2864,N_20074,N_20091);
and UO_2865 (O_2865,N_23809,N_21603);
and UO_2866 (O_2866,N_21517,N_23507);
xnor UO_2867 (O_2867,N_22892,N_22792);
or UO_2868 (O_2868,N_21754,N_24149);
xnor UO_2869 (O_2869,N_22520,N_23205);
xor UO_2870 (O_2870,N_21694,N_20436);
or UO_2871 (O_2871,N_23307,N_20428);
nor UO_2872 (O_2872,N_21966,N_24383);
and UO_2873 (O_2873,N_23029,N_23865);
nor UO_2874 (O_2874,N_23257,N_22584);
or UO_2875 (O_2875,N_22821,N_20665);
nor UO_2876 (O_2876,N_20409,N_23804);
nand UO_2877 (O_2877,N_22346,N_21009);
nand UO_2878 (O_2878,N_24081,N_20474);
xnor UO_2879 (O_2879,N_23615,N_21360);
nand UO_2880 (O_2880,N_24500,N_21887);
xnor UO_2881 (O_2881,N_20257,N_24008);
or UO_2882 (O_2882,N_24879,N_22560);
nor UO_2883 (O_2883,N_23348,N_22561);
xor UO_2884 (O_2884,N_23624,N_24607);
nor UO_2885 (O_2885,N_21943,N_23109);
or UO_2886 (O_2886,N_21740,N_24380);
nor UO_2887 (O_2887,N_20155,N_22874);
and UO_2888 (O_2888,N_24257,N_21032);
and UO_2889 (O_2889,N_22004,N_20159);
and UO_2890 (O_2890,N_22919,N_22336);
xor UO_2891 (O_2891,N_20840,N_23731);
xnor UO_2892 (O_2892,N_20173,N_20705);
xnor UO_2893 (O_2893,N_22774,N_24191);
xor UO_2894 (O_2894,N_24606,N_24344);
and UO_2895 (O_2895,N_21978,N_24271);
or UO_2896 (O_2896,N_24803,N_22639);
nand UO_2897 (O_2897,N_21966,N_22790);
nand UO_2898 (O_2898,N_23028,N_20282);
nand UO_2899 (O_2899,N_20845,N_23330);
xor UO_2900 (O_2900,N_23521,N_23293);
nor UO_2901 (O_2901,N_23322,N_24218);
nor UO_2902 (O_2902,N_20452,N_23060);
nor UO_2903 (O_2903,N_21881,N_22279);
nand UO_2904 (O_2904,N_21688,N_22265);
xor UO_2905 (O_2905,N_20278,N_21171);
xor UO_2906 (O_2906,N_20254,N_23573);
and UO_2907 (O_2907,N_22519,N_22367);
or UO_2908 (O_2908,N_22352,N_24061);
nor UO_2909 (O_2909,N_22724,N_23738);
nor UO_2910 (O_2910,N_21452,N_22119);
or UO_2911 (O_2911,N_20391,N_20952);
xnor UO_2912 (O_2912,N_24563,N_24441);
or UO_2913 (O_2913,N_22797,N_21861);
and UO_2914 (O_2914,N_21534,N_23645);
xnor UO_2915 (O_2915,N_22033,N_21570);
or UO_2916 (O_2916,N_24397,N_20983);
xnor UO_2917 (O_2917,N_20483,N_23363);
xnor UO_2918 (O_2918,N_21710,N_21586);
nor UO_2919 (O_2919,N_23678,N_22331);
or UO_2920 (O_2920,N_21853,N_23463);
and UO_2921 (O_2921,N_23500,N_20461);
nor UO_2922 (O_2922,N_24547,N_20117);
and UO_2923 (O_2923,N_21857,N_23123);
and UO_2924 (O_2924,N_21614,N_23063);
or UO_2925 (O_2925,N_24323,N_20612);
and UO_2926 (O_2926,N_21534,N_22535);
nor UO_2927 (O_2927,N_22667,N_20154);
nand UO_2928 (O_2928,N_20073,N_22920);
nand UO_2929 (O_2929,N_22067,N_21535);
nand UO_2930 (O_2930,N_21101,N_20535);
nor UO_2931 (O_2931,N_24946,N_20306);
nand UO_2932 (O_2932,N_20521,N_21939);
or UO_2933 (O_2933,N_23701,N_23954);
and UO_2934 (O_2934,N_21012,N_20082);
or UO_2935 (O_2935,N_20723,N_20166);
and UO_2936 (O_2936,N_20459,N_20554);
or UO_2937 (O_2937,N_21188,N_24299);
nor UO_2938 (O_2938,N_23283,N_23305);
nand UO_2939 (O_2939,N_24663,N_21275);
nand UO_2940 (O_2940,N_22104,N_23170);
nand UO_2941 (O_2941,N_22148,N_24150);
and UO_2942 (O_2942,N_24297,N_21536);
xnor UO_2943 (O_2943,N_22405,N_21860);
nand UO_2944 (O_2944,N_24994,N_23706);
nand UO_2945 (O_2945,N_21946,N_20464);
or UO_2946 (O_2946,N_21381,N_22460);
nor UO_2947 (O_2947,N_22935,N_23103);
or UO_2948 (O_2948,N_21147,N_22434);
nand UO_2949 (O_2949,N_22097,N_22329);
and UO_2950 (O_2950,N_21666,N_23626);
nand UO_2951 (O_2951,N_21871,N_20310);
xnor UO_2952 (O_2952,N_20424,N_22424);
nand UO_2953 (O_2953,N_20855,N_23337);
nor UO_2954 (O_2954,N_20619,N_22641);
nor UO_2955 (O_2955,N_22727,N_24875);
nor UO_2956 (O_2956,N_20775,N_20086);
nand UO_2957 (O_2957,N_22339,N_23797);
nand UO_2958 (O_2958,N_24844,N_23705);
and UO_2959 (O_2959,N_20061,N_24698);
nor UO_2960 (O_2960,N_20601,N_20093);
and UO_2961 (O_2961,N_21229,N_20064);
or UO_2962 (O_2962,N_21096,N_22070);
xnor UO_2963 (O_2963,N_22970,N_22191);
and UO_2964 (O_2964,N_20147,N_20537);
or UO_2965 (O_2965,N_24877,N_24218);
or UO_2966 (O_2966,N_24600,N_22230);
nand UO_2967 (O_2967,N_24187,N_23208);
xor UO_2968 (O_2968,N_21929,N_23091);
nand UO_2969 (O_2969,N_24656,N_24422);
and UO_2970 (O_2970,N_23167,N_21369);
xnor UO_2971 (O_2971,N_20011,N_22265);
xor UO_2972 (O_2972,N_22236,N_23090);
nor UO_2973 (O_2973,N_20138,N_20586);
nor UO_2974 (O_2974,N_20900,N_20914);
or UO_2975 (O_2975,N_23226,N_23910);
and UO_2976 (O_2976,N_21849,N_20840);
xnor UO_2977 (O_2977,N_23776,N_24175);
or UO_2978 (O_2978,N_21938,N_24738);
and UO_2979 (O_2979,N_23684,N_21190);
or UO_2980 (O_2980,N_24676,N_24135);
nand UO_2981 (O_2981,N_21848,N_24414);
or UO_2982 (O_2982,N_21276,N_21871);
nor UO_2983 (O_2983,N_24509,N_24363);
or UO_2984 (O_2984,N_22706,N_24819);
and UO_2985 (O_2985,N_21472,N_24454);
or UO_2986 (O_2986,N_22864,N_21551);
and UO_2987 (O_2987,N_21728,N_24743);
or UO_2988 (O_2988,N_24022,N_22978);
and UO_2989 (O_2989,N_23690,N_24453);
xnor UO_2990 (O_2990,N_24492,N_21956);
nor UO_2991 (O_2991,N_24493,N_24764);
xnor UO_2992 (O_2992,N_21904,N_20208);
nand UO_2993 (O_2993,N_20826,N_21650);
or UO_2994 (O_2994,N_22373,N_20305);
or UO_2995 (O_2995,N_24855,N_20127);
nand UO_2996 (O_2996,N_20057,N_21025);
nand UO_2997 (O_2997,N_22219,N_20291);
xor UO_2998 (O_2998,N_22271,N_24437);
nor UO_2999 (O_2999,N_24821,N_20425);
endmodule