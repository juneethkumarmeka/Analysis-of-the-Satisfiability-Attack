module basic_750_5000_1000_5_levels_5xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
and U0 (N_0,In_640,In_705);
or U1 (N_1,In_266,In_685);
xnor U2 (N_2,In_115,In_172);
and U3 (N_3,In_26,In_111);
xor U4 (N_4,In_533,In_158);
nand U5 (N_5,In_727,In_149);
and U6 (N_6,In_213,In_692);
and U7 (N_7,In_128,In_617);
nor U8 (N_8,In_670,In_542);
and U9 (N_9,In_463,In_634);
and U10 (N_10,In_50,In_159);
nor U11 (N_11,In_301,In_724);
or U12 (N_12,In_399,In_486);
or U13 (N_13,In_745,In_376);
and U14 (N_14,In_117,In_572);
nor U15 (N_15,In_459,In_269);
or U16 (N_16,In_101,In_56);
or U17 (N_17,In_352,In_652);
or U18 (N_18,In_96,In_252);
and U19 (N_19,In_488,In_249);
nand U20 (N_20,In_503,In_302);
or U21 (N_21,In_458,In_176);
nand U22 (N_22,In_205,In_613);
or U23 (N_23,In_309,In_283);
and U24 (N_24,In_103,In_482);
xnor U25 (N_25,In_448,In_220);
nand U26 (N_26,In_427,In_337);
nand U27 (N_27,In_131,In_61);
nand U28 (N_28,In_528,In_44);
or U29 (N_29,In_304,In_584);
nor U30 (N_30,In_484,In_133);
or U31 (N_31,In_116,In_42);
or U32 (N_32,In_515,In_614);
nor U33 (N_33,In_109,In_168);
nand U34 (N_34,In_255,In_144);
nand U35 (N_35,In_529,In_150);
and U36 (N_36,In_322,In_145);
and U37 (N_37,In_650,In_478);
nand U38 (N_38,In_703,In_135);
nand U39 (N_39,In_643,In_747);
or U40 (N_40,In_59,In_139);
nand U41 (N_41,In_368,In_242);
and U42 (N_42,In_575,In_294);
or U43 (N_43,In_627,In_425);
nor U44 (N_44,In_363,In_430);
nor U45 (N_45,In_718,In_577);
or U46 (N_46,In_21,In_3);
and U47 (N_47,In_34,In_677);
nor U48 (N_48,In_365,In_79);
or U49 (N_49,In_182,In_169);
or U50 (N_50,In_489,In_141);
nor U51 (N_51,In_611,In_244);
nor U52 (N_52,In_393,In_235);
nor U53 (N_53,In_440,In_280);
nand U54 (N_54,In_586,In_497);
nor U55 (N_55,In_237,In_550);
and U56 (N_56,In_271,In_123);
nand U57 (N_57,In_532,In_39);
and U58 (N_58,In_62,In_544);
or U59 (N_59,In_362,In_288);
and U60 (N_60,In_281,In_327);
or U61 (N_61,In_212,In_234);
nor U62 (N_62,In_160,In_349);
or U63 (N_63,In_641,In_218);
nand U64 (N_64,In_635,In_605);
nor U65 (N_65,In_530,In_84);
nor U66 (N_66,In_672,In_462);
or U67 (N_67,In_259,In_667);
and U68 (N_68,In_637,In_574);
or U69 (N_69,In_413,In_582);
nor U70 (N_70,In_130,In_749);
and U71 (N_71,In_183,In_290);
or U72 (N_72,In_28,In_606);
nand U73 (N_73,In_33,In_600);
nand U74 (N_74,In_625,In_329);
or U75 (N_75,In_348,In_711);
and U76 (N_76,In_119,In_70);
and U77 (N_77,In_43,In_706);
and U78 (N_78,In_163,In_728);
or U79 (N_79,In_318,In_320);
and U80 (N_80,In_98,In_653);
nor U81 (N_81,In_668,In_219);
nor U82 (N_82,In_397,In_739);
and U83 (N_83,In_570,In_708);
or U84 (N_84,In_513,In_381);
and U85 (N_85,In_291,In_655);
or U86 (N_86,In_85,In_490);
nor U87 (N_87,In_498,In_125);
and U88 (N_88,In_80,In_569);
and U89 (N_89,In_356,In_394);
nand U90 (N_90,In_373,In_523);
nand U91 (N_91,In_197,In_157);
and U92 (N_92,In_579,In_29);
nand U93 (N_93,In_164,In_618);
nand U94 (N_94,In_541,In_173);
and U95 (N_95,In_270,In_686);
xnor U96 (N_96,In_675,In_60);
and U97 (N_97,In_546,In_260);
and U98 (N_98,In_298,In_94);
xor U99 (N_99,In_4,In_525);
nor U100 (N_100,In_645,In_682);
xor U101 (N_101,In_700,In_562);
and U102 (N_102,In_691,In_69);
nor U103 (N_103,In_622,In_648);
xor U104 (N_104,In_743,In_714);
nand U105 (N_105,In_660,In_306);
nor U106 (N_106,In_537,In_557);
nor U107 (N_107,In_276,In_432);
nor U108 (N_108,In_184,In_419);
nand U109 (N_109,In_639,In_646);
and U110 (N_110,In_684,In_263);
or U111 (N_111,In_375,In_412);
nand U112 (N_112,In_536,In_140);
nor U113 (N_113,In_199,In_704);
or U114 (N_114,In_279,In_722);
xor U115 (N_115,In_75,In_437);
or U116 (N_116,In_253,In_286);
or U117 (N_117,In_312,In_351);
nor U118 (N_118,In_414,In_710);
nor U119 (N_119,In_701,In_204);
or U120 (N_120,In_725,In_509);
and U121 (N_121,In_632,In_734);
nor U122 (N_122,In_284,In_180);
nor U123 (N_123,In_592,In_521);
or U124 (N_124,In_230,In_603);
nand U125 (N_125,In_538,In_468);
nor U126 (N_126,In_347,In_424);
and U127 (N_127,In_407,In_421);
and U128 (N_128,In_656,In_68);
or U129 (N_129,In_494,In_717);
nor U130 (N_130,In_520,In_221);
nor U131 (N_131,In_167,In_387);
nor U132 (N_132,In_341,In_53);
or U133 (N_133,In_18,In_355);
nand U134 (N_134,In_165,In_19);
nand U135 (N_135,In_240,In_372);
nor U136 (N_136,In_662,In_201);
nor U137 (N_137,In_441,In_334);
or U138 (N_138,In_14,In_451);
nand U139 (N_139,In_442,In_594);
nor U140 (N_140,In_607,In_402);
nor U141 (N_141,In_671,In_663);
and U142 (N_142,In_436,In_633);
xor U143 (N_143,In_456,In_154);
or U144 (N_144,In_64,In_738);
and U145 (N_145,In_556,In_181);
and U146 (N_146,In_573,In_619);
xnor U147 (N_147,In_100,In_534);
or U148 (N_148,In_71,In_338);
nand U149 (N_149,In_203,In_207);
or U150 (N_150,In_114,In_483);
nand U151 (N_151,In_24,In_6);
or U152 (N_152,In_251,In_171);
xnor U153 (N_153,In_247,In_364);
and U154 (N_154,In_262,In_323);
and U155 (N_155,In_77,In_2);
and U156 (N_156,In_104,In_517);
and U157 (N_157,In_12,In_241);
xnor U158 (N_158,In_258,In_609);
xnor U159 (N_159,In_325,In_620);
and U160 (N_160,In_514,In_696);
or U161 (N_161,In_687,In_535);
nand U162 (N_162,In_357,In_206);
and U163 (N_163,In_106,In_426);
nand U164 (N_164,In_403,In_423);
nor U165 (N_165,In_31,In_93);
and U166 (N_166,In_474,In_649);
and U167 (N_167,In_510,In_518);
nor U168 (N_168,In_272,In_545);
xnor U169 (N_169,In_688,In_118);
and U170 (N_170,In_449,In_254);
or U171 (N_171,In_112,In_628);
and U172 (N_172,In_335,In_231);
nand U173 (N_173,In_499,In_464);
nand U174 (N_174,In_110,In_328);
nand U175 (N_175,In_720,In_505);
nor U176 (N_176,In_248,In_527);
or U177 (N_177,In_475,In_549);
nand U178 (N_178,In_99,In_319);
nor U179 (N_179,In_553,In_744);
or U180 (N_180,In_560,In_429);
nor U181 (N_181,In_457,In_23);
or U182 (N_182,In_377,In_593);
or U183 (N_183,In_175,In_694);
nand U184 (N_184,In_651,In_623);
or U185 (N_185,In_137,In_602);
or U186 (N_186,In_32,In_41);
nor U187 (N_187,In_400,In_52);
or U188 (N_188,In_243,In_564);
nand U189 (N_189,In_539,In_673);
nand U190 (N_190,In_127,In_88);
xnor U191 (N_191,In_443,In_126);
nor U192 (N_192,In_721,In_477);
or U193 (N_193,In_748,In_732);
or U194 (N_194,In_404,In_78);
xor U195 (N_195,In_487,In_178);
and U196 (N_196,In_416,In_9);
and U197 (N_197,In_151,In_601);
or U198 (N_198,In_152,In_36);
and U199 (N_199,In_588,In_480);
and U200 (N_200,In_519,In_608);
nor U201 (N_201,In_370,In_66);
nor U202 (N_202,In_245,In_492);
and U203 (N_203,In_46,In_47);
nor U204 (N_204,In_174,In_626);
and U205 (N_205,In_709,In_208);
and U206 (N_206,In_354,In_386);
and U207 (N_207,In_679,In_733);
and U208 (N_208,In_310,In_631);
or U209 (N_209,In_689,In_166);
nor U210 (N_210,In_82,In_707);
nand U211 (N_211,In_589,In_344);
or U212 (N_212,In_214,In_124);
or U213 (N_213,In_502,In_305);
nand U214 (N_214,In_339,In_297);
nand U215 (N_215,In_472,In_345);
nand U216 (N_216,In_54,In_49);
nor U217 (N_217,In_236,In_554);
xor U218 (N_218,In_445,In_95);
nor U219 (N_219,In_469,In_378);
or U220 (N_220,In_681,In_332);
nand U221 (N_221,In_223,In_224);
xnor U222 (N_222,In_561,In_741);
or U223 (N_223,In_20,In_274);
nand U224 (N_224,In_142,In_1);
nor U225 (N_225,In_389,In_367);
xor U226 (N_226,In_664,In_303);
nand U227 (N_227,In_239,In_699);
nor U228 (N_228,In_285,In_737);
or U229 (N_229,In_516,In_57);
or U230 (N_230,In_196,In_470);
and U231 (N_231,In_282,In_374);
and U232 (N_232,In_313,In_693);
xor U233 (N_233,In_132,In_384);
nand U234 (N_234,In_250,In_216);
or U235 (N_235,In_390,In_379);
or U236 (N_236,In_485,In_16);
nor U237 (N_237,In_256,In_610);
and U238 (N_238,In_669,In_598);
or U239 (N_239,In_7,In_86);
and U240 (N_240,In_540,In_493);
nand U241 (N_241,In_277,In_331);
or U242 (N_242,In_177,In_15);
or U243 (N_243,In_630,In_326);
or U244 (N_244,In_315,In_278);
nand U245 (N_245,In_559,In_229);
xnor U246 (N_246,In_359,In_555);
nand U247 (N_247,In_83,In_558);
xor U248 (N_248,In_543,In_300);
or U249 (N_249,In_261,In_292);
and U250 (N_250,In_496,In_73);
nor U251 (N_251,In_500,In_287);
and U252 (N_252,In_683,In_435);
or U253 (N_253,In_217,In_148);
and U254 (N_254,In_697,In_120);
nand U255 (N_255,In_391,In_37);
nor U256 (N_256,In_11,In_420);
or U257 (N_257,In_188,In_385);
or U258 (N_258,In_170,In_481);
or U259 (N_259,In_654,In_647);
nand U260 (N_260,In_597,In_674);
nor U261 (N_261,In_371,In_580);
and U262 (N_262,In_105,In_415);
xnor U263 (N_263,In_552,In_460);
nand U264 (N_264,In_726,In_526);
xnor U265 (N_265,In_330,In_202);
nand U266 (N_266,In_129,In_658);
nor U267 (N_267,In_495,In_578);
nand U268 (N_268,In_369,In_522);
or U269 (N_269,In_702,In_102);
nor U270 (N_270,In_38,In_401);
nand U271 (N_271,In_388,In_74);
xnor U272 (N_272,In_343,In_590);
xnor U273 (N_273,In_512,In_246);
nor U274 (N_274,In_746,In_179);
nor U275 (N_275,In_336,In_690);
and U276 (N_276,In_48,In_146);
and U277 (N_277,In_438,In_595);
nor U278 (N_278,In_307,In_238);
nand U279 (N_279,In_531,In_121);
nand U280 (N_280,In_209,In_72);
or U281 (N_281,In_89,In_191);
or U282 (N_282,In_225,In_455);
and U283 (N_283,In_10,In_551);
or U284 (N_284,In_629,In_715);
nand U285 (N_285,In_638,In_511);
and U286 (N_286,In_678,In_90);
xnor U287 (N_287,In_65,In_289);
nand U288 (N_288,In_422,In_273);
nor U289 (N_289,In_107,In_507);
and U290 (N_290,In_113,In_275);
nor U291 (N_291,In_616,In_565);
nor U292 (N_292,In_713,In_396);
nand U293 (N_293,In_333,In_358);
nor U294 (N_294,In_342,In_405);
nor U295 (N_295,In_433,In_680);
or U296 (N_296,In_471,In_740);
nand U297 (N_297,In_308,In_408);
nor U298 (N_298,In_716,In_143);
nor U299 (N_299,In_25,In_317);
xor U300 (N_300,In_742,In_434);
nor U301 (N_301,In_226,In_321);
and U302 (N_302,In_192,In_467);
nand U303 (N_303,In_383,In_504);
nand U304 (N_304,In_644,In_257);
or U305 (N_305,In_439,In_63);
and U306 (N_306,In_35,In_76);
and U307 (N_307,In_566,In_547);
and U308 (N_308,In_228,In_466);
nand U309 (N_309,In_156,In_730);
or U310 (N_310,In_524,In_136);
or U311 (N_311,In_108,In_444);
nand U312 (N_312,In_27,In_162);
or U313 (N_313,In_491,In_581);
xor U314 (N_314,In_731,In_316);
or U315 (N_315,In_479,In_185);
and U316 (N_316,In_729,In_265);
nand U317 (N_317,In_659,In_361);
or U318 (N_318,In_642,In_615);
and U319 (N_319,In_55,In_91);
nor U320 (N_320,In_189,In_293);
and U321 (N_321,In_501,In_360);
xnor U322 (N_322,In_17,In_147);
or U323 (N_323,In_211,In_473);
and U324 (N_324,In_450,In_698);
and U325 (N_325,In_134,In_13);
or U326 (N_326,In_621,In_596);
and U327 (N_327,In_51,In_398);
nor U328 (N_328,In_392,In_81);
xor U329 (N_329,In_657,In_719);
and U330 (N_330,In_431,In_187);
nor U331 (N_331,In_299,In_567);
nand U332 (N_332,In_661,In_380);
and U333 (N_333,In_194,In_604);
or U334 (N_334,In_665,In_453);
nand U335 (N_335,In_264,In_447);
xnor U336 (N_336,In_311,In_410);
or U337 (N_337,In_314,In_233);
xor U338 (N_338,In_200,In_382);
nand U339 (N_339,In_22,In_30);
nor U340 (N_340,In_350,In_723);
or U341 (N_341,In_40,In_712);
nand U342 (N_342,In_295,In_346);
or U343 (N_343,In_296,In_161);
nand U344 (N_344,In_232,In_428);
nand U345 (N_345,In_97,In_406);
nor U346 (N_346,In_268,In_736);
and U347 (N_347,In_576,In_193);
and U348 (N_348,In_67,In_548);
and U349 (N_349,In_636,In_409);
and U350 (N_350,In_92,In_465);
or U351 (N_351,In_195,In_676);
and U352 (N_352,In_571,In_324);
nand U353 (N_353,In_222,In_0);
and U354 (N_354,In_417,In_461);
and U355 (N_355,In_366,In_267);
and U356 (N_356,In_190,In_563);
and U357 (N_357,In_568,In_735);
xnor U358 (N_358,In_138,In_210);
and U359 (N_359,In_612,In_45);
nor U360 (N_360,In_227,In_476);
nand U361 (N_361,In_624,In_215);
nand U362 (N_362,In_340,In_5);
nand U363 (N_363,In_353,In_87);
or U364 (N_364,In_198,In_153);
xor U365 (N_365,In_446,In_411);
nand U366 (N_366,In_395,In_666);
or U367 (N_367,In_591,In_186);
nand U368 (N_368,In_583,In_155);
and U369 (N_369,In_452,In_454);
or U370 (N_370,In_508,In_58);
nor U371 (N_371,In_506,In_585);
or U372 (N_372,In_122,In_418);
xnor U373 (N_373,In_599,In_587);
and U374 (N_374,In_8,In_695);
nand U375 (N_375,In_544,In_25);
and U376 (N_376,In_342,In_341);
or U377 (N_377,In_27,In_464);
or U378 (N_378,In_359,In_544);
nor U379 (N_379,In_257,In_318);
or U380 (N_380,In_576,In_627);
xnor U381 (N_381,In_379,In_519);
nand U382 (N_382,In_614,In_190);
nor U383 (N_383,In_590,In_362);
and U384 (N_384,In_398,In_505);
nor U385 (N_385,In_484,In_273);
nor U386 (N_386,In_255,In_446);
and U387 (N_387,In_713,In_653);
nand U388 (N_388,In_125,In_617);
nor U389 (N_389,In_187,In_695);
and U390 (N_390,In_198,In_670);
and U391 (N_391,In_165,In_566);
and U392 (N_392,In_345,In_330);
nor U393 (N_393,In_237,In_430);
and U394 (N_394,In_337,In_261);
nor U395 (N_395,In_479,In_191);
nor U396 (N_396,In_654,In_193);
and U397 (N_397,In_239,In_60);
and U398 (N_398,In_34,In_506);
and U399 (N_399,In_366,In_363);
nand U400 (N_400,In_186,In_413);
and U401 (N_401,In_385,In_374);
nand U402 (N_402,In_449,In_468);
xor U403 (N_403,In_205,In_359);
nor U404 (N_404,In_485,In_221);
or U405 (N_405,In_162,In_454);
xnor U406 (N_406,In_631,In_72);
nand U407 (N_407,In_460,In_141);
nand U408 (N_408,In_209,In_210);
nand U409 (N_409,In_316,In_30);
nand U410 (N_410,In_582,In_79);
or U411 (N_411,In_41,In_363);
or U412 (N_412,In_143,In_58);
nor U413 (N_413,In_448,In_42);
nor U414 (N_414,In_585,In_508);
and U415 (N_415,In_166,In_343);
and U416 (N_416,In_737,In_174);
nand U417 (N_417,In_344,In_194);
and U418 (N_418,In_96,In_121);
nand U419 (N_419,In_235,In_279);
xnor U420 (N_420,In_365,In_731);
or U421 (N_421,In_580,In_50);
nand U422 (N_422,In_197,In_247);
nor U423 (N_423,In_585,In_279);
nor U424 (N_424,In_662,In_457);
xor U425 (N_425,In_666,In_571);
or U426 (N_426,In_274,In_102);
or U427 (N_427,In_485,In_412);
nor U428 (N_428,In_379,In_647);
and U429 (N_429,In_152,In_77);
and U430 (N_430,In_415,In_570);
or U431 (N_431,In_526,In_530);
nand U432 (N_432,In_535,In_366);
and U433 (N_433,In_315,In_77);
nor U434 (N_434,In_595,In_107);
nand U435 (N_435,In_305,In_457);
and U436 (N_436,In_438,In_659);
nor U437 (N_437,In_317,In_507);
nand U438 (N_438,In_190,In_192);
nor U439 (N_439,In_215,In_512);
and U440 (N_440,In_622,In_681);
or U441 (N_441,In_25,In_413);
nand U442 (N_442,In_96,In_721);
nor U443 (N_443,In_284,In_346);
or U444 (N_444,In_649,In_648);
or U445 (N_445,In_185,In_187);
nor U446 (N_446,In_286,In_186);
nor U447 (N_447,In_119,In_49);
nand U448 (N_448,In_80,In_77);
nand U449 (N_449,In_637,In_288);
or U450 (N_450,In_601,In_687);
or U451 (N_451,In_523,In_563);
and U452 (N_452,In_309,In_7);
and U453 (N_453,In_23,In_392);
xor U454 (N_454,In_556,In_464);
nand U455 (N_455,In_391,In_581);
and U456 (N_456,In_443,In_571);
nor U457 (N_457,In_553,In_587);
and U458 (N_458,In_387,In_103);
or U459 (N_459,In_167,In_318);
or U460 (N_460,In_343,In_390);
and U461 (N_461,In_718,In_405);
and U462 (N_462,In_691,In_493);
and U463 (N_463,In_94,In_41);
xnor U464 (N_464,In_551,In_542);
nor U465 (N_465,In_567,In_113);
nor U466 (N_466,In_227,In_269);
nand U467 (N_467,In_37,In_610);
xor U468 (N_468,In_461,In_626);
nor U469 (N_469,In_287,In_624);
nand U470 (N_470,In_351,In_739);
xnor U471 (N_471,In_468,In_742);
nand U472 (N_472,In_471,In_414);
xor U473 (N_473,In_541,In_487);
xnor U474 (N_474,In_99,In_439);
nor U475 (N_475,In_642,In_260);
or U476 (N_476,In_200,In_122);
xnor U477 (N_477,In_671,In_507);
nand U478 (N_478,In_699,In_300);
nor U479 (N_479,In_284,In_701);
or U480 (N_480,In_509,In_690);
nor U481 (N_481,In_379,In_9);
nor U482 (N_482,In_472,In_524);
or U483 (N_483,In_649,In_607);
xnor U484 (N_484,In_467,In_699);
nor U485 (N_485,In_152,In_671);
nand U486 (N_486,In_366,In_709);
nor U487 (N_487,In_622,In_28);
and U488 (N_488,In_226,In_62);
xnor U489 (N_489,In_595,In_670);
or U490 (N_490,In_596,In_372);
nor U491 (N_491,In_527,In_0);
or U492 (N_492,In_183,In_374);
xnor U493 (N_493,In_706,In_287);
and U494 (N_494,In_600,In_529);
nor U495 (N_495,In_33,In_391);
nor U496 (N_496,In_704,In_660);
nor U497 (N_497,In_131,In_604);
and U498 (N_498,In_239,In_680);
or U499 (N_499,In_531,In_509);
nand U500 (N_500,In_631,In_491);
nand U501 (N_501,In_746,In_507);
nor U502 (N_502,In_641,In_667);
and U503 (N_503,In_350,In_745);
nor U504 (N_504,In_653,In_411);
or U505 (N_505,In_152,In_408);
xnor U506 (N_506,In_142,In_128);
nand U507 (N_507,In_509,In_395);
and U508 (N_508,In_623,In_360);
nor U509 (N_509,In_436,In_188);
and U510 (N_510,In_261,In_696);
and U511 (N_511,In_373,In_6);
or U512 (N_512,In_348,In_319);
nand U513 (N_513,In_101,In_221);
and U514 (N_514,In_124,In_554);
xor U515 (N_515,In_441,In_276);
or U516 (N_516,In_732,In_144);
or U517 (N_517,In_83,In_233);
nand U518 (N_518,In_357,In_232);
nor U519 (N_519,In_427,In_17);
or U520 (N_520,In_225,In_267);
nand U521 (N_521,In_183,In_628);
nor U522 (N_522,In_374,In_191);
or U523 (N_523,In_416,In_549);
or U524 (N_524,In_100,In_652);
nand U525 (N_525,In_380,In_489);
or U526 (N_526,In_608,In_679);
xor U527 (N_527,In_220,In_489);
and U528 (N_528,In_631,In_217);
xnor U529 (N_529,In_498,In_317);
and U530 (N_530,In_619,In_34);
nand U531 (N_531,In_230,In_540);
xnor U532 (N_532,In_16,In_325);
and U533 (N_533,In_745,In_241);
nand U534 (N_534,In_124,In_631);
nand U535 (N_535,In_587,In_54);
nor U536 (N_536,In_88,In_556);
nor U537 (N_537,In_582,In_446);
nor U538 (N_538,In_235,In_154);
nor U539 (N_539,In_481,In_596);
nand U540 (N_540,In_668,In_615);
xor U541 (N_541,In_607,In_413);
nand U542 (N_542,In_129,In_177);
and U543 (N_543,In_55,In_292);
nor U544 (N_544,In_161,In_348);
or U545 (N_545,In_272,In_526);
and U546 (N_546,In_296,In_25);
or U547 (N_547,In_511,In_691);
nand U548 (N_548,In_281,In_560);
nor U549 (N_549,In_279,In_520);
or U550 (N_550,In_575,In_572);
nor U551 (N_551,In_171,In_132);
nor U552 (N_552,In_665,In_57);
or U553 (N_553,In_463,In_163);
nor U554 (N_554,In_526,In_259);
and U555 (N_555,In_67,In_571);
or U556 (N_556,In_734,In_468);
and U557 (N_557,In_269,In_23);
xnor U558 (N_558,In_432,In_660);
nor U559 (N_559,In_76,In_142);
nand U560 (N_560,In_651,In_183);
or U561 (N_561,In_262,In_474);
nor U562 (N_562,In_516,In_513);
nand U563 (N_563,In_435,In_448);
nor U564 (N_564,In_366,In_400);
nand U565 (N_565,In_536,In_199);
or U566 (N_566,In_458,In_114);
or U567 (N_567,In_58,In_265);
nand U568 (N_568,In_621,In_28);
or U569 (N_569,In_655,In_266);
nand U570 (N_570,In_405,In_63);
xnor U571 (N_571,In_679,In_656);
nor U572 (N_572,In_559,In_191);
nand U573 (N_573,In_401,In_420);
nor U574 (N_574,In_339,In_491);
and U575 (N_575,In_296,In_279);
and U576 (N_576,In_607,In_313);
or U577 (N_577,In_481,In_403);
nand U578 (N_578,In_545,In_91);
or U579 (N_579,In_533,In_468);
or U580 (N_580,In_630,In_112);
nor U581 (N_581,In_624,In_728);
nor U582 (N_582,In_190,In_251);
or U583 (N_583,In_537,In_726);
xor U584 (N_584,In_472,In_98);
xnor U585 (N_585,In_212,In_452);
nand U586 (N_586,In_439,In_437);
or U587 (N_587,In_533,In_721);
nand U588 (N_588,In_152,In_56);
xor U589 (N_589,In_598,In_594);
or U590 (N_590,In_100,In_143);
nor U591 (N_591,In_106,In_444);
and U592 (N_592,In_376,In_445);
and U593 (N_593,In_199,In_617);
nand U594 (N_594,In_104,In_214);
nor U595 (N_595,In_399,In_384);
xor U596 (N_596,In_78,In_261);
xnor U597 (N_597,In_700,In_148);
and U598 (N_598,In_502,In_13);
and U599 (N_599,In_601,In_749);
nand U600 (N_600,In_499,In_50);
nor U601 (N_601,In_448,In_449);
and U602 (N_602,In_130,In_414);
and U603 (N_603,In_226,In_6);
or U604 (N_604,In_656,In_156);
nand U605 (N_605,In_297,In_535);
nor U606 (N_606,In_534,In_202);
xor U607 (N_607,In_268,In_357);
nand U608 (N_608,In_290,In_143);
or U609 (N_609,In_702,In_611);
nor U610 (N_610,In_672,In_483);
xnor U611 (N_611,In_209,In_625);
or U612 (N_612,In_401,In_281);
or U613 (N_613,In_442,In_573);
and U614 (N_614,In_681,In_390);
or U615 (N_615,In_392,In_524);
or U616 (N_616,In_581,In_483);
nor U617 (N_617,In_488,In_330);
nor U618 (N_618,In_84,In_125);
or U619 (N_619,In_325,In_388);
nand U620 (N_620,In_593,In_68);
nand U621 (N_621,In_464,In_680);
and U622 (N_622,In_583,In_31);
nand U623 (N_623,In_243,In_540);
or U624 (N_624,In_621,In_98);
nand U625 (N_625,In_570,In_618);
nor U626 (N_626,In_635,In_269);
and U627 (N_627,In_674,In_642);
nor U628 (N_628,In_679,In_695);
or U629 (N_629,In_561,In_468);
or U630 (N_630,In_353,In_688);
and U631 (N_631,In_729,In_642);
xnor U632 (N_632,In_204,In_117);
or U633 (N_633,In_496,In_248);
nand U634 (N_634,In_713,In_59);
and U635 (N_635,In_742,In_498);
or U636 (N_636,In_714,In_310);
nor U637 (N_637,In_540,In_473);
nor U638 (N_638,In_42,In_93);
nand U639 (N_639,In_86,In_132);
or U640 (N_640,In_201,In_175);
or U641 (N_641,In_93,In_692);
xnor U642 (N_642,In_368,In_464);
or U643 (N_643,In_302,In_332);
and U644 (N_644,In_393,In_608);
nand U645 (N_645,In_210,In_691);
xor U646 (N_646,In_378,In_638);
and U647 (N_647,In_566,In_381);
and U648 (N_648,In_261,In_73);
or U649 (N_649,In_493,In_566);
nand U650 (N_650,In_268,In_476);
and U651 (N_651,In_680,In_721);
and U652 (N_652,In_280,In_257);
nand U653 (N_653,In_408,In_261);
nor U654 (N_654,In_463,In_520);
or U655 (N_655,In_103,In_442);
nand U656 (N_656,In_538,In_158);
nand U657 (N_657,In_227,In_40);
or U658 (N_658,In_569,In_645);
or U659 (N_659,In_734,In_159);
nand U660 (N_660,In_418,In_731);
nor U661 (N_661,In_6,In_543);
nand U662 (N_662,In_296,In_107);
and U663 (N_663,In_312,In_359);
nand U664 (N_664,In_39,In_385);
and U665 (N_665,In_532,In_689);
nor U666 (N_666,In_625,In_265);
nor U667 (N_667,In_656,In_508);
nor U668 (N_668,In_663,In_444);
or U669 (N_669,In_302,In_498);
nand U670 (N_670,In_621,In_242);
nand U671 (N_671,In_673,In_262);
or U672 (N_672,In_426,In_29);
or U673 (N_673,In_286,In_211);
xnor U674 (N_674,In_29,In_184);
and U675 (N_675,In_399,In_521);
nand U676 (N_676,In_386,In_307);
nand U677 (N_677,In_1,In_542);
nand U678 (N_678,In_445,In_142);
and U679 (N_679,In_195,In_567);
nand U680 (N_680,In_36,In_181);
nand U681 (N_681,In_456,In_537);
nor U682 (N_682,In_207,In_697);
or U683 (N_683,In_658,In_448);
nor U684 (N_684,In_599,In_569);
and U685 (N_685,In_459,In_399);
nand U686 (N_686,In_639,In_144);
xor U687 (N_687,In_68,In_346);
or U688 (N_688,In_68,In_295);
nor U689 (N_689,In_734,In_5);
nand U690 (N_690,In_185,In_545);
and U691 (N_691,In_612,In_738);
nand U692 (N_692,In_736,In_287);
and U693 (N_693,In_250,In_54);
nor U694 (N_694,In_744,In_479);
or U695 (N_695,In_559,In_747);
nor U696 (N_696,In_356,In_194);
xnor U697 (N_697,In_507,In_302);
or U698 (N_698,In_412,In_635);
or U699 (N_699,In_406,In_331);
nand U700 (N_700,In_6,In_577);
xnor U701 (N_701,In_743,In_280);
nor U702 (N_702,In_463,In_443);
and U703 (N_703,In_580,In_71);
nand U704 (N_704,In_99,In_290);
or U705 (N_705,In_507,In_735);
and U706 (N_706,In_186,In_196);
nand U707 (N_707,In_515,In_746);
or U708 (N_708,In_617,In_185);
nand U709 (N_709,In_32,In_415);
and U710 (N_710,In_713,In_69);
or U711 (N_711,In_346,In_333);
xnor U712 (N_712,In_385,In_531);
nand U713 (N_713,In_48,In_648);
nor U714 (N_714,In_662,In_193);
and U715 (N_715,In_155,In_231);
and U716 (N_716,In_343,In_723);
or U717 (N_717,In_458,In_419);
nand U718 (N_718,In_595,In_307);
nand U719 (N_719,In_511,In_58);
nand U720 (N_720,In_720,In_651);
nand U721 (N_721,In_610,In_293);
nor U722 (N_722,In_322,In_366);
and U723 (N_723,In_374,In_413);
nor U724 (N_724,In_146,In_340);
nand U725 (N_725,In_677,In_705);
or U726 (N_726,In_11,In_109);
and U727 (N_727,In_227,In_211);
or U728 (N_728,In_279,In_350);
nor U729 (N_729,In_490,In_146);
and U730 (N_730,In_467,In_301);
nand U731 (N_731,In_404,In_545);
nor U732 (N_732,In_66,In_299);
and U733 (N_733,In_479,In_699);
nand U734 (N_734,In_497,In_594);
nand U735 (N_735,In_493,In_364);
and U736 (N_736,In_103,In_733);
and U737 (N_737,In_529,In_584);
nor U738 (N_738,In_121,In_412);
nand U739 (N_739,In_465,In_182);
nand U740 (N_740,In_359,In_558);
or U741 (N_741,In_2,In_739);
nand U742 (N_742,In_519,In_18);
nor U743 (N_743,In_505,In_55);
nand U744 (N_744,In_11,In_65);
and U745 (N_745,In_226,In_302);
nand U746 (N_746,In_140,In_653);
nor U747 (N_747,In_354,In_281);
nand U748 (N_748,In_259,In_550);
nor U749 (N_749,In_495,In_389);
nand U750 (N_750,In_213,In_639);
or U751 (N_751,In_22,In_488);
or U752 (N_752,In_136,In_68);
or U753 (N_753,In_91,In_231);
nand U754 (N_754,In_255,In_312);
nand U755 (N_755,In_601,In_111);
and U756 (N_756,In_284,In_716);
or U757 (N_757,In_63,In_707);
or U758 (N_758,In_351,In_435);
or U759 (N_759,In_565,In_469);
or U760 (N_760,In_189,In_331);
nor U761 (N_761,In_427,In_288);
and U762 (N_762,In_176,In_674);
xnor U763 (N_763,In_34,In_325);
xnor U764 (N_764,In_174,In_310);
nor U765 (N_765,In_69,In_280);
nand U766 (N_766,In_469,In_343);
nor U767 (N_767,In_693,In_660);
nor U768 (N_768,In_308,In_42);
and U769 (N_769,In_497,In_386);
nor U770 (N_770,In_286,In_613);
or U771 (N_771,In_555,In_579);
or U772 (N_772,In_504,In_541);
nor U773 (N_773,In_347,In_309);
nand U774 (N_774,In_98,In_226);
or U775 (N_775,In_145,In_469);
xnor U776 (N_776,In_525,In_15);
and U777 (N_777,In_232,In_26);
and U778 (N_778,In_507,In_44);
nor U779 (N_779,In_546,In_530);
nand U780 (N_780,In_372,In_77);
nand U781 (N_781,In_66,In_372);
or U782 (N_782,In_17,In_246);
and U783 (N_783,In_676,In_607);
and U784 (N_784,In_0,In_714);
nor U785 (N_785,In_25,In_530);
or U786 (N_786,In_394,In_206);
nor U787 (N_787,In_376,In_553);
nand U788 (N_788,In_68,In_312);
nor U789 (N_789,In_23,In_489);
nor U790 (N_790,In_569,In_520);
or U791 (N_791,In_691,In_92);
or U792 (N_792,In_170,In_191);
nand U793 (N_793,In_702,In_529);
xnor U794 (N_794,In_581,In_648);
nor U795 (N_795,In_227,In_477);
or U796 (N_796,In_646,In_297);
and U797 (N_797,In_103,In_186);
xnor U798 (N_798,In_367,In_414);
nor U799 (N_799,In_298,In_537);
nor U800 (N_800,In_516,In_59);
and U801 (N_801,In_103,In_315);
xor U802 (N_802,In_269,In_739);
and U803 (N_803,In_402,In_584);
nand U804 (N_804,In_682,In_129);
and U805 (N_805,In_52,In_36);
or U806 (N_806,In_493,In_71);
and U807 (N_807,In_513,In_62);
xnor U808 (N_808,In_670,In_651);
or U809 (N_809,In_167,In_364);
nor U810 (N_810,In_188,In_137);
or U811 (N_811,In_106,In_744);
xor U812 (N_812,In_569,In_260);
nand U813 (N_813,In_251,In_629);
nor U814 (N_814,In_448,In_612);
nor U815 (N_815,In_732,In_412);
and U816 (N_816,In_641,In_331);
nor U817 (N_817,In_45,In_614);
nor U818 (N_818,In_323,In_65);
xnor U819 (N_819,In_17,In_411);
and U820 (N_820,In_391,In_58);
or U821 (N_821,In_388,In_206);
or U822 (N_822,In_677,In_427);
and U823 (N_823,In_157,In_733);
nor U824 (N_824,In_339,In_175);
nand U825 (N_825,In_562,In_252);
xor U826 (N_826,In_683,In_246);
nand U827 (N_827,In_188,In_362);
and U828 (N_828,In_345,In_145);
and U829 (N_829,In_629,In_681);
nor U830 (N_830,In_573,In_51);
xnor U831 (N_831,In_380,In_529);
nand U832 (N_832,In_281,In_597);
xor U833 (N_833,In_186,In_152);
nor U834 (N_834,In_194,In_300);
or U835 (N_835,In_736,In_155);
and U836 (N_836,In_647,In_261);
and U837 (N_837,In_365,In_641);
nor U838 (N_838,In_674,In_489);
and U839 (N_839,In_748,In_124);
xor U840 (N_840,In_411,In_132);
or U841 (N_841,In_285,In_14);
and U842 (N_842,In_382,In_710);
nor U843 (N_843,In_658,In_49);
or U844 (N_844,In_529,In_690);
and U845 (N_845,In_217,In_716);
and U846 (N_846,In_495,In_169);
or U847 (N_847,In_523,In_457);
or U848 (N_848,In_374,In_220);
or U849 (N_849,In_367,In_410);
nor U850 (N_850,In_375,In_639);
nor U851 (N_851,In_179,In_448);
nand U852 (N_852,In_682,In_391);
nor U853 (N_853,In_16,In_507);
or U854 (N_854,In_542,In_280);
nor U855 (N_855,In_378,In_32);
and U856 (N_856,In_132,In_699);
nand U857 (N_857,In_9,In_283);
xor U858 (N_858,In_416,In_530);
nor U859 (N_859,In_239,In_619);
and U860 (N_860,In_483,In_657);
xor U861 (N_861,In_660,In_134);
and U862 (N_862,In_424,In_50);
nand U863 (N_863,In_571,In_370);
nand U864 (N_864,In_513,In_246);
or U865 (N_865,In_125,In_584);
nand U866 (N_866,In_518,In_181);
or U867 (N_867,In_153,In_641);
and U868 (N_868,In_286,In_714);
and U869 (N_869,In_311,In_276);
nand U870 (N_870,In_333,In_536);
nand U871 (N_871,In_326,In_293);
and U872 (N_872,In_318,In_682);
nand U873 (N_873,In_557,In_361);
or U874 (N_874,In_258,In_275);
or U875 (N_875,In_387,In_652);
or U876 (N_876,In_532,In_211);
or U877 (N_877,In_312,In_200);
or U878 (N_878,In_76,In_139);
and U879 (N_879,In_657,In_191);
xor U880 (N_880,In_443,In_160);
xnor U881 (N_881,In_664,In_222);
nand U882 (N_882,In_317,In_65);
and U883 (N_883,In_324,In_160);
nor U884 (N_884,In_401,In_275);
or U885 (N_885,In_660,In_64);
and U886 (N_886,In_493,In_84);
or U887 (N_887,In_303,In_234);
nand U888 (N_888,In_288,In_544);
nand U889 (N_889,In_637,In_616);
nand U890 (N_890,In_388,In_400);
xnor U891 (N_891,In_506,In_137);
or U892 (N_892,In_120,In_121);
and U893 (N_893,In_428,In_234);
nor U894 (N_894,In_285,In_379);
nor U895 (N_895,In_641,In_597);
nand U896 (N_896,In_138,In_426);
or U897 (N_897,In_740,In_515);
nor U898 (N_898,In_520,In_198);
or U899 (N_899,In_402,In_430);
nor U900 (N_900,In_714,In_538);
nor U901 (N_901,In_658,In_449);
or U902 (N_902,In_655,In_408);
xnor U903 (N_903,In_409,In_437);
and U904 (N_904,In_487,In_197);
nor U905 (N_905,In_375,In_372);
xor U906 (N_906,In_480,In_578);
nand U907 (N_907,In_393,In_610);
xor U908 (N_908,In_6,In_400);
or U909 (N_909,In_680,In_479);
nand U910 (N_910,In_270,In_76);
and U911 (N_911,In_309,In_224);
nor U912 (N_912,In_695,In_258);
and U913 (N_913,In_557,In_543);
nor U914 (N_914,In_47,In_231);
nor U915 (N_915,In_414,In_245);
nor U916 (N_916,In_694,In_314);
or U917 (N_917,In_519,In_482);
nand U918 (N_918,In_588,In_6);
or U919 (N_919,In_229,In_604);
nand U920 (N_920,In_488,In_443);
xnor U921 (N_921,In_614,In_460);
or U922 (N_922,In_295,In_364);
or U923 (N_923,In_693,In_53);
xnor U924 (N_924,In_187,In_538);
and U925 (N_925,In_622,In_272);
nand U926 (N_926,In_570,In_118);
or U927 (N_927,In_380,In_193);
nand U928 (N_928,In_371,In_709);
or U929 (N_929,In_588,In_315);
nor U930 (N_930,In_599,In_365);
or U931 (N_931,In_729,In_375);
nand U932 (N_932,In_293,In_33);
nor U933 (N_933,In_730,In_574);
nand U934 (N_934,In_685,In_26);
or U935 (N_935,In_23,In_243);
nor U936 (N_936,In_513,In_117);
or U937 (N_937,In_355,In_680);
nor U938 (N_938,In_140,In_596);
and U939 (N_939,In_76,In_23);
nand U940 (N_940,In_543,In_649);
nor U941 (N_941,In_448,In_7);
or U942 (N_942,In_642,In_533);
or U943 (N_943,In_631,In_101);
nand U944 (N_944,In_709,In_17);
and U945 (N_945,In_113,In_439);
and U946 (N_946,In_36,In_317);
and U947 (N_947,In_167,In_280);
and U948 (N_948,In_278,In_199);
and U949 (N_949,In_612,In_349);
or U950 (N_950,In_238,In_356);
nor U951 (N_951,In_9,In_222);
nand U952 (N_952,In_218,In_194);
or U953 (N_953,In_530,In_252);
or U954 (N_954,In_62,In_268);
nand U955 (N_955,In_337,In_382);
nand U956 (N_956,In_565,In_276);
nor U957 (N_957,In_168,In_121);
nor U958 (N_958,In_613,In_694);
or U959 (N_959,In_233,In_403);
xnor U960 (N_960,In_293,In_4);
nand U961 (N_961,In_56,In_227);
or U962 (N_962,In_512,In_133);
and U963 (N_963,In_592,In_298);
or U964 (N_964,In_443,In_393);
nor U965 (N_965,In_474,In_379);
nand U966 (N_966,In_578,In_84);
nand U967 (N_967,In_675,In_679);
xor U968 (N_968,In_389,In_454);
nand U969 (N_969,In_295,In_430);
nand U970 (N_970,In_682,In_202);
and U971 (N_971,In_208,In_98);
and U972 (N_972,In_296,In_624);
xor U973 (N_973,In_351,In_205);
or U974 (N_974,In_56,In_459);
and U975 (N_975,In_561,In_531);
xnor U976 (N_976,In_479,In_267);
or U977 (N_977,In_691,In_215);
nand U978 (N_978,In_527,In_343);
nand U979 (N_979,In_721,In_70);
and U980 (N_980,In_393,In_549);
or U981 (N_981,In_388,In_714);
and U982 (N_982,In_396,In_634);
and U983 (N_983,In_500,In_533);
and U984 (N_984,In_173,In_389);
nor U985 (N_985,In_248,In_676);
xor U986 (N_986,In_241,In_701);
and U987 (N_987,In_700,In_617);
or U988 (N_988,In_363,In_635);
nand U989 (N_989,In_371,In_73);
nand U990 (N_990,In_385,In_723);
nand U991 (N_991,In_457,In_744);
and U992 (N_992,In_309,In_747);
or U993 (N_993,In_437,In_80);
nor U994 (N_994,In_454,In_276);
nor U995 (N_995,In_352,In_692);
nor U996 (N_996,In_159,In_68);
xnor U997 (N_997,In_598,In_127);
nor U998 (N_998,In_645,In_533);
nor U999 (N_999,In_200,In_522);
xor U1000 (N_1000,N_930,N_119);
or U1001 (N_1001,N_526,N_534);
nand U1002 (N_1002,N_621,N_520);
xnor U1003 (N_1003,N_272,N_984);
or U1004 (N_1004,N_750,N_519);
nor U1005 (N_1005,N_168,N_501);
or U1006 (N_1006,N_493,N_79);
or U1007 (N_1007,N_347,N_226);
nor U1008 (N_1008,N_951,N_708);
nand U1009 (N_1009,N_6,N_723);
or U1010 (N_1010,N_827,N_140);
nor U1011 (N_1011,N_477,N_434);
nand U1012 (N_1012,N_183,N_5);
or U1013 (N_1013,N_910,N_885);
nor U1014 (N_1014,N_73,N_311);
nor U1015 (N_1015,N_688,N_923);
nand U1016 (N_1016,N_27,N_960);
nand U1017 (N_1017,N_985,N_203);
and U1018 (N_1018,N_178,N_93);
or U1019 (N_1019,N_8,N_383);
and U1020 (N_1020,N_23,N_94);
or U1021 (N_1021,N_128,N_897);
and U1022 (N_1022,N_462,N_142);
nor U1023 (N_1023,N_880,N_587);
and U1024 (N_1024,N_934,N_210);
nor U1025 (N_1025,N_883,N_115);
nand U1026 (N_1026,N_891,N_972);
or U1027 (N_1027,N_716,N_539);
or U1028 (N_1028,N_219,N_954);
nand U1029 (N_1029,N_892,N_581);
and U1030 (N_1030,N_285,N_724);
xor U1031 (N_1031,N_822,N_691);
or U1032 (N_1032,N_152,N_784);
nor U1033 (N_1033,N_692,N_382);
and U1034 (N_1034,N_893,N_753);
or U1035 (N_1035,N_940,N_246);
and U1036 (N_1036,N_276,N_683);
nor U1037 (N_1037,N_282,N_346);
or U1038 (N_1038,N_908,N_700);
nor U1039 (N_1039,N_579,N_807);
nand U1040 (N_1040,N_26,N_350);
or U1041 (N_1041,N_832,N_116);
xnor U1042 (N_1042,N_864,N_681);
nand U1043 (N_1043,N_640,N_686);
and U1044 (N_1044,N_196,N_180);
nor U1045 (N_1045,N_679,N_532);
nor U1046 (N_1046,N_889,N_590);
or U1047 (N_1047,N_484,N_460);
and U1048 (N_1048,N_609,N_999);
nor U1049 (N_1049,N_963,N_281);
nor U1050 (N_1050,N_695,N_956);
nand U1051 (N_1051,N_664,N_2);
nand U1052 (N_1052,N_761,N_172);
nor U1053 (N_1053,N_838,N_231);
and U1054 (N_1054,N_192,N_171);
and U1055 (N_1055,N_336,N_261);
nor U1056 (N_1056,N_903,N_987);
or U1057 (N_1057,N_352,N_239);
nand U1058 (N_1058,N_355,N_890);
or U1059 (N_1059,N_645,N_47);
and U1060 (N_1060,N_986,N_97);
or U1061 (N_1061,N_505,N_585);
and U1062 (N_1062,N_390,N_104);
nor U1063 (N_1063,N_666,N_805);
nor U1064 (N_1064,N_961,N_811);
and U1065 (N_1065,N_517,N_829);
or U1066 (N_1066,N_488,N_220);
and U1067 (N_1067,N_411,N_1);
nand U1068 (N_1068,N_33,N_641);
or U1069 (N_1069,N_300,N_546);
nor U1070 (N_1070,N_973,N_450);
and U1071 (N_1071,N_945,N_810);
and U1072 (N_1072,N_323,N_976);
nand U1073 (N_1073,N_980,N_148);
nor U1074 (N_1074,N_101,N_565);
nor U1075 (N_1075,N_249,N_58);
nand U1076 (N_1076,N_943,N_78);
nand U1077 (N_1077,N_179,N_583);
or U1078 (N_1078,N_314,N_952);
nand U1079 (N_1079,N_310,N_372);
xnor U1080 (N_1080,N_169,N_289);
nand U1081 (N_1081,N_126,N_479);
or U1082 (N_1082,N_60,N_461);
xor U1083 (N_1083,N_469,N_67);
nand U1084 (N_1084,N_35,N_250);
or U1085 (N_1085,N_287,N_674);
nor U1086 (N_1086,N_167,N_768);
nor U1087 (N_1087,N_186,N_302);
xnor U1088 (N_1088,N_354,N_907);
and U1089 (N_1089,N_369,N_510);
nand U1090 (N_1090,N_543,N_50);
and U1091 (N_1091,N_22,N_915);
or U1092 (N_1092,N_599,N_266);
and U1093 (N_1093,N_339,N_165);
nand U1094 (N_1094,N_969,N_662);
or U1095 (N_1095,N_362,N_330);
xor U1096 (N_1096,N_797,N_373);
nand U1097 (N_1097,N_495,N_652);
nand U1098 (N_1098,N_854,N_851);
nand U1099 (N_1099,N_759,N_81);
and U1100 (N_1100,N_793,N_427);
xor U1101 (N_1101,N_690,N_243);
and U1102 (N_1102,N_596,N_638);
nand U1103 (N_1103,N_922,N_533);
nand U1104 (N_1104,N_744,N_563);
or U1105 (N_1105,N_475,N_114);
or U1106 (N_1106,N_845,N_559);
or U1107 (N_1107,N_557,N_191);
nand U1108 (N_1108,N_10,N_40);
or U1109 (N_1109,N_727,N_393);
nor U1110 (N_1110,N_994,N_632);
nor U1111 (N_1111,N_800,N_657);
nand U1112 (N_1112,N_595,N_625);
or U1113 (N_1113,N_408,N_284);
nand U1114 (N_1114,N_886,N_392);
nor U1115 (N_1115,N_228,N_491);
xnor U1116 (N_1116,N_366,N_770);
nor U1117 (N_1117,N_574,N_482);
or U1118 (N_1118,N_506,N_646);
nor U1119 (N_1119,N_843,N_749);
or U1120 (N_1120,N_417,N_555);
and U1121 (N_1121,N_798,N_63);
nand U1122 (N_1122,N_857,N_746);
or U1123 (N_1123,N_547,N_942);
nand U1124 (N_1124,N_62,N_421);
and U1125 (N_1125,N_642,N_364);
nor U1126 (N_1126,N_123,N_270);
nor U1127 (N_1127,N_156,N_415);
nand U1128 (N_1128,N_24,N_861);
nor U1129 (N_1129,N_103,N_978);
nor U1130 (N_1130,N_665,N_267);
nand U1131 (N_1131,N_320,N_789);
nand U1132 (N_1132,N_573,N_705);
nand U1133 (N_1133,N_748,N_321);
nor U1134 (N_1134,N_299,N_874);
or U1135 (N_1135,N_28,N_820);
nor U1136 (N_1136,N_176,N_340);
and U1137 (N_1137,N_66,N_702);
nand U1138 (N_1138,N_855,N_668);
nor U1139 (N_1139,N_896,N_388);
xor U1140 (N_1140,N_254,N_410);
or U1141 (N_1141,N_707,N_131);
nor U1142 (N_1142,N_124,N_521);
and U1143 (N_1143,N_568,N_859);
nand U1144 (N_1144,N_296,N_778);
and U1145 (N_1145,N_513,N_255);
or U1146 (N_1146,N_948,N_358);
or U1147 (N_1147,N_997,N_879);
or U1148 (N_1148,N_55,N_663);
nand U1149 (N_1149,N_380,N_420);
nand U1150 (N_1150,N_912,N_122);
nor U1151 (N_1151,N_836,N_18);
nand U1152 (N_1152,N_260,N_75);
and U1153 (N_1153,N_379,N_538);
nand U1154 (N_1154,N_333,N_537);
nor U1155 (N_1155,N_802,N_847);
and U1156 (N_1156,N_556,N_161);
nor U1157 (N_1157,N_763,N_926);
or U1158 (N_1158,N_4,N_713);
or U1159 (N_1159,N_834,N_483);
xor U1160 (N_1160,N_92,N_85);
and U1161 (N_1161,N_840,N_714);
nand U1162 (N_1162,N_865,N_30);
or U1163 (N_1163,N_251,N_207);
or U1164 (N_1164,N_306,N_637);
nand U1165 (N_1165,N_514,N_89);
or U1166 (N_1166,N_858,N_571);
and U1167 (N_1167,N_230,N_584);
nand U1168 (N_1168,N_525,N_830);
nand U1169 (N_1169,N_801,N_529);
nor U1170 (N_1170,N_639,N_360);
nand U1171 (N_1171,N_283,N_215);
or U1172 (N_1172,N_357,N_919);
and U1173 (N_1173,N_471,N_738);
and U1174 (N_1174,N_435,N_911);
or U1175 (N_1175,N_374,N_395);
nor U1176 (N_1176,N_205,N_653);
nor U1177 (N_1177,N_769,N_606);
nor U1178 (N_1178,N_474,N_955);
nor U1179 (N_1179,N_561,N_132);
nor U1180 (N_1180,N_144,N_37);
and U1181 (N_1181,N_737,N_704);
nor U1182 (N_1182,N_470,N_950);
nor U1183 (N_1183,N_967,N_337);
nand U1184 (N_1184,N_887,N_603);
nor U1185 (N_1185,N_562,N_979);
xor U1186 (N_1186,N_643,N_80);
or U1187 (N_1187,N_504,N_57);
or U1188 (N_1188,N_776,N_201);
and U1189 (N_1189,N_386,N_868);
nor U1190 (N_1190,N_279,N_117);
and U1191 (N_1191,N_947,N_20);
or U1192 (N_1192,N_998,N_96);
or U1193 (N_1193,N_338,N_719);
nand U1194 (N_1194,N_188,N_170);
nor U1195 (N_1195,N_105,N_129);
or U1196 (N_1196,N_906,N_490);
and U1197 (N_1197,N_689,N_895);
nand U1198 (N_1198,N_745,N_835);
or U1199 (N_1199,N_757,N_367);
or U1200 (N_1200,N_342,N_673);
nand U1201 (N_1201,N_863,N_617);
nand U1202 (N_1202,N_751,N_275);
nor U1203 (N_1203,N_946,N_499);
nand U1204 (N_1204,N_884,N_157);
and U1205 (N_1205,N_134,N_401);
or U1206 (N_1206,N_160,N_442);
nor U1207 (N_1207,N_438,N_108);
xnor U1208 (N_1208,N_507,N_990);
nand U1209 (N_1209,N_159,N_644);
nand U1210 (N_1210,N_687,N_198);
nand U1211 (N_1211,N_697,N_619);
and U1212 (N_1212,N_828,N_359);
or U1213 (N_1213,N_43,N_651);
nor U1214 (N_1214,N_925,N_677);
nor U1215 (N_1215,N_576,N_781);
nor U1216 (N_1216,N_698,N_402);
nor U1217 (N_1217,N_549,N_523);
nor U1218 (N_1218,N_436,N_9);
nor U1219 (N_1219,N_739,N_597);
or U1220 (N_1220,N_190,N_38);
or U1221 (N_1221,N_909,N_247);
nand U1222 (N_1222,N_837,N_711);
or U1223 (N_1223,N_459,N_849);
xor U1224 (N_1224,N_658,N_368);
nand U1225 (N_1225,N_416,N_194);
nor U1226 (N_1226,N_286,N_515);
nor U1227 (N_1227,N_842,N_240);
or U1228 (N_1228,N_381,N_7);
and U1229 (N_1229,N_343,N_937);
and U1230 (N_1230,N_914,N_536);
or U1231 (N_1231,N_212,N_407);
xnor U1232 (N_1232,N_815,N_613);
nor U1233 (N_1233,N_446,N_14);
nand U1234 (N_1234,N_487,N_413);
and U1235 (N_1235,N_996,N_158);
xor U1236 (N_1236,N_110,N_699);
nor U1237 (N_1237,N_480,N_548);
xor U1238 (N_1238,N_580,N_552);
nor U1239 (N_1239,N_508,N_701);
or U1240 (N_1240,N_959,N_535);
or U1241 (N_1241,N_42,N_983);
nand U1242 (N_1242,N_61,N_65);
nand U1243 (N_1243,N_545,N_263);
nor U1244 (N_1244,N_905,N_709);
or U1245 (N_1245,N_248,N_932);
or U1246 (N_1246,N_349,N_318);
nor U1247 (N_1247,N_703,N_933);
and U1248 (N_1248,N_472,N_592);
nand U1249 (N_1249,N_747,N_64);
or U1250 (N_1250,N_931,N_752);
or U1251 (N_1251,N_649,N_163);
nand U1252 (N_1252,N_672,N_558);
and U1253 (N_1253,N_422,N_418);
and U1254 (N_1254,N_200,N_109);
nand U1255 (N_1255,N_655,N_83);
nand U1256 (N_1256,N_399,N_551);
or U1257 (N_1257,N_432,N_378);
or U1258 (N_1258,N_760,N_607);
and U1259 (N_1259,N_682,N_317);
or U1260 (N_1260,N_804,N_731);
or U1261 (N_1261,N_852,N_918);
nor U1262 (N_1262,N_305,N_694);
xor U1263 (N_1263,N_439,N_308);
and U1264 (N_1264,N_99,N_229);
nor U1265 (N_1265,N_298,N_426);
and U1266 (N_1266,N_670,N_494);
nor U1267 (N_1267,N_944,N_589);
nor U1268 (N_1268,N_503,N_878);
nand U1269 (N_1269,N_732,N_531);
nor U1270 (N_1270,N_385,N_332);
xnor U1271 (N_1271,N_898,N_796);
or U1272 (N_1272,N_913,N_821);
nor U1273 (N_1273,N_775,N_291);
or U1274 (N_1274,N_629,N_611);
nand U1275 (N_1275,N_71,N_363);
nor U1276 (N_1276,N_684,N_154);
nor U1277 (N_1277,N_628,N_222);
xor U1278 (N_1278,N_41,N_975);
nor U1279 (N_1279,N_869,N_569);
xor U1280 (N_1280,N_130,N_817);
or U1281 (N_1281,N_736,N_257);
nand U1282 (N_1282,N_578,N_319);
and U1283 (N_1283,N_680,N_150);
nand U1284 (N_1284,N_166,N_742);
nand U1285 (N_1285,N_862,N_881);
and U1286 (N_1286,N_202,N_882);
and U1287 (N_1287,N_353,N_957);
or U1288 (N_1288,N_232,N_466);
nor U1289 (N_1289,N_217,N_82);
nor U1290 (N_1290,N_256,N_630);
or U1291 (N_1291,N_106,N_204);
nor U1292 (N_1292,N_455,N_788);
nand U1293 (N_1293,N_740,N_920);
xor U1294 (N_1294,N_871,N_540);
or U1295 (N_1295,N_46,N_722);
and U1296 (N_1296,N_924,N_235);
or U1297 (N_1297,N_783,N_988);
and U1298 (N_1298,N_34,N_492);
and U1299 (N_1299,N_712,N_197);
or U1300 (N_1300,N_502,N_635);
and U1301 (N_1301,N_634,N_767);
or U1302 (N_1302,N_147,N_391);
nor U1303 (N_1303,N_334,N_588);
and U1304 (N_1304,N_322,N_258);
and U1305 (N_1305,N_624,N_98);
or U1306 (N_1306,N_327,N_15);
nor U1307 (N_1307,N_777,N_139);
and U1308 (N_1308,N_211,N_825);
nor U1309 (N_1309,N_91,N_660);
nor U1310 (N_1310,N_345,N_107);
nand U1311 (N_1311,N_530,N_982);
nor U1312 (N_1312,N_771,N_389);
xor U1313 (N_1313,N_452,N_456);
nand U1314 (N_1314,N_177,N_457);
nor U1315 (N_1315,N_717,N_964);
nor U1316 (N_1316,N_958,N_111);
nand U1317 (N_1317,N_610,N_19);
and U1318 (N_1318,N_900,N_473);
nand U1319 (N_1319,N_608,N_780);
nor U1320 (N_1320,N_904,N_468);
xor U1321 (N_1321,N_764,N_453);
nand U1322 (N_1322,N_175,N_928);
nand U1323 (N_1323,N_365,N_794);
and U1324 (N_1324,N_516,N_831);
and U1325 (N_1325,N_995,N_447);
nor U1326 (N_1326,N_725,N_400);
nand U1327 (N_1327,N_223,N_974);
nor U1328 (N_1328,N_786,N_39);
xor U1329 (N_1329,N_965,N_600);
nor U1330 (N_1330,N_939,N_143);
nand U1331 (N_1331,N_120,N_290);
nor U1332 (N_1332,N_102,N_84);
and U1333 (N_1333,N_774,N_875);
or U1334 (N_1334,N_315,N_489);
or U1335 (N_1335,N_414,N_155);
and U1336 (N_1336,N_866,N_941);
nand U1337 (N_1337,N_792,N_301);
nor U1338 (N_1338,N_706,N_968);
nand U1339 (N_1339,N_870,N_280);
nand U1340 (N_1340,N_726,N_398);
xnor U1341 (N_1341,N_570,N_485);
nor U1342 (N_1342,N_56,N_465);
xor U1343 (N_1343,N_443,N_331);
and U1344 (N_1344,N_496,N_528);
nand U1345 (N_1345,N_659,N_269);
nand U1346 (N_1346,N_823,N_762);
and U1347 (N_1347,N_500,N_25);
and U1348 (N_1348,N_675,N_478);
nor U1349 (N_1349,N_137,N_497);
and U1350 (N_1350,N_48,N_86);
nand U1351 (N_1351,N_620,N_936);
nand U1352 (N_1352,N_221,N_593);
nand U1353 (N_1353,N_213,N_927);
nand U1354 (N_1354,N_813,N_566);
nand U1355 (N_1355,N_785,N_848);
and U1356 (N_1356,N_68,N_582);
and U1357 (N_1357,N_676,N_735);
or U1358 (N_1358,N_654,N_648);
and U1359 (N_1359,N_758,N_335);
nand U1360 (N_1360,N_187,N_242);
or U1361 (N_1361,N_992,N_541);
or U1362 (N_1362,N_445,N_44);
nand U1363 (N_1363,N_288,N_476);
and U1364 (N_1364,N_463,N_953);
and U1365 (N_1365,N_451,N_431);
and U1366 (N_1366,N_772,N_224);
or U1367 (N_1367,N_52,N_403);
and U1368 (N_1368,N_818,N_803);
nor U1369 (N_1369,N_444,N_650);
nand U1370 (N_1370,N_430,N_575);
xor U1371 (N_1371,N_351,N_227);
or U1372 (N_1372,N_728,N_867);
nor U1373 (N_1373,N_544,N_405);
nand U1374 (N_1374,N_185,N_424);
nor U1375 (N_1375,N_902,N_329);
and U1376 (N_1376,N_127,N_720);
nand U1377 (N_1377,N_522,N_76);
or U1378 (N_1378,N_324,N_295);
nor U1379 (N_1379,N_88,N_604);
and U1380 (N_1380,N_271,N_45);
or U1381 (N_1381,N_949,N_189);
nand U1382 (N_1382,N_146,N_428);
xnor U1383 (N_1383,N_236,N_876);
or U1384 (N_1384,N_586,N_594);
nand U1385 (N_1385,N_844,N_612);
nor U1386 (N_1386,N_138,N_966);
nor U1387 (N_1387,N_577,N_297);
xor U1388 (N_1388,N_375,N_29);
nand U1389 (N_1389,N_993,N_17);
xnor U1390 (N_1390,N_498,N_806);
xnor U1391 (N_1391,N_11,N_809);
nor U1392 (N_1392,N_174,N_356);
nand U1393 (N_1393,N_808,N_633);
and U1394 (N_1394,N_661,N_743);
xnor U1395 (N_1395,N_259,N_787);
nor U1396 (N_1396,N_328,N_182);
nor U1397 (N_1397,N_853,N_293);
or U1398 (N_1398,N_216,N_72);
nand U1399 (N_1399,N_888,N_935);
nor U1400 (N_1400,N_307,N_458);
nand U1401 (N_1401,N_262,N_278);
and U1402 (N_1402,N_618,N_542);
nand U1403 (N_1403,N_782,N_433);
nand U1404 (N_1404,N_326,N_917);
nand U1405 (N_1405,N_371,N_527);
xor U1406 (N_1406,N_100,N_370);
and U1407 (N_1407,N_16,N_512);
nand U1408 (N_1408,N_423,N_846);
nor U1409 (N_1409,N_409,N_481);
nor U1410 (N_1410,N_754,N_729);
nand U1411 (N_1411,N_894,N_162);
or U1412 (N_1412,N_901,N_209);
nand U1413 (N_1413,N_344,N_292);
or U1414 (N_1414,N_509,N_814);
and U1415 (N_1415,N_49,N_348);
nor U1416 (N_1416,N_214,N_733);
nand U1417 (N_1417,N_112,N_397);
nor U1418 (N_1418,N_464,N_626);
or U1419 (N_1419,N_153,N_873);
nand U1420 (N_1420,N_850,N_21);
or U1421 (N_1421,N_826,N_560);
or U1422 (N_1422,N_524,N_233);
or U1423 (N_1423,N_12,N_467);
and U1424 (N_1424,N_425,N_0);
or U1425 (N_1425,N_136,N_615);
xnor U1426 (N_1426,N_572,N_361);
nand U1427 (N_1427,N_567,N_970);
and U1428 (N_1428,N_971,N_773);
nor U1429 (N_1429,N_872,N_437);
or U1430 (N_1430,N_448,N_164);
nor U1431 (N_1431,N_51,N_225);
nor U1432 (N_1432,N_678,N_208);
nor U1433 (N_1433,N_206,N_824);
and U1434 (N_1434,N_133,N_816);
and U1435 (N_1435,N_316,N_730);
nand U1436 (N_1436,N_441,N_718);
or U1437 (N_1437,N_406,N_412);
or U1438 (N_1438,N_294,N_264);
or U1439 (N_1439,N_449,N_627);
nand U1440 (N_1440,N_667,N_87);
or U1441 (N_1441,N_977,N_991);
or U1442 (N_1442,N_125,N_237);
xnor U1443 (N_1443,N_404,N_622);
and U1444 (N_1444,N_899,N_916);
or U1445 (N_1445,N_74,N_693);
or U1446 (N_1446,N_671,N_145);
nand U1447 (N_1447,N_795,N_860);
nor U1448 (N_1448,N_252,N_265);
and U1449 (N_1449,N_396,N_440);
or U1450 (N_1450,N_244,N_696);
nor U1451 (N_1451,N_553,N_181);
and U1452 (N_1452,N_614,N_121);
and U1453 (N_1453,N_454,N_184);
xnor U1454 (N_1454,N_554,N_598);
nand U1455 (N_1455,N_113,N_616);
and U1456 (N_1456,N_376,N_779);
or U1457 (N_1457,N_419,N_53);
nor U1458 (N_1458,N_790,N_36);
or U1459 (N_1459,N_962,N_710);
and U1460 (N_1460,N_69,N_312);
and U1461 (N_1461,N_636,N_812);
nand U1462 (N_1462,N_631,N_765);
or U1463 (N_1463,N_766,N_31);
nor U1464 (N_1464,N_277,N_77);
and U1465 (N_1465,N_149,N_304);
nor U1466 (N_1466,N_791,N_253);
nand U1467 (N_1467,N_70,N_241);
and U1468 (N_1468,N_141,N_601);
or U1469 (N_1469,N_90,N_839);
nand U1470 (N_1470,N_550,N_387);
nor U1471 (N_1471,N_877,N_799);
and U1472 (N_1472,N_95,N_921);
nand U1473 (N_1473,N_341,N_981);
or U1474 (N_1474,N_685,N_303);
nor U1475 (N_1475,N_647,N_13);
and U1476 (N_1476,N_151,N_218);
xnor U1477 (N_1477,N_819,N_273);
and U1478 (N_1478,N_309,N_856);
nand U1479 (N_1479,N_377,N_715);
or U1480 (N_1480,N_118,N_268);
nand U1481 (N_1481,N_833,N_173);
nand U1482 (N_1482,N_195,N_623);
nor U1483 (N_1483,N_59,N_245);
and U1484 (N_1484,N_384,N_234);
and U1485 (N_1485,N_3,N_394);
nor U1486 (N_1486,N_656,N_756);
xnor U1487 (N_1487,N_325,N_605);
or U1488 (N_1488,N_591,N_511);
nand U1489 (N_1489,N_486,N_32);
nor U1490 (N_1490,N_199,N_669);
nand U1491 (N_1491,N_741,N_135);
nand U1492 (N_1492,N_938,N_734);
nand U1493 (N_1493,N_602,N_274);
nor U1494 (N_1494,N_755,N_54);
and U1495 (N_1495,N_238,N_313);
nand U1496 (N_1496,N_564,N_193);
nand U1497 (N_1497,N_518,N_841);
and U1498 (N_1498,N_989,N_429);
and U1499 (N_1499,N_721,N_929);
nand U1500 (N_1500,N_273,N_591);
nand U1501 (N_1501,N_238,N_756);
or U1502 (N_1502,N_560,N_586);
or U1503 (N_1503,N_332,N_275);
or U1504 (N_1504,N_483,N_862);
nor U1505 (N_1505,N_809,N_750);
and U1506 (N_1506,N_217,N_183);
xnor U1507 (N_1507,N_791,N_259);
nand U1508 (N_1508,N_337,N_164);
or U1509 (N_1509,N_337,N_473);
or U1510 (N_1510,N_189,N_399);
xor U1511 (N_1511,N_878,N_431);
nor U1512 (N_1512,N_156,N_449);
and U1513 (N_1513,N_554,N_88);
nand U1514 (N_1514,N_326,N_458);
nor U1515 (N_1515,N_76,N_477);
xnor U1516 (N_1516,N_486,N_841);
or U1517 (N_1517,N_364,N_152);
nand U1518 (N_1518,N_861,N_398);
nand U1519 (N_1519,N_448,N_772);
nor U1520 (N_1520,N_424,N_845);
and U1521 (N_1521,N_607,N_442);
nand U1522 (N_1522,N_247,N_651);
nor U1523 (N_1523,N_614,N_436);
or U1524 (N_1524,N_116,N_342);
and U1525 (N_1525,N_602,N_686);
nor U1526 (N_1526,N_585,N_422);
and U1527 (N_1527,N_927,N_126);
and U1528 (N_1528,N_366,N_875);
nand U1529 (N_1529,N_214,N_975);
nand U1530 (N_1530,N_422,N_189);
nor U1531 (N_1531,N_734,N_982);
nor U1532 (N_1532,N_683,N_206);
nor U1533 (N_1533,N_479,N_311);
or U1534 (N_1534,N_848,N_488);
and U1535 (N_1535,N_642,N_465);
xnor U1536 (N_1536,N_830,N_956);
nand U1537 (N_1537,N_245,N_364);
nand U1538 (N_1538,N_220,N_957);
nor U1539 (N_1539,N_112,N_560);
nor U1540 (N_1540,N_727,N_709);
and U1541 (N_1541,N_690,N_710);
and U1542 (N_1542,N_433,N_460);
or U1543 (N_1543,N_877,N_430);
or U1544 (N_1544,N_621,N_447);
nor U1545 (N_1545,N_800,N_185);
or U1546 (N_1546,N_233,N_457);
nand U1547 (N_1547,N_715,N_408);
and U1548 (N_1548,N_875,N_839);
nand U1549 (N_1549,N_756,N_502);
nand U1550 (N_1550,N_122,N_454);
nand U1551 (N_1551,N_198,N_196);
or U1552 (N_1552,N_931,N_87);
or U1553 (N_1553,N_127,N_902);
or U1554 (N_1554,N_873,N_407);
xor U1555 (N_1555,N_815,N_523);
and U1556 (N_1556,N_302,N_880);
nor U1557 (N_1557,N_16,N_899);
or U1558 (N_1558,N_346,N_527);
nand U1559 (N_1559,N_730,N_425);
and U1560 (N_1560,N_840,N_176);
nor U1561 (N_1561,N_936,N_913);
nand U1562 (N_1562,N_370,N_924);
nor U1563 (N_1563,N_636,N_931);
nor U1564 (N_1564,N_305,N_754);
or U1565 (N_1565,N_452,N_355);
and U1566 (N_1566,N_989,N_746);
nand U1567 (N_1567,N_189,N_152);
nor U1568 (N_1568,N_428,N_79);
nor U1569 (N_1569,N_431,N_687);
xor U1570 (N_1570,N_735,N_758);
and U1571 (N_1571,N_82,N_467);
and U1572 (N_1572,N_218,N_942);
nand U1573 (N_1573,N_573,N_411);
or U1574 (N_1574,N_193,N_185);
and U1575 (N_1575,N_451,N_778);
and U1576 (N_1576,N_524,N_424);
nor U1577 (N_1577,N_957,N_139);
nor U1578 (N_1578,N_599,N_699);
and U1579 (N_1579,N_690,N_122);
nand U1580 (N_1580,N_109,N_381);
nand U1581 (N_1581,N_840,N_822);
and U1582 (N_1582,N_164,N_178);
and U1583 (N_1583,N_203,N_471);
nor U1584 (N_1584,N_183,N_989);
nor U1585 (N_1585,N_247,N_182);
nor U1586 (N_1586,N_734,N_197);
or U1587 (N_1587,N_499,N_257);
nor U1588 (N_1588,N_873,N_712);
and U1589 (N_1589,N_550,N_814);
nor U1590 (N_1590,N_438,N_333);
nand U1591 (N_1591,N_794,N_3);
or U1592 (N_1592,N_151,N_999);
and U1593 (N_1593,N_668,N_580);
or U1594 (N_1594,N_502,N_97);
xnor U1595 (N_1595,N_188,N_607);
or U1596 (N_1596,N_520,N_606);
nand U1597 (N_1597,N_384,N_808);
nand U1598 (N_1598,N_418,N_601);
nand U1599 (N_1599,N_57,N_356);
xor U1600 (N_1600,N_734,N_199);
nand U1601 (N_1601,N_903,N_79);
nor U1602 (N_1602,N_707,N_796);
or U1603 (N_1603,N_224,N_369);
and U1604 (N_1604,N_473,N_59);
or U1605 (N_1605,N_897,N_536);
nor U1606 (N_1606,N_242,N_423);
nor U1607 (N_1607,N_648,N_714);
nand U1608 (N_1608,N_621,N_997);
xnor U1609 (N_1609,N_562,N_85);
nand U1610 (N_1610,N_878,N_698);
and U1611 (N_1611,N_500,N_71);
nor U1612 (N_1612,N_727,N_25);
or U1613 (N_1613,N_863,N_412);
xor U1614 (N_1614,N_865,N_840);
nand U1615 (N_1615,N_747,N_831);
nand U1616 (N_1616,N_404,N_390);
nor U1617 (N_1617,N_328,N_303);
or U1618 (N_1618,N_944,N_297);
or U1619 (N_1619,N_361,N_597);
or U1620 (N_1620,N_972,N_710);
nor U1621 (N_1621,N_426,N_527);
or U1622 (N_1622,N_133,N_330);
xor U1623 (N_1623,N_554,N_468);
and U1624 (N_1624,N_739,N_247);
xor U1625 (N_1625,N_355,N_573);
and U1626 (N_1626,N_297,N_931);
nand U1627 (N_1627,N_374,N_778);
or U1628 (N_1628,N_37,N_131);
nor U1629 (N_1629,N_124,N_592);
nor U1630 (N_1630,N_288,N_346);
and U1631 (N_1631,N_463,N_614);
or U1632 (N_1632,N_86,N_26);
nor U1633 (N_1633,N_821,N_776);
nor U1634 (N_1634,N_715,N_66);
and U1635 (N_1635,N_402,N_59);
nor U1636 (N_1636,N_162,N_102);
and U1637 (N_1637,N_534,N_494);
nand U1638 (N_1638,N_382,N_859);
or U1639 (N_1639,N_823,N_657);
and U1640 (N_1640,N_878,N_380);
nor U1641 (N_1641,N_93,N_352);
nand U1642 (N_1642,N_728,N_53);
or U1643 (N_1643,N_83,N_392);
xnor U1644 (N_1644,N_543,N_621);
nand U1645 (N_1645,N_790,N_583);
xnor U1646 (N_1646,N_698,N_679);
nand U1647 (N_1647,N_457,N_527);
nand U1648 (N_1648,N_593,N_249);
and U1649 (N_1649,N_920,N_322);
nand U1650 (N_1650,N_22,N_179);
nand U1651 (N_1651,N_184,N_984);
nand U1652 (N_1652,N_573,N_902);
and U1653 (N_1653,N_571,N_136);
and U1654 (N_1654,N_298,N_498);
nand U1655 (N_1655,N_215,N_887);
nor U1656 (N_1656,N_458,N_358);
nand U1657 (N_1657,N_647,N_107);
and U1658 (N_1658,N_871,N_710);
or U1659 (N_1659,N_485,N_35);
xnor U1660 (N_1660,N_379,N_414);
and U1661 (N_1661,N_826,N_791);
and U1662 (N_1662,N_298,N_111);
and U1663 (N_1663,N_563,N_338);
nand U1664 (N_1664,N_431,N_972);
nor U1665 (N_1665,N_269,N_32);
nand U1666 (N_1666,N_405,N_366);
or U1667 (N_1667,N_777,N_680);
nand U1668 (N_1668,N_978,N_498);
nand U1669 (N_1669,N_366,N_755);
or U1670 (N_1670,N_266,N_837);
nor U1671 (N_1671,N_997,N_986);
and U1672 (N_1672,N_386,N_211);
nand U1673 (N_1673,N_222,N_116);
nand U1674 (N_1674,N_469,N_221);
nand U1675 (N_1675,N_680,N_883);
or U1676 (N_1676,N_582,N_164);
nor U1677 (N_1677,N_452,N_665);
nor U1678 (N_1678,N_684,N_695);
or U1679 (N_1679,N_413,N_574);
or U1680 (N_1680,N_103,N_626);
nand U1681 (N_1681,N_573,N_378);
and U1682 (N_1682,N_305,N_308);
nand U1683 (N_1683,N_200,N_199);
and U1684 (N_1684,N_415,N_605);
and U1685 (N_1685,N_326,N_264);
or U1686 (N_1686,N_136,N_177);
and U1687 (N_1687,N_496,N_871);
nand U1688 (N_1688,N_491,N_492);
nand U1689 (N_1689,N_32,N_586);
nand U1690 (N_1690,N_223,N_347);
nor U1691 (N_1691,N_439,N_54);
or U1692 (N_1692,N_396,N_301);
and U1693 (N_1693,N_388,N_12);
and U1694 (N_1694,N_816,N_782);
and U1695 (N_1695,N_631,N_28);
nand U1696 (N_1696,N_909,N_402);
and U1697 (N_1697,N_140,N_437);
or U1698 (N_1698,N_314,N_324);
or U1699 (N_1699,N_121,N_456);
nand U1700 (N_1700,N_311,N_674);
and U1701 (N_1701,N_823,N_368);
nand U1702 (N_1702,N_946,N_889);
or U1703 (N_1703,N_194,N_835);
or U1704 (N_1704,N_926,N_179);
nor U1705 (N_1705,N_444,N_131);
nand U1706 (N_1706,N_949,N_224);
nand U1707 (N_1707,N_489,N_607);
nor U1708 (N_1708,N_131,N_829);
or U1709 (N_1709,N_304,N_498);
and U1710 (N_1710,N_458,N_79);
nand U1711 (N_1711,N_62,N_611);
or U1712 (N_1712,N_991,N_663);
nand U1713 (N_1713,N_580,N_886);
nor U1714 (N_1714,N_974,N_851);
or U1715 (N_1715,N_644,N_830);
nand U1716 (N_1716,N_731,N_942);
or U1717 (N_1717,N_508,N_488);
xor U1718 (N_1718,N_217,N_426);
nor U1719 (N_1719,N_834,N_362);
xnor U1720 (N_1720,N_959,N_461);
and U1721 (N_1721,N_934,N_379);
nand U1722 (N_1722,N_278,N_985);
nand U1723 (N_1723,N_28,N_856);
or U1724 (N_1724,N_116,N_553);
nor U1725 (N_1725,N_707,N_509);
and U1726 (N_1726,N_635,N_396);
nand U1727 (N_1727,N_297,N_149);
nor U1728 (N_1728,N_16,N_126);
or U1729 (N_1729,N_142,N_697);
nand U1730 (N_1730,N_526,N_946);
nand U1731 (N_1731,N_703,N_600);
or U1732 (N_1732,N_781,N_577);
xor U1733 (N_1733,N_695,N_793);
or U1734 (N_1734,N_231,N_154);
nand U1735 (N_1735,N_290,N_476);
xnor U1736 (N_1736,N_505,N_20);
nand U1737 (N_1737,N_513,N_263);
xor U1738 (N_1738,N_142,N_746);
nand U1739 (N_1739,N_478,N_701);
and U1740 (N_1740,N_960,N_705);
and U1741 (N_1741,N_446,N_780);
nand U1742 (N_1742,N_136,N_114);
nor U1743 (N_1743,N_694,N_511);
or U1744 (N_1744,N_822,N_544);
nor U1745 (N_1745,N_454,N_5);
xnor U1746 (N_1746,N_268,N_363);
nand U1747 (N_1747,N_23,N_399);
nor U1748 (N_1748,N_66,N_452);
or U1749 (N_1749,N_140,N_250);
and U1750 (N_1750,N_438,N_252);
nand U1751 (N_1751,N_246,N_980);
or U1752 (N_1752,N_712,N_46);
or U1753 (N_1753,N_605,N_69);
and U1754 (N_1754,N_506,N_204);
nand U1755 (N_1755,N_106,N_302);
xor U1756 (N_1756,N_597,N_66);
and U1757 (N_1757,N_234,N_264);
nor U1758 (N_1758,N_927,N_713);
or U1759 (N_1759,N_473,N_882);
or U1760 (N_1760,N_850,N_890);
and U1761 (N_1761,N_957,N_349);
or U1762 (N_1762,N_999,N_120);
nand U1763 (N_1763,N_605,N_995);
nand U1764 (N_1764,N_319,N_200);
nand U1765 (N_1765,N_234,N_846);
nand U1766 (N_1766,N_366,N_783);
nand U1767 (N_1767,N_873,N_269);
nand U1768 (N_1768,N_376,N_81);
or U1769 (N_1769,N_336,N_971);
and U1770 (N_1770,N_603,N_779);
and U1771 (N_1771,N_5,N_639);
nand U1772 (N_1772,N_885,N_178);
or U1773 (N_1773,N_173,N_979);
and U1774 (N_1774,N_887,N_579);
or U1775 (N_1775,N_397,N_791);
and U1776 (N_1776,N_545,N_318);
and U1777 (N_1777,N_490,N_77);
nor U1778 (N_1778,N_954,N_800);
nor U1779 (N_1779,N_895,N_342);
nand U1780 (N_1780,N_426,N_368);
and U1781 (N_1781,N_157,N_626);
and U1782 (N_1782,N_609,N_53);
and U1783 (N_1783,N_83,N_881);
xor U1784 (N_1784,N_722,N_932);
nor U1785 (N_1785,N_14,N_339);
nand U1786 (N_1786,N_521,N_571);
xor U1787 (N_1787,N_728,N_177);
nand U1788 (N_1788,N_890,N_696);
and U1789 (N_1789,N_502,N_875);
nand U1790 (N_1790,N_958,N_158);
xnor U1791 (N_1791,N_702,N_573);
nor U1792 (N_1792,N_570,N_967);
nand U1793 (N_1793,N_825,N_305);
and U1794 (N_1794,N_938,N_337);
nand U1795 (N_1795,N_509,N_663);
nor U1796 (N_1796,N_724,N_892);
or U1797 (N_1797,N_703,N_623);
nand U1798 (N_1798,N_71,N_865);
and U1799 (N_1799,N_824,N_978);
and U1800 (N_1800,N_655,N_807);
nor U1801 (N_1801,N_957,N_12);
nor U1802 (N_1802,N_144,N_747);
nor U1803 (N_1803,N_821,N_309);
and U1804 (N_1804,N_530,N_818);
and U1805 (N_1805,N_869,N_294);
nand U1806 (N_1806,N_76,N_408);
and U1807 (N_1807,N_798,N_900);
and U1808 (N_1808,N_794,N_535);
nand U1809 (N_1809,N_98,N_203);
nor U1810 (N_1810,N_667,N_728);
or U1811 (N_1811,N_673,N_987);
and U1812 (N_1812,N_466,N_396);
and U1813 (N_1813,N_166,N_467);
and U1814 (N_1814,N_869,N_410);
nand U1815 (N_1815,N_688,N_96);
or U1816 (N_1816,N_619,N_149);
nor U1817 (N_1817,N_423,N_103);
nand U1818 (N_1818,N_545,N_473);
or U1819 (N_1819,N_673,N_114);
or U1820 (N_1820,N_152,N_864);
or U1821 (N_1821,N_414,N_275);
nor U1822 (N_1822,N_48,N_870);
nand U1823 (N_1823,N_116,N_224);
or U1824 (N_1824,N_733,N_370);
nand U1825 (N_1825,N_790,N_649);
and U1826 (N_1826,N_769,N_338);
or U1827 (N_1827,N_426,N_285);
or U1828 (N_1828,N_556,N_676);
and U1829 (N_1829,N_805,N_418);
nand U1830 (N_1830,N_858,N_545);
and U1831 (N_1831,N_933,N_122);
xnor U1832 (N_1832,N_91,N_519);
nand U1833 (N_1833,N_186,N_799);
or U1834 (N_1834,N_603,N_110);
and U1835 (N_1835,N_987,N_819);
nand U1836 (N_1836,N_801,N_194);
nor U1837 (N_1837,N_671,N_246);
nor U1838 (N_1838,N_781,N_961);
xor U1839 (N_1839,N_537,N_433);
and U1840 (N_1840,N_779,N_708);
and U1841 (N_1841,N_67,N_25);
nand U1842 (N_1842,N_962,N_131);
nor U1843 (N_1843,N_145,N_689);
and U1844 (N_1844,N_175,N_47);
nor U1845 (N_1845,N_907,N_866);
nor U1846 (N_1846,N_480,N_280);
nor U1847 (N_1847,N_364,N_326);
nand U1848 (N_1848,N_32,N_531);
or U1849 (N_1849,N_216,N_198);
nand U1850 (N_1850,N_154,N_500);
nor U1851 (N_1851,N_788,N_490);
nand U1852 (N_1852,N_829,N_355);
nor U1853 (N_1853,N_431,N_400);
nand U1854 (N_1854,N_862,N_754);
nand U1855 (N_1855,N_448,N_433);
nor U1856 (N_1856,N_690,N_644);
and U1857 (N_1857,N_723,N_684);
nand U1858 (N_1858,N_351,N_534);
or U1859 (N_1859,N_457,N_355);
or U1860 (N_1860,N_212,N_5);
nand U1861 (N_1861,N_668,N_428);
or U1862 (N_1862,N_693,N_769);
or U1863 (N_1863,N_131,N_842);
or U1864 (N_1864,N_936,N_265);
nor U1865 (N_1865,N_702,N_982);
and U1866 (N_1866,N_206,N_820);
nand U1867 (N_1867,N_166,N_337);
and U1868 (N_1868,N_336,N_112);
or U1869 (N_1869,N_949,N_202);
and U1870 (N_1870,N_174,N_30);
or U1871 (N_1871,N_568,N_233);
and U1872 (N_1872,N_475,N_567);
or U1873 (N_1873,N_13,N_556);
nand U1874 (N_1874,N_593,N_285);
or U1875 (N_1875,N_730,N_935);
nand U1876 (N_1876,N_366,N_457);
and U1877 (N_1877,N_344,N_260);
and U1878 (N_1878,N_757,N_250);
and U1879 (N_1879,N_526,N_540);
xnor U1880 (N_1880,N_881,N_985);
and U1881 (N_1881,N_992,N_287);
nand U1882 (N_1882,N_493,N_678);
or U1883 (N_1883,N_996,N_880);
and U1884 (N_1884,N_372,N_525);
xor U1885 (N_1885,N_635,N_450);
or U1886 (N_1886,N_397,N_593);
xnor U1887 (N_1887,N_920,N_106);
nor U1888 (N_1888,N_55,N_46);
nor U1889 (N_1889,N_658,N_895);
or U1890 (N_1890,N_517,N_893);
nor U1891 (N_1891,N_805,N_943);
and U1892 (N_1892,N_641,N_631);
nor U1893 (N_1893,N_819,N_744);
nand U1894 (N_1894,N_479,N_341);
nand U1895 (N_1895,N_215,N_804);
nor U1896 (N_1896,N_871,N_368);
nand U1897 (N_1897,N_782,N_872);
nand U1898 (N_1898,N_863,N_20);
nand U1899 (N_1899,N_150,N_651);
and U1900 (N_1900,N_697,N_918);
xnor U1901 (N_1901,N_278,N_582);
and U1902 (N_1902,N_844,N_62);
nand U1903 (N_1903,N_888,N_779);
or U1904 (N_1904,N_730,N_246);
or U1905 (N_1905,N_207,N_664);
or U1906 (N_1906,N_54,N_978);
nor U1907 (N_1907,N_696,N_767);
and U1908 (N_1908,N_538,N_256);
or U1909 (N_1909,N_483,N_34);
and U1910 (N_1910,N_364,N_232);
or U1911 (N_1911,N_560,N_543);
nor U1912 (N_1912,N_342,N_266);
nand U1913 (N_1913,N_259,N_174);
and U1914 (N_1914,N_671,N_784);
and U1915 (N_1915,N_580,N_251);
nor U1916 (N_1916,N_230,N_720);
and U1917 (N_1917,N_312,N_755);
or U1918 (N_1918,N_945,N_254);
nand U1919 (N_1919,N_923,N_552);
nand U1920 (N_1920,N_778,N_97);
and U1921 (N_1921,N_553,N_828);
nand U1922 (N_1922,N_254,N_112);
nand U1923 (N_1923,N_110,N_451);
nor U1924 (N_1924,N_501,N_486);
nand U1925 (N_1925,N_764,N_649);
or U1926 (N_1926,N_958,N_706);
and U1927 (N_1927,N_422,N_250);
nand U1928 (N_1928,N_132,N_545);
nor U1929 (N_1929,N_555,N_437);
and U1930 (N_1930,N_836,N_600);
and U1931 (N_1931,N_348,N_748);
or U1932 (N_1932,N_957,N_860);
nand U1933 (N_1933,N_454,N_471);
nor U1934 (N_1934,N_616,N_399);
and U1935 (N_1935,N_712,N_988);
xnor U1936 (N_1936,N_61,N_228);
or U1937 (N_1937,N_327,N_1);
nor U1938 (N_1938,N_224,N_563);
and U1939 (N_1939,N_55,N_575);
or U1940 (N_1940,N_91,N_30);
nand U1941 (N_1941,N_415,N_360);
and U1942 (N_1942,N_628,N_703);
xnor U1943 (N_1943,N_331,N_631);
nor U1944 (N_1944,N_356,N_309);
nor U1945 (N_1945,N_431,N_619);
or U1946 (N_1946,N_377,N_876);
and U1947 (N_1947,N_926,N_478);
xnor U1948 (N_1948,N_32,N_577);
nand U1949 (N_1949,N_872,N_767);
xnor U1950 (N_1950,N_18,N_930);
nor U1951 (N_1951,N_236,N_951);
or U1952 (N_1952,N_312,N_832);
or U1953 (N_1953,N_87,N_818);
nand U1954 (N_1954,N_346,N_42);
or U1955 (N_1955,N_285,N_675);
nor U1956 (N_1956,N_801,N_425);
nand U1957 (N_1957,N_376,N_415);
or U1958 (N_1958,N_719,N_936);
or U1959 (N_1959,N_819,N_70);
nand U1960 (N_1960,N_789,N_351);
xnor U1961 (N_1961,N_522,N_624);
nand U1962 (N_1962,N_851,N_351);
or U1963 (N_1963,N_722,N_998);
xnor U1964 (N_1964,N_213,N_492);
or U1965 (N_1965,N_696,N_940);
nand U1966 (N_1966,N_775,N_17);
nor U1967 (N_1967,N_552,N_83);
and U1968 (N_1968,N_650,N_184);
nor U1969 (N_1969,N_830,N_983);
and U1970 (N_1970,N_492,N_757);
nand U1971 (N_1971,N_552,N_42);
nor U1972 (N_1972,N_804,N_737);
nand U1973 (N_1973,N_234,N_665);
and U1974 (N_1974,N_371,N_475);
nor U1975 (N_1975,N_435,N_701);
nand U1976 (N_1976,N_430,N_408);
nor U1977 (N_1977,N_828,N_398);
xnor U1978 (N_1978,N_243,N_971);
and U1979 (N_1979,N_320,N_80);
nand U1980 (N_1980,N_682,N_484);
or U1981 (N_1981,N_876,N_564);
nor U1982 (N_1982,N_407,N_54);
nand U1983 (N_1983,N_124,N_43);
nand U1984 (N_1984,N_910,N_121);
nor U1985 (N_1985,N_605,N_550);
nand U1986 (N_1986,N_618,N_734);
or U1987 (N_1987,N_845,N_589);
nor U1988 (N_1988,N_56,N_748);
nor U1989 (N_1989,N_75,N_745);
or U1990 (N_1990,N_967,N_398);
nor U1991 (N_1991,N_556,N_386);
nand U1992 (N_1992,N_563,N_688);
or U1993 (N_1993,N_661,N_210);
or U1994 (N_1994,N_975,N_660);
nand U1995 (N_1995,N_158,N_545);
nand U1996 (N_1996,N_225,N_273);
or U1997 (N_1997,N_261,N_659);
and U1998 (N_1998,N_510,N_363);
nor U1999 (N_1999,N_93,N_689);
nand U2000 (N_2000,N_1261,N_1738);
or U2001 (N_2001,N_1169,N_1897);
and U2002 (N_2002,N_1836,N_1407);
or U2003 (N_2003,N_1633,N_1337);
nor U2004 (N_2004,N_1865,N_1313);
and U2005 (N_2005,N_1213,N_1410);
or U2006 (N_2006,N_1068,N_1581);
and U2007 (N_2007,N_1302,N_1457);
nor U2008 (N_2008,N_1694,N_1136);
nand U2009 (N_2009,N_1853,N_1929);
nand U2010 (N_2010,N_1587,N_1250);
nor U2011 (N_2011,N_1219,N_1265);
xor U2012 (N_2012,N_1554,N_1324);
nor U2013 (N_2013,N_1533,N_1906);
and U2014 (N_2014,N_1059,N_1875);
xnor U2015 (N_2015,N_1297,N_1513);
nand U2016 (N_2016,N_1128,N_1687);
or U2017 (N_2017,N_1076,N_1989);
or U2018 (N_2018,N_1959,N_1537);
and U2019 (N_2019,N_1448,N_1428);
nand U2020 (N_2020,N_1641,N_1636);
nand U2021 (N_2021,N_1553,N_1386);
nand U2022 (N_2022,N_1007,N_1179);
or U2023 (N_2023,N_1682,N_1237);
xor U2024 (N_2024,N_1119,N_1825);
xor U2025 (N_2025,N_1961,N_1615);
nand U2026 (N_2026,N_1305,N_1318);
nand U2027 (N_2027,N_1765,N_1793);
or U2028 (N_2028,N_1440,N_1882);
xor U2029 (N_2029,N_1538,N_1309);
and U2030 (N_2030,N_1366,N_1917);
nand U2031 (N_2031,N_1647,N_1135);
nor U2032 (N_2032,N_1920,N_1823);
and U2033 (N_2033,N_1167,N_1429);
xnor U2034 (N_2034,N_1288,N_1574);
nor U2035 (N_2035,N_1028,N_1388);
nor U2036 (N_2036,N_1595,N_1002);
and U2037 (N_2037,N_1399,N_1283);
or U2038 (N_2038,N_1982,N_1094);
nor U2039 (N_2039,N_1431,N_1042);
or U2040 (N_2040,N_1604,N_1014);
xnor U2041 (N_2041,N_1634,N_1833);
and U2042 (N_2042,N_1709,N_1078);
nor U2043 (N_2043,N_1990,N_1585);
and U2044 (N_2044,N_1083,N_1969);
nand U2045 (N_2045,N_1215,N_1605);
or U2046 (N_2046,N_1684,N_1455);
nor U2047 (N_2047,N_1693,N_1259);
or U2048 (N_2048,N_1948,N_1072);
xor U2049 (N_2049,N_1450,N_1933);
nand U2050 (N_2050,N_1491,N_1433);
nor U2051 (N_2051,N_1252,N_1027);
xor U2052 (N_2052,N_1644,N_1436);
nand U2053 (N_2053,N_1573,N_1844);
or U2054 (N_2054,N_1396,N_1342);
nand U2055 (N_2055,N_1805,N_1474);
and U2056 (N_2056,N_1086,N_1071);
nand U2057 (N_2057,N_1109,N_1276);
xnor U2058 (N_2058,N_1599,N_1998);
or U2059 (N_2059,N_1626,N_1194);
or U2060 (N_2060,N_1905,N_1150);
xor U2061 (N_2061,N_1876,N_1406);
and U2062 (N_2062,N_1800,N_1935);
nor U2063 (N_2063,N_1787,N_1861);
nand U2064 (N_2064,N_1189,N_1154);
or U2065 (N_2065,N_1839,N_1804);
or U2066 (N_2066,N_1015,N_1488);
or U2067 (N_2067,N_1137,N_1767);
xnor U2068 (N_2068,N_1471,N_1303);
or U2069 (N_2069,N_1162,N_1564);
or U2070 (N_2070,N_1207,N_1245);
nand U2071 (N_2071,N_1067,N_1355);
nor U2072 (N_2072,N_1801,N_1608);
nor U2073 (N_2073,N_1481,N_1343);
nor U2074 (N_2074,N_1953,N_1730);
xor U2075 (N_2075,N_1893,N_1120);
xor U2076 (N_2076,N_1971,N_1936);
or U2077 (N_2077,N_1437,N_1589);
nor U2078 (N_2078,N_1826,N_1795);
and U2079 (N_2079,N_1275,N_1300);
or U2080 (N_2080,N_1361,N_1666);
and U2081 (N_2081,N_1430,N_1409);
or U2082 (N_2082,N_1311,N_1307);
or U2083 (N_2083,N_1523,N_1117);
nand U2084 (N_2084,N_1483,N_1079);
nand U2085 (N_2085,N_1240,N_1568);
and U2086 (N_2086,N_1676,N_1112);
xnor U2087 (N_2087,N_1206,N_1911);
nor U2088 (N_2088,N_1824,N_1695);
nand U2089 (N_2089,N_1308,N_1602);
or U2090 (N_2090,N_1711,N_1988);
xor U2091 (N_2091,N_1187,N_1736);
xnor U2092 (N_2092,N_1609,N_1977);
nand U2093 (N_2093,N_1447,N_1133);
and U2094 (N_2094,N_1758,N_1848);
nand U2095 (N_2095,N_1247,N_1543);
and U2096 (N_2096,N_1441,N_1312);
nand U2097 (N_2097,N_1006,N_1997);
nor U2098 (N_2098,N_1847,N_1732);
or U2099 (N_2099,N_1031,N_1766);
or U2100 (N_2100,N_1299,N_1504);
nor U2101 (N_2101,N_1214,N_1367);
nor U2102 (N_2102,N_1364,N_1351);
or U2103 (N_2103,N_1290,N_1895);
nand U2104 (N_2104,N_1547,N_1658);
nor U2105 (N_2105,N_1753,N_1088);
nand U2106 (N_2106,N_1592,N_1390);
and U2107 (N_2107,N_1418,N_1571);
nand U2108 (N_2108,N_1673,N_1768);
nand U2109 (N_2109,N_1151,N_1975);
and U2110 (N_2110,N_1515,N_1304);
or U2111 (N_2111,N_1268,N_1835);
nand U2112 (N_2112,N_1771,N_1204);
or U2113 (N_2113,N_1191,N_1992);
nor U2114 (N_2114,N_1310,N_1130);
and U2115 (N_2115,N_1968,N_1590);
nor U2116 (N_2116,N_1601,N_1664);
nor U2117 (N_2117,N_1883,N_1501);
and U2118 (N_2118,N_1174,N_1340);
xor U2119 (N_2119,N_1082,N_1570);
xor U2120 (N_2120,N_1889,N_1593);
nand U2121 (N_2121,N_1942,N_1873);
nor U2122 (N_2122,N_1862,N_1872);
or U2123 (N_2123,N_1521,N_1444);
nand U2124 (N_2124,N_1255,N_1257);
or U2125 (N_2125,N_1539,N_1322);
and U2126 (N_2126,N_1211,N_1159);
and U2127 (N_2127,N_1350,N_1256);
nand U2128 (N_2128,N_1496,N_1147);
nand U2129 (N_2129,N_1065,N_1476);
or U2130 (N_2130,N_1212,N_1654);
nor U2131 (N_2131,N_1546,N_1084);
xor U2132 (N_2132,N_1231,N_1054);
or U2133 (N_2133,N_1619,N_1131);
or U2134 (N_2134,N_1482,N_1777);
or U2135 (N_2135,N_1157,N_1220);
or U2136 (N_2136,N_1405,N_1336);
nand U2137 (N_2137,N_1691,N_1620);
nor U2138 (N_2138,N_1728,N_1863);
xnor U2139 (N_2139,N_1545,N_1854);
and U2140 (N_2140,N_1218,N_1815);
or U2141 (N_2141,N_1706,N_1822);
nand U2142 (N_2142,N_1487,N_1505);
nand U2143 (N_2143,N_1026,N_1924);
and U2144 (N_2144,N_1962,N_1722);
or U2145 (N_2145,N_1780,N_1395);
xnor U2146 (N_2146,N_1716,N_1831);
nor U2147 (N_2147,N_1280,N_1281);
or U2148 (N_2148,N_1489,N_1923);
and U2149 (N_2149,N_1560,N_1420);
nor U2150 (N_2150,N_1637,N_1868);
or U2151 (N_2151,N_1566,N_1980);
and U2152 (N_2152,N_1879,N_1675);
nor U2153 (N_2153,N_1463,N_1878);
xor U2154 (N_2154,N_1829,N_1477);
and U2155 (N_2155,N_1049,N_1331);
or U2156 (N_2156,N_1121,N_1392);
and U2157 (N_2157,N_1751,N_1473);
or U2158 (N_2158,N_1421,N_1176);
nand U2159 (N_2159,N_1115,N_1449);
nor U2160 (N_2160,N_1894,N_1165);
and U2161 (N_2161,N_1660,N_1552);
or U2162 (N_2162,N_1458,N_1727);
nand U2163 (N_2163,N_1144,N_1438);
nor U2164 (N_2164,N_1166,N_1970);
nor U2165 (N_2165,N_1346,N_1565);
nand U2166 (N_2166,N_1417,N_1814);
nor U2167 (N_2167,N_1618,N_1271);
nand U2168 (N_2168,N_1472,N_1559);
or U2169 (N_2169,N_1285,N_1202);
nor U2170 (N_2170,N_1485,N_1186);
and U2171 (N_2171,N_1628,N_1649);
and U2172 (N_2172,N_1659,N_1784);
and U2173 (N_2173,N_1680,N_1958);
and U2174 (N_2174,N_1750,N_1129);
nor U2175 (N_2175,N_1264,N_1789);
nor U2176 (N_2176,N_1379,N_1535);
nor U2177 (N_2177,N_1398,N_1293);
nand U2178 (N_2178,N_1323,N_1512);
or U2179 (N_2179,N_1511,N_1851);
nand U2180 (N_2180,N_1575,N_1631);
and U2181 (N_2181,N_1462,N_1389);
or U2182 (N_2182,N_1416,N_1532);
xnor U2183 (N_2183,N_1843,N_1001);
nor U2184 (N_2184,N_1412,N_1029);
or U2185 (N_2185,N_1950,N_1772);
nor U2186 (N_2186,N_1248,N_1762);
or U2187 (N_2187,N_1177,N_1236);
nor U2188 (N_2188,N_1966,N_1170);
nand U2189 (N_2189,N_1233,N_1951);
nor U2190 (N_2190,N_1519,N_1325);
or U2191 (N_2191,N_1500,N_1229);
and U2192 (N_2192,N_1914,N_1005);
xor U2193 (N_2193,N_1153,N_1909);
nor U2194 (N_2194,N_1284,N_1037);
nand U2195 (N_2195,N_1918,N_1080);
nor U2196 (N_2196,N_1465,N_1763);
nor U2197 (N_2197,N_1742,N_1712);
nand U2198 (N_2198,N_1945,N_1315);
or U2199 (N_2199,N_1413,N_1850);
and U2200 (N_2200,N_1880,N_1098);
xor U2201 (N_2201,N_1579,N_1432);
or U2202 (N_2202,N_1734,N_1737);
and U2203 (N_2203,N_1239,N_1104);
nor U2204 (N_2204,N_1341,N_1442);
xor U2205 (N_2205,N_1192,N_1671);
xor U2206 (N_2206,N_1820,N_1516);
or U2207 (N_2207,N_1576,N_1373);
nor U2208 (N_2208,N_1741,N_1749);
nor U2209 (N_2209,N_1612,N_1941);
and U2210 (N_2210,N_1838,N_1955);
nor U2211 (N_2211,N_1607,N_1892);
nand U2212 (N_2212,N_1891,N_1884);
xor U2213 (N_2213,N_1978,N_1902);
nand U2214 (N_2214,N_1118,N_1360);
nor U2215 (N_2215,N_1907,N_1032);
nor U2216 (N_2216,N_1205,N_1306);
or U2217 (N_2217,N_1705,N_1222);
or U2218 (N_2218,N_1164,N_1799);
xnor U2219 (N_2219,N_1099,N_1138);
and U2220 (N_2220,N_1454,N_1611);
and U2221 (N_2221,N_1731,N_1616);
nor U2222 (N_2222,N_1720,N_1258);
nor U2223 (N_2223,N_1755,N_1163);
or U2224 (N_2224,N_1414,N_1846);
nand U2225 (N_2225,N_1286,N_1217);
nor U2226 (N_2226,N_1841,N_1690);
nor U2227 (N_2227,N_1278,N_1209);
nand U2228 (N_2228,N_1445,N_1555);
or U2229 (N_2229,N_1930,N_1655);
nor U2230 (N_2230,N_1494,N_1467);
nand U2231 (N_2231,N_1100,N_1774);
or U2232 (N_2232,N_1996,N_1362);
nor U2233 (N_2233,N_1520,N_1842);
nor U2234 (N_2234,N_1719,N_1885);
nand U2235 (N_2235,N_1542,N_1888);
nand U2236 (N_2236,N_1434,N_1672);
and U2237 (N_2237,N_1044,N_1639);
and U2238 (N_2238,N_1188,N_1740);
and U2239 (N_2239,N_1085,N_1810);
and U2240 (N_2240,N_1073,N_1106);
and U2241 (N_2241,N_1141,N_1794);
nand U2242 (N_2242,N_1677,N_1870);
and U2243 (N_2243,N_1139,N_1613);
nand U2244 (N_2244,N_1499,N_1580);
nand U2245 (N_2245,N_1723,N_1514);
or U2246 (N_2246,N_1643,N_1979);
nor U2247 (N_2247,N_1943,N_1503);
nand U2248 (N_2248,N_1697,N_1277);
nor U2249 (N_2249,N_1715,N_1320);
nor U2250 (N_2250,N_1887,N_1509);
and U2251 (N_2251,N_1175,N_1940);
and U2252 (N_2252,N_1725,N_1289);
xor U2253 (N_2253,N_1156,N_1095);
nand U2254 (N_2254,N_1058,N_1498);
nand U2255 (N_2255,N_1745,N_1426);
nand U2256 (N_2256,N_1551,N_1898);
nand U2257 (N_2257,N_1803,N_1279);
xnor U2258 (N_2258,N_1419,N_1813);
and U2259 (N_2259,N_1965,N_1916);
or U2260 (N_2260,N_1321,N_1928);
nand U2261 (N_2261,N_1852,N_1232);
and U2262 (N_2262,N_1912,N_1267);
and U2263 (N_2263,N_1699,N_1010);
and U2264 (N_2264,N_1017,N_1524);
nand U2265 (N_2265,N_1600,N_1781);
nor U2266 (N_2266,N_1710,N_1123);
or U2267 (N_2267,N_1347,N_1796);
or U2268 (N_2268,N_1773,N_1225);
nor U2269 (N_2269,N_1769,N_1748);
and U2270 (N_2270,N_1060,N_1039);
nand U2271 (N_2271,N_1563,N_1754);
xnor U2272 (N_2272,N_1226,N_1292);
nand U2273 (N_2273,N_1266,N_1077);
nor U2274 (N_2274,N_1466,N_1185);
nand U2275 (N_2275,N_1234,N_1196);
nand U2276 (N_2276,N_1158,N_1908);
nand U2277 (N_2277,N_1770,N_1451);
or U2278 (N_2278,N_1113,N_1263);
nand U2279 (N_2279,N_1807,N_1921);
xnor U2280 (N_2280,N_1886,N_1241);
and U2281 (N_2281,N_1849,N_1103);
or U2282 (N_2282,N_1922,N_1934);
nor U2283 (N_2283,N_1733,N_1013);
and U2284 (N_2284,N_1464,N_1022);
xnor U2285 (N_2285,N_1761,N_1561);
nor U2286 (N_2286,N_1809,N_1183);
nor U2287 (N_2287,N_1759,N_1200);
and U2288 (N_2288,N_1160,N_1714);
nand U2289 (N_2289,N_1506,N_1425);
nor U2290 (N_2290,N_1621,N_1453);
xor U2291 (N_2291,N_1717,N_1785);
and U2292 (N_2292,N_1184,N_1066);
nand U2293 (N_2293,N_1377,N_1370);
or U2294 (N_2294,N_1008,N_1692);
and U2295 (N_2295,N_1021,N_1333);
nand U2296 (N_2296,N_1195,N_1171);
nor U2297 (N_2297,N_1735,N_1662);
nor U2298 (N_2298,N_1915,N_1492);
nand U2299 (N_2299,N_1210,N_1228);
and U2300 (N_2300,N_1287,N_1011);
and U2301 (N_2301,N_1871,N_1480);
nor U2302 (N_2302,N_1125,N_1208);
and U2303 (N_2303,N_1790,N_1630);
nand U2304 (N_2304,N_1557,N_1816);
nor U2305 (N_2305,N_1422,N_1055);
xor U2306 (N_2306,N_1830,N_1925);
nand U2307 (N_2307,N_1376,N_1142);
and U2308 (N_2308,N_1927,N_1316);
nor U2309 (N_2309,N_1627,N_1704);
nand U2310 (N_2310,N_1274,N_1976);
nand U2311 (N_2311,N_1132,N_1269);
and U2312 (N_2312,N_1378,N_1344);
nand U2313 (N_2313,N_1901,N_1069);
and U2314 (N_2314,N_1622,N_1064);
nand U2315 (N_2315,N_1775,N_1262);
nor U2316 (N_2316,N_1363,N_1791);
and U2317 (N_2317,N_1470,N_1629);
or U2318 (N_2318,N_1949,N_1057);
nand U2319 (N_2319,N_1974,N_1798);
nand U2320 (N_2320,N_1954,N_1338);
and U2321 (N_2321,N_1033,N_1148);
xnor U2322 (N_2322,N_1384,N_1349);
or U2323 (N_2323,N_1235,N_1528);
and U2324 (N_2324,N_1686,N_1272);
or U2325 (N_2325,N_1296,N_1572);
nand U2326 (N_2326,N_1030,N_1089);
nor U2327 (N_2327,N_1614,N_1642);
nor U2328 (N_2328,N_1645,N_1653);
or U2329 (N_2329,N_1327,N_1903);
nand U2330 (N_2330,N_1837,N_1536);
nor U2331 (N_2331,N_1696,N_1380);
or U2332 (N_2332,N_1172,N_1294);
xnor U2333 (N_2333,N_1866,N_1701);
and U2334 (N_2334,N_1354,N_1411);
nand U2335 (N_2335,N_1708,N_1531);
nand U2336 (N_2336,N_1840,N_1540);
xor U2337 (N_2337,N_1126,N_1041);
xnor U2338 (N_2338,N_1995,N_1910);
nand U2339 (N_2339,N_1397,N_1238);
nand U2340 (N_2340,N_1385,N_1867);
xnor U2341 (N_2341,N_1502,N_1678);
or U2342 (N_2342,N_1484,N_1534);
or U2343 (N_2343,N_1919,N_1023);
and U2344 (N_2344,N_1063,N_1522);
and U2345 (N_2345,N_1724,N_1960);
and U2346 (N_2346,N_1408,N_1198);
nor U2347 (N_2347,N_1253,N_1778);
nor U2348 (N_2348,N_1375,N_1983);
nor U2349 (N_2349,N_1596,N_1819);
nand U2350 (N_2350,N_1469,N_1097);
nand U2351 (N_2351,N_1947,N_1102);
or U2352 (N_2352,N_1330,N_1591);
and U2353 (N_2353,N_1096,N_1365);
nand U2354 (N_2354,N_1567,N_1973);
or U2355 (N_2355,N_1203,N_1193);
nor U2356 (N_2356,N_1244,N_1981);
or U2357 (N_2357,N_1617,N_1348);
nor U2358 (N_2358,N_1105,N_1702);
nor U2359 (N_2359,N_1400,N_1896);
nor U2360 (N_2360,N_1707,N_1890);
and U2361 (N_2361,N_1757,N_1270);
nand U2362 (N_2362,N_1000,N_1352);
nand U2363 (N_2363,N_1683,N_1404);
or U2364 (N_2364,N_1452,N_1739);
nand U2365 (N_2365,N_1669,N_1254);
nand U2366 (N_2366,N_1070,N_1797);
nand U2367 (N_2367,N_1081,N_1689);
nand U2368 (N_2368,N_1858,N_1549);
or U2369 (N_2369,N_1597,N_1952);
nor U2370 (N_2370,N_1859,N_1374);
nand U2371 (N_2371,N_1319,N_1173);
or U2372 (N_2372,N_1415,N_1756);
or U2373 (N_2373,N_1834,N_1043);
or U2374 (N_2374,N_1273,N_1991);
xor U2375 (N_2375,N_1040,N_1517);
nor U2376 (N_2376,N_1811,N_1776);
and U2377 (N_2377,N_1985,N_1140);
or U2378 (N_2378,N_1821,N_1459);
nor U2379 (N_2379,N_1199,N_1446);
nor U2380 (N_2380,N_1314,N_1510);
nand U2381 (N_2381,N_1074,N_1201);
xor U2382 (N_2382,N_1490,N_1382);
nand U2383 (N_2383,N_1984,N_1899);
nand U2384 (N_2384,N_1881,N_1291);
nor U2385 (N_2385,N_1016,N_1146);
or U2386 (N_2386,N_1004,N_1393);
or U2387 (N_2387,N_1034,N_1178);
and U2388 (N_2388,N_1223,N_1792);
nand U2389 (N_2389,N_1541,N_1588);
nand U2390 (N_2390,N_1053,N_1904);
nor U2391 (N_2391,N_1746,N_1525);
nand U2392 (N_2392,N_1827,N_1391);
nand U2393 (N_2393,N_1703,N_1038);
and U2394 (N_2394,N_1260,N_1443);
and U2395 (N_2395,N_1243,N_1856);
or U2396 (N_2396,N_1817,N_1145);
or U2397 (N_2397,N_1578,N_1635);
and U2398 (N_2398,N_1623,N_1427);
nand U2399 (N_2399,N_1598,N_1946);
nand U2400 (N_2400,N_1012,N_1061);
nor U2401 (N_2401,N_1926,N_1558);
and U2402 (N_2402,N_1665,N_1246);
nor U2403 (N_2403,N_1548,N_1994);
xor U2404 (N_2404,N_1092,N_1874);
nor U2405 (N_2405,N_1045,N_1181);
and U2406 (N_2406,N_1227,N_1582);
nand U2407 (N_2407,N_1050,N_1752);
nand U2408 (N_2408,N_1047,N_1122);
nor U2409 (N_2409,N_1230,N_1329);
and U2410 (N_2410,N_1216,N_1812);
nand U2411 (N_2411,N_1806,N_1134);
and U2412 (N_2412,N_1368,N_1779);
nor U2413 (N_2413,N_1624,N_1544);
or U2414 (N_2414,N_1251,N_1357);
or U2415 (N_2415,N_1845,N_1685);
nor U2416 (N_2416,N_1090,N_1625);
nor U2417 (N_2417,N_1190,N_1650);
nor U2418 (N_2418,N_1486,N_1025);
and U2419 (N_2419,N_1149,N_1584);
xor U2420 (N_2420,N_1298,N_1056);
nor U2421 (N_2421,N_1938,N_1594);
and U2422 (N_2422,N_1124,N_1944);
or U2423 (N_2423,N_1111,N_1802);
and U2424 (N_2424,N_1091,N_1046);
nor U2425 (N_2425,N_1221,N_1718);
and U2426 (N_2426,N_1610,N_1729);
nand U2427 (N_2427,N_1864,N_1497);
and U2428 (N_2428,N_1180,N_1743);
and U2429 (N_2429,N_1024,N_1529);
or U2430 (N_2430,N_1358,N_1661);
or U2431 (N_2431,N_1987,N_1435);
nand U2432 (N_2432,N_1632,N_1108);
nor U2433 (N_2433,N_1857,N_1828);
nand U2434 (N_2434,N_1869,N_1656);
nor U2435 (N_2435,N_1913,N_1093);
xnor U2436 (N_2436,N_1900,N_1479);
nor U2437 (N_2437,N_1155,N_1832);
and U2438 (N_2438,N_1401,N_1999);
and U2439 (N_2439,N_1493,N_1439);
xnor U2440 (N_2440,N_1663,N_1424);
nor U2441 (N_2441,N_1651,N_1667);
xor U2442 (N_2442,N_1688,N_1353);
or U2443 (N_2443,N_1478,N_1224);
or U2444 (N_2444,N_1993,N_1713);
and U2445 (N_2445,N_1606,N_1048);
xnor U2446 (N_2446,N_1957,N_1116);
nand U2447 (N_2447,N_1668,N_1674);
or U2448 (N_2448,N_1698,N_1087);
or U2449 (N_2449,N_1726,N_1670);
or U2450 (N_2450,N_1461,N_1383);
xnor U2451 (N_2451,N_1508,N_1681);
or U2452 (N_2452,N_1402,N_1937);
and U2453 (N_2453,N_1855,N_1507);
and U2454 (N_2454,N_1062,N_1586);
or U2455 (N_2455,N_1956,N_1423);
and U2456 (N_2456,N_1583,N_1550);
or U2457 (N_2457,N_1051,N_1328);
and U2458 (N_2458,N_1019,N_1110);
xor U2459 (N_2459,N_1967,N_1036);
nor U2460 (N_2460,N_1468,N_1760);
and U2461 (N_2461,N_1526,N_1657);
and U2462 (N_2462,N_1475,N_1783);
xor U2463 (N_2463,N_1403,N_1197);
and U2464 (N_2464,N_1527,N_1931);
nor U2465 (N_2465,N_1556,N_1101);
nand U2466 (N_2466,N_1282,N_1652);
and U2467 (N_2467,N_1182,N_1700);
xor U2468 (N_2468,N_1932,N_1371);
and U2469 (N_2469,N_1052,N_1939);
or U2470 (N_2470,N_1114,N_1003);
or U2471 (N_2471,N_1356,N_1679);
nand U2472 (N_2472,N_1877,N_1372);
nand U2473 (N_2473,N_1721,N_1301);
nand U2474 (N_2474,N_1518,N_1638);
and U2475 (N_2475,N_1786,N_1035);
and U2476 (N_2476,N_1335,N_1788);
nor U2477 (N_2477,N_1860,N_1381);
nor U2478 (N_2478,N_1332,N_1562);
or U2479 (N_2479,N_1747,N_1782);
nand U2480 (N_2480,N_1569,N_1744);
and U2481 (N_2481,N_1577,N_1009);
nand U2482 (N_2482,N_1646,N_1818);
and U2483 (N_2483,N_1460,N_1369);
nor U2484 (N_2484,N_1986,N_1242);
nor U2485 (N_2485,N_1972,N_1964);
or U2486 (N_2486,N_1168,N_1394);
or U2487 (N_2487,N_1326,N_1143);
or U2488 (N_2488,N_1456,N_1295);
or U2489 (N_2489,N_1603,N_1648);
nand U2490 (N_2490,N_1018,N_1107);
and U2491 (N_2491,N_1387,N_1334);
or U2492 (N_2492,N_1161,N_1075);
xor U2493 (N_2493,N_1359,N_1530);
nand U2494 (N_2494,N_1495,N_1249);
or U2495 (N_2495,N_1339,N_1764);
nor U2496 (N_2496,N_1020,N_1127);
and U2497 (N_2497,N_1808,N_1317);
nor U2498 (N_2498,N_1640,N_1345);
nor U2499 (N_2499,N_1152,N_1963);
or U2500 (N_2500,N_1025,N_1045);
xor U2501 (N_2501,N_1679,N_1930);
nand U2502 (N_2502,N_1313,N_1153);
nand U2503 (N_2503,N_1637,N_1457);
nor U2504 (N_2504,N_1485,N_1802);
xnor U2505 (N_2505,N_1007,N_1981);
and U2506 (N_2506,N_1046,N_1431);
or U2507 (N_2507,N_1659,N_1561);
and U2508 (N_2508,N_1097,N_1398);
nand U2509 (N_2509,N_1806,N_1456);
and U2510 (N_2510,N_1240,N_1414);
and U2511 (N_2511,N_1275,N_1711);
and U2512 (N_2512,N_1904,N_1723);
nor U2513 (N_2513,N_1032,N_1135);
and U2514 (N_2514,N_1875,N_1002);
nor U2515 (N_2515,N_1369,N_1570);
nand U2516 (N_2516,N_1083,N_1802);
and U2517 (N_2517,N_1051,N_1243);
nand U2518 (N_2518,N_1217,N_1861);
nand U2519 (N_2519,N_1797,N_1182);
nor U2520 (N_2520,N_1598,N_1785);
or U2521 (N_2521,N_1265,N_1360);
nor U2522 (N_2522,N_1040,N_1238);
or U2523 (N_2523,N_1644,N_1410);
nor U2524 (N_2524,N_1426,N_1952);
nor U2525 (N_2525,N_1416,N_1841);
and U2526 (N_2526,N_1776,N_1998);
xnor U2527 (N_2527,N_1127,N_1148);
nor U2528 (N_2528,N_1373,N_1321);
nor U2529 (N_2529,N_1615,N_1652);
nor U2530 (N_2530,N_1826,N_1761);
xor U2531 (N_2531,N_1399,N_1325);
nand U2532 (N_2532,N_1514,N_1323);
nor U2533 (N_2533,N_1384,N_1300);
or U2534 (N_2534,N_1950,N_1241);
nand U2535 (N_2535,N_1935,N_1570);
or U2536 (N_2536,N_1840,N_1725);
or U2537 (N_2537,N_1445,N_1760);
and U2538 (N_2538,N_1298,N_1295);
or U2539 (N_2539,N_1795,N_1747);
or U2540 (N_2540,N_1456,N_1825);
or U2541 (N_2541,N_1404,N_1303);
and U2542 (N_2542,N_1152,N_1642);
xnor U2543 (N_2543,N_1940,N_1928);
nor U2544 (N_2544,N_1795,N_1567);
and U2545 (N_2545,N_1345,N_1644);
and U2546 (N_2546,N_1823,N_1801);
or U2547 (N_2547,N_1738,N_1821);
and U2548 (N_2548,N_1971,N_1442);
nand U2549 (N_2549,N_1300,N_1301);
nand U2550 (N_2550,N_1312,N_1964);
and U2551 (N_2551,N_1147,N_1108);
nor U2552 (N_2552,N_1242,N_1898);
or U2553 (N_2553,N_1237,N_1584);
and U2554 (N_2554,N_1147,N_1034);
nand U2555 (N_2555,N_1246,N_1463);
nand U2556 (N_2556,N_1390,N_1138);
nand U2557 (N_2557,N_1009,N_1348);
and U2558 (N_2558,N_1018,N_1139);
and U2559 (N_2559,N_1967,N_1101);
nand U2560 (N_2560,N_1078,N_1421);
nand U2561 (N_2561,N_1896,N_1961);
nor U2562 (N_2562,N_1286,N_1858);
and U2563 (N_2563,N_1926,N_1471);
nand U2564 (N_2564,N_1452,N_1787);
and U2565 (N_2565,N_1787,N_1596);
and U2566 (N_2566,N_1455,N_1626);
nor U2567 (N_2567,N_1505,N_1041);
or U2568 (N_2568,N_1826,N_1250);
or U2569 (N_2569,N_1370,N_1789);
nor U2570 (N_2570,N_1400,N_1463);
xnor U2571 (N_2571,N_1742,N_1248);
or U2572 (N_2572,N_1349,N_1854);
nor U2573 (N_2573,N_1234,N_1307);
and U2574 (N_2574,N_1755,N_1404);
or U2575 (N_2575,N_1831,N_1028);
nor U2576 (N_2576,N_1397,N_1422);
nor U2577 (N_2577,N_1573,N_1750);
nand U2578 (N_2578,N_1030,N_1473);
or U2579 (N_2579,N_1914,N_1850);
or U2580 (N_2580,N_1778,N_1185);
nor U2581 (N_2581,N_1230,N_1000);
or U2582 (N_2582,N_1515,N_1660);
or U2583 (N_2583,N_1963,N_1768);
xnor U2584 (N_2584,N_1009,N_1901);
nor U2585 (N_2585,N_1002,N_1364);
and U2586 (N_2586,N_1036,N_1458);
and U2587 (N_2587,N_1930,N_1258);
xor U2588 (N_2588,N_1566,N_1493);
nor U2589 (N_2589,N_1545,N_1016);
xnor U2590 (N_2590,N_1867,N_1469);
nor U2591 (N_2591,N_1994,N_1201);
nor U2592 (N_2592,N_1639,N_1747);
xor U2593 (N_2593,N_1185,N_1328);
xor U2594 (N_2594,N_1421,N_1625);
nand U2595 (N_2595,N_1022,N_1557);
and U2596 (N_2596,N_1405,N_1210);
nand U2597 (N_2597,N_1641,N_1420);
nand U2598 (N_2598,N_1180,N_1964);
or U2599 (N_2599,N_1879,N_1844);
or U2600 (N_2600,N_1522,N_1133);
and U2601 (N_2601,N_1906,N_1373);
or U2602 (N_2602,N_1075,N_1013);
nor U2603 (N_2603,N_1308,N_1244);
nor U2604 (N_2604,N_1624,N_1413);
or U2605 (N_2605,N_1983,N_1743);
nor U2606 (N_2606,N_1005,N_1462);
nor U2607 (N_2607,N_1902,N_1226);
or U2608 (N_2608,N_1874,N_1666);
or U2609 (N_2609,N_1585,N_1215);
or U2610 (N_2610,N_1084,N_1802);
or U2611 (N_2611,N_1848,N_1936);
nor U2612 (N_2612,N_1347,N_1756);
and U2613 (N_2613,N_1412,N_1428);
nand U2614 (N_2614,N_1572,N_1242);
or U2615 (N_2615,N_1505,N_1425);
nand U2616 (N_2616,N_1201,N_1762);
xor U2617 (N_2617,N_1971,N_1640);
nor U2618 (N_2618,N_1937,N_1155);
or U2619 (N_2619,N_1376,N_1803);
nand U2620 (N_2620,N_1175,N_1372);
and U2621 (N_2621,N_1640,N_1125);
nor U2622 (N_2622,N_1843,N_1527);
xor U2623 (N_2623,N_1539,N_1310);
nor U2624 (N_2624,N_1175,N_1551);
nor U2625 (N_2625,N_1790,N_1169);
and U2626 (N_2626,N_1675,N_1955);
or U2627 (N_2627,N_1915,N_1513);
and U2628 (N_2628,N_1755,N_1406);
or U2629 (N_2629,N_1222,N_1710);
nand U2630 (N_2630,N_1969,N_1043);
and U2631 (N_2631,N_1710,N_1800);
or U2632 (N_2632,N_1549,N_1289);
nor U2633 (N_2633,N_1289,N_1728);
nor U2634 (N_2634,N_1463,N_1879);
nor U2635 (N_2635,N_1557,N_1104);
xnor U2636 (N_2636,N_1794,N_1819);
nand U2637 (N_2637,N_1019,N_1280);
and U2638 (N_2638,N_1973,N_1379);
xor U2639 (N_2639,N_1793,N_1554);
or U2640 (N_2640,N_1100,N_1533);
nor U2641 (N_2641,N_1166,N_1666);
and U2642 (N_2642,N_1937,N_1150);
and U2643 (N_2643,N_1358,N_1680);
nand U2644 (N_2644,N_1711,N_1660);
nor U2645 (N_2645,N_1936,N_1460);
nand U2646 (N_2646,N_1907,N_1649);
nand U2647 (N_2647,N_1837,N_1212);
and U2648 (N_2648,N_1577,N_1254);
nand U2649 (N_2649,N_1323,N_1568);
and U2650 (N_2650,N_1134,N_1144);
and U2651 (N_2651,N_1426,N_1231);
nor U2652 (N_2652,N_1622,N_1287);
and U2653 (N_2653,N_1070,N_1909);
nor U2654 (N_2654,N_1264,N_1223);
nor U2655 (N_2655,N_1716,N_1925);
nand U2656 (N_2656,N_1929,N_1370);
nor U2657 (N_2657,N_1393,N_1936);
and U2658 (N_2658,N_1201,N_1462);
nand U2659 (N_2659,N_1079,N_1056);
or U2660 (N_2660,N_1450,N_1870);
nor U2661 (N_2661,N_1024,N_1337);
and U2662 (N_2662,N_1330,N_1572);
and U2663 (N_2663,N_1079,N_1262);
or U2664 (N_2664,N_1236,N_1863);
nor U2665 (N_2665,N_1182,N_1905);
xnor U2666 (N_2666,N_1434,N_1794);
nor U2667 (N_2667,N_1408,N_1285);
xor U2668 (N_2668,N_1209,N_1443);
nand U2669 (N_2669,N_1658,N_1582);
nand U2670 (N_2670,N_1615,N_1846);
nand U2671 (N_2671,N_1631,N_1696);
or U2672 (N_2672,N_1378,N_1132);
or U2673 (N_2673,N_1125,N_1965);
nand U2674 (N_2674,N_1068,N_1399);
nor U2675 (N_2675,N_1585,N_1492);
and U2676 (N_2676,N_1423,N_1891);
nor U2677 (N_2677,N_1384,N_1368);
and U2678 (N_2678,N_1976,N_1530);
or U2679 (N_2679,N_1908,N_1684);
and U2680 (N_2680,N_1548,N_1683);
and U2681 (N_2681,N_1026,N_1957);
nand U2682 (N_2682,N_1286,N_1087);
and U2683 (N_2683,N_1915,N_1151);
nand U2684 (N_2684,N_1691,N_1935);
xor U2685 (N_2685,N_1470,N_1951);
nor U2686 (N_2686,N_1254,N_1268);
and U2687 (N_2687,N_1794,N_1953);
nand U2688 (N_2688,N_1608,N_1366);
nor U2689 (N_2689,N_1065,N_1250);
or U2690 (N_2690,N_1684,N_1623);
nor U2691 (N_2691,N_1589,N_1644);
nor U2692 (N_2692,N_1473,N_1003);
nor U2693 (N_2693,N_1219,N_1816);
nand U2694 (N_2694,N_1925,N_1392);
or U2695 (N_2695,N_1891,N_1197);
nor U2696 (N_2696,N_1642,N_1196);
nand U2697 (N_2697,N_1773,N_1024);
nand U2698 (N_2698,N_1735,N_1868);
and U2699 (N_2699,N_1750,N_1807);
nor U2700 (N_2700,N_1370,N_1705);
and U2701 (N_2701,N_1528,N_1562);
or U2702 (N_2702,N_1164,N_1232);
or U2703 (N_2703,N_1366,N_1445);
nand U2704 (N_2704,N_1389,N_1149);
or U2705 (N_2705,N_1621,N_1346);
nand U2706 (N_2706,N_1210,N_1236);
or U2707 (N_2707,N_1837,N_1924);
xnor U2708 (N_2708,N_1616,N_1395);
xor U2709 (N_2709,N_1006,N_1404);
nand U2710 (N_2710,N_1716,N_1584);
nand U2711 (N_2711,N_1387,N_1893);
nor U2712 (N_2712,N_1164,N_1198);
and U2713 (N_2713,N_1499,N_1698);
and U2714 (N_2714,N_1341,N_1160);
nor U2715 (N_2715,N_1013,N_1973);
nand U2716 (N_2716,N_1598,N_1057);
nor U2717 (N_2717,N_1419,N_1197);
nand U2718 (N_2718,N_1816,N_1370);
xor U2719 (N_2719,N_1613,N_1464);
and U2720 (N_2720,N_1618,N_1081);
nor U2721 (N_2721,N_1502,N_1041);
nor U2722 (N_2722,N_1570,N_1872);
and U2723 (N_2723,N_1092,N_1742);
or U2724 (N_2724,N_1088,N_1537);
nand U2725 (N_2725,N_1476,N_1118);
nand U2726 (N_2726,N_1003,N_1044);
or U2727 (N_2727,N_1683,N_1547);
nor U2728 (N_2728,N_1143,N_1664);
or U2729 (N_2729,N_1985,N_1501);
and U2730 (N_2730,N_1074,N_1309);
nor U2731 (N_2731,N_1664,N_1792);
and U2732 (N_2732,N_1430,N_1837);
nor U2733 (N_2733,N_1928,N_1109);
or U2734 (N_2734,N_1607,N_1267);
nor U2735 (N_2735,N_1092,N_1840);
and U2736 (N_2736,N_1731,N_1879);
nor U2737 (N_2737,N_1686,N_1785);
or U2738 (N_2738,N_1833,N_1509);
or U2739 (N_2739,N_1424,N_1770);
and U2740 (N_2740,N_1484,N_1822);
nor U2741 (N_2741,N_1899,N_1377);
nor U2742 (N_2742,N_1764,N_1023);
nor U2743 (N_2743,N_1681,N_1659);
or U2744 (N_2744,N_1853,N_1617);
and U2745 (N_2745,N_1431,N_1006);
xnor U2746 (N_2746,N_1664,N_1807);
xor U2747 (N_2747,N_1571,N_1875);
and U2748 (N_2748,N_1294,N_1779);
and U2749 (N_2749,N_1092,N_1947);
nand U2750 (N_2750,N_1034,N_1488);
nand U2751 (N_2751,N_1153,N_1913);
and U2752 (N_2752,N_1867,N_1374);
and U2753 (N_2753,N_1385,N_1638);
nand U2754 (N_2754,N_1622,N_1255);
nand U2755 (N_2755,N_1629,N_1850);
nand U2756 (N_2756,N_1874,N_1806);
nor U2757 (N_2757,N_1515,N_1068);
nor U2758 (N_2758,N_1058,N_1338);
or U2759 (N_2759,N_1400,N_1909);
nand U2760 (N_2760,N_1491,N_1346);
or U2761 (N_2761,N_1437,N_1526);
nand U2762 (N_2762,N_1613,N_1799);
nand U2763 (N_2763,N_1429,N_1059);
xnor U2764 (N_2764,N_1101,N_1317);
and U2765 (N_2765,N_1884,N_1038);
xor U2766 (N_2766,N_1153,N_1427);
nand U2767 (N_2767,N_1984,N_1281);
xor U2768 (N_2768,N_1859,N_1456);
and U2769 (N_2769,N_1194,N_1112);
nor U2770 (N_2770,N_1530,N_1352);
or U2771 (N_2771,N_1242,N_1233);
nand U2772 (N_2772,N_1452,N_1542);
nand U2773 (N_2773,N_1168,N_1664);
nor U2774 (N_2774,N_1169,N_1992);
nor U2775 (N_2775,N_1783,N_1105);
nor U2776 (N_2776,N_1414,N_1908);
or U2777 (N_2777,N_1384,N_1759);
or U2778 (N_2778,N_1869,N_1466);
xor U2779 (N_2779,N_1687,N_1970);
and U2780 (N_2780,N_1080,N_1779);
nor U2781 (N_2781,N_1788,N_1738);
nand U2782 (N_2782,N_1705,N_1283);
and U2783 (N_2783,N_1267,N_1822);
and U2784 (N_2784,N_1553,N_1396);
or U2785 (N_2785,N_1835,N_1132);
and U2786 (N_2786,N_1974,N_1823);
nand U2787 (N_2787,N_1614,N_1949);
nor U2788 (N_2788,N_1547,N_1061);
nor U2789 (N_2789,N_1661,N_1295);
nand U2790 (N_2790,N_1324,N_1290);
nand U2791 (N_2791,N_1507,N_1032);
xor U2792 (N_2792,N_1915,N_1479);
nand U2793 (N_2793,N_1227,N_1465);
nor U2794 (N_2794,N_1333,N_1975);
and U2795 (N_2795,N_1235,N_1548);
and U2796 (N_2796,N_1473,N_1072);
and U2797 (N_2797,N_1335,N_1169);
nand U2798 (N_2798,N_1621,N_1143);
or U2799 (N_2799,N_1962,N_1272);
and U2800 (N_2800,N_1972,N_1768);
xnor U2801 (N_2801,N_1409,N_1149);
nand U2802 (N_2802,N_1326,N_1054);
nand U2803 (N_2803,N_1507,N_1002);
or U2804 (N_2804,N_1969,N_1668);
nor U2805 (N_2805,N_1313,N_1857);
xor U2806 (N_2806,N_1290,N_1055);
nor U2807 (N_2807,N_1524,N_1736);
and U2808 (N_2808,N_1496,N_1171);
nor U2809 (N_2809,N_1104,N_1593);
nand U2810 (N_2810,N_1264,N_1494);
and U2811 (N_2811,N_1447,N_1958);
nand U2812 (N_2812,N_1912,N_1118);
nand U2813 (N_2813,N_1812,N_1625);
nand U2814 (N_2814,N_1286,N_1928);
and U2815 (N_2815,N_1454,N_1950);
xor U2816 (N_2816,N_1738,N_1178);
nand U2817 (N_2817,N_1047,N_1349);
or U2818 (N_2818,N_1356,N_1931);
nand U2819 (N_2819,N_1075,N_1170);
and U2820 (N_2820,N_1872,N_1031);
nand U2821 (N_2821,N_1211,N_1328);
nor U2822 (N_2822,N_1174,N_1048);
or U2823 (N_2823,N_1323,N_1171);
nand U2824 (N_2824,N_1711,N_1578);
or U2825 (N_2825,N_1473,N_1646);
or U2826 (N_2826,N_1224,N_1019);
nor U2827 (N_2827,N_1163,N_1186);
and U2828 (N_2828,N_1897,N_1375);
and U2829 (N_2829,N_1740,N_1990);
or U2830 (N_2830,N_1883,N_1713);
nand U2831 (N_2831,N_1423,N_1311);
nor U2832 (N_2832,N_1593,N_1887);
nand U2833 (N_2833,N_1849,N_1597);
nor U2834 (N_2834,N_1341,N_1889);
or U2835 (N_2835,N_1890,N_1023);
nor U2836 (N_2836,N_1526,N_1587);
and U2837 (N_2837,N_1036,N_1709);
nand U2838 (N_2838,N_1348,N_1293);
xor U2839 (N_2839,N_1451,N_1692);
nand U2840 (N_2840,N_1755,N_1676);
or U2841 (N_2841,N_1988,N_1725);
or U2842 (N_2842,N_1481,N_1626);
nand U2843 (N_2843,N_1578,N_1484);
and U2844 (N_2844,N_1245,N_1538);
nand U2845 (N_2845,N_1601,N_1572);
nor U2846 (N_2846,N_1767,N_1819);
nand U2847 (N_2847,N_1354,N_1710);
or U2848 (N_2848,N_1371,N_1663);
nand U2849 (N_2849,N_1264,N_1361);
or U2850 (N_2850,N_1881,N_1567);
nor U2851 (N_2851,N_1093,N_1647);
and U2852 (N_2852,N_1285,N_1375);
or U2853 (N_2853,N_1150,N_1859);
nor U2854 (N_2854,N_1382,N_1363);
and U2855 (N_2855,N_1989,N_1715);
nor U2856 (N_2856,N_1986,N_1779);
or U2857 (N_2857,N_1834,N_1724);
or U2858 (N_2858,N_1637,N_1190);
xor U2859 (N_2859,N_1608,N_1635);
and U2860 (N_2860,N_1543,N_1821);
nor U2861 (N_2861,N_1782,N_1628);
or U2862 (N_2862,N_1352,N_1241);
xor U2863 (N_2863,N_1502,N_1727);
and U2864 (N_2864,N_1753,N_1660);
nor U2865 (N_2865,N_1366,N_1529);
or U2866 (N_2866,N_1667,N_1939);
or U2867 (N_2867,N_1241,N_1516);
and U2868 (N_2868,N_1607,N_1392);
nand U2869 (N_2869,N_1458,N_1125);
nor U2870 (N_2870,N_1987,N_1143);
nand U2871 (N_2871,N_1008,N_1885);
nand U2872 (N_2872,N_1764,N_1283);
or U2873 (N_2873,N_1193,N_1564);
and U2874 (N_2874,N_1508,N_1793);
nor U2875 (N_2875,N_1153,N_1224);
nor U2876 (N_2876,N_1776,N_1693);
nand U2877 (N_2877,N_1034,N_1669);
nor U2878 (N_2878,N_1447,N_1832);
or U2879 (N_2879,N_1103,N_1586);
xor U2880 (N_2880,N_1965,N_1143);
xnor U2881 (N_2881,N_1655,N_1500);
xor U2882 (N_2882,N_1489,N_1039);
nor U2883 (N_2883,N_1970,N_1593);
or U2884 (N_2884,N_1888,N_1175);
xor U2885 (N_2885,N_1716,N_1351);
xor U2886 (N_2886,N_1916,N_1032);
xor U2887 (N_2887,N_1426,N_1795);
or U2888 (N_2888,N_1526,N_1706);
nand U2889 (N_2889,N_1836,N_1986);
and U2890 (N_2890,N_1991,N_1362);
xnor U2891 (N_2891,N_1219,N_1451);
or U2892 (N_2892,N_1650,N_1814);
nor U2893 (N_2893,N_1078,N_1759);
or U2894 (N_2894,N_1450,N_1577);
nand U2895 (N_2895,N_1474,N_1338);
or U2896 (N_2896,N_1319,N_1259);
xor U2897 (N_2897,N_1925,N_1400);
or U2898 (N_2898,N_1070,N_1191);
xor U2899 (N_2899,N_1830,N_1177);
nor U2900 (N_2900,N_1727,N_1025);
or U2901 (N_2901,N_1295,N_1224);
or U2902 (N_2902,N_1534,N_1786);
nand U2903 (N_2903,N_1886,N_1396);
or U2904 (N_2904,N_1731,N_1813);
nand U2905 (N_2905,N_1275,N_1316);
or U2906 (N_2906,N_1708,N_1966);
or U2907 (N_2907,N_1949,N_1507);
xnor U2908 (N_2908,N_1642,N_1629);
nand U2909 (N_2909,N_1506,N_1792);
nand U2910 (N_2910,N_1718,N_1852);
nand U2911 (N_2911,N_1640,N_1204);
nand U2912 (N_2912,N_1007,N_1948);
or U2913 (N_2913,N_1441,N_1717);
xor U2914 (N_2914,N_1579,N_1351);
and U2915 (N_2915,N_1547,N_1492);
and U2916 (N_2916,N_1869,N_1208);
nand U2917 (N_2917,N_1650,N_1522);
or U2918 (N_2918,N_1576,N_1852);
or U2919 (N_2919,N_1175,N_1040);
nor U2920 (N_2920,N_1511,N_1462);
and U2921 (N_2921,N_1815,N_1452);
and U2922 (N_2922,N_1462,N_1109);
nand U2923 (N_2923,N_1521,N_1007);
nand U2924 (N_2924,N_1095,N_1484);
and U2925 (N_2925,N_1899,N_1457);
nand U2926 (N_2926,N_1364,N_1618);
and U2927 (N_2927,N_1628,N_1215);
nor U2928 (N_2928,N_1727,N_1202);
or U2929 (N_2929,N_1945,N_1435);
and U2930 (N_2930,N_1713,N_1225);
nand U2931 (N_2931,N_1752,N_1198);
nor U2932 (N_2932,N_1454,N_1988);
nor U2933 (N_2933,N_1496,N_1629);
nand U2934 (N_2934,N_1334,N_1236);
nor U2935 (N_2935,N_1198,N_1404);
nand U2936 (N_2936,N_1941,N_1464);
or U2937 (N_2937,N_1172,N_1924);
or U2938 (N_2938,N_1093,N_1022);
nor U2939 (N_2939,N_1804,N_1907);
xnor U2940 (N_2940,N_1033,N_1369);
and U2941 (N_2941,N_1271,N_1191);
nand U2942 (N_2942,N_1685,N_1586);
nand U2943 (N_2943,N_1110,N_1214);
and U2944 (N_2944,N_1024,N_1626);
nor U2945 (N_2945,N_1403,N_1813);
nand U2946 (N_2946,N_1409,N_1454);
nor U2947 (N_2947,N_1440,N_1640);
xor U2948 (N_2948,N_1305,N_1766);
nand U2949 (N_2949,N_1306,N_1256);
nand U2950 (N_2950,N_1612,N_1957);
nor U2951 (N_2951,N_1286,N_1380);
or U2952 (N_2952,N_1291,N_1551);
and U2953 (N_2953,N_1190,N_1800);
and U2954 (N_2954,N_1507,N_1851);
or U2955 (N_2955,N_1502,N_1354);
nand U2956 (N_2956,N_1468,N_1371);
and U2957 (N_2957,N_1026,N_1834);
or U2958 (N_2958,N_1533,N_1156);
nor U2959 (N_2959,N_1539,N_1767);
nand U2960 (N_2960,N_1730,N_1025);
or U2961 (N_2961,N_1869,N_1233);
and U2962 (N_2962,N_1361,N_1242);
nor U2963 (N_2963,N_1154,N_1195);
and U2964 (N_2964,N_1287,N_1198);
nand U2965 (N_2965,N_1589,N_1482);
or U2966 (N_2966,N_1000,N_1607);
or U2967 (N_2967,N_1915,N_1709);
and U2968 (N_2968,N_1321,N_1378);
nor U2969 (N_2969,N_1315,N_1760);
or U2970 (N_2970,N_1523,N_1045);
nand U2971 (N_2971,N_1782,N_1745);
nor U2972 (N_2972,N_1520,N_1011);
nand U2973 (N_2973,N_1663,N_1833);
nand U2974 (N_2974,N_1523,N_1478);
nor U2975 (N_2975,N_1237,N_1340);
nor U2976 (N_2976,N_1592,N_1950);
nand U2977 (N_2977,N_1988,N_1993);
nor U2978 (N_2978,N_1905,N_1133);
or U2979 (N_2979,N_1063,N_1274);
and U2980 (N_2980,N_1887,N_1477);
nor U2981 (N_2981,N_1294,N_1874);
xnor U2982 (N_2982,N_1914,N_1691);
nand U2983 (N_2983,N_1789,N_1023);
nand U2984 (N_2984,N_1019,N_1966);
xnor U2985 (N_2985,N_1097,N_1843);
nand U2986 (N_2986,N_1840,N_1800);
and U2987 (N_2987,N_1737,N_1532);
xnor U2988 (N_2988,N_1789,N_1497);
nand U2989 (N_2989,N_1881,N_1775);
nor U2990 (N_2990,N_1935,N_1912);
nand U2991 (N_2991,N_1153,N_1851);
nor U2992 (N_2992,N_1244,N_1674);
and U2993 (N_2993,N_1410,N_1729);
xnor U2994 (N_2994,N_1758,N_1125);
xor U2995 (N_2995,N_1487,N_1468);
nand U2996 (N_2996,N_1855,N_1722);
nand U2997 (N_2997,N_1437,N_1916);
nand U2998 (N_2998,N_1301,N_1553);
nor U2999 (N_2999,N_1929,N_1035);
xor U3000 (N_3000,N_2218,N_2911);
xor U3001 (N_3001,N_2702,N_2582);
nor U3002 (N_3002,N_2438,N_2616);
or U3003 (N_3003,N_2774,N_2772);
nor U3004 (N_3004,N_2231,N_2883);
nand U3005 (N_3005,N_2521,N_2551);
and U3006 (N_3006,N_2448,N_2780);
and U3007 (N_3007,N_2281,N_2352);
or U3008 (N_3008,N_2041,N_2668);
and U3009 (N_3009,N_2920,N_2728);
and U3010 (N_3010,N_2028,N_2569);
and U3011 (N_3011,N_2228,N_2366);
xnor U3012 (N_3012,N_2825,N_2539);
nor U3013 (N_3013,N_2017,N_2674);
and U3014 (N_3014,N_2474,N_2770);
xor U3015 (N_3015,N_2221,N_2845);
nand U3016 (N_3016,N_2736,N_2213);
and U3017 (N_3017,N_2425,N_2981);
and U3018 (N_3018,N_2319,N_2758);
or U3019 (N_3019,N_2846,N_2656);
and U3020 (N_3020,N_2907,N_2421);
xnor U3021 (N_3021,N_2235,N_2408);
nand U3022 (N_3022,N_2983,N_2904);
nand U3023 (N_3023,N_2909,N_2196);
xnor U3024 (N_3024,N_2641,N_2267);
xor U3025 (N_3025,N_2717,N_2662);
and U3026 (N_3026,N_2891,N_2445);
xnor U3027 (N_3027,N_2858,N_2234);
xnor U3028 (N_3028,N_2066,N_2779);
or U3029 (N_3029,N_2999,N_2478);
nand U3030 (N_3030,N_2225,N_2581);
nand U3031 (N_3031,N_2878,N_2093);
or U3032 (N_3032,N_2986,N_2627);
nand U3033 (N_3033,N_2354,N_2670);
nand U3034 (N_3034,N_2713,N_2377);
nor U3035 (N_3035,N_2601,N_2476);
nor U3036 (N_3036,N_2716,N_2944);
nand U3037 (N_3037,N_2503,N_2977);
nor U3038 (N_3038,N_2995,N_2519);
nand U3039 (N_3039,N_2921,N_2056);
or U3040 (N_3040,N_2803,N_2444);
or U3041 (N_3041,N_2119,N_2880);
nand U3042 (N_3042,N_2558,N_2651);
nor U3043 (N_3043,N_2429,N_2250);
nand U3044 (N_3044,N_2795,N_2389);
or U3045 (N_3045,N_2181,N_2632);
or U3046 (N_3046,N_2874,N_2039);
and U3047 (N_3047,N_2021,N_2379);
nor U3048 (N_3048,N_2916,N_2435);
and U3049 (N_3049,N_2918,N_2775);
and U3050 (N_3050,N_2208,N_2787);
xor U3051 (N_3051,N_2900,N_2256);
and U3052 (N_3052,N_2295,N_2722);
and U3053 (N_3053,N_2672,N_2811);
or U3054 (N_3054,N_2226,N_2929);
nand U3055 (N_3055,N_2069,N_2763);
nor U3056 (N_3056,N_2494,N_2561);
and U3057 (N_3057,N_2574,N_2404);
nand U3058 (N_3058,N_2931,N_2720);
and U3059 (N_3059,N_2107,N_2524);
xor U3060 (N_3060,N_2784,N_2859);
nand U3061 (N_3061,N_2993,N_2685);
nor U3062 (N_3062,N_2480,N_2358);
and U3063 (N_3063,N_2618,N_2252);
nand U3064 (N_3064,N_2294,N_2441);
nand U3065 (N_3065,N_2351,N_2495);
or U3066 (N_3066,N_2333,N_2417);
nand U3067 (N_3067,N_2792,N_2082);
nor U3068 (N_3068,N_2614,N_2870);
xnor U3069 (N_3069,N_2469,N_2896);
xor U3070 (N_3070,N_2839,N_2262);
and U3071 (N_3071,N_2933,N_2481);
or U3072 (N_3072,N_2095,N_2089);
nand U3073 (N_3073,N_2871,N_2800);
or U3074 (N_3074,N_2482,N_2777);
nor U3075 (N_3075,N_2694,N_2517);
nand U3076 (N_3076,N_2399,N_2598);
xnor U3077 (N_3077,N_2431,N_2301);
xnor U3078 (N_3078,N_2953,N_2141);
xnor U3079 (N_3079,N_2423,N_2745);
xor U3080 (N_3080,N_2375,N_2443);
and U3081 (N_3081,N_2186,N_2655);
nor U3082 (N_3082,N_2688,N_2278);
nor U3083 (N_3083,N_2996,N_2647);
nor U3084 (N_3084,N_2321,N_2285);
nand U3085 (N_3085,N_2762,N_2111);
nand U3086 (N_3086,N_2068,N_2096);
nand U3087 (N_3087,N_2110,N_2755);
or U3088 (N_3088,N_2144,N_2652);
and U3089 (N_3089,N_2862,N_2338);
nor U3090 (N_3090,N_2034,N_2304);
and U3091 (N_3091,N_2092,N_2214);
xnor U3092 (N_3092,N_2698,N_2356);
and U3093 (N_3093,N_2789,N_2552);
nand U3094 (N_3094,N_2057,N_2229);
or U3095 (N_3095,N_2768,N_2619);
or U3096 (N_3096,N_2691,N_2902);
or U3097 (N_3097,N_2557,N_2406);
nor U3098 (N_3098,N_2177,N_2135);
xnor U3099 (N_3099,N_2030,N_2157);
nor U3100 (N_3100,N_2822,N_2254);
or U3101 (N_3101,N_2705,N_2217);
or U3102 (N_3102,N_2283,N_2837);
nor U3103 (N_3103,N_2393,N_2513);
or U3104 (N_3104,N_2675,N_2633);
and U3105 (N_3105,N_2543,N_2807);
nand U3106 (N_3106,N_2426,N_2689);
nand U3107 (N_3107,N_2820,N_2697);
nand U3108 (N_3108,N_2219,N_2279);
nor U3109 (N_3109,N_2361,N_2611);
nor U3110 (N_3110,N_2451,N_2010);
nand U3111 (N_3111,N_2612,N_2345);
or U3112 (N_3112,N_2156,N_2653);
nor U3113 (N_3113,N_2459,N_2497);
and U3114 (N_3114,N_2105,N_2609);
xnor U3115 (N_3115,N_2367,N_2369);
nand U3116 (N_3116,N_2062,N_2123);
and U3117 (N_3117,N_2868,N_2411);
nand U3118 (N_3118,N_2980,N_2751);
and U3119 (N_3119,N_2757,N_2353);
xnor U3120 (N_3120,N_2038,N_2201);
and U3121 (N_3121,N_2037,N_2788);
and U3122 (N_3122,N_2286,N_2915);
nand U3123 (N_3123,N_2244,N_2805);
nor U3124 (N_3124,N_2565,N_2658);
nor U3125 (N_3125,N_2264,N_2885);
or U3126 (N_3126,N_2313,N_2564);
xnor U3127 (N_3127,N_2525,N_2567);
and U3128 (N_3128,N_2850,N_2372);
or U3129 (N_3129,N_2945,N_2311);
nand U3130 (N_3130,N_2085,N_2173);
and U3131 (N_3131,N_2450,N_2280);
and U3132 (N_3132,N_2851,N_2326);
nor U3133 (N_3133,N_2959,N_2391);
nor U3134 (N_3134,N_2491,N_2289);
and U3135 (N_3135,N_2018,N_2116);
xor U3136 (N_3136,N_2591,N_2292);
and U3137 (N_3137,N_2490,N_2606);
nor U3138 (N_3138,N_2288,N_2306);
nor U3139 (N_3139,N_2091,N_2161);
nand U3140 (N_3140,N_2325,N_2479);
xnor U3141 (N_3141,N_2276,N_2886);
nor U3142 (N_3142,N_2468,N_2955);
and U3143 (N_3143,N_2312,N_2409);
or U3144 (N_3144,N_2102,N_2739);
nor U3145 (N_3145,N_2334,N_2101);
or U3146 (N_3146,N_2518,N_2305);
or U3147 (N_3147,N_2589,N_2346);
or U3148 (N_3148,N_2374,N_2938);
nor U3149 (N_3149,N_2984,N_2950);
and U3150 (N_3150,N_2693,N_2013);
xor U3151 (N_3151,N_2852,N_2455);
and U3152 (N_3152,N_2322,N_2873);
or U3153 (N_3153,N_2032,N_2872);
and U3154 (N_3154,N_2195,N_2405);
or U3155 (N_3155,N_2324,N_2723);
nor U3156 (N_3156,N_2982,N_2071);
nand U3157 (N_3157,N_2025,N_2124);
nor U3158 (N_3158,N_2022,N_2638);
or U3159 (N_3159,N_2064,N_2639);
nor U3160 (N_3160,N_2163,N_2621);
nand U3161 (N_3161,N_2882,N_2164);
or U3162 (N_3162,N_2063,N_2155);
or U3163 (N_3163,N_2625,N_2546);
xnor U3164 (N_3164,N_2407,N_2854);
or U3165 (N_3165,N_2470,N_2145);
nand U3166 (N_3166,N_2576,N_2707);
nand U3167 (N_3167,N_2714,N_2336);
nand U3168 (N_3168,N_2258,N_2230);
and U3169 (N_3169,N_2923,N_2106);
and U3170 (N_3170,N_2903,N_2542);
or U3171 (N_3171,N_2452,N_2307);
nor U3172 (N_3172,N_2473,N_2892);
or U3173 (N_3173,N_2579,N_2094);
and U3174 (N_3174,N_2170,N_2831);
or U3175 (N_3175,N_2840,N_2128);
nand U3176 (N_3176,N_2183,N_2791);
xor U3177 (N_3177,N_2097,N_2269);
nor U3178 (N_3178,N_2988,N_2447);
nand U3179 (N_3179,N_2765,N_2752);
nor U3180 (N_3180,N_2149,N_2548);
or U3181 (N_3181,N_2493,N_2860);
nand U3182 (N_3182,N_2750,N_2783);
and U3183 (N_3183,N_2088,N_2340);
nor U3184 (N_3184,N_2948,N_2457);
or U3185 (N_3185,N_2573,N_2744);
or U3186 (N_3186,N_2936,N_2570);
and U3187 (N_3187,N_2659,N_2316);
nand U3188 (N_3188,N_2526,N_2898);
or U3189 (N_3189,N_2175,N_2463);
nand U3190 (N_3190,N_2673,N_2166);
nand U3191 (N_3191,N_2176,N_2547);
xor U3192 (N_3192,N_2575,N_2913);
and U3193 (N_3193,N_2109,N_2814);
xnor U3194 (N_3194,N_2512,N_2958);
nand U3195 (N_3195,N_2593,N_2174);
nand U3196 (N_3196,N_2150,N_2967);
or U3197 (N_3197,N_2472,N_2342);
nor U3198 (N_3198,N_2863,N_2502);
xnor U3199 (N_3199,N_2520,N_2782);
nor U3200 (N_3200,N_2427,N_2626);
xnor U3201 (N_3201,N_2937,N_2255);
nand U3202 (N_3202,N_2696,N_2748);
nand U3203 (N_3203,N_2889,N_2905);
nand U3204 (N_3204,N_2630,N_2687);
and U3205 (N_3205,N_2818,N_2401);
and U3206 (N_3206,N_2162,N_2646);
xor U3207 (N_3207,N_2680,N_2592);
or U3208 (N_3208,N_2615,N_2853);
nand U3209 (N_3209,N_2754,N_2764);
or U3210 (N_3210,N_2099,N_2634);
nor U3211 (N_3211,N_2436,N_2273);
nand U3212 (N_3212,N_2587,N_2500);
or U3213 (N_3213,N_2243,N_2152);
xor U3214 (N_3214,N_2726,N_2585);
and U3215 (N_3215,N_2384,N_2098);
or U3216 (N_3216,N_2743,N_2053);
or U3217 (N_3217,N_2897,N_2260);
or U3218 (N_3218,N_2888,N_2138);
nor U3219 (N_3219,N_2877,N_2079);
or U3220 (N_3220,N_2833,N_2296);
nor U3221 (N_3221,N_2461,N_2908);
or U3222 (N_3222,N_2499,N_2328);
nor U3223 (N_3223,N_2060,N_2061);
nand U3224 (N_3224,N_2810,N_2594);
or U3225 (N_3225,N_2940,N_2396);
and U3226 (N_3226,N_2767,N_2506);
nand U3227 (N_3227,N_2899,N_2185);
nor U3228 (N_3228,N_2972,N_2537);
nor U3229 (N_3229,N_2159,N_2978);
and U3230 (N_3230,N_2036,N_2168);
nand U3231 (N_3231,N_2604,N_2681);
nand U3232 (N_3232,N_2114,N_2003);
or U3233 (N_3233,N_2416,N_2083);
and U3234 (N_3234,N_2151,N_2773);
nand U3235 (N_3235,N_2016,N_2682);
or U3236 (N_3236,N_2419,N_2951);
and U3237 (N_3237,N_2362,N_2265);
nor U3238 (N_3238,N_2290,N_2866);
nor U3239 (N_3239,N_2224,N_2690);
or U3240 (N_3240,N_2090,N_2303);
xnor U3241 (N_3241,N_2695,N_2965);
nand U3242 (N_3242,N_2483,N_2420);
nor U3243 (N_3243,N_2347,N_2317);
and U3244 (N_3244,N_2132,N_2040);
and U3245 (N_3245,N_2654,N_2386);
and U3246 (N_3246,N_2556,N_2033);
nor U3247 (N_3247,N_2934,N_2006);
and U3248 (N_3248,N_2191,N_2394);
nand U3249 (N_3249,N_2719,N_2535);
nor U3250 (N_3250,N_2360,N_2975);
nand U3251 (N_3251,N_2650,N_2223);
and U3252 (N_3252,N_2657,N_2742);
xor U3253 (N_3253,N_2165,N_2732);
nor U3254 (N_3254,N_2320,N_2489);
nor U3255 (N_3255,N_2332,N_2761);
and U3256 (N_3256,N_2644,N_2287);
nand U3257 (N_3257,N_2821,N_2678);
and U3258 (N_3258,N_2180,N_2440);
nor U3259 (N_3259,N_2080,N_2608);
or U3260 (N_3260,N_2596,N_2930);
nand U3261 (N_3261,N_2207,N_2239);
xnor U3262 (N_3262,N_2628,N_2706);
nor U3263 (N_3263,N_2359,N_2241);
and U3264 (N_3264,N_2998,N_2527);
nand U3265 (N_3265,N_2475,N_2487);
nand U3266 (N_3266,N_2893,N_2012);
nand U3267 (N_3267,N_2437,N_2179);
and U3268 (N_3268,N_2636,N_2834);
nor U3269 (N_3269,N_2949,N_2737);
nor U3270 (N_3270,N_2600,N_2631);
and U3271 (N_3271,N_2498,N_2050);
xnor U3272 (N_3272,N_2073,N_2738);
and U3273 (N_3273,N_2588,N_2051);
nor U3274 (N_3274,N_2566,N_2549);
nor U3275 (N_3275,N_2912,N_2890);
and U3276 (N_3276,N_2065,N_2014);
or U3277 (N_3277,N_2291,N_2418);
and U3278 (N_3278,N_2568,N_2414);
or U3279 (N_3279,N_2024,N_2275);
xnor U3280 (N_3280,N_2661,N_2120);
nand U3281 (N_3281,N_2617,N_2086);
and U3282 (N_3282,N_2246,N_2357);
nand U3283 (N_3283,N_2861,N_2058);
or U3284 (N_3284,N_2381,N_2793);
nand U3285 (N_3285,N_2122,N_2067);
nand U3286 (N_3286,N_2153,N_2836);
or U3287 (N_3287,N_2563,N_2299);
nand U3288 (N_3288,N_2209,N_2649);
or U3289 (N_3289,N_2968,N_2160);
xor U3290 (N_3290,N_2530,N_2486);
or U3291 (N_3291,N_2108,N_2462);
nand U3292 (N_3292,N_2348,N_2648);
xor U3293 (N_3293,N_2976,N_2597);
and U3294 (N_3294,N_2496,N_2453);
xnor U3295 (N_3295,N_2365,N_2876);
nand U3296 (N_3296,N_2130,N_2842);
nor U3297 (N_3297,N_2973,N_2613);
and U3298 (N_3298,N_2009,N_2204);
nand U3299 (N_3299,N_2142,N_2640);
nor U3300 (N_3300,N_2799,N_2044);
or U3301 (N_3301,N_2879,N_2623);
and U3302 (N_3302,N_2828,N_2727);
xnor U3303 (N_3303,N_2906,N_2919);
or U3304 (N_3304,N_2449,N_2766);
or U3305 (N_3305,N_2855,N_2865);
or U3306 (N_3306,N_2749,N_2074);
nand U3307 (N_3307,N_2622,N_2113);
or U3308 (N_3308,N_2522,N_2881);
xor U3309 (N_3309,N_2403,N_2712);
nor U3310 (N_3310,N_2684,N_2677);
and U3311 (N_3311,N_2424,N_2927);
and U3312 (N_3312,N_2578,N_2263);
nor U3313 (N_3313,N_2961,N_2344);
xnor U3314 (N_3314,N_2724,N_2599);
or U3315 (N_3315,N_2711,N_2665);
and U3316 (N_3316,N_2055,N_2533);
nor U3317 (N_3317,N_2422,N_2802);
or U3318 (N_3318,N_2309,N_2211);
nor U3319 (N_3319,N_2456,N_2382);
nand U3320 (N_3320,N_2809,N_2154);
xor U3321 (N_3321,N_2314,N_2070);
nor U3322 (N_3322,N_2330,N_2121);
or U3323 (N_3323,N_2428,N_2029);
or U3324 (N_3324,N_2383,N_2869);
or U3325 (N_3325,N_2355,N_2964);
nor U3326 (N_3326,N_2001,N_2284);
xor U3327 (N_3327,N_2077,N_2501);
or U3328 (N_3328,N_2140,N_2703);
nor U3329 (N_3329,N_2718,N_2005);
xnor U3330 (N_3330,N_2942,N_2610);
and U3331 (N_3331,N_2508,N_2467);
xnor U3332 (N_3332,N_2115,N_2242);
or U3333 (N_3333,N_2580,N_2760);
xor U3334 (N_3334,N_2023,N_2676);
or U3335 (N_3335,N_2194,N_2190);
and U3336 (N_3336,N_2434,N_2266);
nand U3337 (N_3337,N_2376,N_2158);
nor U3338 (N_3338,N_2746,N_2371);
or U3339 (N_3339,N_2020,N_2261);
or U3340 (N_3340,N_2710,N_2963);
xor U3341 (N_3341,N_2171,N_2385);
nand U3342 (N_3342,N_2507,N_2637);
and U3343 (N_3343,N_2052,N_2084);
nor U3344 (N_3344,N_2343,N_2560);
or U3345 (N_3345,N_2054,N_2960);
or U3346 (N_3346,N_2031,N_2388);
or U3347 (N_3347,N_2555,N_2813);
xnor U3348 (N_3348,N_2935,N_2740);
or U3349 (N_3349,N_2943,N_2043);
nand U3350 (N_3350,N_2642,N_2620);
and U3351 (N_3351,N_2167,N_2924);
and U3352 (N_3352,N_2484,N_2117);
and U3353 (N_3353,N_2583,N_2026);
nand U3354 (N_3354,N_2753,N_2205);
nand U3355 (N_3355,N_2643,N_2554);
or U3356 (N_3356,N_2395,N_2538);
or U3357 (N_3357,N_2731,N_2794);
and U3358 (N_3358,N_2756,N_2477);
or U3359 (N_3359,N_2917,N_2954);
or U3360 (N_3360,N_2368,N_2605);
nor U3361 (N_3361,N_2991,N_2928);
or U3362 (N_3362,N_2076,N_2541);
or U3363 (N_3363,N_2460,N_2635);
nor U3364 (N_3364,N_2531,N_2838);
nand U3365 (N_3365,N_2433,N_2466);
and U3366 (N_3366,N_2914,N_2143);
and U3367 (N_3367,N_2699,N_2562);
and U3368 (N_3368,N_2227,N_2210);
nand U3369 (N_3369,N_2843,N_2078);
nand U3370 (N_3370,N_2990,N_2222);
or U3371 (N_3371,N_2131,N_2492);
nor U3372 (N_3372,N_2969,N_2237);
nor U3373 (N_3373,N_2559,N_2701);
nand U3374 (N_3374,N_2832,N_2590);
nor U3375 (N_3375,N_2932,N_2830);
and U3376 (N_3376,N_2941,N_2553);
or U3377 (N_3377,N_2586,N_2059);
nand U3378 (N_3378,N_2137,N_2087);
nand U3379 (N_3379,N_2259,N_2187);
nand U3380 (N_3380,N_2532,N_2747);
nor U3381 (N_3381,N_2962,N_2994);
nor U3382 (N_3382,N_2721,N_2816);
nor U3383 (N_3383,N_2798,N_2268);
and U3384 (N_3384,N_2819,N_2516);
nand U3385 (N_3385,N_2257,N_2136);
nor U3386 (N_3386,N_2300,N_2700);
and U3387 (N_3387,N_2759,N_2000);
nand U3388 (N_3388,N_2215,N_2823);
xor U3389 (N_3389,N_2400,N_2146);
or U3390 (N_3390,N_2629,N_2019);
or U3391 (N_3391,N_2464,N_2220);
nor U3392 (N_3392,N_2008,N_2806);
or U3393 (N_3393,N_2997,N_2804);
or U3394 (N_3394,N_2189,N_2236);
xor U3395 (N_3395,N_2572,N_2193);
nor U3396 (N_3396,N_2178,N_2182);
or U3397 (N_3397,N_2926,N_2895);
and U3398 (N_3398,N_2971,N_2318);
and U3399 (N_3399,N_2692,N_2835);
or U3400 (N_3400,N_2607,N_2827);
xnor U3401 (N_3401,N_2946,N_2378);
nor U3402 (N_3402,N_2169,N_2769);
xnor U3403 (N_3403,N_2528,N_2081);
nand U3404 (N_3404,N_2577,N_2042);
or U3405 (N_3405,N_2412,N_2776);
nor U3406 (N_3406,N_2282,N_2002);
nand U3407 (N_3407,N_2432,N_2824);
or U3408 (N_3408,N_2202,N_2349);
and U3409 (N_3409,N_2203,N_2826);
or U3410 (N_3410,N_2200,N_2272);
nor U3411 (N_3411,N_2540,N_2233);
xor U3412 (N_3412,N_2245,N_2595);
or U3413 (N_3413,N_2901,N_2939);
or U3414 (N_3414,N_2232,N_2645);
and U3415 (N_3415,N_2212,N_2442);
nand U3416 (N_3416,N_2602,N_2571);
nand U3417 (N_3417,N_2817,N_2544);
nand U3418 (N_3418,N_2867,N_2801);
nor U3419 (N_3419,N_2534,N_2126);
nor U3420 (N_3420,N_2771,N_2004);
xnor U3421 (N_3421,N_2987,N_2331);
or U3422 (N_3422,N_2297,N_2184);
and U3423 (N_3423,N_2249,N_2125);
nand U3424 (N_3424,N_2100,N_2327);
or U3425 (N_3425,N_2989,N_2709);
or U3426 (N_3426,N_2337,N_2778);
or U3427 (N_3427,N_2216,N_2302);
nor U3428 (N_3428,N_2104,N_2271);
and U3429 (N_3429,N_2148,N_2584);
and U3430 (N_3430,N_2251,N_2274);
or U3431 (N_3431,N_2894,N_2139);
and U3432 (N_3432,N_2849,N_2387);
and U3433 (N_3433,N_2035,N_2733);
and U3434 (N_3434,N_2240,N_2298);
xnor U3435 (N_3435,N_2875,N_2198);
or U3436 (N_3436,N_2514,N_2841);
nor U3437 (N_3437,N_2127,N_2974);
nor U3438 (N_3438,N_2708,N_2458);
nand U3439 (N_3439,N_2172,N_2488);
nand U3440 (N_3440,N_2277,N_2015);
or U3441 (N_3441,N_2329,N_2884);
nor U3442 (N_3442,N_2529,N_2603);
nand U3443 (N_3443,N_2679,N_2666);
nand U3444 (N_3444,N_2363,N_2683);
and U3445 (N_3445,N_2504,N_2545);
nand U3446 (N_3446,N_2864,N_2446);
and U3447 (N_3447,N_2027,N_2047);
nand U3448 (N_3448,N_2729,N_2966);
or U3449 (N_3449,N_2270,N_2247);
xor U3450 (N_3450,N_2844,N_2671);
xnor U3451 (N_3451,N_2007,N_2075);
or U3452 (N_3452,N_2373,N_2197);
and U3453 (N_3453,N_2970,N_2796);
or U3454 (N_3454,N_2660,N_2812);
nand U3455 (N_3455,N_2624,N_2370);
nor U3456 (N_3456,N_2439,N_2103);
or U3457 (N_3457,N_2011,N_2471);
nand U3458 (N_3458,N_2515,N_2686);
nand U3459 (N_3459,N_2397,N_2730);
nor U3460 (N_3460,N_2815,N_2856);
nor U3461 (N_3461,N_2663,N_2922);
nor U3462 (N_3462,N_2715,N_2293);
and U3463 (N_3463,N_2133,N_2315);
and U3464 (N_3464,N_2430,N_2308);
nand U3465 (N_3465,N_2048,N_2335);
or U3466 (N_3466,N_2410,N_2992);
nor U3467 (N_3467,N_2956,N_2485);
or U3468 (N_3468,N_2129,N_2248);
or U3469 (N_3469,N_2413,N_2704);
nand U3470 (N_3470,N_2049,N_2511);
nor U3471 (N_3471,N_2785,N_2797);
or U3472 (N_3472,N_2238,N_2781);
nor U3473 (N_3473,N_2741,N_2323);
or U3474 (N_3474,N_2510,N_2536);
and U3475 (N_3475,N_2310,N_2725);
nor U3476 (N_3476,N_2147,N_2887);
nor U3477 (N_3477,N_2947,N_2509);
and U3478 (N_3478,N_2118,N_2952);
nor U3479 (N_3479,N_2364,N_2134);
nor U3480 (N_3480,N_2985,N_2790);
and U3481 (N_3481,N_2523,N_2341);
nor U3482 (N_3482,N_2398,N_2925);
nor U3483 (N_3483,N_2669,N_2206);
nand U3484 (N_3484,N_2188,N_2112);
xor U3485 (N_3485,N_2192,N_2350);
and U3486 (N_3486,N_2847,N_2808);
and U3487 (N_3487,N_2199,N_2550);
nand U3488 (N_3488,N_2045,N_2390);
or U3489 (N_3489,N_2857,N_2465);
or U3490 (N_3490,N_2253,N_2786);
or U3491 (N_3491,N_2667,N_2664);
nor U3492 (N_3492,N_2957,N_2339);
and U3493 (N_3493,N_2402,N_2072);
xnor U3494 (N_3494,N_2046,N_2454);
nand U3495 (N_3495,N_2415,N_2979);
and U3496 (N_3496,N_2829,N_2380);
xor U3497 (N_3497,N_2392,N_2735);
and U3498 (N_3498,N_2848,N_2505);
and U3499 (N_3499,N_2910,N_2734);
nand U3500 (N_3500,N_2497,N_2472);
or U3501 (N_3501,N_2114,N_2426);
nor U3502 (N_3502,N_2972,N_2685);
and U3503 (N_3503,N_2838,N_2839);
or U3504 (N_3504,N_2828,N_2665);
nor U3505 (N_3505,N_2967,N_2156);
nand U3506 (N_3506,N_2385,N_2803);
or U3507 (N_3507,N_2405,N_2499);
nor U3508 (N_3508,N_2051,N_2758);
or U3509 (N_3509,N_2400,N_2920);
or U3510 (N_3510,N_2323,N_2017);
nand U3511 (N_3511,N_2926,N_2993);
nand U3512 (N_3512,N_2154,N_2250);
nor U3513 (N_3513,N_2767,N_2052);
xor U3514 (N_3514,N_2641,N_2790);
nor U3515 (N_3515,N_2591,N_2413);
and U3516 (N_3516,N_2815,N_2983);
xor U3517 (N_3517,N_2379,N_2403);
or U3518 (N_3518,N_2216,N_2661);
nor U3519 (N_3519,N_2833,N_2560);
nor U3520 (N_3520,N_2425,N_2451);
nand U3521 (N_3521,N_2245,N_2395);
or U3522 (N_3522,N_2357,N_2313);
nor U3523 (N_3523,N_2795,N_2899);
or U3524 (N_3524,N_2114,N_2505);
nor U3525 (N_3525,N_2383,N_2419);
nand U3526 (N_3526,N_2489,N_2336);
and U3527 (N_3527,N_2063,N_2271);
or U3528 (N_3528,N_2881,N_2887);
or U3529 (N_3529,N_2229,N_2567);
or U3530 (N_3530,N_2231,N_2548);
nand U3531 (N_3531,N_2428,N_2839);
nand U3532 (N_3532,N_2598,N_2712);
or U3533 (N_3533,N_2487,N_2087);
nor U3534 (N_3534,N_2578,N_2854);
nor U3535 (N_3535,N_2464,N_2086);
or U3536 (N_3536,N_2727,N_2964);
or U3537 (N_3537,N_2648,N_2554);
or U3538 (N_3538,N_2578,N_2839);
or U3539 (N_3539,N_2657,N_2514);
nand U3540 (N_3540,N_2297,N_2698);
and U3541 (N_3541,N_2882,N_2903);
xnor U3542 (N_3542,N_2723,N_2433);
nor U3543 (N_3543,N_2285,N_2585);
xor U3544 (N_3544,N_2705,N_2915);
nand U3545 (N_3545,N_2042,N_2346);
nor U3546 (N_3546,N_2020,N_2199);
xnor U3547 (N_3547,N_2444,N_2437);
or U3548 (N_3548,N_2749,N_2050);
or U3549 (N_3549,N_2630,N_2792);
and U3550 (N_3550,N_2243,N_2674);
xnor U3551 (N_3551,N_2491,N_2076);
nand U3552 (N_3552,N_2513,N_2669);
and U3553 (N_3553,N_2001,N_2596);
nor U3554 (N_3554,N_2869,N_2165);
nor U3555 (N_3555,N_2645,N_2896);
nor U3556 (N_3556,N_2474,N_2486);
xor U3557 (N_3557,N_2943,N_2463);
nand U3558 (N_3558,N_2118,N_2551);
or U3559 (N_3559,N_2389,N_2846);
xnor U3560 (N_3560,N_2135,N_2484);
nand U3561 (N_3561,N_2488,N_2566);
and U3562 (N_3562,N_2303,N_2392);
and U3563 (N_3563,N_2161,N_2956);
nor U3564 (N_3564,N_2558,N_2970);
xor U3565 (N_3565,N_2749,N_2363);
nor U3566 (N_3566,N_2101,N_2799);
nand U3567 (N_3567,N_2193,N_2780);
nand U3568 (N_3568,N_2546,N_2212);
or U3569 (N_3569,N_2857,N_2493);
and U3570 (N_3570,N_2791,N_2830);
and U3571 (N_3571,N_2729,N_2321);
and U3572 (N_3572,N_2728,N_2141);
or U3573 (N_3573,N_2103,N_2245);
nand U3574 (N_3574,N_2117,N_2824);
nor U3575 (N_3575,N_2256,N_2933);
nor U3576 (N_3576,N_2121,N_2775);
and U3577 (N_3577,N_2695,N_2622);
xnor U3578 (N_3578,N_2286,N_2933);
and U3579 (N_3579,N_2259,N_2285);
nor U3580 (N_3580,N_2979,N_2756);
nor U3581 (N_3581,N_2140,N_2019);
and U3582 (N_3582,N_2645,N_2878);
xnor U3583 (N_3583,N_2827,N_2190);
or U3584 (N_3584,N_2075,N_2428);
and U3585 (N_3585,N_2295,N_2786);
or U3586 (N_3586,N_2086,N_2085);
nor U3587 (N_3587,N_2923,N_2919);
or U3588 (N_3588,N_2372,N_2977);
and U3589 (N_3589,N_2255,N_2768);
and U3590 (N_3590,N_2420,N_2769);
nand U3591 (N_3591,N_2534,N_2012);
or U3592 (N_3592,N_2185,N_2861);
and U3593 (N_3593,N_2599,N_2343);
or U3594 (N_3594,N_2281,N_2824);
nor U3595 (N_3595,N_2458,N_2736);
or U3596 (N_3596,N_2316,N_2873);
or U3597 (N_3597,N_2092,N_2754);
nor U3598 (N_3598,N_2368,N_2728);
or U3599 (N_3599,N_2563,N_2431);
nand U3600 (N_3600,N_2398,N_2779);
or U3601 (N_3601,N_2192,N_2748);
and U3602 (N_3602,N_2581,N_2815);
xnor U3603 (N_3603,N_2623,N_2114);
nand U3604 (N_3604,N_2866,N_2422);
and U3605 (N_3605,N_2152,N_2722);
nand U3606 (N_3606,N_2352,N_2850);
or U3607 (N_3607,N_2632,N_2459);
xor U3608 (N_3608,N_2631,N_2259);
and U3609 (N_3609,N_2352,N_2108);
nor U3610 (N_3610,N_2140,N_2704);
or U3611 (N_3611,N_2078,N_2423);
or U3612 (N_3612,N_2196,N_2790);
nand U3613 (N_3613,N_2564,N_2676);
nor U3614 (N_3614,N_2883,N_2454);
nor U3615 (N_3615,N_2742,N_2361);
and U3616 (N_3616,N_2305,N_2839);
nand U3617 (N_3617,N_2895,N_2020);
xor U3618 (N_3618,N_2118,N_2774);
nor U3619 (N_3619,N_2037,N_2314);
nor U3620 (N_3620,N_2837,N_2895);
and U3621 (N_3621,N_2860,N_2151);
or U3622 (N_3622,N_2330,N_2819);
or U3623 (N_3623,N_2764,N_2430);
and U3624 (N_3624,N_2643,N_2927);
nor U3625 (N_3625,N_2903,N_2006);
nand U3626 (N_3626,N_2062,N_2167);
nand U3627 (N_3627,N_2595,N_2501);
xnor U3628 (N_3628,N_2934,N_2169);
nand U3629 (N_3629,N_2059,N_2827);
nor U3630 (N_3630,N_2092,N_2256);
nor U3631 (N_3631,N_2891,N_2067);
nand U3632 (N_3632,N_2972,N_2057);
xor U3633 (N_3633,N_2601,N_2459);
xor U3634 (N_3634,N_2369,N_2791);
xnor U3635 (N_3635,N_2229,N_2115);
nor U3636 (N_3636,N_2413,N_2120);
or U3637 (N_3637,N_2653,N_2027);
xnor U3638 (N_3638,N_2216,N_2141);
nor U3639 (N_3639,N_2385,N_2010);
xor U3640 (N_3640,N_2953,N_2864);
xnor U3641 (N_3641,N_2379,N_2979);
and U3642 (N_3642,N_2343,N_2939);
xor U3643 (N_3643,N_2462,N_2861);
nor U3644 (N_3644,N_2728,N_2887);
and U3645 (N_3645,N_2053,N_2559);
nor U3646 (N_3646,N_2724,N_2631);
nor U3647 (N_3647,N_2921,N_2055);
nor U3648 (N_3648,N_2264,N_2853);
or U3649 (N_3649,N_2632,N_2801);
or U3650 (N_3650,N_2213,N_2445);
and U3651 (N_3651,N_2030,N_2323);
nor U3652 (N_3652,N_2418,N_2687);
nand U3653 (N_3653,N_2575,N_2674);
nand U3654 (N_3654,N_2529,N_2744);
and U3655 (N_3655,N_2007,N_2383);
and U3656 (N_3656,N_2576,N_2048);
nor U3657 (N_3657,N_2070,N_2929);
nand U3658 (N_3658,N_2893,N_2657);
and U3659 (N_3659,N_2172,N_2624);
and U3660 (N_3660,N_2534,N_2510);
and U3661 (N_3661,N_2608,N_2274);
nor U3662 (N_3662,N_2791,N_2926);
xnor U3663 (N_3663,N_2950,N_2914);
nand U3664 (N_3664,N_2098,N_2115);
and U3665 (N_3665,N_2301,N_2473);
and U3666 (N_3666,N_2867,N_2343);
xor U3667 (N_3667,N_2187,N_2428);
nand U3668 (N_3668,N_2059,N_2147);
and U3669 (N_3669,N_2168,N_2894);
or U3670 (N_3670,N_2611,N_2046);
or U3671 (N_3671,N_2571,N_2641);
nor U3672 (N_3672,N_2058,N_2943);
and U3673 (N_3673,N_2138,N_2429);
or U3674 (N_3674,N_2318,N_2638);
and U3675 (N_3675,N_2496,N_2720);
or U3676 (N_3676,N_2564,N_2204);
and U3677 (N_3677,N_2511,N_2884);
nand U3678 (N_3678,N_2781,N_2557);
and U3679 (N_3679,N_2211,N_2592);
or U3680 (N_3680,N_2823,N_2711);
nand U3681 (N_3681,N_2931,N_2789);
nor U3682 (N_3682,N_2402,N_2196);
nand U3683 (N_3683,N_2163,N_2007);
nor U3684 (N_3684,N_2866,N_2045);
xnor U3685 (N_3685,N_2643,N_2909);
and U3686 (N_3686,N_2198,N_2556);
xor U3687 (N_3687,N_2344,N_2862);
nor U3688 (N_3688,N_2450,N_2597);
and U3689 (N_3689,N_2802,N_2947);
and U3690 (N_3690,N_2945,N_2845);
xor U3691 (N_3691,N_2225,N_2293);
nand U3692 (N_3692,N_2408,N_2096);
or U3693 (N_3693,N_2064,N_2984);
nor U3694 (N_3694,N_2985,N_2376);
and U3695 (N_3695,N_2489,N_2862);
nand U3696 (N_3696,N_2503,N_2673);
or U3697 (N_3697,N_2828,N_2204);
or U3698 (N_3698,N_2045,N_2082);
or U3699 (N_3699,N_2057,N_2811);
and U3700 (N_3700,N_2573,N_2532);
and U3701 (N_3701,N_2327,N_2073);
or U3702 (N_3702,N_2108,N_2082);
nor U3703 (N_3703,N_2059,N_2687);
or U3704 (N_3704,N_2304,N_2387);
or U3705 (N_3705,N_2372,N_2668);
xnor U3706 (N_3706,N_2649,N_2870);
xnor U3707 (N_3707,N_2794,N_2225);
and U3708 (N_3708,N_2276,N_2375);
and U3709 (N_3709,N_2466,N_2644);
and U3710 (N_3710,N_2076,N_2174);
nand U3711 (N_3711,N_2787,N_2321);
and U3712 (N_3712,N_2159,N_2721);
nand U3713 (N_3713,N_2540,N_2923);
or U3714 (N_3714,N_2133,N_2999);
nand U3715 (N_3715,N_2924,N_2128);
and U3716 (N_3716,N_2574,N_2114);
or U3717 (N_3717,N_2024,N_2362);
nand U3718 (N_3718,N_2944,N_2271);
or U3719 (N_3719,N_2161,N_2608);
nor U3720 (N_3720,N_2637,N_2406);
and U3721 (N_3721,N_2576,N_2532);
nand U3722 (N_3722,N_2660,N_2672);
nand U3723 (N_3723,N_2339,N_2673);
and U3724 (N_3724,N_2985,N_2421);
xor U3725 (N_3725,N_2041,N_2039);
or U3726 (N_3726,N_2556,N_2733);
nand U3727 (N_3727,N_2018,N_2014);
nand U3728 (N_3728,N_2655,N_2030);
nor U3729 (N_3729,N_2096,N_2162);
or U3730 (N_3730,N_2139,N_2126);
and U3731 (N_3731,N_2612,N_2870);
nor U3732 (N_3732,N_2156,N_2003);
nor U3733 (N_3733,N_2856,N_2586);
nand U3734 (N_3734,N_2154,N_2821);
and U3735 (N_3735,N_2060,N_2077);
xor U3736 (N_3736,N_2256,N_2573);
and U3737 (N_3737,N_2248,N_2984);
nand U3738 (N_3738,N_2030,N_2247);
or U3739 (N_3739,N_2407,N_2767);
nor U3740 (N_3740,N_2511,N_2174);
nand U3741 (N_3741,N_2273,N_2540);
or U3742 (N_3742,N_2579,N_2882);
nor U3743 (N_3743,N_2622,N_2009);
nand U3744 (N_3744,N_2155,N_2280);
nor U3745 (N_3745,N_2836,N_2625);
and U3746 (N_3746,N_2413,N_2674);
xor U3747 (N_3747,N_2765,N_2515);
nor U3748 (N_3748,N_2497,N_2620);
and U3749 (N_3749,N_2770,N_2914);
nor U3750 (N_3750,N_2577,N_2314);
nor U3751 (N_3751,N_2553,N_2588);
xnor U3752 (N_3752,N_2878,N_2129);
nor U3753 (N_3753,N_2877,N_2380);
nand U3754 (N_3754,N_2838,N_2435);
or U3755 (N_3755,N_2031,N_2916);
xor U3756 (N_3756,N_2150,N_2200);
nand U3757 (N_3757,N_2368,N_2428);
nor U3758 (N_3758,N_2065,N_2890);
nand U3759 (N_3759,N_2416,N_2309);
nand U3760 (N_3760,N_2577,N_2118);
nor U3761 (N_3761,N_2193,N_2944);
xnor U3762 (N_3762,N_2940,N_2727);
and U3763 (N_3763,N_2046,N_2244);
xor U3764 (N_3764,N_2603,N_2354);
or U3765 (N_3765,N_2985,N_2284);
or U3766 (N_3766,N_2771,N_2828);
or U3767 (N_3767,N_2022,N_2195);
or U3768 (N_3768,N_2457,N_2949);
nand U3769 (N_3769,N_2807,N_2890);
nor U3770 (N_3770,N_2983,N_2459);
or U3771 (N_3771,N_2645,N_2558);
and U3772 (N_3772,N_2410,N_2128);
nor U3773 (N_3773,N_2584,N_2230);
and U3774 (N_3774,N_2123,N_2324);
xnor U3775 (N_3775,N_2143,N_2858);
or U3776 (N_3776,N_2410,N_2864);
or U3777 (N_3777,N_2106,N_2625);
or U3778 (N_3778,N_2601,N_2758);
nand U3779 (N_3779,N_2426,N_2812);
nand U3780 (N_3780,N_2662,N_2591);
xor U3781 (N_3781,N_2030,N_2644);
or U3782 (N_3782,N_2046,N_2441);
or U3783 (N_3783,N_2095,N_2868);
and U3784 (N_3784,N_2338,N_2904);
and U3785 (N_3785,N_2344,N_2575);
nand U3786 (N_3786,N_2576,N_2146);
and U3787 (N_3787,N_2543,N_2997);
and U3788 (N_3788,N_2000,N_2696);
or U3789 (N_3789,N_2008,N_2772);
and U3790 (N_3790,N_2156,N_2218);
or U3791 (N_3791,N_2403,N_2274);
nor U3792 (N_3792,N_2249,N_2938);
nor U3793 (N_3793,N_2047,N_2143);
nor U3794 (N_3794,N_2003,N_2415);
and U3795 (N_3795,N_2461,N_2067);
nor U3796 (N_3796,N_2553,N_2948);
nand U3797 (N_3797,N_2581,N_2379);
and U3798 (N_3798,N_2726,N_2229);
xor U3799 (N_3799,N_2734,N_2187);
nor U3800 (N_3800,N_2841,N_2289);
nor U3801 (N_3801,N_2621,N_2470);
nand U3802 (N_3802,N_2913,N_2035);
nand U3803 (N_3803,N_2002,N_2948);
or U3804 (N_3804,N_2442,N_2182);
nor U3805 (N_3805,N_2603,N_2271);
nor U3806 (N_3806,N_2861,N_2331);
xor U3807 (N_3807,N_2432,N_2517);
nand U3808 (N_3808,N_2802,N_2719);
and U3809 (N_3809,N_2535,N_2672);
nand U3810 (N_3810,N_2638,N_2786);
nand U3811 (N_3811,N_2765,N_2961);
or U3812 (N_3812,N_2623,N_2155);
or U3813 (N_3813,N_2822,N_2922);
nand U3814 (N_3814,N_2631,N_2521);
and U3815 (N_3815,N_2169,N_2248);
xnor U3816 (N_3816,N_2166,N_2826);
xnor U3817 (N_3817,N_2099,N_2007);
nand U3818 (N_3818,N_2306,N_2105);
or U3819 (N_3819,N_2449,N_2988);
nand U3820 (N_3820,N_2544,N_2855);
nand U3821 (N_3821,N_2233,N_2789);
or U3822 (N_3822,N_2421,N_2298);
nor U3823 (N_3823,N_2162,N_2472);
and U3824 (N_3824,N_2786,N_2147);
and U3825 (N_3825,N_2433,N_2902);
nand U3826 (N_3826,N_2272,N_2644);
nor U3827 (N_3827,N_2115,N_2374);
nor U3828 (N_3828,N_2753,N_2899);
or U3829 (N_3829,N_2333,N_2580);
nor U3830 (N_3830,N_2754,N_2394);
or U3831 (N_3831,N_2755,N_2461);
and U3832 (N_3832,N_2527,N_2180);
nand U3833 (N_3833,N_2034,N_2442);
nand U3834 (N_3834,N_2235,N_2656);
and U3835 (N_3835,N_2461,N_2782);
nor U3836 (N_3836,N_2529,N_2204);
or U3837 (N_3837,N_2843,N_2057);
or U3838 (N_3838,N_2513,N_2263);
and U3839 (N_3839,N_2431,N_2081);
nor U3840 (N_3840,N_2968,N_2317);
nand U3841 (N_3841,N_2910,N_2794);
nor U3842 (N_3842,N_2740,N_2868);
and U3843 (N_3843,N_2810,N_2490);
nand U3844 (N_3844,N_2395,N_2139);
nand U3845 (N_3845,N_2840,N_2514);
nand U3846 (N_3846,N_2599,N_2440);
nor U3847 (N_3847,N_2107,N_2562);
and U3848 (N_3848,N_2336,N_2528);
nand U3849 (N_3849,N_2823,N_2440);
nand U3850 (N_3850,N_2993,N_2946);
nor U3851 (N_3851,N_2889,N_2629);
or U3852 (N_3852,N_2473,N_2812);
nor U3853 (N_3853,N_2059,N_2708);
nor U3854 (N_3854,N_2845,N_2161);
or U3855 (N_3855,N_2136,N_2678);
xor U3856 (N_3856,N_2252,N_2748);
and U3857 (N_3857,N_2066,N_2551);
nor U3858 (N_3858,N_2497,N_2135);
nor U3859 (N_3859,N_2002,N_2313);
xor U3860 (N_3860,N_2464,N_2574);
nor U3861 (N_3861,N_2899,N_2987);
nand U3862 (N_3862,N_2970,N_2556);
or U3863 (N_3863,N_2479,N_2250);
or U3864 (N_3864,N_2304,N_2894);
xor U3865 (N_3865,N_2686,N_2586);
and U3866 (N_3866,N_2457,N_2632);
and U3867 (N_3867,N_2635,N_2669);
nand U3868 (N_3868,N_2849,N_2901);
or U3869 (N_3869,N_2275,N_2262);
nand U3870 (N_3870,N_2694,N_2211);
nor U3871 (N_3871,N_2571,N_2236);
nor U3872 (N_3872,N_2253,N_2248);
and U3873 (N_3873,N_2880,N_2168);
or U3874 (N_3874,N_2356,N_2232);
nand U3875 (N_3875,N_2017,N_2697);
nand U3876 (N_3876,N_2491,N_2782);
or U3877 (N_3877,N_2200,N_2967);
nand U3878 (N_3878,N_2603,N_2261);
nor U3879 (N_3879,N_2545,N_2040);
xor U3880 (N_3880,N_2005,N_2369);
nand U3881 (N_3881,N_2178,N_2652);
and U3882 (N_3882,N_2195,N_2424);
nand U3883 (N_3883,N_2813,N_2157);
nor U3884 (N_3884,N_2709,N_2133);
nor U3885 (N_3885,N_2841,N_2130);
nand U3886 (N_3886,N_2136,N_2540);
and U3887 (N_3887,N_2304,N_2290);
and U3888 (N_3888,N_2261,N_2269);
nor U3889 (N_3889,N_2883,N_2038);
or U3890 (N_3890,N_2987,N_2622);
xor U3891 (N_3891,N_2298,N_2169);
nor U3892 (N_3892,N_2957,N_2140);
xnor U3893 (N_3893,N_2902,N_2021);
and U3894 (N_3894,N_2303,N_2634);
nor U3895 (N_3895,N_2635,N_2928);
and U3896 (N_3896,N_2594,N_2179);
or U3897 (N_3897,N_2754,N_2566);
and U3898 (N_3898,N_2869,N_2241);
and U3899 (N_3899,N_2897,N_2815);
nand U3900 (N_3900,N_2640,N_2696);
nand U3901 (N_3901,N_2104,N_2874);
and U3902 (N_3902,N_2215,N_2375);
and U3903 (N_3903,N_2647,N_2140);
nand U3904 (N_3904,N_2397,N_2364);
and U3905 (N_3905,N_2260,N_2421);
xnor U3906 (N_3906,N_2637,N_2245);
xnor U3907 (N_3907,N_2917,N_2765);
nor U3908 (N_3908,N_2708,N_2887);
nor U3909 (N_3909,N_2858,N_2788);
nand U3910 (N_3910,N_2734,N_2725);
nand U3911 (N_3911,N_2378,N_2926);
or U3912 (N_3912,N_2451,N_2462);
and U3913 (N_3913,N_2639,N_2701);
xor U3914 (N_3914,N_2033,N_2602);
and U3915 (N_3915,N_2212,N_2853);
nor U3916 (N_3916,N_2668,N_2483);
nor U3917 (N_3917,N_2882,N_2476);
and U3918 (N_3918,N_2760,N_2039);
or U3919 (N_3919,N_2814,N_2842);
or U3920 (N_3920,N_2699,N_2371);
nand U3921 (N_3921,N_2255,N_2091);
and U3922 (N_3922,N_2331,N_2560);
nand U3923 (N_3923,N_2054,N_2449);
and U3924 (N_3924,N_2389,N_2502);
or U3925 (N_3925,N_2395,N_2353);
or U3926 (N_3926,N_2659,N_2754);
xor U3927 (N_3927,N_2473,N_2971);
and U3928 (N_3928,N_2423,N_2796);
or U3929 (N_3929,N_2492,N_2945);
and U3930 (N_3930,N_2537,N_2197);
or U3931 (N_3931,N_2014,N_2960);
nor U3932 (N_3932,N_2271,N_2987);
and U3933 (N_3933,N_2038,N_2146);
or U3934 (N_3934,N_2924,N_2196);
nand U3935 (N_3935,N_2426,N_2919);
and U3936 (N_3936,N_2855,N_2322);
or U3937 (N_3937,N_2013,N_2267);
and U3938 (N_3938,N_2151,N_2092);
or U3939 (N_3939,N_2602,N_2634);
nand U3940 (N_3940,N_2837,N_2712);
nand U3941 (N_3941,N_2749,N_2067);
nand U3942 (N_3942,N_2702,N_2430);
nand U3943 (N_3943,N_2025,N_2701);
or U3944 (N_3944,N_2153,N_2665);
nor U3945 (N_3945,N_2365,N_2664);
and U3946 (N_3946,N_2626,N_2592);
xor U3947 (N_3947,N_2024,N_2643);
or U3948 (N_3948,N_2170,N_2965);
nand U3949 (N_3949,N_2502,N_2237);
or U3950 (N_3950,N_2637,N_2301);
nand U3951 (N_3951,N_2550,N_2806);
nor U3952 (N_3952,N_2126,N_2542);
and U3953 (N_3953,N_2631,N_2758);
xor U3954 (N_3954,N_2080,N_2273);
nor U3955 (N_3955,N_2999,N_2399);
and U3956 (N_3956,N_2638,N_2785);
nor U3957 (N_3957,N_2220,N_2014);
or U3958 (N_3958,N_2542,N_2619);
and U3959 (N_3959,N_2848,N_2077);
and U3960 (N_3960,N_2492,N_2167);
nor U3961 (N_3961,N_2477,N_2884);
nor U3962 (N_3962,N_2259,N_2947);
nand U3963 (N_3963,N_2574,N_2604);
nand U3964 (N_3964,N_2681,N_2379);
and U3965 (N_3965,N_2879,N_2878);
nand U3966 (N_3966,N_2523,N_2831);
nand U3967 (N_3967,N_2199,N_2422);
or U3968 (N_3968,N_2638,N_2355);
and U3969 (N_3969,N_2419,N_2072);
or U3970 (N_3970,N_2465,N_2770);
and U3971 (N_3971,N_2825,N_2612);
or U3972 (N_3972,N_2727,N_2759);
and U3973 (N_3973,N_2059,N_2653);
nor U3974 (N_3974,N_2688,N_2070);
nor U3975 (N_3975,N_2756,N_2331);
and U3976 (N_3976,N_2042,N_2173);
or U3977 (N_3977,N_2084,N_2194);
nand U3978 (N_3978,N_2985,N_2629);
and U3979 (N_3979,N_2144,N_2654);
or U3980 (N_3980,N_2418,N_2989);
xnor U3981 (N_3981,N_2795,N_2301);
and U3982 (N_3982,N_2520,N_2371);
and U3983 (N_3983,N_2290,N_2934);
nand U3984 (N_3984,N_2216,N_2489);
nor U3985 (N_3985,N_2024,N_2143);
or U3986 (N_3986,N_2697,N_2998);
or U3987 (N_3987,N_2445,N_2153);
or U3988 (N_3988,N_2929,N_2554);
and U3989 (N_3989,N_2165,N_2200);
or U3990 (N_3990,N_2515,N_2860);
nor U3991 (N_3991,N_2671,N_2120);
nor U3992 (N_3992,N_2941,N_2731);
nand U3993 (N_3993,N_2329,N_2237);
nand U3994 (N_3994,N_2968,N_2556);
nor U3995 (N_3995,N_2945,N_2364);
and U3996 (N_3996,N_2715,N_2316);
xor U3997 (N_3997,N_2195,N_2558);
or U3998 (N_3998,N_2251,N_2516);
and U3999 (N_3999,N_2658,N_2894);
and U4000 (N_4000,N_3584,N_3628);
xnor U4001 (N_4001,N_3930,N_3894);
or U4002 (N_4002,N_3813,N_3365);
or U4003 (N_4003,N_3201,N_3383);
or U4004 (N_4004,N_3364,N_3717);
nor U4005 (N_4005,N_3072,N_3457);
nand U4006 (N_4006,N_3555,N_3764);
nor U4007 (N_4007,N_3435,N_3922);
or U4008 (N_4008,N_3734,N_3337);
or U4009 (N_4009,N_3344,N_3835);
nor U4010 (N_4010,N_3226,N_3331);
or U4011 (N_4011,N_3990,N_3233);
nand U4012 (N_4012,N_3304,N_3506);
or U4013 (N_4013,N_3247,N_3927);
and U4014 (N_4014,N_3265,N_3287);
nand U4015 (N_4015,N_3864,N_3722);
nor U4016 (N_4016,N_3066,N_3417);
nor U4017 (N_4017,N_3987,N_3549);
or U4018 (N_4018,N_3370,N_3805);
or U4019 (N_4019,N_3491,N_3915);
and U4020 (N_4020,N_3606,N_3034);
or U4021 (N_4021,N_3103,N_3434);
nor U4022 (N_4022,N_3568,N_3751);
and U4023 (N_4023,N_3673,N_3087);
and U4024 (N_4024,N_3063,N_3594);
nand U4025 (N_4025,N_3207,N_3459);
and U4026 (N_4026,N_3322,N_3901);
nor U4027 (N_4027,N_3264,N_3714);
and U4028 (N_4028,N_3105,N_3500);
nand U4029 (N_4029,N_3040,N_3496);
xor U4030 (N_4030,N_3199,N_3870);
nor U4031 (N_4031,N_3368,N_3601);
nor U4032 (N_4032,N_3398,N_3794);
nor U4033 (N_4033,N_3940,N_3412);
or U4034 (N_4034,N_3746,N_3569);
xnor U4035 (N_4035,N_3984,N_3318);
or U4036 (N_4036,N_3334,N_3249);
xnor U4037 (N_4037,N_3503,N_3876);
nand U4038 (N_4038,N_3709,N_3144);
or U4039 (N_4039,N_3176,N_3655);
nand U4040 (N_4040,N_3015,N_3035);
nand U4041 (N_4041,N_3604,N_3613);
and U4042 (N_4042,N_3728,N_3217);
and U4043 (N_4043,N_3428,N_3971);
nor U4044 (N_4044,N_3460,N_3566);
or U4045 (N_4045,N_3638,N_3493);
or U4046 (N_4046,N_3294,N_3809);
nand U4047 (N_4047,N_3501,N_3982);
or U4048 (N_4048,N_3954,N_3684);
and U4049 (N_4049,N_3316,N_3590);
nand U4050 (N_4050,N_3222,N_3981);
or U4051 (N_4051,N_3831,N_3537);
or U4052 (N_4052,N_3856,N_3492);
nor U4053 (N_4053,N_3119,N_3276);
and U4054 (N_4054,N_3818,N_3482);
nand U4055 (N_4055,N_3351,N_3961);
nor U4056 (N_4056,N_3268,N_3596);
or U4057 (N_4057,N_3760,N_3468);
or U4058 (N_4058,N_3490,N_3887);
xor U4059 (N_4059,N_3785,N_3224);
xnor U4060 (N_4060,N_3693,N_3952);
nor U4061 (N_4061,N_3724,N_3524);
nor U4062 (N_4062,N_3907,N_3977);
nand U4063 (N_4063,N_3630,N_3352);
or U4064 (N_4064,N_3719,N_3081);
or U4065 (N_4065,N_3462,N_3485);
or U4066 (N_4066,N_3645,N_3853);
nor U4067 (N_4067,N_3165,N_3789);
nor U4068 (N_4068,N_3725,N_3410);
nand U4069 (N_4069,N_3857,N_3139);
nand U4070 (N_4070,N_3104,N_3966);
nor U4071 (N_4071,N_3649,N_3096);
nand U4072 (N_4072,N_3502,N_3515);
nand U4073 (N_4073,N_3992,N_3350);
nand U4074 (N_4074,N_3202,N_3327);
or U4075 (N_4075,N_3479,N_3585);
xor U4076 (N_4076,N_3499,N_3388);
nand U4077 (N_4077,N_3127,N_3234);
or U4078 (N_4078,N_3427,N_3988);
nand U4079 (N_4079,N_3057,N_3872);
or U4080 (N_4080,N_3092,N_3797);
nand U4081 (N_4081,N_3484,N_3726);
and U4082 (N_4082,N_3054,N_3102);
nand U4083 (N_4083,N_3681,N_3396);
and U4084 (N_4084,N_3145,N_3836);
xnor U4085 (N_4085,N_3259,N_3423);
nor U4086 (N_4086,N_3420,N_3884);
and U4087 (N_4087,N_3178,N_3413);
and U4088 (N_4088,N_3158,N_3972);
or U4089 (N_4089,N_3611,N_3116);
and U4090 (N_4090,N_3041,N_3416);
nand U4091 (N_4091,N_3674,N_3486);
nor U4092 (N_4092,N_3739,N_3752);
nand U4093 (N_4093,N_3577,N_3934);
nor U4094 (N_4094,N_3100,N_3964);
and U4095 (N_4095,N_3529,N_3730);
nor U4096 (N_4096,N_3669,N_3708);
nor U4097 (N_4097,N_3914,N_3407);
nor U4098 (N_4098,N_3778,N_3373);
nand U4099 (N_4099,N_3204,N_3315);
nand U4100 (N_4100,N_3445,N_3540);
nand U4101 (N_4101,N_3855,N_3180);
and U4102 (N_4102,N_3653,N_3393);
nor U4103 (N_4103,N_3754,N_3313);
xnor U4104 (N_4104,N_3497,N_3565);
and U4105 (N_4105,N_3560,N_3523);
nand U4106 (N_4106,N_3402,N_3290);
or U4107 (N_4107,N_3016,N_3146);
or U4108 (N_4108,N_3477,N_3865);
and U4109 (N_4109,N_3161,N_3000);
and U4110 (N_4110,N_3763,N_3195);
and U4111 (N_4111,N_3617,N_3668);
and U4112 (N_4112,N_3414,N_3854);
or U4113 (N_4113,N_3768,N_3859);
or U4114 (N_4114,N_3051,N_3270);
or U4115 (N_4115,N_3359,N_3436);
or U4116 (N_4116,N_3474,N_3661);
and U4117 (N_4117,N_3683,N_3106);
nand U4118 (N_4118,N_3317,N_3473);
nand U4119 (N_4119,N_3633,N_3291);
nand U4120 (N_4120,N_3896,N_3356);
nor U4121 (N_4121,N_3938,N_3732);
or U4122 (N_4122,N_3533,N_3091);
or U4123 (N_4123,N_3571,N_3235);
nor U4124 (N_4124,N_3518,N_3686);
nand U4125 (N_4125,N_3297,N_3862);
and U4126 (N_4126,N_3128,N_3878);
nor U4127 (N_4127,N_3696,N_3505);
nand U4128 (N_4128,N_3059,N_3527);
nor U4129 (N_4129,N_3548,N_3349);
xnor U4130 (N_4130,N_3136,N_3773);
xor U4131 (N_4131,N_3881,N_3030);
nand U4132 (N_4132,N_3399,N_3392);
nor U4133 (N_4133,N_3824,N_3756);
or U4134 (N_4134,N_3419,N_3153);
or U4135 (N_4135,N_3844,N_3847);
and U4136 (N_4136,N_3821,N_3556);
or U4137 (N_4137,N_3196,N_3579);
and U4138 (N_4138,N_3073,N_3775);
and U4139 (N_4139,N_3082,N_3062);
or U4140 (N_4140,N_3888,N_3899);
nor U4141 (N_4141,N_3080,N_3275);
nor U4142 (N_4142,N_3711,N_3037);
nor U4143 (N_4143,N_3135,N_3170);
xor U4144 (N_4144,N_3042,N_3401);
nor U4145 (N_4145,N_3512,N_3767);
or U4146 (N_4146,N_3788,N_3076);
nand U4147 (N_4147,N_3576,N_3437);
nand U4148 (N_4148,N_3454,N_3229);
nor U4149 (N_4149,N_3210,N_3707);
nand U4150 (N_4150,N_3333,N_3892);
and U4151 (N_4151,N_3761,N_3986);
nor U4152 (N_4152,N_3079,N_3691);
and U4153 (N_4153,N_3935,N_3926);
and U4154 (N_4154,N_3308,N_3162);
or U4155 (N_4155,N_3678,N_3979);
or U4156 (N_4156,N_3608,N_3004);
xor U4157 (N_4157,N_3769,N_3721);
or U4158 (N_4158,N_3177,N_3115);
nand U4159 (N_4159,N_3380,N_3480);
or U4160 (N_4160,N_3074,N_3762);
or U4161 (N_4161,N_3044,N_3587);
or U4162 (N_4162,N_3408,N_3531);
or U4163 (N_4163,N_3923,N_3656);
and U4164 (N_4164,N_3543,N_3747);
nand U4165 (N_4165,N_3688,N_3623);
or U4166 (N_4166,N_3298,N_3188);
nor U4167 (N_4167,N_3791,N_3931);
nand U4168 (N_4168,N_3481,N_3559);
and U4169 (N_4169,N_3302,N_3068);
nand U4170 (N_4170,N_3245,N_3248);
xnor U4171 (N_4171,N_3455,N_3895);
nand U4172 (N_4172,N_3622,N_3804);
nand U4173 (N_4173,N_3913,N_3421);
nor U4174 (N_4174,N_3050,N_3672);
nor U4175 (N_4175,N_3009,N_3243);
nand U4176 (N_4176,N_3991,N_3744);
and U4177 (N_4177,N_3305,N_3993);
nand U4178 (N_4178,N_3320,N_3699);
nand U4179 (N_4179,N_3817,N_3637);
and U4180 (N_4180,N_3600,N_3985);
nor U4181 (N_4181,N_3021,N_3173);
or U4182 (N_4182,N_3160,N_3088);
and U4183 (N_4183,N_3731,N_3609);
nand U4184 (N_4184,N_3553,N_3069);
or U4185 (N_4185,N_3363,N_3443);
nor U4186 (N_4186,N_3967,N_3025);
nor U4187 (N_4187,N_3281,N_3369);
xor U4188 (N_4188,N_3727,N_3379);
xor U4189 (N_4189,N_3347,N_3132);
nand U4190 (N_4190,N_3023,N_3592);
nor U4191 (N_4191,N_3598,N_3017);
or U4192 (N_4192,N_3774,N_3692);
nand U4193 (N_4193,N_3883,N_3114);
nor U4194 (N_4194,N_3650,N_3507);
and U4195 (N_4195,N_3012,N_3535);
nand U4196 (N_4196,N_3263,N_3687);
nor U4197 (N_4197,N_3779,N_3659);
or U4198 (N_4198,N_3142,N_3189);
or U4199 (N_4199,N_3504,N_3526);
nand U4200 (N_4200,N_3123,N_3538);
or U4201 (N_4201,N_3710,N_3620);
and U4202 (N_4202,N_3677,N_3124);
nand U4203 (N_4203,N_3869,N_3439);
and U4204 (N_4204,N_3517,N_3530);
nand U4205 (N_4205,N_3858,N_3642);
or U4206 (N_4206,N_3880,N_3022);
or U4207 (N_4207,N_3163,N_3084);
and U4208 (N_4208,N_3346,N_3203);
or U4209 (N_4209,N_3689,N_3932);
or U4210 (N_4210,N_3277,N_3772);
nand U4211 (N_4211,N_3191,N_3282);
nor U4212 (N_4212,N_3822,N_3787);
or U4213 (N_4213,N_3212,N_3406);
or U4214 (N_4214,N_3194,N_3651);
and U4215 (N_4215,N_3269,N_3340);
or U4216 (N_4216,N_3007,N_3885);
nor U4217 (N_4217,N_3395,N_3255);
nand U4218 (N_4218,N_3682,N_3807);
and U4219 (N_4219,N_3953,N_3781);
nor U4220 (N_4220,N_3262,N_3261);
nor U4221 (N_4221,N_3542,N_3371);
and U4222 (N_4222,N_3572,N_3644);
nand U4223 (N_4223,N_3149,N_3336);
or U4224 (N_4224,N_3450,N_3994);
nor U4225 (N_4225,N_3343,N_3841);
or U4226 (N_4226,N_3950,N_3928);
nor U4227 (N_4227,N_3563,N_3740);
nand U4228 (N_4228,N_3698,N_3877);
nand U4229 (N_4229,N_3758,N_3466);
nor U4230 (N_4230,N_3902,N_3815);
or U4231 (N_4231,N_3999,N_3362);
or U4232 (N_4232,N_3842,N_3832);
nand U4233 (N_4233,N_3920,N_3244);
and U4234 (N_4234,N_3546,N_3273);
xnor U4235 (N_4235,N_3765,N_3064);
and U4236 (N_4236,N_3766,N_3010);
nor U4237 (N_4237,N_3378,N_3141);
or U4238 (N_4238,N_3168,N_3400);
nand U4239 (N_4239,N_3975,N_3147);
nor U4240 (N_4240,N_3285,N_3355);
nor U4241 (N_4241,N_3771,N_3770);
nor U4242 (N_4242,N_3676,N_3863);
nand U4243 (N_4243,N_3581,N_3019);
nor U4244 (N_4244,N_3679,N_3487);
nand U4245 (N_4245,N_3615,N_3257);
nor U4246 (N_4246,N_3575,N_3345);
nor U4247 (N_4247,N_3335,N_3516);
and U4248 (N_4248,N_3254,N_3451);
and U4249 (N_4249,N_3834,N_3970);
or U4250 (N_4250,N_3917,N_3792);
nor U4251 (N_4251,N_3939,N_3452);
nor U4252 (N_4252,N_3933,N_3386);
nand U4253 (N_4253,N_3049,N_3467);
nor U4254 (N_4254,N_3715,N_3949);
and U4255 (N_4255,N_3827,N_3806);
nand U4256 (N_4256,N_3394,N_3470);
nor U4257 (N_4257,N_3839,N_3209);
nand U4258 (N_4258,N_3614,N_3219);
or U4259 (N_4259,N_3444,N_3237);
or U4260 (N_4260,N_3955,N_3670);
nor U4261 (N_4261,N_3635,N_3704);
nor U4262 (N_4262,N_3143,N_3820);
nor U4263 (N_4263,N_3110,N_3544);
and U4264 (N_4264,N_3879,N_3152);
nor U4265 (N_4265,N_3641,N_3886);
nand U4266 (N_4266,N_3648,N_3898);
nand U4267 (N_4267,N_3134,N_3280);
and U4268 (N_4268,N_3086,N_3001);
nand U4269 (N_4269,N_3065,N_3242);
nand U4270 (N_4270,N_3403,N_3666);
nand U4271 (N_4271,N_3299,N_3182);
xor U4272 (N_4272,N_3374,N_3547);
and U4273 (N_4273,N_3843,N_3405);
or U4274 (N_4274,N_3018,N_3310);
and U4275 (N_4275,N_3133,N_3108);
or U4276 (N_4276,N_3958,N_3969);
nor U4277 (N_4277,N_3241,N_3258);
or U4278 (N_4278,N_3183,N_3753);
nor U4279 (N_4279,N_3113,N_3833);
or U4280 (N_4280,N_3539,N_3700);
nor U4281 (N_4281,N_3078,N_3083);
and U4282 (N_4282,N_3591,N_3921);
nand U4283 (N_4283,N_3014,N_3384);
or U4284 (N_4284,N_3665,N_3150);
and U4285 (N_4285,N_3438,N_3494);
or U4286 (N_4286,N_3868,N_3912);
nand U4287 (N_4287,N_3157,N_3849);
and U4288 (N_4288,N_3942,N_3819);
xnor U4289 (N_4289,N_3784,N_3941);
or U4290 (N_4290,N_3675,N_3782);
nand U4291 (N_4291,N_3266,N_3140);
nor U4292 (N_4292,N_3122,N_3639);
xnor U4293 (N_4293,N_3441,N_3094);
xnor U4294 (N_4294,N_3227,N_3341);
and U4295 (N_4295,N_3312,N_3861);
nand U4296 (N_4296,N_3520,N_3366);
and U4297 (N_4297,N_3121,N_3002);
nand U4298 (N_4298,N_3742,N_3137);
or U4299 (N_4299,N_3823,N_3573);
and U4300 (N_4300,N_3893,N_3627);
xnor U4301 (N_4301,N_3610,N_3387);
nand U4302 (N_4302,N_3433,N_3154);
nor U4303 (N_4303,N_3796,N_3588);
and U4304 (N_4304,N_3303,N_3013);
and U4305 (N_4305,N_3267,N_3424);
nand U4306 (N_4306,N_3389,N_3089);
nand U4307 (N_4307,N_3070,N_3697);
and U4308 (N_4308,N_3826,N_3440);
and U4309 (N_4309,N_3960,N_3798);
nor U4310 (N_4310,N_3461,N_3447);
nor U4311 (N_4311,N_3032,N_3962);
nand U4312 (N_4312,N_3422,N_3130);
nand U4313 (N_4313,N_3790,N_3866);
xor U4314 (N_4314,N_3456,N_3213);
or U4315 (N_4315,N_3814,N_3442);
and U4316 (N_4316,N_3125,N_3509);
xor U4317 (N_4317,N_3289,N_3028);
or U4318 (N_4318,N_3446,N_3618);
or U4319 (N_4319,N_3671,N_3381);
nand U4320 (N_4320,N_3458,N_3626);
nand U4321 (N_4321,N_3723,N_3253);
nand U4322 (N_4322,N_3712,N_3521);
or U4323 (N_4323,N_3166,N_3075);
and U4324 (N_4324,N_3179,N_3875);
nand U4325 (N_4325,N_3107,N_3514);
nor U4326 (N_4326,N_3471,N_3937);
nor U4327 (N_4327,N_3067,N_3929);
nand U4328 (N_4328,N_3326,N_3031);
nor U4329 (N_4329,N_3956,N_3783);
xnor U4330 (N_4330,N_3580,N_3713);
or U4331 (N_4331,N_3293,N_3348);
nand U4332 (N_4332,N_3251,N_3647);
xnor U4333 (N_4333,N_3228,N_3184);
nand U4334 (N_4334,N_3595,N_3662);
and U4335 (N_4335,N_3936,N_3582);
nand U4336 (N_4336,N_3216,N_3198);
nor U4337 (N_4337,N_3658,N_3567);
nor U4338 (N_4338,N_3328,N_3808);
nor U4339 (N_4339,N_3172,N_3301);
nand U4340 (N_4340,N_3279,N_3570);
and U4341 (N_4341,N_3963,N_3033);
and U4342 (N_4342,N_3519,N_3612);
nor U4343 (N_4343,N_3867,N_3616);
nor U4344 (N_4344,N_3850,N_3957);
and U4345 (N_4345,N_3916,N_3552);
nor U4346 (N_4346,N_3705,N_3685);
and U4347 (N_4347,N_3093,N_3223);
nor U4348 (N_4348,N_3718,N_3632);
or U4349 (N_4349,N_3271,N_3508);
or U4350 (N_4350,N_3260,N_3680);
nor U4351 (N_4351,N_3816,N_3098);
nor U4352 (N_4352,N_3578,N_3541);
or U4353 (N_4353,N_3453,N_3738);
nor U4354 (N_4354,N_3206,N_3488);
nor U4355 (N_4355,N_3636,N_3755);
nand U4356 (N_4356,N_3874,N_3667);
and U4357 (N_4357,N_3562,N_3583);
xor U4358 (N_4358,N_3558,N_3748);
and U4359 (N_4359,N_3968,N_3214);
or U4360 (N_4360,N_3469,N_3510);
xor U4361 (N_4361,N_3976,N_3353);
and U4362 (N_4362,N_3998,N_3882);
nand U4363 (N_4363,N_3904,N_3429);
and U4364 (N_4364,N_3024,N_3288);
nand U4365 (N_4365,N_3360,N_3889);
and U4366 (N_4366,N_3077,N_3274);
nand U4367 (N_4367,N_3174,N_3409);
or U4368 (N_4368,N_3425,N_3621);
nand U4369 (N_4369,N_3483,N_3947);
nor U4370 (N_4370,N_3837,N_3367);
or U4371 (N_4371,N_3812,N_3099);
nand U4372 (N_4372,N_3476,N_3852);
nand U4373 (N_4373,N_3589,N_3238);
and U4374 (N_4374,N_3151,N_3924);
or U4375 (N_4375,N_3250,N_3897);
xnor U4376 (N_4376,N_3786,N_3489);
nor U4377 (N_4377,N_3118,N_3043);
nor U4378 (N_4378,N_3376,N_3300);
and U4379 (N_4379,N_3959,N_3205);
and U4380 (N_4380,N_3735,N_3286);
and U4381 (N_4381,N_3472,N_3586);
nand U4382 (N_4382,N_3185,N_3737);
or U4383 (N_4383,N_3943,N_3664);
and U4384 (N_4384,N_3946,N_3871);
nand U4385 (N_4385,N_3272,N_3382);
or U4386 (N_4386,N_3278,N_3741);
nor U4387 (N_4387,N_3925,N_3169);
nor U4388 (N_4388,N_3003,N_3840);
or U4389 (N_4389,N_3375,N_3148);
nor U4390 (N_4390,N_3495,N_3995);
nor U4391 (N_4391,N_3354,N_3720);
and U4392 (N_4392,N_3605,N_3463);
nand U4393 (N_4393,N_3646,N_3554);
nor U4394 (N_4394,N_3232,N_3906);
nor U4395 (N_4395,N_3706,N_3513);
and U4396 (N_4396,N_3256,N_3625);
and U4397 (N_4397,N_3944,N_3385);
nor U4398 (N_4398,N_3574,N_3187);
nand U4399 (N_4399,N_3095,N_3283);
nand U4400 (N_4400,N_3603,N_3802);
and U4401 (N_4401,N_3339,N_3903);
and U4402 (N_4402,N_3211,N_3631);
nand U4403 (N_4403,N_3101,N_3319);
nor U4404 (N_4404,N_3053,N_3061);
and U4405 (N_4405,N_3431,N_3624);
or U4406 (N_4406,N_3208,N_3749);
nand U4407 (N_4407,N_3052,N_3777);
nor U4408 (N_4408,N_3743,N_3973);
xor U4409 (N_4409,N_3619,N_3989);
or U4410 (N_4410,N_3311,N_3221);
or U4411 (N_4411,N_3757,N_3550);
or U4412 (N_4412,N_3860,N_3323);
nand U4413 (N_4413,N_3090,N_3060);
or U4414 (N_4414,N_3948,N_3006);
or U4415 (N_4415,N_3810,N_3974);
or U4416 (N_4416,N_3186,N_3891);
or U4417 (N_4417,N_3701,N_3129);
nand U4418 (N_4418,N_3338,N_3377);
xor U4419 (N_4419,N_3890,N_3745);
or U4420 (N_4420,N_3663,N_3190);
xor U4421 (N_4421,N_3329,N_3602);
or U4422 (N_4422,N_3131,N_3332);
or U4423 (N_4423,N_3391,N_3545);
nor U4424 (N_4424,N_3225,N_3838);
nor U4425 (N_4425,N_3799,N_3085);
xor U4426 (N_4426,N_3138,N_3164);
nor U4427 (N_4427,N_3008,N_3218);
nand U4428 (N_4428,N_3643,N_3733);
nor U4429 (N_4429,N_3324,N_3900);
or U4430 (N_4430,N_3528,N_3197);
or U4431 (N_4431,N_3246,N_3593);
and U4432 (N_4432,N_3390,N_3951);
and U4433 (N_4433,N_3426,N_3415);
or U4434 (N_4434,N_3607,N_3511);
xnor U4435 (N_4435,N_3561,N_3905);
and U4436 (N_4436,N_3918,N_3236);
xnor U4437 (N_4437,N_3851,N_3800);
xor U4438 (N_4438,N_3846,N_3314);
and U4439 (N_4439,N_3690,N_3361);
and U4440 (N_4440,N_3220,N_3629);
nor U4441 (N_4441,N_3397,N_3534);
nand U4442 (N_4442,N_3181,N_3215);
nand U4443 (N_4443,N_3702,N_3793);
nand U4444 (N_4444,N_3536,N_3156);
xor U4445 (N_4445,N_3111,N_3432);
nand U4446 (N_4446,N_3634,N_3155);
nand U4447 (N_4447,N_3532,N_3945);
nor U4448 (N_4448,N_3703,N_3097);
and U4449 (N_4449,N_3449,N_3047);
xor U4450 (N_4450,N_3026,N_3997);
and U4451 (N_4451,N_3240,N_3252);
and U4452 (N_4452,N_3660,N_3284);
nand U4453 (N_4453,N_3372,N_3039);
or U4454 (N_4454,N_3193,N_3296);
nand U4455 (N_4455,N_3171,N_3759);
nor U4456 (N_4456,N_3848,N_3695);
nand U4457 (N_4457,N_3795,N_3411);
and U4458 (N_4458,N_3230,N_3448);
and U4459 (N_4459,N_3551,N_3597);
nor U4460 (N_4460,N_3776,N_3910);
nor U4461 (N_4461,N_3295,N_3873);
xnor U4462 (N_4462,N_3750,N_3117);
or U4463 (N_4463,N_3657,N_3729);
nand U4464 (N_4464,N_3465,N_3342);
and U4465 (N_4465,N_3475,N_3330);
and U4466 (N_4466,N_3640,N_3803);
and U4467 (N_4467,N_3829,N_3716);
or U4468 (N_4468,N_3564,N_3909);
or U4469 (N_4469,N_3200,N_3306);
or U4470 (N_4470,N_3498,N_3736);
nor U4471 (N_4471,N_3996,N_3464);
nor U4472 (N_4472,N_3978,N_3038);
nand U4473 (N_4473,N_3056,N_3830);
nor U4474 (N_4474,N_3694,N_3321);
nand U4475 (N_4475,N_3522,N_3005);
xor U4476 (N_4476,N_3036,N_3126);
xnor U4477 (N_4477,N_3801,N_3404);
nor U4478 (N_4478,N_3011,N_3965);
and U4479 (N_4479,N_3159,N_3557);
and U4480 (N_4480,N_3055,N_3109);
nor U4481 (N_4481,N_3175,N_3828);
or U4482 (N_4482,N_3020,N_3120);
xor U4483 (N_4483,N_3358,N_3292);
and U4484 (N_4484,N_3780,N_3357);
nor U4485 (N_4485,N_3811,N_3027);
xor U4486 (N_4486,N_3980,N_3845);
or U4487 (N_4487,N_3239,N_3418);
nand U4488 (N_4488,N_3048,N_3908);
or U4489 (N_4489,N_3309,N_3599);
or U4490 (N_4490,N_3029,N_3652);
or U4491 (N_4491,N_3192,N_3983);
nand U4492 (N_4492,N_3825,N_3307);
or U4493 (N_4493,N_3525,N_3046);
nor U4494 (N_4494,N_3911,N_3654);
or U4495 (N_4495,N_3325,N_3045);
xnor U4496 (N_4496,N_3167,N_3231);
nand U4497 (N_4497,N_3071,N_3430);
or U4498 (N_4498,N_3919,N_3112);
or U4499 (N_4499,N_3478,N_3058);
or U4500 (N_4500,N_3149,N_3621);
and U4501 (N_4501,N_3041,N_3372);
or U4502 (N_4502,N_3180,N_3254);
nand U4503 (N_4503,N_3259,N_3756);
xor U4504 (N_4504,N_3463,N_3641);
nor U4505 (N_4505,N_3612,N_3790);
or U4506 (N_4506,N_3497,N_3698);
nor U4507 (N_4507,N_3990,N_3068);
nand U4508 (N_4508,N_3865,N_3008);
or U4509 (N_4509,N_3985,N_3443);
nand U4510 (N_4510,N_3830,N_3431);
and U4511 (N_4511,N_3506,N_3815);
nor U4512 (N_4512,N_3844,N_3333);
nand U4513 (N_4513,N_3088,N_3038);
nand U4514 (N_4514,N_3556,N_3425);
and U4515 (N_4515,N_3445,N_3797);
or U4516 (N_4516,N_3818,N_3856);
nand U4517 (N_4517,N_3906,N_3988);
nand U4518 (N_4518,N_3588,N_3870);
and U4519 (N_4519,N_3233,N_3802);
and U4520 (N_4520,N_3164,N_3137);
and U4521 (N_4521,N_3854,N_3736);
and U4522 (N_4522,N_3091,N_3399);
and U4523 (N_4523,N_3706,N_3758);
and U4524 (N_4524,N_3744,N_3078);
or U4525 (N_4525,N_3933,N_3283);
or U4526 (N_4526,N_3062,N_3656);
and U4527 (N_4527,N_3913,N_3260);
and U4528 (N_4528,N_3861,N_3650);
nor U4529 (N_4529,N_3439,N_3979);
nand U4530 (N_4530,N_3922,N_3025);
nand U4531 (N_4531,N_3908,N_3477);
and U4532 (N_4532,N_3685,N_3596);
nor U4533 (N_4533,N_3315,N_3884);
or U4534 (N_4534,N_3084,N_3503);
nand U4535 (N_4535,N_3406,N_3788);
nand U4536 (N_4536,N_3403,N_3995);
nor U4537 (N_4537,N_3011,N_3407);
nor U4538 (N_4538,N_3191,N_3460);
or U4539 (N_4539,N_3263,N_3856);
or U4540 (N_4540,N_3850,N_3183);
or U4541 (N_4541,N_3840,N_3402);
nand U4542 (N_4542,N_3021,N_3863);
xnor U4543 (N_4543,N_3244,N_3136);
nand U4544 (N_4544,N_3506,N_3176);
or U4545 (N_4545,N_3687,N_3784);
nand U4546 (N_4546,N_3186,N_3246);
or U4547 (N_4547,N_3073,N_3841);
and U4548 (N_4548,N_3801,N_3401);
nor U4549 (N_4549,N_3093,N_3107);
xnor U4550 (N_4550,N_3594,N_3107);
or U4551 (N_4551,N_3586,N_3857);
nor U4552 (N_4552,N_3458,N_3373);
xor U4553 (N_4553,N_3762,N_3979);
nor U4554 (N_4554,N_3027,N_3826);
nor U4555 (N_4555,N_3293,N_3810);
nor U4556 (N_4556,N_3409,N_3567);
nor U4557 (N_4557,N_3450,N_3365);
xnor U4558 (N_4558,N_3497,N_3352);
and U4559 (N_4559,N_3196,N_3867);
or U4560 (N_4560,N_3142,N_3995);
nor U4561 (N_4561,N_3659,N_3248);
xor U4562 (N_4562,N_3821,N_3657);
or U4563 (N_4563,N_3294,N_3152);
and U4564 (N_4564,N_3972,N_3823);
nor U4565 (N_4565,N_3406,N_3905);
and U4566 (N_4566,N_3316,N_3341);
and U4567 (N_4567,N_3187,N_3960);
nand U4568 (N_4568,N_3819,N_3249);
and U4569 (N_4569,N_3592,N_3079);
and U4570 (N_4570,N_3430,N_3874);
or U4571 (N_4571,N_3134,N_3498);
nor U4572 (N_4572,N_3838,N_3952);
nand U4573 (N_4573,N_3465,N_3038);
and U4574 (N_4574,N_3870,N_3545);
nand U4575 (N_4575,N_3368,N_3767);
nand U4576 (N_4576,N_3403,N_3594);
or U4577 (N_4577,N_3437,N_3549);
nand U4578 (N_4578,N_3162,N_3340);
or U4579 (N_4579,N_3726,N_3869);
or U4580 (N_4580,N_3756,N_3806);
nor U4581 (N_4581,N_3235,N_3965);
nand U4582 (N_4582,N_3172,N_3179);
or U4583 (N_4583,N_3329,N_3238);
xor U4584 (N_4584,N_3150,N_3258);
or U4585 (N_4585,N_3750,N_3426);
xor U4586 (N_4586,N_3355,N_3477);
xor U4587 (N_4587,N_3755,N_3044);
nor U4588 (N_4588,N_3923,N_3395);
and U4589 (N_4589,N_3062,N_3414);
or U4590 (N_4590,N_3780,N_3031);
or U4591 (N_4591,N_3074,N_3787);
and U4592 (N_4592,N_3006,N_3823);
nor U4593 (N_4593,N_3145,N_3882);
nor U4594 (N_4594,N_3784,N_3676);
and U4595 (N_4595,N_3112,N_3162);
or U4596 (N_4596,N_3236,N_3248);
and U4597 (N_4597,N_3700,N_3836);
xnor U4598 (N_4598,N_3666,N_3934);
or U4599 (N_4599,N_3165,N_3830);
or U4600 (N_4600,N_3498,N_3805);
nand U4601 (N_4601,N_3817,N_3229);
or U4602 (N_4602,N_3920,N_3771);
nand U4603 (N_4603,N_3072,N_3496);
and U4604 (N_4604,N_3233,N_3454);
nor U4605 (N_4605,N_3160,N_3303);
nand U4606 (N_4606,N_3213,N_3255);
and U4607 (N_4607,N_3206,N_3082);
or U4608 (N_4608,N_3379,N_3329);
xor U4609 (N_4609,N_3523,N_3229);
nor U4610 (N_4610,N_3556,N_3888);
and U4611 (N_4611,N_3232,N_3927);
or U4612 (N_4612,N_3218,N_3155);
or U4613 (N_4613,N_3225,N_3871);
nand U4614 (N_4614,N_3980,N_3956);
or U4615 (N_4615,N_3675,N_3746);
xor U4616 (N_4616,N_3833,N_3060);
or U4617 (N_4617,N_3634,N_3209);
or U4618 (N_4618,N_3014,N_3091);
or U4619 (N_4619,N_3848,N_3209);
nand U4620 (N_4620,N_3841,N_3001);
and U4621 (N_4621,N_3102,N_3362);
nor U4622 (N_4622,N_3628,N_3351);
nor U4623 (N_4623,N_3755,N_3802);
xnor U4624 (N_4624,N_3786,N_3388);
xor U4625 (N_4625,N_3575,N_3459);
and U4626 (N_4626,N_3901,N_3613);
and U4627 (N_4627,N_3165,N_3174);
and U4628 (N_4628,N_3931,N_3720);
or U4629 (N_4629,N_3079,N_3449);
and U4630 (N_4630,N_3333,N_3865);
or U4631 (N_4631,N_3998,N_3330);
nand U4632 (N_4632,N_3031,N_3417);
xnor U4633 (N_4633,N_3985,N_3156);
and U4634 (N_4634,N_3573,N_3285);
nand U4635 (N_4635,N_3920,N_3680);
or U4636 (N_4636,N_3980,N_3963);
nor U4637 (N_4637,N_3854,N_3956);
or U4638 (N_4638,N_3848,N_3100);
xor U4639 (N_4639,N_3302,N_3852);
nand U4640 (N_4640,N_3052,N_3538);
or U4641 (N_4641,N_3996,N_3974);
and U4642 (N_4642,N_3543,N_3533);
nor U4643 (N_4643,N_3614,N_3827);
nor U4644 (N_4644,N_3136,N_3851);
nand U4645 (N_4645,N_3696,N_3551);
xnor U4646 (N_4646,N_3749,N_3176);
and U4647 (N_4647,N_3793,N_3878);
nor U4648 (N_4648,N_3878,N_3414);
nand U4649 (N_4649,N_3454,N_3071);
or U4650 (N_4650,N_3298,N_3917);
nand U4651 (N_4651,N_3054,N_3596);
or U4652 (N_4652,N_3448,N_3091);
xnor U4653 (N_4653,N_3111,N_3222);
nand U4654 (N_4654,N_3728,N_3833);
or U4655 (N_4655,N_3751,N_3385);
and U4656 (N_4656,N_3529,N_3800);
nand U4657 (N_4657,N_3047,N_3668);
or U4658 (N_4658,N_3521,N_3144);
and U4659 (N_4659,N_3201,N_3549);
or U4660 (N_4660,N_3912,N_3949);
or U4661 (N_4661,N_3584,N_3837);
nor U4662 (N_4662,N_3634,N_3205);
nor U4663 (N_4663,N_3011,N_3550);
nand U4664 (N_4664,N_3127,N_3555);
and U4665 (N_4665,N_3187,N_3132);
and U4666 (N_4666,N_3168,N_3453);
and U4667 (N_4667,N_3677,N_3422);
nand U4668 (N_4668,N_3852,N_3861);
nand U4669 (N_4669,N_3964,N_3044);
and U4670 (N_4670,N_3301,N_3679);
and U4671 (N_4671,N_3929,N_3751);
or U4672 (N_4672,N_3280,N_3513);
nor U4673 (N_4673,N_3024,N_3867);
nor U4674 (N_4674,N_3546,N_3355);
and U4675 (N_4675,N_3673,N_3050);
nand U4676 (N_4676,N_3968,N_3805);
nor U4677 (N_4677,N_3450,N_3619);
nand U4678 (N_4678,N_3722,N_3867);
and U4679 (N_4679,N_3926,N_3465);
nand U4680 (N_4680,N_3148,N_3173);
and U4681 (N_4681,N_3698,N_3419);
nor U4682 (N_4682,N_3135,N_3314);
nand U4683 (N_4683,N_3391,N_3015);
or U4684 (N_4684,N_3419,N_3903);
xor U4685 (N_4685,N_3521,N_3455);
nor U4686 (N_4686,N_3542,N_3650);
and U4687 (N_4687,N_3235,N_3751);
or U4688 (N_4688,N_3212,N_3776);
nor U4689 (N_4689,N_3034,N_3929);
and U4690 (N_4690,N_3591,N_3377);
nand U4691 (N_4691,N_3666,N_3988);
and U4692 (N_4692,N_3235,N_3953);
nor U4693 (N_4693,N_3683,N_3412);
or U4694 (N_4694,N_3725,N_3985);
nand U4695 (N_4695,N_3914,N_3710);
and U4696 (N_4696,N_3747,N_3072);
nand U4697 (N_4697,N_3819,N_3056);
nor U4698 (N_4698,N_3973,N_3573);
and U4699 (N_4699,N_3858,N_3006);
and U4700 (N_4700,N_3188,N_3137);
and U4701 (N_4701,N_3940,N_3717);
and U4702 (N_4702,N_3182,N_3043);
or U4703 (N_4703,N_3491,N_3360);
nor U4704 (N_4704,N_3759,N_3680);
or U4705 (N_4705,N_3062,N_3540);
xor U4706 (N_4706,N_3885,N_3335);
or U4707 (N_4707,N_3802,N_3278);
nor U4708 (N_4708,N_3718,N_3281);
nand U4709 (N_4709,N_3601,N_3393);
nand U4710 (N_4710,N_3578,N_3445);
and U4711 (N_4711,N_3502,N_3327);
nor U4712 (N_4712,N_3451,N_3610);
and U4713 (N_4713,N_3078,N_3890);
and U4714 (N_4714,N_3779,N_3286);
nand U4715 (N_4715,N_3102,N_3739);
or U4716 (N_4716,N_3983,N_3382);
or U4717 (N_4717,N_3918,N_3591);
nand U4718 (N_4718,N_3393,N_3898);
nor U4719 (N_4719,N_3509,N_3622);
or U4720 (N_4720,N_3911,N_3082);
and U4721 (N_4721,N_3627,N_3809);
nand U4722 (N_4722,N_3192,N_3562);
and U4723 (N_4723,N_3539,N_3742);
nand U4724 (N_4724,N_3907,N_3675);
nand U4725 (N_4725,N_3478,N_3365);
nor U4726 (N_4726,N_3487,N_3984);
nand U4727 (N_4727,N_3535,N_3026);
nor U4728 (N_4728,N_3238,N_3824);
nor U4729 (N_4729,N_3042,N_3083);
nor U4730 (N_4730,N_3871,N_3095);
nand U4731 (N_4731,N_3560,N_3984);
nand U4732 (N_4732,N_3290,N_3358);
nand U4733 (N_4733,N_3469,N_3068);
nand U4734 (N_4734,N_3145,N_3215);
xor U4735 (N_4735,N_3061,N_3205);
nand U4736 (N_4736,N_3848,N_3681);
and U4737 (N_4737,N_3849,N_3942);
or U4738 (N_4738,N_3843,N_3873);
or U4739 (N_4739,N_3391,N_3229);
nor U4740 (N_4740,N_3499,N_3257);
nand U4741 (N_4741,N_3413,N_3869);
or U4742 (N_4742,N_3977,N_3308);
nand U4743 (N_4743,N_3736,N_3043);
and U4744 (N_4744,N_3079,N_3884);
or U4745 (N_4745,N_3910,N_3889);
or U4746 (N_4746,N_3066,N_3781);
and U4747 (N_4747,N_3708,N_3645);
or U4748 (N_4748,N_3198,N_3815);
and U4749 (N_4749,N_3644,N_3486);
nand U4750 (N_4750,N_3283,N_3354);
or U4751 (N_4751,N_3077,N_3457);
or U4752 (N_4752,N_3891,N_3080);
and U4753 (N_4753,N_3903,N_3600);
nand U4754 (N_4754,N_3573,N_3665);
or U4755 (N_4755,N_3697,N_3401);
nor U4756 (N_4756,N_3141,N_3327);
nand U4757 (N_4757,N_3575,N_3468);
nand U4758 (N_4758,N_3049,N_3526);
nor U4759 (N_4759,N_3642,N_3882);
nor U4760 (N_4760,N_3903,N_3921);
nand U4761 (N_4761,N_3830,N_3187);
or U4762 (N_4762,N_3607,N_3025);
xor U4763 (N_4763,N_3819,N_3854);
or U4764 (N_4764,N_3141,N_3792);
nand U4765 (N_4765,N_3902,N_3403);
nand U4766 (N_4766,N_3646,N_3144);
or U4767 (N_4767,N_3838,N_3574);
or U4768 (N_4768,N_3297,N_3779);
nand U4769 (N_4769,N_3964,N_3870);
and U4770 (N_4770,N_3583,N_3104);
nand U4771 (N_4771,N_3620,N_3974);
nand U4772 (N_4772,N_3748,N_3111);
and U4773 (N_4773,N_3662,N_3856);
nor U4774 (N_4774,N_3792,N_3014);
or U4775 (N_4775,N_3732,N_3184);
nor U4776 (N_4776,N_3726,N_3901);
and U4777 (N_4777,N_3991,N_3284);
and U4778 (N_4778,N_3729,N_3445);
or U4779 (N_4779,N_3855,N_3318);
or U4780 (N_4780,N_3735,N_3646);
xnor U4781 (N_4781,N_3949,N_3995);
nand U4782 (N_4782,N_3161,N_3025);
xor U4783 (N_4783,N_3385,N_3914);
nand U4784 (N_4784,N_3297,N_3667);
nor U4785 (N_4785,N_3684,N_3492);
nor U4786 (N_4786,N_3563,N_3927);
nand U4787 (N_4787,N_3559,N_3996);
xor U4788 (N_4788,N_3853,N_3934);
or U4789 (N_4789,N_3680,N_3925);
and U4790 (N_4790,N_3737,N_3543);
or U4791 (N_4791,N_3457,N_3713);
and U4792 (N_4792,N_3292,N_3959);
nor U4793 (N_4793,N_3143,N_3748);
or U4794 (N_4794,N_3859,N_3907);
or U4795 (N_4795,N_3925,N_3109);
or U4796 (N_4796,N_3019,N_3518);
nand U4797 (N_4797,N_3111,N_3327);
xnor U4798 (N_4798,N_3499,N_3213);
nor U4799 (N_4799,N_3977,N_3199);
nor U4800 (N_4800,N_3512,N_3685);
or U4801 (N_4801,N_3197,N_3536);
nor U4802 (N_4802,N_3725,N_3691);
and U4803 (N_4803,N_3871,N_3821);
and U4804 (N_4804,N_3818,N_3181);
or U4805 (N_4805,N_3367,N_3705);
nand U4806 (N_4806,N_3026,N_3615);
and U4807 (N_4807,N_3256,N_3244);
xor U4808 (N_4808,N_3701,N_3368);
or U4809 (N_4809,N_3108,N_3314);
and U4810 (N_4810,N_3495,N_3052);
and U4811 (N_4811,N_3834,N_3271);
nand U4812 (N_4812,N_3092,N_3791);
xnor U4813 (N_4813,N_3501,N_3793);
or U4814 (N_4814,N_3477,N_3970);
xor U4815 (N_4815,N_3685,N_3657);
and U4816 (N_4816,N_3098,N_3107);
nand U4817 (N_4817,N_3445,N_3631);
nand U4818 (N_4818,N_3032,N_3132);
nor U4819 (N_4819,N_3839,N_3016);
nor U4820 (N_4820,N_3118,N_3046);
and U4821 (N_4821,N_3888,N_3797);
or U4822 (N_4822,N_3596,N_3024);
nand U4823 (N_4823,N_3152,N_3421);
nand U4824 (N_4824,N_3143,N_3066);
nor U4825 (N_4825,N_3273,N_3003);
and U4826 (N_4826,N_3763,N_3420);
nand U4827 (N_4827,N_3872,N_3914);
nor U4828 (N_4828,N_3416,N_3635);
or U4829 (N_4829,N_3902,N_3095);
and U4830 (N_4830,N_3096,N_3552);
nor U4831 (N_4831,N_3682,N_3869);
and U4832 (N_4832,N_3972,N_3206);
nor U4833 (N_4833,N_3483,N_3142);
and U4834 (N_4834,N_3505,N_3601);
xor U4835 (N_4835,N_3563,N_3557);
and U4836 (N_4836,N_3670,N_3447);
or U4837 (N_4837,N_3764,N_3949);
nor U4838 (N_4838,N_3382,N_3000);
xor U4839 (N_4839,N_3367,N_3169);
nand U4840 (N_4840,N_3642,N_3424);
and U4841 (N_4841,N_3203,N_3277);
nand U4842 (N_4842,N_3450,N_3443);
nand U4843 (N_4843,N_3691,N_3914);
or U4844 (N_4844,N_3614,N_3240);
and U4845 (N_4845,N_3250,N_3963);
and U4846 (N_4846,N_3251,N_3010);
nor U4847 (N_4847,N_3076,N_3737);
or U4848 (N_4848,N_3431,N_3047);
and U4849 (N_4849,N_3623,N_3322);
nor U4850 (N_4850,N_3890,N_3439);
and U4851 (N_4851,N_3801,N_3473);
or U4852 (N_4852,N_3856,N_3037);
and U4853 (N_4853,N_3286,N_3709);
xor U4854 (N_4854,N_3165,N_3056);
and U4855 (N_4855,N_3229,N_3378);
nor U4856 (N_4856,N_3644,N_3050);
nor U4857 (N_4857,N_3917,N_3002);
or U4858 (N_4858,N_3049,N_3251);
nand U4859 (N_4859,N_3231,N_3321);
xor U4860 (N_4860,N_3303,N_3276);
xnor U4861 (N_4861,N_3868,N_3869);
or U4862 (N_4862,N_3530,N_3611);
nand U4863 (N_4863,N_3811,N_3578);
xor U4864 (N_4864,N_3438,N_3953);
nand U4865 (N_4865,N_3520,N_3131);
and U4866 (N_4866,N_3213,N_3424);
nand U4867 (N_4867,N_3388,N_3154);
nand U4868 (N_4868,N_3671,N_3908);
nor U4869 (N_4869,N_3730,N_3465);
and U4870 (N_4870,N_3528,N_3852);
and U4871 (N_4871,N_3194,N_3681);
or U4872 (N_4872,N_3330,N_3927);
nor U4873 (N_4873,N_3056,N_3201);
nor U4874 (N_4874,N_3512,N_3594);
xnor U4875 (N_4875,N_3072,N_3168);
nand U4876 (N_4876,N_3752,N_3518);
and U4877 (N_4877,N_3808,N_3409);
and U4878 (N_4878,N_3686,N_3015);
nand U4879 (N_4879,N_3025,N_3239);
or U4880 (N_4880,N_3995,N_3519);
and U4881 (N_4881,N_3464,N_3882);
nor U4882 (N_4882,N_3875,N_3334);
nor U4883 (N_4883,N_3429,N_3517);
or U4884 (N_4884,N_3282,N_3511);
or U4885 (N_4885,N_3541,N_3592);
nor U4886 (N_4886,N_3062,N_3044);
nor U4887 (N_4887,N_3072,N_3660);
xor U4888 (N_4888,N_3043,N_3287);
and U4889 (N_4889,N_3525,N_3377);
nand U4890 (N_4890,N_3505,N_3502);
nor U4891 (N_4891,N_3118,N_3195);
nand U4892 (N_4892,N_3711,N_3175);
nand U4893 (N_4893,N_3434,N_3734);
nand U4894 (N_4894,N_3304,N_3676);
nor U4895 (N_4895,N_3129,N_3511);
or U4896 (N_4896,N_3693,N_3720);
and U4897 (N_4897,N_3331,N_3947);
or U4898 (N_4898,N_3258,N_3873);
nand U4899 (N_4899,N_3068,N_3696);
nand U4900 (N_4900,N_3837,N_3628);
or U4901 (N_4901,N_3473,N_3088);
nand U4902 (N_4902,N_3295,N_3232);
nand U4903 (N_4903,N_3219,N_3057);
or U4904 (N_4904,N_3370,N_3081);
or U4905 (N_4905,N_3933,N_3821);
nor U4906 (N_4906,N_3983,N_3925);
nand U4907 (N_4907,N_3086,N_3918);
nor U4908 (N_4908,N_3168,N_3219);
and U4909 (N_4909,N_3577,N_3522);
nand U4910 (N_4910,N_3203,N_3242);
nand U4911 (N_4911,N_3913,N_3612);
or U4912 (N_4912,N_3109,N_3725);
and U4913 (N_4913,N_3446,N_3528);
nand U4914 (N_4914,N_3146,N_3541);
or U4915 (N_4915,N_3060,N_3753);
and U4916 (N_4916,N_3612,N_3772);
and U4917 (N_4917,N_3364,N_3311);
and U4918 (N_4918,N_3615,N_3910);
nand U4919 (N_4919,N_3278,N_3891);
or U4920 (N_4920,N_3231,N_3481);
and U4921 (N_4921,N_3538,N_3965);
and U4922 (N_4922,N_3399,N_3006);
and U4923 (N_4923,N_3910,N_3535);
nor U4924 (N_4924,N_3604,N_3202);
nand U4925 (N_4925,N_3715,N_3670);
nor U4926 (N_4926,N_3919,N_3840);
xnor U4927 (N_4927,N_3407,N_3960);
or U4928 (N_4928,N_3832,N_3879);
nand U4929 (N_4929,N_3580,N_3919);
nor U4930 (N_4930,N_3872,N_3580);
nand U4931 (N_4931,N_3466,N_3599);
or U4932 (N_4932,N_3257,N_3702);
nand U4933 (N_4933,N_3972,N_3192);
and U4934 (N_4934,N_3130,N_3628);
nand U4935 (N_4935,N_3833,N_3284);
nor U4936 (N_4936,N_3565,N_3860);
nand U4937 (N_4937,N_3400,N_3545);
nand U4938 (N_4938,N_3940,N_3805);
or U4939 (N_4939,N_3720,N_3959);
and U4940 (N_4940,N_3992,N_3266);
nand U4941 (N_4941,N_3511,N_3577);
nand U4942 (N_4942,N_3591,N_3998);
nand U4943 (N_4943,N_3639,N_3458);
or U4944 (N_4944,N_3436,N_3287);
or U4945 (N_4945,N_3156,N_3607);
nor U4946 (N_4946,N_3226,N_3645);
or U4947 (N_4947,N_3746,N_3435);
nand U4948 (N_4948,N_3866,N_3900);
or U4949 (N_4949,N_3584,N_3690);
and U4950 (N_4950,N_3455,N_3965);
nand U4951 (N_4951,N_3819,N_3714);
xnor U4952 (N_4952,N_3122,N_3193);
and U4953 (N_4953,N_3573,N_3163);
or U4954 (N_4954,N_3773,N_3239);
or U4955 (N_4955,N_3440,N_3103);
nand U4956 (N_4956,N_3651,N_3694);
nor U4957 (N_4957,N_3858,N_3542);
and U4958 (N_4958,N_3555,N_3222);
nor U4959 (N_4959,N_3864,N_3935);
or U4960 (N_4960,N_3048,N_3533);
nand U4961 (N_4961,N_3444,N_3301);
and U4962 (N_4962,N_3595,N_3156);
xor U4963 (N_4963,N_3578,N_3444);
or U4964 (N_4964,N_3060,N_3788);
and U4965 (N_4965,N_3232,N_3723);
nand U4966 (N_4966,N_3356,N_3607);
nor U4967 (N_4967,N_3747,N_3863);
and U4968 (N_4968,N_3907,N_3291);
or U4969 (N_4969,N_3035,N_3974);
xor U4970 (N_4970,N_3802,N_3877);
or U4971 (N_4971,N_3772,N_3595);
nand U4972 (N_4972,N_3654,N_3869);
or U4973 (N_4973,N_3539,N_3584);
or U4974 (N_4974,N_3878,N_3687);
and U4975 (N_4975,N_3434,N_3384);
or U4976 (N_4976,N_3315,N_3701);
and U4977 (N_4977,N_3240,N_3027);
or U4978 (N_4978,N_3043,N_3654);
xor U4979 (N_4979,N_3014,N_3221);
xnor U4980 (N_4980,N_3950,N_3087);
xnor U4981 (N_4981,N_3650,N_3316);
nor U4982 (N_4982,N_3307,N_3944);
xor U4983 (N_4983,N_3364,N_3245);
and U4984 (N_4984,N_3600,N_3326);
nor U4985 (N_4985,N_3740,N_3955);
xnor U4986 (N_4986,N_3004,N_3661);
nand U4987 (N_4987,N_3280,N_3931);
and U4988 (N_4988,N_3964,N_3690);
nand U4989 (N_4989,N_3840,N_3436);
nor U4990 (N_4990,N_3665,N_3458);
xor U4991 (N_4991,N_3365,N_3900);
nor U4992 (N_4992,N_3533,N_3107);
nand U4993 (N_4993,N_3506,N_3353);
or U4994 (N_4994,N_3662,N_3027);
or U4995 (N_4995,N_3286,N_3849);
nand U4996 (N_4996,N_3762,N_3566);
nand U4997 (N_4997,N_3411,N_3955);
nand U4998 (N_4998,N_3268,N_3324);
nor U4999 (N_4999,N_3139,N_3176);
nor UO_0 (O_0,N_4648,N_4681);
xor UO_1 (O_1,N_4095,N_4838);
and UO_2 (O_2,N_4378,N_4694);
xnor UO_3 (O_3,N_4672,N_4373);
and UO_4 (O_4,N_4770,N_4527);
nand UO_5 (O_5,N_4932,N_4751);
nor UO_6 (O_6,N_4362,N_4978);
nand UO_7 (O_7,N_4936,N_4557);
nor UO_8 (O_8,N_4486,N_4660);
or UO_9 (O_9,N_4396,N_4997);
or UO_10 (O_10,N_4311,N_4586);
xor UO_11 (O_11,N_4068,N_4577);
or UO_12 (O_12,N_4277,N_4550);
xnor UO_13 (O_13,N_4430,N_4757);
and UO_14 (O_14,N_4031,N_4411);
or UO_15 (O_15,N_4344,N_4874);
nor UO_16 (O_16,N_4444,N_4609);
nand UO_17 (O_17,N_4627,N_4093);
and UO_18 (O_18,N_4345,N_4603);
and UO_19 (O_19,N_4136,N_4434);
and UO_20 (O_20,N_4002,N_4492);
nor UO_21 (O_21,N_4784,N_4354);
or UO_22 (O_22,N_4856,N_4295);
nor UO_23 (O_23,N_4005,N_4613);
nor UO_24 (O_24,N_4118,N_4591);
nor UO_25 (O_25,N_4866,N_4813);
or UO_26 (O_26,N_4168,N_4415);
or UO_27 (O_27,N_4961,N_4296);
nand UO_28 (O_28,N_4710,N_4072);
or UO_29 (O_29,N_4650,N_4985);
nor UO_30 (O_30,N_4477,N_4380);
or UO_31 (O_31,N_4771,N_4863);
or UO_32 (O_32,N_4760,N_4169);
and UO_33 (O_33,N_4558,N_4531);
nor UO_34 (O_34,N_4637,N_4696);
xnor UO_35 (O_35,N_4150,N_4292);
nor UO_36 (O_36,N_4593,N_4585);
nor UO_37 (O_37,N_4673,N_4858);
and UO_38 (O_38,N_4533,N_4748);
nand UO_39 (O_39,N_4847,N_4846);
or UO_40 (O_40,N_4250,N_4474);
or UO_41 (O_41,N_4667,N_4166);
and UO_42 (O_42,N_4922,N_4102);
and UO_43 (O_43,N_4879,N_4392);
nand UO_44 (O_44,N_4211,N_4049);
and UO_45 (O_45,N_4111,N_4853);
xor UO_46 (O_46,N_4205,N_4128);
and UO_47 (O_47,N_4404,N_4873);
nor UO_48 (O_48,N_4545,N_4820);
nand UO_49 (O_49,N_4491,N_4363);
and UO_50 (O_50,N_4259,N_4563);
nor UO_51 (O_51,N_4554,N_4151);
nor UO_52 (O_52,N_4543,N_4897);
and UO_53 (O_53,N_4566,N_4844);
xor UO_54 (O_54,N_4120,N_4747);
nor UO_55 (O_55,N_4061,N_4306);
or UO_56 (O_56,N_4130,N_4678);
nor UO_57 (O_57,N_4862,N_4440);
nor UO_58 (O_58,N_4335,N_4973);
nand UO_59 (O_59,N_4910,N_4903);
and UO_60 (O_60,N_4881,N_4716);
nand UO_61 (O_61,N_4749,N_4988);
or UO_62 (O_62,N_4562,N_4958);
nor UO_63 (O_63,N_4036,N_4200);
and UO_64 (O_64,N_4297,N_4916);
and UO_65 (O_65,N_4991,N_4447);
or UO_66 (O_66,N_4174,N_4657);
nand UO_67 (O_67,N_4412,N_4907);
or UO_68 (O_68,N_4471,N_4164);
nand UO_69 (O_69,N_4171,N_4647);
nand UO_70 (O_70,N_4876,N_4714);
nand UO_71 (O_71,N_4946,N_4548);
xor UO_72 (O_72,N_4407,N_4132);
and UO_73 (O_73,N_4022,N_4811);
and UO_74 (O_74,N_4975,N_4754);
or UO_75 (O_75,N_4940,N_4564);
and UO_76 (O_76,N_4459,N_4107);
or UO_77 (O_77,N_4455,N_4674);
and UO_78 (O_78,N_4268,N_4454);
and UO_79 (O_79,N_4604,N_4112);
or UO_80 (O_80,N_4056,N_4312);
xor UO_81 (O_81,N_4885,N_4789);
nand UO_82 (O_82,N_4688,N_4425);
nor UO_83 (O_83,N_4691,N_4623);
and UO_84 (O_84,N_4815,N_4235);
xor UO_85 (O_85,N_4887,N_4242);
nor UO_86 (O_86,N_4453,N_4030);
and UO_87 (O_87,N_4305,N_4155);
nor UO_88 (O_88,N_4572,N_4989);
and UO_89 (O_89,N_4986,N_4347);
nand UO_90 (O_90,N_4639,N_4385);
and UO_91 (O_91,N_4513,N_4928);
nor UO_92 (O_92,N_4096,N_4063);
and UO_93 (O_93,N_4442,N_4202);
or UO_94 (O_94,N_4935,N_4765);
nand UO_95 (O_95,N_4027,N_4369);
or UO_96 (O_96,N_4656,N_4568);
nor UO_97 (O_97,N_4663,N_4941);
or UO_98 (O_98,N_4618,N_4993);
nand UO_99 (O_99,N_4877,N_4502);
or UO_100 (O_100,N_4511,N_4617);
and UO_101 (O_101,N_4343,N_4619);
nand UO_102 (O_102,N_4826,N_4353);
nor UO_103 (O_103,N_4630,N_4854);
or UO_104 (O_104,N_4512,N_4526);
nand UO_105 (O_105,N_4769,N_4954);
xor UO_106 (O_106,N_4732,N_4115);
and UO_107 (O_107,N_4675,N_4193);
or UO_108 (O_108,N_4508,N_4034);
nand UO_109 (O_109,N_4350,N_4998);
nand UO_110 (O_110,N_4021,N_4349);
xnor UO_111 (O_111,N_4073,N_4341);
nand UO_112 (O_112,N_4763,N_4702);
and UO_113 (O_113,N_4951,N_4984);
xor UO_114 (O_114,N_4949,N_4795);
and UO_115 (O_115,N_4338,N_4701);
or UO_116 (O_116,N_4544,N_4942);
nand UO_117 (O_117,N_4417,N_4255);
nand UO_118 (O_118,N_4651,N_4246);
or UO_119 (O_119,N_4286,N_4836);
nor UO_120 (O_120,N_4461,N_4230);
and UO_121 (O_121,N_4003,N_4231);
and UO_122 (O_122,N_4995,N_4759);
nand UO_123 (O_123,N_4180,N_4181);
and UO_124 (O_124,N_4328,N_4192);
and UO_125 (O_125,N_4662,N_4368);
xnor UO_126 (O_126,N_4573,N_4009);
nand UO_127 (O_127,N_4488,N_4364);
nand UO_128 (O_128,N_4773,N_4621);
nor UO_129 (O_129,N_4176,N_4094);
nand UO_130 (O_130,N_4004,N_4225);
and UO_131 (O_131,N_4584,N_4767);
xor UO_132 (O_132,N_4157,N_4608);
or UO_133 (O_133,N_4865,N_4291);
nand UO_134 (O_134,N_4848,N_4695);
nand UO_135 (O_135,N_4962,N_4163);
nand UO_136 (O_136,N_4708,N_4046);
xnor UO_137 (O_137,N_4085,N_4104);
and UO_138 (O_138,N_4421,N_4287);
or UO_139 (O_139,N_4105,N_4148);
nand UO_140 (O_140,N_4869,N_4933);
xnor UO_141 (O_141,N_4456,N_4926);
nor UO_142 (O_142,N_4886,N_4902);
and UO_143 (O_143,N_4274,N_4642);
or UO_144 (O_144,N_4484,N_4821);
and UO_145 (O_145,N_4616,N_4629);
nor UO_146 (O_146,N_4334,N_4834);
nor UO_147 (O_147,N_4882,N_4390);
xnor UO_148 (O_148,N_4742,N_4361);
nor UO_149 (O_149,N_4515,N_4801);
and UO_150 (O_150,N_4017,N_4685);
nand UO_151 (O_151,N_4794,N_4992);
xor UO_152 (O_152,N_4601,N_4251);
or UO_153 (O_153,N_4313,N_4451);
or UO_154 (O_154,N_4346,N_4920);
and UO_155 (O_155,N_4532,N_4080);
nor UO_156 (O_156,N_4092,N_4842);
and UO_157 (O_157,N_4314,N_4387);
nand UO_158 (O_158,N_4536,N_4495);
or UO_159 (O_159,N_4670,N_4735);
nor UO_160 (O_160,N_4241,N_4374);
and UO_161 (O_161,N_4140,N_4399);
nor UO_162 (O_162,N_4048,N_4884);
and UO_163 (O_163,N_4780,N_4234);
and UO_164 (O_164,N_4283,N_4638);
or UO_165 (O_165,N_4275,N_4414);
nor UO_166 (O_166,N_4590,N_4066);
nor UO_167 (O_167,N_4809,N_4327);
and UO_168 (O_168,N_4693,N_4252);
and UO_169 (O_169,N_4909,N_4805);
or UO_170 (O_170,N_4719,N_4429);
nand UO_171 (O_171,N_4135,N_4162);
nor UO_172 (O_172,N_4041,N_4028);
nor UO_173 (O_173,N_4436,N_4462);
nand UO_174 (O_174,N_4868,N_4952);
and UO_175 (O_175,N_4731,N_4064);
nand UO_176 (O_176,N_4070,N_4724);
xor UO_177 (O_177,N_4139,N_4875);
or UO_178 (O_178,N_4173,N_4547);
and UO_179 (O_179,N_4426,N_4786);
or UO_180 (O_180,N_4463,N_4658);
nor UO_181 (O_181,N_4925,N_4706);
xor UO_182 (O_182,N_4615,N_4131);
and UO_183 (O_183,N_4600,N_4400);
xnor UO_184 (O_184,N_4043,N_4517);
nor UO_185 (O_185,N_4290,N_4753);
xor UO_186 (O_186,N_4703,N_4199);
nor UO_187 (O_187,N_4700,N_4595);
nor UO_188 (O_188,N_4582,N_4071);
and UO_189 (O_189,N_4535,N_4686);
or UO_190 (O_190,N_4445,N_4011);
nand UO_191 (O_191,N_4644,N_4203);
or UO_192 (O_192,N_4342,N_4266);
nor UO_193 (O_193,N_4915,N_4258);
xnor UO_194 (O_194,N_4232,N_4216);
or UO_195 (O_195,N_4010,N_4556);
and UO_196 (O_196,N_4684,N_4037);
and UO_197 (O_197,N_4546,N_4683);
or UO_198 (O_198,N_4588,N_4911);
nand UO_199 (O_199,N_4395,N_4124);
and UO_200 (O_200,N_4496,N_4161);
nor UO_201 (O_201,N_4469,N_4186);
and UO_202 (O_202,N_4740,N_4483);
nor UO_203 (O_203,N_4081,N_4861);
or UO_204 (O_204,N_4552,N_4967);
nor UO_205 (O_205,N_4624,N_4360);
nor UO_206 (O_206,N_4359,N_4806);
nand UO_207 (O_207,N_4825,N_4059);
and UO_208 (O_208,N_4100,N_4109);
or UO_209 (O_209,N_4299,N_4315);
nor UO_210 (O_210,N_4501,N_4116);
or UO_211 (O_211,N_4800,N_4236);
nand UO_212 (O_212,N_4698,N_4507);
nor UO_213 (O_213,N_4626,N_4398);
or UO_214 (O_214,N_4466,N_4792);
nand UO_215 (O_215,N_4224,N_4725);
and UO_216 (O_216,N_4504,N_4244);
and UO_217 (O_217,N_4778,N_4366);
or UO_218 (O_218,N_4752,N_4388);
nand UO_219 (O_219,N_4781,N_4938);
and UO_220 (O_220,N_4728,N_4802);
nor UO_221 (O_221,N_4271,N_4923);
nand UO_222 (O_222,N_4367,N_4518);
xor UO_223 (O_223,N_4288,N_4810);
and UO_224 (O_224,N_4717,N_4891);
or UO_225 (O_225,N_4709,N_4999);
nand UO_226 (O_226,N_4665,N_4147);
and UO_227 (O_227,N_4713,N_4035);
nand UO_228 (O_228,N_4721,N_4329);
nand UO_229 (O_229,N_4798,N_4652);
and UO_230 (O_230,N_4807,N_4676);
nand UO_231 (O_231,N_4079,N_4974);
nand UO_232 (O_232,N_4464,N_4075);
nor UO_233 (O_233,N_4929,N_4405);
and UO_234 (O_234,N_4247,N_4537);
and UO_235 (O_235,N_4175,N_4646);
nor UO_236 (O_236,N_4253,N_4587);
and UO_237 (O_237,N_4029,N_4906);
and UO_238 (O_238,N_4705,N_4260);
and UO_239 (O_239,N_4895,N_4052);
nor UO_240 (O_240,N_4594,N_4014);
or UO_241 (O_241,N_4835,N_4276);
nand UO_242 (O_242,N_4379,N_4177);
nor UO_243 (O_243,N_4076,N_4293);
or UO_244 (O_244,N_4113,N_4322);
nand UO_245 (O_245,N_4823,N_4254);
nor UO_246 (O_246,N_4722,N_4871);
xnor UO_247 (O_247,N_4013,N_4302);
nor UO_248 (O_248,N_4777,N_4976);
or UO_249 (O_249,N_4238,N_4183);
or UO_250 (O_250,N_4032,N_4943);
nand UO_251 (O_251,N_4529,N_4256);
nor UO_252 (O_252,N_4233,N_4808);
and UO_253 (O_253,N_4715,N_4837);
or UO_254 (O_254,N_4240,N_4878);
or UO_255 (O_255,N_4279,N_4448);
and UO_256 (O_256,N_4723,N_4457);
xor UO_257 (O_257,N_4332,N_4990);
nor UO_258 (O_258,N_4620,N_4937);
nand UO_259 (O_259,N_4382,N_4204);
and UO_260 (O_260,N_4077,N_4084);
or UO_261 (O_261,N_4812,N_4160);
and UO_262 (O_262,N_4850,N_4864);
and UO_263 (O_263,N_4833,N_4352);
nor UO_264 (O_264,N_4718,N_4078);
xor UO_265 (O_265,N_4308,N_4386);
or UO_266 (O_266,N_4088,N_4523);
and UO_267 (O_267,N_4487,N_4741);
xor UO_268 (O_268,N_4316,N_4559);
nor UO_269 (O_269,N_4223,N_4972);
nor UO_270 (O_270,N_4679,N_4310);
nand UO_271 (O_271,N_4479,N_4596);
or UO_272 (O_272,N_4008,N_4402);
and UO_273 (O_273,N_4631,N_4215);
nor UO_274 (O_274,N_4282,N_4839);
nand UO_275 (O_275,N_4439,N_4569);
and UO_276 (O_276,N_4510,N_4065);
or UO_277 (O_277,N_4790,N_4924);
xnor UO_278 (O_278,N_4133,N_4237);
and UO_279 (O_279,N_4889,N_4649);
nor UO_280 (O_280,N_4044,N_4278);
nand UO_281 (O_281,N_4689,N_4913);
nand UO_282 (O_282,N_4783,N_4581);
or UO_283 (O_283,N_4191,N_4610);
nand UO_284 (O_284,N_4787,N_4141);
nand UO_285 (O_285,N_4977,N_4045);
and UO_286 (O_286,N_4401,N_4738);
and UO_287 (O_287,N_4154,N_4473);
and UO_288 (O_288,N_4058,N_4890);
nand UO_289 (O_289,N_4475,N_4643);
nand UO_290 (O_290,N_4108,N_4567);
nor UO_291 (O_291,N_4121,N_4153);
and UO_292 (O_292,N_4746,N_4996);
nor UO_293 (O_293,N_4579,N_4745);
nand UO_294 (O_294,N_4730,N_4641);
and UO_295 (O_295,N_4712,N_4653);
nand UO_296 (O_296,N_4827,N_4598);
and UO_297 (O_297,N_4365,N_4356);
or UO_298 (O_298,N_4855,N_4119);
or UO_299 (O_299,N_4575,N_4053);
nand UO_300 (O_300,N_4082,N_4188);
nor UO_301 (O_301,N_4318,N_4570);
xor UO_302 (O_302,N_4525,N_4565);
and UO_303 (O_303,N_4272,N_4633);
nor UO_304 (O_304,N_4772,N_4336);
and UO_305 (O_305,N_4384,N_4146);
nor UO_306 (O_306,N_4489,N_4521);
and UO_307 (O_307,N_4178,N_4645);
or UO_308 (O_308,N_4403,N_4764);
nor UO_309 (O_309,N_4538,N_4602);
nand UO_310 (O_310,N_4899,N_4321);
nor UO_311 (O_311,N_4106,N_4828);
and UO_312 (O_312,N_4138,N_4829);
nand UO_313 (O_313,N_4023,N_4098);
xnor UO_314 (O_314,N_4389,N_4273);
xor UO_315 (O_315,N_4880,N_4142);
nor UO_316 (O_316,N_4228,N_4007);
nor UO_317 (O_317,N_4019,N_4050);
or UO_318 (O_318,N_4607,N_4782);
or UO_319 (O_319,N_4397,N_4062);
nor UO_320 (O_320,N_4468,N_4213);
xnor UO_321 (O_321,N_4265,N_4020);
or UO_322 (O_322,N_4331,N_4497);
nand UO_323 (O_323,N_4428,N_4090);
and UO_324 (O_324,N_4300,N_4210);
nand UO_325 (O_325,N_4774,N_4371);
xnor UO_326 (O_326,N_4091,N_4033);
or UO_327 (O_327,N_4219,N_4611);
xor UO_328 (O_328,N_4304,N_4896);
or UO_329 (O_329,N_4289,N_4221);
nor UO_330 (O_330,N_4632,N_4391);
and UO_331 (O_331,N_4971,N_4214);
xnor UO_332 (O_332,N_4947,N_4883);
or UO_333 (O_333,N_4982,N_4831);
xnor UO_334 (O_334,N_4067,N_4797);
nor UO_335 (O_335,N_4519,N_4432);
nor UO_336 (O_336,N_4539,N_4578);
xor UO_337 (O_337,N_4494,N_4851);
and UO_338 (O_338,N_4955,N_4592);
and UO_339 (O_339,N_4087,N_4097);
nor UO_340 (O_340,N_4888,N_4372);
xnor UO_341 (O_341,N_4325,N_4055);
or UO_342 (O_342,N_4394,N_4375);
or UO_343 (O_343,N_4319,N_4918);
and UO_344 (O_344,N_4571,N_4083);
and UO_345 (O_345,N_4981,N_4420);
and UO_346 (O_346,N_4930,N_4172);
or UO_347 (O_347,N_4931,N_4499);
and UO_348 (O_348,N_4326,N_4452);
nand UO_349 (O_349,N_4666,N_4994);
or UO_350 (O_350,N_4422,N_4498);
nor UO_351 (O_351,N_4743,N_4418);
and UO_352 (O_352,N_4478,N_4333);
or UO_353 (O_353,N_4822,N_4220);
nand UO_354 (O_354,N_4799,N_4330);
and UO_355 (O_355,N_4476,N_4793);
or UO_356 (O_356,N_4419,N_4264);
nand UO_357 (O_357,N_4229,N_4485);
nand UO_358 (O_358,N_4859,N_4317);
nor UO_359 (O_359,N_4553,N_4038);
nand UO_360 (O_360,N_4857,N_4016);
nand UO_361 (O_361,N_4281,N_4791);
nor UO_362 (O_362,N_4860,N_4257);
or UO_363 (O_363,N_4692,N_4549);
nor UO_364 (O_364,N_4503,N_4761);
nand UO_365 (O_365,N_4189,N_4775);
nand UO_366 (O_366,N_4768,N_4437);
nor UO_367 (O_367,N_4054,N_4506);
or UO_368 (O_368,N_4758,N_4149);
or UO_369 (O_369,N_4818,N_4589);
nor UO_370 (O_370,N_4661,N_4438);
or UO_371 (O_371,N_4493,N_4001);
nor UO_372 (O_372,N_4198,N_4788);
or UO_373 (O_373,N_4195,N_4103);
and UO_374 (O_374,N_4561,N_4441);
and UO_375 (O_375,N_4480,N_4423);
nand UO_376 (O_376,N_4534,N_4309);
and UO_377 (O_377,N_4167,N_4816);
nand UO_378 (O_378,N_4051,N_4892);
nand UO_379 (O_379,N_4901,N_4424);
nor UO_380 (O_380,N_4524,N_4249);
or UO_381 (O_381,N_4152,N_4280);
nand UO_382 (O_382,N_4406,N_4298);
nand UO_383 (O_383,N_4129,N_4682);
nor UO_384 (O_384,N_4840,N_4948);
or UO_385 (O_385,N_4697,N_4024);
nor UO_386 (O_386,N_4830,N_4733);
and UO_387 (O_387,N_4750,N_4416);
and UO_388 (O_388,N_4381,N_4190);
nor UO_389 (O_389,N_4912,N_4987);
and UO_390 (O_390,N_4599,N_4137);
and UO_391 (O_391,N_4516,N_4222);
nor UO_392 (O_392,N_4443,N_4006);
or UO_393 (O_393,N_4057,N_4606);
and UO_394 (O_394,N_4000,N_4184);
nor UO_395 (O_395,N_4727,N_4212);
or UO_396 (O_396,N_4597,N_4196);
or UO_397 (O_397,N_4217,N_4377);
nand UO_398 (O_398,N_4458,N_4921);
nor UO_399 (O_399,N_4194,N_4324);
and UO_400 (O_400,N_4509,N_4814);
nand UO_401 (O_401,N_4284,N_4560);
nand UO_402 (O_402,N_4867,N_4159);
nand UO_403 (O_403,N_4207,N_4872);
or UO_404 (O_404,N_4270,N_4209);
nand UO_405 (O_405,N_4522,N_4450);
and UO_406 (O_406,N_4408,N_4025);
or UO_407 (O_407,N_4126,N_4541);
or UO_408 (O_408,N_4968,N_4690);
nor UO_409 (O_409,N_4845,N_4435);
or UO_410 (O_410,N_4677,N_4736);
and UO_411 (O_411,N_4762,N_4980);
nand UO_412 (O_412,N_4785,N_4655);
or UO_413 (O_413,N_4680,N_4945);
or UO_414 (O_414,N_4514,N_4301);
and UO_415 (O_415,N_4303,N_4294);
and UO_416 (O_416,N_4894,N_4500);
and UO_417 (O_417,N_4893,N_4614);
and UO_418 (O_418,N_4963,N_4843);
or UO_419 (O_419,N_4117,N_4635);
or UO_420 (O_420,N_4383,N_4470);
or UO_421 (O_421,N_4012,N_4239);
nand UO_422 (O_422,N_4069,N_4970);
nor UO_423 (O_423,N_4612,N_4427);
or UO_424 (O_424,N_4227,N_4956);
and UO_425 (O_425,N_4852,N_4433);
nor UO_426 (O_426,N_4208,N_4711);
nand UO_427 (O_427,N_4099,N_4393);
and UO_428 (O_428,N_4039,N_4622);
or UO_429 (O_429,N_4520,N_4900);
nand UO_430 (O_430,N_4755,N_4979);
nand UO_431 (O_431,N_4245,N_4530);
nor UO_432 (O_432,N_4320,N_4355);
and UO_433 (O_433,N_4634,N_4348);
nand UO_434 (O_434,N_4934,N_4086);
or UO_435 (O_435,N_4218,N_4449);
nand UO_436 (O_436,N_4156,N_4123);
or UO_437 (O_437,N_4026,N_4720);
nor UO_438 (O_438,N_4351,N_4744);
xnor UO_439 (O_439,N_4505,N_4074);
and UO_440 (O_440,N_4766,N_4944);
nor UO_441 (O_441,N_4243,N_4472);
xor UO_442 (O_442,N_4144,N_4576);
and UO_443 (O_443,N_4410,N_4914);
nand UO_444 (O_444,N_4261,N_4358);
xnor UO_445 (O_445,N_4849,N_4699);
and UO_446 (O_446,N_4125,N_4267);
and UO_447 (O_447,N_4015,N_4555);
nand UO_448 (O_448,N_4654,N_4370);
and UO_449 (O_449,N_4089,N_4182);
nor UO_450 (O_450,N_4898,N_4340);
nor UO_451 (O_451,N_4803,N_4659);
nand UO_452 (O_452,N_4804,N_4460);
nand UO_453 (O_453,N_4170,N_4966);
or UO_454 (O_454,N_4158,N_4841);
xor UO_455 (O_455,N_4542,N_4285);
nor UO_456 (O_456,N_4490,N_4551);
nand UO_457 (O_457,N_4114,N_4756);
nand UO_458 (O_458,N_4707,N_4465);
or UO_459 (O_459,N_4269,N_4939);
or UO_460 (O_460,N_4047,N_4040);
or UO_461 (O_461,N_4263,N_4337);
and UO_462 (O_462,N_4671,N_4669);
or UO_463 (O_463,N_4197,N_4323);
or UO_464 (O_464,N_4904,N_4817);
nor UO_465 (O_465,N_4101,N_4165);
xor UO_466 (O_466,N_4376,N_4965);
nand UO_467 (O_467,N_4969,N_4739);
nor UO_468 (O_468,N_4226,N_4145);
and UO_469 (O_469,N_4640,N_4919);
or UO_470 (O_470,N_4307,N_4467);
and UO_471 (O_471,N_4134,N_4201);
and UO_472 (O_472,N_4110,N_4580);
nand UO_473 (O_473,N_4179,N_4905);
or UO_474 (O_474,N_4583,N_4908);
nor UO_475 (O_475,N_4668,N_4636);
nor UO_476 (O_476,N_4953,N_4431);
nand UO_477 (O_477,N_4339,N_4018);
and UO_478 (O_478,N_4481,N_4917);
nor UO_479 (O_479,N_4413,N_4574);
xnor UO_480 (O_480,N_4779,N_4737);
nand UO_481 (O_481,N_4060,N_4664);
or UO_482 (O_482,N_4960,N_4687);
xor UO_483 (O_483,N_4605,N_4819);
xnor UO_484 (O_484,N_4964,N_4776);
or UO_485 (O_485,N_4950,N_4983);
or UO_486 (O_486,N_4127,N_4528);
or UO_487 (O_487,N_4628,N_4957);
and UO_488 (O_488,N_4409,N_4959);
and UO_489 (O_489,N_4704,N_4185);
xnor UO_490 (O_490,N_4446,N_4143);
xor UO_491 (O_491,N_4357,N_4870);
nor UO_492 (O_492,N_4262,N_4734);
and UO_493 (O_493,N_4122,N_4482);
nor UO_494 (O_494,N_4729,N_4832);
nand UO_495 (O_495,N_4726,N_4248);
nor UO_496 (O_496,N_4540,N_4625);
nor UO_497 (O_497,N_4824,N_4206);
nor UO_498 (O_498,N_4042,N_4796);
and UO_499 (O_499,N_4927,N_4187);
nor UO_500 (O_500,N_4717,N_4454);
or UO_501 (O_501,N_4809,N_4964);
nor UO_502 (O_502,N_4245,N_4986);
or UO_503 (O_503,N_4272,N_4733);
nor UO_504 (O_504,N_4806,N_4712);
nand UO_505 (O_505,N_4741,N_4696);
or UO_506 (O_506,N_4347,N_4251);
or UO_507 (O_507,N_4983,N_4004);
xnor UO_508 (O_508,N_4488,N_4419);
or UO_509 (O_509,N_4137,N_4951);
nor UO_510 (O_510,N_4239,N_4188);
nand UO_511 (O_511,N_4714,N_4650);
and UO_512 (O_512,N_4755,N_4829);
nor UO_513 (O_513,N_4514,N_4730);
or UO_514 (O_514,N_4536,N_4802);
nand UO_515 (O_515,N_4411,N_4730);
and UO_516 (O_516,N_4628,N_4311);
nand UO_517 (O_517,N_4530,N_4730);
and UO_518 (O_518,N_4303,N_4621);
nor UO_519 (O_519,N_4165,N_4779);
nand UO_520 (O_520,N_4843,N_4998);
or UO_521 (O_521,N_4542,N_4920);
and UO_522 (O_522,N_4707,N_4155);
nor UO_523 (O_523,N_4004,N_4492);
and UO_524 (O_524,N_4769,N_4519);
and UO_525 (O_525,N_4527,N_4044);
and UO_526 (O_526,N_4737,N_4749);
or UO_527 (O_527,N_4235,N_4410);
and UO_528 (O_528,N_4187,N_4009);
or UO_529 (O_529,N_4703,N_4431);
and UO_530 (O_530,N_4208,N_4643);
and UO_531 (O_531,N_4874,N_4813);
nor UO_532 (O_532,N_4802,N_4828);
and UO_533 (O_533,N_4185,N_4301);
nor UO_534 (O_534,N_4670,N_4793);
xor UO_535 (O_535,N_4879,N_4652);
or UO_536 (O_536,N_4372,N_4452);
and UO_537 (O_537,N_4895,N_4694);
and UO_538 (O_538,N_4637,N_4663);
nor UO_539 (O_539,N_4364,N_4056);
or UO_540 (O_540,N_4035,N_4862);
nor UO_541 (O_541,N_4521,N_4272);
and UO_542 (O_542,N_4250,N_4366);
nor UO_543 (O_543,N_4148,N_4873);
or UO_544 (O_544,N_4483,N_4844);
or UO_545 (O_545,N_4359,N_4488);
or UO_546 (O_546,N_4135,N_4417);
and UO_547 (O_547,N_4496,N_4328);
and UO_548 (O_548,N_4282,N_4945);
nor UO_549 (O_549,N_4570,N_4503);
nand UO_550 (O_550,N_4108,N_4713);
nand UO_551 (O_551,N_4170,N_4634);
nand UO_552 (O_552,N_4671,N_4330);
nor UO_553 (O_553,N_4889,N_4705);
or UO_554 (O_554,N_4701,N_4509);
nor UO_555 (O_555,N_4690,N_4252);
or UO_556 (O_556,N_4430,N_4012);
nor UO_557 (O_557,N_4927,N_4257);
xor UO_558 (O_558,N_4054,N_4902);
xnor UO_559 (O_559,N_4612,N_4567);
nand UO_560 (O_560,N_4543,N_4703);
nor UO_561 (O_561,N_4088,N_4014);
nor UO_562 (O_562,N_4104,N_4841);
nand UO_563 (O_563,N_4177,N_4621);
and UO_564 (O_564,N_4197,N_4347);
or UO_565 (O_565,N_4604,N_4172);
or UO_566 (O_566,N_4982,N_4600);
nor UO_567 (O_567,N_4470,N_4283);
or UO_568 (O_568,N_4095,N_4374);
nand UO_569 (O_569,N_4181,N_4293);
or UO_570 (O_570,N_4821,N_4210);
nor UO_571 (O_571,N_4878,N_4379);
nor UO_572 (O_572,N_4641,N_4414);
nor UO_573 (O_573,N_4040,N_4758);
nand UO_574 (O_574,N_4036,N_4707);
nor UO_575 (O_575,N_4710,N_4191);
nand UO_576 (O_576,N_4083,N_4635);
xnor UO_577 (O_577,N_4436,N_4429);
nor UO_578 (O_578,N_4990,N_4858);
nand UO_579 (O_579,N_4545,N_4054);
or UO_580 (O_580,N_4569,N_4678);
and UO_581 (O_581,N_4268,N_4491);
nand UO_582 (O_582,N_4088,N_4529);
and UO_583 (O_583,N_4883,N_4018);
xor UO_584 (O_584,N_4759,N_4128);
or UO_585 (O_585,N_4026,N_4993);
and UO_586 (O_586,N_4427,N_4511);
nor UO_587 (O_587,N_4452,N_4070);
nand UO_588 (O_588,N_4630,N_4678);
xnor UO_589 (O_589,N_4158,N_4301);
nand UO_590 (O_590,N_4031,N_4063);
nand UO_591 (O_591,N_4838,N_4971);
or UO_592 (O_592,N_4831,N_4030);
or UO_593 (O_593,N_4504,N_4262);
xor UO_594 (O_594,N_4237,N_4348);
or UO_595 (O_595,N_4889,N_4141);
nor UO_596 (O_596,N_4584,N_4280);
or UO_597 (O_597,N_4569,N_4735);
xnor UO_598 (O_598,N_4672,N_4044);
xnor UO_599 (O_599,N_4404,N_4007);
and UO_600 (O_600,N_4168,N_4553);
and UO_601 (O_601,N_4666,N_4124);
or UO_602 (O_602,N_4934,N_4096);
and UO_603 (O_603,N_4715,N_4683);
and UO_604 (O_604,N_4033,N_4448);
nor UO_605 (O_605,N_4472,N_4916);
nand UO_606 (O_606,N_4560,N_4761);
or UO_607 (O_607,N_4008,N_4228);
or UO_608 (O_608,N_4364,N_4668);
or UO_609 (O_609,N_4936,N_4138);
or UO_610 (O_610,N_4331,N_4083);
nor UO_611 (O_611,N_4792,N_4317);
nor UO_612 (O_612,N_4334,N_4782);
and UO_613 (O_613,N_4212,N_4169);
nand UO_614 (O_614,N_4390,N_4660);
nand UO_615 (O_615,N_4152,N_4391);
nand UO_616 (O_616,N_4183,N_4381);
nor UO_617 (O_617,N_4822,N_4052);
xor UO_618 (O_618,N_4114,N_4031);
and UO_619 (O_619,N_4451,N_4781);
and UO_620 (O_620,N_4934,N_4595);
nand UO_621 (O_621,N_4249,N_4929);
and UO_622 (O_622,N_4650,N_4482);
or UO_623 (O_623,N_4125,N_4536);
xor UO_624 (O_624,N_4761,N_4668);
and UO_625 (O_625,N_4228,N_4016);
or UO_626 (O_626,N_4725,N_4345);
xnor UO_627 (O_627,N_4929,N_4610);
nor UO_628 (O_628,N_4855,N_4918);
xnor UO_629 (O_629,N_4902,N_4791);
nor UO_630 (O_630,N_4544,N_4329);
nand UO_631 (O_631,N_4957,N_4975);
nand UO_632 (O_632,N_4166,N_4589);
or UO_633 (O_633,N_4625,N_4016);
nor UO_634 (O_634,N_4685,N_4561);
nor UO_635 (O_635,N_4248,N_4041);
or UO_636 (O_636,N_4401,N_4979);
nor UO_637 (O_637,N_4188,N_4910);
or UO_638 (O_638,N_4790,N_4182);
nand UO_639 (O_639,N_4204,N_4186);
and UO_640 (O_640,N_4379,N_4843);
nor UO_641 (O_641,N_4402,N_4410);
nand UO_642 (O_642,N_4627,N_4034);
or UO_643 (O_643,N_4289,N_4762);
and UO_644 (O_644,N_4586,N_4061);
nor UO_645 (O_645,N_4075,N_4995);
or UO_646 (O_646,N_4366,N_4591);
xor UO_647 (O_647,N_4931,N_4316);
and UO_648 (O_648,N_4381,N_4016);
or UO_649 (O_649,N_4331,N_4134);
and UO_650 (O_650,N_4924,N_4317);
nand UO_651 (O_651,N_4432,N_4471);
or UO_652 (O_652,N_4045,N_4958);
or UO_653 (O_653,N_4448,N_4218);
or UO_654 (O_654,N_4824,N_4479);
or UO_655 (O_655,N_4302,N_4966);
nor UO_656 (O_656,N_4542,N_4166);
nand UO_657 (O_657,N_4027,N_4596);
nor UO_658 (O_658,N_4544,N_4189);
nor UO_659 (O_659,N_4613,N_4451);
nor UO_660 (O_660,N_4698,N_4263);
or UO_661 (O_661,N_4123,N_4879);
and UO_662 (O_662,N_4558,N_4185);
and UO_663 (O_663,N_4825,N_4729);
nor UO_664 (O_664,N_4776,N_4847);
nand UO_665 (O_665,N_4303,N_4959);
nand UO_666 (O_666,N_4580,N_4361);
and UO_667 (O_667,N_4792,N_4401);
nor UO_668 (O_668,N_4992,N_4677);
and UO_669 (O_669,N_4073,N_4782);
or UO_670 (O_670,N_4942,N_4029);
or UO_671 (O_671,N_4826,N_4854);
nor UO_672 (O_672,N_4095,N_4479);
nor UO_673 (O_673,N_4383,N_4084);
and UO_674 (O_674,N_4804,N_4099);
and UO_675 (O_675,N_4276,N_4008);
and UO_676 (O_676,N_4658,N_4579);
nand UO_677 (O_677,N_4624,N_4696);
nand UO_678 (O_678,N_4137,N_4031);
nand UO_679 (O_679,N_4114,N_4152);
or UO_680 (O_680,N_4769,N_4826);
and UO_681 (O_681,N_4869,N_4980);
or UO_682 (O_682,N_4296,N_4624);
or UO_683 (O_683,N_4710,N_4114);
and UO_684 (O_684,N_4959,N_4834);
nor UO_685 (O_685,N_4533,N_4866);
and UO_686 (O_686,N_4087,N_4151);
or UO_687 (O_687,N_4478,N_4406);
xnor UO_688 (O_688,N_4275,N_4089);
nor UO_689 (O_689,N_4048,N_4361);
and UO_690 (O_690,N_4271,N_4960);
or UO_691 (O_691,N_4685,N_4207);
xnor UO_692 (O_692,N_4656,N_4983);
nand UO_693 (O_693,N_4295,N_4327);
or UO_694 (O_694,N_4709,N_4936);
xnor UO_695 (O_695,N_4929,N_4151);
nand UO_696 (O_696,N_4737,N_4147);
and UO_697 (O_697,N_4319,N_4848);
nor UO_698 (O_698,N_4116,N_4879);
nand UO_699 (O_699,N_4578,N_4626);
or UO_700 (O_700,N_4074,N_4410);
nor UO_701 (O_701,N_4720,N_4441);
or UO_702 (O_702,N_4542,N_4437);
xnor UO_703 (O_703,N_4514,N_4405);
nand UO_704 (O_704,N_4744,N_4169);
nand UO_705 (O_705,N_4766,N_4262);
nand UO_706 (O_706,N_4013,N_4114);
and UO_707 (O_707,N_4570,N_4294);
or UO_708 (O_708,N_4779,N_4671);
nand UO_709 (O_709,N_4713,N_4357);
and UO_710 (O_710,N_4205,N_4046);
nand UO_711 (O_711,N_4800,N_4761);
nand UO_712 (O_712,N_4960,N_4868);
xor UO_713 (O_713,N_4677,N_4755);
nor UO_714 (O_714,N_4006,N_4124);
nand UO_715 (O_715,N_4003,N_4919);
nor UO_716 (O_716,N_4678,N_4375);
xnor UO_717 (O_717,N_4888,N_4601);
nand UO_718 (O_718,N_4467,N_4960);
nor UO_719 (O_719,N_4729,N_4807);
nor UO_720 (O_720,N_4648,N_4999);
nor UO_721 (O_721,N_4025,N_4589);
nand UO_722 (O_722,N_4917,N_4292);
or UO_723 (O_723,N_4010,N_4728);
nand UO_724 (O_724,N_4112,N_4656);
nand UO_725 (O_725,N_4126,N_4891);
or UO_726 (O_726,N_4555,N_4328);
xor UO_727 (O_727,N_4488,N_4138);
and UO_728 (O_728,N_4392,N_4868);
or UO_729 (O_729,N_4222,N_4831);
xnor UO_730 (O_730,N_4636,N_4805);
or UO_731 (O_731,N_4130,N_4191);
or UO_732 (O_732,N_4032,N_4699);
nor UO_733 (O_733,N_4490,N_4017);
nor UO_734 (O_734,N_4969,N_4549);
nand UO_735 (O_735,N_4107,N_4410);
nor UO_736 (O_736,N_4989,N_4560);
or UO_737 (O_737,N_4175,N_4777);
and UO_738 (O_738,N_4494,N_4714);
or UO_739 (O_739,N_4997,N_4909);
or UO_740 (O_740,N_4533,N_4198);
or UO_741 (O_741,N_4502,N_4359);
nand UO_742 (O_742,N_4829,N_4492);
and UO_743 (O_743,N_4163,N_4825);
nand UO_744 (O_744,N_4113,N_4634);
nand UO_745 (O_745,N_4263,N_4666);
nor UO_746 (O_746,N_4050,N_4386);
and UO_747 (O_747,N_4557,N_4799);
nand UO_748 (O_748,N_4635,N_4983);
or UO_749 (O_749,N_4470,N_4989);
and UO_750 (O_750,N_4053,N_4088);
or UO_751 (O_751,N_4279,N_4731);
nor UO_752 (O_752,N_4370,N_4512);
nand UO_753 (O_753,N_4417,N_4033);
nor UO_754 (O_754,N_4274,N_4577);
and UO_755 (O_755,N_4444,N_4792);
or UO_756 (O_756,N_4713,N_4189);
xnor UO_757 (O_757,N_4501,N_4010);
or UO_758 (O_758,N_4543,N_4360);
nand UO_759 (O_759,N_4895,N_4720);
and UO_760 (O_760,N_4168,N_4738);
and UO_761 (O_761,N_4570,N_4792);
and UO_762 (O_762,N_4923,N_4181);
and UO_763 (O_763,N_4796,N_4495);
nand UO_764 (O_764,N_4063,N_4927);
and UO_765 (O_765,N_4442,N_4897);
and UO_766 (O_766,N_4470,N_4538);
nor UO_767 (O_767,N_4562,N_4576);
xor UO_768 (O_768,N_4652,N_4051);
or UO_769 (O_769,N_4887,N_4551);
nor UO_770 (O_770,N_4517,N_4065);
xnor UO_771 (O_771,N_4667,N_4044);
nand UO_772 (O_772,N_4333,N_4536);
nand UO_773 (O_773,N_4427,N_4819);
or UO_774 (O_774,N_4051,N_4910);
and UO_775 (O_775,N_4527,N_4912);
and UO_776 (O_776,N_4627,N_4902);
nor UO_777 (O_777,N_4448,N_4522);
nor UO_778 (O_778,N_4026,N_4891);
nor UO_779 (O_779,N_4811,N_4127);
nor UO_780 (O_780,N_4899,N_4659);
or UO_781 (O_781,N_4205,N_4638);
and UO_782 (O_782,N_4998,N_4690);
or UO_783 (O_783,N_4266,N_4901);
nand UO_784 (O_784,N_4454,N_4541);
xnor UO_785 (O_785,N_4048,N_4723);
nand UO_786 (O_786,N_4844,N_4102);
and UO_787 (O_787,N_4169,N_4851);
and UO_788 (O_788,N_4416,N_4205);
xnor UO_789 (O_789,N_4732,N_4636);
nor UO_790 (O_790,N_4144,N_4617);
and UO_791 (O_791,N_4633,N_4217);
nand UO_792 (O_792,N_4213,N_4438);
or UO_793 (O_793,N_4022,N_4078);
nand UO_794 (O_794,N_4858,N_4074);
nor UO_795 (O_795,N_4514,N_4017);
or UO_796 (O_796,N_4351,N_4872);
nor UO_797 (O_797,N_4112,N_4870);
and UO_798 (O_798,N_4052,N_4156);
nand UO_799 (O_799,N_4124,N_4133);
or UO_800 (O_800,N_4302,N_4837);
and UO_801 (O_801,N_4050,N_4225);
nand UO_802 (O_802,N_4679,N_4065);
or UO_803 (O_803,N_4571,N_4850);
nand UO_804 (O_804,N_4620,N_4244);
or UO_805 (O_805,N_4874,N_4927);
nand UO_806 (O_806,N_4746,N_4972);
or UO_807 (O_807,N_4168,N_4611);
xor UO_808 (O_808,N_4674,N_4980);
and UO_809 (O_809,N_4098,N_4035);
and UO_810 (O_810,N_4665,N_4454);
or UO_811 (O_811,N_4207,N_4373);
and UO_812 (O_812,N_4173,N_4649);
or UO_813 (O_813,N_4494,N_4557);
and UO_814 (O_814,N_4148,N_4327);
or UO_815 (O_815,N_4251,N_4151);
or UO_816 (O_816,N_4010,N_4966);
nand UO_817 (O_817,N_4097,N_4810);
xnor UO_818 (O_818,N_4730,N_4746);
and UO_819 (O_819,N_4175,N_4837);
nor UO_820 (O_820,N_4590,N_4113);
and UO_821 (O_821,N_4351,N_4366);
nand UO_822 (O_822,N_4945,N_4939);
or UO_823 (O_823,N_4629,N_4796);
nand UO_824 (O_824,N_4642,N_4921);
nand UO_825 (O_825,N_4559,N_4359);
nor UO_826 (O_826,N_4648,N_4757);
or UO_827 (O_827,N_4669,N_4439);
and UO_828 (O_828,N_4384,N_4901);
and UO_829 (O_829,N_4219,N_4813);
nand UO_830 (O_830,N_4781,N_4082);
and UO_831 (O_831,N_4287,N_4899);
or UO_832 (O_832,N_4096,N_4495);
or UO_833 (O_833,N_4938,N_4731);
and UO_834 (O_834,N_4950,N_4879);
or UO_835 (O_835,N_4484,N_4078);
nor UO_836 (O_836,N_4298,N_4198);
nor UO_837 (O_837,N_4366,N_4864);
nor UO_838 (O_838,N_4561,N_4071);
nor UO_839 (O_839,N_4415,N_4769);
xnor UO_840 (O_840,N_4229,N_4822);
nand UO_841 (O_841,N_4466,N_4429);
xnor UO_842 (O_842,N_4444,N_4279);
nand UO_843 (O_843,N_4922,N_4168);
or UO_844 (O_844,N_4883,N_4210);
nand UO_845 (O_845,N_4932,N_4857);
nand UO_846 (O_846,N_4363,N_4440);
nor UO_847 (O_847,N_4493,N_4436);
xor UO_848 (O_848,N_4255,N_4151);
nor UO_849 (O_849,N_4249,N_4152);
and UO_850 (O_850,N_4321,N_4273);
nor UO_851 (O_851,N_4168,N_4169);
xnor UO_852 (O_852,N_4057,N_4490);
or UO_853 (O_853,N_4557,N_4465);
nand UO_854 (O_854,N_4228,N_4817);
nand UO_855 (O_855,N_4891,N_4857);
and UO_856 (O_856,N_4343,N_4568);
or UO_857 (O_857,N_4650,N_4859);
and UO_858 (O_858,N_4247,N_4005);
nor UO_859 (O_859,N_4283,N_4668);
xnor UO_860 (O_860,N_4482,N_4794);
nor UO_861 (O_861,N_4630,N_4135);
nor UO_862 (O_862,N_4172,N_4499);
or UO_863 (O_863,N_4147,N_4104);
and UO_864 (O_864,N_4459,N_4458);
and UO_865 (O_865,N_4791,N_4158);
and UO_866 (O_866,N_4341,N_4196);
or UO_867 (O_867,N_4926,N_4367);
and UO_868 (O_868,N_4540,N_4864);
and UO_869 (O_869,N_4509,N_4054);
or UO_870 (O_870,N_4318,N_4593);
nand UO_871 (O_871,N_4704,N_4609);
and UO_872 (O_872,N_4598,N_4864);
or UO_873 (O_873,N_4377,N_4366);
nand UO_874 (O_874,N_4725,N_4753);
nand UO_875 (O_875,N_4858,N_4946);
or UO_876 (O_876,N_4796,N_4175);
xnor UO_877 (O_877,N_4572,N_4107);
or UO_878 (O_878,N_4585,N_4741);
nor UO_879 (O_879,N_4071,N_4797);
or UO_880 (O_880,N_4204,N_4668);
and UO_881 (O_881,N_4211,N_4163);
and UO_882 (O_882,N_4596,N_4803);
or UO_883 (O_883,N_4927,N_4586);
nand UO_884 (O_884,N_4231,N_4394);
nand UO_885 (O_885,N_4626,N_4845);
nor UO_886 (O_886,N_4286,N_4539);
xor UO_887 (O_887,N_4493,N_4698);
and UO_888 (O_888,N_4572,N_4515);
nor UO_889 (O_889,N_4672,N_4590);
nand UO_890 (O_890,N_4219,N_4136);
and UO_891 (O_891,N_4564,N_4023);
nor UO_892 (O_892,N_4297,N_4471);
and UO_893 (O_893,N_4030,N_4779);
nand UO_894 (O_894,N_4764,N_4424);
or UO_895 (O_895,N_4329,N_4743);
xor UO_896 (O_896,N_4408,N_4430);
nand UO_897 (O_897,N_4048,N_4706);
and UO_898 (O_898,N_4652,N_4555);
or UO_899 (O_899,N_4081,N_4599);
xor UO_900 (O_900,N_4067,N_4292);
nor UO_901 (O_901,N_4582,N_4658);
nor UO_902 (O_902,N_4141,N_4538);
nor UO_903 (O_903,N_4968,N_4240);
nor UO_904 (O_904,N_4159,N_4843);
xor UO_905 (O_905,N_4801,N_4134);
nand UO_906 (O_906,N_4160,N_4395);
nor UO_907 (O_907,N_4117,N_4660);
xor UO_908 (O_908,N_4609,N_4702);
and UO_909 (O_909,N_4383,N_4818);
nand UO_910 (O_910,N_4057,N_4075);
nor UO_911 (O_911,N_4832,N_4287);
nor UO_912 (O_912,N_4473,N_4914);
nor UO_913 (O_913,N_4424,N_4647);
or UO_914 (O_914,N_4413,N_4368);
nand UO_915 (O_915,N_4450,N_4901);
nor UO_916 (O_916,N_4690,N_4467);
and UO_917 (O_917,N_4455,N_4704);
nor UO_918 (O_918,N_4062,N_4198);
and UO_919 (O_919,N_4567,N_4539);
nand UO_920 (O_920,N_4980,N_4380);
and UO_921 (O_921,N_4534,N_4206);
xor UO_922 (O_922,N_4465,N_4482);
nor UO_923 (O_923,N_4150,N_4797);
or UO_924 (O_924,N_4390,N_4057);
or UO_925 (O_925,N_4259,N_4094);
and UO_926 (O_926,N_4970,N_4758);
and UO_927 (O_927,N_4230,N_4202);
and UO_928 (O_928,N_4265,N_4357);
nand UO_929 (O_929,N_4659,N_4200);
nand UO_930 (O_930,N_4924,N_4150);
or UO_931 (O_931,N_4535,N_4888);
nor UO_932 (O_932,N_4788,N_4074);
and UO_933 (O_933,N_4803,N_4006);
nor UO_934 (O_934,N_4826,N_4614);
xor UO_935 (O_935,N_4802,N_4722);
and UO_936 (O_936,N_4596,N_4185);
or UO_937 (O_937,N_4711,N_4687);
xor UO_938 (O_938,N_4069,N_4544);
and UO_939 (O_939,N_4128,N_4190);
nor UO_940 (O_940,N_4756,N_4945);
xor UO_941 (O_941,N_4145,N_4661);
nand UO_942 (O_942,N_4915,N_4559);
nand UO_943 (O_943,N_4273,N_4906);
or UO_944 (O_944,N_4305,N_4996);
nand UO_945 (O_945,N_4013,N_4864);
nor UO_946 (O_946,N_4505,N_4304);
nand UO_947 (O_947,N_4179,N_4957);
nand UO_948 (O_948,N_4038,N_4186);
nor UO_949 (O_949,N_4132,N_4577);
xor UO_950 (O_950,N_4961,N_4983);
and UO_951 (O_951,N_4634,N_4436);
and UO_952 (O_952,N_4466,N_4183);
xor UO_953 (O_953,N_4323,N_4919);
or UO_954 (O_954,N_4370,N_4908);
nor UO_955 (O_955,N_4244,N_4555);
nand UO_956 (O_956,N_4572,N_4693);
or UO_957 (O_957,N_4032,N_4890);
nor UO_958 (O_958,N_4150,N_4554);
or UO_959 (O_959,N_4034,N_4370);
nor UO_960 (O_960,N_4594,N_4624);
nor UO_961 (O_961,N_4231,N_4828);
nor UO_962 (O_962,N_4133,N_4244);
and UO_963 (O_963,N_4929,N_4632);
nor UO_964 (O_964,N_4687,N_4677);
nand UO_965 (O_965,N_4661,N_4573);
nor UO_966 (O_966,N_4000,N_4585);
and UO_967 (O_967,N_4637,N_4382);
nand UO_968 (O_968,N_4620,N_4702);
or UO_969 (O_969,N_4103,N_4819);
xnor UO_970 (O_970,N_4386,N_4215);
nand UO_971 (O_971,N_4166,N_4818);
and UO_972 (O_972,N_4230,N_4510);
and UO_973 (O_973,N_4549,N_4598);
nor UO_974 (O_974,N_4014,N_4263);
nand UO_975 (O_975,N_4689,N_4344);
nand UO_976 (O_976,N_4806,N_4613);
nand UO_977 (O_977,N_4246,N_4593);
or UO_978 (O_978,N_4367,N_4442);
and UO_979 (O_979,N_4427,N_4615);
or UO_980 (O_980,N_4856,N_4169);
and UO_981 (O_981,N_4975,N_4805);
nand UO_982 (O_982,N_4667,N_4259);
nand UO_983 (O_983,N_4061,N_4599);
nor UO_984 (O_984,N_4257,N_4577);
and UO_985 (O_985,N_4921,N_4603);
or UO_986 (O_986,N_4133,N_4192);
or UO_987 (O_987,N_4310,N_4273);
xnor UO_988 (O_988,N_4517,N_4113);
or UO_989 (O_989,N_4279,N_4725);
and UO_990 (O_990,N_4791,N_4235);
nor UO_991 (O_991,N_4855,N_4220);
and UO_992 (O_992,N_4548,N_4850);
nor UO_993 (O_993,N_4515,N_4357);
and UO_994 (O_994,N_4645,N_4792);
xor UO_995 (O_995,N_4906,N_4581);
nor UO_996 (O_996,N_4103,N_4140);
and UO_997 (O_997,N_4102,N_4924);
or UO_998 (O_998,N_4905,N_4808);
nand UO_999 (O_999,N_4881,N_4758);
endmodule