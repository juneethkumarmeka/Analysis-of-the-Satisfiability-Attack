module basic_500_3000_500_15_levels_1xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_300,In_380);
nand U1 (N_1,In_112,In_189);
nand U2 (N_2,In_401,In_377);
or U3 (N_3,In_379,In_140);
nor U4 (N_4,In_206,In_292);
nor U5 (N_5,In_194,In_187);
nand U6 (N_6,In_450,In_183);
nor U7 (N_7,In_98,In_313);
and U8 (N_8,In_15,In_352);
nand U9 (N_9,In_257,In_225);
nor U10 (N_10,In_268,In_477);
or U11 (N_11,In_488,In_64);
and U12 (N_12,In_70,In_97);
nand U13 (N_13,In_82,In_472);
and U14 (N_14,In_199,In_163);
nand U15 (N_15,In_246,In_339);
and U16 (N_16,In_141,In_28);
nor U17 (N_17,In_185,In_224);
nor U18 (N_18,In_165,In_443);
and U19 (N_19,In_402,In_137);
or U20 (N_20,In_11,In_394);
and U21 (N_21,In_243,In_494);
and U22 (N_22,In_66,In_440);
and U23 (N_23,In_407,In_170);
and U24 (N_24,In_456,In_188);
and U25 (N_25,In_328,In_279);
and U26 (N_26,In_31,In_209);
nand U27 (N_27,In_434,In_338);
nor U28 (N_28,In_422,In_260);
and U29 (N_29,In_304,In_419);
or U30 (N_30,In_441,In_14);
nand U31 (N_31,In_195,In_463);
nand U32 (N_32,In_453,In_364);
nand U33 (N_33,In_439,In_404);
or U34 (N_34,In_399,In_301);
or U35 (N_35,In_400,In_147);
xnor U36 (N_36,In_219,In_158);
nand U37 (N_37,In_231,In_267);
nand U38 (N_38,In_196,In_480);
nand U39 (N_39,In_376,In_295);
or U40 (N_40,In_266,In_322);
and U41 (N_41,In_424,In_174);
and U42 (N_42,In_86,In_235);
or U43 (N_43,In_412,In_151);
nor U44 (N_44,In_464,In_389);
nand U45 (N_45,In_336,In_121);
or U46 (N_46,In_375,In_294);
or U47 (N_47,In_331,In_208);
or U48 (N_48,In_242,In_438);
nor U49 (N_49,In_349,In_396);
nor U50 (N_50,In_489,In_492);
or U51 (N_51,In_362,In_384);
and U52 (N_52,In_299,In_272);
nand U53 (N_53,In_385,In_34);
nand U54 (N_54,In_214,In_129);
or U55 (N_55,In_393,In_454);
and U56 (N_56,In_499,In_491);
nand U57 (N_57,In_133,In_6);
xor U58 (N_58,In_172,In_43);
and U59 (N_59,In_91,In_126);
nand U60 (N_60,In_146,In_479);
nand U61 (N_61,In_123,In_104);
nand U62 (N_62,In_226,In_35);
nor U63 (N_63,In_96,In_85);
nand U64 (N_64,In_285,In_53);
nand U65 (N_65,In_343,In_127);
nor U66 (N_66,In_405,In_284);
and U67 (N_67,In_144,In_200);
nand U68 (N_68,In_81,In_452);
or U69 (N_69,In_378,In_9);
and U70 (N_70,In_65,In_447);
or U71 (N_71,In_215,In_261);
nand U72 (N_72,In_236,In_397);
nand U73 (N_73,In_40,In_22);
and U74 (N_74,In_56,In_333);
nor U75 (N_75,In_168,In_132);
nand U76 (N_76,In_136,In_288);
nand U77 (N_77,In_18,In_61);
or U78 (N_78,In_448,In_486);
nor U79 (N_79,In_363,In_204);
nand U80 (N_80,In_13,In_446);
or U81 (N_81,In_153,In_345);
nor U82 (N_82,In_36,In_227);
and U83 (N_83,In_234,In_88);
and U84 (N_84,In_125,In_370);
nand U85 (N_85,In_5,In_167);
and U86 (N_86,In_42,In_326);
nor U87 (N_87,In_415,In_83);
or U88 (N_88,In_365,In_203);
and U89 (N_89,In_94,In_179);
or U90 (N_90,In_164,In_390);
or U91 (N_91,In_425,In_131);
or U92 (N_92,In_367,In_223);
nor U93 (N_93,In_344,In_57);
nor U94 (N_94,In_148,In_386);
or U95 (N_95,In_368,In_113);
nand U96 (N_96,In_445,In_449);
or U97 (N_97,In_392,In_0);
and U98 (N_98,In_108,In_103);
and U99 (N_99,In_38,In_232);
nand U100 (N_100,In_319,In_178);
or U101 (N_101,In_433,In_324);
nand U102 (N_102,In_241,In_497);
nor U103 (N_103,In_309,In_411);
and U104 (N_104,In_247,In_150);
nand U105 (N_105,In_408,In_17);
nand U106 (N_106,In_220,In_473);
nor U107 (N_107,In_171,In_250);
nor U108 (N_108,In_459,In_106);
and U109 (N_109,In_277,In_26);
nor U110 (N_110,In_8,In_275);
or U111 (N_111,In_193,In_481);
and U112 (N_112,In_259,In_293);
nor U113 (N_113,In_467,In_84);
nor U114 (N_114,In_240,In_186);
and U115 (N_115,In_342,In_382);
nand U116 (N_116,In_311,In_444);
and U117 (N_117,In_366,In_76);
or U118 (N_118,In_149,In_239);
or U119 (N_119,In_74,In_25);
and U120 (N_120,In_340,In_278);
or U121 (N_121,In_37,In_303);
nand U122 (N_122,In_59,In_471);
nor U123 (N_123,In_205,In_12);
or U124 (N_124,In_460,In_197);
nand U125 (N_125,In_317,In_431);
and U126 (N_126,In_381,In_77);
nand U127 (N_127,In_207,In_255);
and U128 (N_128,In_273,In_281);
and U129 (N_129,In_20,In_361);
and U130 (N_130,In_469,In_3);
nor U131 (N_131,In_184,In_298);
and U132 (N_132,In_156,In_413);
nor U133 (N_133,In_175,In_134);
nor U134 (N_134,In_249,In_201);
nor U135 (N_135,In_45,In_212);
nor U136 (N_136,In_332,In_107);
nor U137 (N_137,In_327,In_198);
or U138 (N_138,In_290,In_258);
and U139 (N_139,In_470,In_166);
nor U140 (N_140,In_182,In_287);
nand U141 (N_141,In_120,In_245);
and U142 (N_142,In_202,In_323);
nor U143 (N_143,In_466,In_16);
nor U144 (N_144,In_346,In_73);
nand U145 (N_145,In_369,In_263);
nand U146 (N_146,In_110,In_359);
nor U147 (N_147,In_173,In_128);
nor U148 (N_148,In_429,In_63);
or U149 (N_149,In_30,In_102);
and U150 (N_150,In_347,In_169);
nand U151 (N_151,In_302,In_253);
and U152 (N_152,In_355,In_305);
and U153 (N_153,In_32,In_130);
nand U154 (N_154,In_181,In_10);
nor U155 (N_155,In_124,In_387);
or U156 (N_156,In_335,In_282);
and U157 (N_157,In_493,In_180);
nor U158 (N_158,In_496,In_348);
nor U159 (N_159,In_67,In_315);
or U160 (N_160,In_62,In_437);
or U161 (N_161,In_116,In_44);
or U162 (N_162,In_270,In_468);
nor U163 (N_163,In_310,In_498);
nor U164 (N_164,In_432,In_2);
or U165 (N_165,In_19,In_230);
and U166 (N_166,In_55,In_353);
and U167 (N_167,In_29,In_90);
nor U168 (N_168,In_118,In_406);
nor U169 (N_169,In_428,In_283);
nor U170 (N_170,In_251,In_47);
xnor U171 (N_171,In_115,In_291);
nor U172 (N_172,In_482,In_92);
nor U173 (N_173,In_487,In_33);
and U174 (N_174,In_75,In_69);
and U175 (N_175,In_418,In_354);
or U176 (N_176,In_229,In_135);
and U177 (N_177,In_60,In_383);
nand U178 (N_178,In_391,In_7);
or U179 (N_179,In_119,In_1);
or U180 (N_180,In_289,In_143);
nand U181 (N_181,In_160,In_161);
or U182 (N_182,In_274,In_142);
nand U183 (N_183,In_276,In_403);
nand U184 (N_184,In_318,In_254);
or U185 (N_185,In_122,In_307);
nor U186 (N_186,In_216,In_49);
or U187 (N_187,In_72,In_217);
nand U188 (N_188,In_192,In_478);
nor U189 (N_189,In_58,In_373);
or U190 (N_190,In_233,In_374);
nor U191 (N_191,In_145,In_21);
nand U192 (N_192,In_337,In_495);
or U193 (N_193,In_341,In_414);
nand U194 (N_194,In_458,In_237);
or U195 (N_195,In_280,In_360);
and U196 (N_196,In_435,In_89);
nand U197 (N_197,In_426,In_117);
nor U198 (N_198,In_330,In_442);
nor U199 (N_199,In_256,In_474);
or U200 (N_200,N_117,In_351);
nand U201 (N_201,N_68,N_28);
nand U202 (N_202,N_153,In_177);
and U203 (N_203,N_190,N_95);
and U204 (N_204,In_211,N_100);
nand U205 (N_205,In_420,In_430);
and U206 (N_206,N_105,N_189);
nand U207 (N_207,N_71,N_111);
and U208 (N_208,N_55,In_334);
and U209 (N_209,N_39,N_193);
nand U210 (N_210,N_154,N_57);
or U211 (N_211,In_176,N_72);
nand U212 (N_212,In_371,In_190);
or U213 (N_213,N_87,N_130);
and U214 (N_214,N_138,N_104);
nor U215 (N_215,N_51,N_126);
nor U216 (N_216,In_485,In_461);
and U217 (N_217,N_41,N_74);
or U218 (N_218,N_120,N_127);
and U219 (N_219,N_1,N_194);
nand U220 (N_220,N_150,In_321);
and U221 (N_221,N_7,In_455);
nand U222 (N_222,N_131,N_93);
nand U223 (N_223,N_158,N_69);
nor U224 (N_224,In_325,In_476);
and U225 (N_225,N_84,N_24);
nand U226 (N_226,N_144,In_286);
or U227 (N_227,N_91,N_73);
nor U228 (N_228,N_60,N_43);
nor U229 (N_229,In_271,N_83);
or U230 (N_230,N_70,In_316);
nor U231 (N_231,In_248,N_192);
or U232 (N_232,N_186,In_423);
nand U233 (N_233,N_159,In_306);
nor U234 (N_234,N_64,N_79);
nor U235 (N_235,N_33,N_183);
nor U236 (N_236,N_181,In_350);
xor U237 (N_237,N_2,N_119);
and U238 (N_238,N_171,N_179);
and U239 (N_239,N_114,N_14);
and U240 (N_240,In_162,N_106);
and U241 (N_241,N_92,N_38);
or U242 (N_242,N_121,In_297);
nor U243 (N_243,N_163,N_12);
nand U244 (N_244,N_11,N_156);
and U245 (N_245,N_56,In_314);
and U246 (N_246,N_97,In_264);
nor U247 (N_247,In_155,In_54);
nand U248 (N_248,N_169,N_35);
nand U249 (N_249,N_184,N_182);
nor U250 (N_250,N_109,In_356);
nand U251 (N_251,N_62,In_262);
or U252 (N_252,In_410,N_99);
nor U253 (N_253,N_174,N_67);
and U254 (N_254,N_40,N_176);
nand U255 (N_255,In_465,N_107);
nor U256 (N_256,N_132,N_167);
and U257 (N_257,N_133,N_52);
nor U258 (N_258,N_145,In_114);
nor U259 (N_259,N_139,N_29);
or U260 (N_260,In_152,In_312);
or U261 (N_261,N_47,N_75);
xor U262 (N_262,N_178,N_78);
and U263 (N_263,In_421,N_198);
and U264 (N_264,In_50,In_238);
xnor U265 (N_265,In_475,N_122);
and U266 (N_266,N_37,N_31);
or U267 (N_267,N_147,N_32);
nor U268 (N_268,In_222,N_23);
nor U269 (N_269,In_388,N_16);
nand U270 (N_270,N_140,N_157);
nand U271 (N_271,In_213,N_103);
nor U272 (N_272,In_157,N_141);
and U273 (N_273,N_30,In_79);
nor U274 (N_274,In_4,In_78);
nand U275 (N_275,In_417,N_102);
nor U276 (N_276,In_296,N_173);
or U277 (N_277,N_108,In_320);
nand U278 (N_278,In_159,N_172);
and U279 (N_279,N_4,In_218);
nor U280 (N_280,In_462,N_5);
nand U281 (N_281,N_170,In_80);
nor U282 (N_282,N_36,In_221);
nand U283 (N_283,N_187,N_129);
or U284 (N_284,N_17,In_27);
and U285 (N_285,In_358,In_451);
nor U286 (N_286,In_416,N_180);
or U287 (N_287,N_3,In_46);
and U288 (N_288,N_96,N_42);
and U289 (N_289,In_51,N_101);
or U290 (N_290,N_177,In_329);
nor U291 (N_291,In_252,In_95);
and U292 (N_292,N_152,In_101);
nor U293 (N_293,In_372,In_138);
nor U294 (N_294,N_63,In_457);
nor U295 (N_295,N_142,N_18);
or U296 (N_296,N_66,N_161);
nor U297 (N_297,N_19,N_50);
or U298 (N_298,N_49,N_6);
or U299 (N_299,N_88,N_149);
and U300 (N_300,In_191,In_357);
nand U301 (N_301,N_48,N_175);
or U302 (N_302,In_395,N_20);
nand U303 (N_303,N_81,In_111);
nand U304 (N_304,In_484,In_100);
nor U305 (N_305,N_197,N_137);
or U306 (N_306,N_80,N_89);
and U307 (N_307,In_244,N_77);
and U308 (N_308,In_483,In_210);
xor U309 (N_309,In_154,In_228);
nand U310 (N_310,In_308,N_45);
nor U311 (N_311,N_98,N_113);
and U312 (N_312,In_269,N_168);
or U313 (N_313,N_135,N_85);
nand U314 (N_314,In_105,N_155);
and U315 (N_315,In_48,N_8);
nand U316 (N_316,In_68,N_166);
or U317 (N_317,N_22,N_116);
nand U318 (N_318,N_10,N_128);
nor U319 (N_319,N_94,N_191);
nand U320 (N_320,N_151,In_139);
and U321 (N_321,In_265,In_490);
nand U322 (N_322,N_134,N_54);
or U323 (N_323,N_196,N_13);
or U324 (N_324,N_125,In_71);
or U325 (N_325,N_26,In_41);
and U326 (N_326,N_0,N_34);
nand U327 (N_327,In_409,In_39);
nand U328 (N_328,N_59,N_27);
nand U329 (N_329,In_52,In_436);
or U330 (N_330,N_148,N_15);
and U331 (N_331,N_195,N_112);
and U332 (N_332,In_93,In_427);
nor U333 (N_333,N_143,N_162);
nand U334 (N_334,N_115,N_110);
nand U335 (N_335,N_165,N_53);
nor U336 (N_336,N_136,N_25);
and U337 (N_337,N_58,N_44);
and U338 (N_338,N_118,N_124);
or U339 (N_339,N_164,N_185);
and U340 (N_340,In_109,N_21);
nor U341 (N_341,N_123,N_46);
nand U342 (N_342,In_24,N_61);
or U343 (N_343,N_146,N_65);
nor U344 (N_344,N_188,In_99);
nor U345 (N_345,N_82,In_398);
nor U346 (N_346,N_76,N_160);
or U347 (N_347,N_9,N_199);
nand U348 (N_348,In_23,In_87);
nor U349 (N_349,N_86,N_90);
and U350 (N_350,N_142,N_58);
nand U351 (N_351,N_95,N_19);
and U352 (N_352,N_56,In_306);
and U353 (N_353,In_296,N_43);
and U354 (N_354,N_161,N_192);
nand U355 (N_355,N_70,N_197);
and U356 (N_356,N_30,N_122);
nor U357 (N_357,In_420,N_98);
and U358 (N_358,N_163,N_192);
nor U359 (N_359,N_6,N_60);
and U360 (N_360,In_139,N_163);
and U361 (N_361,In_436,N_11);
and U362 (N_362,In_244,In_334);
nand U363 (N_363,In_350,N_78);
and U364 (N_364,In_358,N_18);
nand U365 (N_365,N_96,N_36);
nor U366 (N_366,In_308,In_269);
and U367 (N_367,N_23,N_58);
nand U368 (N_368,N_100,N_14);
and U369 (N_369,N_52,In_286);
nor U370 (N_370,In_320,N_92);
nand U371 (N_371,N_73,N_90);
and U372 (N_372,N_2,N_193);
nor U373 (N_373,In_159,N_75);
nor U374 (N_374,In_398,In_485);
or U375 (N_375,In_114,In_111);
and U376 (N_376,N_130,N_173);
and U377 (N_377,In_111,N_160);
or U378 (N_378,N_157,N_195);
nand U379 (N_379,In_78,In_176);
or U380 (N_380,N_192,N_91);
nand U381 (N_381,In_271,N_1);
nand U382 (N_382,N_3,N_0);
and U383 (N_383,N_74,N_34);
nand U384 (N_384,In_114,In_100);
or U385 (N_385,In_222,In_475);
nor U386 (N_386,In_177,N_47);
nand U387 (N_387,N_144,N_136);
nand U388 (N_388,N_111,In_213);
nor U389 (N_389,N_167,N_176);
or U390 (N_390,N_26,N_79);
nand U391 (N_391,N_116,In_114);
or U392 (N_392,In_296,N_45);
nor U393 (N_393,N_109,N_112);
nand U394 (N_394,N_99,In_190);
and U395 (N_395,N_132,N_157);
and U396 (N_396,In_297,N_197);
and U397 (N_397,In_213,In_52);
and U398 (N_398,In_50,N_69);
or U399 (N_399,N_181,N_20);
nand U400 (N_400,N_356,N_387);
or U401 (N_401,N_318,N_280);
nor U402 (N_402,N_323,N_274);
nor U403 (N_403,N_298,N_276);
nor U404 (N_404,N_257,N_374);
nor U405 (N_405,N_287,N_333);
or U406 (N_406,N_368,N_295);
and U407 (N_407,N_212,N_348);
or U408 (N_408,N_320,N_313);
or U409 (N_409,N_273,N_342);
and U410 (N_410,N_345,N_380);
or U411 (N_411,N_346,N_221);
or U412 (N_412,N_247,N_343);
or U413 (N_413,N_326,N_224);
xnor U414 (N_414,N_241,N_250);
and U415 (N_415,N_246,N_354);
nor U416 (N_416,N_294,N_204);
or U417 (N_417,N_265,N_379);
and U418 (N_418,N_338,N_261);
and U419 (N_419,N_200,N_311);
and U420 (N_420,N_330,N_254);
nand U421 (N_421,N_357,N_235);
or U422 (N_422,N_361,N_314);
and U423 (N_423,N_209,N_205);
nand U424 (N_424,N_244,N_266);
nor U425 (N_425,N_281,N_225);
and U426 (N_426,N_251,N_258);
and U427 (N_427,N_301,N_369);
nor U428 (N_428,N_389,N_341);
nand U429 (N_429,N_296,N_291);
or U430 (N_430,N_353,N_384);
and U431 (N_431,N_340,N_292);
or U432 (N_432,N_252,N_390);
nand U433 (N_433,N_271,N_332);
nor U434 (N_434,N_238,N_308);
or U435 (N_435,N_325,N_347);
nand U436 (N_436,N_297,N_371);
or U437 (N_437,N_321,N_370);
or U438 (N_438,N_366,N_226);
nor U439 (N_439,N_222,N_207);
nor U440 (N_440,N_299,N_272);
and U441 (N_441,N_236,N_249);
and U442 (N_442,N_277,N_324);
and U443 (N_443,N_396,N_334);
or U444 (N_444,N_386,N_201);
or U445 (N_445,N_358,N_208);
or U446 (N_446,N_335,N_256);
nor U447 (N_447,N_391,N_383);
or U448 (N_448,N_215,N_203);
or U449 (N_449,N_315,N_220);
and U450 (N_450,N_240,N_372);
or U451 (N_451,N_398,N_286);
and U452 (N_452,N_397,N_278);
and U453 (N_453,N_377,N_259);
and U454 (N_454,N_223,N_243);
or U455 (N_455,N_234,N_337);
and U456 (N_456,N_382,N_309);
nor U457 (N_457,N_206,N_290);
or U458 (N_458,N_305,N_317);
nor U459 (N_459,N_385,N_217);
and U460 (N_460,N_331,N_388);
nor U461 (N_461,N_375,N_216);
or U462 (N_462,N_306,N_351);
nor U463 (N_463,N_365,N_229);
nand U464 (N_464,N_312,N_242);
or U465 (N_465,N_322,N_355);
or U466 (N_466,N_362,N_211);
nor U467 (N_467,N_237,N_394);
nand U468 (N_468,N_231,N_339);
and U469 (N_469,N_393,N_359);
or U470 (N_470,N_336,N_304);
nor U471 (N_471,N_275,N_253);
or U472 (N_472,N_310,N_248);
and U473 (N_473,N_260,N_255);
and U474 (N_474,N_367,N_303);
and U475 (N_475,N_329,N_352);
or U476 (N_476,N_307,N_270);
nand U477 (N_477,N_302,N_213);
nand U478 (N_478,N_344,N_327);
nor U479 (N_479,N_230,N_283);
nor U480 (N_480,N_264,N_328);
nand U481 (N_481,N_267,N_219);
or U482 (N_482,N_279,N_316);
and U483 (N_483,N_289,N_288);
or U484 (N_484,N_285,N_245);
and U485 (N_485,N_350,N_395);
or U486 (N_486,N_218,N_360);
and U487 (N_487,N_363,N_399);
nor U488 (N_488,N_269,N_376);
nand U489 (N_489,N_239,N_300);
or U490 (N_490,N_232,N_319);
and U491 (N_491,N_378,N_227);
nor U492 (N_492,N_282,N_381);
and U493 (N_493,N_214,N_233);
and U494 (N_494,N_228,N_262);
nand U495 (N_495,N_392,N_202);
nor U496 (N_496,N_349,N_293);
nand U497 (N_497,N_210,N_263);
or U498 (N_498,N_373,N_284);
and U499 (N_499,N_268,N_364);
nand U500 (N_500,N_201,N_348);
or U501 (N_501,N_223,N_342);
nor U502 (N_502,N_259,N_238);
nor U503 (N_503,N_346,N_249);
or U504 (N_504,N_258,N_225);
or U505 (N_505,N_305,N_306);
and U506 (N_506,N_242,N_295);
nand U507 (N_507,N_201,N_319);
or U508 (N_508,N_347,N_328);
or U509 (N_509,N_396,N_223);
nand U510 (N_510,N_340,N_217);
nand U511 (N_511,N_306,N_238);
nor U512 (N_512,N_271,N_378);
and U513 (N_513,N_315,N_359);
and U514 (N_514,N_232,N_383);
nor U515 (N_515,N_220,N_229);
nor U516 (N_516,N_223,N_216);
nor U517 (N_517,N_295,N_342);
or U518 (N_518,N_210,N_328);
nand U519 (N_519,N_379,N_328);
nor U520 (N_520,N_273,N_320);
nor U521 (N_521,N_279,N_201);
nor U522 (N_522,N_314,N_225);
nand U523 (N_523,N_268,N_369);
and U524 (N_524,N_320,N_389);
or U525 (N_525,N_205,N_318);
nand U526 (N_526,N_255,N_288);
or U527 (N_527,N_246,N_240);
nor U528 (N_528,N_353,N_203);
and U529 (N_529,N_229,N_246);
and U530 (N_530,N_282,N_386);
nand U531 (N_531,N_312,N_232);
or U532 (N_532,N_257,N_396);
or U533 (N_533,N_327,N_339);
or U534 (N_534,N_385,N_361);
or U535 (N_535,N_232,N_310);
or U536 (N_536,N_346,N_348);
nand U537 (N_537,N_287,N_224);
and U538 (N_538,N_255,N_354);
nand U539 (N_539,N_232,N_362);
and U540 (N_540,N_346,N_223);
or U541 (N_541,N_278,N_232);
or U542 (N_542,N_206,N_251);
nor U543 (N_543,N_200,N_212);
or U544 (N_544,N_353,N_251);
or U545 (N_545,N_287,N_340);
and U546 (N_546,N_308,N_351);
or U547 (N_547,N_351,N_296);
and U548 (N_548,N_245,N_377);
nand U549 (N_549,N_228,N_273);
nand U550 (N_550,N_373,N_357);
or U551 (N_551,N_214,N_326);
nand U552 (N_552,N_294,N_270);
and U553 (N_553,N_310,N_228);
nor U554 (N_554,N_374,N_336);
nand U555 (N_555,N_329,N_376);
and U556 (N_556,N_394,N_232);
nand U557 (N_557,N_397,N_362);
nand U558 (N_558,N_205,N_330);
and U559 (N_559,N_382,N_266);
and U560 (N_560,N_213,N_286);
nand U561 (N_561,N_317,N_384);
and U562 (N_562,N_330,N_317);
nor U563 (N_563,N_306,N_236);
and U564 (N_564,N_318,N_367);
and U565 (N_565,N_370,N_363);
nand U566 (N_566,N_246,N_326);
and U567 (N_567,N_281,N_230);
or U568 (N_568,N_250,N_345);
nor U569 (N_569,N_348,N_388);
nand U570 (N_570,N_231,N_277);
nor U571 (N_571,N_235,N_366);
and U572 (N_572,N_290,N_326);
nand U573 (N_573,N_373,N_312);
and U574 (N_574,N_301,N_226);
nor U575 (N_575,N_262,N_276);
nor U576 (N_576,N_202,N_387);
nand U577 (N_577,N_308,N_243);
nand U578 (N_578,N_334,N_310);
or U579 (N_579,N_247,N_392);
nor U580 (N_580,N_357,N_366);
nor U581 (N_581,N_357,N_244);
nand U582 (N_582,N_369,N_244);
or U583 (N_583,N_328,N_256);
nand U584 (N_584,N_341,N_348);
nand U585 (N_585,N_355,N_228);
or U586 (N_586,N_371,N_212);
and U587 (N_587,N_288,N_349);
and U588 (N_588,N_263,N_368);
and U589 (N_589,N_363,N_233);
nor U590 (N_590,N_352,N_378);
or U591 (N_591,N_265,N_234);
and U592 (N_592,N_209,N_273);
or U593 (N_593,N_301,N_381);
or U594 (N_594,N_369,N_353);
nand U595 (N_595,N_274,N_287);
or U596 (N_596,N_244,N_398);
nand U597 (N_597,N_342,N_222);
nor U598 (N_598,N_244,N_275);
and U599 (N_599,N_315,N_258);
or U600 (N_600,N_531,N_533);
and U601 (N_601,N_445,N_451);
and U602 (N_602,N_447,N_410);
nand U603 (N_603,N_590,N_420);
nand U604 (N_604,N_502,N_488);
or U605 (N_605,N_416,N_406);
or U606 (N_606,N_535,N_570);
or U607 (N_607,N_518,N_465);
nor U608 (N_608,N_558,N_541);
nor U609 (N_609,N_430,N_520);
nand U610 (N_610,N_546,N_461);
or U611 (N_611,N_459,N_584);
and U612 (N_612,N_519,N_515);
nand U613 (N_613,N_555,N_435);
or U614 (N_614,N_462,N_452);
nor U615 (N_615,N_424,N_534);
nand U616 (N_616,N_597,N_592);
nand U617 (N_617,N_510,N_573);
xor U618 (N_618,N_583,N_512);
and U619 (N_619,N_409,N_492);
nor U620 (N_620,N_401,N_526);
nor U621 (N_621,N_438,N_582);
or U622 (N_622,N_446,N_575);
nand U623 (N_623,N_460,N_464);
or U624 (N_624,N_439,N_544);
nor U625 (N_625,N_494,N_405);
nor U626 (N_626,N_580,N_429);
or U627 (N_627,N_469,N_470);
nand U628 (N_628,N_495,N_589);
nand U629 (N_629,N_411,N_566);
or U630 (N_630,N_527,N_486);
nor U631 (N_631,N_467,N_413);
or U632 (N_632,N_521,N_567);
nand U633 (N_633,N_530,N_440);
nand U634 (N_634,N_588,N_581);
nor U635 (N_635,N_565,N_574);
nand U636 (N_636,N_455,N_454);
nand U637 (N_637,N_428,N_499);
and U638 (N_638,N_506,N_417);
or U639 (N_639,N_412,N_436);
nor U640 (N_640,N_538,N_550);
nand U641 (N_641,N_414,N_537);
and U642 (N_642,N_457,N_491);
or U643 (N_643,N_479,N_487);
nand U644 (N_644,N_431,N_579);
nand U645 (N_645,N_482,N_442);
nor U646 (N_646,N_596,N_478);
and U647 (N_647,N_493,N_542);
nand U648 (N_648,N_498,N_554);
and U649 (N_649,N_419,N_556);
and U650 (N_650,N_539,N_423);
and U651 (N_651,N_441,N_514);
or U652 (N_652,N_595,N_594);
nor U653 (N_653,N_540,N_418);
and U654 (N_654,N_528,N_598);
or U655 (N_655,N_517,N_426);
nor U656 (N_656,N_571,N_475);
nor U657 (N_657,N_472,N_415);
nor U658 (N_658,N_402,N_543);
nand U659 (N_659,N_501,N_549);
nand U660 (N_660,N_507,N_545);
nor U661 (N_661,N_557,N_505);
nand U662 (N_662,N_548,N_471);
or U663 (N_663,N_508,N_561);
nor U664 (N_664,N_577,N_504);
nor U665 (N_665,N_587,N_569);
or U666 (N_666,N_425,N_552);
and U667 (N_667,N_568,N_585);
nor U668 (N_668,N_407,N_536);
nor U669 (N_669,N_443,N_403);
nand U670 (N_670,N_497,N_477);
nor U671 (N_671,N_466,N_562);
or U672 (N_672,N_578,N_563);
nor U673 (N_673,N_553,N_532);
nor U674 (N_674,N_458,N_473);
or U675 (N_675,N_513,N_444);
nor U676 (N_676,N_516,N_522);
nand U677 (N_677,N_468,N_422);
nand U678 (N_678,N_551,N_485);
nand U679 (N_679,N_450,N_500);
nor U680 (N_680,N_448,N_576);
and U681 (N_681,N_433,N_404);
nand U682 (N_682,N_564,N_523);
nor U683 (N_683,N_484,N_480);
and U684 (N_684,N_463,N_408);
or U685 (N_685,N_449,N_400);
nor U686 (N_686,N_483,N_591);
xor U687 (N_687,N_453,N_434);
and U688 (N_688,N_560,N_437);
and U689 (N_689,N_456,N_481);
or U690 (N_690,N_427,N_503);
or U691 (N_691,N_547,N_586);
nand U692 (N_692,N_529,N_572);
nor U693 (N_693,N_559,N_525);
nor U694 (N_694,N_511,N_490);
or U695 (N_695,N_524,N_489);
and U696 (N_696,N_593,N_476);
xor U697 (N_697,N_421,N_474);
nand U698 (N_698,N_496,N_432);
and U699 (N_699,N_509,N_599);
nand U700 (N_700,N_484,N_591);
nand U701 (N_701,N_428,N_412);
or U702 (N_702,N_412,N_420);
nor U703 (N_703,N_517,N_537);
nand U704 (N_704,N_485,N_435);
and U705 (N_705,N_564,N_568);
nand U706 (N_706,N_438,N_505);
and U707 (N_707,N_401,N_563);
nor U708 (N_708,N_482,N_473);
and U709 (N_709,N_410,N_409);
and U710 (N_710,N_426,N_503);
nor U711 (N_711,N_470,N_486);
and U712 (N_712,N_596,N_528);
and U713 (N_713,N_404,N_593);
and U714 (N_714,N_537,N_557);
or U715 (N_715,N_597,N_447);
nor U716 (N_716,N_405,N_465);
nor U717 (N_717,N_547,N_474);
nor U718 (N_718,N_579,N_427);
nor U719 (N_719,N_576,N_463);
nor U720 (N_720,N_573,N_413);
or U721 (N_721,N_545,N_490);
nor U722 (N_722,N_558,N_472);
nand U723 (N_723,N_457,N_455);
or U724 (N_724,N_442,N_577);
and U725 (N_725,N_408,N_406);
or U726 (N_726,N_473,N_553);
and U727 (N_727,N_528,N_415);
nand U728 (N_728,N_532,N_442);
nor U729 (N_729,N_429,N_413);
nand U730 (N_730,N_577,N_423);
nor U731 (N_731,N_525,N_560);
nand U732 (N_732,N_499,N_432);
or U733 (N_733,N_513,N_560);
or U734 (N_734,N_559,N_513);
and U735 (N_735,N_400,N_481);
xnor U736 (N_736,N_486,N_450);
and U737 (N_737,N_559,N_515);
or U738 (N_738,N_597,N_540);
nor U739 (N_739,N_553,N_481);
nand U740 (N_740,N_419,N_516);
nor U741 (N_741,N_473,N_582);
nor U742 (N_742,N_540,N_511);
nor U743 (N_743,N_516,N_523);
or U744 (N_744,N_586,N_497);
nand U745 (N_745,N_414,N_545);
nand U746 (N_746,N_434,N_564);
nor U747 (N_747,N_444,N_508);
nor U748 (N_748,N_545,N_589);
or U749 (N_749,N_458,N_403);
nand U750 (N_750,N_533,N_478);
nor U751 (N_751,N_474,N_466);
and U752 (N_752,N_429,N_488);
nand U753 (N_753,N_406,N_510);
nand U754 (N_754,N_565,N_546);
and U755 (N_755,N_542,N_571);
nor U756 (N_756,N_508,N_446);
or U757 (N_757,N_493,N_507);
and U758 (N_758,N_549,N_447);
nor U759 (N_759,N_472,N_407);
nand U760 (N_760,N_521,N_477);
nand U761 (N_761,N_553,N_407);
nand U762 (N_762,N_458,N_420);
nor U763 (N_763,N_414,N_501);
nand U764 (N_764,N_593,N_553);
or U765 (N_765,N_534,N_432);
nor U766 (N_766,N_427,N_483);
nor U767 (N_767,N_525,N_501);
nand U768 (N_768,N_598,N_532);
nand U769 (N_769,N_585,N_499);
and U770 (N_770,N_507,N_523);
and U771 (N_771,N_491,N_515);
and U772 (N_772,N_572,N_521);
and U773 (N_773,N_591,N_513);
nand U774 (N_774,N_540,N_578);
nand U775 (N_775,N_583,N_412);
nand U776 (N_776,N_502,N_478);
or U777 (N_777,N_573,N_462);
nand U778 (N_778,N_497,N_558);
and U779 (N_779,N_504,N_520);
and U780 (N_780,N_550,N_494);
and U781 (N_781,N_461,N_406);
nor U782 (N_782,N_467,N_465);
and U783 (N_783,N_450,N_421);
nand U784 (N_784,N_519,N_575);
or U785 (N_785,N_420,N_476);
or U786 (N_786,N_557,N_599);
or U787 (N_787,N_577,N_461);
or U788 (N_788,N_443,N_502);
nand U789 (N_789,N_590,N_559);
nand U790 (N_790,N_485,N_583);
or U791 (N_791,N_589,N_476);
nor U792 (N_792,N_594,N_562);
and U793 (N_793,N_405,N_541);
or U794 (N_794,N_571,N_478);
nor U795 (N_795,N_510,N_525);
or U796 (N_796,N_540,N_489);
or U797 (N_797,N_451,N_454);
or U798 (N_798,N_516,N_474);
nor U799 (N_799,N_523,N_558);
nor U800 (N_800,N_736,N_770);
or U801 (N_801,N_642,N_685);
nor U802 (N_802,N_647,N_707);
nand U803 (N_803,N_619,N_765);
nand U804 (N_804,N_716,N_625);
nand U805 (N_805,N_792,N_651);
nand U806 (N_806,N_708,N_670);
nor U807 (N_807,N_639,N_652);
nor U808 (N_808,N_641,N_693);
nand U809 (N_809,N_633,N_780);
nand U810 (N_810,N_632,N_630);
nand U811 (N_811,N_705,N_700);
nor U812 (N_812,N_669,N_774);
nand U813 (N_813,N_755,N_745);
nor U814 (N_814,N_614,N_742);
nor U815 (N_815,N_674,N_704);
nor U816 (N_816,N_711,N_724);
and U817 (N_817,N_684,N_794);
and U818 (N_818,N_661,N_601);
nor U819 (N_819,N_662,N_748);
or U820 (N_820,N_753,N_752);
nor U821 (N_821,N_744,N_603);
nor U822 (N_822,N_616,N_648);
nor U823 (N_823,N_714,N_681);
nor U824 (N_824,N_672,N_675);
nand U825 (N_825,N_608,N_760);
nor U826 (N_826,N_718,N_689);
and U827 (N_827,N_605,N_719);
nand U828 (N_828,N_717,N_725);
and U829 (N_829,N_721,N_747);
and U830 (N_830,N_620,N_624);
nand U831 (N_831,N_613,N_627);
and U832 (N_832,N_712,N_754);
or U833 (N_833,N_791,N_631);
nand U834 (N_834,N_715,N_628);
nand U835 (N_835,N_730,N_697);
and U836 (N_836,N_673,N_653);
and U837 (N_837,N_758,N_686);
and U838 (N_838,N_749,N_667);
or U839 (N_839,N_799,N_687);
or U840 (N_840,N_698,N_658);
and U841 (N_841,N_638,N_703);
nand U842 (N_842,N_602,N_699);
or U843 (N_843,N_690,N_635);
or U844 (N_844,N_757,N_696);
nor U845 (N_845,N_727,N_722);
nand U846 (N_846,N_762,N_739);
and U847 (N_847,N_640,N_680);
nand U848 (N_848,N_701,N_751);
nor U849 (N_849,N_789,N_629);
or U850 (N_850,N_797,N_644);
and U851 (N_851,N_604,N_737);
or U852 (N_852,N_679,N_793);
nand U853 (N_853,N_618,N_682);
or U854 (N_854,N_798,N_709);
or U855 (N_855,N_785,N_782);
nor U856 (N_856,N_775,N_694);
nand U857 (N_857,N_645,N_740);
or U858 (N_858,N_607,N_600);
and U859 (N_859,N_676,N_772);
nor U860 (N_860,N_666,N_763);
and U861 (N_861,N_795,N_768);
nor U862 (N_862,N_728,N_710);
nand U863 (N_863,N_621,N_750);
or U864 (N_864,N_706,N_761);
nand U865 (N_865,N_778,N_657);
or U866 (N_866,N_659,N_726);
or U867 (N_867,N_688,N_663);
and U868 (N_868,N_695,N_729);
nor U869 (N_869,N_660,N_769);
and U870 (N_870,N_788,N_790);
and U871 (N_871,N_637,N_720);
or U872 (N_872,N_786,N_735);
nor U873 (N_873,N_610,N_664);
nand U874 (N_874,N_668,N_764);
nand U875 (N_875,N_731,N_756);
and U876 (N_876,N_634,N_615);
nand U877 (N_877,N_617,N_650);
nand U878 (N_878,N_781,N_741);
nand U879 (N_879,N_665,N_783);
or U880 (N_880,N_779,N_609);
or U881 (N_881,N_623,N_636);
nor U882 (N_882,N_759,N_784);
or U883 (N_883,N_646,N_677);
nor U884 (N_884,N_777,N_732);
and U885 (N_885,N_733,N_671);
nand U886 (N_886,N_612,N_766);
nand U887 (N_887,N_771,N_655);
or U888 (N_888,N_692,N_702);
or U889 (N_889,N_787,N_611);
and U890 (N_890,N_767,N_776);
or U891 (N_891,N_626,N_656);
and U892 (N_892,N_678,N_743);
nand U893 (N_893,N_649,N_606);
nand U894 (N_894,N_683,N_738);
and U895 (N_895,N_622,N_723);
nor U896 (N_896,N_746,N_796);
and U897 (N_897,N_713,N_654);
nor U898 (N_898,N_734,N_773);
nor U899 (N_899,N_691,N_643);
or U900 (N_900,N_743,N_770);
nor U901 (N_901,N_788,N_677);
nand U902 (N_902,N_617,N_646);
nor U903 (N_903,N_713,N_689);
nand U904 (N_904,N_607,N_616);
and U905 (N_905,N_641,N_773);
nor U906 (N_906,N_750,N_651);
or U907 (N_907,N_698,N_799);
and U908 (N_908,N_706,N_617);
or U909 (N_909,N_734,N_793);
nor U910 (N_910,N_629,N_632);
nor U911 (N_911,N_606,N_736);
nor U912 (N_912,N_700,N_630);
and U913 (N_913,N_741,N_663);
and U914 (N_914,N_670,N_768);
nand U915 (N_915,N_746,N_648);
or U916 (N_916,N_704,N_752);
or U917 (N_917,N_775,N_753);
nor U918 (N_918,N_797,N_633);
and U919 (N_919,N_685,N_625);
or U920 (N_920,N_642,N_653);
nor U921 (N_921,N_737,N_671);
and U922 (N_922,N_689,N_617);
nor U923 (N_923,N_613,N_744);
and U924 (N_924,N_615,N_606);
nor U925 (N_925,N_758,N_687);
and U926 (N_926,N_688,N_658);
and U927 (N_927,N_601,N_657);
nor U928 (N_928,N_698,N_773);
nand U929 (N_929,N_788,N_697);
or U930 (N_930,N_782,N_628);
and U931 (N_931,N_631,N_711);
nor U932 (N_932,N_668,N_724);
and U933 (N_933,N_665,N_740);
or U934 (N_934,N_654,N_604);
nand U935 (N_935,N_784,N_715);
nor U936 (N_936,N_626,N_687);
nor U937 (N_937,N_619,N_660);
or U938 (N_938,N_765,N_696);
nor U939 (N_939,N_660,N_727);
and U940 (N_940,N_663,N_713);
and U941 (N_941,N_615,N_792);
nand U942 (N_942,N_665,N_690);
and U943 (N_943,N_725,N_756);
nand U944 (N_944,N_645,N_771);
nor U945 (N_945,N_715,N_771);
nand U946 (N_946,N_773,N_786);
nand U947 (N_947,N_608,N_646);
nor U948 (N_948,N_600,N_695);
xor U949 (N_949,N_681,N_751);
or U950 (N_950,N_628,N_681);
xnor U951 (N_951,N_748,N_765);
nor U952 (N_952,N_740,N_622);
or U953 (N_953,N_710,N_789);
or U954 (N_954,N_631,N_648);
and U955 (N_955,N_657,N_753);
nor U956 (N_956,N_740,N_628);
nor U957 (N_957,N_648,N_779);
and U958 (N_958,N_729,N_775);
or U959 (N_959,N_733,N_785);
or U960 (N_960,N_660,N_699);
and U961 (N_961,N_740,N_617);
nor U962 (N_962,N_752,N_692);
and U963 (N_963,N_723,N_625);
and U964 (N_964,N_635,N_617);
or U965 (N_965,N_614,N_621);
xnor U966 (N_966,N_695,N_705);
nand U967 (N_967,N_606,N_739);
nand U968 (N_968,N_667,N_698);
nand U969 (N_969,N_644,N_659);
and U970 (N_970,N_771,N_640);
and U971 (N_971,N_798,N_783);
nand U972 (N_972,N_643,N_635);
or U973 (N_973,N_777,N_776);
nor U974 (N_974,N_746,N_715);
nor U975 (N_975,N_712,N_775);
nor U976 (N_976,N_656,N_645);
and U977 (N_977,N_752,N_712);
nand U978 (N_978,N_729,N_667);
or U979 (N_979,N_664,N_736);
or U980 (N_980,N_664,N_729);
nor U981 (N_981,N_779,N_668);
nor U982 (N_982,N_752,N_624);
or U983 (N_983,N_625,N_759);
and U984 (N_984,N_631,N_709);
and U985 (N_985,N_764,N_727);
or U986 (N_986,N_705,N_613);
nand U987 (N_987,N_781,N_675);
and U988 (N_988,N_790,N_753);
nand U989 (N_989,N_683,N_777);
nor U990 (N_990,N_687,N_746);
nand U991 (N_991,N_763,N_662);
and U992 (N_992,N_721,N_661);
and U993 (N_993,N_706,N_746);
or U994 (N_994,N_681,N_668);
or U995 (N_995,N_748,N_617);
nor U996 (N_996,N_706,N_630);
and U997 (N_997,N_760,N_736);
and U998 (N_998,N_603,N_695);
or U999 (N_999,N_771,N_734);
and U1000 (N_1000,N_959,N_879);
or U1001 (N_1001,N_892,N_838);
nor U1002 (N_1002,N_990,N_968);
or U1003 (N_1003,N_870,N_963);
and U1004 (N_1004,N_818,N_996);
nor U1005 (N_1005,N_806,N_907);
nand U1006 (N_1006,N_826,N_914);
or U1007 (N_1007,N_971,N_932);
or U1008 (N_1008,N_869,N_831);
or U1009 (N_1009,N_832,N_920);
and U1010 (N_1010,N_926,N_897);
and U1011 (N_1011,N_814,N_810);
or U1012 (N_1012,N_816,N_946);
nor U1013 (N_1013,N_976,N_909);
and U1014 (N_1014,N_876,N_967);
nor U1015 (N_1015,N_928,N_827);
and U1016 (N_1016,N_868,N_958);
nand U1017 (N_1017,N_969,N_921);
or U1018 (N_1018,N_995,N_992);
nand U1019 (N_1019,N_880,N_973);
and U1020 (N_1020,N_982,N_993);
and U1021 (N_1021,N_863,N_858);
or U1022 (N_1022,N_917,N_828);
and U1023 (N_1023,N_900,N_804);
nand U1024 (N_1024,N_855,N_867);
nand U1025 (N_1025,N_978,N_985);
nand U1026 (N_1026,N_965,N_801);
nor U1027 (N_1027,N_989,N_925);
nor U1028 (N_1028,N_935,N_964);
and U1029 (N_1029,N_911,N_834);
and U1030 (N_1030,N_934,N_800);
nor U1031 (N_1031,N_918,N_941);
or U1032 (N_1032,N_848,N_987);
nand U1033 (N_1033,N_972,N_830);
and U1034 (N_1034,N_805,N_950);
and U1035 (N_1035,N_860,N_844);
xor U1036 (N_1036,N_984,N_986);
nor U1037 (N_1037,N_952,N_829);
and U1038 (N_1038,N_898,N_874);
nor U1039 (N_1039,N_839,N_991);
nand U1040 (N_1040,N_910,N_877);
nor U1041 (N_1041,N_916,N_923);
or U1042 (N_1042,N_807,N_866);
and U1043 (N_1043,N_882,N_851);
and U1044 (N_1044,N_853,N_891);
or U1045 (N_1045,N_889,N_822);
and U1046 (N_1046,N_942,N_802);
or U1047 (N_1047,N_825,N_861);
nand U1048 (N_1048,N_820,N_803);
and U1049 (N_1049,N_949,N_808);
nor U1050 (N_1050,N_983,N_840);
or U1051 (N_1051,N_864,N_998);
and U1052 (N_1052,N_884,N_981);
nor U1053 (N_1053,N_927,N_899);
and U1054 (N_1054,N_956,N_904);
nand U1055 (N_1055,N_930,N_997);
or U1056 (N_1056,N_811,N_924);
xnor U1057 (N_1057,N_852,N_922);
and U1058 (N_1058,N_948,N_939);
nand U1059 (N_1059,N_843,N_857);
nand U1060 (N_1060,N_962,N_841);
nand U1061 (N_1061,N_951,N_847);
and U1062 (N_1062,N_945,N_999);
nand U1063 (N_1063,N_936,N_929);
and U1064 (N_1064,N_856,N_885);
and U1065 (N_1065,N_966,N_980);
and U1066 (N_1066,N_931,N_994);
xnor U1067 (N_1067,N_835,N_815);
or U1068 (N_1068,N_943,N_854);
or U1069 (N_1069,N_850,N_961);
and U1070 (N_1070,N_893,N_819);
and U1071 (N_1071,N_902,N_817);
or U1072 (N_1072,N_890,N_979);
or U1073 (N_1073,N_974,N_913);
nand U1074 (N_1074,N_912,N_837);
and U1075 (N_1075,N_944,N_905);
nor U1076 (N_1076,N_836,N_938);
and U1077 (N_1077,N_845,N_906);
nand U1078 (N_1078,N_975,N_824);
and U1079 (N_1079,N_812,N_887);
nand U1080 (N_1080,N_937,N_878);
nor U1081 (N_1081,N_903,N_940);
or U1082 (N_1082,N_970,N_859);
nor U1083 (N_1083,N_957,N_875);
nand U1084 (N_1084,N_872,N_919);
nand U1085 (N_1085,N_886,N_895);
nor U1086 (N_1086,N_833,N_908);
and U1087 (N_1087,N_823,N_846);
or U1088 (N_1088,N_873,N_883);
and U1089 (N_1089,N_813,N_849);
and U1090 (N_1090,N_862,N_821);
xor U1091 (N_1091,N_988,N_809);
or U1092 (N_1092,N_888,N_842);
and U1093 (N_1093,N_901,N_977);
nand U1094 (N_1094,N_954,N_871);
or U1095 (N_1095,N_953,N_896);
or U1096 (N_1096,N_881,N_915);
nand U1097 (N_1097,N_955,N_933);
or U1098 (N_1098,N_947,N_960);
nor U1099 (N_1099,N_894,N_865);
or U1100 (N_1100,N_819,N_845);
nor U1101 (N_1101,N_876,N_977);
nor U1102 (N_1102,N_913,N_818);
and U1103 (N_1103,N_928,N_960);
nand U1104 (N_1104,N_911,N_914);
nor U1105 (N_1105,N_857,N_991);
nor U1106 (N_1106,N_871,N_963);
nor U1107 (N_1107,N_952,N_980);
nand U1108 (N_1108,N_987,N_807);
nor U1109 (N_1109,N_930,N_858);
or U1110 (N_1110,N_818,N_900);
and U1111 (N_1111,N_918,N_904);
xor U1112 (N_1112,N_983,N_999);
nor U1113 (N_1113,N_984,N_869);
nor U1114 (N_1114,N_901,N_994);
or U1115 (N_1115,N_902,N_803);
and U1116 (N_1116,N_878,N_974);
nand U1117 (N_1117,N_880,N_840);
nand U1118 (N_1118,N_837,N_875);
or U1119 (N_1119,N_835,N_922);
and U1120 (N_1120,N_843,N_988);
nor U1121 (N_1121,N_994,N_873);
or U1122 (N_1122,N_964,N_869);
or U1123 (N_1123,N_936,N_881);
and U1124 (N_1124,N_981,N_959);
and U1125 (N_1125,N_907,N_883);
nor U1126 (N_1126,N_929,N_914);
nor U1127 (N_1127,N_849,N_888);
and U1128 (N_1128,N_986,N_900);
nor U1129 (N_1129,N_984,N_977);
nor U1130 (N_1130,N_965,N_981);
nor U1131 (N_1131,N_826,N_847);
nor U1132 (N_1132,N_904,N_804);
and U1133 (N_1133,N_966,N_863);
nor U1134 (N_1134,N_908,N_849);
nor U1135 (N_1135,N_996,N_841);
nor U1136 (N_1136,N_835,N_826);
or U1137 (N_1137,N_886,N_814);
or U1138 (N_1138,N_954,N_869);
nand U1139 (N_1139,N_818,N_997);
nor U1140 (N_1140,N_932,N_923);
nor U1141 (N_1141,N_966,N_850);
nand U1142 (N_1142,N_824,N_870);
or U1143 (N_1143,N_891,N_918);
or U1144 (N_1144,N_893,N_838);
and U1145 (N_1145,N_910,N_831);
nor U1146 (N_1146,N_871,N_808);
or U1147 (N_1147,N_818,N_802);
nor U1148 (N_1148,N_802,N_945);
or U1149 (N_1149,N_972,N_898);
nand U1150 (N_1150,N_965,N_929);
or U1151 (N_1151,N_982,N_961);
nor U1152 (N_1152,N_999,N_930);
and U1153 (N_1153,N_885,N_934);
and U1154 (N_1154,N_918,N_920);
and U1155 (N_1155,N_928,N_909);
and U1156 (N_1156,N_822,N_971);
or U1157 (N_1157,N_821,N_988);
or U1158 (N_1158,N_914,N_824);
or U1159 (N_1159,N_924,N_848);
or U1160 (N_1160,N_968,N_995);
and U1161 (N_1161,N_811,N_964);
nand U1162 (N_1162,N_804,N_946);
nor U1163 (N_1163,N_866,N_871);
nor U1164 (N_1164,N_935,N_911);
and U1165 (N_1165,N_976,N_982);
nor U1166 (N_1166,N_967,N_991);
nand U1167 (N_1167,N_851,N_942);
nor U1168 (N_1168,N_969,N_856);
nor U1169 (N_1169,N_849,N_910);
nand U1170 (N_1170,N_935,N_891);
nor U1171 (N_1171,N_997,N_848);
and U1172 (N_1172,N_963,N_874);
and U1173 (N_1173,N_945,N_877);
or U1174 (N_1174,N_940,N_961);
nor U1175 (N_1175,N_850,N_864);
nand U1176 (N_1176,N_917,N_871);
nor U1177 (N_1177,N_812,N_866);
nor U1178 (N_1178,N_835,N_908);
or U1179 (N_1179,N_926,N_892);
nand U1180 (N_1180,N_848,N_862);
nor U1181 (N_1181,N_825,N_857);
and U1182 (N_1182,N_821,N_943);
nand U1183 (N_1183,N_912,N_831);
or U1184 (N_1184,N_875,N_938);
nand U1185 (N_1185,N_891,N_937);
or U1186 (N_1186,N_804,N_923);
nor U1187 (N_1187,N_897,N_855);
or U1188 (N_1188,N_853,N_999);
or U1189 (N_1189,N_961,N_916);
nand U1190 (N_1190,N_954,N_947);
nor U1191 (N_1191,N_969,N_886);
and U1192 (N_1192,N_910,N_816);
or U1193 (N_1193,N_873,N_973);
or U1194 (N_1194,N_900,N_847);
nand U1195 (N_1195,N_927,N_879);
or U1196 (N_1196,N_924,N_982);
nand U1197 (N_1197,N_918,N_987);
and U1198 (N_1198,N_922,N_940);
nor U1199 (N_1199,N_960,N_932);
or U1200 (N_1200,N_1137,N_1111);
nand U1201 (N_1201,N_1021,N_1195);
nand U1202 (N_1202,N_1110,N_1059);
and U1203 (N_1203,N_1047,N_1089);
and U1204 (N_1204,N_1177,N_1186);
or U1205 (N_1205,N_1055,N_1199);
nor U1206 (N_1206,N_1057,N_1116);
and U1207 (N_1207,N_1117,N_1081);
nor U1208 (N_1208,N_1112,N_1158);
or U1209 (N_1209,N_1139,N_1032);
and U1210 (N_1210,N_1051,N_1194);
or U1211 (N_1211,N_1025,N_1093);
and U1212 (N_1212,N_1009,N_1075);
or U1213 (N_1213,N_1187,N_1138);
nand U1214 (N_1214,N_1131,N_1080);
nand U1215 (N_1215,N_1049,N_1133);
nor U1216 (N_1216,N_1058,N_1044);
nand U1217 (N_1217,N_1165,N_1178);
and U1218 (N_1218,N_1061,N_1126);
or U1219 (N_1219,N_1013,N_1119);
nand U1220 (N_1220,N_1070,N_1048);
nor U1221 (N_1221,N_1184,N_1168);
or U1222 (N_1222,N_1114,N_1006);
nand U1223 (N_1223,N_1104,N_1147);
or U1224 (N_1224,N_1105,N_1183);
or U1225 (N_1225,N_1151,N_1094);
nand U1226 (N_1226,N_1159,N_1087);
or U1227 (N_1227,N_1010,N_1102);
nor U1228 (N_1228,N_1078,N_1054);
and U1229 (N_1229,N_1014,N_1115);
and U1230 (N_1230,N_1036,N_1176);
nand U1231 (N_1231,N_1141,N_1196);
nand U1232 (N_1232,N_1103,N_1097);
nand U1233 (N_1233,N_1169,N_1076);
or U1234 (N_1234,N_1012,N_1068);
and U1235 (N_1235,N_1084,N_1164);
nor U1236 (N_1236,N_1192,N_1179);
or U1237 (N_1237,N_1045,N_1030);
or U1238 (N_1238,N_1053,N_1015);
nand U1239 (N_1239,N_1038,N_1002);
or U1240 (N_1240,N_1185,N_1106);
nor U1241 (N_1241,N_1181,N_1129);
and U1242 (N_1242,N_1004,N_1118);
and U1243 (N_1243,N_1092,N_1034);
and U1244 (N_1244,N_1121,N_1050);
or U1245 (N_1245,N_1113,N_1132);
nor U1246 (N_1246,N_1163,N_1144);
nand U1247 (N_1247,N_1069,N_1149);
or U1248 (N_1248,N_1101,N_1017);
nor U1249 (N_1249,N_1091,N_1031);
nand U1250 (N_1250,N_1123,N_1090);
nand U1251 (N_1251,N_1074,N_1088);
and U1252 (N_1252,N_1062,N_1180);
nor U1253 (N_1253,N_1019,N_1124);
nand U1254 (N_1254,N_1077,N_1160);
and U1255 (N_1255,N_1098,N_1046);
nor U1256 (N_1256,N_1100,N_1039);
or U1257 (N_1257,N_1166,N_1150);
or U1258 (N_1258,N_1108,N_1016);
nand U1259 (N_1259,N_1130,N_1174);
nor U1260 (N_1260,N_1198,N_1072);
nand U1261 (N_1261,N_1154,N_1171);
or U1262 (N_1262,N_1056,N_1188);
nand U1263 (N_1263,N_1063,N_1043);
nand U1264 (N_1264,N_1120,N_1155);
and U1265 (N_1265,N_1065,N_1189);
nand U1266 (N_1266,N_1127,N_1005);
nand U1267 (N_1267,N_1128,N_1095);
and U1268 (N_1268,N_1052,N_1041);
or U1269 (N_1269,N_1083,N_1040);
or U1270 (N_1270,N_1190,N_1182);
nand U1271 (N_1271,N_1071,N_1022);
or U1272 (N_1272,N_1007,N_1146);
and U1273 (N_1273,N_1193,N_1122);
nand U1274 (N_1274,N_1008,N_1029);
nand U1275 (N_1275,N_1042,N_1135);
and U1276 (N_1276,N_1136,N_1173);
nand U1277 (N_1277,N_1082,N_1020);
or U1278 (N_1278,N_1197,N_1085);
or U1279 (N_1279,N_1035,N_1099);
nor U1280 (N_1280,N_1191,N_1018);
or U1281 (N_1281,N_1067,N_1011);
and U1282 (N_1282,N_1175,N_1064);
nor U1283 (N_1283,N_1148,N_1153);
nand U1284 (N_1284,N_1170,N_1167);
or U1285 (N_1285,N_1156,N_1073);
nand U1286 (N_1286,N_1066,N_1026);
nor U1287 (N_1287,N_1033,N_1028);
nor U1288 (N_1288,N_1037,N_1086);
nand U1289 (N_1289,N_1060,N_1027);
nand U1290 (N_1290,N_1079,N_1024);
nand U1291 (N_1291,N_1143,N_1107);
or U1292 (N_1292,N_1134,N_1096);
or U1293 (N_1293,N_1023,N_1157);
and U1294 (N_1294,N_1161,N_1172);
and U1295 (N_1295,N_1125,N_1109);
nor U1296 (N_1296,N_1140,N_1152);
nand U1297 (N_1297,N_1145,N_1003);
nand U1298 (N_1298,N_1142,N_1162);
nand U1299 (N_1299,N_1000,N_1001);
and U1300 (N_1300,N_1064,N_1194);
nand U1301 (N_1301,N_1045,N_1124);
nor U1302 (N_1302,N_1190,N_1024);
or U1303 (N_1303,N_1119,N_1197);
and U1304 (N_1304,N_1103,N_1015);
nor U1305 (N_1305,N_1155,N_1034);
and U1306 (N_1306,N_1191,N_1154);
and U1307 (N_1307,N_1083,N_1025);
nand U1308 (N_1308,N_1055,N_1165);
nand U1309 (N_1309,N_1007,N_1101);
nor U1310 (N_1310,N_1189,N_1036);
or U1311 (N_1311,N_1145,N_1159);
nand U1312 (N_1312,N_1195,N_1087);
or U1313 (N_1313,N_1006,N_1074);
or U1314 (N_1314,N_1144,N_1100);
or U1315 (N_1315,N_1072,N_1000);
and U1316 (N_1316,N_1185,N_1144);
or U1317 (N_1317,N_1089,N_1149);
nand U1318 (N_1318,N_1074,N_1011);
or U1319 (N_1319,N_1171,N_1025);
or U1320 (N_1320,N_1179,N_1139);
or U1321 (N_1321,N_1048,N_1196);
nand U1322 (N_1322,N_1150,N_1042);
and U1323 (N_1323,N_1039,N_1161);
nor U1324 (N_1324,N_1015,N_1164);
or U1325 (N_1325,N_1124,N_1179);
and U1326 (N_1326,N_1149,N_1029);
and U1327 (N_1327,N_1089,N_1025);
nand U1328 (N_1328,N_1135,N_1126);
or U1329 (N_1329,N_1134,N_1113);
nor U1330 (N_1330,N_1185,N_1001);
or U1331 (N_1331,N_1076,N_1125);
nor U1332 (N_1332,N_1004,N_1194);
and U1333 (N_1333,N_1078,N_1097);
nand U1334 (N_1334,N_1112,N_1138);
or U1335 (N_1335,N_1050,N_1136);
or U1336 (N_1336,N_1122,N_1158);
or U1337 (N_1337,N_1051,N_1161);
nor U1338 (N_1338,N_1020,N_1037);
nor U1339 (N_1339,N_1135,N_1022);
xor U1340 (N_1340,N_1010,N_1027);
and U1341 (N_1341,N_1024,N_1069);
or U1342 (N_1342,N_1013,N_1126);
or U1343 (N_1343,N_1043,N_1083);
nor U1344 (N_1344,N_1071,N_1117);
nand U1345 (N_1345,N_1118,N_1049);
nand U1346 (N_1346,N_1036,N_1100);
or U1347 (N_1347,N_1007,N_1172);
and U1348 (N_1348,N_1058,N_1131);
or U1349 (N_1349,N_1026,N_1131);
or U1350 (N_1350,N_1135,N_1007);
or U1351 (N_1351,N_1118,N_1174);
nand U1352 (N_1352,N_1194,N_1181);
nor U1353 (N_1353,N_1033,N_1195);
and U1354 (N_1354,N_1010,N_1024);
and U1355 (N_1355,N_1139,N_1153);
nor U1356 (N_1356,N_1091,N_1032);
nor U1357 (N_1357,N_1079,N_1130);
or U1358 (N_1358,N_1179,N_1151);
nand U1359 (N_1359,N_1105,N_1092);
or U1360 (N_1360,N_1025,N_1150);
nor U1361 (N_1361,N_1192,N_1090);
nor U1362 (N_1362,N_1195,N_1068);
nand U1363 (N_1363,N_1111,N_1195);
and U1364 (N_1364,N_1003,N_1038);
nand U1365 (N_1365,N_1033,N_1142);
and U1366 (N_1366,N_1092,N_1018);
nand U1367 (N_1367,N_1152,N_1175);
nor U1368 (N_1368,N_1168,N_1051);
nand U1369 (N_1369,N_1187,N_1108);
or U1370 (N_1370,N_1127,N_1125);
and U1371 (N_1371,N_1058,N_1011);
or U1372 (N_1372,N_1076,N_1135);
nor U1373 (N_1373,N_1078,N_1042);
and U1374 (N_1374,N_1128,N_1087);
nor U1375 (N_1375,N_1019,N_1150);
and U1376 (N_1376,N_1082,N_1196);
nand U1377 (N_1377,N_1132,N_1092);
or U1378 (N_1378,N_1178,N_1161);
nor U1379 (N_1379,N_1157,N_1098);
and U1380 (N_1380,N_1184,N_1076);
nor U1381 (N_1381,N_1114,N_1032);
nand U1382 (N_1382,N_1059,N_1180);
nand U1383 (N_1383,N_1063,N_1093);
xor U1384 (N_1384,N_1135,N_1140);
nand U1385 (N_1385,N_1099,N_1115);
nand U1386 (N_1386,N_1156,N_1107);
or U1387 (N_1387,N_1066,N_1143);
nand U1388 (N_1388,N_1134,N_1102);
nor U1389 (N_1389,N_1163,N_1070);
nand U1390 (N_1390,N_1153,N_1012);
nor U1391 (N_1391,N_1086,N_1144);
nor U1392 (N_1392,N_1012,N_1053);
nor U1393 (N_1393,N_1061,N_1053);
nor U1394 (N_1394,N_1082,N_1093);
nor U1395 (N_1395,N_1124,N_1051);
nand U1396 (N_1396,N_1001,N_1038);
and U1397 (N_1397,N_1146,N_1113);
nand U1398 (N_1398,N_1109,N_1104);
nand U1399 (N_1399,N_1106,N_1159);
and U1400 (N_1400,N_1228,N_1304);
or U1401 (N_1401,N_1212,N_1312);
nand U1402 (N_1402,N_1233,N_1234);
or U1403 (N_1403,N_1295,N_1319);
nor U1404 (N_1404,N_1235,N_1274);
or U1405 (N_1405,N_1358,N_1374);
nand U1406 (N_1406,N_1209,N_1398);
nand U1407 (N_1407,N_1347,N_1381);
and U1408 (N_1408,N_1222,N_1263);
or U1409 (N_1409,N_1213,N_1357);
or U1410 (N_1410,N_1223,N_1253);
and U1411 (N_1411,N_1226,N_1307);
xnor U1412 (N_1412,N_1225,N_1315);
and U1413 (N_1413,N_1217,N_1335);
and U1414 (N_1414,N_1201,N_1279);
and U1415 (N_1415,N_1282,N_1297);
nor U1416 (N_1416,N_1322,N_1311);
or U1417 (N_1417,N_1254,N_1305);
or U1418 (N_1418,N_1382,N_1386);
nor U1419 (N_1419,N_1373,N_1251);
and U1420 (N_1420,N_1390,N_1365);
or U1421 (N_1421,N_1351,N_1215);
nand U1422 (N_1422,N_1264,N_1211);
nor U1423 (N_1423,N_1363,N_1290);
nand U1424 (N_1424,N_1376,N_1393);
or U1425 (N_1425,N_1385,N_1270);
or U1426 (N_1426,N_1291,N_1368);
nor U1427 (N_1427,N_1397,N_1361);
nor U1428 (N_1428,N_1378,N_1289);
nor U1429 (N_1429,N_1370,N_1324);
and U1430 (N_1430,N_1230,N_1210);
or U1431 (N_1431,N_1343,N_1362);
and U1432 (N_1432,N_1298,N_1310);
and U1433 (N_1433,N_1241,N_1281);
nor U1434 (N_1434,N_1349,N_1229);
nand U1435 (N_1435,N_1334,N_1208);
nand U1436 (N_1436,N_1388,N_1238);
or U1437 (N_1437,N_1342,N_1389);
nand U1438 (N_1438,N_1326,N_1272);
nand U1439 (N_1439,N_1301,N_1224);
nand U1440 (N_1440,N_1392,N_1395);
nor U1441 (N_1441,N_1247,N_1308);
nor U1442 (N_1442,N_1339,N_1205);
nand U1443 (N_1443,N_1366,N_1303);
or U1444 (N_1444,N_1354,N_1258);
or U1445 (N_1445,N_1283,N_1330);
or U1446 (N_1446,N_1246,N_1353);
nor U1447 (N_1447,N_1337,N_1250);
nor U1448 (N_1448,N_1317,N_1359);
nor U1449 (N_1449,N_1300,N_1255);
nor U1450 (N_1450,N_1204,N_1329);
nor U1451 (N_1451,N_1273,N_1203);
or U1452 (N_1452,N_1240,N_1399);
nand U1453 (N_1453,N_1276,N_1265);
nor U1454 (N_1454,N_1227,N_1318);
nand U1455 (N_1455,N_1364,N_1261);
or U1456 (N_1456,N_1380,N_1313);
and U1457 (N_1457,N_1341,N_1256);
and U1458 (N_1458,N_1271,N_1360);
or U1459 (N_1459,N_1375,N_1244);
nand U1460 (N_1460,N_1325,N_1287);
and U1461 (N_1461,N_1356,N_1284);
nand U1462 (N_1462,N_1350,N_1396);
nor U1463 (N_1463,N_1232,N_1331);
and U1464 (N_1464,N_1296,N_1387);
and U1465 (N_1465,N_1377,N_1248);
nand U1466 (N_1466,N_1321,N_1278);
nor U1467 (N_1467,N_1237,N_1327);
and U1468 (N_1468,N_1216,N_1383);
and U1469 (N_1469,N_1275,N_1344);
nand U1470 (N_1470,N_1285,N_1268);
and U1471 (N_1471,N_1206,N_1259);
nor U1472 (N_1472,N_1299,N_1391);
nor U1473 (N_1473,N_1286,N_1207);
and U1474 (N_1474,N_1239,N_1336);
nand U1475 (N_1475,N_1394,N_1346);
nor U1476 (N_1476,N_1323,N_1243);
or U1477 (N_1477,N_1294,N_1277);
nand U1478 (N_1478,N_1202,N_1306);
nor U1479 (N_1479,N_1352,N_1316);
or U1480 (N_1480,N_1257,N_1340);
nor U1481 (N_1481,N_1355,N_1372);
or U1482 (N_1482,N_1236,N_1293);
or U1483 (N_1483,N_1302,N_1262);
nand U1484 (N_1484,N_1332,N_1260);
or U1485 (N_1485,N_1371,N_1328);
and U1486 (N_1486,N_1314,N_1220);
nand U1487 (N_1487,N_1221,N_1252);
and U1488 (N_1488,N_1280,N_1249);
and U1489 (N_1489,N_1369,N_1320);
and U1490 (N_1490,N_1309,N_1338);
and U1491 (N_1491,N_1345,N_1348);
or U1492 (N_1492,N_1333,N_1219);
xor U1493 (N_1493,N_1231,N_1214);
and U1494 (N_1494,N_1200,N_1267);
or U1495 (N_1495,N_1288,N_1269);
nor U1496 (N_1496,N_1379,N_1245);
or U1497 (N_1497,N_1384,N_1218);
and U1498 (N_1498,N_1242,N_1292);
or U1499 (N_1499,N_1266,N_1367);
nor U1500 (N_1500,N_1232,N_1308);
nand U1501 (N_1501,N_1353,N_1220);
or U1502 (N_1502,N_1325,N_1310);
nor U1503 (N_1503,N_1259,N_1363);
and U1504 (N_1504,N_1306,N_1305);
and U1505 (N_1505,N_1259,N_1210);
and U1506 (N_1506,N_1306,N_1263);
nor U1507 (N_1507,N_1268,N_1235);
nand U1508 (N_1508,N_1302,N_1272);
or U1509 (N_1509,N_1362,N_1391);
nor U1510 (N_1510,N_1200,N_1398);
nor U1511 (N_1511,N_1237,N_1380);
nor U1512 (N_1512,N_1271,N_1290);
or U1513 (N_1513,N_1375,N_1249);
and U1514 (N_1514,N_1351,N_1269);
nor U1515 (N_1515,N_1317,N_1201);
and U1516 (N_1516,N_1316,N_1376);
or U1517 (N_1517,N_1222,N_1292);
nand U1518 (N_1518,N_1303,N_1332);
nand U1519 (N_1519,N_1293,N_1234);
and U1520 (N_1520,N_1288,N_1254);
and U1521 (N_1521,N_1339,N_1239);
or U1522 (N_1522,N_1364,N_1202);
nand U1523 (N_1523,N_1226,N_1398);
nand U1524 (N_1524,N_1259,N_1263);
nand U1525 (N_1525,N_1226,N_1241);
nor U1526 (N_1526,N_1333,N_1340);
or U1527 (N_1527,N_1366,N_1255);
nor U1528 (N_1528,N_1390,N_1332);
and U1529 (N_1529,N_1330,N_1300);
and U1530 (N_1530,N_1248,N_1218);
and U1531 (N_1531,N_1259,N_1224);
nand U1532 (N_1532,N_1231,N_1389);
nand U1533 (N_1533,N_1253,N_1276);
nor U1534 (N_1534,N_1347,N_1387);
and U1535 (N_1535,N_1278,N_1351);
and U1536 (N_1536,N_1352,N_1290);
and U1537 (N_1537,N_1333,N_1214);
and U1538 (N_1538,N_1226,N_1271);
and U1539 (N_1539,N_1253,N_1380);
or U1540 (N_1540,N_1289,N_1233);
or U1541 (N_1541,N_1235,N_1387);
and U1542 (N_1542,N_1295,N_1308);
xor U1543 (N_1543,N_1331,N_1243);
nor U1544 (N_1544,N_1392,N_1348);
nor U1545 (N_1545,N_1346,N_1335);
and U1546 (N_1546,N_1321,N_1355);
and U1547 (N_1547,N_1214,N_1225);
nand U1548 (N_1548,N_1276,N_1302);
nor U1549 (N_1549,N_1276,N_1298);
nor U1550 (N_1550,N_1329,N_1200);
and U1551 (N_1551,N_1312,N_1220);
or U1552 (N_1552,N_1367,N_1354);
or U1553 (N_1553,N_1348,N_1349);
and U1554 (N_1554,N_1341,N_1332);
nand U1555 (N_1555,N_1259,N_1202);
nor U1556 (N_1556,N_1279,N_1228);
and U1557 (N_1557,N_1379,N_1205);
or U1558 (N_1558,N_1365,N_1347);
and U1559 (N_1559,N_1399,N_1320);
and U1560 (N_1560,N_1370,N_1219);
nand U1561 (N_1561,N_1305,N_1357);
and U1562 (N_1562,N_1344,N_1290);
nor U1563 (N_1563,N_1263,N_1311);
and U1564 (N_1564,N_1203,N_1356);
nor U1565 (N_1565,N_1207,N_1335);
nor U1566 (N_1566,N_1399,N_1247);
or U1567 (N_1567,N_1363,N_1368);
and U1568 (N_1568,N_1360,N_1249);
and U1569 (N_1569,N_1361,N_1307);
or U1570 (N_1570,N_1309,N_1332);
nor U1571 (N_1571,N_1385,N_1290);
or U1572 (N_1572,N_1380,N_1394);
or U1573 (N_1573,N_1362,N_1284);
nand U1574 (N_1574,N_1303,N_1355);
nor U1575 (N_1575,N_1217,N_1301);
nor U1576 (N_1576,N_1273,N_1319);
nor U1577 (N_1577,N_1383,N_1398);
and U1578 (N_1578,N_1373,N_1306);
nor U1579 (N_1579,N_1213,N_1234);
nor U1580 (N_1580,N_1246,N_1382);
and U1581 (N_1581,N_1383,N_1381);
nor U1582 (N_1582,N_1222,N_1392);
nor U1583 (N_1583,N_1323,N_1239);
and U1584 (N_1584,N_1238,N_1300);
nand U1585 (N_1585,N_1288,N_1354);
nand U1586 (N_1586,N_1268,N_1367);
or U1587 (N_1587,N_1268,N_1336);
and U1588 (N_1588,N_1309,N_1241);
and U1589 (N_1589,N_1255,N_1351);
or U1590 (N_1590,N_1330,N_1347);
nor U1591 (N_1591,N_1268,N_1326);
or U1592 (N_1592,N_1283,N_1351);
nand U1593 (N_1593,N_1257,N_1240);
nand U1594 (N_1594,N_1330,N_1343);
nand U1595 (N_1595,N_1304,N_1377);
or U1596 (N_1596,N_1250,N_1379);
or U1597 (N_1597,N_1340,N_1234);
nand U1598 (N_1598,N_1319,N_1244);
nor U1599 (N_1599,N_1335,N_1293);
and U1600 (N_1600,N_1556,N_1552);
nand U1601 (N_1601,N_1442,N_1526);
nor U1602 (N_1602,N_1419,N_1478);
nor U1603 (N_1603,N_1590,N_1426);
and U1604 (N_1604,N_1407,N_1599);
or U1605 (N_1605,N_1542,N_1516);
nand U1606 (N_1606,N_1579,N_1533);
or U1607 (N_1607,N_1432,N_1520);
or U1608 (N_1608,N_1561,N_1548);
and U1609 (N_1609,N_1546,N_1562);
or U1610 (N_1610,N_1462,N_1522);
and U1611 (N_1611,N_1568,N_1457);
and U1612 (N_1612,N_1497,N_1467);
or U1613 (N_1613,N_1483,N_1471);
nand U1614 (N_1614,N_1448,N_1592);
nor U1615 (N_1615,N_1447,N_1591);
or U1616 (N_1616,N_1479,N_1494);
and U1617 (N_1617,N_1539,N_1456);
or U1618 (N_1618,N_1450,N_1530);
or U1619 (N_1619,N_1524,N_1581);
nand U1620 (N_1620,N_1582,N_1434);
or U1621 (N_1621,N_1474,N_1585);
or U1622 (N_1622,N_1482,N_1451);
nor U1623 (N_1623,N_1436,N_1597);
or U1624 (N_1624,N_1584,N_1430);
or U1625 (N_1625,N_1550,N_1502);
nand U1626 (N_1626,N_1423,N_1402);
or U1627 (N_1627,N_1527,N_1574);
or U1628 (N_1628,N_1498,N_1500);
nor U1629 (N_1629,N_1566,N_1560);
nor U1630 (N_1630,N_1421,N_1531);
or U1631 (N_1631,N_1427,N_1578);
or U1632 (N_1632,N_1567,N_1463);
nand U1633 (N_1633,N_1484,N_1464);
nand U1634 (N_1634,N_1535,N_1510);
or U1635 (N_1635,N_1565,N_1557);
nand U1636 (N_1636,N_1460,N_1499);
nor U1637 (N_1637,N_1595,N_1435);
and U1638 (N_1638,N_1587,N_1558);
nand U1639 (N_1639,N_1577,N_1428);
nor U1640 (N_1640,N_1572,N_1505);
or U1641 (N_1641,N_1540,N_1443);
nand U1642 (N_1642,N_1411,N_1404);
nor U1643 (N_1643,N_1525,N_1598);
and U1644 (N_1644,N_1408,N_1521);
or U1645 (N_1645,N_1431,N_1593);
nor U1646 (N_1646,N_1509,N_1424);
or U1647 (N_1647,N_1507,N_1481);
and U1648 (N_1648,N_1555,N_1449);
and U1649 (N_1649,N_1551,N_1454);
or U1650 (N_1650,N_1405,N_1586);
nand U1651 (N_1651,N_1475,N_1594);
nor U1652 (N_1652,N_1512,N_1480);
and U1653 (N_1653,N_1458,N_1536);
nor U1654 (N_1654,N_1420,N_1563);
or U1655 (N_1655,N_1501,N_1487);
nand U1656 (N_1656,N_1476,N_1532);
and U1657 (N_1657,N_1553,N_1439);
nor U1658 (N_1658,N_1415,N_1508);
nor U1659 (N_1659,N_1575,N_1485);
or U1660 (N_1660,N_1490,N_1441);
or U1661 (N_1661,N_1477,N_1570);
or U1662 (N_1662,N_1410,N_1491);
or U1663 (N_1663,N_1406,N_1488);
and U1664 (N_1664,N_1543,N_1496);
nand U1665 (N_1665,N_1489,N_1511);
nor U1666 (N_1666,N_1412,N_1414);
and U1667 (N_1667,N_1400,N_1588);
nor U1668 (N_1668,N_1538,N_1576);
or U1669 (N_1669,N_1418,N_1545);
and U1670 (N_1670,N_1514,N_1569);
and U1671 (N_1671,N_1549,N_1466);
nor U1672 (N_1672,N_1519,N_1438);
and U1673 (N_1673,N_1437,N_1469);
or U1674 (N_1674,N_1495,N_1401);
nor U1675 (N_1675,N_1445,N_1403);
nor U1676 (N_1676,N_1537,N_1573);
and U1677 (N_1677,N_1452,N_1455);
and U1678 (N_1678,N_1515,N_1413);
and U1679 (N_1679,N_1523,N_1417);
and U1680 (N_1680,N_1506,N_1470);
nor U1681 (N_1681,N_1459,N_1583);
nor U1682 (N_1682,N_1461,N_1541);
nand U1683 (N_1683,N_1425,N_1554);
or U1684 (N_1684,N_1547,N_1503);
nor U1685 (N_1685,N_1564,N_1580);
and U1686 (N_1686,N_1409,N_1529);
nand U1687 (N_1687,N_1544,N_1472);
or U1688 (N_1688,N_1517,N_1433);
or U1689 (N_1689,N_1493,N_1473);
and U1690 (N_1690,N_1518,N_1528);
or U1691 (N_1691,N_1422,N_1440);
nand U1692 (N_1692,N_1513,N_1589);
or U1693 (N_1693,N_1596,N_1468);
nand U1694 (N_1694,N_1444,N_1504);
nand U1695 (N_1695,N_1416,N_1446);
or U1696 (N_1696,N_1571,N_1486);
nor U1697 (N_1697,N_1453,N_1534);
or U1698 (N_1698,N_1429,N_1559);
or U1699 (N_1699,N_1465,N_1492);
nor U1700 (N_1700,N_1454,N_1481);
nor U1701 (N_1701,N_1510,N_1582);
nor U1702 (N_1702,N_1573,N_1460);
nand U1703 (N_1703,N_1586,N_1530);
or U1704 (N_1704,N_1448,N_1571);
and U1705 (N_1705,N_1515,N_1566);
nand U1706 (N_1706,N_1528,N_1545);
or U1707 (N_1707,N_1446,N_1528);
nand U1708 (N_1708,N_1485,N_1594);
and U1709 (N_1709,N_1551,N_1475);
nor U1710 (N_1710,N_1415,N_1458);
nor U1711 (N_1711,N_1546,N_1599);
nor U1712 (N_1712,N_1493,N_1577);
or U1713 (N_1713,N_1456,N_1440);
or U1714 (N_1714,N_1454,N_1558);
or U1715 (N_1715,N_1455,N_1424);
or U1716 (N_1716,N_1511,N_1418);
nand U1717 (N_1717,N_1416,N_1466);
nor U1718 (N_1718,N_1465,N_1574);
or U1719 (N_1719,N_1495,N_1564);
nand U1720 (N_1720,N_1491,N_1474);
and U1721 (N_1721,N_1480,N_1495);
or U1722 (N_1722,N_1426,N_1428);
nand U1723 (N_1723,N_1578,N_1405);
and U1724 (N_1724,N_1504,N_1483);
and U1725 (N_1725,N_1583,N_1428);
nor U1726 (N_1726,N_1512,N_1499);
nor U1727 (N_1727,N_1509,N_1560);
nor U1728 (N_1728,N_1549,N_1431);
and U1729 (N_1729,N_1430,N_1484);
and U1730 (N_1730,N_1409,N_1510);
nand U1731 (N_1731,N_1482,N_1582);
or U1732 (N_1732,N_1586,N_1482);
nor U1733 (N_1733,N_1444,N_1483);
and U1734 (N_1734,N_1548,N_1493);
and U1735 (N_1735,N_1440,N_1401);
nor U1736 (N_1736,N_1592,N_1557);
or U1737 (N_1737,N_1429,N_1548);
nor U1738 (N_1738,N_1501,N_1525);
and U1739 (N_1739,N_1536,N_1545);
nor U1740 (N_1740,N_1522,N_1420);
nor U1741 (N_1741,N_1465,N_1593);
nor U1742 (N_1742,N_1592,N_1583);
nand U1743 (N_1743,N_1567,N_1527);
and U1744 (N_1744,N_1443,N_1444);
and U1745 (N_1745,N_1567,N_1459);
nand U1746 (N_1746,N_1474,N_1576);
and U1747 (N_1747,N_1461,N_1588);
nand U1748 (N_1748,N_1558,N_1588);
and U1749 (N_1749,N_1595,N_1457);
or U1750 (N_1750,N_1527,N_1429);
nand U1751 (N_1751,N_1459,N_1505);
nand U1752 (N_1752,N_1481,N_1566);
xnor U1753 (N_1753,N_1484,N_1491);
nand U1754 (N_1754,N_1575,N_1451);
nor U1755 (N_1755,N_1459,N_1599);
and U1756 (N_1756,N_1555,N_1441);
and U1757 (N_1757,N_1401,N_1437);
nor U1758 (N_1758,N_1594,N_1407);
nand U1759 (N_1759,N_1469,N_1407);
nor U1760 (N_1760,N_1401,N_1525);
or U1761 (N_1761,N_1508,N_1443);
or U1762 (N_1762,N_1531,N_1514);
and U1763 (N_1763,N_1563,N_1551);
nor U1764 (N_1764,N_1415,N_1433);
or U1765 (N_1765,N_1557,N_1492);
nor U1766 (N_1766,N_1452,N_1461);
nand U1767 (N_1767,N_1437,N_1426);
or U1768 (N_1768,N_1409,N_1438);
nand U1769 (N_1769,N_1478,N_1552);
or U1770 (N_1770,N_1589,N_1434);
and U1771 (N_1771,N_1425,N_1540);
or U1772 (N_1772,N_1445,N_1438);
nand U1773 (N_1773,N_1462,N_1489);
nor U1774 (N_1774,N_1491,N_1548);
nand U1775 (N_1775,N_1532,N_1474);
nand U1776 (N_1776,N_1543,N_1503);
nor U1777 (N_1777,N_1549,N_1421);
nand U1778 (N_1778,N_1435,N_1423);
or U1779 (N_1779,N_1496,N_1435);
nor U1780 (N_1780,N_1405,N_1419);
and U1781 (N_1781,N_1429,N_1598);
or U1782 (N_1782,N_1503,N_1531);
and U1783 (N_1783,N_1578,N_1552);
nor U1784 (N_1784,N_1552,N_1438);
and U1785 (N_1785,N_1595,N_1528);
and U1786 (N_1786,N_1556,N_1422);
and U1787 (N_1787,N_1589,N_1499);
or U1788 (N_1788,N_1476,N_1464);
nor U1789 (N_1789,N_1566,N_1424);
and U1790 (N_1790,N_1549,N_1457);
nor U1791 (N_1791,N_1432,N_1496);
nor U1792 (N_1792,N_1406,N_1558);
nor U1793 (N_1793,N_1514,N_1547);
nand U1794 (N_1794,N_1540,N_1413);
or U1795 (N_1795,N_1537,N_1433);
nand U1796 (N_1796,N_1548,N_1436);
nand U1797 (N_1797,N_1411,N_1419);
nand U1798 (N_1798,N_1515,N_1502);
nand U1799 (N_1799,N_1523,N_1545);
or U1800 (N_1800,N_1717,N_1764);
or U1801 (N_1801,N_1619,N_1759);
and U1802 (N_1802,N_1701,N_1645);
nor U1803 (N_1803,N_1635,N_1642);
and U1804 (N_1804,N_1602,N_1632);
or U1805 (N_1805,N_1622,N_1731);
nand U1806 (N_1806,N_1762,N_1739);
nor U1807 (N_1807,N_1725,N_1678);
xnor U1808 (N_1808,N_1721,N_1669);
or U1809 (N_1809,N_1750,N_1611);
and U1810 (N_1810,N_1748,N_1790);
and U1811 (N_1811,N_1778,N_1745);
nand U1812 (N_1812,N_1666,N_1636);
nor U1813 (N_1813,N_1641,N_1624);
nor U1814 (N_1814,N_1681,N_1785);
and U1815 (N_1815,N_1737,N_1646);
nor U1816 (N_1816,N_1792,N_1720);
or U1817 (N_1817,N_1671,N_1712);
nor U1818 (N_1818,N_1648,N_1728);
or U1819 (N_1819,N_1652,N_1699);
nand U1820 (N_1820,N_1679,N_1703);
nand U1821 (N_1821,N_1794,N_1664);
or U1822 (N_1822,N_1603,N_1796);
and U1823 (N_1823,N_1684,N_1628);
and U1824 (N_1824,N_1740,N_1688);
or U1825 (N_1825,N_1763,N_1707);
or U1826 (N_1826,N_1673,N_1694);
nor U1827 (N_1827,N_1676,N_1626);
or U1828 (N_1828,N_1781,N_1682);
nand U1829 (N_1829,N_1638,N_1798);
nor U1830 (N_1830,N_1734,N_1690);
nor U1831 (N_1831,N_1680,N_1747);
and U1832 (N_1832,N_1610,N_1647);
and U1833 (N_1833,N_1661,N_1605);
nand U1834 (N_1834,N_1663,N_1692);
nor U1835 (N_1835,N_1755,N_1746);
or U1836 (N_1836,N_1741,N_1633);
nand U1837 (N_1837,N_1713,N_1711);
nand U1838 (N_1838,N_1765,N_1616);
and U1839 (N_1839,N_1674,N_1650);
nor U1840 (N_1840,N_1771,N_1772);
and U1841 (N_1841,N_1716,N_1687);
nor U1842 (N_1842,N_1782,N_1758);
and U1843 (N_1843,N_1789,N_1608);
nand U1844 (N_1844,N_1686,N_1715);
or U1845 (N_1845,N_1620,N_1714);
and U1846 (N_1846,N_1651,N_1660);
or U1847 (N_1847,N_1787,N_1799);
or U1848 (N_1848,N_1606,N_1768);
nor U1849 (N_1849,N_1775,N_1735);
nor U1850 (N_1850,N_1793,N_1655);
or U1851 (N_1851,N_1777,N_1705);
or U1852 (N_1852,N_1662,N_1609);
nor U1853 (N_1853,N_1708,N_1742);
or U1854 (N_1854,N_1779,N_1629);
and U1855 (N_1855,N_1656,N_1723);
nor U1856 (N_1856,N_1640,N_1643);
and U1857 (N_1857,N_1791,N_1776);
or U1858 (N_1858,N_1697,N_1693);
and U1859 (N_1859,N_1700,N_1612);
or U1860 (N_1860,N_1780,N_1774);
or U1861 (N_1861,N_1730,N_1639);
and U1862 (N_1862,N_1753,N_1795);
and U1863 (N_1863,N_1627,N_1736);
nor U1864 (N_1864,N_1649,N_1767);
and U1865 (N_1865,N_1604,N_1657);
nor U1866 (N_1866,N_1786,N_1704);
or U1867 (N_1867,N_1600,N_1691);
or U1868 (N_1868,N_1788,N_1738);
or U1869 (N_1869,N_1769,N_1709);
nand U1870 (N_1870,N_1668,N_1695);
nand U1871 (N_1871,N_1770,N_1653);
or U1872 (N_1872,N_1757,N_1601);
nand U1873 (N_1873,N_1698,N_1743);
and U1874 (N_1874,N_1783,N_1710);
nor U1875 (N_1875,N_1634,N_1670);
or U1876 (N_1876,N_1761,N_1727);
nor U1877 (N_1877,N_1637,N_1702);
and U1878 (N_1878,N_1749,N_1667);
or U1879 (N_1879,N_1752,N_1754);
nor U1880 (N_1880,N_1726,N_1625);
nor U1881 (N_1881,N_1659,N_1654);
nand U1882 (N_1882,N_1706,N_1618);
nor U1883 (N_1883,N_1630,N_1672);
and U1884 (N_1884,N_1685,N_1724);
or U1885 (N_1885,N_1744,N_1617);
or U1886 (N_1886,N_1658,N_1623);
and U1887 (N_1887,N_1683,N_1766);
or U1888 (N_1888,N_1696,N_1631);
nor U1889 (N_1889,N_1718,N_1644);
and U1890 (N_1890,N_1722,N_1729);
nor U1891 (N_1891,N_1733,N_1719);
nor U1892 (N_1892,N_1760,N_1756);
nor U1893 (N_1893,N_1675,N_1621);
and U1894 (N_1894,N_1607,N_1751);
or U1895 (N_1895,N_1677,N_1614);
nand U1896 (N_1896,N_1689,N_1613);
nand U1897 (N_1897,N_1797,N_1615);
nor U1898 (N_1898,N_1732,N_1784);
and U1899 (N_1899,N_1773,N_1665);
nor U1900 (N_1900,N_1768,N_1713);
and U1901 (N_1901,N_1714,N_1651);
or U1902 (N_1902,N_1657,N_1701);
and U1903 (N_1903,N_1657,N_1625);
and U1904 (N_1904,N_1769,N_1749);
nor U1905 (N_1905,N_1740,N_1779);
and U1906 (N_1906,N_1619,N_1758);
nand U1907 (N_1907,N_1722,N_1797);
and U1908 (N_1908,N_1734,N_1780);
nor U1909 (N_1909,N_1673,N_1713);
nor U1910 (N_1910,N_1623,N_1619);
nor U1911 (N_1911,N_1696,N_1760);
and U1912 (N_1912,N_1643,N_1658);
and U1913 (N_1913,N_1698,N_1774);
or U1914 (N_1914,N_1720,N_1707);
or U1915 (N_1915,N_1717,N_1707);
nor U1916 (N_1916,N_1606,N_1634);
nor U1917 (N_1917,N_1686,N_1708);
or U1918 (N_1918,N_1643,N_1752);
or U1919 (N_1919,N_1616,N_1708);
nor U1920 (N_1920,N_1643,N_1691);
or U1921 (N_1921,N_1686,N_1774);
and U1922 (N_1922,N_1601,N_1705);
and U1923 (N_1923,N_1626,N_1775);
nor U1924 (N_1924,N_1737,N_1717);
nor U1925 (N_1925,N_1609,N_1673);
and U1926 (N_1926,N_1712,N_1641);
nand U1927 (N_1927,N_1701,N_1777);
nor U1928 (N_1928,N_1761,N_1759);
nor U1929 (N_1929,N_1630,N_1776);
nand U1930 (N_1930,N_1736,N_1700);
or U1931 (N_1931,N_1764,N_1663);
and U1932 (N_1932,N_1671,N_1685);
or U1933 (N_1933,N_1725,N_1680);
and U1934 (N_1934,N_1620,N_1631);
nand U1935 (N_1935,N_1674,N_1755);
nor U1936 (N_1936,N_1689,N_1771);
or U1937 (N_1937,N_1675,N_1656);
or U1938 (N_1938,N_1777,N_1746);
nand U1939 (N_1939,N_1724,N_1792);
nor U1940 (N_1940,N_1630,N_1675);
nand U1941 (N_1941,N_1744,N_1775);
and U1942 (N_1942,N_1608,N_1621);
nand U1943 (N_1943,N_1611,N_1745);
nor U1944 (N_1944,N_1658,N_1682);
or U1945 (N_1945,N_1776,N_1775);
nand U1946 (N_1946,N_1707,N_1769);
and U1947 (N_1947,N_1680,N_1682);
or U1948 (N_1948,N_1635,N_1737);
and U1949 (N_1949,N_1603,N_1671);
or U1950 (N_1950,N_1673,N_1607);
nor U1951 (N_1951,N_1719,N_1688);
or U1952 (N_1952,N_1655,N_1648);
or U1953 (N_1953,N_1774,N_1772);
nand U1954 (N_1954,N_1743,N_1657);
and U1955 (N_1955,N_1705,N_1608);
or U1956 (N_1956,N_1689,N_1678);
nand U1957 (N_1957,N_1635,N_1628);
nand U1958 (N_1958,N_1776,N_1689);
or U1959 (N_1959,N_1670,N_1725);
nand U1960 (N_1960,N_1632,N_1795);
nor U1961 (N_1961,N_1722,N_1761);
nand U1962 (N_1962,N_1773,N_1733);
and U1963 (N_1963,N_1715,N_1763);
and U1964 (N_1964,N_1760,N_1783);
nor U1965 (N_1965,N_1730,N_1790);
or U1966 (N_1966,N_1791,N_1674);
or U1967 (N_1967,N_1608,N_1638);
or U1968 (N_1968,N_1783,N_1743);
nor U1969 (N_1969,N_1737,N_1638);
nor U1970 (N_1970,N_1606,N_1741);
nand U1971 (N_1971,N_1683,N_1705);
and U1972 (N_1972,N_1766,N_1621);
nand U1973 (N_1973,N_1754,N_1732);
nand U1974 (N_1974,N_1643,N_1606);
and U1975 (N_1975,N_1622,N_1667);
nor U1976 (N_1976,N_1791,N_1757);
nand U1977 (N_1977,N_1786,N_1774);
nor U1978 (N_1978,N_1774,N_1676);
nor U1979 (N_1979,N_1703,N_1795);
and U1980 (N_1980,N_1622,N_1608);
or U1981 (N_1981,N_1797,N_1686);
nand U1982 (N_1982,N_1722,N_1719);
nand U1983 (N_1983,N_1699,N_1615);
nand U1984 (N_1984,N_1731,N_1667);
nor U1985 (N_1985,N_1607,N_1694);
or U1986 (N_1986,N_1739,N_1607);
nand U1987 (N_1987,N_1623,N_1666);
nor U1988 (N_1988,N_1717,N_1791);
xor U1989 (N_1989,N_1693,N_1646);
and U1990 (N_1990,N_1636,N_1767);
or U1991 (N_1991,N_1701,N_1619);
and U1992 (N_1992,N_1616,N_1782);
nand U1993 (N_1993,N_1669,N_1709);
nand U1994 (N_1994,N_1672,N_1736);
nand U1995 (N_1995,N_1622,N_1710);
nand U1996 (N_1996,N_1654,N_1771);
or U1997 (N_1997,N_1785,N_1731);
nand U1998 (N_1998,N_1781,N_1732);
and U1999 (N_1999,N_1742,N_1625);
nand U2000 (N_2000,N_1883,N_1813);
nor U2001 (N_2001,N_1902,N_1833);
nor U2002 (N_2002,N_1839,N_1949);
and U2003 (N_2003,N_1928,N_1858);
nand U2004 (N_2004,N_1952,N_1885);
nor U2005 (N_2005,N_1896,N_1984);
nand U2006 (N_2006,N_1867,N_1815);
and U2007 (N_2007,N_1843,N_1936);
nand U2008 (N_2008,N_1830,N_1929);
nand U2009 (N_2009,N_1947,N_1802);
or U2010 (N_2010,N_1860,N_1958);
nor U2011 (N_2011,N_1868,N_1857);
xor U2012 (N_2012,N_1835,N_1842);
nand U2013 (N_2013,N_1809,N_1906);
nand U2014 (N_2014,N_1878,N_1898);
nand U2015 (N_2015,N_1903,N_1811);
and U2016 (N_2016,N_1998,N_1950);
nand U2017 (N_2017,N_1986,N_1924);
and U2018 (N_2018,N_1819,N_1828);
and U2019 (N_2019,N_1816,N_1920);
and U2020 (N_2020,N_1800,N_1988);
or U2021 (N_2021,N_1915,N_1869);
nand U2022 (N_2022,N_1944,N_1969);
nand U2023 (N_2023,N_1983,N_1873);
nand U2024 (N_2024,N_1976,N_1836);
xor U2025 (N_2025,N_1980,N_1937);
nor U2026 (N_2026,N_1822,N_1901);
nor U2027 (N_2027,N_1957,N_1967);
nand U2028 (N_2028,N_1848,N_1912);
and U2029 (N_2029,N_1991,N_1914);
or U2030 (N_2030,N_1977,N_1876);
nor U2031 (N_2031,N_1872,N_1810);
or U2032 (N_2032,N_1890,N_1817);
nand U2033 (N_2033,N_1993,N_1852);
nor U2034 (N_2034,N_1863,N_1849);
and U2035 (N_2035,N_1905,N_1908);
nand U2036 (N_2036,N_1882,N_1973);
and U2037 (N_2037,N_1968,N_1910);
or U2038 (N_2038,N_1943,N_1922);
nand U2039 (N_2039,N_1856,N_1820);
and U2040 (N_2040,N_1826,N_1989);
and U2041 (N_2041,N_1994,N_1894);
or U2042 (N_2042,N_1909,N_1891);
nor U2043 (N_2043,N_1844,N_1925);
or U2044 (N_2044,N_1970,N_1824);
nand U2045 (N_2045,N_1948,N_1861);
or U2046 (N_2046,N_1854,N_1917);
nor U2047 (N_2047,N_1982,N_1801);
and U2048 (N_2048,N_1840,N_1961);
or U2049 (N_2049,N_1934,N_1834);
nor U2050 (N_2050,N_1975,N_1847);
and U2051 (N_2051,N_1808,N_1942);
nand U2052 (N_2052,N_1837,N_1907);
or U2053 (N_2053,N_1818,N_1827);
or U2054 (N_2054,N_1879,N_1846);
and U2055 (N_2055,N_1951,N_1965);
nand U2056 (N_2056,N_1874,N_1823);
and U2057 (N_2057,N_1803,N_1832);
and U2058 (N_2058,N_1866,N_1918);
and U2059 (N_2059,N_1851,N_1990);
and U2060 (N_2060,N_1995,N_1978);
or U2061 (N_2061,N_1865,N_1931);
nor U2062 (N_2062,N_1881,N_1845);
nand U2063 (N_2063,N_1953,N_1812);
and U2064 (N_2064,N_1859,N_1877);
and U2065 (N_2065,N_1913,N_1959);
or U2066 (N_2066,N_1900,N_1954);
nand U2067 (N_2067,N_1895,N_1938);
nor U2068 (N_2068,N_1940,N_1966);
and U2069 (N_2069,N_1932,N_1825);
nor U2070 (N_2070,N_1855,N_1875);
and U2071 (N_2071,N_1999,N_1829);
or U2072 (N_2072,N_1871,N_1979);
and U2073 (N_2073,N_1939,N_1880);
nand U2074 (N_2074,N_1971,N_1946);
nand U2075 (N_2075,N_1892,N_1972);
nor U2076 (N_2076,N_1956,N_1911);
and U2077 (N_2077,N_1850,N_1974);
nand U2078 (N_2078,N_1889,N_1821);
nor U2079 (N_2079,N_1807,N_1996);
and U2080 (N_2080,N_1945,N_1888);
nand U2081 (N_2081,N_1992,N_1930);
and U2082 (N_2082,N_1893,N_1985);
nor U2083 (N_2083,N_1960,N_1805);
or U2084 (N_2084,N_1933,N_1916);
nor U2085 (N_2085,N_1981,N_1804);
and U2086 (N_2086,N_1919,N_1962);
or U2087 (N_2087,N_1899,N_1870);
nand U2088 (N_2088,N_1886,N_1831);
nand U2089 (N_2089,N_1841,N_1838);
and U2090 (N_2090,N_1862,N_1923);
and U2091 (N_2091,N_1884,N_1853);
or U2092 (N_2092,N_1955,N_1926);
or U2093 (N_2093,N_1864,N_1921);
nor U2094 (N_2094,N_1964,N_1806);
or U2095 (N_2095,N_1814,N_1935);
and U2096 (N_2096,N_1997,N_1927);
or U2097 (N_2097,N_1897,N_1904);
and U2098 (N_2098,N_1941,N_1963);
nor U2099 (N_2099,N_1987,N_1887);
nor U2100 (N_2100,N_1827,N_1970);
or U2101 (N_2101,N_1881,N_1862);
and U2102 (N_2102,N_1901,N_1965);
nor U2103 (N_2103,N_1967,N_1865);
nand U2104 (N_2104,N_1892,N_1926);
nor U2105 (N_2105,N_1894,N_1931);
nand U2106 (N_2106,N_1863,N_1916);
and U2107 (N_2107,N_1966,N_1912);
nor U2108 (N_2108,N_1924,N_1973);
nand U2109 (N_2109,N_1841,N_1844);
nand U2110 (N_2110,N_1873,N_1995);
nor U2111 (N_2111,N_1920,N_1940);
or U2112 (N_2112,N_1832,N_1810);
nand U2113 (N_2113,N_1949,N_1907);
nor U2114 (N_2114,N_1984,N_1879);
or U2115 (N_2115,N_1929,N_1828);
nand U2116 (N_2116,N_1832,N_1872);
or U2117 (N_2117,N_1938,N_1974);
nand U2118 (N_2118,N_1933,N_1883);
or U2119 (N_2119,N_1847,N_1851);
and U2120 (N_2120,N_1955,N_1811);
nand U2121 (N_2121,N_1877,N_1871);
or U2122 (N_2122,N_1983,N_1971);
nand U2123 (N_2123,N_1923,N_1931);
or U2124 (N_2124,N_1941,N_1967);
nor U2125 (N_2125,N_1835,N_1830);
nor U2126 (N_2126,N_1998,N_1893);
nand U2127 (N_2127,N_1977,N_1819);
nor U2128 (N_2128,N_1806,N_1949);
nand U2129 (N_2129,N_1984,N_1935);
nor U2130 (N_2130,N_1815,N_1903);
or U2131 (N_2131,N_1852,N_1909);
nor U2132 (N_2132,N_1992,N_1947);
or U2133 (N_2133,N_1850,N_1824);
or U2134 (N_2134,N_1914,N_1949);
nand U2135 (N_2135,N_1992,N_1951);
and U2136 (N_2136,N_1828,N_1940);
nand U2137 (N_2137,N_1942,N_1839);
nor U2138 (N_2138,N_1817,N_1808);
and U2139 (N_2139,N_1813,N_1922);
nor U2140 (N_2140,N_1974,N_1972);
nor U2141 (N_2141,N_1906,N_1850);
nor U2142 (N_2142,N_1848,N_1868);
nand U2143 (N_2143,N_1838,N_1880);
nor U2144 (N_2144,N_1961,N_1851);
and U2145 (N_2145,N_1867,N_1900);
or U2146 (N_2146,N_1927,N_1921);
nand U2147 (N_2147,N_1998,N_1887);
or U2148 (N_2148,N_1833,N_1873);
and U2149 (N_2149,N_1843,N_1846);
nor U2150 (N_2150,N_1960,N_1947);
nand U2151 (N_2151,N_1866,N_1814);
or U2152 (N_2152,N_1845,N_1972);
nand U2153 (N_2153,N_1970,N_1801);
and U2154 (N_2154,N_1927,N_1869);
nand U2155 (N_2155,N_1829,N_1946);
or U2156 (N_2156,N_1933,N_1850);
or U2157 (N_2157,N_1989,N_1889);
or U2158 (N_2158,N_1936,N_1959);
and U2159 (N_2159,N_1934,N_1819);
nand U2160 (N_2160,N_1888,N_1904);
nand U2161 (N_2161,N_1936,N_1892);
and U2162 (N_2162,N_1871,N_1874);
or U2163 (N_2163,N_1906,N_1916);
nand U2164 (N_2164,N_1983,N_1810);
nand U2165 (N_2165,N_1929,N_1945);
nor U2166 (N_2166,N_1971,N_1823);
xnor U2167 (N_2167,N_1808,N_1898);
nor U2168 (N_2168,N_1805,N_1821);
nand U2169 (N_2169,N_1921,N_1817);
nand U2170 (N_2170,N_1839,N_1983);
and U2171 (N_2171,N_1929,N_1959);
or U2172 (N_2172,N_1967,N_1973);
nor U2173 (N_2173,N_1893,N_1861);
nor U2174 (N_2174,N_1929,N_1878);
and U2175 (N_2175,N_1933,N_1855);
and U2176 (N_2176,N_1908,N_1874);
or U2177 (N_2177,N_1862,N_1921);
nor U2178 (N_2178,N_1829,N_1904);
nand U2179 (N_2179,N_1888,N_1995);
nor U2180 (N_2180,N_1958,N_1825);
nor U2181 (N_2181,N_1906,N_1903);
nor U2182 (N_2182,N_1820,N_1862);
and U2183 (N_2183,N_1874,N_1878);
or U2184 (N_2184,N_1978,N_1853);
nor U2185 (N_2185,N_1923,N_1951);
or U2186 (N_2186,N_1820,N_1919);
nor U2187 (N_2187,N_1820,N_1941);
or U2188 (N_2188,N_1971,N_1812);
and U2189 (N_2189,N_1816,N_1980);
nor U2190 (N_2190,N_1813,N_1828);
and U2191 (N_2191,N_1853,N_1802);
nand U2192 (N_2192,N_1899,N_1902);
or U2193 (N_2193,N_1979,N_1984);
nor U2194 (N_2194,N_1846,N_1985);
or U2195 (N_2195,N_1981,N_1985);
nand U2196 (N_2196,N_1894,N_1868);
or U2197 (N_2197,N_1872,N_1954);
or U2198 (N_2198,N_1968,N_1920);
nand U2199 (N_2199,N_1887,N_1835);
nand U2200 (N_2200,N_2158,N_2051);
or U2201 (N_2201,N_2109,N_2135);
or U2202 (N_2202,N_2008,N_2151);
or U2203 (N_2203,N_2176,N_2027);
nor U2204 (N_2204,N_2056,N_2016);
nand U2205 (N_2205,N_2002,N_2029);
xor U2206 (N_2206,N_2015,N_2144);
nand U2207 (N_2207,N_2065,N_2044);
and U2208 (N_2208,N_2184,N_2145);
or U2209 (N_2209,N_2067,N_2122);
or U2210 (N_2210,N_2028,N_2148);
nand U2211 (N_2211,N_2149,N_2037);
or U2212 (N_2212,N_2115,N_2170);
nor U2213 (N_2213,N_2172,N_2022);
and U2214 (N_2214,N_2023,N_2078);
or U2215 (N_2215,N_2025,N_2005);
nor U2216 (N_2216,N_2179,N_2031);
xnor U2217 (N_2217,N_2033,N_2053);
nand U2218 (N_2218,N_2075,N_2123);
nand U2219 (N_2219,N_2134,N_2105);
or U2220 (N_2220,N_2108,N_2038);
or U2221 (N_2221,N_2054,N_2159);
and U2222 (N_2222,N_2011,N_2048);
nand U2223 (N_2223,N_2086,N_2113);
nand U2224 (N_2224,N_2128,N_2154);
and U2225 (N_2225,N_2132,N_2024);
nor U2226 (N_2226,N_2018,N_2131);
and U2227 (N_2227,N_2125,N_2100);
nor U2228 (N_2228,N_2082,N_2163);
nor U2229 (N_2229,N_2068,N_2007);
or U2230 (N_2230,N_2155,N_2116);
and U2231 (N_2231,N_2032,N_2177);
nor U2232 (N_2232,N_2187,N_2041);
nand U2233 (N_2233,N_2000,N_2112);
and U2234 (N_2234,N_2142,N_2169);
nor U2235 (N_2235,N_2020,N_2039);
and U2236 (N_2236,N_2106,N_2140);
nor U2237 (N_2237,N_2081,N_2175);
or U2238 (N_2238,N_2182,N_2045);
nor U2239 (N_2239,N_2114,N_2192);
nor U2240 (N_2240,N_2070,N_2139);
or U2241 (N_2241,N_2061,N_2183);
or U2242 (N_2242,N_2127,N_2097);
or U2243 (N_2243,N_2107,N_2003);
nand U2244 (N_2244,N_2193,N_2058);
nor U2245 (N_2245,N_2186,N_2143);
or U2246 (N_2246,N_2174,N_2077);
nand U2247 (N_2247,N_2196,N_2060);
nand U2248 (N_2248,N_2085,N_2066);
nor U2249 (N_2249,N_2059,N_2188);
nand U2250 (N_2250,N_2156,N_2194);
or U2251 (N_2251,N_2117,N_2161);
or U2252 (N_2252,N_2035,N_2057);
nand U2253 (N_2253,N_2090,N_2043);
or U2254 (N_2254,N_2167,N_2093);
nor U2255 (N_2255,N_2042,N_2168);
nor U2256 (N_2256,N_2120,N_2162);
nand U2257 (N_2257,N_2195,N_2083);
nand U2258 (N_2258,N_2034,N_2055);
xnor U2259 (N_2259,N_2040,N_2137);
nor U2260 (N_2260,N_2036,N_2073);
and U2261 (N_2261,N_2017,N_2198);
nand U2262 (N_2262,N_2084,N_2052);
nor U2263 (N_2263,N_2178,N_2124);
nor U2264 (N_2264,N_2129,N_2152);
nor U2265 (N_2265,N_2092,N_2050);
nor U2266 (N_2266,N_2133,N_2010);
nand U2267 (N_2267,N_2180,N_2103);
nand U2268 (N_2268,N_2080,N_2079);
nor U2269 (N_2269,N_2104,N_2088);
nor U2270 (N_2270,N_2001,N_2098);
nor U2271 (N_2271,N_2166,N_2064);
nand U2272 (N_2272,N_2019,N_2138);
and U2273 (N_2273,N_2189,N_2130);
or U2274 (N_2274,N_2074,N_2096);
xor U2275 (N_2275,N_2102,N_2095);
nor U2276 (N_2276,N_2047,N_2069);
and U2277 (N_2277,N_2190,N_2091);
nor U2278 (N_2278,N_2006,N_2099);
nand U2279 (N_2279,N_2121,N_2119);
and U2280 (N_2280,N_2199,N_2181);
nor U2281 (N_2281,N_2173,N_2147);
nor U2282 (N_2282,N_2160,N_2063);
nand U2283 (N_2283,N_2165,N_2089);
nor U2284 (N_2284,N_2013,N_2004);
nand U2285 (N_2285,N_2111,N_2094);
nor U2286 (N_2286,N_2046,N_2141);
or U2287 (N_2287,N_2021,N_2071);
and U2288 (N_2288,N_2087,N_2126);
and U2289 (N_2289,N_2191,N_2009);
xnor U2290 (N_2290,N_2118,N_2076);
or U2291 (N_2291,N_2153,N_2101);
or U2292 (N_2292,N_2030,N_2171);
or U2293 (N_2293,N_2014,N_2026);
or U2294 (N_2294,N_2197,N_2136);
nor U2295 (N_2295,N_2110,N_2150);
and U2296 (N_2296,N_2146,N_2012);
nand U2297 (N_2297,N_2185,N_2072);
nor U2298 (N_2298,N_2062,N_2049);
and U2299 (N_2299,N_2164,N_2157);
nand U2300 (N_2300,N_2094,N_2172);
or U2301 (N_2301,N_2115,N_2004);
nor U2302 (N_2302,N_2198,N_2098);
and U2303 (N_2303,N_2172,N_2047);
or U2304 (N_2304,N_2011,N_2080);
or U2305 (N_2305,N_2190,N_2165);
and U2306 (N_2306,N_2148,N_2150);
nand U2307 (N_2307,N_2177,N_2068);
xor U2308 (N_2308,N_2130,N_2135);
nor U2309 (N_2309,N_2146,N_2021);
nor U2310 (N_2310,N_2023,N_2177);
nand U2311 (N_2311,N_2178,N_2108);
and U2312 (N_2312,N_2154,N_2183);
and U2313 (N_2313,N_2006,N_2067);
nor U2314 (N_2314,N_2035,N_2170);
nor U2315 (N_2315,N_2016,N_2078);
nand U2316 (N_2316,N_2044,N_2093);
and U2317 (N_2317,N_2041,N_2004);
and U2318 (N_2318,N_2032,N_2142);
and U2319 (N_2319,N_2171,N_2137);
and U2320 (N_2320,N_2168,N_2185);
nor U2321 (N_2321,N_2010,N_2165);
nor U2322 (N_2322,N_2023,N_2124);
nor U2323 (N_2323,N_2162,N_2082);
or U2324 (N_2324,N_2094,N_2006);
nor U2325 (N_2325,N_2065,N_2069);
nor U2326 (N_2326,N_2192,N_2164);
nand U2327 (N_2327,N_2017,N_2118);
and U2328 (N_2328,N_2180,N_2156);
and U2329 (N_2329,N_2184,N_2048);
nand U2330 (N_2330,N_2011,N_2161);
nand U2331 (N_2331,N_2122,N_2148);
or U2332 (N_2332,N_2025,N_2082);
nand U2333 (N_2333,N_2107,N_2016);
and U2334 (N_2334,N_2140,N_2129);
nor U2335 (N_2335,N_2039,N_2178);
and U2336 (N_2336,N_2120,N_2066);
and U2337 (N_2337,N_2133,N_2035);
or U2338 (N_2338,N_2074,N_2106);
nand U2339 (N_2339,N_2127,N_2150);
nand U2340 (N_2340,N_2165,N_2000);
or U2341 (N_2341,N_2034,N_2056);
nand U2342 (N_2342,N_2090,N_2124);
or U2343 (N_2343,N_2100,N_2140);
or U2344 (N_2344,N_2151,N_2045);
or U2345 (N_2345,N_2004,N_2071);
and U2346 (N_2346,N_2033,N_2052);
nor U2347 (N_2347,N_2154,N_2032);
nor U2348 (N_2348,N_2153,N_2149);
nand U2349 (N_2349,N_2167,N_2104);
nor U2350 (N_2350,N_2117,N_2198);
or U2351 (N_2351,N_2001,N_2060);
nand U2352 (N_2352,N_2103,N_2143);
and U2353 (N_2353,N_2002,N_2136);
nand U2354 (N_2354,N_2106,N_2028);
and U2355 (N_2355,N_2022,N_2045);
nand U2356 (N_2356,N_2193,N_2101);
nor U2357 (N_2357,N_2102,N_2003);
nand U2358 (N_2358,N_2158,N_2175);
and U2359 (N_2359,N_2057,N_2081);
and U2360 (N_2360,N_2008,N_2092);
or U2361 (N_2361,N_2199,N_2115);
nand U2362 (N_2362,N_2028,N_2184);
or U2363 (N_2363,N_2167,N_2053);
or U2364 (N_2364,N_2049,N_2199);
or U2365 (N_2365,N_2032,N_2078);
or U2366 (N_2366,N_2180,N_2020);
nand U2367 (N_2367,N_2064,N_2042);
nor U2368 (N_2368,N_2101,N_2132);
nand U2369 (N_2369,N_2074,N_2052);
nor U2370 (N_2370,N_2008,N_2037);
nand U2371 (N_2371,N_2019,N_2014);
and U2372 (N_2372,N_2132,N_2148);
nor U2373 (N_2373,N_2032,N_2131);
nand U2374 (N_2374,N_2115,N_2133);
or U2375 (N_2375,N_2026,N_2102);
or U2376 (N_2376,N_2186,N_2153);
or U2377 (N_2377,N_2170,N_2124);
nor U2378 (N_2378,N_2043,N_2049);
and U2379 (N_2379,N_2044,N_2103);
and U2380 (N_2380,N_2128,N_2151);
and U2381 (N_2381,N_2184,N_2185);
and U2382 (N_2382,N_2150,N_2006);
nand U2383 (N_2383,N_2105,N_2006);
and U2384 (N_2384,N_2197,N_2004);
nor U2385 (N_2385,N_2182,N_2005);
and U2386 (N_2386,N_2184,N_2057);
nand U2387 (N_2387,N_2084,N_2083);
or U2388 (N_2388,N_2173,N_2015);
nor U2389 (N_2389,N_2156,N_2117);
or U2390 (N_2390,N_2106,N_2158);
and U2391 (N_2391,N_2009,N_2105);
nor U2392 (N_2392,N_2069,N_2026);
and U2393 (N_2393,N_2192,N_2061);
and U2394 (N_2394,N_2063,N_2070);
and U2395 (N_2395,N_2166,N_2000);
or U2396 (N_2396,N_2050,N_2188);
nand U2397 (N_2397,N_2199,N_2198);
or U2398 (N_2398,N_2047,N_2150);
and U2399 (N_2399,N_2079,N_2041);
and U2400 (N_2400,N_2312,N_2263);
and U2401 (N_2401,N_2292,N_2393);
nor U2402 (N_2402,N_2298,N_2359);
nand U2403 (N_2403,N_2234,N_2358);
nor U2404 (N_2404,N_2394,N_2200);
and U2405 (N_2405,N_2217,N_2332);
nand U2406 (N_2406,N_2366,N_2259);
nand U2407 (N_2407,N_2255,N_2220);
or U2408 (N_2408,N_2346,N_2275);
and U2409 (N_2409,N_2376,N_2384);
xnor U2410 (N_2410,N_2385,N_2354);
nand U2411 (N_2411,N_2214,N_2386);
and U2412 (N_2412,N_2301,N_2308);
and U2413 (N_2413,N_2342,N_2328);
nor U2414 (N_2414,N_2233,N_2203);
nor U2415 (N_2415,N_2283,N_2237);
and U2416 (N_2416,N_2262,N_2293);
or U2417 (N_2417,N_2221,N_2218);
nand U2418 (N_2418,N_2258,N_2270);
nor U2419 (N_2419,N_2364,N_2363);
nand U2420 (N_2420,N_2336,N_2252);
and U2421 (N_2421,N_2339,N_2333);
or U2422 (N_2422,N_2313,N_2287);
nand U2423 (N_2423,N_2323,N_2261);
and U2424 (N_2424,N_2243,N_2369);
nand U2425 (N_2425,N_2201,N_2368);
nand U2426 (N_2426,N_2397,N_2314);
nand U2427 (N_2427,N_2331,N_2238);
nor U2428 (N_2428,N_2230,N_2294);
and U2429 (N_2429,N_2399,N_2390);
nor U2430 (N_2430,N_2373,N_2340);
and U2431 (N_2431,N_2318,N_2334);
nor U2432 (N_2432,N_2246,N_2272);
nand U2433 (N_2433,N_2251,N_2355);
nand U2434 (N_2434,N_2360,N_2254);
nor U2435 (N_2435,N_2225,N_2326);
or U2436 (N_2436,N_2281,N_2387);
and U2437 (N_2437,N_2351,N_2231);
or U2438 (N_2438,N_2365,N_2267);
and U2439 (N_2439,N_2296,N_2232);
and U2440 (N_2440,N_2242,N_2250);
and U2441 (N_2441,N_2215,N_2377);
nor U2442 (N_2442,N_2257,N_2286);
or U2443 (N_2443,N_2317,N_2395);
and U2444 (N_2444,N_2343,N_2219);
and U2445 (N_2445,N_2260,N_2362);
nor U2446 (N_2446,N_2239,N_2303);
nor U2447 (N_2447,N_2266,N_2356);
or U2448 (N_2448,N_2227,N_2309);
nor U2449 (N_2449,N_2380,N_2278);
and U2450 (N_2450,N_2273,N_2226);
and U2451 (N_2451,N_2277,N_2335);
nand U2452 (N_2452,N_2322,N_2256);
or U2453 (N_2453,N_2388,N_2229);
and U2454 (N_2454,N_2271,N_2327);
and U2455 (N_2455,N_2265,N_2315);
nand U2456 (N_2456,N_2341,N_2321);
nand U2457 (N_2457,N_2371,N_2381);
and U2458 (N_2458,N_2320,N_2374);
nor U2459 (N_2459,N_2224,N_2204);
nor U2460 (N_2460,N_2205,N_2269);
and U2461 (N_2461,N_2391,N_2357);
nor U2462 (N_2462,N_2383,N_2302);
or U2463 (N_2463,N_2291,N_2244);
xor U2464 (N_2464,N_2382,N_2241);
xnor U2465 (N_2465,N_2347,N_2253);
nor U2466 (N_2466,N_2280,N_2316);
nand U2467 (N_2467,N_2350,N_2311);
and U2468 (N_2468,N_2361,N_2211);
nand U2469 (N_2469,N_2249,N_2213);
or U2470 (N_2470,N_2299,N_2338);
and U2471 (N_2471,N_2370,N_2389);
nand U2472 (N_2472,N_2398,N_2367);
nand U2473 (N_2473,N_2274,N_2236);
and U2474 (N_2474,N_2348,N_2206);
nor U2475 (N_2475,N_2349,N_2288);
or U2476 (N_2476,N_2290,N_2329);
nor U2477 (N_2477,N_2216,N_2297);
or U2478 (N_2478,N_2222,N_2212);
or U2479 (N_2479,N_2247,N_2396);
nand U2480 (N_2480,N_2209,N_2248);
or U2481 (N_2481,N_2324,N_2228);
nand U2482 (N_2482,N_2337,N_2240);
nor U2483 (N_2483,N_2392,N_2276);
or U2484 (N_2484,N_2300,N_2325);
or U2485 (N_2485,N_2310,N_2345);
or U2486 (N_2486,N_2264,N_2306);
and U2487 (N_2487,N_2330,N_2352);
nand U2488 (N_2488,N_2319,N_2279);
and U2489 (N_2489,N_2245,N_2235);
nand U2490 (N_2490,N_2282,N_2268);
nor U2491 (N_2491,N_2353,N_2207);
or U2492 (N_2492,N_2210,N_2378);
nor U2493 (N_2493,N_2375,N_2379);
or U2494 (N_2494,N_2305,N_2284);
or U2495 (N_2495,N_2372,N_2223);
nand U2496 (N_2496,N_2307,N_2344);
and U2497 (N_2497,N_2208,N_2285);
or U2498 (N_2498,N_2289,N_2202);
and U2499 (N_2499,N_2295,N_2304);
and U2500 (N_2500,N_2365,N_2251);
and U2501 (N_2501,N_2308,N_2312);
nand U2502 (N_2502,N_2220,N_2369);
or U2503 (N_2503,N_2208,N_2333);
nand U2504 (N_2504,N_2262,N_2278);
nand U2505 (N_2505,N_2365,N_2367);
and U2506 (N_2506,N_2354,N_2399);
or U2507 (N_2507,N_2207,N_2382);
nor U2508 (N_2508,N_2290,N_2241);
nand U2509 (N_2509,N_2380,N_2327);
nor U2510 (N_2510,N_2256,N_2350);
nand U2511 (N_2511,N_2236,N_2399);
or U2512 (N_2512,N_2252,N_2274);
nor U2513 (N_2513,N_2349,N_2272);
nor U2514 (N_2514,N_2353,N_2259);
nand U2515 (N_2515,N_2269,N_2313);
nand U2516 (N_2516,N_2319,N_2233);
or U2517 (N_2517,N_2246,N_2363);
nand U2518 (N_2518,N_2381,N_2203);
nor U2519 (N_2519,N_2233,N_2310);
nand U2520 (N_2520,N_2299,N_2324);
nand U2521 (N_2521,N_2340,N_2228);
nor U2522 (N_2522,N_2301,N_2392);
or U2523 (N_2523,N_2356,N_2352);
and U2524 (N_2524,N_2201,N_2231);
and U2525 (N_2525,N_2338,N_2314);
nor U2526 (N_2526,N_2271,N_2264);
or U2527 (N_2527,N_2232,N_2388);
or U2528 (N_2528,N_2369,N_2398);
nor U2529 (N_2529,N_2222,N_2219);
nand U2530 (N_2530,N_2386,N_2380);
nand U2531 (N_2531,N_2245,N_2218);
nand U2532 (N_2532,N_2266,N_2204);
nand U2533 (N_2533,N_2367,N_2394);
nand U2534 (N_2534,N_2338,N_2234);
nor U2535 (N_2535,N_2319,N_2313);
and U2536 (N_2536,N_2365,N_2201);
and U2537 (N_2537,N_2289,N_2256);
or U2538 (N_2538,N_2213,N_2209);
and U2539 (N_2539,N_2236,N_2258);
nor U2540 (N_2540,N_2315,N_2258);
and U2541 (N_2541,N_2230,N_2254);
and U2542 (N_2542,N_2370,N_2261);
or U2543 (N_2543,N_2271,N_2212);
nor U2544 (N_2544,N_2323,N_2281);
nor U2545 (N_2545,N_2383,N_2397);
or U2546 (N_2546,N_2281,N_2376);
nand U2547 (N_2547,N_2364,N_2204);
nor U2548 (N_2548,N_2381,N_2383);
nand U2549 (N_2549,N_2355,N_2316);
or U2550 (N_2550,N_2240,N_2221);
and U2551 (N_2551,N_2373,N_2293);
nand U2552 (N_2552,N_2374,N_2219);
nor U2553 (N_2553,N_2311,N_2303);
nor U2554 (N_2554,N_2205,N_2335);
nor U2555 (N_2555,N_2303,N_2314);
or U2556 (N_2556,N_2229,N_2329);
nand U2557 (N_2557,N_2284,N_2234);
nand U2558 (N_2558,N_2261,N_2203);
nand U2559 (N_2559,N_2257,N_2246);
and U2560 (N_2560,N_2314,N_2328);
or U2561 (N_2561,N_2307,N_2336);
nand U2562 (N_2562,N_2379,N_2358);
nor U2563 (N_2563,N_2306,N_2293);
and U2564 (N_2564,N_2277,N_2253);
nor U2565 (N_2565,N_2233,N_2261);
or U2566 (N_2566,N_2233,N_2262);
nor U2567 (N_2567,N_2328,N_2344);
nand U2568 (N_2568,N_2268,N_2399);
or U2569 (N_2569,N_2341,N_2273);
and U2570 (N_2570,N_2285,N_2228);
nor U2571 (N_2571,N_2270,N_2241);
and U2572 (N_2572,N_2302,N_2300);
and U2573 (N_2573,N_2233,N_2301);
and U2574 (N_2574,N_2286,N_2334);
nor U2575 (N_2575,N_2213,N_2370);
nand U2576 (N_2576,N_2251,N_2347);
nand U2577 (N_2577,N_2235,N_2271);
nand U2578 (N_2578,N_2337,N_2273);
nor U2579 (N_2579,N_2289,N_2379);
or U2580 (N_2580,N_2203,N_2382);
or U2581 (N_2581,N_2365,N_2376);
xor U2582 (N_2582,N_2373,N_2237);
nor U2583 (N_2583,N_2372,N_2269);
and U2584 (N_2584,N_2293,N_2389);
nor U2585 (N_2585,N_2200,N_2259);
nand U2586 (N_2586,N_2298,N_2329);
nand U2587 (N_2587,N_2331,N_2305);
nand U2588 (N_2588,N_2224,N_2229);
and U2589 (N_2589,N_2234,N_2272);
and U2590 (N_2590,N_2273,N_2382);
and U2591 (N_2591,N_2315,N_2350);
and U2592 (N_2592,N_2321,N_2324);
or U2593 (N_2593,N_2307,N_2380);
nand U2594 (N_2594,N_2224,N_2271);
and U2595 (N_2595,N_2378,N_2220);
or U2596 (N_2596,N_2397,N_2218);
or U2597 (N_2597,N_2208,N_2382);
or U2598 (N_2598,N_2249,N_2227);
nand U2599 (N_2599,N_2338,N_2369);
nand U2600 (N_2600,N_2595,N_2462);
nand U2601 (N_2601,N_2411,N_2469);
or U2602 (N_2602,N_2549,N_2483);
or U2603 (N_2603,N_2400,N_2529);
and U2604 (N_2604,N_2495,N_2526);
and U2605 (N_2605,N_2512,N_2570);
nor U2606 (N_2606,N_2584,N_2471);
nor U2607 (N_2607,N_2556,N_2456);
nand U2608 (N_2608,N_2494,N_2531);
nor U2609 (N_2609,N_2443,N_2504);
or U2610 (N_2610,N_2503,N_2425);
or U2611 (N_2611,N_2525,N_2438);
xor U2612 (N_2612,N_2442,N_2596);
nand U2613 (N_2613,N_2463,N_2579);
nor U2614 (N_2614,N_2441,N_2533);
or U2615 (N_2615,N_2514,N_2501);
nand U2616 (N_2616,N_2560,N_2588);
or U2617 (N_2617,N_2592,N_2496);
nor U2618 (N_2618,N_2446,N_2573);
and U2619 (N_2619,N_2551,N_2548);
or U2620 (N_2620,N_2591,N_2408);
and U2621 (N_2621,N_2465,N_2594);
or U2622 (N_2622,N_2475,N_2467);
nor U2623 (N_2623,N_2515,N_2405);
nor U2624 (N_2624,N_2497,N_2447);
and U2625 (N_2625,N_2528,N_2586);
nand U2626 (N_2626,N_2566,N_2431);
or U2627 (N_2627,N_2414,N_2485);
or U2628 (N_2628,N_2572,N_2453);
or U2629 (N_2629,N_2564,N_2534);
or U2630 (N_2630,N_2545,N_2415);
nand U2631 (N_2631,N_2519,N_2539);
or U2632 (N_2632,N_2430,N_2454);
or U2633 (N_2633,N_2409,N_2432);
nand U2634 (N_2634,N_2428,N_2412);
or U2635 (N_2635,N_2505,N_2543);
and U2636 (N_2636,N_2582,N_2434);
and U2637 (N_2637,N_2418,N_2520);
and U2638 (N_2638,N_2422,N_2490);
and U2639 (N_2639,N_2563,N_2555);
or U2640 (N_2640,N_2509,N_2502);
or U2641 (N_2641,N_2537,N_2487);
nand U2642 (N_2642,N_2550,N_2488);
nor U2643 (N_2643,N_2511,N_2424);
nand U2644 (N_2644,N_2440,N_2516);
nand U2645 (N_2645,N_2576,N_2419);
and U2646 (N_2646,N_2472,N_2557);
nor U2647 (N_2647,N_2544,N_2553);
or U2648 (N_2648,N_2420,N_2585);
or U2649 (N_2649,N_2464,N_2513);
nand U2650 (N_2650,N_2508,N_2577);
or U2651 (N_2651,N_2590,N_2493);
nor U2652 (N_2652,N_2416,N_2449);
nand U2653 (N_2653,N_2517,N_2506);
xnor U2654 (N_2654,N_2427,N_2451);
nor U2655 (N_2655,N_2522,N_2532);
nand U2656 (N_2656,N_2404,N_2565);
xor U2657 (N_2657,N_2421,N_2507);
or U2658 (N_2658,N_2547,N_2478);
or U2659 (N_2659,N_2561,N_2567);
nand U2660 (N_2660,N_2569,N_2587);
or U2661 (N_2661,N_2536,N_2558);
nand U2662 (N_2662,N_2574,N_2575);
nor U2663 (N_2663,N_2477,N_2562);
nor U2664 (N_2664,N_2476,N_2589);
or U2665 (N_2665,N_2486,N_2429);
xor U2666 (N_2666,N_2457,N_2406);
or U2667 (N_2667,N_2492,N_2530);
nor U2668 (N_2668,N_2417,N_2455);
nor U2669 (N_2669,N_2554,N_2482);
and U2670 (N_2670,N_2401,N_2578);
or U2671 (N_2671,N_2524,N_2439);
nand U2672 (N_2672,N_2426,N_2583);
or U2673 (N_2673,N_2448,N_2559);
nand U2674 (N_2674,N_2597,N_2527);
nand U2675 (N_2675,N_2580,N_2571);
or U2676 (N_2676,N_2479,N_2407);
or U2677 (N_2677,N_2459,N_2433);
nand U2678 (N_2678,N_2480,N_2444);
nor U2679 (N_2679,N_2450,N_2473);
nor U2680 (N_2680,N_2518,N_2435);
nand U2681 (N_2681,N_2510,N_2437);
or U2682 (N_2682,N_2458,N_2402);
nor U2683 (N_2683,N_2423,N_2499);
nand U2684 (N_2684,N_2541,N_2413);
nor U2685 (N_2685,N_2521,N_2452);
or U2686 (N_2686,N_2552,N_2599);
or U2687 (N_2687,N_2546,N_2535);
nand U2688 (N_2688,N_2593,N_2523);
nor U2689 (N_2689,N_2481,N_2491);
nand U2690 (N_2690,N_2460,N_2445);
or U2691 (N_2691,N_2474,N_2484);
xnor U2692 (N_2692,N_2468,N_2489);
nor U2693 (N_2693,N_2498,N_2581);
and U2694 (N_2694,N_2540,N_2538);
or U2695 (N_2695,N_2410,N_2466);
or U2696 (N_2696,N_2542,N_2436);
or U2697 (N_2697,N_2598,N_2461);
nor U2698 (N_2698,N_2568,N_2470);
or U2699 (N_2699,N_2403,N_2500);
nand U2700 (N_2700,N_2471,N_2504);
nor U2701 (N_2701,N_2430,N_2489);
nor U2702 (N_2702,N_2575,N_2453);
nor U2703 (N_2703,N_2444,N_2403);
or U2704 (N_2704,N_2447,N_2453);
and U2705 (N_2705,N_2509,N_2585);
nor U2706 (N_2706,N_2594,N_2409);
nor U2707 (N_2707,N_2521,N_2438);
nor U2708 (N_2708,N_2402,N_2502);
nor U2709 (N_2709,N_2560,N_2564);
nand U2710 (N_2710,N_2487,N_2597);
nand U2711 (N_2711,N_2463,N_2569);
and U2712 (N_2712,N_2580,N_2591);
nand U2713 (N_2713,N_2493,N_2412);
nor U2714 (N_2714,N_2517,N_2559);
nor U2715 (N_2715,N_2519,N_2557);
nor U2716 (N_2716,N_2545,N_2525);
or U2717 (N_2717,N_2518,N_2565);
nand U2718 (N_2718,N_2491,N_2579);
nor U2719 (N_2719,N_2549,N_2564);
nand U2720 (N_2720,N_2559,N_2502);
and U2721 (N_2721,N_2579,N_2416);
or U2722 (N_2722,N_2523,N_2506);
nor U2723 (N_2723,N_2476,N_2418);
or U2724 (N_2724,N_2513,N_2507);
nor U2725 (N_2725,N_2560,N_2468);
and U2726 (N_2726,N_2517,N_2592);
or U2727 (N_2727,N_2572,N_2596);
nor U2728 (N_2728,N_2539,N_2582);
nor U2729 (N_2729,N_2490,N_2518);
nand U2730 (N_2730,N_2464,N_2423);
nor U2731 (N_2731,N_2415,N_2578);
or U2732 (N_2732,N_2555,N_2474);
nor U2733 (N_2733,N_2477,N_2458);
or U2734 (N_2734,N_2559,N_2489);
or U2735 (N_2735,N_2450,N_2579);
or U2736 (N_2736,N_2536,N_2496);
nor U2737 (N_2737,N_2461,N_2439);
nand U2738 (N_2738,N_2569,N_2482);
nor U2739 (N_2739,N_2426,N_2560);
or U2740 (N_2740,N_2491,N_2439);
xor U2741 (N_2741,N_2566,N_2542);
nor U2742 (N_2742,N_2409,N_2477);
or U2743 (N_2743,N_2494,N_2516);
nand U2744 (N_2744,N_2467,N_2476);
or U2745 (N_2745,N_2596,N_2482);
nand U2746 (N_2746,N_2408,N_2490);
nor U2747 (N_2747,N_2539,N_2594);
nand U2748 (N_2748,N_2418,N_2448);
xor U2749 (N_2749,N_2502,N_2421);
nand U2750 (N_2750,N_2497,N_2545);
or U2751 (N_2751,N_2501,N_2542);
nor U2752 (N_2752,N_2441,N_2408);
nor U2753 (N_2753,N_2534,N_2546);
and U2754 (N_2754,N_2510,N_2449);
or U2755 (N_2755,N_2543,N_2570);
nand U2756 (N_2756,N_2531,N_2421);
xnor U2757 (N_2757,N_2504,N_2454);
nand U2758 (N_2758,N_2519,N_2490);
nor U2759 (N_2759,N_2494,N_2415);
or U2760 (N_2760,N_2436,N_2509);
nor U2761 (N_2761,N_2431,N_2458);
nand U2762 (N_2762,N_2511,N_2566);
or U2763 (N_2763,N_2529,N_2573);
or U2764 (N_2764,N_2540,N_2509);
and U2765 (N_2765,N_2519,N_2482);
and U2766 (N_2766,N_2441,N_2496);
or U2767 (N_2767,N_2588,N_2417);
nor U2768 (N_2768,N_2527,N_2532);
and U2769 (N_2769,N_2545,N_2496);
and U2770 (N_2770,N_2412,N_2489);
nor U2771 (N_2771,N_2489,N_2464);
and U2772 (N_2772,N_2476,N_2446);
nand U2773 (N_2773,N_2490,N_2557);
nand U2774 (N_2774,N_2429,N_2472);
nand U2775 (N_2775,N_2599,N_2412);
and U2776 (N_2776,N_2448,N_2446);
nor U2777 (N_2777,N_2501,N_2468);
xor U2778 (N_2778,N_2587,N_2537);
or U2779 (N_2779,N_2414,N_2505);
or U2780 (N_2780,N_2571,N_2431);
or U2781 (N_2781,N_2590,N_2463);
and U2782 (N_2782,N_2455,N_2595);
or U2783 (N_2783,N_2496,N_2482);
nand U2784 (N_2784,N_2421,N_2590);
nor U2785 (N_2785,N_2511,N_2557);
nand U2786 (N_2786,N_2517,N_2516);
nor U2787 (N_2787,N_2400,N_2490);
and U2788 (N_2788,N_2448,N_2508);
nand U2789 (N_2789,N_2598,N_2512);
nor U2790 (N_2790,N_2457,N_2507);
nor U2791 (N_2791,N_2466,N_2487);
nor U2792 (N_2792,N_2410,N_2476);
nand U2793 (N_2793,N_2458,N_2425);
nor U2794 (N_2794,N_2501,N_2515);
nand U2795 (N_2795,N_2476,N_2484);
nor U2796 (N_2796,N_2406,N_2581);
or U2797 (N_2797,N_2490,N_2437);
nor U2798 (N_2798,N_2529,N_2475);
nor U2799 (N_2799,N_2489,N_2562);
or U2800 (N_2800,N_2635,N_2753);
nand U2801 (N_2801,N_2778,N_2600);
and U2802 (N_2802,N_2792,N_2784);
and U2803 (N_2803,N_2739,N_2742);
or U2804 (N_2804,N_2685,N_2617);
or U2805 (N_2805,N_2692,N_2694);
nor U2806 (N_2806,N_2603,N_2726);
nand U2807 (N_2807,N_2632,N_2624);
and U2808 (N_2808,N_2609,N_2645);
and U2809 (N_2809,N_2670,N_2787);
nor U2810 (N_2810,N_2782,N_2691);
and U2811 (N_2811,N_2738,N_2623);
or U2812 (N_2812,N_2788,N_2662);
nand U2813 (N_2813,N_2730,N_2717);
nand U2814 (N_2814,N_2660,N_2735);
and U2815 (N_2815,N_2640,N_2672);
and U2816 (N_2816,N_2716,N_2751);
nand U2817 (N_2817,N_2729,N_2604);
nor U2818 (N_2818,N_2759,N_2736);
nor U2819 (N_2819,N_2762,N_2732);
and U2820 (N_2820,N_2601,N_2744);
or U2821 (N_2821,N_2765,N_2766);
nand U2822 (N_2822,N_2776,N_2728);
and U2823 (N_2823,N_2651,N_2612);
nor U2824 (N_2824,N_2674,N_2629);
or U2825 (N_2825,N_2763,N_2712);
and U2826 (N_2826,N_2610,N_2696);
and U2827 (N_2827,N_2731,N_2681);
nor U2828 (N_2828,N_2769,N_2661);
xor U2829 (N_2829,N_2602,N_2677);
and U2830 (N_2830,N_2680,N_2698);
nor U2831 (N_2831,N_2723,N_2678);
nand U2832 (N_2832,N_2658,N_2613);
and U2833 (N_2833,N_2709,N_2701);
nand U2834 (N_2834,N_2794,N_2684);
nand U2835 (N_2835,N_2772,N_2756);
nor U2836 (N_2836,N_2686,N_2725);
and U2837 (N_2837,N_2687,N_2654);
nand U2838 (N_2838,N_2614,N_2743);
and U2839 (N_2839,N_2775,N_2659);
nand U2840 (N_2840,N_2621,N_2644);
and U2841 (N_2841,N_2734,N_2630);
and U2842 (N_2842,N_2758,N_2703);
nor U2843 (N_2843,N_2707,N_2679);
or U2844 (N_2844,N_2646,N_2608);
and U2845 (N_2845,N_2795,N_2715);
and U2846 (N_2846,N_2675,N_2757);
or U2847 (N_2847,N_2767,N_2690);
or U2848 (N_2848,N_2746,N_2798);
or U2849 (N_2849,N_2627,N_2711);
nand U2850 (N_2850,N_2622,N_2702);
nand U2851 (N_2851,N_2611,N_2619);
nand U2852 (N_2852,N_2656,N_2755);
and U2853 (N_2853,N_2634,N_2704);
and U2854 (N_2854,N_2700,N_2633);
nor U2855 (N_2855,N_2683,N_2747);
and U2856 (N_2856,N_2790,N_2720);
or U2857 (N_2857,N_2628,N_2705);
and U2858 (N_2858,N_2770,N_2733);
nor U2859 (N_2859,N_2780,N_2721);
nand U2860 (N_2860,N_2647,N_2706);
nor U2861 (N_2861,N_2689,N_2641);
and U2862 (N_2862,N_2671,N_2649);
nand U2863 (N_2863,N_2760,N_2663);
nor U2864 (N_2864,N_2748,N_2796);
or U2865 (N_2865,N_2789,N_2718);
nor U2866 (N_2866,N_2676,N_2722);
nor U2867 (N_2867,N_2653,N_2666);
and U2868 (N_2868,N_2688,N_2797);
nor U2869 (N_2869,N_2699,N_2771);
nand U2870 (N_2870,N_2752,N_2638);
or U2871 (N_2871,N_2607,N_2618);
and U2872 (N_2872,N_2615,N_2749);
and U2873 (N_2873,N_2724,N_2673);
and U2874 (N_2874,N_2695,N_2719);
nor U2875 (N_2875,N_2791,N_2793);
or U2876 (N_2876,N_2657,N_2655);
nor U2877 (N_2877,N_2754,N_2697);
and U2878 (N_2878,N_2606,N_2708);
nand U2879 (N_2879,N_2779,N_2761);
nor U2880 (N_2880,N_2773,N_2652);
and U2881 (N_2881,N_2737,N_2665);
and U2882 (N_2882,N_2643,N_2750);
nor U2883 (N_2883,N_2777,N_2785);
nor U2884 (N_2884,N_2648,N_2714);
nand U2885 (N_2885,N_2625,N_2636);
or U2886 (N_2886,N_2745,N_2799);
nor U2887 (N_2887,N_2682,N_2667);
nor U2888 (N_2888,N_2740,N_2639);
and U2889 (N_2889,N_2637,N_2669);
or U2890 (N_2890,N_2764,N_2693);
and U2891 (N_2891,N_2616,N_2664);
nand U2892 (N_2892,N_2783,N_2786);
or U2893 (N_2893,N_2650,N_2626);
nor U2894 (N_2894,N_2668,N_2620);
or U2895 (N_2895,N_2642,N_2741);
nor U2896 (N_2896,N_2710,N_2774);
or U2897 (N_2897,N_2768,N_2713);
nand U2898 (N_2898,N_2781,N_2727);
or U2899 (N_2899,N_2631,N_2605);
nand U2900 (N_2900,N_2600,N_2627);
nand U2901 (N_2901,N_2776,N_2792);
or U2902 (N_2902,N_2629,N_2792);
or U2903 (N_2903,N_2680,N_2797);
or U2904 (N_2904,N_2718,N_2652);
and U2905 (N_2905,N_2770,N_2637);
nor U2906 (N_2906,N_2787,N_2606);
nand U2907 (N_2907,N_2614,N_2755);
nand U2908 (N_2908,N_2740,N_2667);
nand U2909 (N_2909,N_2687,N_2732);
nand U2910 (N_2910,N_2625,N_2780);
nand U2911 (N_2911,N_2605,N_2677);
or U2912 (N_2912,N_2680,N_2729);
nor U2913 (N_2913,N_2716,N_2785);
or U2914 (N_2914,N_2752,N_2703);
or U2915 (N_2915,N_2794,N_2660);
or U2916 (N_2916,N_2773,N_2711);
or U2917 (N_2917,N_2618,N_2648);
or U2918 (N_2918,N_2735,N_2624);
nor U2919 (N_2919,N_2744,N_2746);
nand U2920 (N_2920,N_2692,N_2795);
nor U2921 (N_2921,N_2784,N_2785);
nor U2922 (N_2922,N_2736,N_2677);
nand U2923 (N_2923,N_2768,N_2650);
nand U2924 (N_2924,N_2641,N_2781);
or U2925 (N_2925,N_2756,N_2642);
nand U2926 (N_2926,N_2727,N_2747);
and U2927 (N_2927,N_2650,N_2683);
nor U2928 (N_2928,N_2601,N_2731);
and U2929 (N_2929,N_2620,N_2762);
nor U2930 (N_2930,N_2696,N_2601);
and U2931 (N_2931,N_2749,N_2619);
nor U2932 (N_2932,N_2615,N_2798);
nand U2933 (N_2933,N_2667,N_2699);
or U2934 (N_2934,N_2649,N_2760);
nand U2935 (N_2935,N_2766,N_2629);
or U2936 (N_2936,N_2613,N_2790);
and U2937 (N_2937,N_2757,N_2753);
nor U2938 (N_2938,N_2667,N_2619);
nand U2939 (N_2939,N_2742,N_2653);
and U2940 (N_2940,N_2732,N_2609);
nor U2941 (N_2941,N_2779,N_2682);
or U2942 (N_2942,N_2781,N_2640);
nor U2943 (N_2943,N_2699,N_2657);
nand U2944 (N_2944,N_2660,N_2669);
or U2945 (N_2945,N_2635,N_2682);
and U2946 (N_2946,N_2628,N_2798);
or U2947 (N_2947,N_2613,N_2738);
and U2948 (N_2948,N_2790,N_2653);
and U2949 (N_2949,N_2768,N_2674);
nor U2950 (N_2950,N_2606,N_2734);
nand U2951 (N_2951,N_2709,N_2610);
nor U2952 (N_2952,N_2778,N_2760);
nand U2953 (N_2953,N_2671,N_2770);
or U2954 (N_2954,N_2641,N_2762);
nand U2955 (N_2955,N_2625,N_2708);
nand U2956 (N_2956,N_2766,N_2747);
nand U2957 (N_2957,N_2757,N_2761);
and U2958 (N_2958,N_2758,N_2604);
or U2959 (N_2959,N_2743,N_2671);
and U2960 (N_2960,N_2768,N_2766);
or U2961 (N_2961,N_2605,N_2796);
nand U2962 (N_2962,N_2773,N_2606);
and U2963 (N_2963,N_2713,N_2672);
or U2964 (N_2964,N_2753,N_2622);
and U2965 (N_2965,N_2757,N_2653);
nor U2966 (N_2966,N_2744,N_2689);
and U2967 (N_2967,N_2681,N_2625);
nand U2968 (N_2968,N_2760,N_2733);
or U2969 (N_2969,N_2750,N_2700);
and U2970 (N_2970,N_2625,N_2640);
or U2971 (N_2971,N_2638,N_2635);
and U2972 (N_2972,N_2707,N_2744);
nor U2973 (N_2973,N_2642,N_2656);
and U2974 (N_2974,N_2724,N_2623);
xor U2975 (N_2975,N_2676,N_2710);
and U2976 (N_2976,N_2603,N_2678);
nand U2977 (N_2977,N_2648,N_2696);
and U2978 (N_2978,N_2717,N_2736);
and U2979 (N_2979,N_2784,N_2668);
nor U2980 (N_2980,N_2760,N_2616);
nor U2981 (N_2981,N_2637,N_2699);
and U2982 (N_2982,N_2740,N_2615);
and U2983 (N_2983,N_2720,N_2649);
nand U2984 (N_2984,N_2715,N_2692);
and U2985 (N_2985,N_2668,N_2680);
nor U2986 (N_2986,N_2657,N_2611);
nor U2987 (N_2987,N_2755,N_2747);
or U2988 (N_2988,N_2743,N_2730);
and U2989 (N_2989,N_2760,N_2714);
nand U2990 (N_2990,N_2711,N_2601);
or U2991 (N_2991,N_2726,N_2750);
nor U2992 (N_2992,N_2679,N_2796);
nand U2993 (N_2993,N_2619,N_2655);
nand U2994 (N_2994,N_2723,N_2634);
or U2995 (N_2995,N_2653,N_2731);
nor U2996 (N_2996,N_2731,N_2667);
nor U2997 (N_2997,N_2774,N_2664);
nand U2998 (N_2998,N_2704,N_2738);
or U2999 (N_2999,N_2740,N_2715);
nor UO_0 (O_0,N_2832,N_2924);
or UO_1 (O_1,N_2979,N_2822);
nor UO_2 (O_2,N_2894,N_2930);
or UO_3 (O_3,N_2851,N_2810);
and UO_4 (O_4,N_2978,N_2986);
and UO_5 (O_5,N_2952,N_2813);
and UO_6 (O_6,N_2990,N_2836);
nand UO_7 (O_7,N_2937,N_2829);
and UO_8 (O_8,N_2866,N_2935);
or UO_9 (O_9,N_2834,N_2989);
nor UO_10 (O_10,N_2828,N_2971);
and UO_11 (O_11,N_2925,N_2812);
nand UO_12 (O_12,N_2948,N_2831);
nand UO_13 (O_13,N_2868,N_2840);
or UO_14 (O_14,N_2926,N_2929);
nand UO_15 (O_15,N_2886,N_2833);
and UO_16 (O_16,N_2872,N_2910);
nand UO_17 (O_17,N_2966,N_2975);
xnor UO_18 (O_18,N_2958,N_2950);
nor UO_19 (O_19,N_2913,N_2887);
or UO_20 (O_20,N_2988,N_2903);
nor UO_21 (O_21,N_2911,N_2964);
and UO_22 (O_22,N_2977,N_2854);
and UO_23 (O_23,N_2867,N_2998);
and UO_24 (O_24,N_2853,N_2839);
or UO_25 (O_25,N_2818,N_2876);
xnor UO_26 (O_26,N_2972,N_2819);
or UO_27 (O_27,N_2938,N_2820);
nor UO_28 (O_28,N_2920,N_2947);
or UO_29 (O_29,N_2904,N_2817);
and UO_30 (O_30,N_2804,N_2893);
nor UO_31 (O_31,N_2995,N_2803);
nand UO_32 (O_32,N_2885,N_2928);
and UO_33 (O_33,N_2870,N_2891);
or UO_34 (O_34,N_2888,N_2914);
nand UO_35 (O_35,N_2905,N_2902);
and UO_36 (O_36,N_2862,N_2835);
nor UO_37 (O_37,N_2823,N_2941);
nor UO_38 (O_38,N_2908,N_2883);
and UO_39 (O_39,N_2996,N_2847);
and UO_40 (O_40,N_2940,N_2841);
or UO_41 (O_41,N_2848,N_2884);
or UO_42 (O_42,N_2889,N_2955);
nand UO_43 (O_43,N_2982,N_2967);
and UO_44 (O_44,N_2997,N_2943);
or UO_45 (O_45,N_2849,N_2965);
nor UO_46 (O_46,N_2846,N_2949);
or UO_47 (O_47,N_2875,N_2946);
or UO_48 (O_48,N_2932,N_2918);
and UO_49 (O_49,N_2954,N_2973);
or UO_50 (O_50,N_2800,N_2827);
nor UO_51 (O_51,N_2980,N_2921);
nand UO_52 (O_52,N_2923,N_2882);
or UO_53 (O_53,N_2927,N_2900);
or UO_54 (O_54,N_2821,N_2805);
and UO_55 (O_55,N_2994,N_2806);
and UO_56 (O_56,N_2814,N_2944);
and UO_57 (O_57,N_2976,N_2916);
and UO_58 (O_58,N_2811,N_2871);
nand UO_59 (O_59,N_2991,N_2815);
nand UO_60 (O_60,N_2890,N_2942);
or UO_61 (O_61,N_2933,N_2951);
nor UO_62 (O_62,N_2808,N_2878);
nor UO_63 (O_63,N_2961,N_2983);
or UO_64 (O_64,N_2859,N_2824);
xor UO_65 (O_65,N_2917,N_2960);
and UO_66 (O_66,N_2934,N_2969);
and UO_67 (O_67,N_2957,N_2802);
and UO_68 (O_68,N_2864,N_2830);
and UO_69 (O_69,N_2974,N_2838);
or UO_70 (O_70,N_2993,N_2809);
nand UO_71 (O_71,N_2880,N_2919);
nand UO_72 (O_72,N_2992,N_2899);
nor UO_73 (O_73,N_2881,N_2843);
nor UO_74 (O_74,N_2865,N_2915);
and UO_75 (O_75,N_2936,N_2855);
and UO_76 (O_76,N_2963,N_2896);
nand UO_77 (O_77,N_2922,N_2906);
or UO_78 (O_78,N_2858,N_2897);
or UO_79 (O_79,N_2845,N_2844);
and UO_80 (O_80,N_2850,N_2912);
nor UO_81 (O_81,N_2863,N_2984);
nor UO_82 (O_82,N_2945,N_2895);
and UO_83 (O_83,N_2968,N_2852);
and UO_84 (O_84,N_2909,N_2962);
or UO_85 (O_85,N_2999,N_2939);
and UO_86 (O_86,N_2874,N_2879);
and UO_87 (O_87,N_2857,N_2807);
and UO_88 (O_88,N_2860,N_2892);
xnor UO_89 (O_89,N_2856,N_2907);
or UO_90 (O_90,N_2873,N_2837);
or UO_91 (O_91,N_2981,N_2959);
or UO_92 (O_92,N_2953,N_2826);
nand UO_93 (O_93,N_2816,N_2985);
nand UO_94 (O_94,N_2898,N_2931);
nand UO_95 (O_95,N_2877,N_2987);
nand UO_96 (O_96,N_2861,N_2825);
and UO_97 (O_97,N_2842,N_2901);
nor UO_98 (O_98,N_2801,N_2869);
nand UO_99 (O_99,N_2970,N_2956);
or UO_100 (O_100,N_2865,N_2972);
or UO_101 (O_101,N_2842,N_2808);
and UO_102 (O_102,N_2922,N_2862);
or UO_103 (O_103,N_2859,N_2802);
nor UO_104 (O_104,N_2914,N_2843);
or UO_105 (O_105,N_2815,N_2974);
nor UO_106 (O_106,N_2873,N_2911);
nor UO_107 (O_107,N_2868,N_2917);
nand UO_108 (O_108,N_2890,N_2918);
and UO_109 (O_109,N_2865,N_2885);
nand UO_110 (O_110,N_2914,N_2822);
or UO_111 (O_111,N_2954,N_2812);
nor UO_112 (O_112,N_2885,N_2849);
or UO_113 (O_113,N_2816,N_2881);
or UO_114 (O_114,N_2976,N_2947);
or UO_115 (O_115,N_2843,N_2938);
nand UO_116 (O_116,N_2984,N_2915);
or UO_117 (O_117,N_2943,N_2933);
nor UO_118 (O_118,N_2994,N_2817);
nand UO_119 (O_119,N_2872,N_2904);
nor UO_120 (O_120,N_2893,N_2928);
or UO_121 (O_121,N_2952,N_2928);
nand UO_122 (O_122,N_2829,N_2978);
or UO_123 (O_123,N_2902,N_2937);
nand UO_124 (O_124,N_2996,N_2851);
nor UO_125 (O_125,N_2866,N_2819);
nand UO_126 (O_126,N_2956,N_2957);
nor UO_127 (O_127,N_2881,N_2862);
or UO_128 (O_128,N_2922,N_2870);
nand UO_129 (O_129,N_2917,N_2851);
and UO_130 (O_130,N_2858,N_2904);
nor UO_131 (O_131,N_2940,N_2881);
or UO_132 (O_132,N_2929,N_2886);
nor UO_133 (O_133,N_2816,N_2906);
nand UO_134 (O_134,N_2950,N_2954);
nor UO_135 (O_135,N_2821,N_2817);
and UO_136 (O_136,N_2976,N_2807);
nor UO_137 (O_137,N_2849,N_2933);
nand UO_138 (O_138,N_2904,N_2823);
or UO_139 (O_139,N_2923,N_2835);
nand UO_140 (O_140,N_2957,N_2815);
nand UO_141 (O_141,N_2985,N_2948);
nor UO_142 (O_142,N_2992,N_2976);
nand UO_143 (O_143,N_2913,N_2830);
and UO_144 (O_144,N_2928,N_2880);
nor UO_145 (O_145,N_2848,N_2839);
nand UO_146 (O_146,N_2854,N_2824);
nand UO_147 (O_147,N_2927,N_2851);
or UO_148 (O_148,N_2809,N_2944);
or UO_149 (O_149,N_2934,N_2860);
or UO_150 (O_150,N_2902,N_2917);
or UO_151 (O_151,N_2843,N_2915);
or UO_152 (O_152,N_2858,N_2848);
and UO_153 (O_153,N_2838,N_2950);
nor UO_154 (O_154,N_2859,N_2990);
or UO_155 (O_155,N_2811,N_2927);
or UO_156 (O_156,N_2880,N_2960);
or UO_157 (O_157,N_2991,N_2877);
nor UO_158 (O_158,N_2860,N_2908);
or UO_159 (O_159,N_2857,N_2880);
or UO_160 (O_160,N_2818,N_2886);
nand UO_161 (O_161,N_2833,N_2867);
and UO_162 (O_162,N_2916,N_2914);
nor UO_163 (O_163,N_2944,N_2839);
nor UO_164 (O_164,N_2801,N_2841);
or UO_165 (O_165,N_2914,N_2973);
nor UO_166 (O_166,N_2912,N_2945);
xor UO_167 (O_167,N_2888,N_2927);
nor UO_168 (O_168,N_2872,N_2847);
nor UO_169 (O_169,N_2866,N_2884);
and UO_170 (O_170,N_2863,N_2958);
or UO_171 (O_171,N_2961,N_2996);
nand UO_172 (O_172,N_2978,N_2950);
or UO_173 (O_173,N_2969,N_2809);
or UO_174 (O_174,N_2892,N_2997);
nor UO_175 (O_175,N_2899,N_2815);
and UO_176 (O_176,N_2885,N_2974);
and UO_177 (O_177,N_2973,N_2807);
or UO_178 (O_178,N_2800,N_2802);
or UO_179 (O_179,N_2933,N_2821);
or UO_180 (O_180,N_2972,N_2934);
xnor UO_181 (O_181,N_2934,N_2839);
nor UO_182 (O_182,N_2884,N_2852);
or UO_183 (O_183,N_2970,N_2821);
and UO_184 (O_184,N_2894,N_2897);
nand UO_185 (O_185,N_2882,N_2877);
and UO_186 (O_186,N_2939,N_2954);
nand UO_187 (O_187,N_2959,N_2852);
xnor UO_188 (O_188,N_2802,N_2818);
or UO_189 (O_189,N_2893,N_2823);
and UO_190 (O_190,N_2997,N_2949);
or UO_191 (O_191,N_2994,N_2804);
nor UO_192 (O_192,N_2843,N_2800);
nand UO_193 (O_193,N_2871,N_2998);
or UO_194 (O_194,N_2924,N_2869);
nand UO_195 (O_195,N_2802,N_2833);
or UO_196 (O_196,N_2881,N_2807);
xnor UO_197 (O_197,N_2984,N_2816);
or UO_198 (O_198,N_2992,N_2844);
or UO_199 (O_199,N_2801,N_2978);
nor UO_200 (O_200,N_2923,N_2881);
nand UO_201 (O_201,N_2802,N_2881);
and UO_202 (O_202,N_2968,N_2919);
nand UO_203 (O_203,N_2809,N_2983);
and UO_204 (O_204,N_2845,N_2825);
nor UO_205 (O_205,N_2860,N_2910);
or UO_206 (O_206,N_2874,N_2969);
or UO_207 (O_207,N_2858,N_2923);
nor UO_208 (O_208,N_2930,N_2916);
nor UO_209 (O_209,N_2903,N_2933);
or UO_210 (O_210,N_2893,N_2841);
or UO_211 (O_211,N_2881,N_2951);
nand UO_212 (O_212,N_2997,N_2811);
nand UO_213 (O_213,N_2850,N_2932);
nor UO_214 (O_214,N_2972,N_2812);
nor UO_215 (O_215,N_2918,N_2814);
and UO_216 (O_216,N_2833,N_2964);
or UO_217 (O_217,N_2921,N_2805);
or UO_218 (O_218,N_2952,N_2925);
and UO_219 (O_219,N_2822,N_2952);
or UO_220 (O_220,N_2974,N_2850);
and UO_221 (O_221,N_2827,N_2801);
and UO_222 (O_222,N_2982,N_2910);
nand UO_223 (O_223,N_2915,N_2817);
and UO_224 (O_224,N_2846,N_2901);
or UO_225 (O_225,N_2923,N_2824);
or UO_226 (O_226,N_2946,N_2956);
nand UO_227 (O_227,N_2801,N_2837);
nor UO_228 (O_228,N_2864,N_2850);
nor UO_229 (O_229,N_2859,N_2907);
or UO_230 (O_230,N_2889,N_2931);
nor UO_231 (O_231,N_2971,N_2949);
and UO_232 (O_232,N_2889,N_2930);
nand UO_233 (O_233,N_2987,N_2989);
nor UO_234 (O_234,N_2955,N_2823);
or UO_235 (O_235,N_2986,N_2853);
and UO_236 (O_236,N_2975,N_2926);
nand UO_237 (O_237,N_2888,N_2958);
nor UO_238 (O_238,N_2989,N_2844);
or UO_239 (O_239,N_2818,N_2857);
nor UO_240 (O_240,N_2874,N_2904);
or UO_241 (O_241,N_2847,N_2963);
and UO_242 (O_242,N_2891,N_2854);
and UO_243 (O_243,N_2927,N_2889);
or UO_244 (O_244,N_2939,N_2827);
and UO_245 (O_245,N_2990,N_2963);
and UO_246 (O_246,N_2894,N_2946);
nor UO_247 (O_247,N_2877,N_2899);
nand UO_248 (O_248,N_2992,N_2846);
nor UO_249 (O_249,N_2888,N_2912);
and UO_250 (O_250,N_2818,N_2919);
nor UO_251 (O_251,N_2957,N_2999);
nand UO_252 (O_252,N_2999,N_2882);
nand UO_253 (O_253,N_2918,N_2870);
nand UO_254 (O_254,N_2957,N_2854);
or UO_255 (O_255,N_2810,N_2968);
or UO_256 (O_256,N_2930,N_2948);
nand UO_257 (O_257,N_2858,N_2993);
nand UO_258 (O_258,N_2864,N_2838);
and UO_259 (O_259,N_2975,N_2907);
nand UO_260 (O_260,N_2875,N_2867);
nor UO_261 (O_261,N_2857,N_2912);
nor UO_262 (O_262,N_2922,N_2953);
nand UO_263 (O_263,N_2829,N_2802);
nor UO_264 (O_264,N_2847,N_2874);
nand UO_265 (O_265,N_2809,N_2857);
and UO_266 (O_266,N_2941,N_2820);
nand UO_267 (O_267,N_2818,N_2825);
and UO_268 (O_268,N_2992,N_2923);
and UO_269 (O_269,N_2925,N_2941);
and UO_270 (O_270,N_2940,N_2809);
nand UO_271 (O_271,N_2965,N_2907);
nand UO_272 (O_272,N_2994,N_2920);
nor UO_273 (O_273,N_2816,N_2828);
or UO_274 (O_274,N_2987,N_2961);
nor UO_275 (O_275,N_2911,N_2956);
and UO_276 (O_276,N_2915,N_2881);
nor UO_277 (O_277,N_2908,N_2980);
nor UO_278 (O_278,N_2953,N_2918);
nor UO_279 (O_279,N_2873,N_2856);
and UO_280 (O_280,N_2880,N_2869);
nor UO_281 (O_281,N_2910,N_2818);
nand UO_282 (O_282,N_2862,N_2875);
and UO_283 (O_283,N_2935,N_2905);
nand UO_284 (O_284,N_2808,N_2832);
or UO_285 (O_285,N_2881,N_2933);
nor UO_286 (O_286,N_2831,N_2874);
and UO_287 (O_287,N_2806,N_2998);
and UO_288 (O_288,N_2976,N_2834);
and UO_289 (O_289,N_2977,N_2877);
or UO_290 (O_290,N_2806,N_2961);
nand UO_291 (O_291,N_2953,N_2856);
and UO_292 (O_292,N_2846,N_2933);
nand UO_293 (O_293,N_2805,N_2996);
or UO_294 (O_294,N_2881,N_2984);
or UO_295 (O_295,N_2890,N_2862);
and UO_296 (O_296,N_2892,N_2833);
nor UO_297 (O_297,N_2988,N_2855);
nand UO_298 (O_298,N_2998,N_2949);
or UO_299 (O_299,N_2947,N_2999);
and UO_300 (O_300,N_2996,N_2869);
or UO_301 (O_301,N_2824,N_2833);
nor UO_302 (O_302,N_2948,N_2887);
nor UO_303 (O_303,N_2811,N_2998);
and UO_304 (O_304,N_2838,N_2888);
nand UO_305 (O_305,N_2952,N_2823);
nand UO_306 (O_306,N_2902,N_2961);
nand UO_307 (O_307,N_2873,N_2914);
or UO_308 (O_308,N_2888,N_2977);
nand UO_309 (O_309,N_2990,N_2996);
or UO_310 (O_310,N_2966,N_2884);
nand UO_311 (O_311,N_2980,N_2880);
or UO_312 (O_312,N_2884,N_2947);
or UO_313 (O_313,N_2911,N_2994);
nor UO_314 (O_314,N_2982,N_2987);
and UO_315 (O_315,N_2865,N_2826);
nor UO_316 (O_316,N_2830,N_2916);
or UO_317 (O_317,N_2852,N_2920);
or UO_318 (O_318,N_2939,N_2981);
or UO_319 (O_319,N_2930,N_2897);
nor UO_320 (O_320,N_2867,N_2812);
nor UO_321 (O_321,N_2861,N_2801);
nor UO_322 (O_322,N_2813,N_2812);
nor UO_323 (O_323,N_2841,N_2883);
nor UO_324 (O_324,N_2863,N_2852);
and UO_325 (O_325,N_2895,N_2972);
or UO_326 (O_326,N_2817,N_2997);
or UO_327 (O_327,N_2968,N_2883);
or UO_328 (O_328,N_2848,N_2981);
nor UO_329 (O_329,N_2866,N_2834);
nand UO_330 (O_330,N_2876,N_2816);
nand UO_331 (O_331,N_2884,N_2833);
and UO_332 (O_332,N_2901,N_2942);
and UO_333 (O_333,N_2817,N_2917);
or UO_334 (O_334,N_2892,N_2981);
and UO_335 (O_335,N_2884,N_2942);
nand UO_336 (O_336,N_2801,N_2828);
nand UO_337 (O_337,N_2986,N_2884);
nand UO_338 (O_338,N_2891,N_2820);
nor UO_339 (O_339,N_2999,N_2986);
or UO_340 (O_340,N_2985,N_2895);
nor UO_341 (O_341,N_2830,N_2891);
nand UO_342 (O_342,N_2965,N_2824);
nor UO_343 (O_343,N_2968,N_2879);
nor UO_344 (O_344,N_2840,N_2941);
or UO_345 (O_345,N_2810,N_2834);
nand UO_346 (O_346,N_2997,N_2862);
nor UO_347 (O_347,N_2855,N_2847);
or UO_348 (O_348,N_2974,N_2968);
xor UO_349 (O_349,N_2898,N_2962);
xnor UO_350 (O_350,N_2821,N_2990);
nand UO_351 (O_351,N_2857,N_2866);
or UO_352 (O_352,N_2955,N_2975);
nor UO_353 (O_353,N_2978,N_2927);
nor UO_354 (O_354,N_2803,N_2993);
nor UO_355 (O_355,N_2979,N_2921);
or UO_356 (O_356,N_2897,N_2883);
nand UO_357 (O_357,N_2869,N_2949);
xor UO_358 (O_358,N_2995,N_2991);
nor UO_359 (O_359,N_2803,N_2806);
nand UO_360 (O_360,N_2811,N_2875);
or UO_361 (O_361,N_2940,N_2944);
or UO_362 (O_362,N_2895,N_2877);
nor UO_363 (O_363,N_2878,N_2952);
nor UO_364 (O_364,N_2995,N_2949);
nor UO_365 (O_365,N_2812,N_2825);
nor UO_366 (O_366,N_2943,N_2835);
nor UO_367 (O_367,N_2831,N_2955);
or UO_368 (O_368,N_2828,N_2872);
and UO_369 (O_369,N_2913,N_2818);
or UO_370 (O_370,N_2989,N_2821);
nor UO_371 (O_371,N_2983,N_2873);
nand UO_372 (O_372,N_2978,N_2918);
nand UO_373 (O_373,N_2977,N_2884);
nand UO_374 (O_374,N_2965,N_2927);
or UO_375 (O_375,N_2831,N_2873);
and UO_376 (O_376,N_2951,N_2853);
nand UO_377 (O_377,N_2928,N_2818);
and UO_378 (O_378,N_2987,N_2805);
nand UO_379 (O_379,N_2951,N_2994);
nor UO_380 (O_380,N_2969,N_2900);
or UO_381 (O_381,N_2940,N_2840);
nand UO_382 (O_382,N_2980,N_2962);
or UO_383 (O_383,N_2877,N_2859);
nor UO_384 (O_384,N_2984,N_2967);
nor UO_385 (O_385,N_2843,N_2922);
or UO_386 (O_386,N_2848,N_2905);
and UO_387 (O_387,N_2850,N_2976);
nand UO_388 (O_388,N_2846,N_2969);
and UO_389 (O_389,N_2873,N_2889);
nor UO_390 (O_390,N_2998,N_2923);
or UO_391 (O_391,N_2808,N_2915);
and UO_392 (O_392,N_2864,N_2940);
nand UO_393 (O_393,N_2959,N_2811);
and UO_394 (O_394,N_2923,N_2928);
and UO_395 (O_395,N_2924,N_2843);
or UO_396 (O_396,N_2969,N_2828);
nand UO_397 (O_397,N_2801,N_2918);
or UO_398 (O_398,N_2810,N_2887);
and UO_399 (O_399,N_2938,N_2924);
nor UO_400 (O_400,N_2914,N_2943);
nor UO_401 (O_401,N_2913,N_2915);
nand UO_402 (O_402,N_2970,N_2850);
and UO_403 (O_403,N_2974,N_2830);
nand UO_404 (O_404,N_2898,N_2963);
nor UO_405 (O_405,N_2808,N_2947);
and UO_406 (O_406,N_2997,N_2968);
nand UO_407 (O_407,N_2937,N_2813);
nor UO_408 (O_408,N_2870,N_2945);
nand UO_409 (O_409,N_2966,N_2878);
or UO_410 (O_410,N_2998,N_2839);
or UO_411 (O_411,N_2911,N_2849);
or UO_412 (O_412,N_2831,N_2848);
or UO_413 (O_413,N_2865,N_2833);
nand UO_414 (O_414,N_2982,N_2836);
nand UO_415 (O_415,N_2931,N_2922);
or UO_416 (O_416,N_2856,N_2906);
and UO_417 (O_417,N_2995,N_2951);
or UO_418 (O_418,N_2996,N_2952);
or UO_419 (O_419,N_2936,N_2912);
and UO_420 (O_420,N_2946,N_2992);
and UO_421 (O_421,N_2851,N_2893);
nand UO_422 (O_422,N_2948,N_2931);
nand UO_423 (O_423,N_2841,N_2947);
and UO_424 (O_424,N_2848,N_2947);
xor UO_425 (O_425,N_2854,N_2850);
nor UO_426 (O_426,N_2828,N_2808);
or UO_427 (O_427,N_2993,N_2863);
and UO_428 (O_428,N_2970,N_2963);
nand UO_429 (O_429,N_2854,N_2862);
or UO_430 (O_430,N_2896,N_2856);
and UO_431 (O_431,N_2970,N_2994);
or UO_432 (O_432,N_2938,N_2991);
and UO_433 (O_433,N_2932,N_2833);
or UO_434 (O_434,N_2840,N_2965);
nor UO_435 (O_435,N_2973,N_2857);
or UO_436 (O_436,N_2905,N_2895);
nand UO_437 (O_437,N_2890,N_2936);
nor UO_438 (O_438,N_2833,N_2845);
and UO_439 (O_439,N_2942,N_2866);
or UO_440 (O_440,N_2906,N_2874);
nor UO_441 (O_441,N_2989,N_2904);
nand UO_442 (O_442,N_2840,N_2919);
nand UO_443 (O_443,N_2817,N_2992);
xor UO_444 (O_444,N_2924,N_2814);
nand UO_445 (O_445,N_2966,N_2983);
nor UO_446 (O_446,N_2959,N_2889);
and UO_447 (O_447,N_2854,N_2881);
nand UO_448 (O_448,N_2938,N_2966);
nand UO_449 (O_449,N_2925,N_2855);
or UO_450 (O_450,N_2877,N_2842);
and UO_451 (O_451,N_2954,N_2800);
nand UO_452 (O_452,N_2817,N_2855);
nand UO_453 (O_453,N_2951,N_2993);
or UO_454 (O_454,N_2879,N_2960);
and UO_455 (O_455,N_2836,N_2857);
nand UO_456 (O_456,N_2962,N_2914);
or UO_457 (O_457,N_2850,N_2885);
and UO_458 (O_458,N_2988,N_2912);
nor UO_459 (O_459,N_2806,N_2809);
nor UO_460 (O_460,N_2839,N_2979);
nor UO_461 (O_461,N_2921,N_2981);
or UO_462 (O_462,N_2883,N_2873);
nor UO_463 (O_463,N_2813,N_2959);
nand UO_464 (O_464,N_2907,N_2920);
and UO_465 (O_465,N_2990,N_2993);
and UO_466 (O_466,N_2886,N_2876);
nor UO_467 (O_467,N_2954,N_2932);
or UO_468 (O_468,N_2823,N_2804);
nor UO_469 (O_469,N_2801,N_2885);
nor UO_470 (O_470,N_2814,N_2895);
nor UO_471 (O_471,N_2881,N_2886);
nor UO_472 (O_472,N_2890,N_2885);
and UO_473 (O_473,N_2933,N_2845);
or UO_474 (O_474,N_2906,N_2992);
nand UO_475 (O_475,N_2853,N_2929);
and UO_476 (O_476,N_2813,N_2899);
nand UO_477 (O_477,N_2918,N_2894);
and UO_478 (O_478,N_2930,N_2938);
or UO_479 (O_479,N_2837,N_2824);
and UO_480 (O_480,N_2812,N_2986);
nor UO_481 (O_481,N_2969,N_2842);
and UO_482 (O_482,N_2995,N_2875);
or UO_483 (O_483,N_2823,N_2894);
nor UO_484 (O_484,N_2825,N_2826);
nand UO_485 (O_485,N_2995,N_2976);
nor UO_486 (O_486,N_2802,N_2844);
and UO_487 (O_487,N_2858,N_2991);
and UO_488 (O_488,N_2801,N_2812);
and UO_489 (O_489,N_2904,N_2923);
nand UO_490 (O_490,N_2969,N_2889);
or UO_491 (O_491,N_2867,N_2972);
or UO_492 (O_492,N_2838,N_2980);
nand UO_493 (O_493,N_2982,N_2884);
and UO_494 (O_494,N_2955,N_2966);
nand UO_495 (O_495,N_2885,N_2956);
nand UO_496 (O_496,N_2950,N_2939);
or UO_497 (O_497,N_2942,N_2860);
nor UO_498 (O_498,N_2906,N_2847);
nor UO_499 (O_499,N_2992,N_2984);
endmodule