module basic_1500_15000_2000_50_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
and U0 (N_0,In_1383,In_62);
or U1 (N_1,In_584,In_378);
nand U2 (N_2,In_253,In_274);
nand U3 (N_3,In_638,In_314);
nand U4 (N_4,In_566,In_693);
nand U5 (N_5,In_731,In_417);
nor U6 (N_6,In_825,In_1237);
nor U7 (N_7,In_1281,In_1413);
nand U8 (N_8,In_17,In_1041);
and U9 (N_9,In_541,In_330);
or U10 (N_10,In_1066,In_1444);
and U11 (N_11,In_604,In_1007);
and U12 (N_12,In_1389,In_783);
and U13 (N_13,In_1165,In_1278);
xor U14 (N_14,In_1173,In_1141);
xnor U15 (N_15,In_726,In_1397);
nor U16 (N_16,In_876,In_997);
nor U17 (N_17,In_340,In_602);
or U18 (N_18,In_794,In_1283);
or U19 (N_19,In_152,In_1108);
nor U20 (N_20,In_925,In_847);
nor U21 (N_21,In_712,In_349);
xor U22 (N_22,In_1109,In_1057);
or U23 (N_23,In_20,In_108);
and U24 (N_24,In_213,In_494);
xor U25 (N_25,In_963,In_411);
xnor U26 (N_26,In_1097,In_1002);
nand U27 (N_27,In_236,In_905);
xnor U28 (N_28,In_127,In_579);
xnor U29 (N_29,In_697,In_316);
or U30 (N_30,In_1169,In_1287);
nand U31 (N_31,In_436,In_715);
or U32 (N_32,In_767,In_1220);
or U33 (N_33,In_772,In_1305);
and U34 (N_34,In_775,In_99);
nand U35 (N_35,In_728,In_1028);
or U36 (N_36,In_509,In_1496);
or U37 (N_37,In_1225,In_52);
nor U38 (N_38,In_35,In_974);
xor U39 (N_39,In_1341,In_359);
or U40 (N_40,In_81,In_1000);
nand U41 (N_41,In_448,In_771);
and U42 (N_42,In_678,In_55);
and U43 (N_43,In_1010,In_705);
and U44 (N_44,In_112,In_495);
and U45 (N_45,In_1029,In_1259);
nand U46 (N_46,In_839,In_600);
and U47 (N_47,In_1032,In_254);
or U48 (N_48,In_123,In_396);
and U49 (N_49,In_1103,In_118);
nor U50 (N_50,In_1150,In_1497);
or U51 (N_51,In_1133,In_734);
or U52 (N_52,In_1250,In_1113);
nor U53 (N_53,In_559,In_523);
or U54 (N_54,In_986,In_246);
and U55 (N_55,In_507,In_286);
xor U56 (N_56,In_1375,In_545);
or U57 (N_57,In_674,In_784);
nand U58 (N_58,In_1062,In_1298);
nand U59 (N_59,In_1263,In_603);
xnor U60 (N_60,In_700,In_1494);
or U61 (N_61,In_419,In_162);
and U62 (N_62,In_1132,In_40);
or U63 (N_63,In_1112,In_1477);
and U64 (N_64,In_337,In_363);
nand U65 (N_65,In_489,In_623);
nor U66 (N_66,In_570,In_1221);
xor U67 (N_67,In_1411,In_1234);
nor U68 (N_68,In_307,In_553);
nor U69 (N_69,In_93,In_513);
and U70 (N_70,In_1034,In_763);
xnor U71 (N_71,In_774,In_1364);
nand U72 (N_72,In_1125,In_61);
or U73 (N_73,In_104,In_1303);
xor U74 (N_74,In_131,In_1243);
or U75 (N_75,In_1058,In_1345);
or U76 (N_76,In_999,In_711);
nand U77 (N_77,In_1242,In_922);
nor U78 (N_78,In_423,In_251);
nor U79 (N_79,In_1377,In_450);
nor U80 (N_80,In_919,In_1363);
xor U81 (N_81,In_399,In_814);
and U82 (N_82,In_90,In_850);
and U83 (N_83,In_446,In_568);
nor U84 (N_84,In_585,In_1027);
or U85 (N_85,In_272,In_1333);
xnor U86 (N_86,In_439,In_231);
xor U87 (N_87,In_1198,In_1235);
or U88 (N_88,In_583,In_629);
or U89 (N_89,In_1154,In_689);
xnor U90 (N_90,In_696,In_838);
nand U91 (N_91,In_680,In_66);
nand U92 (N_92,In_287,In_822);
and U93 (N_93,In_199,In_373);
nor U94 (N_94,In_531,In_1460);
and U95 (N_95,In_658,In_407);
and U96 (N_96,In_950,In_1473);
or U97 (N_97,In_1446,In_572);
nand U98 (N_98,In_1428,In_854);
xor U99 (N_99,In_842,In_1139);
or U100 (N_100,In_1459,In_1328);
and U101 (N_101,In_483,In_857);
and U102 (N_102,In_485,In_292);
xor U103 (N_103,In_1137,In_1213);
nand U104 (N_104,In_145,In_518);
and U105 (N_105,In_683,In_719);
or U106 (N_106,In_270,In_377);
nor U107 (N_107,In_969,In_358);
nand U108 (N_108,In_1212,In_339);
nor U109 (N_109,In_1246,In_334);
or U110 (N_110,In_1081,In_170);
and U111 (N_111,In_1055,In_67);
nor U112 (N_112,In_621,In_74);
or U113 (N_113,In_470,In_1130);
and U114 (N_114,In_1370,In_453);
and U115 (N_115,In_46,In_57);
nor U116 (N_116,In_1270,In_125);
xor U117 (N_117,In_452,In_532);
and U118 (N_118,In_1189,In_1366);
nand U119 (N_119,In_150,In_322);
nand U120 (N_120,In_1082,In_889);
or U121 (N_121,In_1048,In_207);
and U122 (N_122,In_191,In_1174);
nor U123 (N_123,In_317,In_757);
and U124 (N_124,In_752,In_515);
and U125 (N_125,In_1493,In_1431);
nand U126 (N_126,In_174,In_329);
and U127 (N_127,In_652,In_987);
nand U128 (N_128,In_790,In_39);
nor U129 (N_129,In_1215,In_1261);
and U130 (N_130,In_724,In_973);
and U131 (N_131,In_1110,In_1443);
or U132 (N_132,In_806,In_1047);
xor U133 (N_133,In_302,In_321);
nand U134 (N_134,In_224,In_424);
nor U135 (N_135,In_43,In_480);
nand U136 (N_136,In_308,In_894);
nand U137 (N_137,In_832,In_1438);
nand U138 (N_138,In_122,In_1092);
nor U139 (N_139,In_1396,In_533);
nand U140 (N_140,In_467,In_409);
or U141 (N_141,In_617,In_1437);
xnor U142 (N_142,In_759,In_964);
nand U143 (N_143,In_63,In_5);
nor U144 (N_144,In_594,In_676);
nor U145 (N_145,In_812,In_1197);
xor U146 (N_146,In_1104,In_173);
and U147 (N_147,In_786,In_240);
nor U148 (N_148,In_156,In_427);
and U149 (N_149,In_718,In_1023);
or U150 (N_150,In_178,In_1005);
and U151 (N_151,In_1188,In_433);
nand U152 (N_152,In_1295,In_1052);
and U153 (N_153,In_1211,In_1316);
xnor U154 (N_154,In_606,In_547);
nand U155 (N_155,In_1408,In_114);
nand U156 (N_156,In_0,In_855);
or U157 (N_157,In_1071,In_295);
and U158 (N_158,In_1138,In_931);
nor U159 (N_159,In_918,In_745);
nor U160 (N_160,In_391,In_1084);
and U161 (N_161,In_1367,In_1284);
nand U162 (N_162,In_687,In_1180);
nand U163 (N_163,In_578,In_827);
and U164 (N_164,In_1120,In_761);
or U165 (N_165,In_1267,In_1335);
xor U166 (N_166,In_78,In_1471);
xor U167 (N_167,In_714,In_1244);
and U168 (N_168,In_1353,In_465);
and U169 (N_169,In_851,In_498);
xnor U170 (N_170,In_196,In_506);
nand U171 (N_171,In_1480,In_168);
and U172 (N_172,In_1076,In_1067);
xnor U173 (N_173,In_546,In_1483);
or U174 (N_174,In_462,In_1035);
xor U175 (N_175,In_810,In_672);
xor U176 (N_176,In_1166,In_900);
xnor U177 (N_177,In_1468,In_552);
xor U178 (N_178,In_344,In_1222);
nor U179 (N_179,In_628,In_482);
nand U180 (N_180,In_1190,In_1300);
and U181 (N_181,In_777,In_141);
xor U182 (N_182,In_1272,In_10);
or U183 (N_183,In_819,In_798);
and U184 (N_184,In_941,In_34);
and U185 (N_185,In_338,In_1230);
nand U186 (N_186,In_796,In_225);
xnor U187 (N_187,In_912,In_370);
or U188 (N_188,In_657,In_177);
and U189 (N_189,In_475,In_520);
and U190 (N_190,In_549,In_103);
xor U191 (N_191,In_536,In_1127);
nand U192 (N_192,In_204,In_1193);
xnor U193 (N_193,In_1122,In_468);
nor U194 (N_194,In_1085,In_497);
or U195 (N_195,In_356,In_743);
nor U196 (N_196,In_981,In_4);
xor U197 (N_197,In_312,In_51);
or U198 (N_198,In_1184,In_166);
xnor U199 (N_199,In_47,In_195);
and U200 (N_200,In_948,In_829);
xor U201 (N_201,In_284,In_400);
or U202 (N_202,In_245,In_631);
nor U203 (N_203,In_25,In_146);
or U204 (N_204,In_350,In_186);
and U205 (N_205,In_1365,In_930);
and U206 (N_206,In_1340,In_266);
xor U207 (N_207,In_1489,In_741);
xnor U208 (N_208,In_33,In_1465);
nor U209 (N_209,In_778,In_342);
xnor U210 (N_210,In_770,In_116);
nor U211 (N_211,In_1192,In_610);
nor U212 (N_212,In_362,In_1297);
and U213 (N_213,In_663,In_1275);
xor U214 (N_214,In_488,In_472);
nor U215 (N_215,In_12,In_1183);
nand U216 (N_216,In_867,In_1347);
or U217 (N_217,In_210,In_445);
and U218 (N_218,In_521,In_179);
and U219 (N_219,In_1388,In_1487);
nor U220 (N_220,In_1216,In_679);
xor U221 (N_221,In_31,In_1282);
xor U222 (N_222,In_815,In_319);
nor U223 (N_223,In_632,In_1121);
nor U224 (N_224,In_802,In_1181);
nand U225 (N_225,In_820,In_1256);
and U226 (N_226,In_1466,In_1185);
or U227 (N_227,In_1075,In_1485);
or U228 (N_228,In_526,In_230);
or U229 (N_229,In_435,In_985);
nor U230 (N_230,In_92,In_1436);
and U231 (N_231,In_525,In_296);
nor U232 (N_232,In_285,In_431);
and U233 (N_233,In_686,In_1355);
xor U234 (N_234,In_206,In_704);
xor U235 (N_235,In_1254,In_79);
and U236 (N_236,In_458,In_1306);
or U237 (N_237,In_682,In_897);
nor U238 (N_238,In_248,In_1145);
and U239 (N_239,In_325,In_1046);
xor U240 (N_240,In_664,In_1404);
nor U241 (N_241,In_165,In_404);
xnor U242 (N_242,In_535,In_333);
or U243 (N_243,In_1126,In_534);
xnor U244 (N_244,In_713,In_702);
or U245 (N_245,In_949,In_1315);
and U246 (N_246,In_343,In_639);
nor U247 (N_247,In_1382,In_590);
or U248 (N_248,In_1311,In_951);
nor U249 (N_249,In_164,In_76);
xnor U250 (N_250,In_128,In_216);
nand U251 (N_251,In_866,In_365);
nor U252 (N_252,In_68,In_1476);
xnor U253 (N_253,In_1146,In_1020);
or U254 (N_254,In_271,In_1031);
xor U255 (N_255,In_989,In_959);
xnor U256 (N_256,In_643,In_268);
or U257 (N_257,In_229,In_803);
and U258 (N_258,In_1412,In_1409);
nand U259 (N_259,In_1202,In_782);
xnor U260 (N_260,In_612,In_1495);
xor U261 (N_261,In_909,In_1239);
nor U262 (N_262,In_1218,In_1490);
nor U263 (N_263,In_1167,In_263);
and U264 (N_264,In_1274,In_920);
xnor U265 (N_265,In_273,In_269);
and U266 (N_266,In_1338,In_1271);
xnor U267 (N_267,In_364,In_878);
and U268 (N_268,In_110,In_1406);
and U269 (N_269,In_1417,In_281);
nor U270 (N_270,In_801,In_15);
and U271 (N_271,In_389,In_360);
or U272 (N_272,In_1260,In_1314);
and U273 (N_273,In_300,In_598);
or U274 (N_274,In_609,In_481);
nor U275 (N_275,In_1253,In_858);
or U276 (N_276,In_187,In_1499);
and U277 (N_277,In_887,In_1403);
or U278 (N_278,In_1276,In_935);
or U279 (N_279,In_383,In_161);
or U280 (N_280,In_1323,In_403);
xor U281 (N_281,In_587,In_1114);
and U282 (N_282,In_768,In_818);
nand U283 (N_283,In_556,In_1105);
or U284 (N_284,In_916,In_730);
nor U285 (N_285,In_841,In_554);
nor U286 (N_286,In_394,In_1474);
nor U287 (N_287,In_1107,In_27);
or U288 (N_288,In_201,In_218);
and U289 (N_289,In_1326,In_157);
or U290 (N_290,In_873,In_1098);
nand U291 (N_291,In_754,In_1458);
and U292 (N_292,In_1044,In_1163);
nand U293 (N_293,In_901,In_619);
nand U294 (N_294,In_82,In_1091);
and U295 (N_295,In_1042,In_352);
and U296 (N_296,In_297,In_1384);
or U297 (N_297,In_326,In_1293);
or U298 (N_298,In_1380,In_514);
nor U299 (N_299,In_660,In_926);
or U300 (N_300,N_224,N_214);
nand U301 (N_301,In_992,N_221);
or U302 (N_302,In_1013,In_659);
xnor U303 (N_303,In_1083,In_1290);
xnor U304 (N_304,In_903,In_557);
nor U305 (N_305,In_1117,In_1159);
xnor U306 (N_306,In_382,N_111);
or U307 (N_307,In_142,N_237);
nand U308 (N_308,N_293,In_1451);
and U309 (N_309,In_132,N_71);
xnor U310 (N_310,In_890,In_421);
xnor U311 (N_311,In_1461,N_90);
or U312 (N_312,N_119,In_978);
xnor U313 (N_313,N_278,In_461);
and U314 (N_314,In_567,In_1140);
nor U315 (N_315,N_117,In_908);
nand U316 (N_316,In_666,N_124);
or U317 (N_317,N_180,In_414);
and U318 (N_318,N_216,In_418);
or U319 (N_319,In_1414,In_137);
xnor U320 (N_320,In_23,N_290);
nor U321 (N_321,N_168,In_1080);
and U322 (N_322,N_175,In_217);
nand U323 (N_323,In_256,In_747);
nor U324 (N_324,In_871,N_115);
or U325 (N_325,N_140,In_739);
nor U326 (N_326,N_107,N_193);
and U327 (N_327,In_473,In_698);
and U328 (N_328,In_764,In_1424);
nor U329 (N_329,In_831,In_94);
xor U330 (N_330,In_1427,In_648);
nor U331 (N_331,In_654,N_63);
or U332 (N_332,In_1068,In_875);
and U333 (N_333,In_944,In_1472);
nor U334 (N_334,N_79,N_15);
nand U335 (N_335,In_222,N_80);
nor U336 (N_336,In_1312,In_924);
nand U337 (N_337,N_10,In_744);
nand U338 (N_338,In_571,In_869);
and U339 (N_339,In_906,In_670);
xnor U340 (N_340,In_1093,In_484);
xnor U341 (N_341,In_1177,In_940);
nor U342 (N_342,In_1207,In_740);
or U343 (N_343,In_324,In_107);
xor U344 (N_344,In_60,In_1350);
nor U345 (N_345,In_220,N_260);
nand U346 (N_346,In_991,In_490);
and U347 (N_347,In_21,In_1361);
or U348 (N_348,In_582,In_561);
or U349 (N_349,N_202,In_422);
or U350 (N_350,N_69,In_1462);
or U351 (N_351,In_1484,In_595);
xor U352 (N_352,In_392,N_41);
nand U353 (N_353,In_192,In_447);
nor U354 (N_354,In_907,N_160);
nor U355 (N_355,N_267,In_426);
nor U356 (N_356,In_402,In_1371);
and U357 (N_357,In_1131,In_574);
or U358 (N_358,In_834,In_977);
nor U359 (N_359,N_158,In_212);
nand U360 (N_360,In_1392,In_758);
and U361 (N_361,In_265,In_279);
nor U362 (N_362,In_884,In_932);
xnor U363 (N_363,In_1191,In_1401);
or U364 (N_364,In_811,In_160);
and U365 (N_365,In_486,In_1011);
xnor U366 (N_366,In_1024,In_98);
or U367 (N_367,N_33,In_956);
and U368 (N_368,In_725,In_1241);
nor U369 (N_369,N_13,N_211);
or U370 (N_370,N_252,In_859);
xor U371 (N_371,In_742,N_299);
and U372 (N_372,N_44,In_24);
or U373 (N_373,N_96,In_65);
or U374 (N_374,In_821,In_190);
or U375 (N_375,N_34,N_19);
nor U376 (N_376,In_258,In_1478);
xor U377 (N_377,N_207,In_48);
or U378 (N_378,In_1410,N_289);
nor U379 (N_379,In_381,In_892);
nor U380 (N_380,N_146,In_1224);
or U381 (N_381,In_881,In_1329);
and U382 (N_382,N_61,In_1425);
nor U383 (N_383,In_1030,In_1226);
nor U384 (N_384,In_115,In_1060);
nor U385 (N_385,N_222,In_252);
nor U386 (N_386,In_53,In_684);
nor U387 (N_387,In_1336,N_236);
or U388 (N_388,N_12,N_186);
xor U389 (N_389,In_70,N_257);
nor U390 (N_390,In_1343,In_1186);
xnor U391 (N_391,In_1026,N_94);
or U392 (N_392,N_39,In_91);
or U393 (N_393,N_192,In_618);
or U394 (N_394,N_151,In_727);
and U395 (N_395,In_1456,In_111);
nand U396 (N_396,In_885,In_299);
and U397 (N_397,In_184,In_477);
and U398 (N_398,In_1018,In_1320);
and U399 (N_399,In_649,In_524);
nor U400 (N_400,N_253,In_645);
nor U401 (N_401,In_625,In_675);
nand U402 (N_402,In_586,In_301);
or U403 (N_403,In_1349,N_109);
or U404 (N_404,In_1175,In_563);
nor U405 (N_405,In_277,N_273);
nor U406 (N_406,In_369,In_1398);
xnor U407 (N_407,In_936,N_228);
xor U408 (N_408,In_1432,N_25);
nand U409 (N_409,In_627,N_241);
nor U410 (N_410,In_817,In_1025);
and U411 (N_411,N_134,In_149);
or U412 (N_412,In_163,In_685);
nand U413 (N_413,In_406,In_544);
nor U414 (N_414,N_298,In_387);
or U415 (N_415,N_72,In_1142);
xor U416 (N_416,N_20,In_722);
and U417 (N_417,In_1168,In_332);
nor U418 (N_418,In_1294,N_37);
and U419 (N_419,In_1454,In_124);
or U420 (N_420,N_29,In_681);
xor U421 (N_421,In_1149,In_1072);
or U422 (N_422,In_888,In_310);
or U423 (N_423,In_345,In_1321);
and U424 (N_424,In_793,N_194);
nand U425 (N_425,In_3,In_1457);
nand U426 (N_426,In_694,In_813);
xnor U427 (N_427,In_278,N_159);
nor U428 (N_428,In_723,N_284);
or U429 (N_429,N_65,In_1433);
xnor U430 (N_430,In_393,In_1426);
nor U431 (N_431,In_868,In_182);
or U432 (N_432,In_189,In_255);
and U433 (N_433,In_139,In_237);
or U434 (N_434,N_116,N_36);
xnor U435 (N_435,In_7,N_254);
and U436 (N_436,In_1206,In_710);
and U437 (N_437,In_1160,In_1017);
xor U438 (N_438,In_1469,In_914);
and U439 (N_439,In_938,In_416);
nor U440 (N_440,In_1299,N_43);
xnor U441 (N_441,In_729,In_543);
nand U442 (N_442,N_70,In_856);
and U443 (N_443,In_1087,In_1399);
and U444 (N_444,In_996,In_6);
nor U445 (N_445,N_145,In_1325);
nor U446 (N_446,In_902,In_454);
nand U447 (N_447,In_998,In_1227);
xor U448 (N_448,In_955,In_1136);
or U449 (N_449,N_269,N_259);
and U450 (N_450,In_569,In_519);
and U451 (N_451,In_367,In_466);
xor U452 (N_452,N_0,In_347);
or U453 (N_453,In_836,N_181);
nor U454 (N_454,In_575,In_917);
or U455 (N_455,In_646,In_870);
and U456 (N_456,N_120,In_200);
nand U457 (N_457,N_282,N_68);
nand U458 (N_458,In_848,In_967);
nand U459 (N_459,N_67,In_947);
nand U460 (N_460,In_96,In_751);
and U461 (N_461,In_667,N_191);
or U462 (N_462,In_1178,N_195);
and U463 (N_463,In_1452,In_1036);
xor U464 (N_464,In_117,N_132);
and U465 (N_465,In_980,N_106);
xnor U466 (N_466,In_954,In_785);
nand U467 (N_467,In_573,N_239);
nor U468 (N_468,In_1106,N_66);
nand U469 (N_469,In_318,N_189);
xnor U470 (N_470,N_261,N_59);
nor U471 (N_471,In_510,In_637);
nand U472 (N_472,In_233,In_133);
xnor U473 (N_473,In_30,In_361);
xnor U474 (N_474,In_80,In_500);
xnor U475 (N_475,In_910,In_939);
xnor U476 (N_476,N_104,In_366);
nand U477 (N_477,N_234,In_564);
xnor U478 (N_478,In_214,In_443);
or U479 (N_479,N_22,N_38);
or U480 (N_480,In_241,N_210);
and U481 (N_481,In_833,In_376);
nand U482 (N_482,In_106,In_1481);
or U483 (N_483,N_139,In_580);
or U484 (N_484,In_749,N_64);
xnor U485 (N_485,In_1376,In_1147);
or U486 (N_486,N_58,N_198);
xnor U487 (N_487,In_290,In_708);
xnor U488 (N_488,In_807,In_1003);
xor U489 (N_489,In_677,In_1199);
xor U490 (N_490,In_1176,In_1236);
nor U491 (N_491,In_451,In_1077);
or U492 (N_492,In_493,N_242);
or U493 (N_493,In_323,In_756);
nand U494 (N_494,In_44,In_1279);
nand U495 (N_495,In_952,N_156);
xnor U496 (N_496,In_845,In_1289);
and U497 (N_497,N_102,N_1);
xor U498 (N_498,N_174,N_170);
nor U499 (N_499,N_206,In_1086);
xor U500 (N_500,In_1123,In_1187);
or U501 (N_501,In_1344,In_242);
or U502 (N_502,In_257,In_59);
nand U503 (N_503,In_799,In_504);
nor U504 (N_504,In_957,In_1196);
nand U505 (N_505,In_795,In_843);
and U506 (N_506,In_605,N_3);
nand U507 (N_507,In_895,In_1339);
or U508 (N_508,In_1088,In_1022);
nor U509 (N_509,In_1153,In_456);
nand U510 (N_510,In_805,In_375);
or U511 (N_511,In_1358,In_592);
xnor U512 (N_512,In_551,In_1449);
nor U513 (N_513,N_203,N_135);
and U514 (N_514,In_968,In_800);
or U515 (N_515,In_809,In_1357);
or U516 (N_516,In_1313,In_158);
nor U517 (N_517,In_85,In_1129);
or U518 (N_518,In_853,In_384);
or U519 (N_519,In_597,In_762);
nand U520 (N_520,In_701,In_471);
xor U521 (N_521,N_110,In_1247);
and U522 (N_522,N_274,In_984);
xnor U523 (N_523,In_650,In_966);
nor U524 (N_524,In_1492,In_765);
nor U525 (N_525,In_1151,In_613);
or U526 (N_526,In_1292,In_840);
nor U527 (N_527,In_501,N_131);
or U528 (N_528,In_596,In_1441);
xnor U529 (N_529,In_577,N_204);
nand U530 (N_530,In_1381,In_780);
nor U531 (N_531,In_642,In_865);
nor U532 (N_532,In_335,N_280);
or U533 (N_533,N_213,In_1001);
nand U534 (N_534,In_1208,In_915);
nand U535 (N_535,In_826,N_75);
nand U536 (N_536,N_275,N_57);
xnor U537 (N_537,In_508,In_1322);
and U538 (N_538,In_234,In_1447);
or U539 (N_539,In_934,In_662);
or U540 (N_540,N_232,In_1285);
xnor U541 (N_541,In_636,In_401);
or U542 (N_542,In_593,In_615);
nor U543 (N_543,N_138,N_114);
or U544 (N_544,In_291,In_1228);
nand U545 (N_545,N_126,In_1201);
and U546 (N_546,In_983,In_185);
nor U547 (N_547,In_692,In_1095);
or U548 (N_548,In_175,In_1245);
nand U549 (N_549,In_893,In_971);
nand U550 (N_550,In_1099,In_368);
and U551 (N_551,N_2,In_503);
and U552 (N_552,In_101,In_1407);
and U553 (N_553,In_1373,In_249);
nand U554 (N_554,In_669,N_287);
xor U555 (N_555,In_634,In_49);
xnor U556 (N_556,N_182,In_1400);
nand U557 (N_557,In_425,In_264);
xor U558 (N_558,In_1249,In_371);
nor U559 (N_559,In_429,In_1262);
nor U560 (N_560,In_144,In_315);
xnor U561 (N_561,In_589,In_8);
or U562 (N_562,N_54,N_153);
nand U563 (N_563,N_248,In_1498);
or U564 (N_564,N_223,In_83);
or U565 (N_565,N_296,N_103);
nor U566 (N_566,In_769,In_313);
and U567 (N_567,In_655,In_517);
nor U568 (N_568,In_641,N_6);
and U569 (N_569,In_1391,N_255);
nor U570 (N_570,In_1265,In_434);
and U571 (N_571,N_179,N_251);
and U572 (N_572,In_147,In_1049);
nor U573 (N_573,N_98,N_85);
nor U574 (N_574,N_281,In_988);
and U575 (N_575,N_208,N_74);
xnor U576 (N_576,In_886,N_276);
nand U577 (N_577,In_540,In_976);
nor U578 (N_578,In_937,N_133);
and U579 (N_579,N_185,In_267);
or U580 (N_580,In_1061,In_1051);
nor U581 (N_581,In_823,In_197);
nand U582 (N_582,In_496,N_28);
nor U583 (N_583,In_348,In_961);
nor U584 (N_584,In_1009,N_26);
xnor U585 (N_585,In_1378,In_537);
nor U586 (N_586,N_167,In_899);
or U587 (N_587,N_51,In_766);
xnor U588 (N_588,In_1394,In_331);
and U589 (N_589,In_933,In_760);
and U590 (N_590,N_82,In_644);
xor U591 (N_591,In_804,In_1359);
nor U592 (N_592,In_1124,In_491);
nor U593 (N_593,In_105,N_270);
xnor U594 (N_594,In_864,In_294);
nand U595 (N_595,In_1301,In_946);
and U596 (N_596,N_5,In_1337);
or U597 (N_597,N_112,In_2);
xor U598 (N_598,In_1453,In_154);
and U599 (N_599,In_235,In_211);
nor U600 (N_600,In_736,N_256);
or U601 (N_601,In_1450,N_559);
xnor U602 (N_602,N_231,N_402);
nand U603 (N_603,In_1308,In_1219);
nand U604 (N_604,N_442,N_328);
or U605 (N_605,N_488,In_1014);
and U606 (N_606,In_505,In_611);
nor U607 (N_607,N_78,N_31);
nor U608 (N_608,N_157,In_459);
xor U609 (N_609,In_432,In_1385);
nand U610 (N_610,In_183,In_395);
and U611 (N_611,In_262,In_1264);
nor U612 (N_612,N_149,N_121);
nand U613 (N_613,N_567,N_348);
or U614 (N_614,N_53,N_453);
or U615 (N_615,In_720,N_454);
nand U616 (N_616,N_365,N_499);
and U617 (N_617,N_339,N_574);
nor U618 (N_618,In_1334,In_420);
xor U619 (N_619,N_587,In_54);
and U620 (N_620,In_244,In_209);
and U621 (N_621,In_261,N_409);
or U622 (N_622,In_913,N_577);
xnor U623 (N_623,N_533,In_565);
nor U624 (N_624,In_1439,In_208);
nor U625 (N_625,In_354,N_524);
or U626 (N_626,In_408,N_105);
nand U627 (N_627,In_1442,In_703);
or U628 (N_628,In_695,In_219);
nor U629 (N_629,In_1346,N_432);
nand U630 (N_630,In_72,In_1162);
xnor U631 (N_631,N_262,In_1065);
nand U632 (N_632,N_143,N_319);
or U633 (N_633,N_285,N_586);
nand U634 (N_634,N_445,N_336);
and U635 (N_635,N_347,In_1054);
and U636 (N_636,N_32,N_42);
and U637 (N_637,In_1094,N_52);
xor U638 (N_638,In_153,In_1327);
or U639 (N_639,N_526,In_620);
or U640 (N_640,In_1229,N_383);
xnor U641 (N_641,N_505,In_1422);
nor U642 (N_642,In_750,In_1415);
xor U643 (N_643,In_1430,In_527);
nor U644 (N_644,N_434,In_22);
nor U645 (N_645,N_459,N_472);
nand U646 (N_646,N_521,N_363);
or U647 (N_647,N_486,In_591);
nor U648 (N_648,N_77,N_399);
xnor U649 (N_649,In_1379,N_7);
nand U650 (N_650,In_120,In_353);
nor U651 (N_651,N_447,In_1070);
nand U652 (N_652,N_422,In_753);
xnor U653 (N_653,In_1251,N_469);
nor U654 (N_654,N_50,N_502);
nor U655 (N_655,In_921,In_126);
nor U656 (N_656,N_349,N_455);
xor U657 (N_657,N_108,N_199);
nand U658 (N_658,N_327,In_1369);
and U659 (N_659,N_147,N_35);
nand U660 (N_660,N_529,In_633);
or U661 (N_661,N_345,N_288);
or U662 (N_662,In_460,N_27);
xor U663 (N_663,N_437,In_1164);
or U664 (N_664,N_342,N_583);
nand U665 (N_665,In_336,N_297);
nor U666 (N_666,In_327,N_405);
xor U667 (N_667,N_95,N_129);
and U668 (N_668,N_312,N_475);
nor U669 (N_669,In_1331,N_364);
nor U670 (N_670,In_71,In_437);
or U671 (N_671,In_119,In_1342);
nand U672 (N_672,In_882,N_142);
nor U673 (N_673,N_426,In_298);
and U674 (N_674,N_373,N_398);
and U675 (N_675,N_563,In_707);
and U676 (N_676,N_429,In_1362);
nor U677 (N_677,N_581,In_478);
xor U678 (N_678,N_118,N_400);
nand U679 (N_679,In_502,N_215);
nor U680 (N_680,In_1419,In_721);
xor U681 (N_681,In_476,In_651);
or U682 (N_682,N_391,In_1037);
xnor U683 (N_683,N_295,In_1064);
xor U684 (N_684,N_322,N_310);
or U685 (N_685,In_1310,In_883);
xnor U686 (N_686,In_1158,In_1296);
nor U687 (N_687,In_134,N_243);
and U688 (N_688,N_517,In_28);
nand U689 (N_689,N_161,In_1288);
nor U690 (N_690,N_238,N_263);
and U691 (N_691,In_1351,In_171);
nand U692 (N_692,N_561,N_233);
or U693 (N_693,N_317,N_47);
and U694 (N_694,In_283,N_318);
nor U695 (N_695,N_177,N_425);
nor U696 (N_696,N_380,N_320);
and U697 (N_697,N_585,In_306);
xnor U698 (N_698,In_138,N_440);
xnor U699 (N_699,N_197,In_42);
or U700 (N_700,In_440,In_1390);
or U701 (N_701,In_247,In_1491);
nor U702 (N_702,N_408,N_375);
xor U703 (N_703,In_788,N_21);
and U704 (N_704,In_282,N_362);
xor U705 (N_705,In_304,N_128);
nor U706 (N_706,In_781,N_438);
and U707 (N_707,N_531,N_576);
xnor U708 (N_708,In_844,In_1420);
or U709 (N_709,In_1118,N_393);
and U710 (N_710,In_1440,In_1038);
or U711 (N_711,N_18,In_1280);
nor U712 (N_712,N_356,N_492);
and U713 (N_713,N_394,In_69);
or U714 (N_714,N_592,In_309);
nor U715 (N_715,In_1209,In_159);
xnor U716 (N_716,N_172,In_1214);
and U717 (N_717,In_19,In_442);
or U718 (N_718,N_87,In_41);
xnor U719 (N_719,N_519,N_166);
and U720 (N_720,N_101,N_451);
nand U721 (N_721,In_194,N_389);
xnor U722 (N_722,In_1156,In_320);
nor U723 (N_723,N_331,N_565);
nand U724 (N_724,N_247,In_668);
xor U725 (N_725,In_614,N_360);
and U726 (N_726,N_99,N_562);
xor U727 (N_727,N_494,N_89);
nand U728 (N_728,N_523,N_335);
or U729 (N_729,N_176,N_127);
nor U730 (N_730,N_230,In_140);
and U731 (N_731,In_1238,In_188);
xor U732 (N_732,N_100,N_265);
xor U733 (N_733,In_415,In_1015);
nor U734 (N_734,N_582,In_990);
nand U735 (N_735,In_136,In_86);
nor U736 (N_736,N_300,N_546);
xor U737 (N_737,In_449,In_1317);
or U738 (N_738,N_554,In_243);
and U739 (N_739,N_379,In_576);
and U740 (N_740,In_1100,N_16);
nor U741 (N_741,In_1302,In_1356);
and U742 (N_742,N_11,In_1016);
xnor U743 (N_743,In_943,In_671);
or U744 (N_744,N_465,In_341);
nor U745 (N_745,N_534,In_202);
xor U746 (N_746,In_1332,N_184);
xor U747 (N_747,N_506,N_444);
xnor U748 (N_748,N_589,In_1006);
nand U749 (N_749,In_380,In_455);
nor U750 (N_750,N_307,N_346);
nor U751 (N_751,N_550,In_390);
or U752 (N_752,N_23,N_420);
nand U753 (N_753,In_193,In_75);
and U754 (N_754,N_370,N_309);
or U755 (N_755,In_1179,N_544);
nor U756 (N_756,N_476,In_1059);
xor U757 (N_757,In_1257,N_286);
or U758 (N_758,In_1152,N_359);
and U759 (N_759,N_512,N_569);
nor U760 (N_760,In_289,N_395);
and U761 (N_761,N_169,In_1423);
xor U762 (N_762,N_498,In_746);
and U763 (N_763,In_1008,In_463);
nor U764 (N_764,N_46,In_1);
or U765 (N_765,In_1056,In_1210);
or U766 (N_766,N_495,In_555);
xnor U767 (N_767,N_240,In_1387);
or U768 (N_768,In_1050,N_88);
and U769 (N_769,In_1360,In_239);
or U770 (N_770,In_167,N_547);
or U771 (N_771,N_17,N_418);
nand U772 (N_772,In_45,N_162);
xor U773 (N_773,In_1448,In_970);
nand U774 (N_774,In_787,N_479);
xnor U775 (N_775,In_647,In_1157);
or U776 (N_776,In_877,In_16);
nor U777 (N_777,In_1204,N_548);
nand U778 (N_778,In_1102,N_543);
nor U779 (N_779,N_514,In_102);
xor U780 (N_780,N_510,In_979);
and U781 (N_781,N_468,N_340);
and U782 (N_782,N_163,N_564);
nand U783 (N_783,N_480,In_1004);
and U784 (N_784,N_183,N_466);
nand U785 (N_785,N_386,N_478);
nand U786 (N_786,In_738,In_1101);
and U787 (N_787,N_62,In_962);
and U788 (N_788,N_150,N_188);
xor U789 (N_789,N_421,N_518);
or U790 (N_790,In_1161,N_406);
nand U791 (N_791,In_911,In_1319);
nor U792 (N_792,N_303,N_558);
or U793 (N_793,In_624,In_357);
nand U794 (N_794,N_598,N_441);
nand U795 (N_795,In_1435,In_1200);
or U796 (N_796,In_1324,N_381);
xor U797 (N_797,In_169,In_879);
nor U798 (N_798,N_93,In_1368);
or U799 (N_799,In_732,N_424);
nand U800 (N_800,N_477,N_246);
xor U801 (N_801,N_374,N_474);
nand U802 (N_802,N_430,N_575);
nand U803 (N_803,In_1240,In_374);
and U804 (N_804,In_232,N_24);
and U805 (N_805,N_200,In_151);
nor U806 (N_806,N_545,N_496);
nor U807 (N_807,In_64,N_450);
nor U808 (N_808,In_622,N_201);
xnor U809 (N_809,In_18,In_155);
nor U810 (N_810,N_413,In_1148);
nor U811 (N_811,N_377,N_357);
xor U812 (N_812,In_755,In_789);
and U813 (N_813,In_203,In_538);
and U814 (N_814,N_217,In_1488);
xor U815 (N_815,In_457,N_568);
or U816 (N_816,N_504,N_209);
or U817 (N_817,In_428,N_588);
nand U818 (N_818,In_487,In_953);
xnor U819 (N_819,In_923,In_172);
and U820 (N_820,N_404,N_154);
xor U821 (N_821,In_1255,N_334);
nor U822 (N_822,N_354,N_461);
nor U823 (N_823,N_458,N_448);
and U824 (N_824,In_898,N_411);
or U825 (N_825,N_258,N_361);
nand U826 (N_826,N_333,N_136);
nor U827 (N_827,N_489,N_81);
nor U828 (N_828,In_1395,In_305);
xor U829 (N_829,In_221,In_372);
nand U830 (N_830,N_225,In_1172);
and U831 (N_831,In_288,In_1039);
nand U832 (N_832,In_1135,In_260);
nor U833 (N_833,N_178,In_558);
nand U834 (N_834,In_1405,N_302);
or U835 (N_835,N_460,In_735);
and U836 (N_836,N_555,In_965);
xnor U837 (N_837,N_330,N_509);
and U838 (N_838,In_773,N_539);
xor U839 (N_839,In_846,In_982);
xnor U840 (N_840,N_56,In_479);
nor U841 (N_841,In_1203,N_137);
or U842 (N_842,N_196,In_1021);
or U843 (N_843,In_95,In_872);
or U844 (N_844,N_86,N_516);
nand U845 (N_845,In_1119,N_60);
nand U846 (N_846,In_776,In_1063);
or U847 (N_847,N_556,In_748);
nor U848 (N_848,In_13,In_1445);
or U849 (N_849,N_249,In_1352);
xor U850 (N_850,In_716,In_512);
xor U851 (N_851,In_492,N_387);
nand U852 (N_852,In_1273,In_1012);
or U853 (N_853,N_73,N_326);
xnor U854 (N_854,In_608,In_1053);
and U855 (N_855,In_1455,In_635);
xnor U856 (N_856,N_205,N_308);
xor U857 (N_857,In_205,In_665);
nor U858 (N_858,N_122,In_995);
nor U859 (N_859,N_272,In_276);
and U860 (N_860,N_491,In_530);
or U861 (N_861,In_346,In_958);
and U862 (N_862,In_97,In_88);
and U863 (N_863,N_532,N_599);
nand U864 (N_864,N_325,In_410);
and U865 (N_865,N_552,In_880);
nand U866 (N_866,In_38,N_452);
xnor U867 (N_867,N_511,In_528);
nand U868 (N_868,N_292,In_143);
nand U869 (N_869,N_549,N_113);
and U870 (N_870,In_1134,N_4);
or U871 (N_871,In_1182,In_1269);
or U872 (N_872,In_849,N_493);
nor U873 (N_873,In_1421,In_1479);
xor U874 (N_874,N_353,In_1043);
nand U875 (N_875,In_640,N_123);
nor U876 (N_876,In_994,In_874);
xor U877 (N_877,N_305,In_1416);
xnor U878 (N_878,N_219,In_397);
nand U879 (N_879,N_304,N_423);
nand U880 (N_880,In_89,N_462);
nand U881 (N_881,N_173,In_1143);
xnor U882 (N_882,In_542,In_180);
xor U883 (N_883,In_293,In_1019);
or U884 (N_884,In_1291,N_415);
nor U885 (N_885,N_431,In_1393);
and U886 (N_886,In_1286,In_1429);
and U887 (N_887,In_9,N_390);
xnor U888 (N_888,In_1223,N_8);
xor U889 (N_889,N_14,N_314);
nand U890 (N_890,In_808,In_1318);
nor U891 (N_891,N_435,N_40);
or U892 (N_892,In_11,In_1252);
or U893 (N_893,In_438,In_588);
and U894 (N_894,In_626,N_316);
nand U895 (N_895,In_835,N_385);
or U896 (N_896,N_218,N_584);
or U897 (N_897,In_1418,N_306);
nor U898 (N_898,In_942,In_1069);
nor U899 (N_899,In_109,In_355);
and U900 (N_900,N_893,N_828);
nand U901 (N_901,In_413,N_806);
nor U902 (N_902,N_605,N_323);
and U903 (N_903,N_679,In_50);
nand U904 (N_904,N_226,N_741);
xor U905 (N_905,In_699,N_485);
or U906 (N_906,In_599,N_700);
or U907 (N_907,In_37,In_860);
nor U908 (N_908,In_511,In_469);
nor U909 (N_909,N_652,N_714);
nor U910 (N_910,N_481,N_757);
nand U911 (N_911,N_865,N_672);
or U912 (N_912,N_751,N_542);
nor U913 (N_913,N_752,N_403);
nor U914 (N_914,N_351,In_1486);
xor U915 (N_915,N_484,In_779);
xnor U916 (N_916,N_781,In_228);
or U917 (N_917,N_845,N_753);
or U918 (N_918,N_626,N_321);
and U919 (N_919,N_407,N_730);
xnor U920 (N_920,N_874,N_775);
xnor U921 (N_921,N_637,N_849);
nor U922 (N_922,N_810,In_733);
nor U923 (N_923,N_647,N_683);
or U924 (N_924,N_834,N_392);
and U925 (N_925,N_693,N_449);
and U926 (N_926,N_710,N_780);
xor U927 (N_927,N_770,In_1195);
and U928 (N_928,N_746,N_83);
or U929 (N_929,In_1464,N_368);
xnor U930 (N_930,N_329,N_663);
nor U931 (N_931,N_732,In_690);
xor U932 (N_932,N_358,N_500);
or U933 (N_933,In_1374,N_571);
nor U934 (N_934,N_776,N_527);
and U935 (N_935,N_786,N_660);
and U936 (N_936,N_838,In_560);
xor U937 (N_937,N_875,In_379);
or U938 (N_938,N_867,N_635);
nor U939 (N_939,N_654,N_673);
nand U940 (N_940,N_621,N_763);
nor U941 (N_941,N_687,N_851);
xor U942 (N_942,N_725,In_1096);
nor U943 (N_943,In_36,N_646);
or U944 (N_944,N_439,In_58);
xor U945 (N_945,In_927,In_1233);
xnor U946 (N_946,N_600,N_528);
nor U947 (N_947,N_846,N_648);
or U948 (N_948,In_852,N_863);
and U949 (N_949,N_665,N_839);
xnor U950 (N_950,In_516,N_680);
or U951 (N_951,N_388,In_388);
nor U952 (N_952,N_737,In_1074);
or U953 (N_953,N_313,N_848);
or U954 (N_954,N_212,N_617);
nand U955 (N_955,In_1348,N_401);
or U956 (N_956,In_1217,N_742);
or U957 (N_957,N_551,N_827);
or U958 (N_958,N_844,N_9);
xnor U959 (N_959,N_877,N_688);
nand U960 (N_960,In_135,N_711);
nand U961 (N_961,In_176,N_410);
nand U962 (N_962,N_164,N_835);
and U963 (N_963,N_557,In_56);
and U964 (N_964,N_879,In_993);
xor U965 (N_965,N_376,N_804);
xor U966 (N_966,In_601,N_535);
xor U967 (N_967,In_223,N_756);
nor U968 (N_968,N_595,In_227);
nor U969 (N_969,N_782,N_91);
or U970 (N_970,N_774,N_823);
or U971 (N_971,N_525,N_634);
nor U972 (N_972,N_664,In_1078);
and U973 (N_973,N_803,In_385);
nor U974 (N_974,In_837,N_337);
nor U975 (N_975,N_490,N_832);
or U976 (N_976,N_817,N_613);
or U977 (N_977,N_866,N_704);
nor U978 (N_978,N_45,N_638);
and U979 (N_979,N_144,N_812);
xnor U980 (N_980,N_833,N_707);
nand U981 (N_981,N_669,N_792);
xor U982 (N_982,N_894,N_859);
xnor U983 (N_983,N_235,N_624);
nor U984 (N_984,In_26,N_887);
or U985 (N_985,N_895,In_1155);
nor U986 (N_986,In_328,In_673);
or U987 (N_987,N_630,In_661);
xnor U988 (N_988,N_315,N_734);
and U989 (N_989,N_743,N_890);
or U990 (N_990,N_716,N_606);
or U991 (N_991,In_928,In_1111);
xor U992 (N_992,In_691,N_779);
and U993 (N_993,N_662,In_100);
xnor U994 (N_994,In_1470,N_573);
or U995 (N_995,N_187,N_324);
nand U996 (N_996,N_837,N_815);
and U997 (N_997,N_591,In_1304);
nand U998 (N_998,In_441,In_1386);
and U999 (N_999,N_807,In_862);
and U1000 (N_1000,N_790,N_869);
xnor U1001 (N_1001,N_332,N_721);
nand U1002 (N_1002,N_596,N_857);
xnor U1003 (N_1003,N_777,N_513);
and U1004 (N_1004,N_854,N_609);
or U1005 (N_1005,N_748,In_828);
nand U1006 (N_1006,N_873,N_855);
nand U1007 (N_1007,N_897,In_1258);
xnor U1008 (N_1008,N_503,In_960);
xor U1009 (N_1009,N_783,N_892);
xnor U1010 (N_1010,N_229,N_698);
nor U1011 (N_1011,N_728,In_896);
xor U1012 (N_1012,In_130,In_303);
and U1013 (N_1013,In_1171,In_1040);
nand U1014 (N_1014,N_881,N_868);
and U1015 (N_1015,In_1232,N_764);
or U1016 (N_1016,N_870,In_522);
and U1017 (N_1017,N_771,N_642);
nor U1018 (N_1018,N_824,In_198);
or U1019 (N_1019,N_702,N_808);
nand U1020 (N_1020,N_655,N_729);
and U1021 (N_1021,N_853,N_607);
and U1022 (N_1022,N_722,N_457);
and U1023 (N_1023,In_474,In_215);
and U1024 (N_1024,In_398,In_706);
and U1025 (N_1025,N_378,N_668);
and U1026 (N_1026,N_816,N_141);
and U1027 (N_1027,N_850,In_891);
xor U1028 (N_1028,In_29,N_371);
and U1029 (N_1029,N_899,N_841);
nor U1030 (N_1030,N_541,N_836);
or U1031 (N_1031,N_819,In_975);
nand U1032 (N_1032,In_1170,N_520);
xnor U1033 (N_1033,N_482,In_972);
xor U1034 (N_1034,N_463,N_831);
and U1035 (N_1035,N_703,N_822);
or U1036 (N_1036,N_636,N_628);
nor U1037 (N_1037,N_311,In_1372);
nand U1038 (N_1038,N_657,In_1090);
and U1039 (N_1039,In_1463,N_656);
nand U1040 (N_1040,N_483,N_612);
and U1041 (N_1041,N_747,N_125);
xor U1042 (N_1042,N_653,N_355);
nor U1043 (N_1043,N_681,N_876);
or U1044 (N_1044,N_338,In_1089);
nor U1045 (N_1045,In_1079,N_697);
nor U1046 (N_1046,N_473,N_593);
and U1047 (N_1047,N_341,N_759);
and U1048 (N_1048,N_802,N_427);
nor U1049 (N_1049,N_758,In_1467);
nand U1050 (N_1050,In_121,N_676);
xnor U1051 (N_1051,N_553,N_889);
or U1052 (N_1052,N_366,N_797);
nand U1053 (N_1053,N_623,N_745);
xor U1054 (N_1054,N_661,N_884);
or U1055 (N_1055,N_659,N_794);
xor U1056 (N_1056,N_433,N_898);
or U1057 (N_1057,N_580,N_724);
and U1058 (N_1058,N_744,N_896);
and U1059 (N_1059,N_694,N_190);
nor U1060 (N_1060,In_1115,N_619);
or U1061 (N_1061,N_244,N_540);
xnor U1062 (N_1062,In_529,N_640);
nand U1063 (N_1063,N_871,N_464);
nand U1064 (N_1064,N_97,N_604);
or U1065 (N_1065,N_726,N_762);
or U1066 (N_1066,N_674,In_1194);
or U1067 (N_1067,In_386,N_736);
nor U1068 (N_1068,N_627,N_840);
or U1069 (N_1069,N_675,N_497);
nor U1070 (N_1070,N_615,N_291);
nor U1071 (N_1071,N_671,In_791);
and U1072 (N_1072,N_419,In_824);
nor U1073 (N_1073,In_830,N_620);
and U1074 (N_1074,N_727,In_539);
or U1075 (N_1075,N_508,In_1116);
nand U1076 (N_1076,N_755,N_861);
and U1077 (N_1077,N_670,N_611);
or U1078 (N_1078,In_709,In_607);
or U1079 (N_1079,N_712,N_883);
or U1080 (N_1080,N_152,N_891);
nand U1081 (N_1081,N_677,N_800);
and U1082 (N_1082,N_689,N_165);
and U1083 (N_1083,N_487,N_749);
and U1084 (N_1084,N_515,N_814);
xnor U1085 (N_1085,N_631,N_739);
or U1086 (N_1086,N_826,N_536);
or U1087 (N_1087,N_695,In_1231);
nor U1088 (N_1088,N_733,N_76);
nor U1089 (N_1089,N_862,N_436);
nor U1090 (N_1090,N_843,N_412);
and U1091 (N_1091,N_842,N_760);
and U1092 (N_1092,N_530,N_537);
and U1093 (N_1093,N_829,In_1434);
and U1094 (N_1094,N_650,N_414);
xnor U1095 (N_1095,N_872,N_788);
xor U1096 (N_1096,N_708,N_860);
and U1097 (N_1097,N_417,N_227);
xnor U1098 (N_1098,N_692,N_769);
xnor U1099 (N_1099,In_32,N_886);
or U1100 (N_1100,N_597,In_14);
and U1101 (N_1101,N_761,N_813);
xnor U1102 (N_1102,In_1402,In_259);
or U1103 (N_1103,N_685,N_632);
nor U1104 (N_1104,N_682,N_789);
or U1105 (N_1105,In_581,N_608);
nor U1106 (N_1106,N_245,N_384);
or U1107 (N_1107,N_507,In_226);
and U1108 (N_1108,N_878,N_590);
nor U1109 (N_1109,N_821,N_602);
and U1110 (N_1110,N_818,N_301);
and U1111 (N_1111,N_277,N_271);
nor U1112 (N_1112,N_641,In_1128);
xnor U1113 (N_1113,N_772,N_610);
or U1114 (N_1114,N_787,N_416);
nor U1115 (N_1115,In_797,N_856);
and U1116 (N_1116,N_678,In_238);
nor U1117 (N_1117,N_805,N_522);
nand U1118 (N_1118,In_129,N_649);
xnor U1119 (N_1119,N_778,In_405);
and U1120 (N_1120,In_861,N_268);
and U1121 (N_1121,In_1033,N_572);
nor U1122 (N_1122,N_731,N_344);
and U1123 (N_1123,N_717,N_171);
nor U1124 (N_1124,N_791,In_412);
xor U1125 (N_1125,N_690,In_792);
and U1126 (N_1126,N_443,N_382);
nand U1127 (N_1127,In_550,N_765);
nand U1128 (N_1128,N_718,N_754);
and U1129 (N_1129,In_904,N_811);
and U1130 (N_1130,N_148,N_735);
nand U1131 (N_1131,N_651,In_688);
nor U1132 (N_1132,N_643,In_929);
xnor U1133 (N_1133,N_705,In_1482);
or U1134 (N_1134,N_666,In_113);
nor U1135 (N_1135,In_1248,N_684);
and U1136 (N_1136,In_77,In_351);
nor U1137 (N_1137,N_250,N_396);
and U1138 (N_1138,In_816,In_444);
and U1139 (N_1139,N_428,N_691);
or U1140 (N_1140,In_1309,N_467);
or U1141 (N_1141,N_352,In_464);
nand U1142 (N_1142,In_148,N_773);
and U1143 (N_1143,N_30,N_603);
xnor U1144 (N_1144,N_616,In_311);
and U1145 (N_1145,N_852,N_709);
and U1146 (N_1146,N_49,N_130);
and U1147 (N_1147,N_538,N_501);
nor U1148 (N_1148,N_830,N_367);
and U1149 (N_1149,N_578,In_430);
nor U1150 (N_1150,N_801,In_1045);
or U1151 (N_1151,In_1268,N_84);
xor U1152 (N_1152,In_653,N_471);
nor U1153 (N_1153,N_614,In_280);
or U1154 (N_1154,N_796,N_456);
nor U1155 (N_1155,N_799,N_350);
nand U1156 (N_1156,In_1266,In_1277);
xnor U1157 (N_1157,N_369,N_784);
nand U1158 (N_1158,N_864,N_768);
nand U1159 (N_1159,In_1205,N_446);
nand U1160 (N_1160,N_888,N_795);
or U1161 (N_1161,In_1144,In_616);
nand U1162 (N_1162,In_656,N_715);
and U1163 (N_1163,N_155,In_737);
and U1164 (N_1164,N_639,N_294);
nand U1165 (N_1165,In_73,N_220);
nand U1166 (N_1166,In_562,N_809);
and U1167 (N_1167,In_499,In_84);
nor U1168 (N_1168,N_847,N_397);
nand U1169 (N_1169,N_645,In_863);
or U1170 (N_1170,N_793,In_717);
nand U1171 (N_1171,N_343,N_618);
nand U1172 (N_1172,N_283,N_723);
nand U1173 (N_1173,In_548,N_719);
or U1174 (N_1174,N_825,N_798);
nand U1175 (N_1175,N_767,N_785);
and U1176 (N_1176,N_766,In_1475);
xnor U1177 (N_1177,N_55,N_372);
nor U1178 (N_1178,In_87,N_880);
nand U1179 (N_1179,N_625,N_658);
xor U1180 (N_1180,In_630,N_622);
nor U1181 (N_1181,N_686,N_92);
or U1182 (N_1182,N_885,N_560);
or U1183 (N_1183,N_706,In_181);
nand U1184 (N_1184,N_570,In_275);
xnor U1185 (N_1185,N_266,In_1330);
xnor U1186 (N_1186,N_858,N_594);
and U1187 (N_1187,In_1073,N_701);
xnor U1188 (N_1188,N_264,In_1307);
xnor U1189 (N_1189,N_579,N_48);
xor U1190 (N_1190,N_740,N_667);
nor U1191 (N_1191,N_629,N_633);
nand U1192 (N_1192,In_250,N_699);
xnor U1193 (N_1193,N_601,N_644);
xnor U1194 (N_1194,N_696,N_566);
and U1195 (N_1195,N_882,N_820);
or U1196 (N_1196,In_1354,N_720);
xnor U1197 (N_1197,In_945,N_750);
xnor U1198 (N_1198,N_470,N_713);
xor U1199 (N_1199,N_738,N_279);
and U1200 (N_1200,N_1199,N_1060);
nand U1201 (N_1201,N_983,N_1140);
or U1202 (N_1202,N_996,N_966);
or U1203 (N_1203,N_1059,N_1083);
or U1204 (N_1204,N_1165,N_1058);
nor U1205 (N_1205,N_1158,N_1073);
nand U1206 (N_1206,N_1181,N_920);
nand U1207 (N_1207,N_980,N_1193);
or U1208 (N_1208,N_1101,N_1196);
nor U1209 (N_1209,N_1135,N_1157);
and U1210 (N_1210,N_1166,N_1098);
nor U1211 (N_1211,N_1141,N_1033);
xnor U1212 (N_1212,N_1048,N_937);
or U1213 (N_1213,N_1075,N_1085);
xnor U1214 (N_1214,N_1138,N_1168);
nand U1215 (N_1215,N_919,N_934);
and U1216 (N_1216,N_961,N_984);
nor U1217 (N_1217,N_1137,N_970);
nor U1218 (N_1218,N_924,N_985);
and U1219 (N_1219,N_1045,N_1142);
nor U1220 (N_1220,N_979,N_1162);
nand U1221 (N_1221,N_1034,N_1038);
nand U1222 (N_1222,N_1008,N_1072);
or U1223 (N_1223,N_935,N_910);
or U1224 (N_1224,N_1068,N_986);
or U1225 (N_1225,N_989,N_1029);
nor U1226 (N_1226,N_906,N_1129);
and U1227 (N_1227,N_1039,N_965);
or U1228 (N_1228,N_959,N_1103);
and U1229 (N_1229,N_1180,N_947);
and U1230 (N_1230,N_921,N_1081);
nor U1231 (N_1231,N_1118,N_929);
nor U1232 (N_1232,N_915,N_1169);
and U1233 (N_1233,N_1106,N_1100);
and U1234 (N_1234,N_1119,N_1025);
or U1235 (N_1235,N_954,N_990);
or U1236 (N_1236,N_1177,N_1107);
nand U1237 (N_1237,N_1050,N_1056);
nand U1238 (N_1238,N_963,N_1197);
xnor U1239 (N_1239,N_1104,N_1126);
and U1240 (N_1240,N_952,N_1128);
or U1241 (N_1241,N_1071,N_976);
xor U1242 (N_1242,N_987,N_1148);
and U1243 (N_1243,N_1080,N_943);
nand U1244 (N_1244,N_1067,N_930);
or U1245 (N_1245,N_1145,N_1091);
nand U1246 (N_1246,N_1120,N_997);
nor U1247 (N_1247,N_1020,N_1078);
nor U1248 (N_1248,N_1144,N_1095);
xnor U1249 (N_1249,N_1046,N_1190);
and U1250 (N_1250,N_1160,N_993);
xor U1251 (N_1251,N_1149,N_1174);
xor U1252 (N_1252,N_1179,N_1093);
nor U1253 (N_1253,N_956,N_1032);
nor U1254 (N_1254,N_1176,N_971);
nand U1255 (N_1255,N_1178,N_1003);
and U1256 (N_1256,N_1125,N_1043);
nand U1257 (N_1257,N_936,N_975);
and U1258 (N_1258,N_1163,N_1051);
and U1259 (N_1259,N_926,N_918);
xnor U1260 (N_1260,N_1031,N_1132);
and U1261 (N_1261,N_1055,N_1122);
xnor U1262 (N_1262,N_974,N_945);
or U1263 (N_1263,N_1156,N_969);
nand U1264 (N_1264,N_1005,N_904);
nand U1265 (N_1265,N_940,N_1155);
and U1266 (N_1266,N_1110,N_1198);
nand U1267 (N_1267,N_1184,N_1147);
nand U1268 (N_1268,N_1009,N_933);
or U1269 (N_1269,N_1172,N_1109);
nor U1270 (N_1270,N_1134,N_1052);
and U1271 (N_1271,N_953,N_1014);
xnor U1272 (N_1272,N_1066,N_1111);
nand U1273 (N_1273,N_1112,N_1099);
xor U1274 (N_1274,N_1164,N_922);
or U1275 (N_1275,N_962,N_1154);
and U1276 (N_1276,N_1006,N_1105);
nand U1277 (N_1277,N_1023,N_948);
or U1278 (N_1278,N_1139,N_1062);
xor U1279 (N_1279,N_958,N_1016);
nor U1280 (N_1280,N_1017,N_1108);
nor U1281 (N_1281,N_911,N_1047);
nand U1282 (N_1282,N_1030,N_1044);
nor U1283 (N_1283,N_1136,N_1012);
nor U1284 (N_1284,N_1040,N_1028);
and U1285 (N_1285,N_1127,N_1074);
or U1286 (N_1286,N_1121,N_1175);
xnor U1287 (N_1287,N_1013,N_992);
and U1288 (N_1288,N_916,N_967);
nor U1289 (N_1289,N_955,N_1057);
nor U1290 (N_1290,N_1082,N_1036);
nand U1291 (N_1291,N_1114,N_1084);
nand U1292 (N_1292,N_900,N_941);
and U1293 (N_1293,N_912,N_1173);
and U1294 (N_1294,N_1041,N_928);
xor U1295 (N_1295,N_902,N_1102);
nor U1296 (N_1296,N_1117,N_923);
nor U1297 (N_1297,N_1010,N_938);
and U1298 (N_1298,N_1061,N_973);
nor U1299 (N_1299,N_1194,N_1087);
nor U1300 (N_1300,N_1159,N_1079);
nand U1301 (N_1301,N_1187,N_1113);
nand U1302 (N_1302,N_1186,N_1185);
nand U1303 (N_1303,N_1130,N_995);
or U1304 (N_1304,N_1131,N_939);
and U1305 (N_1305,N_1022,N_944);
or U1306 (N_1306,N_972,N_908);
nor U1307 (N_1307,N_1092,N_1183);
nor U1308 (N_1308,N_994,N_1086);
xnor U1309 (N_1309,N_1011,N_1037);
xor U1310 (N_1310,N_1133,N_988);
nor U1311 (N_1311,N_1001,N_1123);
or U1312 (N_1312,N_1150,N_1143);
or U1313 (N_1313,N_1026,N_1096);
nand U1314 (N_1314,N_1182,N_1064);
and U1315 (N_1315,N_1054,N_991);
nand U1316 (N_1316,N_978,N_1189);
or U1317 (N_1317,N_1094,N_931);
and U1318 (N_1318,N_1153,N_1195);
nor U1319 (N_1319,N_946,N_982);
xor U1320 (N_1320,N_1090,N_932);
xor U1321 (N_1321,N_1049,N_1018);
and U1322 (N_1322,N_1146,N_1188);
xor U1323 (N_1323,N_1089,N_977);
nor U1324 (N_1324,N_1171,N_1007);
xor U1325 (N_1325,N_1024,N_950);
or U1326 (N_1326,N_1192,N_1076);
xnor U1327 (N_1327,N_1116,N_1167);
nor U1328 (N_1328,N_1151,N_949);
nor U1329 (N_1329,N_1035,N_1019);
xor U1330 (N_1330,N_1027,N_964);
xor U1331 (N_1331,N_1170,N_903);
nand U1332 (N_1332,N_1002,N_957);
and U1333 (N_1333,N_1015,N_917);
or U1334 (N_1334,N_1000,N_1042);
and U1335 (N_1335,N_1152,N_914);
nand U1336 (N_1336,N_1161,N_925);
or U1337 (N_1337,N_1004,N_1088);
and U1338 (N_1338,N_909,N_1053);
or U1339 (N_1339,N_968,N_998);
and U1340 (N_1340,N_1065,N_1115);
or U1341 (N_1341,N_907,N_1063);
or U1342 (N_1342,N_960,N_1191);
nand U1343 (N_1343,N_927,N_1124);
nor U1344 (N_1344,N_942,N_981);
nor U1345 (N_1345,N_1077,N_913);
xor U1346 (N_1346,N_1097,N_1021);
and U1347 (N_1347,N_951,N_1070);
nand U1348 (N_1348,N_1069,N_901);
or U1349 (N_1349,N_999,N_905);
xor U1350 (N_1350,N_900,N_1154);
or U1351 (N_1351,N_1081,N_997);
nor U1352 (N_1352,N_1171,N_927);
nand U1353 (N_1353,N_936,N_1057);
nor U1354 (N_1354,N_921,N_1022);
nand U1355 (N_1355,N_969,N_998);
and U1356 (N_1356,N_967,N_1078);
nand U1357 (N_1357,N_1147,N_1030);
nand U1358 (N_1358,N_1098,N_1084);
xnor U1359 (N_1359,N_946,N_942);
nor U1360 (N_1360,N_1068,N_923);
nand U1361 (N_1361,N_1033,N_973);
and U1362 (N_1362,N_919,N_986);
nand U1363 (N_1363,N_1122,N_1132);
or U1364 (N_1364,N_1154,N_926);
xnor U1365 (N_1365,N_909,N_1014);
and U1366 (N_1366,N_1162,N_963);
nor U1367 (N_1367,N_1079,N_935);
nor U1368 (N_1368,N_1060,N_995);
nor U1369 (N_1369,N_1053,N_1161);
and U1370 (N_1370,N_992,N_1036);
or U1371 (N_1371,N_912,N_922);
and U1372 (N_1372,N_1022,N_1099);
nor U1373 (N_1373,N_1066,N_1006);
nand U1374 (N_1374,N_1197,N_941);
or U1375 (N_1375,N_1122,N_1103);
xnor U1376 (N_1376,N_1092,N_918);
nand U1377 (N_1377,N_1064,N_1007);
nand U1378 (N_1378,N_1110,N_915);
nand U1379 (N_1379,N_1166,N_1103);
and U1380 (N_1380,N_998,N_922);
or U1381 (N_1381,N_1152,N_938);
xor U1382 (N_1382,N_939,N_1078);
xor U1383 (N_1383,N_1100,N_945);
xor U1384 (N_1384,N_931,N_916);
and U1385 (N_1385,N_964,N_1053);
nor U1386 (N_1386,N_920,N_1137);
or U1387 (N_1387,N_962,N_944);
nand U1388 (N_1388,N_1083,N_962);
nor U1389 (N_1389,N_959,N_1169);
and U1390 (N_1390,N_1176,N_1025);
nand U1391 (N_1391,N_988,N_1122);
and U1392 (N_1392,N_992,N_915);
and U1393 (N_1393,N_1009,N_1039);
xor U1394 (N_1394,N_961,N_1169);
nor U1395 (N_1395,N_923,N_1197);
and U1396 (N_1396,N_904,N_1181);
nand U1397 (N_1397,N_1083,N_901);
xnor U1398 (N_1398,N_951,N_1198);
and U1399 (N_1399,N_1146,N_1043);
or U1400 (N_1400,N_969,N_1017);
xnor U1401 (N_1401,N_1073,N_1023);
xnor U1402 (N_1402,N_1119,N_1121);
nand U1403 (N_1403,N_1183,N_912);
xnor U1404 (N_1404,N_1002,N_924);
nand U1405 (N_1405,N_997,N_943);
or U1406 (N_1406,N_1018,N_987);
or U1407 (N_1407,N_961,N_970);
xnor U1408 (N_1408,N_973,N_1194);
xor U1409 (N_1409,N_1032,N_1089);
or U1410 (N_1410,N_1021,N_1051);
or U1411 (N_1411,N_969,N_1033);
xnor U1412 (N_1412,N_1156,N_1108);
nor U1413 (N_1413,N_1113,N_1164);
and U1414 (N_1414,N_978,N_1112);
nor U1415 (N_1415,N_1057,N_966);
nand U1416 (N_1416,N_914,N_954);
or U1417 (N_1417,N_1004,N_1002);
and U1418 (N_1418,N_986,N_982);
and U1419 (N_1419,N_1186,N_1166);
or U1420 (N_1420,N_909,N_1021);
or U1421 (N_1421,N_1161,N_1188);
xnor U1422 (N_1422,N_944,N_1100);
nand U1423 (N_1423,N_1189,N_1038);
nor U1424 (N_1424,N_907,N_926);
or U1425 (N_1425,N_997,N_998);
and U1426 (N_1426,N_1078,N_1128);
and U1427 (N_1427,N_927,N_948);
nand U1428 (N_1428,N_900,N_1067);
nand U1429 (N_1429,N_917,N_1065);
or U1430 (N_1430,N_1091,N_1199);
and U1431 (N_1431,N_934,N_1147);
xor U1432 (N_1432,N_1048,N_1185);
or U1433 (N_1433,N_1022,N_1153);
xor U1434 (N_1434,N_1169,N_1029);
xnor U1435 (N_1435,N_1199,N_908);
xor U1436 (N_1436,N_946,N_1033);
and U1437 (N_1437,N_1182,N_1082);
nor U1438 (N_1438,N_1148,N_1040);
nand U1439 (N_1439,N_1175,N_925);
or U1440 (N_1440,N_1053,N_970);
xor U1441 (N_1441,N_1034,N_1178);
nand U1442 (N_1442,N_1047,N_1092);
and U1443 (N_1443,N_1082,N_1141);
nand U1444 (N_1444,N_1133,N_967);
nand U1445 (N_1445,N_1145,N_916);
nor U1446 (N_1446,N_1015,N_1059);
or U1447 (N_1447,N_982,N_992);
or U1448 (N_1448,N_1107,N_987);
nand U1449 (N_1449,N_1098,N_957);
nor U1450 (N_1450,N_925,N_942);
or U1451 (N_1451,N_1191,N_1032);
or U1452 (N_1452,N_1124,N_1011);
xnor U1453 (N_1453,N_1138,N_977);
nand U1454 (N_1454,N_1198,N_1114);
and U1455 (N_1455,N_1048,N_984);
nand U1456 (N_1456,N_966,N_920);
nand U1457 (N_1457,N_1089,N_990);
nor U1458 (N_1458,N_1000,N_1172);
nand U1459 (N_1459,N_1124,N_982);
nand U1460 (N_1460,N_1050,N_1020);
nor U1461 (N_1461,N_1065,N_1075);
nor U1462 (N_1462,N_955,N_1142);
or U1463 (N_1463,N_1088,N_1121);
or U1464 (N_1464,N_961,N_1197);
and U1465 (N_1465,N_1146,N_1126);
or U1466 (N_1466,N_1077,N_1149);
nor U1467 (N_1467,N_1053,N_1091);
and U1468 (N_1468,N_1110,N_911);
or U1469 (N_1469,N_928,N_1033);
nor U1470 (N_1470,N_1017,N_1121);
xor U1471 (N_1471,N_957,N_1049);
or U1472 (N_1472,N_945,N_1054);
nand U1473 (N_1473,N_927,N_1161);
nor U1474 (N_1474,N_967,N_938);
xnor U1475 (N_1475,N_921,N_935);
nor U1476 (N_1476,N_1021,N_1082);
nor U1477 (N_1477,N_1019,N_1006);
nand U1478 (N_1478,N_1138,N_1149);
nand U1479 (N_1479,N_983,N_1036);
xnor U1480 (N_1480,N_1098,N_979);
xnor U1481 (N_1481,N_942,N_1144);
nor U1482 (N_1482,N_1079,N_947);
nand U1483 (N_1483,N_950,N_1054);
or U1484 (N_1484,N_993,N_1154);
xnor U1485 (N_1485,N_1060,N_1094);
and U1486 (N_1486,N_1052,N_924);
nor U1487 (N_1487,N_1004,N_1073);
and U1488 (N_1488,N_1078,N_1188);
nand U1489 (N_1489,N_959,N_1022);
nand U1490 (N_1490,N_957,N_965);
nor U1491 (N_1491,N_1106,N_1142);
xor U1492 (N_1492,N_1087,N_1059);
or U1493 (N_1493,N_1102,N_1069);
or U1494 (N_1494,N_1158,N_906);
and U1495 (N_1495,N_957,N_1093);
xnor U1496 (N_1496,N_1159,N_1185);
xor U1497 (N_1497,N_993,N_1009);
nand U1498 (N_1498,N_1016,N_990);
or U1499 (N_1499,N_1162,N_1032);
nor U1500 (N_1500,N_1396,N_1421);
xor U1501 (N_1501,N_1432,N_1465);
or U1502 (N_1502,N_1361,N_1373);
nand U1503 (N_1503,N_1382,N_1410);
nor U1504 (N_1504,N_1428,N_1457);
nand U1505 (N_1505,N_1366,N_1328);
xnor U1506 (N_1506,N_1468,N_1487);
nor U1507 (N_1507,N_1417,N_1242);
nor U1508 (N_1508,N_1284,N_1354);
and U1509 (N_1509,N_1339,N_1258);
nand U1510 (N_1510,N_1244,N_1498);
xor U1511 (N_1511,N_1293,N_1255);
nand U1512 (N_1512,N_1494,N_1357);
and U1513 (N_1513,N_1451,N_1402);
nand U1514 (N_1514,N_1492,N_1379);
nor U1515 (N_1515,N_1345,N_1299);
xnor U1516 (N_1516,N_1356,N_1360);
or U1517 (N_1517,N_1227,N_1460);
xor U1518 (N_1518,N_1349,N_1476);
xor U1519 (N_1519,N_1479,N_1423);
nor U1520 (N_1520,N_1403,N_1438);
nand U1521 (N_1521,N_1369,N_1298);
nand U1522 (N_1522,N_1474,N_1208);
and U1523 (N_1523,N_1325,N_1201);
or U1524 (N_1524,N_1367,N_1384);
or U1525 (N_1525,N_1297,N_1320);
xnor U1526 (N_1526,N_1401,N_1383);
nand U1527 (N_1527,N_1287,N_1407);
nand U1528 (N_1528,N_1425,N_1265);
or U1529 (N_1529,N_1362,N_1351);
xor U1530 (N_1530,N_1217,N_1453);
nand U1531 (N_1531,N_1427,N_1279);
xnor U1532 (N_1532,N_1283,N_1415);
and U1533 (N_1533,N_1497,N_1480);
or U1534 (N_1534,N_1323,N_1378);
and U1535 (N_1535,N_1355,N_1385);
or U1536 (N_1536,N_1414,N_1314);
xor U1537 (N_1537,N_1470,N_1332);
xor U1538 (N_1538,N_1335,N_1266);
or U1539 (N_1539,N_1271,N_1285);
nand U1540 (N_1540,N_1368,N_1202);
xnor U1541 (N_1541,N_1463,N_1338);
xor U1542 (N_1542,N_1426,N_1329);
or U1543 (N_1543,N_1459,N_1397);
nand U1544 (N_1544,N_1377,N_1203);
nor U1545 (N_1545,N_1495,N_1493);
or U1546 (N_1546,N_1386,N_1376);
nand U1547 (N_1547,N_1394,N_1481);
and U1548 (N_1548,N_1239,N_1257);
nor U1549 (N_1549,N_1380,N_1461);
nand U1550 (N_1550,N_1234,N_1443);
and U1551 (N_1551,N_1301,N_1393);
nand U1552 (N_1552,N_1340,N_1353);
nand U1553 (N_1553,N_1315,N_1365);
xor U1554 (N_1554,N_1422,N_1250);
and U1555 (N_1555,N_1350,N_1464);
nor U1556 (N_1556,N_1249,N_1218);
or U1557 (N_1557,N_1486,N_1359);
nor U1558 (N_1558,N_1441,N_1260);
nor U1559 (N_1559,N_1295,N_1209);
and U1560 (N_1560,N_1324,N_1482);
xor U1561 (N_1561,N_1232,N_1433);
nor U1562 (N_1562,N_1216,N_1289);
nor U1563 (N_1563,N_1471,N_1302);
or U1564 (N_1564,N_1446,N_1319);
nor U1565 (N_1565,N_1313,N_1404);
and U1566 (N_1566,N_1306,N_1304);
xor U1567 (N_1567,N_1445,N_1455);
xor U1568 (N_1568,N_1224,N_1262);
xor U1569 (N_1569,N_1381,N_1326);
xor U1570 (N_1570,N_1400,N_1429);
nand U1571 (N_1571,N_1375,N_1267);
xor U1572 (N_1572,N_1264,N_1363);
xor U1573 (N_1573,N_1277,N_1496);
nand U1574 (N_1574,N_1406,N_1372);
nor U1575 (N_1575,N_1200,N_1300);
and U1576 (N_1576,N_1269,N_1473);
and U1577 (N_1577,N_1392,N_1488);
nor U1578 (N_1578,N_1472,N_1256);
or U1579 (N_1579,N_1499,N_1272);
nand U1580 (N_1580,N_1276,N_1305);
nor U1581 (N_1581,N_1437,N_1466);
and U1582 (N_1582,N_1390,N_1282);
and U1583 (N_1583,N_1204,N_1412);
xnor U1584 (N_1584,N_1225,N_1247);
nand U1585 (N_1585,N_1251,N_1228);
nor U1586 (N_1586,N_1248,N_1222);
nand U1587 (N_1587,N_1374,N_1364);
nor U1588 (N_1588,N_1442,N_1337);
or U1589 (N_1589,N_1274,N_1205);
xor U1590 (N_1590,N_1278,N_1254);
and U1591 (N_1591,N_1398,N_1409);
nor U1592 (N_1592,N_1296,N_1292);
nor U1593 (N_1593,N_1456,N_1483);
xor U1594 (N_1594,N_1237,N_1344);
nand U1595 (N_1595,N_1316,N_1341);
and U1596 (N_1596,N_1334,N_1405);
nor U1597 (N_1597,N_1230,N_1408);
nand U1598 (N_1598,N_1221,N_1245);
xor U1599 (N_1599,N_1310,N_1318);
and U1600 (N_1600,N_1347,N_1358);
nand U1601 (N_1601,N_1210,N_1321);
nor U1602 (N_1602,N_1458,N_1240);
nand U1603 (N_1603,N_1327,N_1447);
or U1604 (N_1604,N_1462,N_1434);
or U1605 (N_1605,N_1387,N_1330);
or U1606 (N_1606,N_1490,N_1223);
xor U1607 (N_1607,N_1439,N_1233);
or U1608 (N_1608,N_1211,N_1317);
or U1609 (N_1609,N_1273,N_1261);
or U1610 (N_1610,N_1238,N_1475);
nand U1611 (N_1611,N_1389,N_1342);
or U1612 (N_1612,N_1370,N_1491);
and U1613 (N_1613,N_1419,N_1207);
and U1614 (N_1614,N_1399,N_1435);
nand U1615 (N_1615,N_1308,N_1450);
or U1616 (N_1616,N_1280,N_1212);
and U1617 (N_1617,N_1235,N_1275);
or U1618 (N_1618,N_1252,N_1449);
or U1619 (N_1619,N_1303,N_1219);
nor U1620 (N_1620,N_1452,N_1418);
nand U1621 (N_1621,N_1268,N_1294);
nor U1622 (N_1622,N_1286,N_1241);
xor U1623 (N_1623,N_1454,N_1484);
nand U1624 (N_1624,N_1290,N_1288);
xor U1625 (N_1625,N_1312,N_1214);
or U1626 (N_1626,N_1246,N_1231);
nand U1627 (N_1627,N_1206,N_1352);
nand U1628 (N_1628,N_1395,N_1477);
nor U1629 (N_1629,N_1411,N_1469);
nor U1630 (N_1630,N_1431,N_1413);
nand U1631 (N_1631,N_1436,N_1348);
nor U1632 (N_1632,N_1263,N_1226);
xnor U1633 (N_1633,N_1467,N_1430);
nand U1634 (N_1634,N_1281,N_1388);
or U1635 (N_1635,N_1259,N_1343);
nor U1636 (N_1636,N_1448,N_1420);
nand U1637 (N_1637,N_1371,N_1322);
nor U1638 (N_1638,N_1416,N_1391);
or U1639 (N_1639,N_1270,N_1311);
nand U1640 (N_1640,N_1309,N_1331);
nand U1641 (N_1641,N_1243,N_1440);
nor U1642 (N_1642,N_1229,N_1485);
nor U1643 (N_1643,N_1424,N_1336);
xor U1644 (N_1644,N_1220,N_1333);
nor U1645 (N_1645,N_1291,N_1307);
or U1646 (N_1646,N_1213,N_1236);
and U1647 (N_1647,N_1444,N_1489);
nand U1648 (N_1648,N_1253,N_1478);
and U1649 (N_1649,N_1346,N_1215);
nor U1650 (N_1650,N_1294,N_1412);
nand U1651 (N_1651,N_1357,N_1200);
and U1652 (N_1652,N_1373,N_1452);
nand U1653 (N_1653,N_1461,N_1320);
nor U1654 (N_1654,N_1314,N_1449);
nor U1655 (N_1655,N_1303,N_1304);
and U1656 (N_1656,N_1322,N_1367);
xor U1657 (N_1657,N_1345,N_1461);
or U1658 (N_1658,N_1423,N_1287);
nor U1659 (N_1659,N_1494,N_1200);
nand U1660 (N_1660,N_1211,N_1302);
or U1661 (N_1661,N_1493,N_1444);
and U1662 (N_1662,N_1363,N_1270);
nor U1663 (N_1663,N_1246,N_1335);
nor U1664 (N_1664,N_1266,N_1303);
and U1665 (N_1665,N_1488,N_1290);
xnor U1666 (N_1666,N_1436,N_1329);
or U1667 (N_1667,N_1358,N_1247);
xnor U1668 (N_1668,N_1252,N_1282);
nor U1669 (N_1669,N_1264,N_1202);
or U1670 (N_1670,N_1270,N_1428);
and U1671 (N_1671,N_1335,N_1494);
nor U1672 (N_1672,N_1232,N_1227);
and U1673 (N_1673,N_1431,N_1289);
xnor U1674 (N_1674,N_1268,N_1364);
xor U1675 (N_1675,N_1251,N_1343);
xor U1676 (N_1676,N_1478,N_1432);
nand U1677 (N_1677,N_1361,N_1227);
xor U1678 (N_1678,N_1409,N_1471);
xnor U1679 (N_1679,N_1425,N_1313);
nand U1680 (N_1680,N_1444,N_1447);
and U1681 (N_1681,N_1448,N_1249);
nor U1682 (N_1682,N_1256,N_1228);
and U1683 (N_1683,N_1204,N_1212);
xnor U1684 (N_1684,N_1461,N_1398);
or U1685 (N_1685,N_1206,N_1382);
nand U1686 (N_1686,N_1220,N_1491);
nor U1687 (N_1687,N_1421,N_1466);
or U1688 (N_1688,N_1238,N_1383);
xor U1689 (N_1689,N_1445,N_1436);
and U1690 (N_1690,N_1455,N_1490);
or U1691 (N_1691,N_1391,N_1267);
nand U1692 (N_1692,N_1417,N_1266);
xor U1693 (N_1693,N_1496,N_1413);
nor U1694 (N_1694,N_1269,N_1230);
and U1695 (N_1695,N_1214,N_1301);
nor U1696 (N_1696,N_1227,N_1425);
nand U1697 (N_1697,N_1495,N_1256);
xor U1698 (N_1698,N_1297,N_1263);
and U1699 (N_1699,N_1390,N_1219);
nand U1700 (N_1700,N_1430,N_1429);
nand U1701 (N_1701,N_1366,N_1316);
nor U1702 (N_1702,N_1315,N_1254);
or U1703 (N_1703,N_1276,N_1394);
nand U1704 (N_1704,N_1373,N_1346);
and U1705 (N_1705,N_1360,N_1322);
xor U1706 (N_1706,N_1403,N_1202);
or U1707 (N_1707,N_1371,N_1458);
nand U1708 (N_1708,N_1457,N_1369);
nor U1709 (N_1709,N_1446,N_1318);
nor U1710 (N_1710,N_1279,N_1438);
nor U1711 (N_1711,N_1426,N_1216);
xor U1712 (N_1712,N_1420,N_1314);
and U1713 (N_1713,N_1287,N_1296);
or U1714 (N_1714,N_1305,N_1421);
or U1715 (N_1715,N_1380,N_1464);
nor U1716 (N_1716,N_1246,N_1270);
nand U1717 (N_1717,N_1262,N_1391);
and U1718 (N_1718,N_1402,N_1218);
nor U1719 (N_1719,N_1246,N_1348);
and U1720 (N_1720,N_1348,N_1469);
nor U1721 (N_1721,N_1464,N_1433);
xnor U1722 (N_1722,N_1218,N_1352);
xor U1723 (N_1723,N_1263,N_1281);
nand U1724 (N_1724,N_1374,N_1344);
or U1725 (N_1725,N_1437,N_1480);
nand U1726 (N_1726,N_1390,N_1368);
xor U1727 (N_1727,N_1360,N_1485);
and U1728 (N_1728,N_1397,N_1250);
and U1729 (N_1729,N_1315,N_1277);
and U1730 (N_1730,N_1424,N_1235);
nor U1731 (N_1731,N_1351,N_1426);
and U1732 (N_1732,N_1329,N_1324);
nand U1733 (N_1733,N_1225,N_1452);
xor U1734 (N_1734,N_1224,N_1229);
xor U1735 (N_1735,N_1472,N_1417);
and U1736 (N_1736,N_1242,N_1375);
nand U1737 (N_1737,N_1425,N_1275);
and U1738 (N_1738,N_1316,N_1413);
or U1739 (N_1739,N_1357,N_1458);
nand U1740 (N_1740,N_1465,N_1278);
xor U1741 (N_1741,N_1256,N_1476);
nor U1742 (N_1742,N_1426,N_1403);
nor U1743 (N_1743,N_1442,N_1417);
nor U1744 (N_1744,N_1221,N_1383);
nor U1745 (N_1745,N_1472,N_1461);
nor U1746 (N_1746,N_1203,N_1437);
and U1747 (N_1747,N_1430,N_1454);
or U1748 (N_1748,N_1342,N_1382);
nand U1749 (N_1749,N_1342,N_1324);
or U1750 (N_1750,N_1392,N_1265);
nor U1751 (N_1751,N_1476,N_1370);
nor U1752 (N_1752,N_1358,N_1254);
nand U1753 (N_1753,N_1348,N_1234);
nand U1754 (N_1754,N_1248,N_1377);
and U1755 (N_1755,N_1486,N_1261);
nor U1756 (N_1756,N_1342,N_1287);
nand U1757 (N_1757,N_1450,N_1494);
nor U1758 (N_1758,N_1409,N_1376);
nor U1759 (N_1759,N_1342,N_1486);
xnor U1760 (N_1760,N_1455,N_1200);
nand U1761 (N_1761,N_1407,N_1256);
nand U1762 (N_1762,N_1232,N_1369);
nor U1763 (N_1763,N_1251,N_1256);
or U1764 (N_1764,N_1268,N_1434);
and U1765 (N_1765,N_1391,N_1402);
or U1766 (N_1766,N_1265,N_1249);
and U1767 (N_1767,N_1464,N_1494);
xnor U1768 (N_1768,N_1466,N_1224);
and U1769 (N_1769,N_1304,N_1475);
xor U1770 (N_1770,N_1347,N_1348);
and U1771 (N_1771,N_1416,N_1352);
nor U1772 (N_1772,N_1330,N_1384);
and U1773 (N_1773,N_1354,N_1419);
nor U1774 (N_1774,N_1289,N_1226);
or U1775 (N_1775,N_1439,N_1327);
xnor U1776 (N_1776,N_1237,N_1281);
and U1777 (N_1777,N_1474,N_1226);
nor U1778 (N_1778,N_1287,N_1456);
nor U1779 (N_1779,N_1431,N_1202);
nor U1780 (N_1780,N_1354,N_1367);
and U1781 (N_1781,N_1398,N_1311);
nor U1782 (N_1782,N_1461,N_1325);
nand U1783 (N_1783,N_1373,N_1257);
nand U1784 (N_1784,N_1451,N_1272);
or U1785 (N_1785,N_1315,N_1322);
nand U1786 (N_1786,N_1255,N_1214);
and U1787 (N_1787,N_1412,N_1206);
or U1788 (N_1788,N_1268,N_1357);
and U1789 (N_1789,N_1389,N_1457);
nand U1790 (N_1790,N_1439,N_1365);
and U1791 (N_1791,N_1219,N_1460);
and U1792 (N_1792,N_1476,N_1244);
xnor U1793 (N_1793,N_1437,N_1266);
nor U1794 (N_1794,N_1278,N_1393);
xor U1795 (N_1795,N_1454,N_1475);
or U1796 (N_1796,N_1376,N_1483);
nor U1797 (N_1797,N_1476,N_1494);
or U1798 (N_1798,N_1443,N_1332);
nor U1799 (N_1799,N_1346,N_1359);
nor U1800 (N_1800,N_1791,N_1519);
or U1801 (N_1801,N_1688,N_1756);
or U1802 (N_1802,N_1629,N_1727);
nand U1803 (N_1803,N_1511,N_1732);
nand U1804 (N_1804,N_1643,N_1521);
and U1805 (N_1805,N_1589,N_1799);
nand U1806 (N_1806,N_1648,N_1744);
xor U1807 (N_1807,N_1579,N_1628);
nand U1808 (N_1808,N_1785,N_1552);
or U1809 (N_1809,N_1584,N_1750);
and U1810 (N_1810,N_1696,N_1792);
or U1811 (N_1811,N_1630,N_1562);
or U1812 (N_1812,N_1613,N_1522);
nand U1813 (N_1813,N_1678,N_1534);
or U1814 (N_1814,N_1614,N_1617);
or U1815 (N_1815,N_1590,N_1777);
xnor U1816 (N_1816,N_1707,N_1671);
nand U1817 (N_1817,N_1760,N_1669);
nand U1818 (N_1818,N_1660,N_1586);
and U1819 (N_1819,N_1743,N_1788);
nand U1820 (N_1820,N_1507,N_1553);
nor U1821 (N_1821,N_1639,N_1758);
nand U1822 (N_1822,N_1625,N_1506);
xnor U1823 (N_1823,N_1631,N_1615);
or U1824 (N_1824,N_1704,N_1626);
and U1825 (N_1825,N_1599,N_1752);
nor U1826 (N_1826,N_1555,N_1773);
or U1827 (N_1827,N_1702,N_1762);
nor U1828 (N_1828,N_1650,N_1528);
and U1829 (N_1829,N_1588,N_1646);
xnor U1830 (N_1830,N_1776,N_1537);
nor U1831 (N_1831,N_1736,N_1547);
nand U1832 (N_1832,N_1708,N_1618);
nor U1833 (N_1833,N_1602,N_1544);
xnor U1834 (N_1834,N_1711,N_1719);
and U1835 (N_1835,N_1716,N_1573);
and U1836 (N_1836,N_1748,N_1657);
xor U1837 (N_1837,N_1763,N_1582);
nand U1838 (N_1838,N_1782,N_1606);
nand U1839 (N_1839,N_1765,N_1778);
nor U1840 (N_1840,N_1523,N_1500);
and U1841 (N_1841,N_1635,N_1638);
nor U1842 (N_1842,N_1786,N_1718);
nand U1843 (N_1843,N_1580,N_1572);
xor U1844 (N_1844,N_1520,N_1661);
nand U1845 (N_1845,N_1633,N_1510);
nor U1846 (N_1846,N_1681,N_1566);
xnor U1847 (N_1847,N_1608,N_1738);
or U1848 (N_1848,N_1766,N_1609);
nand U1849 (N_1849,N_1714,N_1593);
nand U1850 (N_1850,N_1749,N_1710);
nor U1851 (N_1851,N_1601,N_1793);
or U1852 (N_1852,N_1790,N_1612);
or U1853 (N_1853,N_1787,N_1538);
nor U1854 (N_1854,N_1774,N_1771);
nand U1855 (N_1855,N_1649,N_1619);
or U1856 (N_1856,N_1616,N_1622);
xnor U1857 (N_1857,N_1741,N_1742);
nand U1858 (N_1858,N_1662,N_1699);
xnor U1859 (N_1859,N_1533,N_1740);
nand U1860 (N_1860,N_1642,N_1715);
nand U1861 (N_1861,N_1682,N_1583);
nor U1862 (N_1862,N_1685,N_1739);
xor U1863 (N_1863,N_1693,N_1755);
or U1864 (N_1864,N_1564,N_1529);
nor U1865 (N_1865,N_1568,N_1632);
nor U1866 (N_1866,N_1652,N_1559);
or U1867 (N_1867,N_1546,N_1605);
and U1868 (N_1868,N_1517,N_1666);
xnor U1869 (N_1869,N_1581,N_1737);
and U1870 (N_1870,N_1717,N_1607);
nand U1871 (N_1871,N_1767,N_1587);
xnor U1872 (N_1872,N_1591,N_1541);
or U1873 (N_1873,N_1677,N_1734);
xnor U1874 (N_1874,N_1508,N_1745);
nor U1875 (N_1875,N_1668,N_1723);
and U1876 (N_1876,N_1620,N_1576);
xnor U1877 (N_1877,N_1664,N_1751);
and U1878 (N_1878,N_1563,N_1554);
nand U1879 (N_1879,N_1504,N_1784);
or U1880 (N_1880,N_1575,N_1543);
or U1881 (N_1881,N_1595,N_1753);
xor U1882 (N_1882,N_1536,N_1781);
nor U1883 (N_1883,N_1574,N_1644);
xnor U1884 (N_1884,N_1675,N_1689);
nand U1885 (N_1885,N_1789,N_1700);
and U1886 (N_1886,N_1663,N_1641);
and U1887 (N_1887,N_1516,N_1721);
xnor U1888 (N_1888,N_1526,N_1501);
and U1889 (N_1889,N_1532,N_1513);
or U1890 (N_1890,N_1694,N_1712);
and U1891 (N_1891,N_1597,N_1687);
nor U1892 (N_1892,N_1656,N_1515);
or U1893 (N_1893,N_1690,N_1624);
nand U1894 (N_1894,N_1684,N_1670);
and U1895 (N_1895,N_1735,N_1542);
or U1896 (N_1896,N_1540,N_1557);
nand U1897 (N_1897,N_1713,N_1621);
xnor U1898 (N_1898,N_1747,N_1779);
and U1899 (N_1899,N_1565,N_1505);
nand U1900 (N_1900,N_1610,N_1550);
xor U1901 (N_1901,N_1794,N_1725);
nor U1902 (N_1902,N_1764,N_1724);
nor U1903 (N_1903,N_1667,N_1640);
and U1904 (N_1904,N_1634,N_1659);
and U1905 (N_1905,N_1592,N_1509);
xnor U1906 (N_1906,N_1775,N_1558);
nand U1907 (N_1907,N_1623,N_1604);
nand U1908 (N_1908,N_1705,N_1706);
xnor U1909 (N_1909,N_1731,N_1754);
and U1910 (N_1910,N_1654,N_1759);
nand U1911 (N_1911,N_1655,N_1549);
and U1912 (N_1912,N_1698,N_1561);
nand U1913 (N_1913,N_1795,N_1567);
xor U1914 (N_1914,N_1676,N_1535);
or U1915 (N_1915,N_1530,N_1701);
or U1916 (N_1916,N_1672,N_1556);
xnor U1917 (N_1917,N_1729,N_1545);
nand U1918 (N_1918,N_1658,N_1636);
or U1919 (N_1919,N_1524,N_1578);
or U1920 (N_1920,N_1673,N_1514);
xnor U1921 (N_1921,N_1570,N_1611);
and U1922 (N_1922,N_1730,N_1502);
and U1923 (N_1923,N_1598,N_1772);
nand U1924 (N_1924,N_1695,N_1637);
nand U1925 (N_1925,N_1674,N_1770);
nor U1926 (N_1926,N_1525,N_1569);
or U1927 (N_1927,N_1577,N_1518);
xnor U1928 (N_1928,N_1722,N_1703);
nand U1929 (N_1929,N_1798,N_1680);
xnor U1930 (N_1930,N_1548,N_1728);
nor U1931 (N_1931,N_1603,N_1757);
xor U1932 (N_1932,N_1665,N_1683);
and U1933 (N_1933,N_1761,N_1653);
or U1934 (N_1934,N_1697,N_1679);
nand U1935 (N_1935,N_1746,N_1780);
nand U1936 (N_1936,N_1600,N_1551);
and U1937 (N_1937,N_1594,N_1691);
or U1938 (N_1938,N_1797,N_1571);
nor U1939 (N_1939,N_1783,N_1627);
or U1940 (N_1940,N_1709,N_1512);
and U1941 (N_1941,N_1596,N_1527);
nand U1942 (N_1942,N_1720,N_1769);
and U1943 (N_1943,N_1692,N_1585);
or U1944 (N_1944,N_1733,N_1503);
nand U1945 (N_1945,N_1539,N_1686);
and U1946 (N_1946,N_1796,N_1560);
xor U1947 (N_1947,N_1647,N_1531);
or U1948 (N_1948,N_1651,N_1768);
nand U1949 (N_1949,N_1645,N_1726);
xnor U1950 (N_1950,N_1768,N_1753);
nor U1951 (N_1951,N_1573,N_1622);
nor U1952 (N_1952,N_1530,N_1548);
nor U1953 (N_1953,N_1734,N_1724);
or U1954 (N_1954,N_1766,N_1532);
or U1955 (N_1955,N_1752,N_1538);
or U1956 (N_1956,N_1601,N_1650);
nand U1957 (N_1957,N_1564,N_1596);
xnor U1958 (N_1958,N_1506,N_1551);
nand U1959 (N_1959,N_1733,N_1589);
nor U1960 (N_1960,N_1577,N_1635);
and U1961 (N_1961,N_1541,N_1662);
and U1962 (N_1962,N_1562,N_1665);
nand U1963 (N_1963,N_1691,N_1766);
nand U1964 (N_1964,N_1663,N_1690);
nor U1965 (N_1965,N_1577,N_1746);
xnor U1966 (N_1966,N_1526,N_1574);
or U1967 (N_1967,N_1625,N_1693);
nor U1968 (N_1968,N_1613,N_1695);
nor U1969 (N_1969,N_1634,N_1520);
nor U1970 (N_1970,N_1666,N_1510);
or U1971 (N_1971,N_1648,N_1729);
nor U1972 (N_1972,N_1550,N_1504);
or U1973 (N_1973,N_1681,N_1512);
nand U1974 (N_1974,N_1506,N_1679);
or U1975 (N_1975,N_1601,N_1778);
xor U1976 (N_1976,N_1764,N_1512);
or U1977 (N_1977,N_1591,N_1536);
xnor U1978 (N_1978,N_1535,N_1662);
or U1979 (N_1979,N_1761,N_1652);
xnor U1980 (N_1980,N_1540,N_1675);
nor U1981 (N_1981,N_1734,N_1592);
nor U1982 (N_1982,N_1626,N_1672);
and U1983 (N_1983,N_1787,N_1572);
xnor U1984 (N_1984,N_1698,N_1668);
or U1985 (N_1985,N_1563,N_1589);
and U1986 (N_1986,N_1651,N_1608);
nor U1987 (N_1987,N_1586,N_1509);
and U1988 (N_1988,N_1543,N_1651);
or U1989 (N_1989,N_1594,N_1510);
or U1990 (N_1990,N_1689,N_1592);
nand U1991 (N_1991,N_1501,N_1721);
nor U1992 (N_1992,N_1502,N_1749);
and U1993 (N_1993,N_1715,N_1678);
or U1994 (N_1994,N_1797,N_1651);
or U1995 (N_1995,N_1792,N_1740);
nand U1996 (N_1996,N_1757,N_1652);
or U1997 (N_1997,N_1661,N_1681);
nand U1998 (N_1998,N_1581,N_1519);
nand U1999 (N_1999,N_1617,N_1644);
or U2000 (N_2000,N_1511,N_1515);
or U2001 (N_2001,N_1556,N_1666);
nand U2002 (N_2002,N_1590,N_1769);
and U2003 (N_2003,N_1625,N_1538);
nor U2004 (N_2004,N_1637,N_1545);
nand U2005 (N_2005,N_1545,N_1506);
and U2006 (N_2006,N_1744,N_1597);
nor U2007 (N_2007,N_1552,N_1677);
or U2008 (N_2008,N_1797,N_1706);
nor U2009 (N_2009,N_1667,N_1783);
xnor U2010 (N_2010,N_1537,N_1746);
nand U2011 (N_2011,N_1781,N_1552);
nor U2012 (N_2012,N_1567,N_1544);
and U2013 (N_2013,N_1505,N_1553);
nand U2014 (N_2014,N_1718,N_1607);
xnor U2015 (N_2015,N_1556,N_1733);
nor U2016 (N_2016,N_1628,N_1580);
xnor U2017 (N_2017,N_1518,N_1655);
nor U2018 (N_2018,N_1526,N_1711);
nor U2019 (N_2019,N_1640,N_1643);
nor U2020 (N_2020,N_1724,N_1617);
and U2021 (N_2021,N_1623,N_1570);
nor U2022 (N_2022,N_1706,N_1718);
nor U2023 (N_2023,N_1595,N_1780);
or U2024 (N_2024,N_1736,N_1779);
and U2025 (N_2025,N_1757,N_1722);
nor U2026 (N_2026,N_1773,N_1521);
or U2027 (N_2027,N_1692,N_1631);
xor U2028 (N_2028,N_1790,N_1575);
and U2029 (N_2029,N_1797,N_1616);
nand U2030 (N_2030,N_1512,N_1743);
xor U2031 (N_2031,N_1710,N_1673);
or U2032 (N_2032,N_1692,N_1604);
xor U2033 (N_2033,N_1738,N_1505);
or U2034 (N_2034,N_1774,N_1707);
or U2035 (N_2035,N_1769,N_1733);
xor U2036 (N_2036,N_1737,N_1723);
and U2037 (N_2037,N_1508,N_1733);
nor U2038 (N_2038,N_1515,N_1645);
or U2039 (N_2039,N_1539,N_1591);
or U2040 (N_2040,N_1626,N_1512);
and U2041 (N_2041,N_1523,N_1708);
nor U2042 (N_2042,N_1579,N_1521);
nand U2043 (N_2043,N_1690,N_1661);
nand U2044 (N_2044,N_1765,N_1757);
xnor U2045 (N_2045,N_1535,N_1741);
or U2046 (N_2046,N_1547,N_1683);
nand U2047 (N_2047,N_1630,N_1525);
nand U2048 (N_2048,N_1622,N_1721);
and U2049 (N_2049,N_1640,N_1588);
xnor U2050 (N_2050,N_1763,N_1663);
or U2051 (N_2051,N_1791,N_1574);
or U2052 (N_2052,N_1637,N_1770);
nor U2053 (N_2053,N_1531,N_1773);
xnor U2054 (N_2054,N_1658,N_1702);
xor U2055 (N_2055,N_1526,N_1628);
or U2056 (N_2056,N_1682,N_1726);
nand U2057 (N_2057,N_1762,N_1607);
or U2058 (N_2058,N_1768,N_1535);
or U2059 (N_2059,N_1606,N_1674);
nand U2060 (N_2060,N_1589,N_1734);
nand U2061 (N_2061,N_1560,N_1583);
and U2062 (N_2062,N_1685,N_1553);
nor U2063 (N_2063,N_1516,N_1581);
and U2064 (N_2064,N_1763,N_1600);
or U2065 (N_2065,N_1633,N_1677);
and U2066 (N_2066,N_1611,N_1723);
nor U2067 (N_2067,N_1593,N_1627);
or U2068 (N_2068,N_1659,N_1721);
xnor U2069 (N_2069,N_1567,N_1578);
and U2070 (N_2070,N_1518,N_1670);
and U2071 (N_2071,N_1746,N_1774);
nor U2072 (N_2072,N_1501,N_1707);
nand U2073 (N_2073,N_1617,N_1616);
xor U2074 (N_2074,N_1526,N_1557);
and U2075 (N_2075,N_1731,N_1503);
xor U2076 (N_2076,N_1589,N_1507);
and U2077 (N_2077,N_1623,N_1688);
or U2078 (N_2078,N_1597,N_1609);
xnor U2079 (N_2079,N_1588,N_1775);
or U2080 (N_2080,N_1759,N_1532);
and U2081 (N_2081,N_1660,N_1512);
nand U2082 (N_2082,N_1776,N_1528);
nand U2083 (N_2083,N_1684,N_1583);
or U2084 (N_2084,N_1677,N_1684);
nor U2085 (N_2085,N_1632,N_1635);
nand U2086 (N_2086,N_1555,N_1556);
xor U2087 (N_2087,N_1660,N_1526);
or U2088 (N_2088,N_1525,N_1733);
nand U2089 (N_2089,N_1779,N_1700);
xnor U2090 (N_2090,N_1587,N_1739);
and U2091 (N_2091,N_1622,N_1525);
xor U2092 (N_2092,N_1532,N_1640);
and U2093 (N_2093,N_1680,N_1706);
nand U2094 (N_2094,N_1748,N_1572);
nor U2095 (N_2095,N_1713,N_1659);
nor U2096 (N_2096,N_1754,N_1672);
or U2097 (N_2097,N_1724,N_1684);
or U2098 (N_2098,N_1757,N_1771);
nor U2099 (N_2099,N_1648,N_1550);
and U2100 (N_2100,N_1801,N_1914);
nand U2101 (N_2101,N_1804,N_2093);
nor U2102 (N_2102,N_2007,N_2045);
nor U2103 (N_2103,N_1937,N_2022);
and U2104 (N_2104,N_2037,N_2038);
nor U2105 (N_2105,N_2089,N_1839);
xnor U2106 (N_2106,N_1819,N_2086);
nand U2107 (N_2107,N_2071,N_1959);
and U2108 (N_2108,N_2051,N_1889);
nor U2109 (N_2109,N_1953,N_2061);
and U2110 (N_2110,N_2048,N_2033);
nor U2111 (N_2111,N_2063,N_2017);
xor U2112 (N_2112,N_2015,N_1882);
and U2113 (N_2113,N_2013,N_1848);
xnor U2114 (N_2114,N_2006,N_1925);
xor U2115 (N_2115,N_1960,N_1892);
nor U2116 (N_2116,N_1815,N_2052);
nand U2117 (N_2117,N_1850,N_1931);
xnor U2118 (N_2118,N_1821,N_1946);
or U2119 (N_2119,N_1849,N_1825);
and U2120 (N_2120,N_1814,N_1807);
xor U2121 (N_2121,N_1993,N_1928);
xnor U2122 (N_2122,N_1813,N_2055);
xnor U2123 (N_2123,N_1851,N_1836);
nand U2124 (N_2124,N_1843,N_1981);
xnor U2125 (N_2125,N_1955,N_1888);
xor U2126 (N_2126,N_1929,N_1861);
and U2127 (N_2127,N_1958,N_1980);
xor U2128 (N_2128,N_1846,N_1820);
xor U2129 (N_2129,N_2040,N_1844);
nor U2130 (N_2130,N_1969,N_2011);
nand U2131 (N_2131,N_2036,N_1853);
or U2132 (N_2132,N_1874,N_1833);
and U2133 (N_2133,N_1965,N_1950);
nand U2134 (N_2134,N_1999,N_2009);
nand U2135 (N_2135,N_2059,N_2034);
nand U2136 (N_2136,N_2004,N_1816);
nor U2137 (N_2137,N_1904,N_1824);
xnor U2138 (N_2138,N_1898,N_1802);
nand U2139 (N_2139,N_2088,N_1913);
and U2140 (N_2140,N_1910,N_1989);
nor U2141 (N_2141,N_1970,N_2054);
or U2142 (N_2142,N_1978,N_1944);
xor U2143 (N_2143,N_2049,N_2066);
or U2144 (N_2144,N_2095,N_2041);
nand U2145 (N_2145,N_2075,N_1936);
and U2146 (N_2146,N_1922,N_2029);
or U2147 (N_2147,N_1903,N_1962);
nand U2148 (N_2148,N_2050,N_1876);
or U2149 (N_2149,N_1890,N_1964);
nand U2150 (N_2150,N_1905,N_1859);
nor U2151 (N_2151,N_2043,N_1941);
nand U2152 (N_2152,N_1883,N_2053);
or U2153 (N_2153,N_2035,N_2062);
and U2154 (N_2154,N_1995,N_1907);
nor U2155 (N_2155,N_1900,N_1948);
and U2156 (N_2156,N_1939,N_1854);
nand U2157 (N_2157,N_2042,N_1826);
and U2158 (N_2158,N_2039,N_1996);
xnor U2159 (N_2159,N_2069,N_2008);
or U2160 (N_2160,N_1871,N_1856);
xnor U2161 (N_2161,N_2012,N_1884);
xnor U2162 (N_2162,N_1855,N_1829);
nor U2163 (N_2163,N_1986,N_1895);
and U2164 (N_2164,N_1915,N_2091);
or U2165 (N_2165,N_1886,N_2000);
and U2166 (N_2166,N_2047,N_1831);
nand U2167 (N_2167,N_1911,N_2057);
xnor U2168 (N_2168,N_2014,N_1908);
nand U2169 (N_2169,N_1998,N_2090);
nor U2170 (N_2170,N_1835,N_1817);
or U2171 (N_2171,N_1988,N_2072);
and U2172 (N_2172,N_1920,N_1943);
and U2173 (N_2173,N_1896,N_2077);
nor U2174 (N_2174,N_1897,N_2074);
nand U2175 (N_2175,N_1982,N_1909);
and U2176 (N_2176,N_1935,N_1881);
or U2177 (N_2177,N_1997,N_1860);
nor U2178 (N_2178,N_2030,N_1879);
or U2179 (N_2179,N_1869,N_1934);
and U2180 (N_2180,N_2031,N_1901);
and U2181 (N_2181,N_2098,N_1923);
nor U2182 (N_2182,N_1880,N_1838);
and U2183 (N_2183,N_1985,N_1976);
nand U2184 (N_2184,N_1891,N_1823);
nor U2185 (N_2185,N_2070,N_2094);
and U2186 (N_2186,N_1974,N_2080);
xor U2187 (N_2187,N_1906,N_1872);
and U2188 (N_2188,N_1811,N_1868);
xnor U2189 (N_2189,N_1864,N_1977);
xor U2190 (N_2190,N_1847,N_2068);
or U2191 (N_2191,N_2056,N_1966);
or U2192 (N_2192,N_1822,N_2084);
or U2193 (N_2193,N_1887,N_2092);
nand U2194 (N_2194,N_1912,N_1806);
nor U2195 (N_2195,N_2067,N_2099);
nor U2196 (N_2196,N_1952,N_2073);
nor U2197 (N_2197,N_1875,N_2005);
or U2198 (N_2198,N_1932,N_2018);
or U2199 (N_2199,N_1899,N_1991);
xnor U2200 (N_2200,N_1885,N_1916);
xnor U2201 (N_2201,N_2020,N_2058);
and U2202 (N_2202,N_1862,N_1963);
and U2203 (N_2203,N_1968,N_1921);
nor U2204 (N_2204,N_1990,N_2024);
xnor U2205 (N_2205,N_2082,N_2096);
nor U2206 (N_2206,N_1930,N_1878);
nand U2207 (N_2207,N_1834,N_1832);
xnor U2208 (N_2208,N_1947,N_1902);
or U2209 (N_2209,N_1873,N_2003);
or U2210 (N_2210,N_1945,N_1992);
or U2211 (N_2211,N_2046,N_1877);
nand U2212 (N_2212,N_1987,N_1949);
nor U2213 (N_2213,N_2079,N_1830);
nand U2214 (N_2214,N_1857,N_2081);
or U2215 (N_2215,N_1867,N_1866);
nand U2216 (N_2216,N_1973,N_1810);
nand U2217 (N_2217,N_1858,N_2032);
or U2218 (N_2218,N_1800,N_2097);
nor U2219 (N_2219,N_2044,N_1961);
or U2220 (N_2220,N_1942,N_2064);
and U2221 (N_2221,N_1852,N_2016);
nor U2222 (N_2222,N_1803,N_1926);
xnor U2223 (N_2223,N_2023,N_1828);
xnor U2224 (N_2224,N_2028,N_2083);
xor U2225 (N_2225,N_1972,N_1924);
and U2226 (N_2226,N_1983,N_1984);
nand U2227 (N_2227,N_1840,N_1956);
or U2228 (N_2228,N_1933,N_2019);
nor U2229 (N_2229,N_1805,N_1827);
or U2230 (N_2230,N_2026,N_1918);
nand U2231 (N_2231,N_1870,N_2025);
xor U2232 (N_2232,N_2085,N_2021);
and U2233 (N_2233,N_1837,N_1954);
xor U2234 (N_2234,N_1841,N_1809);
nor U2235 (N_2235,N_2060,N_1842);
or U2236 (N_2236,N_1975,N_1994);
nand U2237 (N_2237,N_2087,N_1893);
nor U2238 (N_2238,N_1808,N_1865);
or U2239 (N_2239,N_2001,N_2002);
nand U2240 (N_2240,N_1971,N_2065);
nand U2241 (N_2241,N_1957,N_1917);
nand U2242 (N_2242,N_2078,N_1863);
nand U2243 (N_2243,N_1919,N_1938);
or U2244 (N_2244,N_1979,N_1812);
nand U2245 (N_2245,N_1894,N_1845);
nand U2246 (N_2246,N_2027,N_2010);
xnor U2247 (N_2247,N_1940,N_1951);
or U2248 (N_2248,N_1927,N_1967);
nand U2249 (N_2249,N_2076,N_1818);
or U2250 (N_2250,N_1822,N_1813);
nor U2251 (N_2251,N_1934,N_1817);
nor U2252 (N_2252,N_1876,N_2015);
xor U2253 (N_2253,N_2035,N_2047);
and U2254 (N_2254,N_1979,N_2025);
and U2255 (N_2255,N_1882,N_1937);
nor U2256 (N_2256,N_2012,N_1952);
xor U2257 (N_2257,N_1801,N_1972);
and U2258 (N_2258,N_1880,N_1832);
nand U2259 (N_2259,N_1831,N_1935);
and U2260 (N_2260,N_2070,N_1958);
xor U2261 (N_2261,N_1888,N_1811);
or U2262 (N_2262,N_2066,N_1902);
and U2263 (N_2263,N_1884,N_1978);
xnor U2264 (N_2264,N_2096,N_1892);
nand U2265 (N_2265,N_1895,N_1838);
nand U2266 (N_2266,N_2001,N_2040);
or U2267 (N_2267,N_1943,N_1887);
or U2268 (N_2268,N_1894,N_2000);
nor U2269 (N_2269,N_1973,N_2047);
or U2270 (N_2270,N_1812,N_2094);
or U2271 (N_2271,N_2027,N_2062);
xor U2272 (N_2272,N_1885,N_2010);
xor U2273 (N_2273,N_1835,N_1958);
nor U2274 (N_2274,N_2094,N_1909);
and U2275 (N_2275,N_2073,N_1840);
nor U2276 (N_2276,N_1853,N_1870);
xor U2277 (N_2277,N_2068,N_1971);
nand U2278 (N_2278,N_2023,N_1857);
nand U2279 (N_2279,N_1863,N_1988);
nand U2280 (N_2280,N_1978,N_1998);
xor U2281 (N_2281,N_2018,N_2016);
and U2282 (N_2282,N_1989,N_2093);
nand U2283 (N_2283,N_1871,N_1970);
or U2284 (N_2284,N_2000,N_1948);
and U2285 (N_2285,N_2051,N_2095);
nand U2286 (N_2286,N_2007,N_2035);
nor U2287 (N_2287,N_1944,N_2065);
xor U2288 (N_2288,N_2013,N_1876);
and U2289 (N_2289,N_1840,N_2077);
and U2290 (N_2290,N_1940,N_2022);
nor U2291 (N_2291,N_1832,N_2069);
and U2292 (N_2292,N_2016,N_1929);
xor U2293 (N_2293,N_1805,N_1826);
or U2294 (N_2294,N_2093,N_1988);
or U2295 (N_2295,N_1965,N_2091);
xnor U2296 (N_2296,N_2015,N_2090);
xor U2297 (N_2297,N_2021,N_1847);
or U2298 (N_2298,N_1997,N_1973);
nor U2299 (N_2299,N_1815,N_1980);
nor U2300 (N_2300,N_1951,N_1903);
xor U2301 (N_2301,N_2069,N_1863);
and U2302 (N_2302,N_2024,N_1911);
or U2303 (N_2303,N_1851,N_1827);
or U2304 (N_2304,N_1995,N_1809);
and U2305 (N_2305,N_2057,N_1842);
or U2306 (N_2306,N_2030,N_1942);
nor U2307 (N_2307,N_1906,N_1810);
and U2308 (N_2308,N_2040,N_1875);
or U2309 (N_2309,N_1925,N_2049);
or U2310 (N_2310,N_1989,N_2080);
nand U2311 (N_2311,N_1977,N_2064);
nand U2312 (N_2312,N_2048,N_1832);
and U2313 (N_2313,N_2032,N_2083);
or U2314 (N_2314,N_1867,N_1970);
xor U2315 (N_2315,N_2066,N_1989);
or U2316 (N_2316,N_1891,N_1901);
nand U2317 (N_2317,N_1961,N_1856);
or U2318 (N_2318,N_1922,N_1967);
nand U2319 (N_2319,N_2027,N_1940);
nand U2320 (N_2320,N_1893,N_1827);
or U2321 (N_2321,N_1999,N_1959);
nand U2322 (N_2322,N_2023,N_1921);
nand U2323 (N_2323,N_1822,N_1915);
xnor U2324 (N_2324,N_2093,N_1822);
xnor U2325 (N_2325,N_1835,N_1924);
or U2326 (N_2326,N_2091,N_1866);
nor U2327 (N_2327,N_1947,N_1879);
nand U2328 (N_2328,N_2004,N_2081);
nor U2329 (N_2329,N_2050,N_1962);
nor U2330 (N_2330,N_2064,N_2020);
and U2331 (N_2331,N_1817,N_1908);
nand U2332 (N_2332,N_2018,N_1923);
xnor U2333 (N_2333,N_2074,N_1931);
nor U2334 (N_2334,N_1945,N_1969);
nand U2335 (N_2335,N_1990,N_2007);
xor U2336 (N_2336,N_1883,N_2023);
nand U2337 (N_2337,N_1869,N_1865);
or U2338 (N_2338,N_2098,N_1943);
nor U2339 (N_2339,N_1917,N_1978);
xnor U2340 (N_2340,N_2080,N_1905);
xor U2341 (N_2341,N_1827,N_2018);
or U2342 (N_2342,N_1942,N_1906);
and U2343 (N_2343,N_1934,N_1995);
xor U2344 (N_2344,N_1993,N_1951);
nand U2345 (N_2345,N_1888,N_1953);
nand U2346 (N_2346,N_1970,N_2005);
nand U2347 (N_2347,N_1931,N_2006);
nand U2348 (N_2348,N_2091,N_1820);
and U2349 (N_2349,N_1904,N_1801);
xor U2350 (N_2350,N_1979,N_1949);
and U2351 (N_2351,N_2008,N_1910);
xor U2352 (N_2352,N_1839,N_1861);
nand U2353 (N_2353,N_2023,N_1940);
nor U2354 (N_2354,N_1996,N_1852);
or U2355 (N_2355,N_1974,N_1923);
nand U2356 (N_2356,N_2003,N_1910);
or U2357 (N_2357,N_2008,N_1856);
or U2358 (N_2358,N_1861,N_1977);
nand U2359 (N_2359,N_1880,N_1800);
or U2360 (N_2360,N_1839,N_2099);
and U2361 (N_2361,N_1989,N_2070);
and U2362 (N_2362,N_1974,N_1949);
nor U2363 (N_2363,N_1892,N_1950);
xor U2364 (N_2364,N_1884,N_1803);
xor U2365 (N_2365,N_2007,N_1886);
and U2366 (N_2366,N_1928,N_2077);
or U2367 (N_2367,N_1984,N_2017);
xnor U2368 (N_2368,N_1835,N_1956);
nand U2369 (N_2369,N_1996,N_2091);
nor U2370 (N_2370,N_1844,N_1995);
nor U2371 (N_2371,N_2056,N_1809);
nor U2372 (N_2372,N_1858,N_2006);
nor U2373 (N_2373,N_1927,N_1943);
nor U2374 (N_2374,N_1925,N_2066);
nand U2375 (N_2375,N_2088,N_1942);
and U2376 (N_2376,N_1930,N_1817);
or U2377 (N_2377,N_1971,N_1872);
nor U2378 (N_2378,N_1843,N_1884);
nor U2379 (N_2379,N_1968,N_1941);
nand U2380 (N_2380,N_1862,N_1970);
nand U2381 (N_2381,N_1954,N_1931);
nand U2382 (N_2382,N_1968,N_1987);
or U2383 (N_2383,N_2074,N_1954);
or U2384 (N_2384,N_2051,N_1893);
and U2385 (N_2385,N_1827,N_2060);
and U2386 (N_2386,N_2052,N_1823);
nor U2387 (N_2387,N_1891,N_1914);
nor U2388 (N_2388,N_1838,N_1918);
and U2389 (N_2389,N_1970,N_1854);
and U2390 (N_2390,N_1940,N_2085);
nor U2391 (N_2391,N_1979,N_2078);
and U2392 (N_2392,N_1908,N_1953);
nand U2393 (N_2393,N_2063,N_1918);
xnor U2394 (N_2394,N_1927,N_2008);
xnor U2395 (N_2395,N_1950,N_2089);
and U2396 (N_2396,N_1865,N_1835);
and U2397 (N_2397,N_2036,N_1824);
or U2398 (N_2398,N_1980,N_1874);
nor U2399 (N_2399,N_1952,N_1946);
nor U2400 (N_2400,N_2317,N_2152);
nor U2401 (N_2401,N_2339,N_2290);
nand U2402 (N_2402,N_2258,N_2250);
and U2403 (N_2403,N_2223,N_2108);
or U2404 (N_2404,N_2120,N_2213);
nand U2405 (N_2405,N_2107,N_2170);
xor U2406 (N_2406,N_2142,N_2364);
nor U2407 (N_2407,N_2115,N_2116);
or U2408 (N_2408,N_2201,N_2230);
nand U2409 (N_2409,N_2200,N_2157);
or U2410 (N_2410,N_2246,N_2355);
or U2411 (N_2411,N_2352,N_2338);
xnor U2412 (N_2412,N_2191,N_2153);
and U2413 (N_2413,N_2242,N_2117);
and U2414 (N_2414,N_2212,N_2381);
or U2415 (N_2415,N_2249,N_2244);
or U2416 (N_2416,N_2394,N_2268);
xor U2417 (N_2417,N_2270,N_2390);
nand U2418 (N_2418,N_2294,N_2332);
nand U2419 (N_2419,N_2251,N_2276);
or U2420 (N_2420,N_2101,N_2374);
nor U2421 (N_2421,N_2112,N_2126);
nand U2422 (N_2422,N_2285,N_2214);
nand U2423 (N_2423,N_2102,N_2243);
nand U2424 (N_2424,N_2344,N_2316);
nand U2425 (N_2425,N_2202,N_2193);
nor U2426 (N_2426,N_2347,N_2354);
or U2427 (N_2427,N_2398,N_2129);
xor U2428 (N_2428,N_2369,N_2122);
and U2429 (N_2429,N_2124,N_2211);
nor U2430 (N_2430,N_2391,N_2334);
xnor U2431 (N_2431,N_2240,N_2169);
nor U2432 (N_2432,N_2386,N_2209);
nand U2433 (N_2433,N_2280,N_2205);
xnor U2434 (N_2434,N_2306,N_2283);
nand U2435 (N_2435,N_2143,N_2395);
nand U2436 (N_2436,N_2301,N_2151);
or U2437 (N_2437,N_2217,N_2207);
or U2438 (N_2438,N_2293,N_2133);
nand U2439 (N_2439,N_2172,N_2300);
or U2440 (N_2440,N_2125,N_2262);
and U2441 (N_2441,N_2164,N_2229);
nand U2442 (N_2442,N_2315,N_2127);
xnor U2443 (N_2443,N_2247,N_2224);
and U2444 (N_2444,N_2330,N_2357);
xor U2445 (N_2445,N_2148,N_2239);
or U2446 (N_2446,N_2171,N_2254);
xnor U2447 (N_2447,N_2371,N_2144);
or U2448 (N_2448,N_2118,N_2376);
nand U2449 (N_2449,N_2296,N_2181);
nor U2450 (N_2450,N_2324,N_2168);
xor U2451 (N_2451,N_2277,N_2389);
xor U2452 (N_2452,N_2308,N_2110);
nand U2453 (N_2453,N_2311,N_2342);
nand U2454 (N_2454,N_2208,N_2196);
or U2455 (N_2455,N_2165,N_2192);
nor U2456 (N_2456,N_2138,N_2275);
and U2457 (N_2457,N_2333,N_2385);
nor U2458 (N_2458,N_2360,N_2139);
and U2459 (N_2459,N_2287,N_2366);
or U2460 (N_2460,N_2237,N_2348);
xor U2461 (N_2461,N_2216,N_2248);
and U2462 (N_2462,N_2255,N_2182);
and U2463 (N_2463,N_2372,N_2259);
or U2464 (N_2464,N_2264,N_2174);
or U2465 (N_2465,N_2187,N_2314);
or U2466 (N_2466,N_2121,N_2161);
nor U2467 (N_2467,N_2197,N_2384);
or U2468 (N_2468,N_2309,N_2323);
or U2469 (N_2469,N_2328,N_2377);
or U2470 (N_2470,N_2286,N_2111);
nor U2471 (N_2471,N_2104,N_2326);
nor U2472 (N_2472,N_2325,N_2396);
nor U2473 (N_2473,N_2199,N_2253);
nor U2474 (N_2474,N_2362,N_2319);
and U2475 (N_2475,N_2204,N_2278);
and U2476 (N_2476,N_2173,N_2341);
and U2477 (N_2477,N_2265,N_2281);
nor U2478 (N_2478,N_2299,N_2130);
and U2479 (N_2479,N_2186,N_2267);
xor U2480 (N_2480,N_2318,N_2156);
and U2481 (N_2481,N_2154,N_2257);
nand U2482 (N_2482,N_2131,N_2236);
nand U2483 (N_2483,N_2105,N_2358);
xnor U2484 (N_2484,N_2279,N_2393);
or U2485 (N_2485,N_2103,N_2179);
xor U2486 (N_2486,N_2215,N_2128);
nor U2487 (N_2487,N_2382,N_2114);
and U2488 (N_2488,N_2194,N_2252);
nor U2489 (N_2489,N_2167,N_2176);
or U2490 (N_2490,N_2145,N_2274);
nand U2491 (N_2491,N_2313,N_2260);
or U2492 (N_2492,N_2206,N_2232);
or U2493 (N_2493,N_2177,N_2288);
nand U2494 (N_2494,N_2349,N_2353);
or U2495 (N_2495,N_2383,N_2305);
and U2496 (N_2496,N_2135,N_2261);
nand U2497 (N_2497,N_2210,N_2387);
nand U2498 (N_2498,N_2310,N_2373);
nand U2499 (N_2499,N_2123,N_2375);
and U2500 (N_2500,N_2368,N_2365);
nand U2501 (N_2501,N_2163,N_2329);
nor U2502 (N_2502,N_2113,N_2351);
and U2503 (N_2503,N_2235,N_2241);
nand U2504 (N_2504,N_2304,N_2343);
or U2505 (N_2505,N_2337,N_2225);
nand U2506 (N_2506,N_2189,N_2340);
nand U2507 (N_2507,N_2256,N_2228);
or U2508 (N_2508,N_2284,N_2233);
nand U2509 (N_2509,N_2188,N_2175);
or U2510 (N_2510,N_2361,N_2147);
nor U2511 (N_2511,N_2291,N_2345);
xor U2512 (N_2512,N_2141,N_2321);
and U2513 (N_2513,N_2227,N_2307);
or U2514 (N_2514,N_2335,N_2203);
or U2515 (N_2515,N_2136,N_2184);
or U2516 (N_2516,N_2327,N_2271);
and U2517 (N_2517,N_2183,N_2119);
nor U2518 (N_2518,N_2190,N_2269);
and U2519 (N_2519,N_2218,N_2166);
and U2520 (N_2520,N_2302,N_2222);
nor U2521 (N_2521,N_2198,N_2221);
xor U2522 (N_2522,N_2149,N_2226);
xnor U2523 (N_2523,N_2238,N_2100);
nand U2524 (N_2524,N_2132,N_2263);
nand U2525 (N_2525,N_2292,N_2370);
nand U2526 (N_2526,N_2134,N_2245);
xnor U2527 (N_2527,N_2150,N_2158);
xor U2528 (N_2528,N_2336,N_2331);
nand U2529 (N_2529,N_2231,N_2195);
or U2530 (N_2530,N_2346,N_2178);
or U2531 (N_2531,N_2392,N_2320);
xnor U2532 (N_2532,N_2137,N_2220);
and U2533 (N_2533,N_2356,N_2272);
nand U2534 (N_2534,N_2380,N_2295);
nor U2535 (N_2535,N_2234,N_2322);
nand U2536 (N_2536,N_2180,N_2379);
nor U2537 (N_2537,N_2350,N_2378);
and U2538 (N_2538,N_2219,N_2106);
or U2539 (N_2539,N_2297,N_2266);
or U2540 (N_2540,N_2160,N_2303);
nand U2541 (N_2541,N_2155,N_2399);
or U2542 (N_2542,N_2397,N_2273);
and U2543 (N_2543,N_2289,N_2162);
xnor U2544 (N_2544,N_2312,N_2109);
nor U2545 (N_2545,N_2367,N_2298);
nor U2546 (N_2546,N_2146,N_2359);
and U2547 (N_2547,N_2363,N_2140);
xnor U2548 (N_2548,N_2185,N_2159);
and U2549 (N_2549,N_2388,N_2282);
nor U2550 (N_2550,N_2122,N_2334);
nor U2551 (N_2551,N_2208,N_2185);
nor U2552 (N_2552,N_2272,N_2289);
and U2553 (N_2553,N_2328,N_2260);
xor U2554 (N_2554,N_2313,N_2323);
xnor U2555 (N_2555,N_2260,N_2155);
or U2556 (N_2556,N_2367,N_2379);
or U2557 (N_2557,N_2236,N_2161);
or U2558 (N_2558,N_2151,N_2384);
and U2559 (N_2559,N_2324,N_2229);
xnor U2560 (N_2560,N_2334,N_2220);
and U2561 (N_2561,N_2171,N_2353);
or U2562 (N_2562,N_2164,N_2241);
xor U2563 (N_2563,N_2261,N_2199);
or U2564 (N_2564,N_2175,N_2369);
nor U2565 (N_2565,N_2181,N_2188);
nand U2566 (N_2566,N_2166,N_2122);
xnor U2567 (N_2567,N_2210,N_2394);
or U2568 (N_2568,N_2194,N_2383);
and U2569 (N_2569,N_2282,N_2369);
or U2570 (N_2570,N_2360,N_2174);
and U2571 (N_2571,N_2345,N_2397);
or U2572 (N_2572,N_2219,N_2324);
and U2573 (N_2573,N_2130,N_2208);
nor U2574 (N_2574,N_2392,N_2276);
nand U2575 (N_2575,N_2179,N_2119);
and U2576 (N_2576,N_2237,N_2190);
and U2577 (N_2577,N_2325,N_2294);
and U2578 (N_2578,N_2147,N_2119);
and U2579 (N_2579,N_2302,N_2109);
xor U2580 (N_2580,N_2189,N_2247);
and U2581 (N_2581,N_2334,N_2369);
xor U2582 (N_2582,N_2267,N_2222);
xor U2583 (N_2583,N_2159,N_2271);
or U2584 (N_2584,N_2343,N_2371);
xnor U2585 (N_2585,N_2390,N_2289);
or U2586 (N_2586,N_2366,N_2321);
nand U2587 (N_2587,N_2256,N_2377);
or U2588 (N_2588,N_2283,N_2144);
or U2589 (N_2589,N_2246,N_2190);
or U2590 (N_2590,N_2256,N_2169);
nand U2591 (N_2591,N_2345,N_2248);
and U2592 (N_2592,N_2245,N_2258);
nor U2593 (N_2593,N_2337,N_2385);
and U2594 (N_2594,N_2396,N_2189);
nand U2595 (N_2595,N_2223,N_2244);
xnor U2596 (N_2596,N_2263,N_2126);
xor U2597 (N_2597,N_2206,N_2342);
or U2598 (N_2598,N_2152,N_2119);
nor U2599 (N_2599,N_2379,N_2318);
nor U2600 (N_2600,N_2312,N_2263);
nand U2601 (N_2601,N_2393,N_2352);
and U2602 (N_2602,N_2227,N_2192);
and U2603 (N_2603,N_2148,N_2321);
nor U2604 (N_2604,N_2353,N_2294);
nand U2605 (N_2605,N_2249,N_2271);
and U2606 (N_2606,N_2219,N_2113);
nor U2607 (N_2607,N_2342,N_2289);
or U2608 (N_2608,N_2335,N_2260);
and U2609 (N_2609,N_2331,N_2159);
nand U2610 (N_2610,N_2199,N_2319);
or U2611 (N_2611,N_2199,N_2247);
or U2612 (N_2612,N_2158,N_2338);
nand U2613 (N_2613,N_2159,N_2274);
or U2614 (N_2614,N_2302,N_2304);
xnor U2615 (N_2615,N_2360,N_2285);
nor U2616 (N_2616,N_2393,N_2320);
xnor U2617 (N_2617,N_2354,N_2345);
and U2618 (N_2618,N_2379,N_2279);
nor U2619 (N_2619,N_2259,N_2174);
nor U2620 (N_2620,N_2311,N_2338);
or U2621 (N_2621,N_2237,N_2220);
nand U2622 (N_2622,N_2355,N_2124);
and U2623 (N_2623,N_2175,N_2332);
nand U2624 (N_2624,N_2118,N_2203);
and U2625 (N_2625,N_2138,N_2364);
nand U2626 (N_2626,N_2137,N_2158);
nor U2627 (N_2627,N_2284,N_2243);
nor U2628 (N_2628,N_2232,N_2306);
or U2629 (N_2629,N_2277,N_2325);
nor U2630 (N_2630,N_2176,N_2130);
and U2631 (N_2631,N_2370,N_2118);
nand U2632 (N_2632,N_2351,N_2329);
and U2633 (N_2633,N_2372,N_2154);
xor U2634 (N_2634,N_2117,N_2397);
or U2635 (N_2635,N_2306,N_2139);
or U2636 (N_2636,N_2293,N_2130);
or U2637 (N_2637,N_2326,N_2374);
nor U2638 (N_2638,N_2375,N_2109);
nand U2639 (N_2639,N_2348,N_2227);
and U2640 (N_2640,N_2364,N_2115);
and U2641 (N_2641,N_2295,N_2374);
and U2642 (N_2642,N_2110,N_2155);
nand U2643 (N_2643,N_2293,N_2290);
xnor U2644 (N_2644,N_2243,N_2328);
nor U2645 (N_2645,N_2197,N_2297);
xor U2646 (N_2646,N_2345,N_2210);
nor U2647 (N_2647,N_2322,N_2238);
or U2648 (N_2648,N_2227,N_2309);
and U2649 (N_2649,N_2216,N_2110);
or U2650 (N_2650,N_2161,N_2353);
xor U2651 (N_2651,N_2364,N_2329);
nand U2652 (N_2652,N_2220,N_2390);
nand U2653 (N_2653,N_2196,N_2143);
xor U2654 (N_2654,N_2298,N_2120);
or U2655 (N_2655,N_2112,N_2229);
nor U2656 (N_2656,N_2267,N_2210);
xor U2657 (N_2657,N_2367,N_2251);
nor U2658 (N_2658,N_2301,N_2256);
nor U2659 (N_2659,N_2329,N_2326);
nor U2660 (N_2660,N_2290,N_2213);
and U2661 (N_2661,N_2372,N_2187);
nand U2662 (N_2662,N_2394,N_2368);
or U2663 (N_2663,N_2156,N_2334);
and U2664 (N_2664,N_2157,N_2286);
nand U2665 (N_2665,N_2182,N_2175);
nand U2666 (N_2666,N_2147,N_2213);
nor U2667 (N_2667,N_2397,N_2286);
or U2668 (N_2668,N_2120,N_2116);
nand U2669 (N_2669,N_2287,N_2336);
and U2670 (N_2670,N_2381,N_2196);
or U2671 (N_2671,N_2321,N_2198);
xnor U2672 (N_2672,N_2281,N_2345);
and U2673 (N_2673,N_2277,N_2131);
and U2674 (N_2674,N_2201,N_2226);
nand U2675 (N_2675,N_2146,N_2297);
xor U2676 (N_2676,N_2366,N_2368);
and U2677 (N_2677,N_2250,N_2152);
or U2678 (N_2678,N_2231,N_2184);
xnor U2679 (N_2679,N_2379,N_2142);
nand U2680 (N_2680,N_2350,N_2364);
xor U2681 (N_2681,N_2217,N_2154);
xor U2682 (N_2682,N_2225,N_2343);
xor U2683 (N_2683,N_2265,N_2278);
xnor U2684 (N_2684,N_2303,N_2223);
or U2685 (N_2685,N_2317,N_2261);
xnor U2686 (N_2686,N_2109,N_2347);
nand U2687 (N_2687,N_2286,N_2185);
or U2688 (N_2688,N_2394,N_2346);
nor U2689 (N_2689,N_2183,N_2175);
and U2690 (N_2690,N_2183,N_2180);
nand U2691 (N_2691,N_2367,N_2164);
nor U2692 (N_2692,N_2271,N_2195);
or U2693 (N_2693,N_2371,N_2236);
nor U2694 (N_2694,N_2367,N_2235);
or U2695 (N_2695,N_2321,N_2231);
xor U2696 (N_2696,N_2194,N_2124);
and U2697 (N_2697,N_2353,N_2315);
xor U2698 (N_2698,N_2126,N_2261);
or U2699 (N_2699,N_2348,N_2339);
or U2700 (N_2700,N_2547,N_2423);
and U2701 (N_2701,N_2599,N_2511);
or U2702 (N_2702,N_2503,N_2415);
xor U2703 (N_2703,N_2455,N_2551);
nor U2704 (N_2704,N_2490,N_2431);
nor U2705 (N_2705,N_2563,N_2608);
or U2706 (N_2706,N_2546,N_2458);
nand U2707 (N_2707,N_2642,N_2521);
and U2708 (N_2708,N_2403,N_2532);
nand U2709 (N_2709,N_2435,N_2456);
or U2710 (N_2710,N_2537,N_2556);
or U2711 (N_2711,N_2595,N_2478);
and U2712 (N_2712,N_2497,N_2533);
nor U2713 (N_2713,N_2668,N_2679);
or U2714 (N_2714,N_2657,N_2651);
nand U2715 (N_2715,N_2680,N_2466);
xnor U2716 (N_2716,N_2512,N_2585);
and U2717 (N_2717,N_2422,N_2420);
xnor U2718 (N_2718,N_2436,N_2504);
nor U2719 (N_2719,N_2450,N_2622);
or U2720 (N_2720,N_2439,N_2550);
nand U2721 (N_2721,N_2640,N_2631);
nor U2722 (N_2722,N_2688,N_2535);
nand U2723 (N_2723,N_2624,N_2612);
and U2724 (N_2724,N_2582,N_2502);
and U2725 (N_2725,N_2566,N_2655);
xnor U2726 (N_2726,N_2685,N_2570);
nand U2727 (N_2727,N_2540,N_2643);
nand U2728 (N_2728,N_2462,N_2616);
and U2729 (N_2729,N_2492,N_2613);
and U2730 (N_2730,N_2488,N_2609);
nor U2731 (N_2731,N_2467,N_2638);
and U2732 (N_2732,N_2457,N_2611);
or U2733 (N_2733,N_2565,N_2667);
nand U2734 (N_2734,N_2578,N_2621);
or U2735 (N_2735,N_2670,N_2634);
xor U2736 (N_2736,N_2654,N_2418);
nand U2737 (N_2737,N_2548,N_2579);
and U2738 (N_2738,N_2482,N_2639);
nand U2739 (N_2739,N_2445,N_2587);
nand U2740 (N_2740,N_2693,N_2689);
and U2741 (N_2741,N_2493,N_2401);
and U2742 (N_2742,N_2427,N_2692);
or U2743 (N_2743,N_2553,N_2597);
xor U2744 (N_2744,N_2662,N_2414);
or U2745 (N_2745,N_2460,N_2614);
nand U2746 (N_2746,N_2416,N_2494);
or U2747 (N_2747,N_2652,N_2446);
and U2748 (N_2748,N_2541,N_2659);
nand U2749 (N_2749,N_2618,N_2602);
and U2750 (N_2750,N_2690,N_2538);
nand U2751 (N_2751,N_2687,N_2632);
and U2752 (N_2752,N_2684,N_2586);
and U2753 (N_2753,N_2525,N_2577);
nand U2754 (N_2754,N_2649,N_2426);
or U2755 (N_2755,N_2592,N_2646);
nor U2756 (N_2756,N_2672,N_2665);
nand U2757 (N_2757,N_2411,N_2477);
nor U2758 (N_2758,N_2628,N_2475);
nor U2759 (N_2759,N_2453,N_2417);
and U2760 (N_2760,N_2454,N_2437);
or U2761 (N_2761,N_2440,N_2678);
nand U2762 (N_2762,N_2552,N_2676);
or U2763 (N_2763,N_2469,N_2584);
nand U2764 (N_2764,N_2653,N_2580);
nand U2765 (N_2765,N_2451,N_2656);
nand U2766 (N_2766,N_2664,N_2574);
xor U2767 (N_2767,N_2523,N_2515);
nor U2768 (N_2768,N_2402,N_2575);
xnor U2769 (N_2769,N_2698,N_2645);
and U2770 (N_2770,N_2562,N_2471);
nand U2771 (N_2771,N_2675,N_2677);
nor U2772 (N_2772,N_2543,N_2428);
nor U2773 (N_2773,N_2476,N_2491);
nor U2774 (N_2774,N_2444,N_2573);
nand U2775 (N_2775,N_2473,N_2430);
nor U2776 (N_2776,N_2633,N_2530);
or U2777 (N_2777,N_2480,N_2669);
nor U2778 (N_2778,N_2560,N_2498);
nor U2779 (N_2779,N_2429,N_2516);
and U2780 (N_2780,N_2590,N_2410);
nor U2781 (N_2781,N_2527,N_2559);
xor U2782 (N_2782,N_2594,N_2518);
nor U2783 (N_2783,N_2620,N_2557);
nand U2784 (N_2784,N_2539,N_2526);
or U2785 (N_2785,N_2554,N_2536);
nand U2786 (N_2786,N_2641,N_2583);
xor U2787 (N_2787,N_2419,N_2408);
nand U2788 (N_2788,N_2528,N_2561);
xor U2789 (N_2789,N_2500,N_2404);
nand U2790 (N_2790,N_2581,N_2569);
xor U2791 (N_2791,N_2441,N_2406);
xor U2792 (N_2792,N_2671,N_2572);
and U2793 (N_2793,N_2697,N_2424);
or U2794 (N_2794,N_2483,N_2625);
xnor U2795 (N_2795,N_2448,N_2682);
nor U2796 (N_2796,N_2508,N_2470);
or U2797 (N_2797,N_2558,N_2650);
nor U2798 (N_2798,N_2647,N_2567);
or U2799 (N_2799,N_2610,N_2673);
and U2800 (N_2800,N_2501,N_2635);
and U2801 (N_2801,N_2630,N_2576);
nor U2802 (N_2802,N_2615,N_2617);
and U2803 (N_2803,N_2443,N_2555);
or U2804 (N_2804,N_2531,N_2637);
nand U2805 (N_2805,N_2449,N_2468);
xnor U2806 (N_2806,N_2513,N_2452);
and U2807 (N_2807,N_2607,N_2571);
or U2808 (N_2808,N_2568,N_2589);
nand U2809 (N_2809,N_2660,N_2564);
nand U2810 (N_2810,N_2699,N_2606);
xnor U2811 (N_2811,N_2604,N_2683);
xor U2812 (N_2812,N_2461,N_2434);
and U2813 (N_2813,N_2432,N_2534);
nand U2814 (N_2814,N_2619,N_2520);
xnor U2815 (N_2815,N_2524,N_2514);
or U2816 (N_2816,N_2433,N_2605);
and U2817 (N_2817,N_2472,N_2666);
xor U2818 (N_2818,N_2479,N_2484);
xor U2819 (N_2819,N_2627,N_2506);
or U2820 (N_2820,N_2438,N_2636);
nor U2821 (N_2821,N_2686,N_2623);
nand U2822 (N_2822,N_2691,N_2485);
nand U2823 (N_2823,N_2529,N_2405);
xor U2824 (N_2824,N_2412,N_2644);
or U2825 (N_2825,N_2495,N_2593);
or U2826 (N_2826,N_2681,N_2519);
nor U2827 (N_2827,N_2626,N_2409);
nor U2828 (N_2828,N_2601,N_2510);
nand U2829 (N_2829,N_2695,N_2596);
nor U2830 (N_2830,N_2499,N_2486);
nand U2831 (N_2831,N_2544,N_2603);
nand U2832 (N_2832,N_2507,N_2545);
or U2833 (N_2833,N_2694,N_2463);
and U2834 (N_2834,N_2522,N_2648);
or U2835 (N_2835,N_2487,N_2489);
nor U2836 (N_2836,N_2465,N_2658);
and U2837 (N_2837,N_2588,N_2549);
or U2838 (N_2838,N_2598,N_2509);
or U2839 (N_2839,N_2629,N_2400);
nor U2840 (N_2840,N_2542,N_2464);
and U2841 (N_2841,N_2474,N_2696);
nand U2842 (N_2842,N_2591,N_2481);
nor U2843 (N_2843,N_2661,N_2425);
nor U2844 (N_2844,N_2421,N_2459);
nor U2845 (N_2845,N_2600,N_2663);
nor U2846 (N_2846,N_2442,N_2674);
or U2847 (N_2847,N_2505,N_2407);
nand U2848 (N_2848,N_2496,N_2517);
xnor U2849 (N_2849,N_2447,N_2413);
nand U2850 (N_2850,N_2452,N_2566);
and U2851 (N_2851,N_2571,N_2509);
xnor U2852 (N_2852,N_2643,N_2541);
xor U2853 (N_2853,N_2607,N_2573);
nor U2854 (N_2854,N_2573,N_2425);
xnor U2855 (N_2855,N_2635,N_2664);
or U2856 (N_2856,N_2499,N_2684);
nor U2857 (N_2857,N_2690,N_2618);
nand U2858 (N_2858,N_2490,N_2500);
or U2859 (N_2859,N_2601,N_2676);
nor U2860 (N_2860,N_2560,N_2586);
and U2861 (N_2861,N_2455,N_2434);
and U2862 (N_2862,N_2563,N_2690);
xor U2863 (N_2863,N_2696,N_2475);
nand U2864 (N_2864,N_2436,N_2505);
xnor U2865 (N_2865,N_2644,N_2433);
or U2866 (N_2866,N_2683,N_2430);
nand U2867 (N_2867,N_2402,N_2669);
or U2868 (N_2868,N_2674,N_2548);
and U2869 (N_2869,N_2586,N_2434);
or U2870 (N_2870,N_2591,N_2625);
and U2871 (N_2871,N_2480,N_2659);
and U2872 (N_2872,N_2541,N_2596);
or U2873 (N_2873,N_2605,N_2635);
or U2874 (N_2874,N_2647,N_2486);
xnor U2875 (N_2875,N_2523,N_2541);
xnor U2876 (N_2876,N_2627,N_2541);
nand U2877 (N_2877,N_2404,N_2582);
and U2878 (N_2878,N_2417,N_2612);
or U2879 (N_2879,N_2610,N_2552);
nor U2880 (N_2880,N_2462,N_2619);
and U2881 (N_2881,N_2483,N_2683);
and U2882 (N_2882,N_2497,N_2441);
xor U2883 (N_2883,N_2445,N_2696);
and U2884 (N_2884,N_2412,N_2598);
or U2885 (N_2885,N_2541,N_2537);
nand U2886 (N_2886,N_2508,N_2532);
nand U2887 (N_2887,N_2677,N_2680);
nand U2888 (N_2888,N_2616,N_2458);
nand U2889 (N_2889,N_2650,N_2546);
nand U2890 (N_2890,N_2486,N_2654);
xor U2891 (N_2891,N_2472,N_2561);
xor U2892 (N_2892,N_2669,N_2693);
nor U2893 (N_2893,N_2622,N_2413);
nand U2894 (N_2894,N_2694,N_2516);
nor U2895 (N_2895,N_2674,N_2668);
or U2896 (N_2896,N_2607,N_2484);
or U2897 (N_2897,N_2481,N_2574);
nand U2898 (N_2898,N_2514,N_2579);
nor U2899 (N_2899,N_2645,N_2676);
or U2900 (N_2900,N_2542,N_2661);
or U2901 (N_2901,N_2471,N_2547);
or U2902 (N_2902,N_2581,N_2535);
or U2903 (N_2903,N_2671,N_2660);
xnor U2904 (N_2904,N_2666,N_2676);
xor U2905 (N_2905,N_2616,N_2488);
xnor U2906 (N_2906,N_2539,N_2422);
nand U2907 (N_2907,N_2689,N_2556);
xor U2908 (N_2908,N_2414,N_2458);
nand U2909 (N_2909,N_2679,N_2491);
nand U2910 (N_2910,N_2672,N_2433);
xnor U2911 (N_2911,N_2663,N_2690);
xnor U2912 (N_2912,N_2414,N_2601);
nand U2913 (N_2913,N_2426,N_2632);
and U2914 (N_2914,N_2567,N_2595);
and U2915 (N_2915,N_2482,N_2573);
and U2916 (N_2916,N_2435,N_2634);
xor U2917 (N_2917,N_2494,N_2612);
or U2918 (N_2918,N_2516,N_2620);
nor U2919 (N_2919,N_2521,N_2474);
and U2920 (N_2920,N_2618,N_2476);
xor U2921 (N_2921,N_2480,N_2414);
nand U2922 (N_2922,N_2611,N_2449);
nor U2923 (N_2923,N_2409,N_2466);
nand U2924 (N_2924,N_2444,N_2440);
nor U2925 (N_2925,N_2575,N_2578);
nand U2926 (N_2926,N_2460,N_2608);
nand U2927 (N_2927,N_2500,N_2401);
xnor U2928 (N_2928,N_2471,N_2464);
and U2929 (N_2929,N_2563,N_2656);
or U2930 (N_2930,N_2419,N_2452);
and U2931 (N_2931,N_2637,N_2677);
xor U2932 (N_2932,N_2613,N_2669);
and U2933 (N_2933,N_2445,N_2457);
xor U2934 (N_2934,N_2643,N_2697);
nand U2935 (N_2935,N_2546,N_2678);
and U2936 (N_2936,N_2691,N_2461);
or U2937 (N_2937,N_2507,N_2484);
xnor U2938 (N_2938,N_2566,N_2632);
nand U2939 (N_2939,N_2588,N_2511);
and U2940 (N_2940,N_2570,N_2630);
nand U2941 (N_2941,N_2474,N_2593);
nor U2942 (N_2942,N_2576,N_2502);
xnor U2943 (N_2943,N_2424,N_2692);
nand U2944 (N_2944,N_2471,N_2479);
and U2945 (N_2945,N_2581,N_2401);
and U2946 (N_2946,N_2457,N_2651);
nor U2947 (N_2947,N_2618,N_2550);
xnor U2948 (N_2948,N_2553,N_2554);
nor U2949 (N_2949,N_2607,N_2604);
nand U2950 (N_2950,N_2463,N_2588);
nor U2951 (N_2951,N_2610,N_2575);
nand U2952 (N_2952,N_2422,N_2496);
nor U2953 (N_2953,N_2551,N_2558);
nor U2954 (N_2954,N_2567,N_2531);
nor U2955 (N_2955,N_2550,N_2608);
xnor U2956 (N_2956,N_2572,N_2563);
or U2957 (N_2957,N_2489,N_2560);
xor U2958 (N_2958,N_2669,N_2680);
nor U2959 (N_2959,N_2619,N_2552);
and U2960 (N_2960,N_2593,N_2411);
or U2961 (N_2961,N_2428,N_2657);
and U2962 (N_2962,N_2493,N_2464);
nor U2963 (N_2963,N_2691,N_2483);
or U2964 (N_2964,N_2598,N_2424);
nand U2965 (N_2965,N_2412,N_2415);
nand U2966 (N_2966,N_2578,N_2611);
xnor U2967 (N_2967,N_2548,N_2552);
nor U2968 (N_2968,N_2469,N_2493);
xnor U2969 (N_2969,N_2423,N_2544);
xor U2970 (N_2970,N_2468,N_2672);
nand U2971 (N_2971,N_2553,N_2664);
nand U2972 (N_2972,N_2438,N_2642);
nand U2973 (N_2973,N_2584,N_2450);
nand U2974 (N_2974,N_2556,N_2664);
and U2975 (N_2975,N_2619,N_2447);
nor U2976 (N_2976,N_2480,N_2655);
or U2977 (N_2977,N_2560,N_2644);
nor U2978 (N_2978,N_2517,N_2514);
nor U2979 (N_2979,N_2610,N_2661);
and U2980 (N_2980,N_2596,N_2647);
or U2981 (N_2981,N_2485,N_2539);
nor U2982 (N_2982,N_2602,N_2660);
nor U2983 (N_2983,N_2520,N_2688);
nand U2984 (N_2984,N_2590,N_2572);
nand U2985 (N_2985,N_2676,N_2491);
nand U2986 (N_2986,N_2525,N_2444);
or U2987 (N_2987,N_2443,N_2421);
nand U2988 (N_2988,N_2639,N_2684);
and U2989 (N_2989,N_2593,N_2562);
or U2990 (N_2990,N_2472,N_2627);
or U2991 (N_2991,N_2621,N_2566);
xor U2992 (N_2992,N_2615,N_2690);
xnor U2993 (N_2993,N_2438,N_2472);
xor U2994 (N_2994,N_2684,N_2561);
nor U2995 (N_2995,N_2567,N_2683);
or U2996 (N_2996,N_2443,N_2452);
nor U2997 (N_2997,N_2417,N_2462);
nor U2998 (N_2998,N_2623,N_2613);
or U2999 (N_2999,N_2517,N_2560);
xnor U3000 (N_3000,N_2819,N_2789);
or U3001 (N_3001,N_2749,N_2797);
or U3002 (N_3002,N_2932,N_2814);
nor U3003 (N_3003,N_2760,N_2981);
or U3004 (N_3004,N_2842,N_2708);
nand U3005 (N_3005,N_2852,N_2897);
and U3006 (N_3006,N_2765,N_2731);
nand U3007 (N_3007,N_2737,N_2905);
or U3008 (N_3008,N_2886,N_2702);
nand U3009 (N_3009,N_2748,N_2803);
nand U3010 (N_3010,N_2945,N_2917);
or U3011 (N_3011,N_2841,N_2959);
or U3012 (N_3012,N_2856,N_2986);
xor U3013 (N_3013,N_2700,N_2937);
or U3014 (N_3014,N_2824,N_2881);
or U3015 (N_3015,N_2723,N_2785);
xor U3016 (N_3016,N_2781,N_2880);
nand U3017 (N_3017,N_2736,N_2719);
or U3018 (N_3018,N_2929,N_2858);
xor U3019 (N_3019,N_2851,N_2954);
nor U3020 (N_3020,N_2712,N_2786);
and U3021 (N_3021,N_2701,N_2909);
nand U3022 (N_3022,N_2919,N_2924);
xor U3023 (N_3023,N_2928,N_2831);
or U3024 (N_3024,N_2949,N_2808);
nor U3025 (N_3025,N_2714,N_2792);
nand U3026 (N_3026,N_2735,N_2835);
or U3027 (N_3027,N_2816,N_2796);
nor U3028 (N_3028,N_2873,N_2862);
nand U3029 (N_3029,N_2742,N_2982);
nor U3030 (N_3030,N_2899,N_2952);
nor U3031 (N_3031,N_2948,N_2745);
nand U3032 (N_3032,N_2746,N_2703);
xor U3033 (N_3033,N_2992,N_2989);
nor U3034 (N_3034,N_2947,N_2974);
xor U3035 (N_3035,N_2894,N_2713);
or U3036 (N_3036,N_2990,N_2844);
nand U3037 (N_3037,N_2732,N_2978);
xor U3038 (N_3038,N_2729,N_2747);
nand U3039 (N_3039,N_2788,N_2941);
or U3040 (N_3040,N_2846,N_2991);
nand U3041 (N_3041,N_2942,N_2925);
xnor U3042 (N_3042,N_2743,N_2825);
nand U3043 (N_3043,N_2717,N_2812);
and U3044 (N_3044,N_2798,N_2836);
nand U3045 (N_3045,N_2854,N_2775);
and U3046 (N_3046,N_2969,N_2870);
or U3047 (N_3047,N_2810,N_2716);
nand U3048 (N_3048,N_2984,N_2995);
and U3049 (N_3049,N_2802,N_2906);
or U3050 (N_3050,N_2787,N_2916);
nor U3051 (N_3051,N_2751,N_2908);
nand U3052 (N_3052,N_2963,N_2939);
xnor U3053 (N_3053,N_2800,N_2815);
and U3054 (N_3054,N_2869,N_2965);
and U3055 (N_3055,N_2931,N_2892);
and U3056 (N_3056,N_2875,N_2795);
nor U3057 (N_3057,N_2759,N_2985);
and U3058 (N_3058,N_2706,N_2843);
nor U3059 (N_3059,N_2915,N_2935);
nor U3060 (N_3060,N_2857,N_2801);
or U3061 (N_3061,N_2956,N_2754);
nand U3062 (N_3062,N_2890,N_2794);
xor U3063 (N_3063,N_2987,N_2888);
and U3064 (N_3064,N_2711,N_2829);
nand U3065 (N_3065,N_2896,N_2864);
nor U3066 (N_3066,N_2849,N_2780);
xnor U3067 (N_3067,N_2720,N_2715);
and U3068 (N_3068,N_2766,N_2763);
nand U3069 (N_3069,N_2980,N_2821);
nand U3070 (N_3070,N_2926,N_2927);
xor U3071 (N_3071,N_2868,N_2828);
or U3072 (N_3072,N_2953,N_2764);
nor U3073 (N_3073,N_2898,N_2839);
and U3074 (N_3074,N_2818,N_2960);
nand U3075 (N_3075,N_2883,N_2838);
nor U3076 (N_3076,N_2921,N_2877);
nand U3077 (N_3077,N_2940,N_2772);
xnor U3078 (N_3078,N_2866,N_2867);
and U3079 (N_3079,N_2734,N_2721);
nand U3080 (N_3080,N_2855,N_2791);
nor U3081 (N_3081,N_2770,N_2961);
nand U3082 (N_3082,N_2777,N_2914);
nor U3083 (N_3083,N_2827,N_2790);
and U3084 (N_3084,N_2972,N_2901);
xnor U3085 (N_3085,N_2865,N_2776);
nor U3086 (N_3086,N_2799,N_2891);
and U3087 (N_3087,N_2761,N_2994);
nand U3088 (N_3088,N_2957,N_2755);
nor U3089 (N_3089,N_2837,N_2912);
and U3090 (N_3090,N_2861,N_2977);
nor U3091 (N_3091,N_2840,N_2728);
xor U3092 (N_3092,N_2903,N_2975);
nand U3093 (N_3093,N_2725,N_2740);
and U3094 (N_3094,N_2750,N_2923);
nand U3095 (N_3095,N_2834,N_2902);
xnor U3096 (N_3096,N_2756,N_2758);
nand U3097 (N_3097,N_2704,N_2907);
nand U3098 (N_3098,N_2934,N_2885);
xor U3099 (N_3099,N_2806,N_2900);
xnor U3100 (N_3100,N_2832,N_2913);
nor U3101 (N_3101,N_2733,N_2904);
and U3102 (N_3102,N_2762,N_2946);
or U3103 (N_3103,N_2833,N_2850);
xor U3104 (N_3104,N_2860,N_2933);
nor U3105 (N_3105,N_2738,N_2709);
and U3106 (N_3106,N_2782,N_2805);
and U3107 (N_3107,N_2893,N_2936);
nand U3108 (N_3108,N_2938,N_2970);
and U3109 (N_3109,N_2853,N_2830);
xnor U3110 (N_3110,N_2967,N_2922);
or U3111 (N_3111,N_2918,N_2848);
or U3112 (N_3112,N_2889,N_2774);
nor U3113 (N_3113,N_2813,N_2878);
nor U3114 (N_3114,N_2847,N_2811);
nand U3115 (N_3115,N_2988,N_2882);
and U3116 (N_3116,N_2778,N_2817);
nand U3117 (N_3117,N_2920,N_2710);
or U3118 (N_3118,N_2726,N_2845);
nand U3119 (N_3119,N_2718,N_2999);
nor U3120 (N_3120,N_2753,N_2996);
or U3121 (N_3121,N_2730,N_2971);
or U3122 (N_3122,N_2752,N_2783);
nor U3123 (N_3123,N_2943,N_2784);
nor U3124 (N_3124,N_2822,N_2998);
nor U3125 (N_3125,N_2884,N_2872);
and U3126 (N_3126,N_2807,N_2958);
and U3127 (N_3127,N_2859,N_2979);
and U3128 (N_3128,N_2769,N_2722);
nor U3129 (N_3129,N_2950,N_2962);
nor U3130 (N_3130,N_2951,N_2879);
nand U3131 (N_3131,N_2911,N_2826);
xnor U3132 (N_3132,N_2993,N_2895);
or U3133 (N_3133,N_2809,N_2757);
and U3134 (N_3134,N_2768,N_2705);
nor U3135 (N_3135,N_2727,N_2887);
nor U3136 (N_3136,N_2741,N_2773);
nor U3137 (N_3137,N_2707,N_2997);
xor U3138 (N_3138,N_2964,N_2983);
or U3139 (N_3139,N_2820,N_2966);
nand U3140 (N_3140,N_2724,N_2804);
nand U3141 (N_3141,N_2744,N_2968);
and U3142 (N_3142,N_2767,N_2823);
xor U3143 (N_3143,N_2876,N_2874);
nor U3144 (N_3144,N_2779,N_2973);
nand U3145 (N_3145,N_2976,N_2739);
and U3146 (N_3146,N_2871,N_2771);
or U3147 (N_3147,N_2944,N_2910);
nand U3148 (N_3148,N_2793,N_2930);
and U3149 (N_3149,N_2863,N_2955);
and U3150 (N_3150,N_2712,N_2784);
nor U3151 (N_3151,N_2847,N_2713);
nor U3152 (N_3152,N_2992,N_2819);
or U3153 (N_3153,N_2875,N_2742);
nand U3154 (N_3154,N_2876,N_2806);
xor U3155 (N_3155,N_2798,N_2906);
xnor U3156 (N_3156,N_2826,N_2982);
nor U3157 (N_3157,N_2818,N_2880);
nor U3158 (N_3158,N_2790,N_2993);
nor U3159 (N_3159,N_2917,N_2821);
or U3160 (N_3160,N_2710,N_2834);
nor U3161 (N_3161,N_2942,N_2901);
nor U3162 (N_3162,N_2724,N_2955);
and U3163 (N_3163,N_2911,N_2852);
and U3164 (N_3164,N_2757,N_2797);
xnor U3165 (N_3165,N_2958,N_2865);
nand U3166 (N_3166,N_2989,N_2933);
xor U3167 (N_3167,N_2985,N_2791);
xnor U3168 (N_3168,N_2980,N_2764);
nor U3169 (N_3169,N_2825,N_2832);
and U3170 (N_3170,N_2872,N_2866);
and U3171 (N_3171,N_2810,N_2719);
and U3172 (N_3172,N_2858,N_2874);
nor U3173 (N_3173,N_2757,N_2791);
and U3174 (N_3174,N_2859,N_2872);
xor U3175 (N_3175,N_2949,N_2857);
and U3176 (N_3176,N_2914,N_2712);
and U3177 (N_3177,N_2780,N_2706);
nand U3178 (N_3178,N_2858,N_2992);
nand U3179 (N_3179,N_2872,N_2927);
xnor U3180 (N_3180,N_2807,N_2765);
or U3181 (N_3181,N_2840,N_2763);
or U3182 (N_3182,N_2788,N_2936);
nand U3183 (N_3183,N_2708,N_2974);
nand U3184 (N_3184,N_2886,N_2723);
xnor U3185 (N_3185,N_2997,N_2867);
or U3186 (N_3186,N_2852,N_2869);
xor U3187 (N_3187,N_2838,N_2744);
xnor U3188 (N_3188,N_2935,N_2840);
or U3189 (N_3189,N_2776,N_2825);
or U3190 (N_3190,N_2991,N_2750);
xor U3191 (N_3191,N_2923,N_2898);
xnor U3192 (N_3192,N_2992,N_2902);
nand U3193 (N_3193,N_2948,N_2819);
or U3194 (N_3194,N_2987,N_2778);
xnor U3195 (N_3195,N_2848,N_2866);
and U3196 (N_3196,N_2833,N_2743);
or U3197 (N_3197,N_2925,N_2829);
nor U3198 (N_3198,N_2989,N_2925);
or U3199 (N_3199,N_2806,N_2820);
nor U3200 (N_3200,N_2841,N_2971);
nor U3201 (N_3201,N_2730,N_2992);
and U3202 (N_3202,N_2950,N_2763);
nand U3203 (N_3203,N_2834,N_2813);
and U3204 (N_3204,N_2976,N_2918);
nor U3205 (N_3205,N_2772,N_2808);
or U3206 (N_3206,N_2805,N_2775);
nand U3207 (N_3207,N_2775,N_2733);
nor U3208 (N_3208,N_2987,N_2978);
nor U3209 (N_3209,N_2704,N_2817);
or U3210 (N_3210,N_2733,N_2752);
nand U3211 (N_3211,N_2837,N_2727);
and U3212 (N_3212,N_2971,N_2831);
and U3213 (N_3213,N_2763,N_2910);
nand U3214 (N_3214,N_2937,N_2852);
xnor U3215 (N_3215,N_2848,N_2747);
or U3216 (N_3216,N_2847,N_2941);
nor U3217 (N_3217,N_2765,N_2903);
nand U3218 (N_3218,N_2859,N_2853);
xor U3219 (N_3219,N_2869,N_2885);
or U3220 (N_3220,N_2793,N_2733);
and U3221 (N_3221,N_2893,N_2709);
xnor U3222 (N_3222,N_2724,N_2877);
nand U3223 (N_3223,N_2806,N_2849);
nor U3224 (N_3224,N_2768,N_2987);
nand U3225 (N_3225,N_2719,N_2955);
nor U3226 (N_3226,N_2968,N_2990);
nand U3227 (N_3227,N_2923,N_2782);
and U3228 (N_3228,N_2923,N_2947);
xor U3229 (N_3229,N_2821,N_2929);
or U3230 (N_3230,N_2816,N_2916);
nand U3231 (N_3231,N_2995,N_2870);
or U3232 (N_3232,N_2718,N_2821);
nand U3233 (N_3233,N_2727,N_2854);
or U3234 (N_3234,N_2718,N_2883);
nor U3235 (N_3235,N_2953,N_2708);
xor U3236 (N_3236,N_2986,N_2940);
or U3237 (N_3237,N_2809,N_2769);
or U3238 (N_3238,N_2777,N_2994);
or U3239 (N_3239,N_2716,N_2962);
and U3240 (N_3240,N_2992,N_2744);
nor U3241 (N_3241,N_2987,N_2968);
nand U3242 (N_3242,N_2905,N_2741);
and U3243 (N_3243,N_2862,N_2876);
nor U3244 (N_3244,N_2918,N_2795);
and U3245 (N_3245,N_2977,N_2943);
xor U3246 (N_3246,N_2818,N_2840);
or U3247 (N_3247,N_2986,N_2907);
nand U3248 (N_3248,N_2746,N_2854);
nor U3249 (N_3249,N_2836,N_2856);
nor U3250 (N_3250,N_2753,N_2884);
and U3251 (N_3251,N_2908,N_2849);
nor U3252 (N_3252,N_2815,N_2740);
or U3253 (N_3253,N_2745,N_2753);
nor U3254 (N_3254,N_2841,N_2850);
xor U3255 (N_3255,N_2743,N_2797);
xor U3256 (N_3256,N_2812,N_2870);
nand U3257 (N_3257,N_2715,N_2752);
nand U3258 (N_3258,N_2853,N_2847);
xnor U3259 (N_3259,N_2710,N_2981);
or U3260 (N_3260,N_2705,N_2872);
nor U3261 (N_3261,N_2816,N_2872);
xor U3262 (N_3262,N_2962,N_2705);
or U3263 (N_3263,N_2890,N_2915);
or U3264 (N_3264,N_2891,N_2930);
nor U3265 (N_3265,N_2938,N_2823);
xor U3266 (N_3266,N_2808,N_2797);
and U3267 (N_3267,N_2806,N_2807);
and U3268 (N_3268,N_2745,N_2904);
xor U3269 (N_3269,N_2845,N_2980);
xnor U3270 (N_3270,N_2758,N_2735);
nand U3271 (N_3271,N_2949,N_2852);
nor U3272 (N_3272,N_2837,N_2813);
nand U3273 (N_3273,N_2721,N_2791);
xor U3274 (N_3274,N_2735,N_2834);
and U3275 (N_3275,N_2743,N_2706);
or U3276 (N_3276,N_2753,N_2768);
xor U3277 (N_3277,N_2707,N_2948);
nand U3278 (N_3278,N_2979,N_2707);
or U3279 (N_3279,N_2960,N_2824);
or U3280 (N_3280,N_2902,N_2751);
or U3281 (N_3281,N_2984,N_2706);
and U3282 (N_3282,N_2790,N_2976);
nor U3283 (N_3283,N_2756,N_2987);
xor U3284 (N_3284,N_2737,N_2839);
nand U3285 (N_3285,N_2703,N_2800);
xnor U3286 (N_3286,N_2821,N_2892);
nor U3287 (N_3287,N_2806,N_2797);
or U3288 (N_3288,N_2773,N_2940);
nand U3289 (N_3289,N_2730,N_2732);
and U3290 (N_3290,N_2971,N_2733);
or U3291 (N_3291,N_2988,N_2851);
xor U3292 (N_3292,N_2916,N_2705);
nor U3293 (N_3293,N_2723,N_2889);
or U3294 (N_3294,N_2739,N_2857);
nor U3295 (N_3295,N_2946,N_2882);
nor U3296 (N_3296,N_2986,N_2830);
nor U3297 (N_3297,N_2842,N_2870);
xnor U3298 (N_3298,N_2989,N_2803);
xnor U3299 (N_3299,N_2821,N_2780);
and U3300 (N_3300,N_3270,N_3205);
xor U3301 (N_3301,N_3024,N_3218);
nor U3302 (N_3302,N_3103,N_3107);
nor U3303 (N_3303,N_3058,N_3274);
nor U3304 (N_3304,N_3296,N_3215);
nand U3305 (N_3305,N_3233,N_3166);
xnor U3306 (N_3306,N_3179,N_3172);
nand U3307 (N_3307,N_3036,N_3294);
nand U3308 (N_3308,N_3008,N_3245);
or U3309 (N_3309,N_3134,N_3113);
xnor U3310 (N_3310,N_3141,N_3148);
nand U3311 (N_3311,N_3127,N_3212);
and U3312 (N_3312,N_3007,N_3120);
nand U3313 (N_3313,N_3189,N_3226);
xor U3314 (N_3314,N_3262,N_3059);
xnor U3315 (N_3315,N_3298,N_3152);
and U3316 (N_3316,N_3019,N_3197);
or U3317 (N_3317,N_3288,N_3228);
and U3318 (N_3318,N_3185,N_3266);
nor U3319 (N_3319,N_3225,N_3170);
nor U3320 (N_3320,N_3022,N_3214);
and U3321 (N_3321,N_3249,N_3081);
and U3322 (N_3322,N_3279,N_3039);
xor U3323 (N_3323,N_3167,N_3133);
or U3324 (N_3324,N_3153,N_3235);
nor U3325 (N_3325,N_3063,N_3162);
or U3326 (N_3326,N_3043,N_3032);
xor U3327 (N_3327,N_3010,N_3090);
xor U3328 (N_3328,N_3201,N_3042);
nor U3329 (N_3329,N_3251,N_3057);
nor U3330 (N_3330,N_3267,N_3048);
xor U3331 (N_3331,N_3031,N_3020);
or U3332 (N_3332,N_3281,N_3100);
nand U3333 (N_3333,N_3102,N_3015);
or U3334 (N_3334,N_3291,N_3142);
and U3335 (N_3335,N_3150,N_3250);
xnor U3336 (N_3336,N_3154,N_3068);
nor U3337 (N_3337,N_3222,N_3053);
nand U3338 (N_3338,N_3180,N_3181);
and U3339 (N_3339,N_3295,N_3175);
nand U3340 (N_3340,N_3091,N_3040);
or U3341 (N_3341,N_3144,N_3160);
nor U3342 (N_3342,N_3105,N_3123);
nand U3343 (N_3343,N_3098,N_3033);
xor U3344 (N_3344,N_3078,N_3023);
nor U3345 (N_3345,N_3055,N_3116);
nor U3346 (N_3346,N_3268,N_3163);
nor U3347 (N_3347,N_3217,N_3194);
and U3348 (N_3348,N_3095,N_3232);
and U3349 (N_3349,N_3129,N_3017);
xnor U3350 (N_3350,N_3004,N_3130);
and U3351 (N_3351,N_3248,N_3271);
nor U3352 (N_3352,N_3038,N_3277);
or U3353 (N_3353,N_3049,N_3069);
and U3354 (N_3354,N_3051,N_3168);
nor U3355 (N_3355,N_3157,N_3165);
and U3356 (N_3356,N_3261,N_3178);
or U3357 (N_3357,N_3210,N_3276);
xor U3358 (N_3358,N_3109,N_3062);
nor U3359 (N_3359,N_3275,N_3190);
xor U3360 (N_3360,N_3187,N_3080);
nor U3361 (N_3361,N_3083,N_3026);
xnor U3362 (N_3362,N_3230,N_3151);
or U3363 (N_3363,N_3241,N_3050);
nand U3364 (N_3364,N_3115,N_3034);
nand U3365 (N_3365,N_3240,N_3182);
and U3366 (N_3366,N_3072,N_3287);
nor U3367 (N_3367,N_3079,N_3227);
or U3368 (N_3368,N_3138,N_3280);
xnor U3369 (N_3369,N_3136,N_3088);
nor U3370 (N_3370,N_3066,N_3285);
or U3371 (N_3371,N_3132,N_3067);
nand U3372 (N_3372,N_3099,N_3236);
xnor U3373 (N_3373,N_3253,N_3244);
xor U3374 (N_3374,N_3076,N_3199);
or U3375 (N_3375,N_3077,N_3211);
xor U3376 (N_3376,N_3025,N_3065);
and U3377 (N_3377,N_3035,N_3147);
nand U3378 (N_3378,N_3156,N_3044);
xor U3379 (N_3379,N_3169,N_3299);
nand U3380 (N_3380,N_3257,N_3202);
or U3381 (N_3381,N_3106,N_3247);
or U3382 (N_3382,N_3269,N_3243);
or U3383 (N_3383,N_3085,N_3121);
nor U3384 (N_3384,N_3101,N_3238);
and U3385 (N_3385,N_3117,N_3278);
or U3386 (N_3386,N_3173,N_3272);
or U3387 (N_3387,N_3258,N_3092);
nand U3388 (N_3388,N_3028,N_3061);
or U3389 (N_3389,N_3139,N_3140);
and U3390 (N_3390,N_3149,N_3111);
and U3391 (N_3391,N_3094,N_3096);
nand U3392 (N_3392,N_3084,N_3221);
xnor U3393 (N_3393,N_3131,N_3012);
nor U3394 (N_3394,N_3209,N_3122);
xor U3395 (N_3395,N_3071,N_3263);
and U3396 (N_3396,N_3193,N_3186);
xnor U3397 (N_3397,N_3073,N_3198);
xnor U3398 (N_3398,N_3125,N_3260);
nand U3399 (N_3399,N_3070,N_3196);
and U3400 (N_3400,N_3158,N_3011);
and U3401 (N_3401,N_3045,N_3112);
xnor U3402 (N_3402,N_3283,N_3014);
nand U3403 (N_3403,N_3009,N_3030);
xor U3404 (N_3404,N_3137,N_3146);
nand U3405 (N_3405,N_3119,N_3041);
nor U3406 (N_3406,N_3093,N_3126);
xor U3407 (N_3407,N_3074,N_3229);
nor U3408 (N_3408,N_3003,N_3124);
xor U3409 (N_3409,N_3108,N_3087);
nor U3410 (N_3410,N_3016,N_3056);
and U3411 (N_3411,N_3110,N_3265);
nor U3412 (N_3412,N_3234,N_3286);
xnor U3413 (N_3413,N_3237,N_3086);
xor U3414 (N_3414,N_3282,N_3224);
nand U3415 (N_3415,N_3289,N_3052);
or U3416 (N_3416,N_3155,N_3213);
xor U3417 (N_3417,N_3246,N_3029);
nor U3418 (N_3418,N_3046,N_3002);
nor U3419 (N_3419,N_3220,N_3223);
xnor U3420 (N_3420,N_3013,N_3161);
xnor U3421 (N_3421,N_3216,N_3254);
or U3422 (N_3422,N_3188,N_3171);
xor U3423 (N_3423,N_3184,N_3192);
nor U3424 (N_3424,N_3208,N_3135);
or U3425 (N_3425,N_3054,N_3206);
xor U3426 (N_3426,N_3200,N_3242);
nor U3427 (N_3427,N_3000,N_3195);
nor U3428 (N_3428,N_3143,N_3060);
xnor U3429 (N_3429,N_3128,N_3021);
and U3430 (N_3430,N_3207,N_3082);
nand U3431 (N_3431,N_3005,N_3018);
nor U3432 (N_3432,N_3297,N_3145);
xor U3433 (N_3433,N_3203,N_3001);
and U3434 (N_3434,N_3097,N_3293);
or U3435 (N_3435,N_3252,N_3164);
nand U3436 (N_3436,N_3273,N_3264);
and U3437 (N_3437,N_3089,N_3292);
nand U3438 (N_3438,N_3006,N_3231);
nor U3439 (N_3439,N_3159,N_3118);
and U3440 (N_3440,N_3219,N_3174);
and U3441 (N_3441,N_3075,N_3177);
xnor U3442 (N_3442,N_3114,N_3176);
and U3443 (N_3443,N_3255,N_3104);
nor U3444 (N_3444,N_3183,N_3290);
and U3445 (N_3445,N_3047,N_3204);
nor U3446 (N_3446,N_3191,N_3284);
xnor U3447 (N_3447,N_3064,N_3259);
and U3448 (N_3448,N_3027,N_3239);
or U3449 (N_3449,N_3256,N_3037);
nand U3450 (N_3450,N_3031,N_3027);
or U3451 (N_3451,N_3158,N_3116);
or U3452 (N_3452,N_3221,N_3287);
or U3453 (N_3453,N_3186,N_3052);
nand U3454 (N_3454,N_3030,N_3156);
xnor U3455 (N_3455,N_3209,N_3187);
xnor U3456 (N_3456,N_3201,N_3228);
nand U3457 (N_3457,N_3153,N_3156);
xor U3458 (N_3458,N_3062,N_3032);
and U3459 (N_3459,N_3085,N_3298);
nand U3460 (N_3460,N_3275,N_3005);
and U3461 (N_3461,N_3165,N_3138);
nand U3462 (N_3462,N_3205,N_3149);
nand U3463 (N_3463,N_3223,N_3102);
or U3464 (N_3464,N_3208,N_3189);
or U3465 (N_3465,N_3124,N_3030);
and U3466 (N_3466,N_3204,N_3165);
and U3467 (N_3467,N_3206,N_3168);
xnor U3468 (N_3468,N_3117,N_3291);
nor U3469 (N_3469,N_3244,N_3239);
or U3470 (N_3470,N_3281,N_3067);
xnor U3471 (N_3471,N_3040,N_3285);
and U3472 (N_3472,N_3236,N_3036);
xor U3473 (N_3473,N_3179,N_3104);
xor U3474 (N_3474,N_3012,N_3194);
xnor U3475 (N_3475,N_3232,N_3253);
or U3476 (N_3476,N_3143,N_3139);
xnor U3477 (N_3477,N_3002,N_3102);
or U3478 (N_3478,N_3094,N_3286);
nand U3479 (N_3479,N_3141,N_3078);
nand U3480 (N_3480,N_3185,N_3046);
nor U3481 (N_3481,N_3247,N_3251);
xor U3482 (N_3482,N_3022,N_3105);
and U3483 (N_3483,N_3172,N_3055);
nor U3484 (N_3484,N_3226,N_3269);
or U3485 (N_3485,N_3118,N_3072);
nand U3486 (N_3486,N_3263,N_3018);
nor U3487 (N_3487,N_3139,N_3249);
nor U3488 (N_3488,N_3262,N_3189);
xnor U3489 (N_3489,N_3117,N_3299);
nand U3490 (N_3490,N_3100,N_3222);
nor U3491 (N_3491,N_3089,N_3093);
or U3492 (N_3492,N_3054,N_3029);
nor U3493 (N_3493,N_3246,N_3205);
nand U3494 (N_3494,N_3161,N_3035);
nor U3495 (N_3495,N_3018,N_3196);
xnor U3496 (N_3496,N_3134,N_3197);
and U3497 (N_3497,N_3272,N_3253);
nand U3498 (N_3498,N_3034,N_3178);
xor U3499 (N_3499,N_3033,N_3142);
and U3500 (N_3500,N_3123,N_3249);
and U3501 (N_3501,N_3218,N_3000);
or U3502 (N_3502,N_3265,N_3206);
nand U3503 (N_3503,N_3147,N_3093);
and U3504 (N_3504,N_3037,N_3209);
and U3505 (N_3505,N_3107,N_3098);
and U3506 (N_3506,N_3098,N_3263);
nand U3507 (N_3507,N_3170,N_3072);
xor U3508 (N_3508,N_3032,N_3061);
nand U3509 (N_3509,N_3285,N_3280);
xor U3510 (N_3510,N_3264,N_3259);
nand U3511 (N_3511,N_3062,N_3025);
and U3512 (N_3512,N_3274,N_3185);
and U3513 (N_3513,N_3088,N_3100);
nor U3514 (N_3514,N_3176,N_3093);
and U3515 (N_3515,N_3234,N_3041);
nor U3516 (N_3516,N_3066,N_3229);
nor U3517 (N_3517,N_3224,N_3168);
nor U3518 (N_3518,N_3229,N_3096);
nor U3519 (N_3519,N_3128,N_3223);
nor U3520 (N_3520,N_3007,N_3189);
or U3521 (N_3521,N_3195,N_3136);
and U3522 (N_3522,N_3152,N_3151);
nand U3523 (N_3523,N_3030,N_3121);
nor U3524 (N_3524,N_3068,N_3130);
or U3525 (N_3525,N_3126,N_3131);
or U3526 (N_3526,N_3098,N_3197);
and U3527 (N_3527,N_3113,N_3178);
nand U3528 (N_3528,N_3109,N_3009);
nor U3529 (N_3529,N_3298,N_3158);
xnor U3530 (N_3530,N_3045,N_3001);
xor U3531 (N_3531,N_3258,N_3023);
xor U3532 (N_3532,N_3104,N_3292);
and U3533 (N_3533,N_3058,N_3201);
nand U3534 (N_3534,N_3123,N_3164);
nor U3535 (N_3535,N_3168,N_3021);
nand U3536 (N_3536,N_3071,N_3191);
xor U3537 (N_3537,N_3099,N_3188);
xnor U3538 (N_3538,N_3283,N_3238);
xnor U3539 (N_3539,N_3084,N_3231);
and U3540 (N_3540,N_3095,N_3122);
or U3541 (N_3541,N_3156,N_3157);
nor U3542 (N_3542,N_3105,N_3215);
nor U3543 (N_3543,N_3241,N_3258);
or U3544 (N_3544,N_3032,N_3091);
and U3545 (N_3545,N_3220,N_3117);
or U3546 (N_3546,N_3295,N_3102);
and U3547 (N_3547,N_3000,N_3151);
and U3548 (N_3548,N_3296,N_3061);
nand U3549 (N_3549,N_3244,N_3095);
xor U3550 (N_3550,N_3036,N_3143);
nor U3551 (N_3551,N_3127,N_3235);
or U3552 (N_3552,N_3213,N_3069);
xnor U3553 (N_3553,N_3202,N_3011);
nand U3554 (N_3554,N_3021,N_3009);
nor U3555 (N_3555,N_3240,N_3226);
and U3556 (N_3556,N_3118,N_3222);
and U3557 (N_3557,N_3296,N_3129);
or U3558 (N_3558,N_3173,N_3172);
nor U3559 (N_3559,N_3009,N_3053);
xnor U3560 (N_3560,N_3027,N_3085);
xor U3561 (N_3561,N_3277,N_3161);
nor U3562 (N_3562,N_3224,N_3144);
nand U3563 (N_3563,N_3053,N_3111);
and U3564 (N_3564,N_3115,N_3286);
xnor U3565 (N_3565,N_3159,N_3224);
and U3566 (N_3566,N_3116,N_3234);
xnor U3567 (N_3567,N_3017,N_3224);
or U3568 (N_3568,N_3127,N_3209);
or U3569 (N_3569,N_3093,N_3060);
nand U3570 (N_3570,N_3049,N_3243);
nand U3571 (N_3571,N_3040,N_3115);
xnor U3572 (N_3572,N_3247,N_3201);
nand U3573 (N_3573,N_3116,N_3097);
xor U3574 (N_3574,N_3194,N_3220);
and U3575 (N_3575,N_3044,N_3103);
or U3576 (N_3576,N_3114,N_3175);
and U3577 (N_3577,N_3085,N_3296);
and U3578 (N_3578,N_3010,N_3234);
nand U3579 (N_3579,N_3272,N_3120);
nand U3580 (N_3580,N_3088,N_3050);
xnor U3581 (N_3581,N_3195,N_3205);
xnor U3582 (N_3582,N_3126,N_3285);
and U3583 (N_3583,N_3282,N_3100);
xor U3584 (N_3584,N_3162,N_3253);
and U3585 (N_3585,N_3236,N_3160);
nand U3586 (N_3586,N_3106,N_3262);
nor U3587 (N_3587,N_3056,N_3074);
nand U3588 (N_3588,N_3210,N_3293);
and U3589 (N_3589,N_3095,N_3263);
and U3590 (N_3590,N_3040,N_3097);
or U3591 (N_3591,N_3003,N_3243);
xor U3592 (N_3592,N_3066,N_3195);
nor U3593 (N_3593,N_3289,N_3268);
and U3594 (N_3594,N_3134,N_3234);
or U3595 (N_3595,N_3241,N_3150);
nand U3596 (N_3596,N_3248,N_3231);
or U3597 (N_3597,N_3295,N_3172);
nor U3598 (N_3598,N_3009,N_3167);
xnor U3599 (N_3599,N_3298,N_3214);
and U3600 (N_3600,N_3498,N_3333);
and U3601 (N_3601,N_3534,N_3416);
nand U3602 (N_3602,N_3320,N_3451);
or U3603 (N_3603,N_3395,N_3472);
nor U3604 (N_3604,N_3542,N_3474);
and U3605 (N_3605,N_3371,N_3506);
and U3606 (N_3606,N_3501,N_3400);
xor U3607 (N_3607,N_3379,N_3438);
nor U3608 (N_3608,N_3316,N_3512);
or U3609 (N_3609,N_3563,N_3556);
and U3610 (N_3610,N_3356,N_3423);
and U3611 (N_3611,N_3490,N_3419);
nor U3612 (N_3612,N_3377,N_3365);
nand U3613 (N_3613,N_3524,N_3574);
nand U3614 (N_3614,N_3376,N_3595);
or U3615 (N_3615,N_3433,N_3315);
and U3616 (N_3616,N_3483,N_3437);
or U3617 (N_3617,N_3560,N_3578);
nand U3618 (N_3618,N_3361,N_3328);
and U3619 (N_3619,N_3525,N_3552);
nand U3620 (N_3620,N_3541,N_3477);
and U3621 (N_3621,N_3457,N_3439);
and U3622 (N_3622,N_3460,N_3344);
nor U3623 (N_3623,N_3456,N_3367);
nor U3624 (N_3624,N_3455,N_3346);
or U3625 (N_3625,N_3493,N_3470);
nor U3626 (N_3626,N_3468,N_3485);
xor U3627 (N_3627,N_3504,N_3445);
or U3628 (N_3628,N_3325,N_3406);
or U3629 (N_3629,N_3467,N_3586);
xor U3630 (N_3630,N_3517,N_3374);
and U3631 (N_3631,N_3454,N_3546);
nand U3632 (N_3632,N_3398,N_3394);
nor U3633 (N_3633,N_3370,N_3413);
xnor U3634 (N_3634,N_3307,N_3348);
nand U3635 (N_3635,N_3469,N_3597);
nor U3636 (N_3636,N_3463,N_3588);
and U3637 (N_3637,N_3473,N_3547);
nand U3638 (N_3638,N_3415,N_3475);
nand U3639 (N_3639,N_3570,N_3554);
nor U3640 (N_3640,N_3324,N_3514);
nand U3641 (N_3641,N_3411,N_3354);
or U3642 (N_3642,N_3382,N_3491);
and U3643 (N_3643,N_3311,N_3424);
and U3644 (N_3644,N_3532,N_3562);
nand U3645 (N_3645,N_3579,N_3386);
or U3646 (N_3646,N_3568,N_3387);
and U3647 (N_3647,N_3596,N_3323);
or U3648 (N_3648,N_3511,N_3355);
nand U3649 (N_3649,N_3599,N_3375);
xnor U3650 (N_3650,N_3434,N_3378);
or U3651 (N_3651,N_3566,N_3304);
xnor U3652 (N_3652,N_3340,N_3435);
nand U3653 (N_3653,N_3523,N_3426);
nand U3654 (N_3654,N_3543,N_3381);
or U3655 (N_3655,N_3580,N_3393);
xor U3656 (N_3656,N_3336,N_3352);
and U3657 (N_3657,N_3521,N_3519);
nor U3658 (N_3658,N_3332,N_3510);
xor U3659 (N_3659,N_3412,N_3572);
or U3660 (N_3660,N_3430,N_3421);
xor U3661 (N_3661,N_3507,N_3418);
and U3662 (N_3662,N_3341,N_3312);
nand U3663 (N_3663,N_3571,N_3366);
xor U3664 (N_3664,N_3487,N_3347);
xnor U3665 (N_3665,N_3446,N_3389);
nand U3666 (N_3666,N_3591,N_3520);
xor U3667 (N_3667,N_3453,N_3497);
and U3668 (N_3668,N_3443,N_3334);
nand U3669 (N_3669,N_3442,N_3399);
and U3670 (N_3670,N_3544,N_3515);
xor U3671 (N_3671,N_3590,N_3425);
and U3672 (N_3672,N_3372,N_3585);
and U3673 (N_3673,N_3549,N_3531);
and U3674 (N_3674,N_3569,N_3353);
nand U3675 (N_3675,N_3397,N_3561);
and U3676 (N_3676,N_3499,N_3404);
or U3677 (N_3677,N_3441,N_3494);
and U3678 (N_3678,N_3300,N_3500);
nor U3679 (N_3679,N_3318,N_3385);
and U3680 (N_3680,N_3310,N_3535);
nand U3681 (N_3681,N_3509,N_3301);
or U3682 (N_3682,N_3537,N_3350);
or U3683 (N_3683,N_3440,N_3528);
nand U3684 (N_3684,N_3388,N_3536);
and U3685 (N_3685,N_3558,N_3427);
nand U3686 (N_3686,N_3409,N_3380);
or U3687 (N_3687,N_3584,N_3429);
or U3688 (N_3688,N_3464,N_3466);
xor U3689 (N_3689,N_3349,N_3502);
xnor U3690 (N_3690,N_3327,N_3436);
nand U3691 (N_3691,N_3471,N_3476);
nand U3692 (N_3692,N_3577,N_3326);
and U3693 (N_3693,N_3548,N_3593);
nor U3694 (N_3694,N_3362,N_3410);
nand U3695 (N_3695,N_3305,N_3539);
or U3696 (N_3696,N_3363,N_3486);
nor U3697 (N_3697,N_3383,N_3308);
xnor U3698 (N_3698,N_3351,N_3496);
nand U3699 (N_3699,N_3321,N_3575);
nor U3700 (N_3700,N_3422,N_3581);
nand U3701 (N_3701,N_3302,N_3503);
or U3702 (N_3702,N_3533,N_3331);
or U3703 (N_3703,N_3319,N_3565);
xor U3704 (N_3704,N_3551,N_3492);
nor U3705 (N_3705,N_3358,N_3407);
nor U3706 (N_3706,N_3432,N_3545);
nor U3707 (N_3707,N_3309,N_3317);
nor U3708 (N_3708,N_3369,N_3417);
nor U3709 (N_3709,N_3522,N_3553);
xnor U3710 (N_3710,N_3480,N_3306);
nor U3711 (N_3711,N_3555,N_3414);
nor U3712 (N_3712,N_3530,N_3390);
or U3713 (N_3713,N_3465,N_3489);
xor U3714 (N_3714,N_3484,N_3482);
nand U3715 (N_3715,N_3529,N_3357);
xor U3716 (N_3716,N_3458,N_3462);
nand U3717 (N_3717,N_3364,N_3505);
and U3718 (N_3718,N_3527,N_3401);
nor U3719 (N_3719,N_3559,N_3449);
nand U3720 (N_3720,N_3342,N_3587);
and U3721 (N_3721,N_3448,N_3391);
and U3722 (N_3722,N_3329,N_3508);
xnor U3723 (N_3723,N_3481,N_3360);
or U3724 (N_3724,N_3330,N_3478);
and U3725 (N_3725,N_3550,N_3582);
xnor U3726 (N_3726,N_3459,N_3479);
xnor U3727 (N_3727,N_3567,N_3538);
xor U3728 (N_3728,N_3573,N_3518);
xor U3729 (N_3729,N_3513,N_3339);
xor U3730 (N_3730,N_3598,N_3405);
and U3731 (N_3731,N_3420,N_3576);
nor U3732 (N_3732,N_3526,N_3540);
or U3733 (N_3733,N_3313,N_3392);
and U3734 (N_3734,N_3335,N_3396);
nand U3735 (N_3735,N_3444,N_3589);
xor U3736 (N_3736,N_3495,N_3408);
nor U3737 (N_3737,N_3428,N_3431);
or U3738 (N_3738,N_3384,N_3368);
and U3739 (N_3739,N_3338,N_3359);
xnor U3740 (N_3740,N_3564,N_3303);
xor U3741 (N_3741,N_3461,N_3583);
nor U3742 (N_3742,N_3373,N_3322);
nor U3743 (N_3743,N_3557,N_3314);
or U3744 (N_3744,N_3337,N_3345);
and U3745 (N_3745,N_3516,N_3592);
nor U3746 (N_3746,N_3343,N_3403);
and U3747 (N_3747,N_3594,N_3488);
nand U3748 (N_3748,N_3452,N_3450);
or U3749 (N_3749,N_3447,N_3402);
nor U3750 (N_3750,N_3452,N_3411);
nand U3751 (N_3751,N_3484,N_3589);
xnor U3752 (N_3752,N_3344,N_3423);
nor U3753 (N_3753,N_3372,N_3425);
nor U3754 (N_3754,N_3392,N_3550);
nand U3755 (N_3755,N_3316,N_3340);
nand U3756 (N_3756,N_3473,N_3421);
or U3757 (N_3757,N_3385,N_3507);
nand U3758 (N_3758,N_3442,N_3324);
nor U3759 (N_3759,N_3540,N_3376);
nand U3760 (N_3760,N_3418,N_3590);
nor U3761 (N_3761,N_3582,N_3310);
nor U3762 (N_3762,N_3413,N_3500);
or U3763 (N_3763,N_3440,N_3521);
nand U3764 (N_3764,N_3390,N_3325);
or U3765 (N_3765,N_3543,N_3420);
xor U3766 (N_3766,N_3474,N_3436);
or U3767 (N_3767,N_3381,N_3511);
nor U3768 (N_3768,N_3330,N_3383);
and U3769 (N_3769,N_3536,N_3514);
or U3770 (N_3770,N_3475,N_3361);
xnor U3771 (N_3771,N_3471,N_3342);
nand U3772 (N_3772,N_3561,N_3301);
xor U3773 (N_3773,N_3458,N_3586);
nor U3774 (N_3774,N_3339,N_3480);
or U3775 (N_3775,N_3422,N_3557);
and U3776 (N_3776,N_3315,N_3332);
nor U3777 (N_3777,N_3300,N_3399);
and U3778 (N_3778,N_3528,N_3385);
xor U3779 (N_3779,N_3412,N_3335);
nor U3780 (N_3780,N_3480,N_3407);
and U3781 (N_3781,N_3526,N_3480);
nor U3782 (N_3782,N_3347,N_3406);
nand U3783 (N_3783,N_3434,N_3306);
or U3784 (N_3784,N_3322,N_3528);
or U3785 (N_3785,N_3569,N_3413);
xor U3786 (N_3786,N_3393,N_3544);
nor U3787 (N_3787,N_3539,N_3595);
nor U3788 (N_3788,N_3598,N_3567);
and U3789 (N_3789,N_3492,N_3306);
and U3790 (N_3790,N_3537,N_3489);
or U3791 (N_3791,N_3406,N_3523);
nand U3792 (N_3792,N_3388,N_3366);
nor U3793 (N_3793,N_3422,N_3475);
and U3794 (N_3794,N_3419,N_3539);
nor U3795 (N_3795,N_3561,N_3549);
nand U3796 (N_3796,N_3427,N_3319);
xnor U3797 (N_3797,N_3368,N_3375);
or U3798 (N_3798,N_3454,N_3404);
and U3799 (N_3799,N_3400,N_3425);
or U3800 (N_3800,N_3514,N_3542);
nor U3801 (N_3801,N_3536,N_3371);
nand U3802 (N_3802,N_3320,N_3311);
and U3803 (N_3803,N_3377,N_3304);
nand U3804 (N_3804,N_3384,N_3400);
xnor U3805 (N_3805,N_3487,N_3447);
xnor U3806 (N_3806,N_3400,N_3508);
nor U3807 (N_3807,N_3495,N_3537);
nor U3808 (N_3808,N_3310,N_3509);
nor U3809 (N_3809,N_3537,N_3430);
nand U3810 (N_3810,N_3509,N_3452);
xnor U3811 (N_3811,N_3442,N_3323);
xor U3812 (N_3812,N_3483,N_3597);
nand U3813 (N_3813,N_3361,N_3457);
or U3814 (N_3814,N_3366,N_3544);
xnor U3815 (N_3815,N_3324,N_3558);
and U3816 (N_3816,N_3486,N_3310);
xnor U3817 (N_3817,N_3456,N_3492);
and U3818 (N_3818,N_3382,N_3423);
or U3819 (N_3819,N_3360,N_3485);
or U3820 (N_3820,N_3384,N_3401);
or U3821 (N_3821,N_3566,N_3517);
and U3822 (N_3822,N_3307,N_3598);
and U3823 (N_3823,N_3558,N_3592);
and U3824 (N_3824,N_3321,N_3322);
xor U3825 (N_3825,N_3356,N_3436);
or U3826 (N_3826,N_3338,N_3334);
nor U3827 (N_3827,N_3449,N_3578);
nor U3828 (N_3828,N_3588,N_3582);
nor U3829 (N_3829,N_3326,N_3462);
or U3830 (N_3830,N_3427,N_3554);
nand U3831 (N_3831,N_3528,N_3495);
nor U3832 (N_3832,N_3468,N_3510);
and U3833 (N_3833,N_3561,N_3328);
nand U3834 (N_3834,N_3435,N_3443);
or U3835 (N_3835,N_3411,N_3563);
or U3836 (N_3836,N_3356,N_3303);
nor U3837 (N_3837,N_3409,N_3447);
nand U3838 (N_3838,N_3510,N_3304);
and U3839 (N_3839,N_3311,N_3412);
xor U3840 (N_3840,N_3520,N_3537);
and U3841 (N_3841,N_3406,N_3388);
nand U3842 (N_3842,N_3505,N_3331);
and U3843 (N_3843,N_3432,N_3553);
or U3844 (N_3844,N_3345,N_3482);
or U3845 (N_3845,N_3355,N_3415);
nand U3846 (N_3846,N_3353,N_3529);
nand U3847 (N_3847,N_3541,N_3330);
and U3848 (N_3848,N_3301,N_3399);
nor U3849 (N_3849,N_3490,N_3354);
nor U3850 (N_3850,N_3517,N_3472);
xor U3851 (N_3851,N_3311,N_3367);
xnor U3852 (N_3852,N_3360,N_3368);
nor U3853 (N_3853,N_3510,N_3379);
nor U3854 (N_3854,N_3473,N_3433);
nand U3855 (N_3855,N_3537,N_3538);
or U3856 (N_3856,N_3425,N_3515);
xor U3857 (N_3857,N_3570,N_3418);
xor U3858 (N_3858,N_3318,N_3592);
and U3859 (N_3859,N_3516,N_3436);
nand U3860 (N_3860,N_3505,N_3373);
and U3861 (N_3861,N_3470,N_3448);
or U3862 (N_3862,N_3525,N_3563);
and U3863 (N_3863,N_3596,N_3487);
or U3864 (N_3864,N_3301,N_3381);
or U3865 (N_3865,N_3390,N_3589);
or U3866 (N_3866,N_3302,N_3433);
nand U3867 (N_3867,N_3570,N_3595);
nand U3868 (N_3868,N_3384,N_3430);
or U3869 (N_3869,N_3310,N_3454);
nor U3870 (N_3870,N_3360,N_3384);
xnor U3871 (N_3871,N_3343,N_3556);
nand U3872 (N_3872,N_3332,N_3457);
and U3873 (N_3873,N_3497,N_3362);
or U3874 (N_3874,N_3335,N_3417);
and U3875 (N_3875,N_3365,N_3376);
or U3876 (N_3876,N_3300,N_3509);
nor U3877 (N_3877,N_3554,N_3309);
nor U3878 (N_3878,N_3417,N_3543);
nor U3879 (N_3879,N_3483,N_3457);
nor U3880 (N_3880,N_3535,N_3322);
xor U3881 (N_3881,N_3414,N_3575);
nor U3882 (N_3882,N_3387,N_3340);
nand U3883 (N_3883,N_3566,N_3406);
xnor U3884 (N_3884,N_3440,N_3598);
or U3885 (N_3885,N_3356,N_3409);
or U3886 (N_3886,N_3314,N_3403);
or U3887 (N_3887,N_3307,N_3316);
nand U3888 (N_3888,N_3508,N_3433);
nand U3889 (N_3889,N_3459,N_3554);
xor U3890 (N_3890,N_3462,N_3474);
nand U3891 (N_3891,N_3335,N_3389);
or U3892 (N_3892,N_3483,N_3325);
or U3893 (N_3893,N_3363,N_3536);
or U3894 (N_3894,N_3337,N_3545);
xnor U3895 (N_3895,N_3359,N_3485);
nor U3896 (N_3896,N_3432,N_3352);
and U3897 (N_3897,N_3426,N_3499);
or U3898 (N_3898,N_3571,N_3516);
nor U3899 (N_3899,N_3357,N_3449);
nor U3900 (N_3900,N_3808,N_3869);
nor U3901 (N_3901,N_3717,N_3874);
and U3902 (N_3902,N_3616,N_3889);
nor U3903 (N_3903,N_3658,N_3673);
nor U3904 (N_3904,N_3685,N_3784);
or U3905 (N_3905,N_3881,N_3709);
and U3906 (N_3906,N_3842,N_3640);
and U3907 (N_3907,N_3660,N_3830);
and U3908 (N_3908,N_3811,N_3780);
xnor U3909 (N_3909,N_3634,N_3679);
nand U3910 (N_3910,N_3666,N_3703);
and U3911 (N_3911,N_3769,N_3623);
or U3912 (N_3912,N_3814,N_3887);
nor U3913 (N_3913,N_3740,N_3799);
nand U3914 (N_3914,N_3846,N_3826);
or U3915 (N_3915,N_3820,N_3608);
xor U3916 (N_3916,N_3661,N_3773);
nand U3917 (N_3917,N_3641,N_3655);
nand U3918 (N_3918,N_3771,N_3859);
and U3919 (N_3919,N_3809,N_3768);
nor U3920 (N_3920,N_3840,N_3801);
or U3921 (N_3921,N_3677,N_3795);
and U3922 (N_3922,N_3860,N_3630);
nand U3923 (N_3923,N_3624,N_3744);
and U3924 (N_3924,N_3650,N_3878);
nor U3925 (N_3925,N_3631,N_3725);
or U3926 (N_3926,N_3837,N_3804);
nor U3927 (N_3927,N_3705,N_3712);
xor U3928 (N_3928,N_3827,N_3745);
nor U3929 (N_3929,N_3733,N_3895);
and U3930 (N_3930,N_3606,N_3607);
nor U3931 (N_3931,N_3684,N_3806);
nor U3932 (N_3932,N_3824,N_3766);
nor U3933 (N_3933,N_3721,N_3877);
nor U3934 (N_3934,N_3767,N_3639);
and U3935 (N_3935,N_3803,N_3702);
nand U3936 (N_3936,N_3752,N_3861);
and U3937 (N_3937,N_3776,N_3671);
xnor U3938 (N_3938,N_3855,N_3600);
nand U3939 (N_3939,N_3815,N_3839);
nor U3940 (N_3940,N_3646,N_3796);
nand U3941 (N_3941,N_3612,N_3680);
and U3942 (N_3942,N_3864,N_3831);
and U3943 (N_3943,N_3753,N_3619);
or U3944 (N_3944,N_3694,N_3622);
xor U3945 (N_3945,N_3833,N_3629);
and U3946 (N_3946,N_3708,N_3763);
xnor U3947 (N_3947,N_3618,N_3838);
xnor U3948 (N_3948,N_3720,N_3603);
nand U3949 (N_3949,N_3653,N_3649);
xnor U3950 (N_3950,N_3698,N_3664);
and U3951 (N_3951,N_3888,N_3870);
nand U3952 (N_3952,N_3893,N_3690);
and U3953 (N_3953,N_3798,N_3851);
and U3954 (N_3954,N_3693,N_3691);
and U3955 (N_3955,N_3689,N_3627);
or U3956 (N_3956,N_3852,N_3654);
nand U3957 (N_3957,N_3880,N_3682);
nand U3958 (N_3958,N_3797,N_3626);
xnor U3959 (N_3959,N_3734,N_3657);
nor U3960 (N_3960,N_3778,N_3710);
nand U3961 (N_3961,N_3670,N_3873);
or U3962 (N_3962,N_3628,N_3754);
nand U3963 (N_3963,N_3621,N_3807);
and U3964 (N_3964,N_3747,N_3835);
xor U3965 (N_3965,N_3805,N_3735);
nand U3966 (N_3966,N_3697,N_3772);
nand U3967 (N_3967,N_3704,N_3898);
and U3968 (N_3968,N_3821,N_3891);
xor U3969 (N_3969,N_3847,N_3637);
nor U3970 (N_3970,N_3786,N_3722);
or U3971 (N_3971,N_3866,N_3739);
and U3972 (N_3972,N_3897,N_3848);
nor U3973 (N_3973,N_3668,N_3858);
or U3974 (N_3974,N_3755,N_3865);
or U3975 (N_3975,N_3609,N_3647);
or U3976 (N_3976,N_3794,N_3672);
nor U3977 (N_3977,N_3743,N_3765);
xor U3978 (N_3978,N_3706,N_3883);
and U3979 (N_3979,N_3802,N_3890);
and U3980 (N_3980,N_3678,N_3882);
or U3981 (N_3981,N_3764,N_3617);
or U3982 (N_3982,N_3719,N_3762);
nor U3983 (N_3983,N_3834,N_3662);
nand U3984 (N_3984,N_3812,N_3711);
nand U3985 (N_3985,N_3876,N_3688);
nor U3986 (N_3986,N_3669,N_3868);
nand U3987 (N_3987,N_3714,N_3791);
xnor U3988 (N_3988,N_3885,N_3867);
and U3989 (N_3989,N_3856,N_3849);
nor U3990 (N_3990,N_3850,N_3782);
nor U3991 (N_3991,N_3665,N_3686);
nand U3992 (N_3992,N_3775,N_3793);
or U3993 (N_3993,N_3853,N_3841);
xor U3994 (N_3994,N_3800,N_3718);
or U3995 (N_3995,N_3854,N_3728);
nand U3996 (N_3996,N_3816,N_3746);
nand U3997 (N_3997,N_3643,N_3674);
or U3998 (N_3998,N_3894,N_3723);
and U3999 (N_3999,N_3749,N_3620);
or U4000 (N_4000,N_3611,N_3737);
or U4001 (N_4001,N_3632,N_3615);
and U4002 (N_4002,N_3695,N_3651);
or U4003 (N_4003,N_3787,N_3604);
and U4004 (N_4004,N_3879,N_3758);
xor U4005 (N_4005,N_3727,N_3692);
nand U4006 (N_4006,N_3843,N_3642);
and U4007 (N_4007,N_3610,N_3715);
and U4008 (N_4008,N_3732,N_3681);
nand U4009 (N_4009,N_3687,N_3676);
or U4010 (N_4010,N_3770,N_3817);
nor U4011 (N_4011,N_3818,N_3748);
and U4012 (N_4012,N_3648,N_3844);
nor U4013 (N_4013,N_3731,N_3699);
and U4014 (N_4014,N_3810,N_3667);
nand U4015 (N_4015,N_3845,N_3638);
and U4016 (N_4016,N_3783,N_3781);
nor U4017 (N_4017,N_3823,N_3701);
and U4018 (N_4018,N_3777,N_3605);
and U4019 (N_4019,N_3892,N_3863);
nand U4020 (N_4020,N_3713,N_3785);
and U4021 (N_4021,N_3790,N_3871);
and U4022 (N_4022,N_3614,N_3645);
xnor U4023 (N_4023,N_3724,N_3736);
xor U4024 (N_4024,N_3601,N_3716);
or U4025 (N_4025,N_3774,N_3779);
xnor U4026 (N_4026,N_3625,N_3886);
xor U4027 (N_4027,N_3750,N_3696);
nand U4028 (N_4028,N_3875,N_3822);
or U4029 (N_4029,N_3683,N_3644);
and U4030 (N_4030,N_3899,N_3741);
nand U4031 (N_4031,N_3659,N_3700);
or U4032 (N_4032,N_3759,N_3896);
nand U4033 (N_4033,N_3829,N_3836);
xor U4034 (N_4034,N_3636,N_3788);
nor U4035 (N_4035,N_3635,N_3862);
nand U4036 (N_4036,N_3884,N_3789);
nor U4037 (N_4037,N_3792,N_3613);
nand U4038 (N_4038,N_3813,N_3602);
and U4039 (N_4039,N_3832,N_3760);
or U4040 (N_4040,N_3633,N_3675);
xor U4041 (N_4041,N_3857,N_3730);
nor U4042 (N_4042,N_3656,N_3726);
nor U4043 (N_4043,N_3825,N_3756);
or U4044 (N_4044,N_3729,N_3872);
nand U4045 (N_4045,N_3819,N_3663);
nand U4046 (N_4046,N_3761,N_3751);
and U4047 (N_4047,N_3757,N_3652);
xnor U4048 (N_4048,N_3707,N_3828);
nor U4049 (N_4049,N_3742,N_3738);
xnor U4050 (N_4050,N_3678,N_3690);
and U4051 (N_4051,N_3827,N_3753);
nor U4052 (N_4052,N_3781,N_3695);
and U4053 (N_4053,N_3697,N_3802);
xnor U4054 (N_4054,N_3617,N_3826);
xor U4055 (N_4055,N_3850,N_3724);
nor U4056 (N_4056,N_3741,N_3772);
nand U4057 (N_4057,N_3742,N_3689);
or U4058 (N_4058,N_3720,N_3714);
nor U4059 (N_4059,N_3631,N_3893);
and U4060 (N_4060,N_3832,N_3863);
nor U4061 (N_4061,N_3600,N_3720);
and U4062 (N_4062,N_3664,N_3714);
nor U4063 (N_4063,N_3702,N_3853);
nand U4064 (N_4064,N_3794,N_3677);
xor U4065 (N_4065,N_3671,N_3647);
nor U4066 (N_4066,N_3630,N_3610);
xor U4067 (N_4067,N_3833,N_3809);
and U4068 (N_4068,N_3816,N_3687);
nor U4069 (N_4069,N_3771,N_3789);
nand U4070 (N_4070,N_3697,N_3637);
nor U4071 (N_4071,N_3891,N_3830);
xnor U4072 (N_4072,N_3809,N_3849);
and U4073 (N_4073,N_3749,N_3728);
and U4074 (N_4074,N_3899,N_3646);
nand U4075 (N_4075,N_3697,N_3602);
or U4076 (N_4076,N_3666,N_3804);
xor U4077 (N_4077,N_3756,N_3729);
and U4078 (N_4078,N_3884,N_3637);
or U4079 (N_4079,N_3665,N_3728);
and U4080 (N_4080,N_3853,N_3611);
nand U4081 (N_4081,N_3689,N_3841);
or U4082 (N_4082,N_3683,N_3669);
nor U4083 (N_4083,N_3851,N_3838);
nand U4084 (N_4084,N_3606,N_3780);
nor U4085 (N_4085,N_3885,N_3897);
nand U4086 (N_4086,N_3644,N_3619);
and U4087 (N_4087,N_3687,N_3749);
nand U4088 (N_4088,N_3799,N_3719);
nand U4089 (N_4089,N_3652,N_3853);
nand U4090 (N_4090,N_3694,N_3771);
nand U4091 (N_4091,N_3737,N_3766);
xor U4092 (N_4092,N_3642,N_3780);
and U4093 (N_4093,N_3742,N_3752);
or U4094 (N_4094,N_3892,N_3836);
and U4095 (N_4095,N_3821,N_3892);
or U4096 (N_4096,N_3761,N_3875);
and U4097 (N_4097,N_3854,N_3860);
nor U4098 (N_4098,N_3894,N_3801);
nand U4099 (N_4099,N_3777,N_3845);
nor U4100 (N_4100,N_3659,N_3899);
nor U4101 (N_4101,N_3772,N_3779);
nor U4102 (N_4102,N_3642,N_3600);
and U4103 (N_4103,N_3728,N_3604);
nor U4104 (N_4104,N_3711,N_3851);
nor U4105 (N_4105,N_3822,N_3850);
and U4106 (N_4106,N_3659,N_3877);
nand U4107 (N_4107,N_3791,N_3612);
xor U4108 (N_4108,N_3800,N_3676);
and U4109 (N_4109,N_3762,N_3881);
and U4110 (N_4110,N_3674,N_3739);
nand U4111 (N_4111,N_3638,N_3741);
xor U4112 (N_4112,N_3650,N_3699);
or U4113 (N_4113,N_3813,N_3710);
or U4114 (N_4114,N_3690,N_3697);
xnor U4115 (N_4115,N_3721,N_3831);
nor U4116 (N_4116,N_3751,N_3651);
and U4117 (N_4117,N_3614,N_3621);
nand U4118 (N_4118,N_3633,N_3710);
xor U4119 (N_4119,N_3678,N_3687);
nand U4120 (N_4120,N_3730,N_3869);
or U4121 (N_4121,N_3817,N_3607);
and U4122 (N_4122,N_3825,N_3735);
nand U4123 (N_4123,N_3686,N_3672);
nand U4124 (N_4124,N_3745,N_3672);
nor U4125 (N_4125,N_3638,N_3766);
or U4126 (N_4126,N_3844,N_3625);
nand U4127 (N_4127,N_3827,N_3788);
nand U4128 (N_4128,N_3695,N_3870);
xnor U4129 (N_4129,N_3754,N_3679);
xnor U4130 (N_4130,N_3667,N_3622);
nand U4131 (N_4131,N_3688,N_3627);
nand U4132 (N_4132,N_3677,N_3734);
nand U4133 (N_4133,N_3750,N_3804);
nor U4134 (N_4134,N_3612,N_3730);
nand U4135 (N_4135,N_3655,N_3637);
and U4136 (N_4136,N_3799,N_3663);
and U4137 (N_4137,N_3788,N_3810);
xor U4138 (N_4138,N_3849,N_3630);
nor U4139 (N_4139,N_3788,N_3659);
nand U4140 (N_4140,N_3863,N_3660);
nor U4141 (N_4141,N_3838,N_3834);
and U4142 (N_4142,N_3869,N_3740);
or U4143 (N_4143,N_3802,N_3648);
and U4144 (N_4144,N_3686,N_3661);
and U4145 (N_4145,N_3701,N_3778);
xor U4146 (N_4146,N_3794,N_3686);
nor U4147 (N_4147,N_3733,N_3690);
or U4148 (N_4148,N_3790,N_3724);
and U4149 (N_4149,N_3744,N_3727);
nor U4150 (N_4150,N_3878,N_3868);
and U4151 (N_4151,N_3762,N_3731);
nor U4152 (N_4152,N_3832,N_3636);
or U4153 (N_4153,N_3822,N_3676);
and U4154 (N_4154,N_3739,N_3786);
nor U4155 (N_4155,N_3875,N_3824);
nor U4156 (N_4156,N_3783,N_3610);
and U4157 (N_4157,N_3654,N_3608);
xor U4158 (N_4158,N_3863,N_3782);
xor U4159 (N_4159,N_3744,N_3709);
and U4160 (N_4160,N_3622,N_3829);
and U4161 (N_4161,N_3667,N_3821);
or U4162 (N_4162,N_3852,N_3764);
or U4163 (N_4163,N_3682,N_3785);
and U4164 (N_4164,N_3844,N_3893);
or U4165 (N_4165,N_3825,N_3629);
and U4166 (N_4166,N_3657,N_3680);
and U4167 (N_4167,N_3721,N_3696);
nor U4168 (N_4168,N_3687,N_3693);
xor U4169 (N_4169,N_3888,N_3604);
and U4170 (N_4170,N_3890,N_3877);
nor U4171 (N_4171,N_3606,N_3675);
nand U4172 (N_4172,N_3750,N_3651);
or U4173 (N_4173,N_3699,N_3634);
or U4174 (N_4174,N_3675,N_3611);
or U4175 (N_4175,N_3755,N_3748);
nand U4176 (N_4176,N_3861,N_3718);
and U4177 (N_4177,N_3888,N_3805);
nand U4178 (N_4178,N_3692,N_3716);
xor U4179 (N_4179,N_3816,N_3765);
nor U4180 (N_4180,N_3832,N_3662);
and U4181 (N_4181,N_3802,N_3646);
or U4182 (N_4182,N_3676,N_3757);
and U4183 (N_4183,N_3685,N_3611);
xnor U4184 (N_4184,N_3828,N_3815);
or U4185 (N_4185,N_3695,N_3814);
nand U4186 (N_4186,N_3696,N_3859);
nor U4187 (N_4187,N_3857,N_3803);
or U4188 (N_4188,N_3661,N_3662);
xor U4189 (N_4189,N_3652,N_3884);
xor U4190 (N_4190,N_3802,N_3891);
or U4191 (N_4191,N_3755,N_3897);
or U4192 (N_4192,N_3633,N_3666);
and U4193 (N_4193,N_3844,N_3776);
nand U4194 (N_4194,N_3865,N_3783);
or U4195 (N_4195,N_3786,N_3748);
and U4196 (N_4196,N_3838,N_3638);
and U4197 (N_4197,N_3770,N_3665);
or U4198 (N_4198,N_3660,N_3805);
or U4199 (N_4199,N_3794,N_3897);
and U4200 (N_4200,N_3909,N_3943);
and U4201 (N_4201,N_3926,N_4009);
nand U4202 (N_4202,N_3934,N_3942);
and U4203 (N_4203,N_4188,N_4068);
or U4204 (N_4204,N_4138,N_4089);
and U4205 (N_4205,N_4081,N_4056);
and U4206 (N_4206,N_4106,N_3974);
xor U4207 (N_4207,N_4173,N_4163);
or U4208 (N_4208,N_3948,N_4184);
xor U4209 (N_4209,N_4029,N_4050);
nand U4210 (N_4210,N_4170,N_3947);
or U4211 (N_4211,N_4164,N_4146);
or U4212 (N_4212,N_4072,N_4123);
nor U4213 (N_4213,N_4167,N_3922);
nor U4214 (N_4214,N_3977,N_3937);
xnor U4215 (N_4215,N_4044,N_3995);
and U4216 (N_4216,N_4011,N_4093);
xor U4217 (N_4217,N_4113,N_4136);
nor U4218 (N_4218,N_3960,N_4076);
nand U4219 (N_4219,N_4122,N_4031);
or U4220 (N_4220,N_3908,N_3971);
xor U4221 (N_4221,N_3933,N_4128);
xor U4222 (N_4222,N_3915,N_3967);
or U4223 (N_4223,N_4153,N_4114);
or U4224 (N_4224,N_3999,N_3986);
xnor U4225 (N_4225,N_4067,N_4149);
xnor U4226 (N_4226,N_4144,N_3904);
nor U4227 (N_4227,N_4186,N_4079);
nor U4228 (N_4228,N_4018,N_4196);
nor U4229 (N_4229,N_4185,N_3975);
and U4230 (N_4230,N_3913,N_4100);
nand U4231 (N_4231,N_3970,N_4054);
and U4232 (N_4232,N_4063,N_3984);
or U4233 (N_4233,N_4193,N_4069);
or U4234 (N_4234,N_3928,N_3939);
xor U4235 (N_4235,N_4105,N_4126);
nor U4236 (N_4236,N_4133,N_3907);
nand U4237 (N_4237,N_4108,N_3921);
xnor U4238 (N_4238,N_3936,N_3954);
or U4239 (N_4239,N_4092,N_4074);
nand U4240 (N_4240,N_4012,N_3955);
or U4241 (N_4241,N_4145,N_4116);
nand U4242 (N_4242,N_3953,N_4065);
xor U4243 (N_4243,N_3962,N_3978);
or U4244 (N_4244,N_3959,N_3989);
nand U4245 (N_4245,N_4060,N_4005);
and U4246 (N_4246,N_4125,N_4198);
nand U4247 (N_4247,N_4179,N_4160);
and U4248 (N_4248,N_4039,N_4032);
nand U4249 (N_4249,N_4037,N_3930);
nor U4250 (N_4250,N_3966,N_4038);
nor U4251 (N_4251,N_4099,N_4157);
nand U4252 (N_4252,N_3929,N_3964);
nor U4253 (N_4253,N_4177,N_4152);
xnor U4254 (N_4254,N_4033,N_3914);
nand U4255 (N_4255,N_3982,N_3988);
or U4256 (N_4256,N_4066,N_4082);
xnor U4257 (N_4257,N_4021,N_3997);
nor U4258 (N_4258,N_4194,N_4023);
nor U4259 (N_4259,N_3935,N_4174);
and U4260 (N_4260,N_4134,N_4040);
nor U4261 (N_4261,N_4142,N_4191);
or U4262 (N_4262,N_4150,N_3945);
or U4263 (N_4263,N_3979,N_3910);
nand U4264 (N_4264,N_4169,N_3920);
nand U4265 (N_4265,N_4071,N_4045);
nand U4266 (N_4266,N_4176,N_3938);
or U4267 (N_4267,N_4052,N_4083);
or U4268 (N_4268,N_3996,N_4156);
or U4269 (N_4269,N_4182,N_4102);
xnor U4270 (N_4270,N_4112,N_4086);
or U4271 (N_4271,N_3927,N_3993);
nand U4272 (N_4272,N_3991,N_4129);
nor U4273 (N_4273,N_3923,N_4006);
xnor U4274 (N_4274,N_4127,N_4026);
and U4275 (N_4275,N_4141,N_4140);
nor U4276 (N_4276,N_4027,N_4183);
nor U4277 (N_4277,N_3906,N_4130);
or U4278 (N_4278,N_4178,N_4014);
nand U4279 (N_4279,N_4028,N_4043);
or U4280 (N_4280,N_3902,N_4137);
nor U4281 (N_4281,N_4107,N_3998);
xnor U4282 (N_4282,N_4120,N_4084);
and U4283 (N_4283,N_4022,N_3957);
xnor U4284 (N_4284,N_4077,N_3987);
and U4285 (N_4285,N_4020,N_4002);
and U4286 (N_4286,N_4162,N_4124);
and U4287 (N_4287,N_4197,N_4088);
nor U4288 (N_4288,N_3916,N_4013);
and U4289 (N_4289,N_4016,N_3949);
or U4290 (N_4290,N_4103,N_3918);
and U4291 (N_4291,N_4041,N_4048);
nand U4292 (N_4292,N_4189,N_4192);
nor U4293 (N_4293,N_3980,N_4121);
nand U4294 (N_4294,N_4042,N_4035);
xor U4295 (N_4295,N_3951,N_4015);
and U4296 (N_4296,N_3965,N_4061);
and U4297 (N_4297,N_4132,N_4117);
and U4298 (N_4298,N_3992,N_4019);
xor U4299 (N_4299,N_4057,N_4159);
nor U4300 (N_4300,N_4104,N_4118);
nor U4301 (N_4301,N_4175,N_4053);
nand U4302 (N_4302,N_4058,N_4154);
xnor U4303 (N_4303,N_3990,N_4199);
xor U4304 (N_4304,N_3972,N_4155);
and U4305 (N_4305,N_3981,N_3968);
and U4306 (N_4306,N_4007,N_4010);
nor U4307 (N_4307,N_4181,N_3944);
nand U4308 (N_4308,N_4135,N_4075);
nand U4309 (N_4309,N_4017,N_4090);
xor U4310 (N_4310,N_3905,N_4111);
nor U4311 (N_4311,N_4151,N_4062);
or U4312 (N_4312,N_4098,N_3958);
xor U4313 (N_4313,N_3925,N_3917);
nor U4314 (N_4314,N_4109,N_4049);
nor U4315 (N_4315,N_4166,N_4008);
xor U4316 (N_4316,N_3900,N_3983);
nand U4317 (N_4317,N_4110,N_3940);
or U4318 (N_4318,N_4165,N_3903);
or U4319 (N_4319,N_3932,N_3952);
and U4320 (N_4320,N_4143,N_4001);
or U4321 (N_4321,N_3912,N_4158);
xor U4322 (N_4322,N_4004,N_3976);
and U4323 (N_4323,N_4172,N_4095);
xnor U4324 (N_4324,N_4051,N_4147);
nand U4325 (N_4325,N_3950,N_3901);
xnor U4326 (N_4326,N_4097,N_3911);
nand U4327 (N_4327,N_4161,N_3931);
xnor U4328 (N_4328,N_3985,N_4139);
and U4329 (N_4329,N_4000,N_4003);
nor U4330 (N_4330,N_4087,N_3973);
nor U4331 (N_4331,N_4094,N_4180);
xor U4332 (N_4332,N_4064,N_3956);
nor U4333 (N_4333,N_4059,N_3961);
nand U4334 (N_4334,N_3963,N_3946);
xnor U4335 (N_4335,N_4085,N_4073);
nor U4336 (N_4336,N_4091,N_4030);
nand U4337 (N_4337,N_4024,N_4101);
nor U4338 (N_4338,N_4190,N_4025);
nor U4339 (N_4339,N_4046,N_4070);
nand U4340 (N_4340,N_4047,N_3919);
and U4341 (N_4341,N_3969,N_4036);
xnor U4342 (N_4342,N_4187,N_4080);
xor U4343 (N_4343,N_4115,N_4055);
nor U4344 (N_4344,N_4131,N_4119);
xor U4345 (N_4345,N_3994,N_4096);
or U4346 (N_4346,N_4168,N_4078);
nand U4347 (N_4347,N_4148,N_4195);
or U4348 (N_4348,N_4171,N_3924);
xor U4349 (N_4349,N_4034,N_3941);
xor U4350 (N_4350,N_4195,N_4161);
nor U4351 (N_4351,N_3941,N_4016);
or U4352 (N_4352,N_4005,N_4191);
xnor U4353 (N_4353,N_3962,N_4164);
and U4354 (N_4354,N_4120,N_3995);
and U4355 (N_4355,N_4094,N_3905);
and U4356 (N_4356,N_4148,N_4035);
or U4357 (N_4357,N_3952,N_3976);
or U4358 (N_4358,N_4053,N_3945);
or U4359 (N_4359,N_3904,N_4184);
nor U4360 (N_4360,N_3969,N_3923);
or U4361 (N_4361,N_4159,N_4007);
or U4362 (N_4362,N_3971,N_3959);
nor U4363 (N_4363,N_4090,N_4093);
nand U4364 (N_4364,N_4146,N_4188);
nor U4365 (N_4365,N_3912,N_3970);
or U4366 (N_4366,N_4018,N_3928);
xnor U4367 (N_4367,N_4166,N_4192);
or U4368 (N_4368,N_4106,N_3941);
nor U4369 (N_4369,N_3907,N_3975);
nor U4370 (N_4370,N_4018,N_4099);
nand U4371 (N_4371,N_4024,N_4027);
xor U4372 (N_4372,N_4039,N_4132);
or U4373 (N_4373,N_4136,N_4160);
nor U4374 (N_4374,N_3986,N_4160);
xor U4375 (N_4375,N_4167,N_4017);
nor U4376 (N_4376,N_4147,N_4141);
and U4377 (N_4377,N_4098,N_4083);
and U4378 (N_4378,N_4007,N_4034);
nor U4379 (N_4379,N_4150,N_4005);
or U4380 (N_4380,N_4140,N_4135);
nand U4381 (N_4381,N_4119,N_4157);
xnor U4382 (N_4382,N_4138,N_3927);
xnor U4383 (N_4383,N_3947,N_4095);
or U4384 (N_4384,N_3947,N_4023);
and U4385 (N_4385,N_4047,N_4143);
or U4386 (N_4386,N_3964,N_4166);
nand U4387 (N_4387,N_4048,N_4087);
nand U4388 (N_4388,N_4182,N_3915);
nand U4389 (N_4389,N_4025,N_3950);
or U4390 (N_4390,N_4162,N_3979);
nor U4391 (N_4391,N_4152,N_4014);
and U4392 (N_4392,N_4023,N_4038);
nand U4393 (N_4393,N_3931,N_4025);
or U4394 (N_4394,N_3939,N_4143);
nand U4395 (N_4395,N_4087,N_3924);
nor U4396 (N_4396,N_3949,N_4091);
nor U4397 (N_4397,N_3925,N_4055);
or U4398 (N_4398,N_3920,N_3950);
nor U4399 (N_4399,N_4064,N_4145);
nand U4400 (N_4400,N_4009,N_4072);
nor U4401 (N_4401,N_4084,N_4072);
and U4402 (N_4402,N_3969,N_3905);
or U4403 (N_4403,N_4122,N_4178);
nor U4404 (N_4404,N_3958,N_3922);
nor U4405 (N_4405,N_4083,N_4139);
nand U4406 (N_4406,N_4094,N_4185);
xor U4407 (N_4407,N_4143,N_3991);
or U4408 (N_4408,N_3922,N_4164);
and U4409 (N_4409,N_4167,N_4189);
nor U4410 (N_4410,N_4029,N_4051);
nand U4411 (N_4411,N_4143,N_4061);
and U4412 (N_4412,N_3969,N_4028);
nand U4413 (N_4413,N_3984,N_4018);
nor U4414 (N_4414,N_4187,N_4052);
nand U4415 (N_4415,N_4088,N_4022);
and U4416 (N_4416,N_3999,N_4021);
or U4417 (N_4417,N_4020,N_4058);
nand U4418 (N_4418,N_4041,N_3984);
nor U4419 (N_4419,N_4176,N_4008);
xnor U4420 (N_4420,N_4052,N_4182);
nor U4421 (N_4421,N_4008,N_4189);
xnor U4422 (N_4422,N_4012,N_4147);
xor U4423 (N_4423,N_3907,N_4077);
and U4424 (N_4424,N_4058,N_4059);
or U4425 (N_4425,N_4069,N_4173);
nor U4426 (N_4426,N_3981,N_4047);
and U4427 (N_4427,N_3977,N_3947);
nor U4428 (N_4428,N_3935,N_4161);
or U4429 (N_4429,N_4133,N_4173);
nand U4430 (N_4430,N_4007,N_4000);
xor U4431 (N_4431,N_4168,N_3947);
nor U4432 (N_4432,N_4089,N_4046);
nand U4433 (N_4433,N_4085,N_3938);
nand U4434 (N_4434,N_4059,N_4067);
nand U4435 (N_4435,N_4197,N_4020);
xnor U4436 (N_4436,N_4072,N_4079);
nand U4437 (N_4437,N_4004,N_4119);
or U4438 (N_4438,N_4131,N_4137);
or U4439 (N_4439,N_4130,N_4072);
or U4440 (N_4440,N_4193,N_4010);
xnor U4441 (N_4441,N_4135,N_3936);
and U4442 (N_4442,N_3978,N_4016);
or U4443 (N_4443,N_4182,N_4143);
nand U4444 (N_4444,N_4016,N_4108);
nor U4445 (N_4445,N_4095,N_3912);
nor U4446 (N_4446,N_4053,N_4110);
and U4447 (N_4447,N_4036,N_4116);
and U4448 (N_4448,N_3950,N_4147);
or U4449 (N_4449,N_4041,N_4004);
and U4450 (N_4450,N_3947,N_3926);
and U4451 (N_4451,N_3931,N_4162);
nor U4452 (N_4452,N_4141,N_3912);
nand U4453 (N_4453,N_3940,N_4170);
or U4454 (N_4454,N_3953,N_4021);
or U4455 (N_4455,N_4193,N_4060);
and U4456 (N_4456,N_4117,N_3961);
nor U4457 (N_4457,N_4004,N_4142);
nor U4458 (N_4458,N_4168,N_3911);
or U4459 (N_4459,N_3942,N_4183);
xor U4460 (N_4460,N_4123,N_4033);
and U4461 (N_4461,N_4145,N_4005);
or U4462 (N_4462,N_3953,N_4043);
nand U4463 (N_4463,N_4050,N_4132);
and U4464 (N_4464,N_3964,N_3938);
xor U4465 (N_4465,N_4063,N_4102);
nand U4466 (N_4466,N_3997,N_3974);
xnor U4467 (N_4467,N_4055,N_3946);
or U4468 (N_4468,N_4064,N_4104);
nand U4469 (N_4469,N_3912,N_3915);
nor U4470 (N_4470,N_4115,N_3967);
and U4471 (N_4471,N_3906,N_3929);
and U4472 (N_4472,N_3911,N_3905);
nor U4473 (N_4473,N_4141,N_4035);
xnor U4474 (N_4474,N_3994,N_4015);
xor U4475 (N_4475,N_3979,N_3916);
xor U4476 (N_4476,N_4052,N_4115);
nand U4477 (N_4477,N_3936,N_4006);
and U4478 (N_4478,N_4146,N_3969);
nand U4479 (N_4479,N_3927,N_3939);
xnor U4480 (N_4480,N_4170,N_4191);
or U4481 (N_4481,N_3985,N_4077);
and U4482 (N_4482,N_4055,N_4122);
and U4483 (N_4483,N_4016,N_3975);
and U4484 (N_4484,N_4191,N_4151);
nor U4485 (N_4485,N_3924,N_4020);
or U4486 (N_4486,N_4129,N_4177);
or U4487 (N_4487,N_4084,N_3927);
or U4488 (N_4488,N_4138,N_3982);
and U4489 (N_4489,N_3980,N_4118);
or U4490 (N_4490,N_4144,N_4087);
nor U4491 (N_4491,N_4095,N_4139);
and U4492 (N_4492,N_4122,N_3985);
nor U4493 (N_4493,N_3999,N_4155);
xnor U4494 (N_4494,N_4181,N_4011);
nand U4495 (N_4495,N_3948,N_4022);
or U4496 (N_4496,N_3986,N_3982);
nand U4497 (N_4497,N_3999,N_3928);
nand U4498 (N_4498,N_4004,N_4081);
xnor U4499 (N_4499,N_4188,N_4017);
and U4500 (N_4500,N_4289,N_4438);
or U4501 (N_4501,N_4445,N_4277);
or U4502 (N_4502,N_4399,N_4215);
nand U4503 (N_4503,N_4404,N_4390);
nand U4504 (N_4504,N_4379,N_4315);
nand U4505 (N_4505,N_4260,N_4381);
and U4506 (N_4506,N_4339,N_4374);
and U4507 (N_4507,N_4240,N_4375);
nor U4508 (N_4508,N_4239,N_4410);
xnor U4509 (N_4509,N_4452,N_4446);
or U4510 (N_4510,N_4456,N_4286);
and U4511 (N_4511,N_4394,N_4480);
or U4512 (N_4512,N_4376,N_4494);
or U4513 (N_4513,N_4299,N_4405);
nand U4514 (N_4514,N_4217,N_4397);
and U4515 (N_4515,N_4245,N_4327);
and U4516 (N_4516,N_4280,N_4499);
or U4517 (N_4517,N_4326,N_4235);
xor U4518 (N_4518,N_4265,N_4242);
and U4519 (N_4519,N_4443,N_4266);
nand U4520 (N_4520,N_4343,N_4473);
or U4521 (N_4521,N_4284,N_4457);
xor U4522 (N_4522,N_4449,N_4264);
xor U4523 (N_4523,N_4487,N_4482);
and U4524 (N_4524,N_4303,N_4252);
nor U4525 (N_4525,N_4477,N_4476);
nand U4526 (N_4526,N_4291,N_4253);
or U4527 (N_4527,N_4391,N_4305);
xor U4528 (N_4528,N_4454,N_4232);
or U4529 (N_4529,N_4226,N_4358);
nor U4530 (N_4530,N_4488,N_4336);
xor U4531 (N_4531,N_4342,N_4356);
nand U4532 (N_4532,N_4436,N_4380);
nor U4533 (N_4533,N_4371,N_4203);
nor U4534 (N_4534,N_4248,N_4442);
and U4535 (N_4535,N_4278,N_4366);
nor U4536 (N_4536,N_4218,N_4311);
nand U4537 (N_4537,N_4316,N_4431);
xor U4538 (N_4538,N_4200,N_4417);
nor U4539 (N_4539,N_4341,N_4418);
or U4540 (N_4540,N_4261,N_4302);
xnor U4541 (N_4541,N_4458,N_4415);
nand U4542 (N_4542,N_4466,N_4227);
xor U4543 (N_4543,N_4257,N_4497);
nand U4544 (N_4544,N_4401,N_4396);
and U4545 (N_4545,N_4387,N_4212);
nand U4546 (N_4546,N_4292,N_4463);
or U4547 (N_4547,N_4223,N_4451);
or U4548 (N_4548,N_4484,N_4392);
xnor U4549 (N_4549,N_4495,N_4268);
nand U4550 (N_4550,N_4414,N_4363);
or U4551 (N_4551,N_4453,N_4350);
nand U4552 (N_4552,N_4238,N_4309);
and U4553 (N_4553,N_4330,N_4262);
or U4554 (N_4554,N_4283,N_4447);
nor U4555 (N_4555,N_4352,N_4307);
or U4556 (N_4556,N_4317,N_4498);
xor U4557 (N_4557,N_4409,N_4353);
nand U4558 (N_4558,N_4419,N_4365);
xnor U4559 (N_4559,N_4279,N_4472);
and U4560 (N_4560,N_4301,N_4259);
xnor U4561 (N_4561,N_4355,N_4398);
xor U4562 (N_4562,N_4430,N_4220);
and U4563 (N_4563,N_4205,N_4389);
xor U4564 (N_4564,N_4319,N_4273);
or U4565 (N_4565,N_4496,N_4294);
xor U4566 (N_4566,N_4288,N_4337);
or U4567 (N_4567,N_4403,N_4439);
nand U4568 (N_4568,N_4465,N_4441);
xor U4569 (N_4569,N_4360,N_4384);
or U4570 (N_4570,N_4271,N_4471);
nand U4571 (N_4571,N_4435,N_4335);
xnor U4572 (N_4572,N_4267,N_4256);
nor U4573 (N_4573,N_4493,N_4450);
nor U4574 (N_4574,N_4462,N_4386);
and U4575 (N_4575,N_4269,N_4272);
xnor U4576 (N_4576,N_4425,N_4400);
xor U4577 (N_4577,N_4479,N_4328);
nor U4578 (N_4578,N_4312,N_4385);
nand U4579 (N_4579,N_4408,N_4411);
nor U4580 (N_4580,N_4448,N_4306);
or U4581 (N_4581,N_4320,N_4346);
nand U4582 (N_4582,N_4333,N_4206);
nand U4583 (N_4583,N_4370,N_4334);
nor U4584 (N_4584,N_4444,N_4427);
nand U4585 (N_4585,N_4491,N_4244);
xor U4586 (N_4586,N_4347,N_4406);
or U4587 (N_4587,N_4323,N_4331);
nor U4588 (N_4588,N_4231,N_4393);
or U4589 (N_4589,N_4359,N_4221);
nor U4590 (N_4590,N_4470,N_4233);
and U4591 (N_4591,N_4383,N_4255);
and U4592 (N_4592,N_4377,N_4300);
and U4593 (N_4593,N_4219,N_4357);
and U4594 (N_4594,N_4354,N_4237);
nand U4595 (N_4595,N_4468,N_4481);
nor U4596 (N_4596,N_4422,N_4276);
nor U4597 (N_4597,N_4246,N_4251);
nand U4598 (N_4598,N_4367,N_4423);
xnor U4599 (N_4599,N_4369,N_4426);
and U4600 (N_4600,N_4459,N_4329);
or U4601 (N_4601,N_4213,N_4361);
xnor U4602 (N_4602,N_4424,N_4208);
nand U4603 (N_4603,N_4460,N_4432);
xnor U4604 (N_4604,N_4467,N_4314);
and U4605 (N_4605,N_4372,N_4204);
nor U4606 (N_4606,N_4407,N_4464);
and U4607 (N_4607,N_4373,N_4348);
or U4608 (N_4608,N_4247,N_4485);
and U4609 (N_4609,N_4338,N_4402);
nand U4610 (N_4610,N_4270,N_4388);
and U4611 (N_4611,N_4413,N_4428);
nand U4612 (N_4612,N_4322,N_4275);
nand U4613 (N_4613,N_4475,N_4321);
xor U4614 (N_4614,N_4201,N_4224);
nand U4615 (N_4615,N_4304,N_4281);
xor U4616 (N_4616,N_4416,N_4230);
or U4617 (N_4617,N_4461,N_4297);
and U4618 (N_4618,N_4296,N_4455);
and U4619 (N_4619,N_4349,N_4282);
nor U4620 (N_4620,N_4258,N_4243);
and U4621 (N_4621,N_4351,N_4249);
and U4622 (N_4622,N_4313,N_4395);
nand U4623 (N_4623,N_4324,N_4241);
and U4624 (N_4624,N_4483,N_4474);
or U4625 (N_4625,N_4214,N_4437);
xnor U4626 (N_4626,N_4234,N_4378);
nor U4627 (N_4627,N_4364,N_4202);
xor U4628 (N_4628,N_4216,N_4382);
nand U4629 (N_4629,N_4325,N_4228);
xnor U4630 (N_4630,N_4263,N_4222);
nor U4631 (N_4631,N_4368,N_4344);
and U4632 (N_4632,N_4421,N_4229);
nand U4633 (N_4633,N_4254,N_4236);
xor U4634 (N_4634,N_4345,N_4429);
or U4635 (N_4635,N_4285,N_4490);
or U4636 (N_4636,N_4340,N_4211);
nor U4637 (N_4637,N_4207,N_4318);
nor U4638 (N_4638,N_4420,N_4287);
nor U4639 (N_4639,N_4308,N_4250);
nor U4640 (N_4640,N_4290,N_4293);
or U4641 (N_4641,N_4210,N_4492);
nand U4642 (N_4642,N_4412,N_4332);
xor U4643 (N_4643,N_4469,N_4274);
nand U4644 (N_4644,N_4362,N_4433);
or U4645 (N_4645,N_4298,N_4209);
nor U4646 (N_4646,N_4489,N_4310);
xnor U4647 (N_4647,N_4478,N_4295);
and U4648 (N_4648,N_4440,N_4434);
nor U4649 (N_4649,N_4486,N_4225);
nor U4650 (N_4650,N_4366,N_4279);
nor U4651 (N_4651,N_4423,N_4460);
and U4652 (N_4652,N_4399,N_4390);
nand U4653 (N_4653,N_4482,N_4266);
xor U4654 (N_4654,N_4396,N_4342);
and U4655 (N_4655,N_4414,N_4294);
xnor U4656 (N_4656,N_4322,N_4350);
xor U4657 (N_4657,N_4242,N_4250);
xnor U4658 (N_4658,N_4206,N_4478);
nand U4659 (N_4659,N_4445,N_4256);
nand U4660 (N_4660,N_4343,N_4321);
and U4661 (N_4661,N_4310,N_4473);
nor U4662 (N_4662,N_4272,N_4207);
xor U4663 (N_4663,N_4330,N_4391);
or U4664 (N_4664,N_4478,N_4486);
nor U4665 (N_4665,N_4364,N_4345);
nand U4666 (N_4666,N_4300,N_4253);
and U4667 (N_4667,N_4390,N_4415);
and U4668 (N_4668,N_4221,N_4369);
xor U4669 (N_4669,N_4248,N_4404);
nand U4670 (N_4670,N_4433,N_4274);
and U4671 (N_4671,N_4444,N_4374);
nand U4672 (N_4672,N_4285,N_4368);
and U4673 (N_4673,N_4251,N_4410);
nand U4674 (N_4674,N_4458,N_4432);
or U4675 (N_4675,N_4261,N_4425);
nor U4676 (N_4676,N_4295,N_4456);
nor U4677 (N_4677,N_4491,N_4354);
and U4678 (N_4678,N_4255,N_4382);
or U4679 (N_4679,N_4372,N_4364);
nand U4680 (N_4680,N_4437,N_4470);
nand U4681 (N_4681,N_4325,N_4416);
xor U4682 (N_4682,N_4351,N_4364);
or U4683 (N_4683,N_4455,N_4316);
or U4684 (N_4684,N_4344,N_4469);
xor U4685 (N_4685,N_4463,N_4436);
or U4686 (N_4686,N_4388,N_4252);
nand U4687 (N_4687,N_4408,N_4374);
nor U4688 (N_4688,N_4412,N_4364);
nand U4689 (N_4689,N_4365,N_4251);
and U4690 (N_4690,N_4302,N_4272);
and U4691 (N_4691,N_4276,N_4362);
xnor U4692 (N_4692,N_4263,N_4441);
nor U4693 (N_4693,N_4375,N_4402);
and U4694 (N_4694,N_4435,N_4307);
xnor U4695 (N_4695,N_4309,N_4326);
nor U4696 (N_4696,N_4224,N_4350);
or U4697 (N_4697,N_4215,N_4258);
or U4698 (N_4698,N_4385,N_4224);
and U4699 (N_4699,N_4335,N_4330);
or U4700 (N_4700,N_4369,N_4252);
nand U4701 (N_4701,N_4237,N_4476);
or U4702 (N_4702,N_4304,N_4228);
xor U4703 (N_4703,N_4363,N_4298);
nand U4704 (N_4704,N_4311,N_4366);
or U4705 (N_4705,N_4456,N_4461);
nor U4706 (N_4706,N_4322,N_4441);
or U4707 (N_4707,N_4441,N_4359);
xor U4708 (N_4708,N_4422,N_4495);
nand U4709 (N_4709,N_4472,N_4310);
or U4710 (N_4710,N_4433,N_4490);
and U4711 (N_4711,N_4384,N_4368);
xor U4712 (N_4712,N_4494,N_4285);
and U4713 (N_4713,N_4322,N_4266);
nor U4714 (N_4714,N_4362,N_4454);
nand U4715 (N_4715,N_4230,N_4355);
or U4716 (N_4716,N_4222,N_4331);
nor U4717 (N_4717,N_4250,N_4481);
xor U4718 (N_4718,N_4425,N_4366);
xor U4719 (N_4719,N_4315,N_4461);
nor U4720 (N_4720,N_4308,N_4273);
or U4721 (N_4721,N_4459,N_4359);
or U4722 (N_4722,N_4369,N_4393);
nor U4723 (N_4723,N_4316,N_4372);
nor U4724 (N_4724,N_4285,N_4205);
nand U4725 (N_4725,N_4489,N_4378);
nor U4726 (N_4726,N_4498,N_4440);
xor U4727 (N_4727,N_4471,N_4465);
xor U4728 (N_4728,N_4423,N_4383);
nand U4729 (N_4729,N_4457,N_4438);
xnor U4730 (N_4730,N_4386,N_4459);
or U4731 (N_4731,N_4475,N_4415);
nand U4732 (N_4732,N_4481,N_4406);
nor U4733 (N_4733,N_4283,N_4246);
xor U4734 (N_4734,N_4236,N_4423);
nor U4735 (N_4735,N_4201,N_4312);
xnor U4736 (N_4736,N_4328,N_4487);
and U4737 (N_4737,N_4215,N_4275);
and U4738 (N_4738,N_4440,N_4315);
nand U4739 (N_4739,N_4210,N_4458);
nand U4740 (N_4740,N_4311,N_4265);
xor U4741 (N_4741,N_4439,N_4252);
nor U4742 (N_4742,N_4394,N_4352);
nand U4743 (N_4743,N_4341,N_4245);
xor U4744 (N_4744,N_4220,N_4382);
nor U4745 (N_4745,N_4250,N_4214);
or U4746 (N_4746,N_4262,N_4465);
nor U4747 (N_4747,N_4465,N_4430);
nand U4748 (N_4748,N_4413,N_4317);
or U4749 (N_4749,N_4489,N_4275);
and U4750 (N_4750,N_4379,N_4435);
or U4751 (N_4751,N_4207,N_4405);
xnor U4752 (N_4752,N_4253,N_4337);
nand U4753 (N_4753,N_4224,N_4444);
nand U4754 (N_4754,N_4449,N_4322);
nor U4755 (N_4755,N_4478,N_4402);
or U4756 (N_4756,N_4243,N_4266);
nand U4757 (N_4757,N_4469,N_4452);
and U4758 (N_4758,N_4389,N_4243);
or U4759 (N_4759,N_4314,N_4224);
nor U4760 (N_4760,N_4367,N_4312);
and U4761 (N_4761,N_4300,N_4432);
nand U4762 (N_4762,N_4422,N_4402);
xnor U4763 (N_4763,N_4467,N_4380);
xor U4764 (N_4764,N_4393,N_4237);
nand U4765 (N_4765,N_4468,N_4203);
or U4766 (N_4766,N_4444,N_4415);
or U4767 (N_4767,N_4436,N_4275);
and U4768 (N_4768,N_4366,N_4265);
nand U4769 (N_4769,N_4464,N_4429);
nand U4770 (N_4770,N_4418,N_4484);
xnor U4771 (N_4771,N_4234,N_4461);
and U4772 (N_4772,N_4347,N_4305);
nand U4773 (N_4773,N_4487,N_4457);
nor U4774 (N_4774,N_4275,N_4226);
xnor U4775 (N_4775,N_4440,N_4212);
xor U4776 (N_4776,N_4272,N_4432);
nand U4777 (N_4777,N_4301,N_4461);
and U4778 (N_4778,N_4293,N_4224);
xnor U4779 (N_4779,N_4371,N_4387);
nand U4780 (N_4780,N_4367,N_4378);
nand U4781 (N_4781,N_4374,N_4235);
and U4782 (N_4782,N_4244,N_4295);
and U4783 (N_4783,N_4333,N_4229);
nand U4784 (N_4784,N_4366,N_4457);
nor U4785 (N_4785,N_4313,N_4351);
xor U4786 (N_4786,N_4347,N_4374);
nand U4787 (N_4787,N_4347,N_4270);
or U4788 (N_4788,N_4364,N_4459);
or U4789 (N_4789,N_4437,N_4269);
nor U4790 (N_4790,N_4217,N_4307);
xnor U4791 (N_4791,N_4314,N_4222);
nor U4792 (N_4792,N_4321,N_4469);
nand U4793 (N_4793,N_4233,N_4226);
and U4794 (N_4794,N_4213,N_4390);
xor U4795 (N_4795,N_4498,N_4379);
nand U4796 (N_4796,N_4243,N_4319);
xor U4797 (N_4797,N_4386,N_4240);
nand U4798 (N_4798,N_4458,N_4427);
and U4799 (N_4799,N_4455,N_4476);
or U4800 (N_4800,N_4797,N_4708);
nor U4801 (N_4801,N_4678,N_4647);
nor U4802 (N_4802,N_4666,N_4706);
or U4803 (N_4803,N_4560,N_4772);
nand U4804 (N_4804,N_4684,N_4532);
xnor U4805 (N_4805,N_4509,N_4661);
xnor U4806 (N_4806,N_4612,N_4773);
xnor U4807 (N_4807,N_4575,N_4671);
xnor U4808 (N_4808,N_4534,N_4585);
or U4809 (N_4809,N_4637,N_4528);
nor U4810 (N_4810,N_4531,N_4530);
nand U4811 (N_4811,N_4511,N_4595);
nor U4812 (N_4812,N_4655,N_4710);
nor U4813 (N_4813,N_4519,N_4747);
nor U4814 (N_4814,N_4593,N_4728);
xor U4815 (N_4815,N_4787,N_4729);
or U4816 (N_4816,N_4604,N_4645);
and U4817 (N_4817,N_4626,N_4611);
xnor U4818 (N_4818,N_4629,N_4759);
nand U4819 (N_4819,N_4529,N_4641);
nand U4820 (N_4820,N_4658,N_4725);
or U4821 (N_4821,N_4798,N_4781);
nand U4822 (N_4822,N_4712,N_4685);
xnor U4823 (N_4823,N_4619,N_4782);
and U4824 (N_4824,N_4628,N_4724);
nand U4825 (N_4825,N_4714,N_4700);
xor U4826 (N_4826,N_4523,N_4635);
and U4827 (N_4827,N_4646,N_4653);
or U4828 (N_4828,N_4587,N_4761);
nor U4829 (N_4829,N_4561,N_4766);
and U4830 (N_4830,N_4662,N_4721);
xnor U4831 (N_4831,N_4640,N_4506);
and U4832 (N_4832,N_4623,N_4672);
xor U4833 (N_4833,N_4794,N_4517);
xor U4834 (N_4834,N_4715,N_4664);
or U4835 (N_4835,N_4631,N_4739);
and U4836 (N_4836,N_4775,N_4636);
xor U4837 (N_4837,N_4756,N_4581);
nor U4838 (N_4838,N_4745,N_4736);
nor U4839 (N_4839,N_4771,N_4633);
and U4840 (N_4840,N_4525,N_4565);
and U4841 (N_4841,N_4608,N_4606);
xnor U4842 (N_4842,N_4770,N_4702);
and U4843 (N_4843,N_4505,N_4597);
xor U4844 (N_4844,N_4716,N_4768);
and U4845 (N_4845,N_4727,N_4624);
and U4846 (N_4846,N_4555,N_4546);
or U4847 (N_4847,N_4785,N_4726);
nand U4848 (N_4848,N_4699,N_4669);
xor U4849 (N_4849,N_4730,N_4746);
xnor U4850 (N_4850,N_4676,N_4796);
xnor U4851 (N_4851,N_4535,N_4694);
and U4852 (N_4852,N_4698,N_4570);
nand U4853 (N_4853,N_4731,N_4553);
nor U4854 (N_4854,N_4552,N_4690);
nor U4855 (N_4855,N_4639,N_4542);
nand U4856 (N_4856,N_4783,N_4568);
or U4857 (N_4857,N_4670,N_4737);
xnor U4858 (N_4858,N_4501,N_4757);
nor U4859 (N_4859,N_4650,N_4701);
xor U4860 (N_4860,N_4563,N_4686);
xor U4861 (N_4861,N_4649,N_4742);
nor U4862 (N_4862,N_4679,N_4677);
nor U4863 (N_4863,N_4579,N_4668);
nor U4864 (N_4864,N_4614,N_4634);
xor U4865 (N_4865,N_4513,N_4516);
nor U4866 (N_4866,N_4704,N_4642);
xnor U4867 (N_4867,N_4550,N_4557);
and U4868 (N_4868,N_4718,N_4697);
nor U4869 (N_4869,N_4687,N_4691);
nor U4870 (N_4870,N_4693,N_4695);
or U4871 (N_4871,N_4682,N_4524);
nand U4872 (N_4872,N_4654,N_4776);
and U4873 (N_4873,N_4594,N_4507);
xor U4874 (N_4874,N_4564,N_4514);
and U4875 (N_4875,N_4765,N_4733);
or U4876 (N_4876,N_4567,N_4569);
and U4877 (N_4877,N_4589,N_4692);
and U4878 (N_4878,N_4738,N_4526);
nor U4879 (N_4879,N_4571,N_4707);
and U4880 (N_4880,N_4651,N_4625);
xnor U4881 (N_4881,N_4790,N_4777);
or U4882 (N_4882,N_4621,N_4543);
and U4883 (N_4883,N_4659,N_4675);
xnor U4884 (N_4884,N_4603,N_4780);
xor U4885 (N_4885,N_4591,N_4769);
nor U4886 (N_4886,N_4644,N_4763);
xnor U4887 (N_4887,N_4792,N_4610);
or U4888 (N_4888,N_4544,N_4599);
xor U4889 (N_4889,N_4627,N_4577);
and U4890 (N_4890,N_4576,N_4521);
xor U4891 (N_4891,N_4504,N_4598);
and U4892 (N_4892,N_4590,N_4774);
or U4893 (N_4893,N_4559,N_4795);
nor U4894 (N_4894,N_4788,N_4667);
nand U4895 (N_4895,N_4572,N_4566);
or U4896 (N_4896,N_4580,N_4749);
nor U4897 (N_4897,N_4503,N_4750);
xor U4898 (N_4898,N_4540,N_4784);
nand U4899 (N_4899,N_4615,N_4713);
nor U4900 (N_4900,N_4574,N_4789);
and U4901 (N_4901,N_4723,N_4538);
nor U4902 (N_4902,N_4793,N_4748);
and U4903 (N_4903,N_4510,N_4660);
nor U4904 (N_4904,N_4573,N_4630);
xnor U4905 (N_4905,N_4549,N_4512);
nand U4906 (N_4906,N_4681,N_4722);
and U4907 (N_4907,N_4734,N_4539);
xor U4908 (N_4908,N_4584,N_4583);
xor U4909 (N_4909,N_4717,N_4711);
or U4910 (N_4910,N_4764,N_4541);
nand U4911 (N_4911,N_4683,N_4720);
and U4912 (N_4912,N_4786,N_4663);
and U4913 (N_4913,N_4582,N_4588);
and U4914 (N_4914,N_4735,N_4609);
and U4915 (N_4915,N_4578,N_4547);
xnor U4916 (N_4916,N_4620,N_4502);
or U4917 (N_4917,N_4778,N_4508);
or U4918 (N_4918,N_4696,N_4741);
or U4919 (N_4919,N_4767,N_4703);
or U4920 (N_4920,N_4605,N_4613);
xnor U4921 (N_4921,N_4657,N_4536);
nor U4922 (N_4922,N_4751,N_4688);
nor U4923 (N_4923,N_4520,N_4622);
nand U4924 (N_4924,N_4616,N_4709);
or U4925 (N_4925,N_4545,N_4607);
xnor U4926 (N_4926,N_4558,N_4522);
or U4927 (N_4927,N_4500,N_4537);
xor U4928 (N_4928,N_4548,N_4648);
or U4929 (N_4929,N_4596,N_4719);
xnor U4930 (N_4930,N_4652,N_4779);
or U4931 (N_4931,N_4600,N_4760);
and U4932 (N_4932,N_4656,N_4518);
xnor U4933 (N_4933,N_4592,N_4732);
xor U4934 (N_4934,N_4527,N_4533);
xor U4935 (N_4935,N_4515,N_4643);
and U4936 (N_4936,N_4673,N_4740);
nor U4937 (N_4937,N_4743,N_4665);
nand U4938 (N_4938,N_4791,N_4617);
or U4939 (N_4939,N_4601,N_4689);
or U4940 (N_4940,N_4680,N_4554);
or U4941 (N_4941,N_4754,N_4618);
and U4942 (N_4942,N_4551,N_4762);
nand U4943 (N_4943,N_4744,N_4632);
and U4944 (N_4944,N_4755,N_4758);
xnor U4945 (N_4945,N_4602,N_4556);
and U4946 (N_4946,N_4752,N_4799);
and U4947 (N_4947,N_4638,N_4562);
or U4948 (N_4948,N_4674,N_4753);
xnor U4949 (N_4949,N_4705,N_4586);
xnor U4950 (N_4950,N_4583,N_4511);
nor U4951 (N_4951,N_4712,N_4798);
and U4952 (N_4952,N_4686,N_4507);
nor U4953 (N_4953,N_4755,N_4785);
nor U4954 (N_4954,N_4694,N_4538);
nor U4955 (N_4955,N_4559,N_4654);
xor U4956 (N_4956,N_4799,N_4606);
and U4957 (N_4957,N_4787,N_4771);
or U4958 (N_4958,N_4670,N_4760);
nor U4959 (N_4959,N_4731,N_4500);
or U4960 (N_4960,N_4769,N_4532);
nor U4961 (N_4961,N_4616,N_4556);
xnor U4962 (N_4962,N_4509,N_4570);
nor U4963 (N_4963,N_4787,N_4520);
nand U4964 (N_4964,N_4606,N_4740);
nor U4965 (N_4965,N_4659,N_4554);
xnor U4966 (N_4966,N_4635,N_4786);
nor U4967 (N_4967,N_4627,N_4792);
nor U4968 (N_4968,N_4696,N_4677);
or U4969 (N_4969,N_4640,N_4789);
nand U4970 (N_4970,N_4679,N_4716);
nand U4971 (N_4971,N_4786,N_4675);
and U4972 (N_4972,N_4666,N_4552);
nand U4973 (N_4973,N_4600,N_4553);
xor U4974 (N_4974,N_4614,N_4550);
and U4975 (N_4975,N_4785,N_4617);
nor U4976 (N_4976,N_4739,N_4781);
nor U4977 (N_4977,N_4698,N_4585);
or U4978 (N_4978,N_4506,N_4505);
or U4979 (N_4979,N_4635,N_4597);
xor U4980 (N_4980,N_4633,N_4774);
nor U4981 (N_4981,N_4581,N_4720);
nor U4982 (N_4982,N_4763,N_4607);
or U4983 (N_4983,N_4687,N_4755);
or U4984 (N_4984,N_4538,N_4522);
nor U4985 (N_4985,N_4602,N_4799);
nand U4986 (N_4986,N_4663,N_4535);
or U4987 (N_4987,N_4671,N_4780);
nor U4988 (N_4988,N_4725,N_4687);
nand U4989 (N_4989,N_4735,N_4797);
xor U4990 (N_4990,N_4704,N_4776);
or U4991 (N_4991,N_4698,N_4677);
nand U4992 (N_4992,N_4776,N_4528);
and U4993 (N_4993,N_4611,N_4687);
nor U4994 (N_4994,N_4740,N_4504);
xor U4995 (N_4995,N_4514,N_4761);
and U4996 (N_4996,N_4688,N_4538);
xor U4997 (N_4997,N_4547,N_4764);
xor U4998 (N_4998,N_4576,N_4556);
nand U4999 (N_4999,N_4768,N_4788);
xor U5000 (N_5000,N_4642,N_4677);
and U5001 (N_5001,N_4760,N_4588);
nor U5002 (N_5002,N_4639,N_4642);
xnor U5003 (N_5003,N_4585,N_4652);
or U5004 (N_5004,N_4584,N_4674);
nor U5005 (N_5005,N_4575,N_4735);
nand U5006 (N_5006,N_4516,N_4546);
and U5007 (N_5007,N_4763,N_4672);
nor U5008 (N_5008,N_4535,N_4612);
or U5009 (N_5009,N_4575,N_4621);
xnor U5010 (N_5010,N_4772,N_4717);
xnor U5011 (N_5011,N_4617,N_4716);
and U5012 (N_5012,N_4750,N_4680);
or U5013 (N_5013,N_4526,N_4713);
or U5014 (N_5014,N_4734,N_4789);
xnor U5015 (N_5015,N_4665,N_4790);
nand U5016 (N_5016,N_4724,N_4608);
nor U5017 (N_5017,N_4548,N_4689);
nand U5018 (N_5018,N_4653,N_4777);
or U5019 (N_5019,N_4536,N_4734);
and U5020 (N_5020,N_4770,N_4577);
nor U5021 (N_5021,N_4566,N_4696);
nand U5022 (N_5022,N_4600,N_4799);
or U5023 (N_5023,N_4660,N_4629);
or U5024 (N_5024,N_4502,N_4656);
and U5025 (N_5025,N_4780,N_4570);
nand U5026 (N_5026,N_4611,N_4760);
nor U5027 (N_5027,N_4618,N_4727);
or U5028 (N_5028,N_4508,N_4684);
nand U5029 (N_5029,N_4785,N_4741);
and U5030 (N_5030,N_4544,N_4716);
and U5031 (N_5031,N_4610,N_4592);
xor U5032 (N_5032,N_4502,N_4714);
and U5033 (N_5033,N_4757,N_4517);
nand U5034 (N_5034,N_4534,N_4663);
nand U5035 (N_5035,N_4689,N_4711);
xnor U5036 (N_5036,N_4509,N_4581);
and U5037 (N_5037,N_4795,N_4778);
nand U5038 (N_5038,N_4777,N_4708);
xnor U5039 (N_5039,N_4748,N_4693);
nand U5040 (N_5040,N_4644,N_4611);
or U5041 (N_5041,N_4727,N_4601);
and U5042 (N_5042,N_4725,N_4559);
nor U5043 (N_5043,N_4697,N_4598);
nand U5044 (N_5044,N_4642,N_4662);
xor U5045 (N_5045,N_4736,N_4655);
nand U5046 (N_5046,N_4763,N_4657);
nor U5047 (N_5047,N_4742,N_4708);
xor U5048 (N_5048,N_4587,N_4606);
xnor U5049 (N_5049,N_4651,N_4763);
xor U5050 (N_5050,N_4787,N_4668);
and U5051 (N_5051,N_4594,N_4751);
and U5052 (N_5052,N_4652,N_4753);
and U5053 (N_5053,N_4717,N_4550);
or U5054 (N_5054,N_4518,N_4524);
nor U5055 (N_5055,N_4648,N_4756);
or U5056 (N_5056,N_4517,N_4650);
nand U5057 (N_5057,N_4583,N_4789);
nor U5058 (N_5058,N_4593,N_4631);
nor U5059 (N_5059,N_4665,N_4779);
nor U5060 (N_5060,N_4712,N_4634);
and U5061 (N_5061,N_4700,N_4554);
nand U5062 (N_5062,N_4575,N_4796);
nor U5063 (N_5063,N_4649,N_4712);
and U5064 (N_5064,N_4533,N_4657);
nor U5065 (N_5065,N_4587,N_4531);
or U5066 (N_5066,N_4502,N_4516);
and U5067 (N_5067,N_4737,N_4651);
or U5068 (N_5068,N_4580,N_4657);
nand U5069 (N_5069,N_4514,N_4692);
and U5070 (N_5070,N_4667,N_4608);
nand U5071 (N_5071,N_4616,N_4711);
nor U5072 (N_5072,N_4641,N_4527);
nor U5073 (N_5073,N_4719,N_4565);
nand U5074 (N_5074,N_4544,N_4764);
or U5075 (N_5075,N_4641,N_4541);
nor U5076 (N_5076,N_4511,N_4562);
nand U5077 (N_5077,N_4780,N_4531);
or U5078 (N_5078,N_4737,N_4726);
xnor U5079 (N_5079,N_4712,N_4529);
xnor U5080 (N_5080,N_4690,N_4702);
or U5081 (N_5081,N_4574,N_4570);
or U5082 (N_5082,N_4743,N_4752);
xor U5083 (N_5083,N_4703,N_4505);
and U5084 (N_5084,N_4558,N_4680);
or U5085 (N_5085,N_4678,N_4618);
nor U5086 (N_5086,N_4676,N_4661);
nand U5087 (N_5087,N_4598,N_4562);
or U5088 (N_5088,N_4642,N_4730);
nand U5089 (N_5089,N_4722,N_4723);
nand U5090 (N_5090,N_4609,N_4672);
or U5091 (N_5091,N_4586,N_4679);
nor U5092 (N_5092,N_4533,N_4550);
or U5093 (N_5093,N_4765,N_4631);
nor U5094 (N_5094,N_4554,N_4719);
xor U5095 (N_5095,N_4771,N_4716);
nand U5096 (N_5096,N_4754,N_4558);
and U5097 (N_5097,N_4521,N_4798);
nor U5098 (N_5098,N_4521,N_4714);
nor U5099 (N_5099,N_4612,N_4506);
nor U5100 (N_5100,N_5004,N_5020);
xor U5101 (N_5101,N_4947,N_5043);
and U5102 (N_5102,N_4981,N_4854);
nand U5103 (N_5103,N_4980,N_5016);
nor U5104 (N_5104,N_5014,N_4979);
nor U5105 (N_5105,N_5099,N_4826);
nor U5106 (N_5106,N_4823,N_4946);
xor U5107 (N_5107,N_4861,N_5056);
nor U5108 (N_5108,N_5076,N_4897);
or U5109 (N_5109,N_4887,N_4879);
nor U5110 (N_5110,N_4857,N_4840);
xor U5111 (N_5111,N_5002,N_5059);
and U5112 (N_5112,N_4881,N_4802);
nor U5113 (N_5113,N_5054,N_4808);
or U5114 (N_5114,N_4974,N_5079);
nor U5115 (N_5115,N_4984,N_5071);
or U5116 (N_5116,N_5049,N_4805);
nor U5117 (N_5117,N_5098,N_4912);
and U5118 (N_5118,N_4916,N_4999);
xor U5119 (N_5119,N_4870,N_4875);
and U5120 (N_5120,N_4913,N_4819);
nor U5121 (N_5121,N_5025,N_4859);
nand U5122 (N_5122,N_5035,N_4919);
nand U5123 (N_5123,N_5068,N_4872);
xnor U5124 (N_5124,N_4934,N_4945);
xor U5125 (N_5125,N_4830,N_4853);
nand U5126 (N_5126,N_4836,N_4973);
or U5127 (N_5127,N_4824,N_4977);
nor U5128 (N_5128,N_5042,N_4894);
or U5129 (N_5129,N_4993,N_4917);
or U5130 (N_5130,N_4985,N_4860);
nand U5131 (N_5131,N_5073,N_4991);
nand U5132 (N_5132,N_4965,N_4856);
xor U5133 (N_5133,N_4890,N_4838);
and U5134 (N_5134,N_4882,N_4992);
or U5135 (N_5135,N_4904,N_4954);
nand U5136 (N_5136,N_5061,N_4800);
nand U5137 (N_5137,N_4978,N_5069);
and U5138 (N_5138,N_5058,N_5087);
nand U5139 (N_5139,N_5015,N_5018);
nor U5140 (N_5140,N_5096,N_4814);
nor U5141 (N_5141,N_4813,N_4982);
or U5142 (N_5142,N_5036,N_4817);
and U5143 (N_5143,N_5041,N_5029);
xnor U5144 (N_5144,N_4943,N_5037);
or U5145 (N_5145,N_4833,N_4848);
or U5146 (N_5146,N_5011,N_4921);
nand U5147 (N_5147,N_4927,N_5050);
nand U5148 (N_5148,N_4878,N_4987);
and U5149 (N_5149,N_4990,N_4818);
nor U5150 (N_5150,N_4914,N_4988);
xor U5151 (N_5151,N_4835,N_4806);
and U5152 (N_5152,N_5077,N_4936);
nor U5153 (N_5153,N_5009,N_5052);
nor U5154 (N_5154,N_4942,N_5083);
xor U5155 (N_5155,N_5026,N_5013);
or U5156 (N_5156,N_5092,N_5053);
nor U5157 (N_5157,N_4803,N_4962);
nor U5158 (N_5158,N_4901,N_5008);
nand U5159 (N_5159,N_4964,N_4995);
and U5160 (N_5160,N_4847,N_4828);
xor U5161 (N_5161,N_4972,N_5017);
or U5162 (N_5162,N_4834,N_4874);
nand U5163 (N_5163,N_5030,N_5031);
xnor U5164 (N_5164,N_5046,N_5048);
nor U5165 (N_5165,N_4967,N_5062);
or U5166 (N_5166,N_4850,N_4843);
xnor U5167 (N_5167,N_5074,N_5097);
xnor U5168 (N_5168,N_5078,N_4825);
nor U5169 (N_5169,N_4829,N_4845);
nor U5170 (N_5170,N_4876,N_4944);
nand U5171 (N_5171,N_4996,N_4810);
nor U5172 (N_5172,N_4948,N_4905);
or U5173 (N_5173,N_4966,N_4846);
or U5174 (N_5174,N_5090,N_4832);
and U5175 (N_5175,N_4883,N_4940);
and U5176 (N_5176,N_5024,N_5040);
xnor U5177 (N_5177,N_4893,N_4938);
and U5178 (N_5178,N_5051,N_4997);
nor U5179 (N_5179,N_4931,N_4935);
nand U5180 (N_5180,N_4820,N_4900);
nor U5181 (N_5181,N_4960,N_4892);
or U5182 (N_5182,N_5019,N_5003);
or U5183 (N_5183,N_4867,N_4852);
xor U5184 (N_5184,N_4811,N_4831);
xnor U5185 (N_5185,N_4908,N_5063);
xnor U5186 (N_5186,N_4804,N_4949);
or U5187 (N_5187,N_4928,N_4841);
and U5188 (N_5188,N_4862,N_4815);
and U5189 (N_5189,N_4963,N_4986);
xor U5190 (N_5190,N_4923,N_5085);
nand U5191 (N_5191,N_4865,N_4961);
nand U5192 (N_5192,N_5022,N_5088);
xor U5193 (N_5193,N_4827,N_4971);
and U5194 (N_5194,N_5039,N_4816);
xnor U5195 (N_5195,N_4937,N_4842);
nand U5196 (N_5196,N_4920,N_4873);
xnor U5197 (N_5197,N_5086,N_4930);
nor U5198 (N_5198,N_4925,N_4998);
nand U5199 (N_5199,N_4933,N_4915);
and U5200 (N_5200,N_4958,N_4822);
nand U5201 (N_5201,N_4807,N_4871);
and U5202 (N_5202,N_5027,N_4896);
xor U5203 (N_5203,N_4863,N_4886);
xnor U5204 (N_5204,N_4821,N_4959);
and U5205 (N_5205,N_4951,N_5000);
xor U5206 (N_5206,N_5012,N_4910);
nor U5207 (N_5207,N_4922,N_5044);
or U5208 (N_5208,N_4911,N_5091);
nand U5209 (N_5209,N_4891,N_5093);
and U5210 (N_5210,N_5067,N_5089);
nand U5211 (N_5211,N_4812,N_4953);
and U5212 (N_5212,N_4955,N_4866);
nand U5213 (N_5213,N_4952,N_4864);
xnor U5214 (N_5214,N_5095,N_5033);
or U5215 (N_5215,N_5032,N_4903);
xnor U5216 (N_5216,N_4976,N_5047);
and U5217 (N_5217,N_4906,N_4924);
nand U5218 (N_5218,N_4844,N_4939);
nand U5219 (N_5219,N_4989,N_5007);
and U5220 (N_5220,N_4899,N_4918);
nand U5221 (N_5221,N_4889,N_4907);
and U5222 (N_5222,N_5045,N_5084);
nand U5223 (N_5223,N_5066,N_5057);
nand U5224 (N_5224,N_5075,N_5072);
nor U5225 (N_5225,N_4970,N_5028);
xor U5226 (N_5226,N_4969,N_4855);
or U5227 (N_5227,N_4868,N_4909);
and U5228 (N_5228,N_5005,N_5081);
and U5229 (N_5229,N_5064,N_4851);
or U5230 (N_5230,N_4837,N_4994);
nor U5231 (N_5231,N_5055,N_5065);
nor U5232 (N_5232,N_4869,N_5038);
nor U5233 (N_5233,N_4926,N_4929);
xnor U5234 (N_5234,N_4975,N_4809);
and U5235 (N_5235,N_4950,N_5070);
nor U5236 (N_5236,N_5034,N_5021);
or U5237 (N_5237,N_4849,N_4983);
xor U5238 (N_5238,N_4877,N_4941);
nand U5239 (N_5239,N_4885,N_4956);
nand U5240 (N_5240,N_4858,N_5060);
nand U5241 (N_5241,N_4801,N_4902);
nor U5242 (N_5242,N_4895,N_4888);
and U5243 (N_5243,N_4884,N_5080);
nor U5244 (N_5244,N_4880,N_4968);
nor U5245 (N_5245,N_4957,N_4932);
or U5246 (N_5246,N_5094,N_4839);
and U5247 (N_5247,N_4898,N_5001);
nand U5248 (N_5248,N_5023,N_5006);
nand U5249 (N_5249,N_5082,N_5010);
nand U5250 (N_5250,N_4879,N_4884);
and U5251 (N_5251,N_4875,N_4962);
and U5252 (N_5252,N_4975,N_5018);
or U5253 (N_5253,N_5080,N_4883);
and U5254 (N_5254,N_5001,N_4804);
nand U5255 (N_5255,N_4829,N_4912);
nor U5256 (N_5256,N_5063,N_5077);
xnor U5257 (N_5257,N_5053,N_4835);
or U5258 (N_5258,N_4804,N_5020);
or U5259 (N_5259,N_4831,N_4844);
nor U5260 (N_5260,N_4899,N_4955);
nor U5261 (N_5261,N_4946,N_5012);
xor U5262 (N_5262,N_4919,N_4985);
xnor U5263 (N_5263,N_4871,N_4932);
nand U5264 (N_5264,N_4810,N_4848);
or U5265 (N_5265,N_4819,N_4846);
and U5266 (N_5266,N_4816,N_4825);
or U5267 (N_5267,N_4834,N_4920);
and U5268 (N_5268,N_4963,N_4898);
nand U5269 (N_5269,N_5073,N_5019);
nand U5270 (N_5270,N_4928,N_4939);
xnor U5271 (N_5271,N_4808,N_4815);
or U5272 (N_5272,N_5090,N_5052);
nand U5273 (N_5273,N_4954,N_5016);
nor U5274 (N_5274,N_5016,N_5031);
and U5275 (N_5275,N_4878,N_5083);
xnor U5276 (N_5276,N_4886,N_4925);
nor U5277 (N_5277,N_4877,N_5058);
or U5278 (N_5278,N_4911,N_4910);
nor U5279 (N_5279,N_4921,N_5056);
and U5280 (N_5280,N_5042,N_5041);
xor U5281 (N_5281,N_4981,N_4940);
and U5282 (N_5282,N_5012,N_4937);
and U5283 (N_5283,N_4831,N_5022);
and U5284 (N_5284,N_5044,N_4821);
or U5285 (N_5285,N_4837,N_4818);
or U5286 (N_5286,N_5065,N_4882);
nor U5287 (N_5287,N_4979,N_4971);
or U5288 (N_5288,N_4867,N_5050);
xnor U5289 (N_5289,N_4844,N_4808);
nand U5290 (N_5290,N_5063,N_4809);
or U5291 (N_5291,N_4851,N_5028);
nand U5292 (N_5292,N_4856,N_5082);
or U5293 (N_5293,N_4831,N_4884);
or U5294 (N_5294,N_5021,N_4915);
or U5295 (N_5295,N_4991,N_4939);
xnor U5296 (N_5296,N_4827,N_4810);
xnor U5297 (N_5297,N_5062,N_5054);
and U5298 (N_5298,N_5038,N_4971);
xor U5299 (N_5299,N_4970,N_4953);
nand U5300 (N_5300,N_4836,N_4997);
or U5301 (N_5301,N_5048,N_5072);
xnor U5302 (N_5302,N_4939,N_5016);
xnor U5303 (N_5303,N_4911,N_4967);
and U5304 (N_5304,N_4974,N_4973);
nand U5305 (N_5305,N_5030,N_4849);
nor U5306 (N_5306,N_4938,N_4923);
xor U5307 (N_5307,N_4902,N_5066);
xnor U5308 (N_5308,N_4934,N_4871);
nor U5309 (N_5309,N_5087,N_4998);
or U5310 (N_5310,N_4989,N_5085);
or U5311 (N_5311,N_4966,N_4951);
and U5312 (N_5312,N_5038,N_5008);
nor U5313 (N_5313,N_4826,N_4805);
xor U5314 (N_5314,N_4990,N_4960);
nor U5315 (N_5315,N_5020,N_4914);
nand U5316 (N_5316,N_4967,N_4931);
or U5317 (N_5317,N_4909,N_4900);
nor U5318 (N_5318,N_5079,N_5074);
or U5319 (N_5319,N_4937,N_4849);
or U5320 (N_5320,N_4999,N_4930);
or U5321 (N_5321,N_4864,N_5056);
nor U5322 (N_5322,N_4826,N_4973);
nor U5323 (N_5323,N_5054,N_5086);
nor U5324 (N_5324,N_4953,N_4994);
or U5325 (N_5325,N_4887,N_4837);
nand U5326 (N_5326,N_5068,N_4811);
or U5327 (N_5327,N_5076,N_4978);
xor U5328 (N_5328,N_4868,N_4942);
or U5329 (N_5329,N_5043,N_4825);
nor U5330 (N_5330,N_4924,N_4952);
nor U5331 (N_5331,N_4829,N_5007);
and U5332 (N_5332,N_4828,N_5002);
nand U5333 (N_5333,N_4822,N_5093);
nand U5334 (N_5334,N_4903,N_5092);
xnor U5335 (N_5335,N_4970,N_4968);
and U5336 (N_5336,N_4853,N_5033);
nand U5337 (N_5337,N_4989,N_4861);
nor U5338 (N_5338,N_4916,N_4933);
xor U5339 (N_5339,N_4985,N_5020);
nor U5340 (N_5340,N_4916,N_5065);
nand U5341 (N_5341,N_4976,N_5079);
and U5342 (N_5342,N_4953,N_4896);
and U5343 (N_5343,N_4919,N_5076);
nor U5344 (N_5344,N_5011,N_4801);
nor U5345 (N_5345,N_4987,N_4908);
or U5346 (N_5346,N_5084,N_5078);
and U5347 (N_5347,N_4836,N_4889);
xnor U5348 (N_5348,N_4853,N_4964);
nand U5349 (N_5349,N_4880,N_4820);
nor U5350 (N_5350,N_4826,N_4837);
xor U5351 (N_5351,N_4817,N_4809);
and U5352 (N_5352,N_4965,N_5043);
and U5353 (N_5353,N_4997,N_4960);
and U5354 (N_5354,N_5000,N_4966);
nand U5355 (N_5355,N_5096,N_5020);
and U5356 (N_5356,N_5074,N_4872);
nor U5357 (N_5357,N_5003,N_4882);
or U5358 (N_5358,N_5075,N_4880);
or U5359 (N_5359,N_4965,N_5040);
xnor U5360 (N_5360,N_4936,N_5031);
and U5361 (N_5361,N_5009,N_4896);
nor U5362 (N_5362,N_4928,N_5097);
and U5363 (N_5363,N_5097,N_5088);
nor U5364 (N_5364,N_4977,N_4989);
xor U5365 (N_5365,N_4990,N_5008);
and U5366 (N_5366,N_4877,N_4922);
and U5367 (N_5367,N_4805,N_4841);
and U5368 (N_5368,N_4853,N_4820);
xor U5369 (N_5369,N_5013,N_4847);
xor U5370 (N_5370,N_5001,N_5010);
and U5371 (N_5371,N_5031,N_4904);
nand U5372 (N_5372,N_4818,N_4805);
and U5373 (N_5373,N_4850,N_5037);
nand U5374 (N_5374,N_5001,N_4859);
nand U5375 (N_5375,N_4846,N_4874);
nor U5376 (N_5376,N_4937,N_4865);
nor U5377 (N_5377,N_4919,N_4821);
nand U5378 (N_5378,N_4989,N_4826);
xnor U5379 (N_5379,N_5084,N_5029);
xnor U5380 (N_5380,N_4962,N_4920);
or U5381 (N_5381,N_4936,N_5054);
nand U5382 (N_5382,N_5026,N_5089);
and U5383 (N_5383,N_4986,N_5016);
xor U5384 (N_5384,N_4818,N_4800);
nand U5385 (N_5385,N_5073,N_4901);
xnor U5386 (N_5386,N_5066,N_4994);
xor U5387 (N_5387,N_5030,N_4874);
xnor U5388 (N_5388,N_4924,N_5083);
and U5389 (N_5389,N_4853,N_4916);
nand U5390 (N_5390,N_4996,N_4990);
and U5391 (N_5391,N_5064,N_4992);
xor U5392 (N_5392,N_5040,N_4936);
xor U5393 (N_5393,N_4940,N_5027);
nor U5394 (N_5394,N_5097,N_5087);
nand U5395 (N_5395,N_4873,N_4944);
and U5396 (N_5396,N_4927,N_5099);
or U5397 (N_5397,N_4858,N_5088);
or U5398 (N_5398,N_4828,N_4997);
nand U5399 (N_5399,N_5055,N_5071);
nand U5400 (N_5400,N_5177,N_5130);
and U5401 (N_5401,N_5333,N_5326);
nand U5402 (N_5402,N_5224,N_5207);
nand U5403 (N_5403,N_5141,N_5373);
nor U5404 (N_5404,N_5263,N_5379);
nand U5405 (N_5405,N_5228,N_5367);
or U5406 (N_5406,N_5168,N_5174);
nand U5407 (N_5407,N_5305,N_5233);
nor U5408 (N_5408,N_5231,N_5131);
xor U5409 (N_5409,N_5162,N_5129);
nand U5410 (N_5410,N_5176,N_5293);
nand U5411 (N_5411,N_5299,N_5111);
and U5412 (N_5412,N_5113,N_5268);
nand U5413 (N_5413,N_5192,N_5374);
xnor U5414 (N_5414,N_5262,N_5167);
and U5415 (N_5415,N_5296,N_5185);
and U5416 (N_5416,N_5390,N_5127);
or U5417 (N_5417,N_5285,N_5393);
and U5418 (N_5418,N_5140,N_5109);
xnor U5419 (N_5419,N_5363,N_5232);
or U5420 (N_5420,N_5237,N_5317);
nor U5421 (N_5421,N_5249,N_5352);
nor U5422 (N_5422,N_5202,N_5205);
and U5423 (N_5423,N_5230,N_5256);
or U5424 (N_5424,N_5220,N_5314);
and U5425 (N_5425,N_5124,N_5276);
or U5426 (N_5426,N_5375,N_5143);
nand U5427 (N_5427,N_5308,N_5284);
nand U5428 (N_5428,N_5105,N_5280);
nand U5429 (N_5429,N_5351,N_5337);
nand U5430 (N_5430,N_5304,N_5366);
nand U5431 (N_5431,N_5336,N_5264);
or U5432 (N_5432,N_5196,N_5195);
nand U5433 (N_5433,N_5139,N_5189);
nand U5434 (N_5434,N_5138,N_5252);
nand U5435 (N_5435,N_5211,N_5241);
nand U5436 (N_5436,N_5135,N_5161);
xnor U5437 (N_5437,N_5165,N_5267);
and U5438 (N_5438,N_5312,N_5272);
nand U5439 (N_5439,N_5319,N_5221);
nor U5440 (N_5440,N_5137,N_5219);
or U5441 (N_5441,N_5259,N_5112);
and U5442 (N_5442,N_5387,N_5398);
xor U5443 (N_5443,N_5370,N_5186);
nand U5444 (N_5444,N_5247,N_5157);
and U5445 (N_5445,N_5101,N_5238);
or U5446 (N_5446,N_5273,N_5171);
and U5447 (N_5447,N_5368,N_5327);
or U5448 (N_5448,N_5320,N_5147);
and U5449 (N_5449,N_5248,N_5321);
and U5450 (N_5450,N_5132,N_5110);
and U5451 (N_5451,N_5356,N_5206);
or U5452 (N_5452,N_5369,N_5297);
nand U5453 (N_5453,N_5155,N_5229);
or U5454 (N_5454,N_5134,N_5385);
nand U5455 (N_5455,N_5331,N_5234);
and U5456 (N_5456,N_5316,N_5244);
nor U5457 (N_5457,N_5274,N_5378);
xor U5458 (N_5458,N_5120,N_5322);
nor U5459 (N_5459,N_5144,N_5114);
nand U5460 (N_5460,N_5216,N_5246);
nor U5461 (N_5461,N_5125,N_5159);
and U5462 (N_5462,N_5344,N_5384);
nand U5463 (N_5463,N_5225,N_5235);
nor U5464 (N_5464,N_5173,N_5382);
or U5465 (N_5465,N_5332,N_5146);
or U5466 (N_5466,N_5371,N_5275);
xnor U5467 (N_5467,N_5180,N_5377);
nand U5468 (N_5468,N_5123,N_5266);
nor U5469 (N_5469,N_5106,N_5397);
and U5470 (N_5470,N_5239,N_5353);
and U5471 (N_5471,N_5270,N_5212);
xnor U5472 (N_5472,N_5283,N_5359);
and U5473 (N_5473,N_5289,N_5193);
xor U5474 (N_5474,N_5118,N_5278);
and U5475 (N_5475,N_5396,N_5295);
and U5476 (N_5476,N_5178,N_5100);
and U5477 (N_5477,N_5175,N_5136);
nor U5478 (N_5478,N_5222,N_5226);
nand U5479 (N_5479,N_5355,N_5343);
nor U5480 (N_5480,N_5291,N_5313);
xnor U5481 (N_5481,N_5342,N_5203);
xor U5482 (N_5482,N_5346,N_5362);
xnor U5483 (N_5483,N_5151,N_5279);
nor U5484 (N_5484,N_5345,N_5164);
and U5485 (N_5485,N_5376,N_5158);
nor U5486 (N_5486,N_5198,N_5341);
nor U5487 (N_5487,N_5133,N_5236);
xor U5488 (N_5488,N_5302,N_5349);
nor U5489 (N_5489,N_5301,N_5354);
and U5490 (N_5490,N_5142,N_5218);
nor U5491 (N_5491,N_5395,N_5357);
or U5492 (N_5492,N_5204,N_5380);
or U5493 (N_5493,N_5340,N_5102);
nor U5494 (N_5494,N_5152,N_5148);
and U5495 (N_5495,N_5288,N_5339);
and U5496 (N_5496,N_5290,N_5126);
nand U5497 (N_5497,N_5181,N_5242);
xnor U5498 (N_5498,N_5149,N_5169);
nor U5499 (N_5499,N_5104,N_5254);
or U5500 (N_5500,N_5217,N_5122);
or U5501 (N_5501,N_5315,N_5309);
nor U5502 (N_5502,N_5121,N_5303);
nand U5503 (N_5503,N_5245,N_5323);
and U5504 (N_5504,N_5328,N_5311);
nor U5505 (N_5505,N_5310,N_5389);
or U5506 (N_5506,N_5160,N_5128);
and U5507 (N_5507,N_5227,N_5282);
xnor U5508 (N_5508,N_5240,N_5117);
and U5509 (N_5509,N_5388,N_5338);
or U5510 (N_5510,N_5200,N_5277);
nand U5511 (N_5511,N_5243,N_5335);
and U5512 (N_5512,N_5119,N_5300);
nand U5513 (N_5513,N_5250,N_5394);
or U5514 (N_5514,N_5201,N_5358);
nor U5515 (N_5515,N_5265,N_5179);
nand U5516 (N_5516,N_5163,N_5150);
and U5517 (N_5517,N_5108,N_5360);
nor U5518 (N_5518,N_5381,N_5383);
nor U5519 (N_5519,N_5399,N_5208);
nand U5520 (N_5520,N_5223,N_5116);
nor U5521 (N_5521,N_5209,N_5298);
nor U5522 (N_5522,N_5318,N_5188);
nand U5523 (N_5523,N_5348,N_5292);
xor U5524 (N_5524,N_5251,N_5329);
nand U5525 (N_5525,N_5213,N_5391);
xnor U5526 (N_5526,N_5294,N_5306);
and U5527 (N_5527,N_5115,N_5287);
nor U5528 (N_5528,N_5334,N_5182);
and U5529 (N_5529,N_5214,N_5210);
and U5530 (N_5530,N_5255,N_5170);
and U5531 (N_5531,N_5361,N_5154);
or U5532 (N_5532,N_5330,N_5392);
nand U5533 (N_5533,N_5107,N_5166);
xnor U5534 (N_5534,N_5153,N_5145);
nor U5535 (N_5535,N_5324,N_5364);
and U5536 (N_5536,N_5156,N_5386);
nor U5537 (N_5537,N_5307,N_5372);
or U5538 (N_5538,N_5257,N_5187);
xor U5539 (N_5539,N_5271,N_5260);
and U5540 (N_5540,N_5281,N_5286);
and U5541 (N_5541,N_5347,N_5325);
nor U5542 (N_5542,N_5215,N_5197);
nand U5543 (N_5543,N_5199,N_5269);
xnor U5544 (N_5544,N_5103,N_5172);
or U5545 (N_5545,N_5183,N_5261);
xor U5546 (N_5546,N_5258,N_5190);
nor U5547 (N_5547,N_5194,N_5191);
xnor U5548 (N_5548,N_5253,N_5365);
xor U5549 (N_5549,N_5350,N_5184);
or U5550 (N_5550,N_5178,N_5238);
and U5551 (N_5551,N_5166,N_5202);
and U5552 (N_5552,N_5285,N_5203);
or U5553 (N_5553,N_5144,N_5354);
or U5554 (N_5554,N_5110,N_5272);
nor U5555 (N_5555,N_5320,N_5366);
and U5556 (N_5556,N_5194,N_5290);
nor U5557 (N_5557,N_5315,N_5126);
or U5558 (N_5558,N_5330,N_5360);
xnor U5559 (N_5559,N_5286,N_5381);
or U5560 (N_5560,N_5231,N_5172);
xor U5561 (N_5561,N_5372,N_5212);
xnor U5562 (N_5562,N_5183,N_5168);
nor U5563 (N_5563,N_5181,N_5172);
nor U5564 (N_5564,N_5237,N_5127);
xor U5565 (N_5565,N_5333,N_5189);
or U5566 (N_5566,N_5296,N_5223);
nor U5567 (N_5567,N_5187,N_5138);
and U5568 (N_5568,N_5158,N_5304);
nor U5569 (N_5569,N_5242,N_5261);
or U5570 (N_5570,N_5282,N_5390);
or U5571 (N_5571,N_5170,N_5310);
nor U5572 (N_5572,N_5105,N_5227);
xnor U5573 (N_5573,N_5191,N_5391);
xor U5574 (N_5574,N_5382,N_5153);
xnor U5575 (N_5575,N_5185,N_5254);
or U5576 (N_5576,N_5318,N_5194);
nor U5577 (N_5577,N_5140,N_5398);
or U5578 (N_5578,N_5218,N_5221);
nand U5579 (N_5579,N_5146,N_5333);
nor U5580 (N_5580,N_5279,N_5177);
or U5581 (N_5581,N_5356,N_5173);
xnor U5582 (N_5582,N_5266,N_5393);
xnor U5583 (N_5583,N_5162,N_5248);
xor U5584 (N_5584,N_5180,N_5200);
nor U5585 (N_5585,N_5179,N_5241);
nand U5586 (N_5586,N_5261,N_5266);
nand U5587 (N_5587,N_5111,N_5387);
xor U5588 (N_5588,N_5313,N_5272);
or U5589 (N_5589,N_5351,N_5116);
xnor U5590 (N_5590,N_5368,N_5277);
or U5591 (N_5591,N_5299,N_5150);
xor U5592 (N_5592,N_5253,N_5105);
nor U5593 (N_5593,N_5124,N_5398);
or U5594 (N_5594,N_5271,N_5365);
and U5595 (N_5595,N_5391,N_5393);
nor U5596 (N_5596,N_5273,N_5202);
nor U5597 (N_5597,N_5244,N_5371);
and U5598 (N_5598,N_5102,N_5202);
or U5599 (N_5599,N_5363,N_5239);
nand U5600 (N_5600,N_5197,N_5222);
nand U5601 (N_5601,N_5125,N_5294);
xor U5602 (N_5602,N_5355,N_5148);
nor U5603 (N_5603,N_5396,N_5289);
nand U5604 (N_5604,N_5102,N_5171);
nor U5605 (N_5605,N_5244,N_5164);
or U5606 (N_5606,N_5154,N_5282);
nand U5607 (N_5607,N_5276,N_5229);
nor U5608 (N_5608,N_5350,N_5187);
and U5609 (N_5609,N_5148,N_5168);
nand U5610 (N_5610,N_5380,N_5215);
and U5611 (N_5611,N_5349,N_5315);
xor U5612 (N_5612,N_5274,N_5143);
and U5613 (N_5613,N_5156,N_5384);
nand U5614 (N_5614,N_5199,N_5398);
nor U5615 (N_5615,N_5293,N_5195);
nor U5616 (N_5616,N_5110,N_5291);
nor U5617 (N_5617,N_5150,N_5302);
xnor U5618 (N_5618,N_5227,N_5141);
xnor U5619 (N_5619,N_5169,N_5255);
xor U5620 (N_5620,N_5341,N_5161);
or U5621 (N_5621,N_5373,N_5168);
nand U5622 (N_5622,N_5392,N_5324);
or U5623 (N_5623,N_5139,N_5169);
nor U5624 (N_5624,N_5261,N_5211);
xor U5625 (N_5625,N_5158,N_5146);
nand U5626 (N_5626,N_5310,N_5323);
and U5627 (N_5627,N_5383,N_5145);
or U5628 (N_5628,N_5274,N_5167);
and U5629 (N_5629,N_5333,N_5291);
or U5630 (N_5630,N_5124,N_5378);
and U5631 (N_5631,N_5260,N_5320);
or U5632 (N_5632,N_5364,N_5227);
or U5633 (N_5633,N_5332,N_5379);
and U5634 (N_5634,N_5208,N_5385);
nand U5635 (N_5635,N_5304,N_5278);
nor U5636 (N_5636,N_5198,N_5260);
nor U5637 (N_5637,N_5359,N_5318);
nor U5638 (N_5638,N_5135,N_5164);
and U5639 (N_5639,N_5342,N_5244);
and U5640 (N_5640,N_5126,N_5301);
nand U5641 (N_5641,N_5283,N_5313);
and U5642 (N_5642,N_5325,N_5219);
and U5643 (N_5643,N_5333,N_5306);
nor U5644 (N_5644,N_5152,N_5222);
nor U5645 (N_5645,N_5263,N_5105);
nor U5646 (N_5646,N_5342,N_5109);
and U5647 (N_5647,N_5176,N_5342);
or U5648 (N_5648,N_5394,N_5240);
and U5649 (N_5649,N_5399,N_5170);
nand U5650 (N_5650,N_5175,N_5326);
or U5651 (N_5651,N_5221,N_5173);
xnor U5652 (N_5652,N_5107,N_5267);
and U5653 (N_5653,N_5283,N_5395);
nand U5654 (N_5654,N_5208,N_5352);
nor U5655 (N_5655,N_5180,N_5143);
nor U5656 (N_5656,N_5280,N_5193);
and U5657 (N_5657,N_5139,N_5339);
nor U5658 (N_5658,N_5190,N_5153);
or U5659 (N_5659,N_5181,N_5301);
xnor U5660 (N_5660,N_5163,N_5126);
nor U5661 (N_5661,N_5115,N_5196);
nor U5662 (N_5662,N_5351,N_5300);
or U5663 (N_5663,N_5233,N_5296);
xor U5664 (N_5664,N_5157,N_5228);
nand U5665 (N_5665,N_5189,N_5295);
nand U5666 (N_5666,N_5131,N_5246);
nor U5667 (N_5667,N_5186,N_5373);
and U5668 (N_5668,N_5373,N_5275);
xnor U5669 (N_5669,N_5166,N_5362);
nand U5670 (N_5670,N_5115,N_5250);
nand U5671 (N_5671,N_5340,N_5361);
nor U5672 (N_5672,N_5392,N_5318);
nor U5673 (N_5673,N_5102,N_5176);
nor U5674 (N_5674,N_5352,N_5200);
nor U5675 (N_5675,N_5340,N_5308);
nand U5676 (N_5676,N_5329,N_5131);
or U5677 (N_5677,N_5306,N_5156);
nor U5678 (N_5678,N_5344,N_5205);
xor U5679 (N_5679,N_5319,N_5336);
nor U5680 (N_5680,N_5237,N_5259);
or U5681 (N_5681,N_5325,N_5333);
nor U5682 (N_5682,N_5251,N_5123);
nand U5683 (N_5683,N_5175,N_5161);
and U5684 (N_5684,N_5222,N_5288);
nand U5685 (N_5685,N_5289,N_5121);
nand U5686 (N_5686,N_5162,N_5192);
nand U5687 (N_5687,N_5374,N_5238);
xnor U5688 (N_5688,N_5346,N_5233);
nand U5689 (N_5689,N_5162,N_5376);
xnor U5690 (N_5690,N_5213,N_5125);
or U5691 (N_5691,N_5300,N_5366);
xor U5692 (N_5692,N_5159,N_5175);
xnor U5693 (N_5693,N_5209,N_5391);
xor U5694 (N_5694,N_5318,N_5267);
and U5695 (N_5695,N_5131,N_5160);
xnor U5696 (N_5696,N_5139,N_5119);
and U5697 (N_5697,N_5303,N_5126);
or U5698 (N_5698,N_5219,N_5250);
and U5699 (N_5699,N_5265,N_5177);
xor U5700 (N_5700,N_5673,N_5597);
nand U5701 (N_5701,N_5650,N_5476);
and U5702 (N_5702,N_5502,N_5660);
and U5703 (N_5703,N_5684,N_5469);
or U5704 (N_5704,N_5631,N_5470);
and U5705 (N_5705,N_5690,N_5570);
nor U5706 (N_5706,N_5537,N_5675);
nor U5707 (N_5707,N_5698,N_5444);
nor U5708 (N_5708,N_5509,N_5401);
nor U5709 (N_5709,N_5475,N_5495);
xnor U5710 (N_5710,N_5462,N_5605);
or U5711 (N_5711,N_5487,N_5588);
or U5712 (N_5712,N_5686,N_5543);
or U5713 (N_5713,N_5593,N_5474);
or U5714 (N_5714,N_5621,N_5435);
or U5715 (N_5715,N_5546,N_5434);
and U5716 (N_5716,N_5425,N_5654);
xnor U5717 (N_5717,N_5594,N_5516);
xnor U5718 (N_5718,N_5436,N_5582);
nand U5719 (N_5719,N_5524,N_5608);
and U5720 (N_5720,N_5672,N_5480);
nor U5721 (N_5721,N_5424,N_5533);
nand U5722 (N_5722,N_5527,N_5633);
and U5723 (N_5723,N_5587,N_5497);
nand U5724 (N_5724,N_5630,N_5699);
and U5725 (N_5725,N_5664,N_5590);
nand U5726 (N_5726,N_5421,N_5467);
or U5727 (N_5727,N_5648,N_5433);
or U5728 (N_5728,N_5490,N_5586);
xnor U5729 (N_5729,N_5507,N_5519);
nor U5730 (N_5730,N_5472,N_5418);
nor U5731 (N_5731,N_5610,N_5641);
nor U5732 (N_5732,N_5625,N_5419);
or U5733 (N_5733,N_5529,N_5693);
nand U5734 (N_5734,N_5437,N_5429);
and U5735 (N_5735,N_5554,N_5563);
xor U5736 (N_5736,N_5620,N_5541);
or U5737 (N_5737,N_5657,N_5409);
or U5738 (N_5738,N_5580,N_5477);
nor U5739 (N_5739,N_5432,N_5493);
xnor U5740 (N_5740,N_5518,N_5456);
xor U5741 (N_5741,N_5674,N_5651);
or U5742 (N_5742,N_5676,N_5611);
and U5743 (N_5743,N_5565,N_5410);
or U5744 (N_5744,N_5540,N_5679);
xor U5745 (N_5745,N_5647,N_5431);
nor U5746 (N_5746,N_5569,N_5691);
and U5747 (N_5747,N_5468,N_5417);
or U5748 (N_5748,N_5656,N_5501);
and U5749 (N_5749,N_5685,N_5411);
and U5750 (N_5750,N_5413,N_5426);
and U5751 (N_5751,N_5515,N_5451);
nand U5752 (N_5752,N_5430,N_5688);
xnor U5753 (N_5753,N_5552,N_5615);
xnor U5754 (N_5754,N_5579,N_5535);
or U5755 (N_5755,N_5655,N_5407);
nor U5756 (N_5756,N_5643,N_5466);
nor U5757 (N_5757,N_5689,N_5481);
xnor U5758 (N_5758,N_5640,N_5616);
nor U5759 (N_5759,N_5498,N_5403);
and U5760 (N_5760,N_5405,N_5559);
and U5761 (N_5761,N_5613,N_5578);
xor U5762 (N_5762,N_5601,N_5662);
and U5763 (N_5763,N_5568,N_5575);
and U5764 (N_5764,N_5439,N_5683);
nor U5765 (N_5765,N_5634,N_5652);
or U5766 (N_5766,N_5596,N_5528);
nand U5767 (N_5767,N_5557,N_5551);
nand U5768 (N_5768,N_5423,N_5471);
xor U5769 (N_5769,N_5682,N_5549);
nand U5770 (N_5770,N_5681,N_5504);
or U5771 (N_5771,N_5520,N_5473);
xor U5772 (N_5772,N_5523,N_5526);
or U5773 (N_5773,N_5503,N_5677);
and U5774 (N_5774,N_5428,N_5452);
or U5775 (N_5775,N_5584,N_5442);
xor U5776 (N_5776,N_5463,N_5482);
nand U5777 (N_5777,N_5623,N_5458);
nor U5778 (N_5778,N_5694,N_5408);
or U5779 (N_5779,N_5619,N_5485);
nor U5780 (N_5780,N_5602,N_5511);
xor U5781 (N_5781,N_5658,N_5595);
or U5782 (N_5782,N_5618,N_5448);
and U5783 (N_5783,N_5598,N_5667);
nor U5784 (N_5784,N_5457,N_5538);
and U5785 (N_5785,N_5505,N_5659);
xnor U5786 (N_5786,N_5514,N_5669);
xnor U5787 (N_5787,N_5612,N_5464);
nand U5788 (N_5788,N_5697,N_5488);
nor U5789 (N_5789,N_5609,N_5500);
xnor U5790 (N_5790,N_5402,N_5695);
xnor U5791 (N_5791,N_5492,N_5406);
nand U5792 (N_5792,N_5599,N_5440);
nand U5793 (N_5793,N_5517,N_5522);
or U5794 (N_5794,N_5531,N_5627);
or U5795 (N_5795,N_5574,N_5553);
or U5796 (N_5796,N_5521,N_5532);
nor U5797 (N_5797,N_5663,N_5499);
and U5798 (N_5798,N_5628,N_5585);
or U5799 (N_5799,N_5646,N_5513);
nand U5800 (N_5800,N_5454,N_5583);
or U5801 (N_5801,N_5642,N_5668);
nor U5802 (N_5802,N_5560,N_5606);
nor U5803 (N_5803,N_5441,N_5486);
xor U5804 (N_5804,N_5412,N_5455);
xor U5805 (N_5805,N_5550,N_5591);
or U5806 (N_5806,N_5489,N_5508);
or U5807 (N_5807,N_5576,N_5561);
nand U5808 (N_5808,N_5645,N_5446);
and U5809 (N_5809,N_5624,N_5422);
nand U5810 (N_5810,N_5453,N_5414);
or U5811 (N_5811,N_5506,N_5692);
nor U5812 (N_5812,N_5427,N_5678);
or U5813 (N_5813,N_5661,N_5644);
or U5814 (N_5814,N_5534,N_5562);
and U5815 (N_5815,N_5617,N_5567);
and U5816 (N_5816,N_5639,N_5600);
nand U5817 (N_5817,N_5450,N_5512);
nand U5818 (N_5818,N_5449,N_5438);
nor U5819 (N_5819,N_5629,N_5547);
nand U5820 (N_5820,N_5573,N_5510);
or U5821 (N_5821,N_5404,N_5530);
nand U5822 (N_5822,N_5459,N_5556);
nand U5823 (N_5823,N_5670,N_5483);
nand U5824 (N_5824,N_5665,N_5555);
and U5825 (N_5825,N_5496,N_5622);
xor U5826 (N_5826,N_5636,N_5589);
nand U5827 (N_5827,N_5525,N_5671);
nor U5828 (N_5828,N_5687,N_5416);
and U5829 (N_5829,N_5544,N_5545);
nor U5830 (N_5830,N_5581,N_5494);
nor U5831 (N_5831,N_5491,N_5680);
nand U5832 (N_5832,N_5536,N_5447);
nor U5833 (N_5833,N_5571,N_5566);
nand U5834 (N_5834,N_5484,N_5653);
xor U5835 (N_5835,N_5415,N_5420);
nand U5836 (N_5836,N_5626,N_5548);
or U5837 (N_5837,N_5539,N_5572);
or U5838 (N_5838,N_5696,N_5465);
or U5839 (N_5839,N_5445,N_5479);
nor U5840 (N_5840,N_5632,N_5592);
nand U5841 (N_5841,N_5542,N_5638);
nor U5842 (N_5842,N_5649,N_5558);
nor U5843 (N_5843,N_5400,N_5577);
and U5844 (N_5844,N_5443,N_5603);
xnor U5845 (N_5845,N_5666,N_5635);
xnor U5846 (N_5846,N_5637,N_5478);
nand U5847 (N_5847,N_5607,N_5461);
or U5848 (N_5848,N_5604,N_5460);
and U5849 (N_5849,N_5614,N_5564);
xor U5850 (N_5850,N_5560,N_5494);
nor U5851 (N_5851,N_5575,N_5606);
xnor U5852 (N_5852,N_5669,N_5591);
nor U5853 (N_5853,N_5568,N_5591);
nand U5854 (N_5854,N_5472,N_5680);
nand U5855 (N_5855,N_5524,N_5590);
xor U5856 (N_5856,N_5672,N_5650);
or U5857 (N_5857,N_5513,N_5699);
nand U5858 (N_5858,N_5659,N_5478);
nor U5859 (N_5859,N_5422,N_5634);
xnor U5860 (N_5860,N_5562,N_5663);
nor U5861 (N_5861,N_5637,N_5599);
nor U5862 (N_5862,N_5575,N_5623);
nor U5863 (N_5863,N_5652,N_5635);
xnor U5864 (N_5864,N_5475,N_5409);
or U5865 (N_5865,N_5407,N_5411);
and U5866 (N_5866,N_5536,N_5401);
nand U5867 (N_5867,N_5480,N_5555);
or U5868 (N_5868,N_5662,N_5632);
xnor U5869 (N_5869,N_5533,N_5502);
and U5870 (N_5870,N_5413,N_5542);
and U5871 (N_5871,N_5448,N_5425);
nand U5872 (N_5872,N_5689,N_5457);
nor U5873 (N_5873,N_5617,N_5671);
nor U5874 (N_5874,N_5639,N_5566);
or U5875 (N_5875,N_5418,N_5550);
nand U5876 (N_5876,N_5529,N_5490);
and U5877 (N_5877,N_5548,N_5577);
nor U5878 (N_5878,N_5654,N_5570);
xnor U5879 (N_5879,N_5457,N_5401);
xnor U5880 (N_5880,N_5692,N_5411);
nor U5881 (N_5881,N_5457,N_5634);
and U5882 (N_5882,N_5403,N_5555);
and U5883 (N_5883,N_5494,N_5507);
and U5884 (N_5884,N_5580,N_5566);
and U5885 (N_5885,N_5485,N_5649);
nand U5886 (N_5886,N_5454,N_5530);
nand U5887 (N_5887,N_5697,N_5551);
nor U5888 (N_5888,N_5425,N_5612);
xor U5889 (N_5889,N_5621,N_5477);
nor U5890 (N_5890,N_5587,N_5646);
xnor U5891 (N_5891,N_5619,N_5428);
xnor U5892 (N_5892,N_5493,N_5471);
xor U5893 (N_5893,N_5612,N_5677);
nand U5894 (N_5894,N_5632,N_5415);
nor U5895 (N_5895,N_5650,N_5610);
xor U5896 (N_5896,N_5673,N_5493);
nand U5897 (N_5897,N_5576,N_5632);
nand U5898 (N_5898,N_5455,N_5597);
xnor U5899 (N_5899,N_5644,N_5498);
and U5900 (N_5900,N_5458,N_5430);
nand U5901 (N_5901,N_5635,N_5535);
nand U5902 (N_5902,N_5563,N_5459);
nand U5903 (N_5903,N_5520,N_5531);
nand U5904 (N_5904,N_5464,N_5592);
or U5905 (N_5905,N_5429,N_5502);
or U5906 (N_5906,N_5585,N_5414);
nor U5907 (N_5907,N_5624,N_5661);
nand U5908 (N_5908,N_5485,N_5666);
nor U5909 (N_5909,N_5676,N_5478);
and U5910 (N_5910,N_5506,N_5693);
or U5911 (N_5911,N_5547,N_5580);
or U5912 (N_5912,N_5590,N_5412);
or U5913 (N_5913,N_5437,N_5424);
xor U5914 (N_5914,N_5625,N_5514);
xor U5915 (N_5915,N_5514,N_5433);
and U5916 (N_5916,N_5628,N_5668);
and U5917 (N_5917,N_5638,N_5614);
or U5918 (N_5918,N_5473,N_5554);
nor U5919 (N_5919,N_5530,N_5450);
nand U5920 (N_5920,N_5569,N_5520);
xor U5921 (N_5921,N_5616,N_5696);
nor U5922 (N_5922,N_5589,N_5657);
nor U5923 (N_5923,N_5678,N_5504);
xnor U5924 (N_5924,N_5507,N_5464);
or U5925 (N_5925,N_5445,N_5414);
xnor U5926 (N_5926,N_5539,N_5662);
and U5927 (N_5927,N_5669,N_5496);
xnor U5928 (N_5928,N_5454,N_5423);
and U5929 (N_5929,N_5519,N_5603);
nand U5930 (N_5930,N_5534,N_5672);
nor U5931 (N_5931,N_5615,N_5601);
xnor U5932 (N_5932,N_5624,N_5553);
and U5933 (N_5933,N_5400,N_5442);
or U5934 (N_5934,N_5556,N_5603);
nand U5935 (N_5935,N_5581,N_5627);
and U5936 (N_5936,N_5652,N_5646);
nor U5937 (N_5937,N_5429,N_5525);
xor U5938 (N_5938,N_5417,N_5425);
xnor U5939 (N_5939,N_5450,N_5585);
xor U5940 (N_5940,N_5431,N_5651);
xor U5941 (N_5941,N_5434,N_5627);
and U5942 (N_5942,N_5684,N_5581);
nor U5943 (N_5943,N_5568,N_5516);
xnor U5944 (N_5944,N_5498,N_5523);
xor U5945 (N_5945,N_5564,N_5517);
and U5946 (N_5946,N_5557,N_5472);
nand U5947 (N_5947,N_5501,N_5697);
and U5948 (N_5948,N_5437,N_5413);
nand U5949 (N_5949,N_5414,N_5462);
xnor U5950 (N_5950,N_5579,N_5676);
xor U5951 (N_5951,N_5514,N_5401);
xor U5952 (N_5952,N_5664,N_5649);
and U5953 (N_5953,N_5449,N_5531);
xor U5954 (N_5954,N_5476,N_5522);
xnor U5955 (N_5955,N_5629,N_5428);
nand U5956 (N_5956,N_5689,N_5600);
or U5957 (N_5957,N_5584,N_5488);
xor U5958 (N_5958,N_5590,N_5596);
xnor U5959 (N_5959,N_5431,N_5588);
nand U5960 (N_5960,N_5537,N_5445);
nor U5961 (N_5961,N_5682,N_5678);
or U5962 (N_5962,N_5519,N_5671);
or U5963 (N_5963,N_5443,N_5525);
nor U5964 (N_5964,N_5595,N_5402);
nor U5965 (N_5965,N_5468,N_5693);
nor U5966 (N_5966,N_5471,N_5694);
nor U5967 (N_5967,N_5486,N_5468);
nor U5968 (N_5968,N_5491,N_5504);
nor U5969 (N_5969,N_5422,N_5447);
xor U5970 (N_5970,N_5677,N_5618);
and U5971 (N_5971,N_5645,N_5686);
nand U5972 (N_5972,N_5600,N_5592);
xnor U5973 (N_5973,N_5427,N_5411);
nor U5974 (N_5974,N_5465,N_5656);
xnor U5975 (N_5975,N_5519,N_5567);
xor U5976 (N_5976,N_5539,N_5689);
or U5977 (N_5977,N_5582,N_5600);
nor U5978 (N_5978,N_5494,N_5439);
nor U5979 (N_5979,N_5444,N_5635);
and U5980 (N_5980,N_5460,N_5668);
or U5981 (N_5981,N_5412,N_5679);
or U5982 (N_5982,N_5442,N_5594);
nor U5983 (N_5983,N_5626,N_5611);
and U5984 (N_5984,N_5549,N_5587);
nand U5985 (N_5985,N_5694,N_5487);
or U5986 (N_5986,N_5563,N_5643);
and U5987 (N_5987,N_5435,N_5641);
or U5988 (N_5988,N_5544,N_5595);
xnor U5989 (N_5989,N_5648,N_5678);
nand U5990 (N_5990,N_5542,N_5421);
xnor U5991 (N_5991,N_5479,N_5553);
and U5992 (N_5992,N_5679,N_5665);
and U5993 (N_5993,N_5543,N_5665);
xnor U5994 (N_5994,N_5695,N_5459);
and U5995 (N_5995,N_5400,N_5449);
or U5996 (N_5996,N_5689,N_5534);
and U5997 (N_5997,N_5542,N_5538);
nor U5998 (N_5998,N_5432,N_5610);
nand U5999 (N_5999,N_5420,N_5557);
or U6000 (N_6000,N_5924,N_5943);
and U6001 (N_6001,N_5766,N_5751);
and U6002 (N_6002,N_5722,N_5901);
nand U6003 (N_6003,N_5890,N_5716);
nor U6004 (N_6004,N_5739,N_5831);
or U6005 (N_6005,N_5755,N_5863);
xnor U6006 (N_6006,N_5908,N_5797);
or U6007 (N_6007,N_5931,N_5784);
and U6008 (N_6008,N_5788,N_5760);
or U6009 (N_6009,N_5852,N_5795);
nor U6010 (N_6010,N_5824,N_5830);
nand U6011 (N_6011,N_5894,N_5954);
xor U6012 (N_6012,N_5922,N_5854);
and U6013 (N_6013,N_5891,N_5871);
nor U6014 (N_6014,N_5750,N_5771);
xnor U6015 (N_6015,N_5999,N_5861);
or U6016 (N_6016,N_5879,N_5906);
and U6017 (N_6017,N_5970,N_5735);
and U6018 (N_6018,N_5897,N_5713);
or U6019 (N_6019,N_5940,N_5947);
nor U6020 (N_6020,N_5944,N_5780);
xor U6021 (N_6021,N_5717,N_5859);
xor U6022 (N_6022,N_5878,N_5742);
nor U6023 (N_6023,N_5885,N_5787);
nor U6024 (N_6024,N_5992,N_5703);
nor U6025 (N_6025,N_5734,N_5721);
xnor U6026 (N_6026,N_5952,N_5864);
xnor U6027 (N_6027,N_5958,N_5994);
or U6028 (N_6028,N_5802,N_5911);
and U6029 (N_6029,N_5786,N_5855);
xnor U6030 (N_6030,N_5728,N_5828);
nand U6031 (N_6031,N_5840,N_5715);
xnor U6032 (N_6032,N_5711,N_5837);
or U6033 (N_6033,N_5835,N_5892);
xnor U6034 (N_6034,N_5929,N_5932);
and U6035 (N_6035,N_5991,N_5986);
nor U6036 (N_6036,N_5977,N_5939);
or U6037 (N_6037,N_5978,N_5895);
or U6038 (N_6038,N_5925,N_5997);
nor U6039 (N_6039,N_5832,N_5720);
or U6040 (N_6040,N_5725,N_5950);
nand U6041 (N_6041,N_5983,N_5822);
and U6042 (N_6042,N_5921,N_5814);
or U6043 (N_6043,N_5708,N_5752);
and U6044 (N_6044,N_5769,N_5846);
nor U6045 (N_6045,N_5733,N_5710);
or U6046 (N_6046,N_5873,N_5872);
xor U6047 (N_6047,N_5881,N_5746);
or U6048 (N_6048,N_5763,N_5800);
nor U6049 (N_6049,N_5756,N_5839);
nor U6050 (N_6050,N_5900,N_5823);
nor U6051 (N_6051,N_5903,N_5914);
nor U6052 (N_6052,N_5731,N_5794);
nor U6053 (N_6053,N_5841,N_5730);
or U6054 (N_6054,N_5803,N_5963);
nor U6055 (N_6055,N_5806,N_5880);
nor U6056 (N_6056,N_5777,N_5928);
or U6057 (N_6057,N_5812,N_5704);
xnor U6058 (N_6058,N_5969,N_5792);
and U6059 (N_6059,N_5945,N_5876);
or U6060 (N_6060,N_5745,N_5799);
and U6061 (N_6061,N_5882,N_5816);
nor U6062 (N_6062,N_5920,N_5813);
nor U6063 (N_6063,N_5818,N_5853);
nor U6064 (N_6064,N_5966,N_5836);
nor U6065 (N_6065,N_5990,N_5738);
and U6066 (N_6066,N_5982,N_5727);
nor U6067 (N_6067,N_5916,N_5865);
or U6068 (N_6068,N_5793,N_5754);
and U6069 (N_6069,N_5807,N_5987);
or U6070 (N_6070,N_5709,N_5706);
xor U6071 (N_6071,N_5961,N_5765);
nand U6072 (N_6072,N_5953,N_5757);
xnor U6073 (N_6073,N_5967,N_5849);
xnor U6074 (N_6074,N_5741,N_5843);
nand U6075 (N_6075,N_5789,N_5949);
or U6076 (N_6076,N_5926,N_5888);
xor U6077 (N_6077,N_5848,N_5874);
and U6078 (N_6078,N_5886,N_5956);
nor U6079 (N_6079,N_5779,N_5829);
nor U6080 (N_6080,N_5842,N_5775);
nand U6081 (N_6081,N_5898,N_5860);
nor U6082 (N_6082,N_5905,N_5783);
or U6083 (N_6083,N_5942,N_5762);
or U6084 (N_6084,N_5917,N_5737);
and U6085 (N_6085,N_5913,N_5866);
nor U6086 (N_6086,N_5838,N_5781);
nand U6087 (N_6087,N_5770,N_5985);
xnor U6088 (N_6088,N_5971,N_5896);
or U6089 (N_6089,N_5912,N_5851);
nand U6090 (N_6090,N_5764,N_5868);
xnor U6091 (N_6091,N_5700,N_5753);
nor U6092 (N_6092,N_5815,N_5858);
and U6093 (N_6093,N_5941,N_5948);
or U6094 (N_6094,N_5826,N_5981);
nor U6095 (N_6095,N_5960,N_5732);
nor U6096 (N_6096,N_5810,N_5712);
xnor U6097 (N_6097,N_5736,N_5778);
nand U6098 (N_6098,N_5936,N_5959);
or U6099 (N_6099,N_5877,N_5974);
nor U6100 (N_6100,N_5834,N_5951);
and U6101 (N_6101,N_5904,N_5776);
xor U6102 (N_6102,N_5809,N_5980);
xnor U6103 (N_6103,N_5790,N_5935);
nor U6104 (N_6104,N_5869,N_5930);
and U6105 (N_6105,N_5782,N_5759);
and U6106 (N_6106,N_5850,N_5938);
or U6107 (N_6107,N_5862,N_5923);
xnor U6108 (N_6108,N_5743,N_5804);
and U6109 (N_6109,N_5899,N_5937);
or U6110 (N_6110,N_5976,N_5856);
or U6111 (N_6111,N_5744,N_5748);
or U6112 (N_6112,N_5749,N_5984);
and U6113 (N_6113,N_5933,N_5965);
or U6114 (N_6114,N_5719,N_5772);
and U6115 (N_6115,N_5988,N_5867);
xor U6116 (N_6116,N_5893,N_5827);
and U6117 (N_6117,N_5902,N_5909);
and U6118 (N_6118,N_5791,N_5844);
nand U6119 (N_6119,N_5998,N_5968);
xor U6120 (N_6120,N_5767,N_5973);
and U6121 (N_6121,N_5889,N_5714);
or U6122 (N_6122,N_5724,N_5975);
and U6123 (N_6123,N_5758,N_5884);
nor U6124 (N_6124,N_5915,N_5723);
nand U6125 (N_6125,N_5740,N_5768);
and U6126 (N_6126,N_5955,N_5996);
nor U6127 (N_6127,N_5907,N_5707);
nand U6128 (N_6128,N_5887,N_5819);
nand U6129 (N_6129,N_5847,N_5773);
xor U6130 (N_6130,N_5833,N_5701);
and U6131 (N_6131,N_5726,N_5875);
nor U6132 (N_6132,N_5870,N_5817);
or U6133 (N_6133,N_5995,N_5808);
nor U6134 (N_6134,N_5919,N_5979);
xnor U6135 (N_6135,N_5857,N_5934);
nor U6136 (N_6136,N_5927,N_5962);
nand U6137 (N_6137,N_5993,N_5946);
or U6138 (N_6138,N_5957,N_5796);
nor U6139 (N_6139,N_5798,N_5747);
and U6140 (N_6140,N_5825,N_5811);
nand U6141 (N_6141,N_5705,N_5964);
and U6142 (N_6142,N_5910,N_5729);
nor U6143 (N_6143,N_5805,N_5821);
or U6144 (N_6144,N_5883,N_5801);
and U6145 (N_6145,N_5785,N_5774);
nor U6146 (N_6146,N_5702,N_5845);
nor U6147 (N_6147,N_5918,N_5972);
and U6148 (N_6148,N_5989,N_5718);
and U6149 (N_6149,N_5820,N_5761);
nor U6150 (N_6150,N_5713,N_5916);
nor U6151 (N_6151,N_5769,N_5887);
xnor U6152 (N_6152,N_5969,N_5828);
or U6153 (N_6153,N_5857,N_5709);
nand U6154 (N_6154,N_5722,N_5721);
xor U6155 (N_6155,N_5989,N_5991);
xnor U6156 (N_6156,N_5762,N_5748);
nand U6157 (N_6157,N_5838,N_5731);
and U6158 (N_6158,N_5989,N_5776);
and U6159 (N_6159,N_5746,N_5831);
and U6160 (N_6160,N_5808,N_5926);
xnor U6161 (N_6161,N_5875,N_5966);
nor U6162 (N_6162,N_5912,N_5911);
and U6163 (N_6163,N_5941,N_5860);
xor U6164 (N_6164,N_5888,N_5752);
xor U6165 (N_6165,N_5973,N_5985);
and U6166 (N_6166,N_5933,N_5993);
and U6167 (N_6167,N_5864,N_5725);
and U6168 (N_6168,N_5728,N_5802);
nand U6169 (N_6169,N_5907,N_5909);
xnor U6170 (N_6170,N_5832,N_5721);
nor U6171 (N_6171,N_5721,N_5896);
or U6172 (N_6172,N_5848,N_5753);
xor U6173 (N_6173,N_5884,N_5738);
or U6174 (N_6174,N_5857,N_5953);
nor U6175 (N_6175,N_5946,N_5730);
xor U6176 (N_6176,N_5871,N_5832);
and U6177 (N_6177,N_5866,N_5975);
or U6178 (N_6178,N_5789,N_5925);
nand U6179 (N_6179,N_5839,N_5971);
or U6180 (N_6180,N_5700,N_5968);
xor U6181 (N_6181,N_5928,N_5751);
and U6182 (N_6182,N_5911,N_5948);
xnor U6183 (N_6183,N_5932,N_5898);
and U6184 (N_6184,N_5702,N_5948);
nor U6185 (N_6185,N_5934,N_5769);
and U6186 (N_6186,N_5880,N_5918);
and U6187 (N_6187,N_5731,N_5773);
nand U6188 (N_6188,N_5744,N_5941);
nand U6189 (N_6189,N_5769,N_5778);
xnor U6190 (N_6190,N_5987,N_5936);
nand U6191 (N_6191,N_5967,N_5826);
nand U6192 (N_6192,N_5746,N_5855);
and U6193 (N_6193,N_5903,N_5726);
nand U6194 (N_6194,N_5848,N_5975);
or U6195 (N_6195,N_5750,N_5751);
nor U6196 (N_6196,N_5857,N_5899);
and U6197 (N_6197,N_5763,N_5831);
nor U6198 (N_6198,N_5755,N_5985);
nor U6199 (N_6199,N_5972,N_5767);
nand U6200 (N_6200,N_5915,N_5886);
or U6201 (N_6201,N_5909,N_5823);
xnor U6202 (N_6202,N_5852,N_5799);
nor U6203 (N_6203,N_5895,N_5746);
and U6204 (N_6204,N_5910,N_5883);
nand U6205 (N_6205,N_5864,N_5796);
xnor U6206 (N_6206,N_5752,N_5795);
xor U6207 (N_6207,N_5951,N_5807);
xor U6208 (N_6208,N_5777,N_5999);
and U6209 (N_6209,N_5803,N_5709);
and U6210 (N_6210,N_5997,N_5905);
xnor U6211 (N_6211,N_5977,N_5864);
nor U6212 (N_6212,N_5972,N_5992);
or U6213 (N_6213,N_5930,N_5852);
nand U6214 (N_6214,N_5862,N_5982);
and U6215 (N_6215,N_5705,N_5801);
or U6216 (N_6216,N_5754,N_5994);
or U6217 (N_6217,N_5891,N_5716);
and U6218 (N_6218,N_5789,N_5992);
nor U6219 (N_6219,N_5937,N_5801);
nor U6220 (N_6220,N_5967,N_5715);
nand U6221 (N_6221,N_5921,N_5891);
or U6222 (N_6222,N_5770,N_5874);
nand U6223 (N_6223,N_5757,N_5854);
nor U6224 (N_6224,N_5785,N_5726);
nor U6225 (N_6225,N_5922,N_5753);
or U6226 (N_6226,N_5758,N_5877);
or U6227 (N_6227,N_5947,N_5822);
nor U6228 (N_6228,N_5980,N_5778);
or U6229 (N_6229,N_5985,N_5738);
xor U6230 (N_6230,N_5848,N_5832);
nor U6231 (N_6231,N_5913,N_5947);
or U6232 (N_6232,N_5945,N_5852);
xor U6233 (N_6233,N_5946,N_5816);
xor U6234 (N_6234,N_5872,N_5805);
and U6235 (N_6235,N_5894,N_5835);
or U6236 (N_6236,N_5798,N_5880);
or U6237 (N_6237,N_5715,N_5960);
nor U6238 (N_6238,N_5805,N_5816);
nand U6239 (N_6239,N_5738,N_5752);
nor U6240 (N_6240,N_5816,N_5817);
nand U6241 (N_6241,N_5861,N_5993);
nor U6242 (N_6242,N_5793,N_5953);
and U6243 (N_6243,N_5899,N_5835);
or U6244 (N_6244,N_5888,N_5970);
and U6245 (N_6245,N_5714,N_5720);
xor U6246 (N_6246,N_5921,N_5710);
or U6247 (N_6247,N_5877,N_5936);
nor U6248 (N_6248,N_5881,N_5758);
and U6249 (N_6249,N_5813,N_5773);
nand U6250 (N_6250,N_5874,N_5903);
nand U6251 (N_6251,N_5883,N_5742);
xor U6252 (N_6252,N_5915,N_5758);
nor U6253 (N_6253,N_5934,N_5807);
nand U6254 (N_6254,N_5761,N_5841);
nand U6255 (N_6255,N_5753,N_5718);
and U6256 (N_6256,N_5760,N_5823);
or U6257 (N_6257,N_5944,N_5738);
nor U6258 (N_6258,N_5701,N_5993);
xor U6259 (N_6259,N_5720,N_5771);
or U6260 (N_6260,N_5953,N_5866);
and U6261 (N_6261,N_5767,N_5791);
nor U6262 (N_6262,N_5755,N_5775);
or U6263 (N_6263,N_5847,N_5997);
xnor U6264 (N_6264,N_5700,N_5770);
xnor U6265 (N_6265,N_5806,N_5799);
or U6266 (N_6266,N_5972,N_5788);
nand U6267 (N_6267,N_5767,N_5906);
nor U6268 (N_6268,N_5754,N_5781);
xor U6269 (N_6269,N_5860,N_5779);
nor U6270 (N_6270,N_5986,N_5900);
xor U6271 (N_6271,N_5728,N_5701);
xor U6272 (N_6272,N_5823,N_5938);
nand U6273 (N_6273,N_5734,N_5998);
nand U6274 (N_6274,N_5788,N_5891);
nor U6275 (N_6275,N_5972,N_5810);
or U6276 (N_6276,N_5724,N_5731);
nand U6277 (N_6277,N_5740,N_5830);
nor U6278 (N_6278,N_5887,N_5960);
and U6279 (N_6279,N_5828,N_5966);
and U6280 (N_6280,N_5865,N_5958);
xor U6281 (N_6281,N_5729,N_5980);
and U6282 (N_6282,N_5777,N_5961);
xnor U6283 (N_6283,N_5913,N_5833);
xor U6284 (N_6284,N_5978,N_5879);
nand U6285 (N_6285,N_5700,N_5726);
nor U6286 (N_6286,N_5786,N_5898);
nor U6287 (N_6287,N_5914,N_5714);
nor U6288 (N_6288,N_5959,N_5822);
and U6289 (N_6289,N_5902,N_5787);
nor U6290 (N_6290,N_5985,N_5828);
nand U6291 (N_6291,N_5854,N_5998);
xor U6292 (N_6292,N_5876,N_5774);
xor U6293 (N_6293,N_5814,N_5751);
xnor U6294 (N_6294,N_5960,N_5817);
nor U6295 (N_6295,N_5700,N_5960);
xnor U6296 (N_6296,N_5983,N_5958);
and U6297 (N_6297,N_5988,N_5874);
and U6298 (N_6298,N_5700,N_5756);
or U6299 (N_6299,N_5971,N_5937);
xnor U6300 (N_6300,N_6258,N_6187);
or U6301 (N_6301,N_6201,N_6195);
nor U6302 (N_6302,N_6124,N_6016);
and U6303 (N_6303,N_6086,N_6058);
xnor U6304 (N_6304,N_6205,N_6213);
or U6305 (N_6305,N_6169,N_6050);
xnor U6306 (N_6306,N_6104,N_6222);
or U6307 (N_6307,N_6223,N_6102);
or U6308 (N_6308,N_6158,N_6293);
xor U6309 (N_6309,N_6005,N_6051);
and U6310 (N_6310,N_6029,N_6143);
nor U6311 (N_6311,N_6239,N_6139);
or U6312 (N_6312,N_6234,N_6163);
or U6313 (N_6313,N_6170,N_6210);
xor U6314 (N_6314,N_6140,N_6200);
nor U6315 (N_6315,N_6262,N_6072);
and U6316 (N_6316,N_6007,N_6238);
xor U6317 (N_6317,N_6218,N_6098);
nand U6318 (N_6318,N_6261,N_6144);
nor U6319 (N_6319,N_6003,N_6099);
or U6320 (N_6320,N_6209,N_6105);
and U6321 (N_6321,N_6033,N_6198);
nand U6322 (N_6322,N_6228,N_6037);
or U6323 (N_6323,N_6287,N_6097);
and U6324 (N_6324,N_6288,N_6224);
xor U6325 (N_6325,N_6275,N_6285);
nor U6326 (N_6326,N_6156,N_6214);
nor U6327 (N_6327,N_6296,N_6061);
nor U6328 (N_6328,N_6250,N_6260);
or U6329 (N_6329,N_6088,N_6043);
or U6330 (N_6330,N_6253,N_6161);
and U6331 (N_6331,N_6215,N_6101);
and U6332 (N_6332,N_6068,N_6094);
nand U6333 (N_6333,N_6113,N_6123);
and U6334 (N_6334,N_6028,N_6015);
nand U6335 (N_6335,N_6090,N_6064);
or U6336 (N_6336,N_6298,N_6035);
or U6337 (N_6337,N_6217,N_6268);
or U6338 (N_6338,N_6063,N_6208);
and U6339 (N_6339,N_6236,N_6245);
nand U6340 (N_6340,N_6079,N_6020);
nor U6341 (N_6341,N_6083,N_6279);
or U6342 (N_6342,N_6175,N_6254);
and U6343 (N_6343,N_6100,N_6025);
xor U6344 (N_6344,N_6087,N_6202);
nor U6345 (N_6345,N_6181,N_6011);
or U6346 (N_6346,N_6179,N_6023);
nand U6347 (N_6347,N_6248,N_6030);
nor U6348 (N_6348,N_6045,N_6067);
and U6349 (N_6349,N_6075,N_6252);
and U6350 (N_6350,N_6182,N_6199);
and U6351 (N_6351,N_6203,N_6273);
nor U6352 (N_6352,N_6138,N_6162);
and U6353 (N_6353,N_6227,N_6013);
xnor U6354 (N_6354,N_6184,N_6065);
xor U6355 (N_6355,N_6267,N_6019);
xnor U6356 (N_6356,N_6055,N_6168);
nand U6357 (N_6357,N_6039,N_6080);
and U6358 (N_6358,N_6294,N_6119);
nor U6359 (N_6359,N_6062,N_6111);
xor U6360 (N_6360,N_6042,N_6241);
nand U6361 (N_6361,N_6150,N_6036);
or U6362 (N_6362,N_6280,N_6220);
xor U6363 (N_6363,N_6165,N_6272);
nor U6364 (N_6364,N_6112,N_6106);
or U6365 (N_6365,N_6136,N_6177);
or U6366 (N_6366,N_6004,N_6026);
nand U6367 (N_6367,N_6017,N_6266);
or U6368 (N_6368,N_6257,N_6115);
nor U6369 (N_6369,N_6070,N_6010);
nor U6370 (N_6370,N_6290,N_6247);
and U6371 (N_6371,N_6056,N_6282);
or U6372 (N_6372,N_6071,N_6259);
and U6373 (N_6373,N_6270,N_6103);
nor U6374 (N_6374,N_6242,N_6151);
nand U6375 (N_6375,N_6012,N_6231);
xnor U6376 (N_6376,N_6192,N_6076);
nand U6377 (N_6377,N_6134,N_6135);
xor U6378 (N_6378,N_6281,N_6000);
and U6379 (N_6379,N_6255,N_6246);
and U6380 (N_6380,N_6173,N_6074);
nand U6381 (N_6381,N_6131,N_6263);
nand U6382 (N_6382,N_6093,N_6141);
nand U6383 (N_6383,N_6194,N_6240);
nand U6384 (N_6384,N_6142,N_6292);
and U6385 (N_6385,N_6001,N_6171);
and U6386 (N_6386,N_6132,N_6052);
xnor U6387 (N_6387,N_6256,N_6044);
and U6388 (N_6388,N_6006,N_6225);
nand U6389 (N_6389,N_6002,N_6277);
nor U6390 (N_6390,N_6166,N_6077);
nand U6391 (N_6391,N_6160,N_6085);
nor U6392 (N_6392,N_6137,N_6146);
nor U6393 (N_6393,N_6147,N_6244);
xnor U6394 (N_6394,N_6278,N_6159);
nand U6395 (N_6395,N_6049,N_6289);
and U6396 (N_6396,N_6078,N_6060);
xnor U6397 (N_6397,N_6233,N_6283);
nand U6398 (N_6398,N_6174,N_6186);
xor U6399 (N_6399,N_6054,N_6206);
or U6400 (N_6400,N_6121,N_6073);
nand U6401 (N_6401,N_6107,N_6297);
nand U6402 (N_6402,N_6109,N_6024);
nor U6403 (N_6403,N_6172,N_6133);
xor U6404 (N_6404,N_6230,N_6110);
and U6405 (N_6405,N_6180,N_6092);
nand U6406 (N_6406,N_6114,N_6034);
or U6407 (N_6407,N_6128,N_6229);
or U6408 (N_6408,N_6221,N_6095);
and U6409 (N_6409,N_6040,N_6153);
and U6410 (N_6410,N_6149,N_6126);
nor U6411 (N_6411,N_6021,N_6243);
nor U6412 (N_6412,N_6249,N_6053);
xor U6413 (N_6413,N_6235,N_6108);
and U6414 (N_6414,N_6117,N_6027);
xor U6415 (N_6415,N_6127,N_6274);
or U6416 (N_6416,N_6008,N_6091);
xor U6417 (N_6417,N_6154,N_6059);
or U6418 (N_6418,N_6167,N_6189);
or U6419 (N_6419,N_6069,N_6032);
nor U6420 (N_6420,N_6193,N_6084);
and U6421 (N_6421,N_6145,N_6031);
or U6422 (N_6422,N_6155,N_6157);
or U6423 (N_6423,N_6183,N_6299);
or U6424 (N_6424,N_6178,N_6286);
xnor U6425 (N_6425,N_6265,N_6276);
nand U6426 (N_6426,N_6190,N_6152);
and U6427 (N_6427,N_6219,N_6014);
nand U6428 (N_6428,N_6148,N_6057);
xnor U6429 (N_6429,N_6176,N_6164);
nor U6430 (N_6430,N_6232,N_6116);
or U6431 (N_6431,N_6120,N_6226);
and U6432 (N_6432,N_6048,N_6237);
nand U6433 (N_6433,N_6197,N_6271);
and U6434 (N_6434,N_6047,N_6082);
nand U6435 (N_6435,N_6129,N_6212);
or U6436 (N_6436,N_6204,N_6196);
xnor U6437 (N_6437,N_6207,N_6089);
nor U6438 (N_6438,N_6125,N_6118);
and U6439 (N_6439,N_6269,N_6251);
xor U6440 (N_6440,N_6211,N_6038);
nand U6441 (N_6441,N_6122,N_6291);
nor U6442 (N_6442,N_6264,N_6216);
nor U6443 (N_6443,N_6191,N_6009);
xnor U6444 (N_6444,N_6284,N_6096);
xor U6445 (N_6445,N_6066,N_6081);
or U6446 (N_6446,N_6046,N_6018);
nor U6447 (N_6447,N_6022,N_6185);
or U6448 (N_6448,N_6295,N_6188);
or U6449 (N_6449,N_6041,N_6130);
xnor U6450 (N_6450,N_6269,N_6150);
or U6451 (N_6451,N_6179,N_6036);
nor U6452 (N_6452,N_6217,N_6074);
nand U6453 (N_6453,N_6158,N_6277);
or U6454 (N_6454,N_6043,N_6152);
nor U6455 (N_6455,N_6024,N_6201);
and U6456 (N_6456,N_6046,N_6019);
nand U6457 (N_6457,N_6029,N_6231);
or U6458 (N_6458,N_6117,N_6023);
xnor U6459 (N_6459,N_6054,N_6293);
or U6460 (N_6460,N_6157,N_6132);
and U6461 (N_6461,N_6236,N_6077);
and U6462 (N_6462,N_6286,N_6166);
and U6463 (N_6463,N_6013,N_6298);
nor U6464 (N_6464,N_6233,N_6230);
nand U6465 (N_6465,N_6224,N_6208);
nor U6466 (N_6466,N_6101,N_6049);
nor U6467 (N_6467,N_6233,N_6272);
and U6468 (N_6468,N_6201,N_6093);
or U6469 (N_6469,N_6155,N_6080);
and U6470 (N_6470,N_6291,N_6097);
or U6471 (N_6471,N_6137,N_6071);
xor U6472 (N_6472,N_6151,N_6012);
xnor U6473 (N_6473,N_6072,N_6225);
xor U6474 (N_6474,N_6112,N_6226);
xor U6475 (N_6475,N_6191,N_6130);
and U6476 (N_6476,N_6205,N_6170);
nor U6477 (N_6477,N_6023,N_6106);
nand U6478 (N_6478,N_6122,N_6034);
nand U6479 (N_6479,N_6135,N_6190);
xnor U6480 (N_6480,N_6084,N_6296);
nand U6481 (N_6481,N_6078,N_6153);
nand U6482 (N_6482,N_6168,N_6102);
or U6483 (N_6483,N_6283,N_6051);
or U6484 (N_6484,N_6152,N_6179);
or U6485 (N_6485,N_6157,N_6299);
nand U6486 (N_6486,N_6000,N_6069);
nand U6487 (N_6487,N_6005,N_6191);
nand U6488 (N_6488,N_6195,N_6015);
nand U6489 (N_6489,N_6212,N_6054);
xor U6490 (N_6490,N_6058,N_6029);
nor U6491 (N_6491,N_6149,N_6134);
or U6492 (N_6492,N_6020,N_6220);
nor U6493 (N_6493,N_6068,N_6049);
nand U6494 (N_6494,N_6185,N_6032);
nor U6495 (N_6495,N_6269,N_6215);
nor U6496 (N_6496,N_6098,N_6293);
nand U6497 (N_6497,N_6013,N_6250);
nand U6498 (N_6498,N_6027,N_6197);
xnor U6499 (N_6499,N_6036,N_6041);
or U6500 (N_6500,N_6080,N_6210);
xnor U6501 (N_6501,N_6090,N_6281);
nor U6502 (N_6502,N_6109,N_6072);
nor U6503 (N_6503,N_6238,N_6248);
nor U6504 (N_6504,N_6111,N_6236);
or U6505 (N_6505,N_6231,N_6110);
and U6506 (N_6506,N_6185,N_6056);
xor U6507 (N_6507,N_6241,N_6054);
or U6508 (N_6508,N_6068,N_6268);
xnor U6509 (N_6509,N_6109,N_6067);
or U6510 (N_6510,N_6279,N_6230);
xnor U6511 (N_6511,N_6051,N_6115);
or U6512 (N_6512,N_6036,N_6189);
xnor U6513 (N_6513,N_6117,N_6103);
nor U6514 (N_6514,N_6166,N_6169);
or U6515 (N_6515,N_6136,N_6227);
nand U6516 (N_6516,N_6019,N_6268);
xnor U6517 (N_6517,N_6047,N_6296);
and U6518 (N_6518,N_6232,N_6283);
and U6519 (N_6519,N_6044,N_6116);
xor U6520 (N_6520,N_6121,N_6192);
or U6521 (N_6521,N_6066,N_6254);
nand U6522 (N_6522,N_6260,N_6295);
and U6523 (N_6523,N_6104,N_6265);
nor U6524 (N_6524,N_6040,N_6260);
nand U6525 (N_6525,N_6104,N_6060);
nor U6526 (N_6526,N_6000,N_6122);
nor U6527 (N_6527,N_6029,N_6134);
nor U6528 (N_6528,N_6273,N_6210);
nor U6529 (N_6529,N_6000,N_6106);
xnor U6530 (N_6530,N_6282,N_6223);
nor U6531 (N_6531,N_6098,N_6183);
nand U6532 (N_6532,N_6149,N_6217);
and U6533 (N_6533,N_6095,N_6250);
xnor U6534 (N_6534,N_6254,N_6007);
or U6535 (N_6535,N_6220,N_6231);
xor U6536 (N_6536,N_6202,N_6024);
and U6537 (N_6537,N_6084,N_6107);
or U6538 (N_6538,N_6012,N_6265);
or U6539 (N_6539,N_6147,N_6092);
or U6540 (N_6540,N_6194,N_6051);
xnor U6541 (N_6541,N_6166,N_6248);
xnor U6542 (N_6542,N_6054,N_6254);
nor U6543 (N_6543,N_6263,N_6088);
or U6544 (N_6544,N_6236,N_6260);
nor U6545 (N_6545,N_6157,N_6128);
and U6546 (N_6546,N_6173,N_6213);
nor U6547 (N_6547,N_6024,N_6172);
or U6548 (N_6548,N_6208,N_6018);
or U6549 (N_6549,N_6297,N_6272);
xor U6550 (N_6550,N_6094,N_6164);
and U6551 (N_6551,N_6240,N_6079);
nand U6552 (N_6552,N_6219,N_6292);
nor U6553 (N_6553,N_6086,N_6123);
and U6554 (N_6554,N_6237,N_6268);
xnor U6555 (N_6555,N_6211,N_6271);
or U6556 (N_6556,N_6063,N_6097);
xnor U6557 (N_6557,N_6160,N_6295);
and U6558 (N_6558,N_6045,N_6113);
xnor U6559 (N_6559,N_6229,N_6294);
and U6560 (N_6560,N_6043,N_6228);
and U6561 (N_6561,N_6251,N_6078);
or U6562 (N_6562,N_6278,N_6150);
and U6563 (N_6563,N_6143,N_6134);
or U6564 (N_6564,N_6180,N_6299);
or U6565 (N_6565,N_6127,N_6118);
and U6566 (N_6566,N_6242,N_6194);
nand U6567 (N_6567,N_6123,N_6281);
nor U6568 (N_6568,N_6039,N_6011);
and U6569 (N_6569,N_6009,N_6254);
xnor U6570 (N_6570,N_6136,N_6272);
and U6571 (N_6571,N_6009,N_6087);
nand U6572 (N_6572,N_6296,N_6242);
or U6573 (N_6573,N_6057,N_6077);
nor U6574 (N_6574,N_6091,N_6299);
xor U6575 (N_6575,N_6140,N_6051);
or U6576 (N_6576,N_6263,N_6156);
xnor U6577 (N_6577,N_6228,N_6164);
and U6578 (N_6578,N_6055,N_6135);
and U6579 (N_6579,N_6282,N_6062);
or U6580 (N_6580,N_6075,N_6091);
xor U6581 (N_6581,N_6119,N_6032);
or U6582 (N_6582,N_6113,N_6114);
and U6583 (N_6583,N_6088,N_6122);
nor U6584 (N_6584,N_6213,N_6245);
nand U6585 (N_6585,N_6010,N_6171);
and U6586 (N_6586,N_6251,N_6253);
and U6587 (N_6587,N_6136,N_6159);
and U6588 (N_6588,N_6058,N_6121);
and U6589 (N_6589,N_6085,N_6255);
xnor U6590 (N_6590,N_6274,N_6227);
and U6591 (N_6591,N_6212,N_6118);
and U6592 (N_6592,N_6057,N_6127);
nor U6593 (N_6593,N_6031,N_6102);
and U6594 (N_6594,N_6020,N_6260);
or U6595 (N_6595,N_6216,N_6251);
xor U6596 (N_6596,N_6218,N_6222);
and U6597 (N_6597,N_6001,N_6152);
and U6598 (N_6598,N_6025,N_6126);
and U6599 (N_6599,N_6112,N_6003);
xor U6600 (N_6600,N_6315,N_6549);
nor U6601 (N_6601,N_6550,N_6562);
or U6602 (N_6602,N_6453,N_6538);
or U6603 (N_6603,N_6513,N_6536);
or U6604 (N_6604,N_6370,N_6392);
nor U6605 (N_6605,N_6532,N_6400);
nand U6606 (N_6606,N_6357,N_6423);
nor U6607 (N_6607,N_6335,N_6345);
and U6608 (N_6608,N_6484,N_6332);
and U6609 (N_6609,N_6403,N_6514);
xnor U6610 (N_6610,N_6451,N_6348);
xor U6611 (N_6611,N_6408,N_6437);
nor U6612 (N_6612,N_6316,N_6346);
or U6613 (N_6613,N_6544,N_6504);
xnor U6614 (N_6614,N_6405,N_6509);
nor U6615 (N_6615,N_6448,N_6493);
nand U6616 (N_6616,N_6520,N_6318);
nand U6617 (N_6617,N_6441,N_6341);
and U6618 (N_6618,N_6547,N_6569);
and U6619 (N_6619,N_6465,N_6312);
and U6620 (N_6620,N_6596,N_6548);
or U6621 (N_6621,N_6308,N_6480);
nand U6622 (N_6622,N_6476,N_6352);
and U6623 (N_6623,N_6522,N_6380);
and U6624 (N_6624,N_6545,N_6416);
xor U6625 (N_6625,N_6533,N_6521);
nor U6626 (N_6626,N_6478,N_6310);
nor U6627 (N_6627,N_6580,N_6489);
nor U6628 (N_6628,N_6443,N_6359);
or U6629 (N_6629,N_6563,N_6376);
nor U6630 (N_6630,N_6450,N_6397);
and U6631 (N_6631,N_6436,N_6495);
xor U6632 (N_6632,N_6576,N_6415);
and U6633 (N_6633,N_6586,N_6377);
nor U6634 (N_6634,N_6553,N_6507);
or U6635 (N_6635,N_6502,N_6425);
nor U6636 (N_6636,N_6498,N_6575);
nand U6637 (N_6637,N_6344,N_6467);
nand U6638 (N_6638,N_6428,N_6460);
and U6639 (N_6639,N_6599,N_6390);
and U6640 (N_6640,N_6475,N_6573);
or U6641 (N_6641,N_6379,N_6592);
nor U6642 (N_6642,N_6469,N_6561);
and U6643 (N_6643,N_6517,N_6383);
or U6644 (N_6644,N_6378,N_6358);
and U6645 (N_6645,N_6585,N_6393);
or U6646 (N_6646,N_6481,N_6323);
nand U6647 (N_6647,N_6477,N_6527);
or U6648 (N_6648,N_6395,N_6452);
nand U6649 (N_6649,N_6399,N_6572);
nand U6650 (N_6650,N_6331,N_6447);
and U6651 (N_6651,N_6363,N_6394);
nand U6652 (N_6652,N_6389,N_6410);
nor U6653 (N_6653,N_6307,N_6388);
xor U6654 (N_6654,N_6426,N_6326);
nand U6655 (N_6655,N_6325,N_6472);
nand U6656 (N_6656,N_6420,N_6566);
nor U6657 (N_6657,N_6361,N_6551);
nor U6658 (N_6658,N_6531,N_6558);
xnor U6659 (N_6659,N_6427,N_6540);
and U6660 (N_6660,N_6313,N_6353);
xnor U6661 (N_6661,N_6539,N_6567);
xnor U6662 (N_6662,N_6304,N_6589);
xnor U6663 (N_6663,N_6327,N_6314);
nor U6664 (N_6664,N_6442,N_6446);
or U6665 (N_6665,N_6463,N_6364);
xnor U6666 (N_6666,N_6305,N_6583);
nor U6667 (N_6667,N_6369,N_6356);
nor U6668 (N_6668,N_6497,N_6515);
or U6669 (N_6669,N_6482,N_6577);
nand U6670 (N_6670,N_6508,N_6387);
nor U6671 (N_6671,N_6386,N_6365);
or U6672 (N_6672,N_6505,N_6391);
and U6673 (N_6673,N_6546,N_6320);
nor U6674 (N_6674,N_6457,N_6578);
and U6675 (N_6675,N_6554,N_6455);
and U6676 (N_6676,N_6409,N_6511);
or U6677 (N_6677,N_6375,N_6598);
or U6678 (N_6678,N_6339,N_6584);
and U6679 (N_6679,N_6303,N_6440);
or U6680 (N_6680,N_6556,N_6471);
nand U6681 (N_6681,N_6591,N_6501);
and U6682 (N_6682,N_6535,N_6491);
nor U6683 (N_6683,N_6373,N_6368);
nor U6684 (N_6684,N_6382,N_6581);
nand U6685 (N_6685,N_6338,N_6328);
nor U6686 (N_6686,N_6431,N_6552);
xnor U6687 (N_6687,N_6500,N_6490);
nand U6688 (N_6688,N_6385,N_6433);
or U6689 (N_6689,N_6523,N_6559);
or U6690 (N_6690,N_6530,N_6412);
nor U6691 (N_6691,N_6483,N_6430);
and U6692 (N_6692,N_6496,N_6355);
and U6693 (N_6693,N_6384,N_6449);
xor U6694 (N_6694,N_6454,N_6524);
nand U6695 (N_6695,N_6537,N_6317);
nand U6696 (N_6696,N_6444,N_6518);
and U6697 (N_6697,N_6300,N_6371);
xor U6698 (N_6698,N_6404,N_6564);
nand U6699 (N_6699,N_6445,N_6333);
nand U6700 (N_6700,N_6595,N_6439);
nor U6701 (N_6701,N_6486,N_6506);
or U6702 (N_6702,N_6343,N_6407);
nand U6703 (N_6703,N_6503,N_6555);
and U6704 (N_6704,N_6417,N_6340);
xnor U6705 (N_6705,N_6458,N_6597);
and U6706 (N_6706,N_6485,N_6396);
and U6707 (N_6707,N_6593,N_6588);
and U6708 (N_6708,N_6319,N_6411);
and U6709 (N_6709,N_6324,N_6374);
nor U6710 (N_6710,N_6438,N_6422);
or U6711 (N_6711,N_6462,N_6579);
nand U6712 (N_6712,N_6349,N_6424);
and U6713 (N_6713,N_6487,N_6337);
or U6714 (N_6714,N_6570,N_6526);
xor U6715 (N_6715,N_6429,N_6435);
and U6716 (N_6716,N_6468,N_6510);
nor U6717 (N_6717,N_6329,N_6470);
xnor U6718 (N_6718,N_6402,N_6414);
and U6719 (N_6719,N_6574,N_6499);
nor U6720 (N_6720,N_6366,N_6587);
xor U6721 (N_6721,N_6519,N_6398);
nand U6722 (N_6722,N_6473,N_6354);
xor U6723 (N_6723,N_6434,N_6492);
nand U6724 (N_6724,N_6322,N_6309);
or U6725 (N_6725,N_6419,N_6512);
nor U6726 (N_6726,N_6311,N_6418);
or U6727 (N_6727,N_6456,N_6381);
and U6728 (N_6728,N_6406,N_6565);
and U6729 (N_6729,N_6541,N_6302);
xor U6730 (N_6730,N_6362,N_6543);
xnor U6731 (N_6731,N_6528,N_6474);
xnor U6732 (N_6732,N_6334,N_6571);
or U6733 (N_6733,N_6488,N_6494);
and U6734 (N_6734,N_6367,N_6330);
xnor U6735 (N_6735,N_6432,N_6479);
xnor U6736 (N_6736,N_6568,N_6560);
nand U6737 (N_6737,N_6516,N_6464);
and U6738 (N_6738,N_6401,N_6321);
or U6739 (N_6739,N_6413,N_6557);
and U6740 (N_6740,N_6590,N_6534);
or U6741 (N_6741,N_6360,N_6529);
nor U6742 (N_6742,N_6306,N_6421);
nand U6743 (N_6743,N_6350,N_6542);
xor U6744 (N_6744,N_6466,N_6582);
nor U6745 (N_6745,N_6347,N_6594);
nand U6746 (N_6746,N_6342,N_6525);
nand U6747 (N_6747,N_6301,N_6459);
nor U6748 (N_6748,N_6372,N_6351);
and U6749 (N_6749,N_6336,N_6461);
or U6750 (N_6750,N_6578,N_6539);
and U6751 (N_6751,N_6512,N_6498);
or U6752 (N_6752,N_6567,N_6444);
xor U6753 (N_6753,N_6382,N_6527);
or U6754 (N_6754,N_6496,N_6304);
nand U6755 (N_6755,N_6379,N_6575);
xnor U6756 (N_6756,N_6509,N_6344);
and U6757 (N_6757,N_6591,N_6520);
nor U6758 (N_6758,N_6306,N_6440);
nor U6759 (N_6759,N_6497,N_6549);
or U6760 (N_6760,N_6370,N_6574);
xnor U6761 (N_6761,N_6532,N_6418);
or U6762 (N_6762,N_6495,N_6340);
or U6763 (N_6763,N_6506,N_6443);
and U6764 (N_6764,N_6480,N_6309);
nand U6765 (N_6765,N_6425,N_6304);
nor U6766 (N_6766,N_6515,N_6304);
and U6767 (N_6767,N_6504,N_6586);
nand U6768 (N_6768,N_6492,N_6557);
and U6769 (N_6769,N_6568,N_6306);
and U6770 (N_6770,N_6362,N_6467);
nand U6771 (N_6771,N_6570,N_6490);
and U6772 (N_6772,N_6462,N_6488);
xor U6773 (N_6773,N_6351,N_6404);
or U6774 (N_6774,N_6525,N_6353);
nand U6775 (N_6775,N_6463,N_6441);
and U6776 (N_6776,N_6399,N_6389);
or U6777 (N_6777,N_6434,N_6502);
nor U6778 (N_6778,N_6311,N_6403);
nand U6779 (N_6779,N_6330,N_6541);
or U6780 (N_6780,N_6300,N_6537);
and U6781 (N_6781,N_6318,N_6353);
nand U6782 (N_6782,N_6567,N_6463);
and U6783 (N_6783,N_6494,N_6504);
nor U6784 (N_6784,N_6331,N_6365);
and U6785 (N_6785,N_6450,N_6548);
nor U6786 (N_6786,N_6369,N_6368);
or U6787 (N_6787,N_6529,N_6511);
nor U6788 (N_6788,N_6595,N_6552);
nand U6789 (N_6789,N_6486,N_6461);
and U6790 (N_6790,N_6526,N_6473);
xnor U6791 (N_6791,N_6418,N_6366);
xnor U6792 (N_6792,N_6485,N_6521);
nand U6793 (N_6793,N_6371,N_6516);
xor U6794 (N_6794,N_6350,N_6343);
nand U6795 (N_6795,N_6317,N_6318);
nor U6796 (N_6796,N_6329,N_6575);
and U6797 (N_6797,N_6471,N_6308);
xnor U6798 (N_6798,N_6557,N_6572);
xnor U6799 (N_6799,N_6326,N_6470);
or U6800 (N_6800,N_6472,N_6465);
xor U6801 (N_6801,N_6454,N_6341);
or U6802 (N_6802,N_6490,N_6447);
nor U6803 (N_6803,N_6568,N_6445);
nor U6804 (N_6804,N_6545,N_6593);
nor U6805 (N_6805,N_6528,N_6553);
nand U6806 (N_6806,N_6508,N_6505);
nor U6807 (N_6807,N_6418,N_6500);
nand U6808 (N_6808,N_6467,N_6492);
and U6809 (N_6809,N_6423,N_6410);
nand U6810 (N_6810,N_6539,N_6409);
xor U6811 (N_6811,N_6506,N_6467);
xor U6812 (N_6812,N_6506,N_6569);
xor U6813 (N_6813,N_6542,N_6473);
nand U6814 (N_6814,N_6313,N_6567);
xnor U6815 (N_6815,N_6476,N_6396);
xor U6816 (N_6816,N_6580,N_6410);
xor U6817 (N_6817,N_6361,N_6477);
and U6818 (N_6818,N_6402,N_6466);
nand U6819 (N_6819,N_6484,N_6428);
and U6820 (N_6820,N_6387,N_6474);
xnor U6821 (N_6821,N_6337,N_6524);
nor U6822 (N_6822,N_6591,N_6551);
or U6823 (N_6823,N_6542,N_6372);
xnor U6824 (N_6824,N_6373,N_6443);
nor U6825 (N_6825,N_6332,N_6477);
nor U6826 (N_6826,N_6519,N_6518);
nand U6827 (N_6827,N_6473,N_6323);
xnor U6828 (N_6828,N_6457,N_6303);
or U6829 (N_6829,N_6477,N_6358);
or U6830 (N_6830,N_6392,N_6321);
nor U6831 (N_6831,N_6599,N_6590);
xor U6832 (N_6832,N_6374,N_6378);
nor U6833 (N_6833,N_6567,N_6333);
or U6834 (N_6834,N_6378,N_6311);
or U6835 (N_6835,N_6428,N_6423);
nor U6836 (N_6836,N_6392,N_6376);
xor U6837 (N_6837,N_6525,N_6387);
nand U6838 (N_6838,N_6557,N_6527);
and U6839 (N_6839,N_6432,N_6472);
or U6840 (N_6840,N_6302,N_6326);
nand U6841 (N_6841,N_6358,N_6394);
nand U6842 (N_6842,N_6494,N_6498);
xnor U6843 (N_6843,N_6558,N_6476);
nor U6844 (N_6844,N_6546,N_6326);
nor U6845 (N_6845,N_6569,N_6596);
nor U6846 (N_6846,N_6486,N_6368);
and U6847 (N_6847,N_6342,N_6454);
nor U6848 (N_6848,N_6439,N_6388);
or U6849 (N_6849,N_6405,N_6514);
xnor U6850 (N_6850,N_6493,N_6411);
xor U6851 (N_6851,N_6348,N_6464);
or U6852 (N_6852,N_6501,N_6544);
nor U6853 (N_6853,N_6529,N_6598);
xor U6854 (N_6854,N_6398,N_6471);
or U6855 (N_6855,N_6359,N_6337);
nand U6856 (N_6856,N_6456,N_6414);
nand U6857 (N_6857,N_6546,N_6332);
nor U6858 (N_6858,N_6344,N_6334);
and U6859 (N_6859,N_6474,N_6370);
and U6860 (N_6860,N_6535,N_6315);
xor U6861 (N_6861,N_6435,N_6378);
or U6862 (N_6862,N_6557,N_6411);
and U6863 (N_6863,N_6577,N_6559);
and U6864 (N_6864,N_6518,N_6389);
nor U6865 (N_6865,N_6454,N_6470);
and U6866 (N_6866,N_6435,N_6558);
or U6867 (N_6867,N_6517,N_6439);
and U6868 (N_6868,N_6599,N_6589);
nor U6869 (N_6869,N_6345,N_6476);
or U6870 (N_6870,N_6567,N_6322);
and U6871 (N_6871,N_6595,N_6401);
or U6872 (N_6872,N_6395,N_6380);
nand U6873 (N_6873,N_6367,N_6410);
nand U6874 (N_6874,N_6579,N_6373);
and U6875 (N_6875,N_6379,N_6337);
or U6876 (N_6876,N_6585,N_6495);
and U6877 (N_6877,N_6384,N_6558);
nor U6878 (N_6878,N_6566,N_6427);
xnor U6879 (N_6879,N_6385,N_6328);
nor U6880 (N_6880,N_6515,N_6548);
nor U6881 (N_6881,N_6305,N_6467);
or U6882 (N_6882,N_6598,N_6503);
xnor U6883 (N_6883,N_6553,N_6546);
xnor U6884 (N_6884,N_6436,N_6581);
and U6885 (N_6885,N_6365,N_6349);
or U6886 (N_6886,N_6400,N_6513);
xor U6887 (N_6887,N_6328,N_6376);
nand U6888 (N_6888,N_6498,N_6360);
and U6889 (N_6889,N_6344,N_6321);
or U6890 (N_6890,N_6343,N_6546);
xnor U6891 (N_6891,N_6386,N_6471);
nor U6892 (N_6892,N_6448,N_6537);
and U6893 (N_6893,N_6450,N_6419);
or U6894 (N_6894,N_6352,N_6416);
and U6895 (N_6895,N_6595,N_6357);
xor U6896 (N_6896,N_6574,N_6529);
xnor U6897 (N_6897,N_6545,N_6318);
and U6898 (N_6898,N_6395,N_6324);
nor U6899 (N_6899,N_6352,N_6415);
xnor U6900 (N_6900,N_6618,N_6602);
xnor U6901 (N_6901,N_6712,N_6798);
xor U6902 (N_6902,N_6747,N_6858);
and U6903 (N_6903,N_6878,N_6720);
or U6904 (N_6904,N_6845,N_6795);
or U6905 (N_6905,N_6663,N_6743);
and U6906 (N_6906,N_6695,N_6642);
or U6907 (N_6907,N_6761,N_6862);
xor U6908 (N_6908,N_6813,N_6716);
nor U6909 (N_6909,N_6652,N_6792);
and U6910 (N_6910,N_6880,N_6802);
or U6911 (N_6911,N_6861,N_6779);
or U6912 (N_6912,N_6699,N_6814);
nand U6913 (N_6913,N_6824,N_6776);
nor U6914 (N_6914,N_6848,N_6696);
nor U6915 (N_6915,N_6611,N_6883);
or U6916 (N_6916,N_6751,N_6809);
and U6917 (N_6917,N_6886,N_6619);
and U6918 (N_6918,N_6650,N_6781);
xor U6919 (N_6919,N_6784,N_6614);
nor U6920 (N_6920,N_6896,N_6885);
and U6921 (N_6921,N_6752,N_6756);
nor U6922 (N_6922,N_6662,N_6853);
or U6923 (N_6923,N_6797,N_6732);
or U6924 (N_6924,N_6622,N_6887);
nor U6925 (N_6925,N_6729,N_6874);
or U6926 (N_6926,N_6616,N_6791);
or U6927 (N_6927,N_6839,N_6893);
or U6928 (N_6928,N_6777,N_6855);
and U6929 (N_6929,N_6664,N_6669);
xnor U6930 (N_6930,N_6681,N_6897);
nand U6931 (N_6931,N_6682,N_6725);
xor U6932 (N_6932,N_6627,N_6649);
nand U6933 (N_6933,N_6694,N_6804);
nor U6934 (N_6934,N_6786,N_6709);
or U6935 (N_6935,N_6608,N_6647);
nand U6936 (N_6936,N_6692,N_6783);
or U6937 (N_6937,N_6688,N_6875);
nor U6938 (N_6938,N_6676,N_6641);
nand U6939 (N_6939,N_6705,N_6758);
nand U6940 (N_6940,N_6631,N_6739);
xnor U6941 (N_6941,N_6854,N_6634);
nand U6942 (N_6942,N_6717,N_6640);
or U6943 (N_6943,N_6668,N_6762);
nand U6944 (N_6944,N_6866,N_6841);
or U6945 (N_6945,N_6749,N_6811);
or U6946 (N_6946,N_6844,N_6852);
nor U6947 (N_6947,N_6726,N_6721);
nand U6948 (N_6948,N_6819,N_6630);
nand U6949 (N_6949,N_6706,N_6697);
and U6950 (N_6950,N_6693,N_6778);
xor U6951 (N_6951,N_6701,N_6617);
xor U6952 (N_6952,N_6863,N_6680);
xor U6953 (N_6953,N_6864,N_6820);
xnor U6954 (N_6954,N_6823,N_6628);
or U6955 (N_6955,N_6757,N_6765);
nand U6956 (N_6956,N_6808,N_6801);
and U6957 (N_6957,N_6828,N_6713);
and U6958 (N_6958,N_6655,N_6629);
or U6959 (N_6959,N_6737,N_6719);
or U6960 (N_6960,N_6633,N_6736);
xor U6961 (N_6961,N_6796,N_6788);
nand U6962 (N_6962,N_6755,N_6715);
xnor U6963 (N_6963,N_6645,N_6759);
and U6964 (N_6964,N_6888,N_6865);
and U6965 (N_6965,N_6800,N_6790);
nor U6966 (N_6966,N_6637,N_6882);
or U6967 (N_6967,N_6687,N_6621);
xor U6968 (N_6968,N_6700,N_6689);
or U6969 (N_6969,N_6607,N_6876);
xnor U6970 (N_6970,N_6771,N_6683);
xnor U6971 (N_6971,N_6872,N_6895);
xor U6972 (N_6972,N_6812,N_6856);
xor U6973 (N_6973,N_6685,N_6774);
or U6974 (N_6974,N_6821,N_6766);
xor U6975 (N_6975,N_6837,N_6710);
or U6976 (N_6976,N_6723,N_6834);
nor U6977 (N_6977,N_6859,N_6659);
xor U6978 (N_6978,N_6750,N_6738);
and U6979 (N_6979,N_6868,N_6632);
nand U6980 (N_6980,N_6870,N_6826);
nor U6981 (N_6981,N_6773,N_6780);
or U6982 (N_6982,N_6609,N_6840);
nand U6983 (N_6983,N_6770,N_6742);
xnor U6984 (N_6984,N_6799,N_6711);
nor U6985 (N_6985,N_6782,N_6651);
and U6986 (N_6986,N_6601,N_6829);
xor U6987 (N_6987,N_6772,N_6636);
xnor U6988 (N_6988,N_6658,N_6623);
xor U6989 (N_6989,N_6787,N_6753);
or U6990 (N_6990,N_6625,N_6793);
nand U6991 (N_6991,N_6600,N_6832);
and U6992 (N_6992,N_6830,N_6661);
or U6993 (N_6993,N_6789,N_6892);
xnor U6994 (N_6994,N_6653,N_6794);
nand U6995 (N_6995,N_6679,N_6889);
nor U6996 (N_6996,N_6842,N_6718);
nand U6997 (N_6997,N_6702,N_6769);
or U6998 (N_6998,N_6672,N_6741);
and U6999 (N_6999,N_6724,N_6833);
or U7000 (N_7000,N_6644,N_6894);
nand U7001 (N_7001,N_6815,N_6740);
and U7002 (N_7002,N_6704,N_6860);
nand U7003 (N_7003,N_6635,N_6898);
nor U7004 (N_7004,N_6703,N_6657);
nor U7005 (N_7005,N_6646,N_6639);
or U7006 (N_7006,N_6825,N_6744);
nand U7007 (N_7007,N_6890,N_6691);
and U7008 (N_7008,N_6831,N_6748);
or U7009 (N_7009,N_6822,N_6670);
and U7010 (N_7010,N_6728,N_6610);
and U7011 (N_7011,N_6764,N_6730);
or U7012 (N_7012,N_6722,N_6899);
nand U7013 (N_7013,N_6674,N_6612);
xnor U7014 (N_7014,N_6684,N_6806);
and U7015 (N_7015,N_6671,N_6768);
nand U7016 (N_7016,N_6817,N_6707);
and U7017 (N_7017,N_6869,N_6698);
or U7018 (N_7018,N_6775,N_6803);
and U7019 (N_7019,N_6615,N_6656);
or U7020 (N_7020,N_6818,N_6603);
nand U7021 (N_7021,N_6624,N_6708);
xor U7022 (N_7022,N_6849,N_6666);
or U7023 (N_7023,N_6827,N_6835);
nand U7024 (N_7024,N_6760,N_6648);
or U7025 (N_7025,N_6667,N_6604);
or U7026 (N_7026,N_6626,N_6733);
xor U7027 (N_7027,N_6620,N_6785);
xnor U7028 (N_7028,N_6665,N_6810);
xnor U7029 (N_7029,N_6884,N_6605);
nor U7030 (N_7030,N_6838,N_6678);
nand U7031 (N_7031,N_6686,N_6843);
nor U7032 (N_7032,N_6727,N_6613);
nor U7033 (N_7033,N_6871,N_6731);
or U7034 (N_7034,N_6735,N_6654);
nor U7035 (N_7035,N_6879,N_6606);
or U7036 (N_7036,N_6805,N_6877);
nor U7037 (N_7037,N_6660,N_6675);
nor U7038 (N_7038,N_6690,N_6836);
nor U7039 (N_7039,N_6847,N_6857);
and U7040 (N_7040,N_6673,N_6846);
and U7041 (N_7041,N_6891,N_6643);
or U7042 (N_7042,N_6867,N_6807);
and U7043 (N_7043,N_6714,N_6763);
and U7044 (N_7044,N_6734,N_6850);
xor U7045 (N_7045,N_6767,N_6754);
xnor U7046 (N_7046,N_6881,N_6851);
nand U7047 (N_7047,N_6873,N_6745);
xnor U7048 (N_7048,N_6677,N_6746);
nor U7049 (N_7049,N_6638,N_6816);
xor U7050 (N_7050,N_6731,N_6720);
nand U7051 (N_7051,N_6714,N_6601);
xor U7052 (N_7052,N_6725,N_6832);
nand U7053 (N_7053,N_6796,N_6676);
and U7054 (N_7054,N_6834,N_6884);
and U7055 (N_7055,N_6682,N_6777);
xnor U7056 (N_7056,N_6863,N_6641);
nand U7057 (N_7057,N_6726,N_6627);
xnor U7058 (N_7058,N_6836,N_6703);
nand U7059 (N_7059,N_6776,N_6663);
nand U7060 (N_7060,N_6846,N_6768);
nor U7061 (N_7061,N_6762,N_6658);
nand U7062 (N_7062,N_6685,N_6749);
nor U7063 (N_7063,N_6784,N_6602);
nand U7064 (N_7064,N_6652,N_6676);
xor U7065 (N_7065,N_6632,N_6711);
and U7066 (N_7066,N_6648,N_6886);
or U7067 (N_7067,N_6766,N_6780);
nor U7068 (N_7068,N_6643,N_6721);
xnor U7069 (N_7069,N_6678,N_6655);
nand U7070 (N_7070,N_6804,N_6677);
and U7071 (N_7071,N_6730,N_6645);
nand U7072 (N_7072,N_6809,N_6640);
and U7073 (N_7073,N_6784,N_6832);
nor U7074 (N_7074,N_6611,N_6683);
or U7075 (N_7075,N_6625,N_6629);
xnor U7076 (N_7076,N_6788,N_6828);
nor U7077 (N_7077,N_6755,N_6639);
nor U7078 (N_7078,N_6722,N_6836);
nor U7079 (N_7079,N_6657,N_6753);
xor U7080 (N_7080,N_6818,N_6765);
nand U7081 (N_7081,N_6801,N_6790);
xor U7082 (N_7082,N_6682,N_6808);
nand U7083 (N_7083,N_6626,N_6631);
and U7084 (N_7084,N_6776,N_6734);
and U7085 (N_7085,N_6653,N_6835);
or U7086 (N_7086,N_6798,N_6739);
nand U7087 (N_7087,N_6804,N_6798);
nor U7088 (N_7088,N_6607,N_6869);
and U7089 (N_7089,N_6768,N_6826);
nor U7090 (N_7090,N_6811,N_6875);
nand U7091 (N_7091,N_6727,N_6607);
nand U7092 (N_7092,N_6736,N_6804);
or U7093 (N_7093,N_6858,N_6625);
or U7094 (N_7094,N_6781,N_6655);
xnor U7095 (N_7095,N_6873,N_6601);
nor U7096 (N_7096,N_6849,N_6732);
and U7097 (N_7097,N_6764,N_6697);
nor U7098 (N_7098,N_6773,N_6602);
and U7099 (N_7099,N_6671,N_6601);
or U7100 (N_7100,N_6853,N_6765);
nand U7101 (N_7101,N_6600,N_6866);
and U7102 (N_7102,N_6852,N_6745);
xnor U7103 (N_7103,N_6851,N_6825);
or U7104 (N_7104,N_6680,N_6782);
xnor U7105 (N_7105,N_6749,N_6728);
xor U7106 (N_7106,N_6863,N_6878);
nor U7107 (N_7107,N_6897,N_6872);
nand U7108 (N_7108,N_6616,N_6656);
nor U7109 (N_7109,N_6640,N_6790);
nor U7110 (N_7110,N_6791,N_6856);
or U7111 (N_7111,N_6704,N_6749);
nand U7112 (N_7112,N_6793,N_6893);
or U7113 (N_7113,N_6604,N_6854);
xor U7114 (N_7114,N_6841,N_6855);
xnor U7115 (N_7115,N_6698,N_6753);
nor U7116 (N_7116,N_6733,N_6717);
and U7117 (N_7117,N_6877,N_6754);
xor U7118 (N_7118,N_6829,N_6690);
nand U7119 (N_7119,N_6823,N_6873);
nand U7120 (N_7120,N_6623,N_6826);
nand U7121 (N_7121,N_6770,N_6799);
nor U7122 (N_7122,N_6746,N_6798);
and U7123 (N_7123,N_6882,N_6838);
or U7124 (N_7124,N_6849,N_6706);
nand U7125 (N_7125,N_6794,N_6609);
and U7126 (N_7126,N_6847,N_6698);
xor U7127 (N_7127,N_6709,N_6653);
nor U7128 (N_7128,N_6845,N_6666);
or U7129 (N_7129,N_6769,N_6745);
nor U7130 (N_7130,N_6899,N_6881);
nand U7131 (N_7131,N_6604,N_6600);
nor U7132 (N_7132,N_6612,N_6889);
xnor U7133 (N_7133,N_6820,N_6636);
and U7134 (N_7134,N_6781,N_6735);
or U7135 (N_7135,N_6637,N_6782);
nand U7136 (N_7136,N_6671,N_6778);
nor U7137 (N_7137,N_6675,N_6777);
nand U7138 (N_7138,N_6881,N_6810);
and U7139 (N_7139,N_6898,N_6784);
and U7140 (N_7140,N_6797,N_6883);
or U7141 (N_7141,N_6767,N_6691);
xnor U7142 (N_7142,N_6870,N_6874);
nor U7143 (N_7143,N_6688,N_6670);
nand U7144 (N_7144,N_6714,N_6855);
nor U7145 (N_7145,N_6614,N_6731);
xnor U7146 (N_7146,N_6671,N_6871);
xor U7147 (N_7147,N_6885,N_6672);
xnor U7148 (N_7148,N_6771,N_6883);
nor U7149 (N_7149,N_6637,N_6869);
xnor U7150 (N_7150,N_6879,N_6757);
nor U7151 (N_7151,N_6749,N_6898);
xnor U7152 (N_7152,N_6620,N_6699);
or U7153 (N_7153,N_6761,N_6753);
nand U7154 (N_7154,N_6850,N_6888);
and U7155 (N_7155,N_6884,N_6613);
or U7156 (N_7156,N_6691,N_6754);
and U7157 (N_7157,N_6687,N_6638);
and U7158 (N_7158,N_6621,N_6688);
nor U7159 (N_7159,N_6861,N_6618);
and U7160 (N_7160,N_6731,N_6752);
nor U7161 (N_7161,N_6825,N_6868);
and U7162 (N_7162,N_6718,N_6774);
or U7163 (N_7163,N_6820,N_6712);
or U7164 (N_7164,N_6618,N_6879);
nor U7165 (N_7165,N_6639,N_6863);
nand U7166 (N_7166,N_6725,N_6660);
nor U7167 (N_7167,N_6813,N_6759);
or U7168 (N_7168,N_6810,N_6877);
xor U7169 (N_7169,N_6690,N_6882);
xnor U7170 (N_7170,N_6876,N_6706);
or U7171 (N_7171,N_6635,N_6665);
or U7172 (N_7172,N_6891,N_6719);
or U7173 (N_7173,N_6762,N_6815);
xor U7174 (N_7174,N_6808,N_6857);
nor U7175 (N_7175,N_6847,N_6763);
nand U7176 (N_7176,N_6681,N_6614);
nor U7177 (N_7177,N_6868,N_6607);
nor U7178 (N_7178,N_6646,N_6669);
nor U7179 (N_7179,N_6871,N_6844);
and U7180 (N_7180,N_6634,N_6876);
xor U7181 (N_7181,N_6679,N_6817);
nand U7182 (N_7182,N_6787,N_6659);
nand U7183 (N_7183,N_6622,N_6643);
xnor U7184 (N_7184,N_6780,N_6852);
xnor U7185 (N_7185,N_6774,N_6819);
xnor U7186 (N_7186,N_6659,N_6843);
and U7187 (N_7187,N_6639,N_6762);
nor U7188 (N_7188,N_6669,N_6827);
nand U7189 (N_7189,N_6811,N_6790);
and U7190 (N_7190,N_6720,N_6747);
and U7191 (N_7191,N_6653,N_6854);
xnor U7192 (N_7192,N_6874,N_6780);
nor U7193 (N_7193,N_6849,N_6709);
and U7194 (N_7194,N_6863,N_6708);
nor U7195 (N_7195,N_6746,N_6827);
or U7196 (N_7196,N_6668,N_6767);
or U7197 (N_7197,N_6712,N_6898);
xnor U7198 (N_7198,N_6712,N_6698);
nand U7199 (N_7199,N_6765,N_6600);
nor U7200 (N_7200,N_7135,N_6965);
nand U7201 (N_7201,N_6996,N_7072);
or U7202 (N_7202,N_6946,N_7086);
xor U7203 (N_7203,N_7159,N_6909);
nor U7204 (N_7204,N_7031,N_6939);
nor U7205 (N_7205,N_6984,N_7105);
and U7206 (N_7206,N_6917,N_7060);
xnor U7207 (N_7207,N_7134,N_7172);
xor U7208 (N_7208,N_6948,N_7011);
nand U7209 (N_7209,N_7118,N_7010);
nor U7210 (N_7210,N_7085,N_7115);
xnor U7211 (N_7211,N_6980,N_6911);
nand U7212 (N_7212,N_7145,N_7052);
xnor U7213 (N_7213,N_7157,N_7186);
or U7214 (N_7214,N_7065,N_6925);
and U7215 (N_7215,N_7035,N_7191);
nand U7216 (N_7216,N_7196,N_7067);
or U7217 (N_7217,N_6972,N_6924);
nor U7218 (N_7218,N_7198,N_7151);
nor U7219 (N_7219,N_7043,N_6932);
xnor U7220 (N_7220,N_7189,N_7055);
nor U7221 (N_7221,N_7032,N_6971);
or U7222 (N_7222,N_6906,N_7082);
and U7223 (N_7223,N_6966,N_6983);
and U7224 (N_7224,N_6926,N_6931);
nor U7225 (N_7225,N_7113,N_6910);
xnor U7226 (N_7226,N_7136,N_7155);
or U7227 (N_7227,N_7164,N_7027);
xor U7228 (N_7228,N_7018,N_7139);
xnor U7229 (N_7229,N_7161,N_7039);
or U7230 (N_7230,N_7014,N_7061);
and U7231 (N_7231,N_6991,N_7177);
nor U7232 (N_7232,N_6944,N_7071);
xor U7233 (N_7233,N_7131,N_7003);
nand U7234 (N_7234,N_7179,N_6901);
xor U7235 (N_7235,N_6949,N_7128);
xnor U7236 (N_7236,N_7048,N_6973);
nor U7237 (N_7237,N_6905,N_7079);
or U7238 (N_7238,N_6958,N_7144);
nor U7239 (N_7239,N_6954,N_7021);
or U7240 (N_7240,N_7044,N_7034);
nand U7241 (N_7241,N_7025,N_7049);
xor U7242 (N_7242,N_7023,N_7024);
xnor U7243 (N_7243,N_7175,N_7037);
nand U7244 (N_7244,N_6968,N_6908);
or U7245 (N_7245,N_7167,N_7080);
and U7246 (N_7246,N_6959,N_6900);
xor U7247 (N_7247,N_7069,N_7095);
nor U7248 (N_7248,N_7009,N_7109);
or U7249 (N_7249,N_7162,N_7087);
nor U7250 (N_7250,N_7042,N_6919);
nor U7251 (N_7251,N_6930,N_7022);
nor U7252 (N_7252,N_7068,N_6953);
or U7253 (N_7253,N_6995,N_7070);
xnor U7254 (N_7254,N_7020,N_6975);
or U7255 (N_7255,N_7094,N_6903);
nor U7256 (N_7256,N_6934,N_7148);
or U7257 (N_7257,N_6982,N_7103);
nor U7258 (N_7258,N_6981,N_7053);
nand U7259 (N_7259,N_7193,N_7182);
nor U7260 (N_7260,N_7093,N_7026);
and U7261 (N_7261,N_6902,N_6988);
nand U7262 (N_7262,N_7168,N_6912);
xor U7263 (N_7263,N_7058,N_7047);
and U7264 (N_7264,N_6913,N_7013);
nand U7265 (N_7265,N_7123,N_6969);
xnor U7266 (N_7266,N_6951,N_7045);
nor U7267 (N_7267,N_7000,N_6952);
and U7268 (N_7268,N_7074,N_6941);
nor U7269 (N_7269,N_7137,N_7108);
xor U7270 (N_7270,N_7028,N_7064);
and U7271 (N_7271,N_7110,N_7119);
nor U7272 (N_7272,N_7130,N_7019);
or U7273 (N_7273,N_7180,N_7176);
or U7274 (N_7274,N_7138,N_7133);
xor U7275 (N_7275,N_7102,N_7008);
nand U7276 (N_7276,N_6938,N_7152);
and U7277 (N_7277,N_6997,N_7017);
xor U7278 (N_7278,N_7001,N_7147);
and U7279 (N_7279,N_7101,N_7190);
or U7280 (N_7280,N_7051,N_6955);
and U7281 (N_7281,N_7050,N_6937);
nor U7282 (N_7282,N_6921,N_7142);
xnor U7283 (N_7283,N_6950,N_7059);
xor U7284 (N_7284,N_6945,N_7041);
and U7285 (N_7285,N_6956,N_7156);
nand U7286 (N_7286,N_7170,N_7036);
nor U7287 (N_7287,N_6947,N_6923);
nor U7288 (N_7288,N_7088,N_6993);
nand U7289 (N_7289,N_6986,N_6967);
nor U7290 (N_7290,N_7154,N_6994);
nand U7291 (N_7291,N_7063,N_7120);
or U7292 (N_7292,N_7054,N_7140);
nor U7293 (N_7293,N_6920,N_7089);
xor U7294 (N_7294,N_7184,N_7197);
or U7295 (N_7295,N_6987,N_7038);
xor U7296 (N_7296,N_6915,N_7153);
xor U7297 (N_7297,N_7199,N_6914);
nor U7298 (N_7298,N_7016,N_7073);
or U7299 (N_7299,N_6974,N_6977);
nor U7300 (N_7300,N_7158,N_7097);
nand U7301 (N_7301,N_6998,N_6929);
nand U7302 (N_7302,N_7090,N_7132);
nand U7303 (N_7303,N_7091,N_7005);
and U7304 (N_7304,N_6961,N_7185);
nor U7305 (N_7305,N_6999,N_6927);
and U7306 (N_7306,N_6916,N_6935);
and U7307 (N_7307,N_7124,N_7116);
nor U7308 (N_7308,N_6989,N_6940);
or U7309 (N_7309,N_7057,N_7081);
and U7310 (N_7310,N_7015,N_7146);
or U7311 (N_7311,N_7117,N_7149);
nand U7312 (N_7312,N_7127,N_7173);
nand U7313 (N_7313,N_7106,N_7046);
nand U7314 (N_7314,N_7030,N_7084);
nor U7315 (N_7315,N_6942,N_7078);
xor U7316 (N_7316,N_7029,N_7112);
nor U7317 (N_7317,N_7100,N_7040);
nand U7318 (N_7318,N_7181,N_6907);
xnor U7319 (N_7319,N_7096,N_7092);
nand U7320 (N_7320,N_7006,N_7150);
or U7321 (N_7321,N_7122,N_7076);
nor U7322 (N_7322,N_7194,N_7174);
and U7323 (N_7323,N_7114,N_7099);
and U7324 (N_7324,N_7187,N_6970);
nand U7325 (N_7325,N_7125,N_7160);
nand U7326 (N_7326,N_6963,N_7007);
xor U7327 (N_7327,N_7066,N_6943);
xnor U7328 (N_7328,N_6979,N_6918);
nand U7329 (N_7329,N_7056,N_7012);
nand U7330 (N_7330,N_7083,N_7107);
xnor U7331 (N_7331,N_6904,N_7126);
nor U7332 (N_7332,N_6933,N_7129);
or U7333 (N_7333,N_7171,N_7192);
xor U7334 (N_7334,N_7002,N_7111);
nor U7335 (N_7335,N_7163,N_7141);
or U7336 (N_7336,N_6985,N_6960);
nand U7337 (N_7337,N_7104,N_6922);
and U7338 (N_7338,N_7166,N_7183);
and U7339 (N_7339,N_7169,N_7033);
xor U7340 (N_7340,N_7004,N_6962);
or U7341 (N_7341,N_7075,N_7143);
xor U7342 (N_7342,N_6990,N_7165);
and U7343 (N_7343,N_6976,N_7077);
nor U7344 (N_7344,N_6928,N_6978);
nand U7345 (N_7345,N_7062,N_7188);
nor U7346 (N_7346,N_6964,N_6957);
or U7347 (N_7347,N_6936,N_7121);
nor U7348 (N_7348,N_7195,N_6992);
nand U7349 (N_7349,N_7098,N_7178);
nor U7350 (N_7350,N_6959,N_7070);
and U7351 (N_7351,N_7161,N_7072);
nor U7352 (N_7352,N_7151,N_6933);
or U7353 (N_7353,N_7020,N_6989);
xor U7354 (N_7354,N_7154,N_6931);
xnor U7355 (N_7355,N_6976,N_6934);
or U7356 (N_7356,N_7164,N_7053);
or U7357 (N_7357,N_7087,N_7180);
nor U7358 (N_7358,N_7094,N_7195);
nand U7359 (N_7359,N_6938,N_7118);
nor U7360 (N_7360,N_7107,N_7094);
or U7361 (N_7361,N_7003,N_7125);
nor U7362 (N_7362,N_7032,N_6979);
nand U7363 (N_7363,N_6915,N_7001);
or U7364 (N_7364,N_6956,N_6963);
and U7365 (N_7365,N_7041,N_6981);
nand U7366 (N_7366,N_6930,N_6932);
and U7367 (N_7367,N_7062,N_6905);
or U7368 (N_7368,N_7142,N_7120);
and U7369 (N_7369,N_6965,N_6928);
nand U7370 (N_7370,N_7060,N_6989);
nor U7371 (N_7371,N_7019,N_7076);
and U7372 (N_7372,N_7030,N_6951);
nand U7373 (N_7373,N_7055,N_6917);
nor U7374 (N_7374,N_6982,N_7186);
nor U7375 (N_7375,N_7148,N_6933);
nor U7376 (N_7376,N_6972,N_6994);
nor U7377 (N_7377,N_6940,N_6924);
xnor U7378 (N_7378,N_6941,N_7072);
nor U7379 (N_7379,N_6910,N_7191);
nor U7380 (N_7380,N_7183,N_6952);
nand U7381 (N_7381,N_6955,N_6988);
and U7382 (N_7382,N_7139,N_6983);
nor U7383 (N_7383,N_6919,N_7005);
xnor U7384 (N_7384,N_7110,N_7002);
and U7385 (N_7385,N_6932,N_6902);
xor U7386 (N_7386,N_7039,N_6935);
xor U7387 (N_7387,N_7185,N_6944);
and U7388 (N_7388,N_7043,N_6981);
and U7389 (N_7389,N_7189,N_6913);
nand U7390 (N_7390,N_7149,N_6924);
xnor U7391 (N_7391,N_7003,N_7197);
or U7392 (N_7392,N_7133,N_6982);
nor U7393 (N_7393,N_7157,N_6984);
nor U7394 (N_7394,N_7039,N_6990);
nor U7395 (N_7395,N_7068,N_7031);
xnor U7396 (N_7396,N_7189,N_7012);
or U7397 (N_7397,N_7132,N_7039);
and U7398 (N_7398,N_7132,N_7168);
and U7399 (N_7399,N_7040,N_7043);
nor U7400 (N_7400,N_7173,N_6994);
or U7401 (N_7401,N_6901,N_7094);
or U7402 (N_7402,N_7192,N_7022);
xnor U7403 (N_7403,N_7004,N_7060);
nor U7404 (N_7404,N_6998,N_6995);
xnor U7405 (N_7405,N_6955,N_7166);
nand U7406 (N_7406,N_7058,N_6969);
or U7407 (N_7407,N_7136,N_6937);
and U7408 (N_7408,N_6948,N_7017);
and U7409 (N_7409,N_7146,N_6961);
nand U7410 (N_7410,N_7021,N_6943);
xnor U7411 (N_7411,N_6964,N_6952);
or U7412 (N_7412,N_6918,N_6966);
nand U7413 (N_7413,N_6926,N_6978);
or U7414 (N_7414,N_7096,N_7136);
xnor U7415 (N_7415,N_6952,N_7084);
xor U7416 (N_7416,N_6904,N_7103);
or U7417 (N_7417,N_7002,N_7115);
or U7418 (N_7418,N_6918,N_6947);
or U7419 (N_7419,N_7057,N_7026);
or U7420 (N_7420,N_6937,N_6985);
and U7421 (N_7421,N_6917,N_7135);
nand U7422 (N_7422,N_7017,N_7115);
nor U7423 (N_7423,N_6988,N_7164);
nor U7424 (N_7424,N_7090,N_7080);
xor U7425 (N_7425,N_6991,N_7044);
or U7426 (N_7426,N_7090,N_7176);
nand U7427 (N_7427,N_6967,N_7064);
and U7428 (N_7428,N_7015,N_7005);
nand U7429 (N_7429,N_7142,N_6961);
nor U7430 (N_7430,N_7083,N_7135);
nor U7431 (N_7431,N_7055,N_6983);
nand U7432 (N_7432,N_6995,N_7163);
nand U7433 (N_7433,N_6998,N_7110);
nor U7434 (N_7434,N_7157,N_6964);
xnor U7435 (N_7435,N_7149,N_7012);
or U7436 (N_7436,N_6927,N_7086);
xnor U7437 (N_7437,N_6949,N_7124);
xor U7438 (N_7438,N_6981,N_7144);
and U7439 (N_7439,N_7103,N_7030);
xor U7440 (N_7440,N_7017,N_7111);
or U7441 (N_7441,N_7108,N_6931);
or U7442 (N_7442,N_7122,N_7140);
and U7443 (N_7443,N_7067,N_7014);
nor U7444 (N_7444,N_7167,N_7034);
or U7445 (N_7445,N_7020,N_6958);
nor U7446 (N_7446,N_6965,N_7090);
and U7447 (N_7447,N_6956,N_6998);
xnor U7448 (N_7448,N_7078,N_7045);
nor U7449 (N_7449,N_6913,N_7029);
or U7450 (N_7450,N_6965,N_7080);
nor U7451 (N_7451,N_6983,N_7192);
and U7452 (N_7452,N_6919,N_6920);
or U7453 (N_7453,N_7029,N_7155);
xnor U7454 (N_7454,N_6935,N_7002);
and U7455 (N_7455,N_6945,N_7114);
xnor U7456 (N_7456,N_7154,N_7054);
and U7457 (N_7457,N_7146,N_7026);
nand U7458 (N_7458,N_6994,N_6984);
or U7459 (N_7459,N_6918,N_7004);
nor U7460 (N_7460,N_6964,N_7172);
xor U7461 (N_7461,N_7009,N_7149);
or U7462 (N_7462,N_6960,N_7044);
xnor U7463 (N_7463,N_7145,N_7122);
nand U7464 (N_7464,N_6903,N_7098);
nor U7465 (N_7465,N_6998,N_7086);
nand U7466 (N_7466,N_6902,N_7102);
xor U7467 (N_7467,N_7117,N_6976);
nor U7468 (N_7468,N_6993,N_7083);
and U7469 (N_7469,N_7111,N_7022);
nand U7470 (N_7470,N_7120,N_7070);
and U7471 (N_7471,N_7065,N_7121);
nand U7472 (N_7472,N_7068,N_7077);
nor U7473 (N_7473,N_6913,N_7041);
or U7474 (N_7474,N_7142,N_7088);
and U7475 (N_7475,N_6905,N_7049);
xnor U7476 (N_7476,N_6925,N_7043);
nor U7477 (N_7477,N_6988,N_7123);
nand U7478 (N_7478,N_7002,N_6948);
xor U7479 (N_7479,N_7096,N_7012);
xor U7480 (N_7480,N_7157,N_7032);
or U7481 (N_7481,N_6978,N_6962);
nand U7482 (N_7482,N_6945,N_6905);
nor U7483 (N_7483,N_7094,N_7130);
and U7484 (N_7484,N_7018,N_7192);
nor U7485 (N_7485,N_7129,N_7123);
or U7486 (N_7486,N_7070,N_6956);
xor U7487 (N_7487,N_7192,N_7099);
nor U7488 (N_7488,N_7027,N_6923);
or U7489 (N_7489,N_7039,N_7122);
nor U7490 (N_7490,N_6963,N_7019);
nor U7491 (N_7491,N_6961,N_6972);
nand U7492 (N_7492,N_6913,N_6912);
nor U7493 (N_7493,N_6923,N_7053);
nor U7494 (N_7494,N_6946,N_7056);
or U7495 (N_7495,N_6918,N_6932);
or U7496 (N_7496,N_7086,N_7119);
and U7497 (N_7497,N_6972,N_7187);
or U7498 (N_7498,N_6987,N_7109);
nand U7499 (N_7499,N_7031,N_7136);
and U7500 (N_7500,N_7443,N_7334);
nand U7501 (N_7501,N_7260,N_7491);
or U7502 (N_7502,N_7423,N_7418);
xor U7503 (N_7503,N_7247,N_7290);
xnor U7504 (N_7504,N_7495,N_7279);
nand U7505 (N_7505,N_7313,N_7322);
and U7506 (N_7506,N_7365,N_7340);
and U7507 (N_7507,N_7343,N_7346);
and U7508 (N_7508,N_7381,N_7351);
and U7509 (N_7509,N_7405,N_7296);
and U7510 (N_7510,N_7314,N_7325);
xnor U7511 (N_7511,N_7398,N_7306);
nand U7512 (N_7512,N_7295,N_7361);
nand U7513 (N_7513,N_7344,N_7387);
nor U7514 (N_7514,N_7372,N_7476);
nand U7515 (N_7515,N_7428,N_7268);
nor U7516 (N_7516,N_7465,N_7499);
nand U7517 (N_7517,N_7201,N_7480);
nor U7518 (N_7518,N_7464,N_7248);
and U7519 (N_7519,N_7458,N_7249);
xor U7520 (N_7520,N_7326,N_7388);
and U7521 (N_7521,N_7481,N_7277);
nand U7522 (N_7522,N_7218,N_7427);
and U7523 (N_7523,N_7444,N_7225);
nand U7524 (N_7524,N_7456,N_7489);
xnor U7525 (N_7525,N_7370,N_7312);
or U7526 (N_7526,N_7224,N_7377);
nor U7527 (N_7527,N_7236,N_7274);
nand U7528 (N_7528,N_7397,N_7374);
nor U7529 (N_7529,N_7259,N_7229);
nor U7530 (N_7530,N_7331,N_7301);
xnor U7531 (N_7531,N_7333,N_7478);
xor U7532 (N_7532,N_7293,N_7422);
and U7533 (N_7533,N_7251,N_7366);
and U7534 (N_7534,N_7396,N_7239);
and U7535 (N_7535,N_7309,N_7291);
or U7536 (N_7536,N_7400,N_7451);
or U7537 (N_7537,N_7276,N_7206);
nand U7538 (N_7538,N_7283,N_7307);
or U7539 (N_7539,N_7359,N_7261);
and U7540 (N_7540,N_7319,N_7490);
and U7541 (N_7541,N_7357,N_7262);
or U7542 (N_7542,N_7273,N_7350);
nor U7543 (N_7543,N_7373,N_7415);
and U7544 (N_7544,N_7399,N_7233);
and U7545 (N_7545,N_7482,N_7231);
or U7546 (N_7546,N_7226,N_7311);
nand U7547 (N_7547,N_7452,N_7498);
xor U7548 (N_7548,N_7385,N_7448);
nand U7549 (N_7549,N_7235,N_7256);
nor U7550 (N_7550,N_7342,N_7230);
xor U7551 (N_7551,N_7460,N_7441);
and U7552 (N_7552,N_7287,N_7485);
nand U7553 (N_7553,N_7300,N_7475);
nor U7554 (N_7554,N_7329,N_7434);
and U7555 (N_7555,N_7375,N_7281);
nand U7556 (N_7556,N_7403,N_7417);
nand U7557 (N_7557,N_7432,N_7217);
xnor U7558 (N_7558,N_7227,N_7416);
nor U7559 (N_7559,N_7446,N_7292);
xor U7560 (N_7560,N_7459,N_7462);
or U7561 (N_7561,N_7393,N_7404);
and U7562 (N_7562,N_7243,N_7320);
nor U7563 (N_7563,N_7264,N_7376);
nand U7564 (N_7564,N_7339,N_7254);
and U7565 (N_7565,N_7488,N_7278);
nor U7566 (N_7566,N_7210,N_7440);
nand U7567 (N_7567,N_7355,N_7285);
nand U7568 (N_7568,N_7271,N_7461);
nor U7569 (N_7569,N_7242,N_7246);
xnor U7570 (N_7570,N_7299,N_7380);
and U7571 (N_7571,N_7297,N_7431);
xnor U7572 (N_7572,N_7335,N_7282);
nor U7573 (N_7573,N_7445,N_7321);
xor U7574 (N_7574,N_7202,N_7353);
or U7575 (N_7575,N_7252,N_7436);
or U7576 (N_7576,N_7263,N_7369);
nor U7577 (N_7577,N_7303,N_7241);
nand U7578 (N_7578,N_7487,N_7472);
nand U7579 (N_7579,N_7269,N_7215);
nor U7580 (N_7580,N_7338,N_7430);
nand U7581 (N_7581,N_7479,N_7395);
xor U7582 (N_7582,N_7337,N_7341);
or U7583 (N_7583,N_7204,N_7409);
or U7584 (N_7584,N_7267,N_7429);
and U7585 (N_7585,N_7474,N_7200);
and U7586 (N_7586,N_7356,N_7466);
xor U7587 (N_7587,N_7253,N_7494);
and U7588 (N_7588,N_7435,N_7392);
and U7589 (N_7589,N_7412,N_7463);
or U7590 (N_7590,N_7424,N_7315);
and U7591 (N_7591,N_7228,N_7327);
nand U7592 (N_7592,N_7382,N_7330);
xnor U7593 (N_7593,N_7238,N_7232);
nand U7594 (N_7594,N_7305,N_7216);
nand U7595 (N_7595,N_7389,N_7410);
or U7596 (N_7596,N_7371,N_7349);
xor U7597 (N_7597,N_7209,N_7394);
xnor U7598 (N_7598,N_7368,N_7250);
nand U7599 (N_7599,N_7265,N_7237);
xnor U7600 (N_7600,N_7390,N_7450);
or U7601 (N_7601,N_7294,N_7310);
nor U7602 (N_7602,N_7421,N_7288);
nor U7603 (N_7603,N_7266,N_7214);
nor U7604 (N_7604,N_7477,N_7280);
nand U7605 (N_7605,N_7298,N_7496);
and U7606 (N_7606,N_7419,N_7208);
nand U7607 (N_7607,N_7244,N_7408);
xnor U7608 (N_7608,N_7347,N_7470);
nand U7609 (N_7609,N_7220,N_7272);
xnor U7610 (N_7610,N_7289,N_7401);
xor U7611 (N_7611,N_7258,N_7453);
and U7612 (N_7612,N_7437,N_7454);
nor U7613 (N_7613,N_7402,N_7467);
or U7614 (N_7614,N_7492,N_7364);
or U7615 (N_7615,N_7336,N_7447);
nand U7616 (N_7616,N_7317,N_7486);
or U7617 (N_7617,N_7442,N_7348);
nand U7618 (N_7618,N_7302,N_7379);
and U7619 (N_7619,N_7345,N_7358);
or U7620 (N_7620,N_7406,N_7221);
or U7621 (N_7621,N_7203,N_7449);
or U7622 (N_7622,N_7386,N_7328);
xor U7623 (N_7623,N_7425,N_7275);
or U7624 (N_7624,N_7219,N_7438);
xnor U7625 (N_7625,N_7211,N_7457);
nor U7626 (N_7626,N_7484,N_7363);
and U7627 (N_7627,N_7270,N_7362);
xnor U7628 (N_7628,N_7414,N_7426);
nor U7629 (N_7629,N_7471,N_7316);
or U7630 (N_7630,N_7255,N_7407);
nor U7631 (N_7631,N_7439,N_7497);
or U7632 (N_7632,N_7493,N_7383);
nand U7633 (N_7633,N_7205,N_7360);
nor U7634 (N_7634,N_7308,N_7222);
or U7635 (N_7635,N_7286,N_7473);
and U7636 (N_7636,N_7391,N_7433);
and U7637 (N_7637,N_7420,N_7413);
and U7638 (N_7638,N_7332,N_7234);
nor U7639 (N_7639,N_7367,N_7455);
nand U7640 (N_7640,N_7318,N_7223);
nand U7641 (N_7641,N_7245,N_7378);
nor U7642 (N_7642,N_7411,N_7469);
and U7643 (N_7643,N_7213,N_7384);
nor U7644 (N_7644,N_7323,N_7304);
xor U7645 (N_7645,N_7483,N_7240);
and U7646 (N_7646,N_7257,N_7284);
and U7647 (N_7647,N_7324,N_7354);
and U7648 (N_7648,N_7212,N_7352);
and U7649 (N_7649,N_7207,N_7468);
nor U7650 (N_7650,N_7223,N_7382);
xor U7651 (N_7651,N_7349,N_7481);
and U7652 (N_7652,N_7320,N_7446);
nor U7653 (N_7653,N_7414,N_7361);
or U7654 (N_7654,N_7221,N_7456);
nand U7655 (N_7655,N_7336,N_7489);
xor U7656 (N_7656,N_7253,N_7374);
and U7657 (N_7657,N_7216,N_7235);
or U7658 (N_7658,N_7443,N_7473);
nand U7659 (N_7659,N_7245,N_7397);
xor U7660 (N_7660,N_7458,N_7334);
and U7661 (N_7661,N_7242,N_7218);
xnor U7662 (N_7662,N_7443,N_7361);
and U7663 (N_7663,N_7213,N_7366);
or U7664 (N_7664,N_7424,N_7346);
nand U7665 (N_7665,N_7499,N_7266);
xor U7666 (N_7666,N_7231,N_7444);
nor U7667 (N_7667,N_7220,N_7293);
and U7668 (N_7668,N_7492,N_7282);
xnor U7669 (N_7669,N_7453,N_7309);
nor U7670 (N_7670,N_7219,N_7334);
nor U7671 (N_7671,N_7486,N_7219);
xnor U7672 (N_7672,N_7434,N_7216);
or U7673 (N_7673,N_7206,N_7340);
nor U7674 (N_7674,N_7267,N_7453);
and U7675 (N_7675,N_7330,N_7229);
xnor U7676 (N_7676,N_7340,N_7274);
nand U7677 (N_7677,N_7263,N_7403);
nor U7678 (N_7678,N_7453,N_7248);
or U7679 (N_7679,N_7469,N_7218);
xor U7680 (N_7680,N_7343,N_7270);
or U7681 (N_7681,N_7247,N_7315);
or U7682 (N_7682,N_7372,N_7302);
nand U7683 (N_7683,N_7331,N_7485);
nand U7684 (N_7684,N_7441,N_7449);
nor U7685 (N_7685,N_7402,N_7310);
or U7686 (N_7686,N_7203,N_7348);
nand U7687 (N_7687,N_7222,N_7204);
and U7688 (N_7688,N_7365,N_7218);
and U7689 (N_7689,N_7411,N_7286);
or U7690 (N_7690,N_7289,N_7426);
nor U7691 (N_7691,N_7439,N_7264);
nand U7692 (N_7692,N_7232,N_7292);
xnor U7693 (N_7693,N_7483,N_7418);
nand U7694 (N_7694,N_7333,N_7350);
nor U7695 (N_7695,N_7265,N_7348);
nand U7696 (N_7696,N_7421,N_7488);
and U7697 (N_7697,N_7402,N_7373);
xor U7698 (N_7698,N_7384,N_7239);
nor U7699 (N_7699,N_7398,N_7360);
or U7700 (N_7700,N_7497,N_7426);
or U7701 (N_7701,N_7277,N_7419);
nand U7702 (N_7702,N_7329,N_7441);
xnor U7703 (N_7703,N_7432,N_7313);
or U7704 (N_7704,N_7211,N_7317);
nor U7705 (N_7705,N_7237,N_7343);
and U7706 (N_7706,N_7361,N_7353);
or U7707 (N_7707,N_7275,N_7236);
nor U7708 (N_7708,N_7391,N_7384);
xor U7709 (N_7709,N_7495,N_7441);
and U7710 (N_7710,N_7282,N_7435);
xor U7711 (N_7711,N_7236,N_7367);
nand U7712 (N_7712,N_7414,N_7373);
nor U7713 (N_7713,N_7454,N_7364);
nand U7714 (N_7714,N_7489,N_7338);
nor U7715 (N_7715,N_7341,N_7338);
and U7716 (N_7716,N_7362,N_7456);
nor U7717 (N_7717,N_7360,N_7275);
and U7718 (N_7718,N_7452,N_7345);
nor U7719 (N_7719,N_7318,N_7402);
and U7720 (N_7720,N_7380,N_7314);
or U7721 (N_7721,N_7235,N_7325);
xor U7722 (N_7722,N_7330,N_7293);
xor U7723 (N_7723,N_7408,N_7252);
nand U7724 (N_7724,N_7213,N_7226);
nand U7725 (N_7725,N_7473,N_7313);
xor U7726 (N_7726,N_7466,N_7440);
nand U7727 (N_7727,N_7343,N_7282);
nor U7728 (N_7728,N_7368,N_7265);
and U7729 (N_7729,N_7468,N_7295);
nor U7730 (N_7730,N_7457,N_7494);
or U7731 (N_7731,N_7336,N_7235);
or U7732 (N_7732,N_7311,N_7442);
nor U7733 (N_7733,N_7495,N_7494);
or U7734 (N_7734,N_7304,N_7344);
and U7735 (N_7735,N_7411,N_7201);
xor U7736 (N_7736,N_7257,N_7475);
nand U7737 (N_7737,N_7285,N_7238);
nand U7738 (N_7738,N_7352,N_7209);
or U7739 (N_7739,N_7356,N_7387);
nand U7740 (N_7740,N_7453,N_7314);
xor U7741 (N_7741,N_7237,N_7318);
nand U7742 (N_7742,N_7319,N_7392);
xnor U7743 (N_7743,N_7444,N_7213);
or U7744 (N_7744,N_7428,N_7352);
nand U7745 (N_7745,N_7266,N_7457);
nand U7746 (N_7746,N_7422,N_7429);
or U7747 (N_7747,N_7240,N_7360);
xnor U7748 (N_7748,N_7347,N_7242);
xor U7749 (N_7749,N_7447,N_7302);
or U7750 (N_7750,N_7392,N_7477);
xor U7751 (N_7751,N_7463,N_7388);
xnor U7752 (N_7752,N_7444,N_7363);
or U7753 (N_7753,N_7309,N_7460);
nand U7754 (N_7754,N_7235,N_7419);
nor U7755 (N_7755,N_7279,N_7307);
or U7756 (N_7756,N_7329,N_7249);
nand U7757 (N_7757,N_7463,N_7461);
nor U7758 (N_7758,N_7380,N_7205);
nand U7759 (N_7759,N_7343,N_7301);
nand U7760 (N_7760,N_7434,N_7435);
or U7761 (N_7761,N_7475,N_7386);
or U7762 (N_7762,N_7470,N_7329);
nand U7763 (N_7763,N_7210,N_7467);
nor U7764 (N_7764,N_7458,N_7255);
nor U7765 (N_7765,N_7351,N_7294);
and U7766 (N_7766,N_7282,N_7270);
or U7767 (N_7767,N_7354,N_7428);
nor U7768 (N_7768,N_7395,N_7309);
or U7769 (N_7769,N_7243,N_7208);
and U7770 (N_7770,N_7394,N_7349);
or U7771 (N_7771,N_7274,N_7484);
nor U7772 (N_7772,N_7238,N_7454);
nand U7773 (N_7773,N_7344,N_7484);
and U7774 (N_7774,N_7415,N_7214);
nand U7775 (N_7775,N_7403,N_7419);
nor U7776 (N_7776,N_7303,N_7235);
xnor U7777 (N_7777,N_7421,N_7436);
nor U7778 (N_7778,N_7313,N_7297);
nand U7779 (N_7779,N_7480,N_7345);
xor U7780 (N_7780,N_7271,N_7409);
xnor U7781 (N_7781,N_7475,N_7246);
xor U7782 (N_7782,N_7284,N_7248);
xor U7783 (N_7783,N_7408,N_7350);
nand U7784 (N_7784,N_7284,N_7373);
nand U7785 (N_7785,N_7333,N_7380);
and U7786 (N_7786,N_7476,N_7473);
or U7787 (N_7787,N_7363,N_7204);
xnor U7788 (N_7788,N_7366,N_7216);
or U7789 (N_7789,N_7264,N_7308);
nand U7790 (N_7790,N_7457,N_7267);
and U7791 (N_7791,N_7312,N_7226);
xor U7792 (N_7792,N_7217,N_7276);
xor U7793 (N_7793,N_7384,N_7335);
nor U7794 (N_7794,N_7216,N_7308);
nor U7795 (N_7795,N_7428,N_7418);
xnor U7796 (N_7796,N_7302,N_7351);
or U7797 (N_7797,N_7422,N_7407);
nor U7798 (N_7798,N_7427,N_7343);
xnor U7799 (N_7799,N_7224,N_7247);
xnor U7800 (N_7800,N_7749,N_7655);
nor U7801 (N_7801,N_7608,N_7777);
nor U7802 (N_7802,N_7609,N_7747);
or U7803 (N_7803,N_7526,N_7599);
nor U7804 (N_7804,N_7778,N_7576);
and U7805 (N_7805,N_7657,N_7536);
nor U7806 (N_7806,N_7764,N_7742);
nand U7807 (N_7807,N_7773,N_7504);
and U7808 (N_7808,N_7568,N_7787);
xnor U7809 (N_7809,N_7701,N_7666);
nor U7810 (N_7810,N_7769,N_7685);
and U7811 (N_7811,N_7614,N_7798);
nand U7812 (N_7812,N_7616,N_7706);
or U7813 (N_7813,N_7687,N_7751);
nor U7814 (N_7814,N_7535,N_7733);
nand U7815 (N_7815,N_7668,N_7513);
or U7816 (N_7816,N_7652,N_7712);
or U7817 (N_7817,N_7705,N_7528);
nor U7818 (N_7818,N_7692,N_7761);
and U7819 (N_7819,N_7691,N_7781);
xnor U7820 (N_7820,N_7543,N_7713);
nand U7821 (N_7821,N_7647,N_7618);
and U7822 (N_7822,N_7678,N_7532);
xnor U7823 (N_7823,N_7745,N_7520);
xor U7824 (N_7824,N_7631,N_7728);
xnor U7825 (N_7825,N_7621,N_7667);
xnor U7826 (N_7826,N_7675,N_7771);
nand U7827 (N_7827,N_7661,N_7559);
nand U7828 (N_7828,N_7753,N_7649);
nor U7829 (N_7829,N_7715,N_7774);
nand U7830 (N_7830,N_7736,N_7522);
xnor U7831 (N_7831,N_7629,N_7596);
nand U7832 (N_7832,N_7780,N_7542);
nor U7833 (N_7833,N_7799,N_7592);
or U7834 (N_7834,N_7517,N_7540);
nor U7835 (N_7835,N_7703,N_7502);
nor U7836 (N_7836,N_7597,N_7775);
nor U7837 (N_7837,N_7622,N_7562);
nand U7838 (N_7838,N_7791,N_7602);
nand U7839 (N_7839,N_7730,N_7610);
xor U7840 (N_7840,N_7611,N_7653);
and U7841 (N_7841,N_7690,N_7527);
or U7842 (N_7842,N_7548,N_7590);
and U7843 (N_7843,N_7663,N_7697);
xnor U7844 (N_7844,N_7577,N_7752);
and U7845 (N_7845,N_7630,N_7595);
nor U7846 (N_7846,N_7534,N_7579);
and U7847 (N_7847,N_7735,N_7759);
nor U7848 (N_7848,N_7533,N_7546);
nand U7849 (N_7849,N_7555,N_7686);
nor U7850 (N_7850,N_7672,N_7662);
and U7851 (N_7851,N_7605,N_7665);
xnor U7852 (N_7852,N_7537,N_7669);
xor U7853 (N_7853,N_7566,N_7628);
xnor U7854 (N_7854,N_7714,N_7716);
and U7855 (N_7855,N_7793,N_7746);
xor U7856 (N_7856,N_7623,N_7788);
nand U7857 (N_7857,N_7547,N_7737);
xor U7858 (N_7858,N_7738,N_7565);
nor U7859 (N_7859,N_7754,N_7569);
xor U7860 (N_7860,N_7766,N_7510);
nand U7861 (N_7861,N_7606,N_7689);
nand U7862 (N_7862,N_7765,N_7589);
or U7863 (N_7863,N_7585,N_7594);
xnor U7864 (N_7864,N_7664,N_7556);
xor U7865 (N_7865,N_7636,N_7500);
or U7866 (N_7866,N_7524,N_7554);
nand U7867 (N_7867,N_7545,N_7726);
nand U7868 (N_7868,N_7511,N_7587);
and U7869 (N_7869,N_7583,N_7708);
or U7870 (N_7870,N_7743,N_7683);
nand U7871 (N_7871,N_7702,N_7581);
and U7872 (N_7872,N_7523,N_7563);
nand U7873 (N_7873,N_7682,N_7707);
or U7874 (N_7874,N_7684,N_7725);
xor U7875 (N_7875,N_7603,N_7709);
or U7876 (N_7876,N_7501,N_7792);
nand U7877 (N_7877,N_7627,N_7696);
xnor U7878 (N_7878,N_7763,N_7558);
or U7879 (N_7879,N_7541,N_7643);
xnor U7880 (N_7880,N_7508,N_7518);
xnor U7881 (N_7881,N_7758,N_7586);
or U7882 (N_7882,N_7637,N_7561);
xnor U7883 (N_7883,N_7695,N_7784);
or U7884 (N_7884,N_7525,N_7711);
xnor U7885 (N_7885,N_7721,N_7794);
or U7886 (N_7886,N_7538,N_7507);
nand U7887 (N_7887,N_7646,N_7676);
nand U7888 (N_7888,N_7724,N_7617);
and U7889 (N_7889,N_7505,N_7607);
and U7890 (N_7890,N_7723,N_7734);
and U7891 (N_7891,N_7674,N_7748);
or U7892 (N_7892,N_7509,N_7620);
or U7893 (N_7893,N_7519,N_7544);
xor U7894 (N_7894,N_7710,N_7694);
nor U7895 (N_7895,N_7762,N_7521);
xnor U7896 (N_7896,N_7591,N_7550);
nor U7897 (N_7897,N_7626,N_7633);
nor U7898 (N_7898,N_7670,N_7727);
or U7899 (N_7899,N_7514,N_7580);
nand U7900 (N_7900,N_7744,N_7634);
xor U7901 (N_7901,N_7729,N_7575);
nand U7902 (N_7902,N_7601,N_7718);
nor U7903 (N_7903,N_7755,N_7739);
xor U7904 (N_7904,N_7767,N_7776);
nand U7905 (N_7905,N_7688,N_7516);
or U7906 (N_7906,N_7573,N_7677);
or U7907 (N_7907,N_7756,N_7604);
nand U7908 (N_7908,N_7635,N_7785);
xnor U7909 (N_7909,N_7770,N_7564);
nor U7910 (N_7910,N_7772,N_7717);
nand U7911 (N_7911,N_7741,N_7557);
nand U7912 (N_7912,N_7660,N_7644);
nand U7913 (N_7913,N_7584,N_7615);
xor U7914 (N_7914,N_7640,N_7624);
xnor U7915 (N_7915,N_7567,N_7704);
nor U7916 (N_7916,N_7673,N_7651);
nor U7917 (N_7917,N_7760,N_7570);
and U7918 (N_7918,N_7699,N_7797);
xor U7919 (N_7919,N_7529,N_7553);
nor U7920 (N_7920,N_7531,N_7588);
nand U7921 (N_7921,N_7698,N_7732);
xnor U7922 (N_7922,N_7572,N_7790);
or U7923 (N_7923,N_7530,N_7549);
or U7924 (N_7924,N_7795,N_7593);
nand U7925 (N_7925,N_7740,N_7693);
xnor U7926 (N_7926,N_7720,N_7632);
or U7927 (N_7927,N_7552,N_7700);
xor U7928 (N_7928,N_7782,N_7551);
xor U7929 (N_7929,N_7783,N_7796);
and U7930 (N_7930,N_7679,N_7654);
or U7931 (N_7931,N_7578,N_7731);
xnor U7932 (N_7932,N_7650,N_7722);
nand U7933 (N_7933,N_7625,N_7515);
or U7934 (N_7934,N_7571,N_7681);
nand U7935 (N_7935,N_7658,N_7612);
nor U7936 (N_7936,N_7750,N_7757);
or U7937 (N_7937,N_7506,N_7648);
xor U7938 (N_7938,N_7598,N_7560);
nand U7939 (N_7939,N_7642,N_7786);
xnor U7940 (N_7940,N_7613,N_7680);
or U7941 (N_7941,N_7574,N_7503);
or U7942 (N_7942,N_7638,N_7656);
or U7943 (N_7943,N_7619,N_7768);
or U7944 (N_7944,N_7539,N_7671);
or U7945 (N_7945,N_7641,N_7645);
nand U7946 (N_7946,N_7779,N_7789);
nand U7947 (N_7947,N_7639,N_7512);
xnor U7948 (N_7948,N_7600,N_7659);
xnor U7949 (N_7949,N_7582,N_7719);
or U7950 (N_7950,N_7728,N_7618);
xnor U7951 (N_7951,N_7521,N_7587);
nor U7952 (N_7952,N_7553,N_7662);
xor U7953 (N_7953,N_7707,N_7747);
and U7954 (N_7954,N_7659,N_7528);
nand U7955 (N_7955,N_7662,N_7548);
nand U7956 (N_7956,N_7530,N_7726);
xnor U7957 (N_7957,N_7656,N_7511);
nor U7958 (N_7958,N_7713,N_7591);
or U7959 (N_7959,N_7576,N_7640);
nor U7960 (N_7960,N_7660,N_7511);
and U7961 (N_7961,N_7533,N_7793);
xnor U7962 (N_7962,N_7709,N_7563);
or U7963 (N_7963,N_7797,N_7777);
and U7964 (N_7964,N_7645,N_7699);
nor U7965 (N_7965,N_7767,N_7651);
or U7966 (N_7966,N_7599,N_7696);
nor U7967 (N_7967,N_7500,N_7607);
nor U7968 (N_7968,N_7609,N_7799);
nand U7969 (N_7969,N_7531,N_7506);
or U7970 (N_7970,N_7543,N_7511);
and U7971 (N_7971,N_7757,N_7701);
nand U7972 (N_7972,N_7672,N_7683);
and U7973 (N_7973,N_7757,N_7793);
or U7974 (N_7974,N_7651,N_7721);
xnor U7975 (N_7975,N_7603,N_7758);
or U7976 (N_7976,N_7735,N_7649);
or U7977 (N_7977,N_7625,N_7616);
nor U7978 (N_7978,N_7696,N_7690);
nor U7979 (N_7979,N_7603,N_7501);
or U7980 (N_7980,N_7521,N_7665);
xor U7981 (N_7981,N_7628,N_7575);
or U7982 (N_7982,N_7560,N_7625);
nand U7983 (N_7983,N_7757,N_7592);
xor U7984 (N_7984,N_7547,N_7677);
or U7985 (N_7985,N_7712,N_7523);
nand U7986 (N_7986,N_7663,N_7538);
xnor U7987 (N_7987,N_7791,N_7740);
or U7988 (N_7988,N_7575,N_7603);
nor U7989 (N_7989,N_7749,N_7607);
and U7990 (N_7990,N_7544,N_7644);
nor U7991 (N_7991,N_7655,N_7584);
and U7992 (N_7992,N_7743,N_7563);
and U7993 (N_7993,N_7683,N_7778);
and U7994 (N_7994,N_7781,N_7789);
or U7995 (N_7995,N_7758,N_7505);
and U7996 (N_7996,N_7728,N_7779);
or U7997 (N_7997,N_7547,N_7691);
xnor U7998 (N_7998,N_7546,N_7624);
or U7999 (N_7999,N_7774,N_7782);
nor U8000 (N_8000,N_7734,N_7598);
nand U8001 (N_8001,N_7699,N_7554);
and U8002 (N_8002,N_7585,N_7534);
nand U8003 (N_8003,N_7634,N_7741);
nand U8004 (N_8004,N_7668,N_7599);
nor U8005 (N_8005,N_7681,N_7738);
xnor U8006 (N_8006,N_7571,N_7502);
xnor U8007 (N_8007,N_7778,N_7740);
xor U8008 (N_8008,N_7721,N_7748);
nor U8009 (N_8009,N_7653,N_7601);
nor U8010 (N_8010,N_7603,N_7534);
xor U8011 (N_8011,N_7755,N_7551);
or U8012 (N_8012,N_7588,N_7698);
and U8013 (N_8013,N_7792,N_7742);
or U8014 (N_8014,N_7642,N_7591);
and U8015 (N_8015,N_7660,N_7713);
nand U8016 (N_8016,N_7698,N_7584);
and U8017 (N_8017,N_7762,N_7754);
xnor U8018 (N_8018,N_7503,N_7742);
xnor U8019 (N_8019,N_7554,N_7526);
nand U8020 (N_8020,N_7784,N_7697);
nand U8021 (N_8021,N_7598,N_7771);
and U8022 (N_8022,N_7790,N_7686);
xnor U8023 (N_8023,N_7572,N_7686);
nor U8024 (N_8024,N_7677,N_7623);
nor U8025 (N_8025,N_7581,N_7734);
nand U8026 (N_8026,N_7682,N_7555);
xor U8027 (N_8027,N_7511,N_7776);
or U8028 (N_8028,N_7535,N_7676);
nand U8029 (N_8029,N_7672,N_7593);
xnor U8030 (N_8030,N_7794,N_7715);
and U8031 (N_8031,N_7593,N_7586);
nor U8032 (N_8032,N_7587,N_7633);
xor U8033 (N_8033,N_7614,N_7776);
and U8034 (N_8034,N_7748,N_7513);
and U8035 (N_8035,N_7649,N_7575);
and U8036 (N_8036,N_7697,N_7689);
xnor U8037 (N_8037,N_7689,N_7506);
and U8038 (N_8038,N_7564,N_7519);
xor U8039 (N_8039,N_7581,N_7546);
and U8040 (N_8040,N_7707,N_7670);
or U8041 (N_8041,N_7625,N_7672);
nand U8042 (N_8042,N_7548,N_7591);
and U8043 (N_8043,N_7578,N_7518);
or U8044 (N_8044,N_7649,N_7541);
nor U8045 (N_8045,N_7695,N_7638);
nand U8046 (N_8046,N_7706,N_7696);
nor U8047 (N_8047,N_7519,N_7518);
nor U8048 (N_8048,N_7774,N_7795);
and U8049 (N_8049,N_7511,N_7748);
and U8050 (N_8050,N_7581,N_7502);
and U8051 (N_8051,N_7710,N_7706);
and U8052 (N_8052,N_7744,N_7706);
nor U8053 (N_8053,N_7778,N_7533);
or U8054 (N_8054,N_7585,N_7573);
or U8055 (N_8055,N_7532,N_7727);
and U8056 (N_8056,N_7691,N_7579);
nor U8057 (N_8057,N_7638,N_7798);
nor U8058 (N_8058,N_7759,N_7751);
nor U8059 (N_8059,N_7773,N_7593);
nor U8060 (N_8060,N_7773,N_7723);
xnor U8061 (N_8061,N_7770,N_7659);
or U8062 (N_8062,N_7614,N_7568);
nor U8063 (N_8063,N_7559,N_7535);
and U8064 (N_8064,N_7543,N_7503);
nand U8065 (N_8065,N_7700,N_7563);
xnor U8066 (N_8066,N_7750,N_7570);
or U8067 (N_8067,N_7632,N_7699);
xnor U8068 (N_8068,N_7573,N_7736);
or U8069 (N_8069,N_7716,N_7632);
nand U8070 (N_8070,N_7708,N_7518);
nor U8071 (N_8071,N_7672,N_7646);
nand U8072 (N_8072,N_7794,N_7618);
and U8073 (N_8073,N_7567,N_7597);
or U8074 (N_8074,N_7650,N_7707);
xnor U8075 (N_8075,N_7644,N_7540);
nor U8076 (N_8076,N_7642,N_7549);
nand U8077 (N_8077,N_7778,N_7516);
xor U8078 (N_8078,N_7681,N_7650);
nor U8079 (N_8079,N_7705,N_7778);
xnor U8080 (N_8080,N_7577,N_7723);
xnor U8081 (N_8081,N_7654,N_7557);
and U8082 (N_8082,N_7760,N_7739);
or U8083 (N_8083,N_7654,N_7677);
and U8084 (N_8084,N_7795,N_7675);
nand U8085 (N_8085,N_7595,N_7723);
or U8086 (N_8086,N_7616,N_7680);
nand U8087 (N_8087,N_7662,N_7655);
and U8088 (N_8088,N_7718,N_7644);
xor U8089 (N_8089,N_7692,N_7755);
nand U8090 (N_8090,N_7750,N_7602);
nor U8091 (N_8091,N_7634,N_7509);
nand U8092 (N_8092,N_7742,N_7676);
or U8093 (N_8093,N_7698,N_7675);
xor U8094 (N_8094,N_7505,N_7777);
nand U8095 (N_8095,N_7666,N_7738);
and U8096 (N_8096,N_7728,N_7733);
or U8097 (N_8097,N_7531,N_7732);
and U8098 (N_8098,N_7742,N_7644);
nor U8099 (N_8099,N_7677,N_7620);
xor U8100 (N_8100,N_7860,N_7847);
nand U8101 (N_8101,N_8022,N_7911);
nor U8102 (N_8102,N_7835,N_7937);
nor U8103 (N_8103,N_7842,N_7935);
and U8104 (N_8104,N_7976,N_8092);
nor U8105 (N_8105,N_8080,N_7925);
or U8106 (N_8106,N_7804,N_7802);
or U8107 (N_8107,N_8064,N_8077);
nor U8108 (N_8108,N_7829,N_7917);
nand U8109 (N_8109,N_7866,N_7856);
nor U8110 (N_8110,N_8025,N_7904);
xor U8111 (N_8111,N_7965,N_8086);
nand U8112 (N_8112,N_7843,N_7882);
xnor U8113 (N_8113,N_7826,N_7845);
or U8114 (N_8114,N_8062,N_7938);
nand U8115 (N_8115,N_8051,N_8040);
or U8116 (N_8116,N_7898,N_7915);
and U8117 (N_8117,N_7852,N_7810);
and U8118 (N_8118,N_8052,N_8019);
nor U8119 (N_8119,N_8050,N_7908);
nand U8120 (N_8120,N_8012,N_8097);
and U8121 (N_8121,N_7889,N_7834);
or U8122 (N_8122,N_7982,N_8038);
nand U8123 (N_8123,N_7920,N_7959);
xor U8124 (N_8124,N_7998,N_8029);
and U8125 (N_8125,N_8057,N_8046);
xnor U8126 (N_8126,N_8009,N_8008);
nor U8127 (N_8127,N_7929,N_7903);
nor U8128 (N_8128,N_7836,N_8091);
xor U8129 (N_8129,N_8079,N_8094);
nor U8130 (N_8130,N_8018,N_7864);
nand U8131 (N_8131,N_7883,N_7857);
nor U8132 (N_8132,N_7841,N_8082);
nor U8133 (N_8133,N_7913,N_7919);
or U8134 (N_8134,N_7894,N_7936);
xnor U8135 (N_8135,N_8081,N_7850);
or U8136 (N_8136,N_7906,N_7806);
or U8137 (N_8137,N_8072,N_8068);
or U8138 (N_8138,N_7941,N_7820);
or U8139 (N_8139,N_8049,N_7888);
or U8140 (N_8140,N_8039,N_8016);
or U8141 (N_8141,N_8036,N_7805);
and U8142 (N_8142,N_8048,N_7944);
xnor U8143 (N_8143,N_7816,N_8067);
nand U8144 (N_8144,N_7817,N_7876);
and U8145 (N_8145,N_7973,N_8075);
and U8146 (N_8146,N_7962,N_7961);
nand U8147 (N_8147,N_7803,N_7971);
xor U8148 (N_8148,N_7995,N_8010);
and U8149 (N_8149,N_7943,N_7951);
nand U8150 (N_8150,N_8047,N_7887);
xor U8151 (N_8151,N_7809,N_7892);
or U8152 (N_8152,N_7890,N_7838);
nand U8153 (N_8153,N_7879,N_7886);
nand U8154 (N_8154,N_8017,N_7993);
and U8155 (N_8155,N_7862,N_7932);
nand U8156 (N_8156,N_8063,N_8034);
or U8157 (N_8157,N_8028,N_7955);
xor U8158 (N_8158,N_7916,N_8053);
nand U8159 (N_8159,N_7927,N_7855);
or U8160 (N_8160,N_7827,N_7884);
nor U8161 (N_8161,N_7865,N_7873);
and U8162 (N_8162,N_7861,N_7940);
nor U8163 (N_8163,N_7914,N_7996);
and U8164 (N_8164,N_7956,N_7885);
and U8165 (N_8165,N_7905,N_8044);
or U8166 (N_8166,N_8045,N_8021);
xnor U8167 (N_8167,N_8001,N_8088);
nor U8168 (N_8168,N_7828,N_7949);
nand U8169 (N_8169,N_8070,N_7990);
xor U8170 (N_8170,N_8033,N_7831);
and U8171 (N_8171,N_7837,N_7954);
or U8172 (N_8172,N_7822,N_7896);
nor U8173 (N_8173,N_8098,N_7969);
nor U8174 (N_8174,N_7849,N_8059);
xnor U8175 (N_8175,N_8015,N_8020);
nand U8176 (N_8176,N_7840,N_7874);
xor U8177 (N_8177,N_8006,N_7891);
nor U8178 (N_8178,N_7984,N_7881);
nand U8179 (N_8179,N_8099,N_7931);
nor U8180 (N_8180,N_8037,N_8014);
nand U8181 (N_8181,N_7947,N_8089);
nor U8182 (N_8182,N_7991,N_8071);
nor U8183 (N_8183,N_8087,N_7833);
nand U8184 (N_8184,N_7946,N_7912);
or U8185 (N_8185,N_7978,N_7808);
nand U8186 (N_8186,N_7986,N_8076);
nor U8187 (N_8187,N_7968,N_7846);
xnor U8188 (N_8188,N_7981,N_7979);
xnor U8189 (N_8189,N_7985,N_7963);
nor U8190 (N_8190,N_7839,N_8002);
and U8191 (N_8191,N_7933,N_7923);
nor U8192 (N_8192,N_7950,N_7854);
and U8193 (N_8193,N_8056,N_7921);
xor U8194 (N_8194,N_8030,N_8061);
or U8195 (N_8195,N_7825,N_7859);
nand U8196 (N_8196,N_7983,N_7812);
and U8197 (N_8197,N_7989,N_7972);
nor U8198 (N_8198,N_7823,N_7928);
nand U8199 (N_8199,N_7880,N_7900);
and U8200 (N_8200,N_7964,N_8035);
and U8201 (N_8201,N_7818,N_7930);
xnor U8202 (N_8202,N_7878,N_7952);
and U8203 (N_8203,N_8027,N_7848);
or U8204 (N_8204,N_7858,N_7815);
nor U8205 (N_8205,N_7853,N_8055);
xor U8206 (N_8206,N_8058,N_8031);
and U8207 (N_8207,N_8005,N_7868);
and U8208 (N_8208,N_8096,N_7970);
nand U8209 (N_8209,N_7851,N_7801);
nand U8210 (N_8210,N_8090,N_8011);
nand U8211 (N_8211,N_7975,N_7872);
or U8212 (N_8212,N_7807,N_7902);
xnor U8213 (N_8213,N_8032,N_8000);
nand U8214 (N_8214,N_8054,N_7832);
or U8215 (N_8215,N_7988,N_7871);
xor U8216 (N_8216,N_8041,N_8095);
xnor U8217 (N_8217,N_7957,N_8024);
xor U8218 (N_8218,N_8043,N_8074);
nand U8219 (N_8219,N_7945,N_7869);
nor U8220 (N_8220,N_8069,N_7977);
and U8221 (N_8221,N_7863,N_7844);
xor U8222 (N_8222,N_7800,N_8003);
and U8223 (N_8223,N_8085,N_7918);
xor U8224 (N_8224,N_8042,N_7987);
xnor U8225 (N_8225,N_7997,N_7907);
and U8226 (N_8226,N_7958,N_7967);
nor U8227 (N_8227,N_8066,N_8073);
nand U8228 (N_8228,N_7999,N_8078);
nand U8229 (N_8229,N_7974,N_7953);
nand U8230 (N_8230,N_7870,N_8083);
xnor U8231 (N_8231,N_8013,N_7811);
and U8232 (N_8232,N_8084,N_7934);
xnor U8233 (N_8233,N_7867,N_7814);
or U8234 (N_8234,N_8060,N_7966);
xor U8235 (N_8235,N_7939,N_8026);
nor U8236 (N_8236,N_7922,N_7821);
nor U8237 (N_8237,N_8065,N_8023);
and U8238 (N_8238,N_7893,N_7819);
and U8239 (N_8239,N_7992,N_7926);
or U8240 (N_8240,N_8007,N_7875);
xnor U8241 (N_8241,N_7813,N_8004);
xor U8242 (N_8242,N_7994,N_7901);
nor U8243 (N_8243,N_7960,N_7899);
and U8244 (N_8244,N_7877,N_7830);
and U8245 (N_8245,N_7909,N_7910);
nand U8246 (N_8246,N_8093,N_7895);
nor U8247 (N_8247,N_7924,N_7897);
xnor U8248 (N_8248,N_7948,N_7942);
nand U8249 (N_8249,N_7980,N_7824);
and U8250 (N_8250,N_8088,N_7937);
nor U8251 (N_8251,N_7954,N_7919);
nor U8252 (N_8252,N_7955,N_8064);
nand U8253 (N_8253,N_7859,N_7993);
nand U8254 (N_8254,N_7930,N_8099);
or U8255 (N_8255,N_8014,N_7874);
xnor U8256 (N_8256,N_8060,N_7987);
and U8257 (N_8257,N_7913,N_7876);
xnor U8258 (N_8258,N_8058,N_7823);
or U8259 (N_8259,N_7933,N_7973);
or U8260 (N_8260,N_7815,N_7856);
and U8261 (N_8261,N_8085,N_7810);
and U8262 (N_8262,N_8073,N_7801);
xnor U8263 (N_8263,N_7985,N_8005);
and U8264 (N_8264,N_8025,N_7867);
nor U8265 (N_8265,N_7809,N_8006);
and U8266 (N_8266,N_7928,N_8052);
or U8267 (N_8267,N_8004,N_7991);
xor U8268 (N_8268,N_8064,N_7957);
nor U8269 (N_8269,N_7992,N_8010);
nand U8270 (N_8270,N_8074,N_7919);
or U8271 (N_8271,N_7800,N_7841);
and U8272 (N_8272,N_7852,N_8047);
or U8273 (N_8273,N_8066,N_7885);
xor U8274 (N_8274,N_8040,N_7942);
nor U8275 (N_8275,N_7963,N_7833);
nor U8276 (N_8276,N_7963,N_7892);
or U8277 (N_8277,N_7881,N_8065);
nor U8278 (N_8278,N_8019,N_7905);
or U8279 (N_8279,N_7964,N_8066);
or U8280 (N_8280,N_7960,N_8032);
nand U8281 (N_8281,N_7980,N_7891);
and U8282 (N_8282,N_8074,N_7900);
nand U8283 (N_8283,N_7827,N_7936);
or U8284 (N_8284,N_8046,N_7999);
xor U8285 (N_8285,N_7830,N_8087);
xor U8286 (N_8286,N_7915,N_7926);
xnor U8287 (N_8287,N_7928,N_7870);
and U8288 (N_8288,N_7922,N_7944);
nor U8289 (N_8289,N_8015,N_8009);
nand U8290 (N_8290,N_8005,N_7827);
or U8291 (N_8291,N_7905,N_8075);
nand U8292 (N_8292,N_7927,N_7918);
or U8293 (N_8293,N_7804,N_7920);
nand U8294 (N_8294,N_8048,N_8086);
nand U8295 (N_8295,N_7806,N_7952);
xnor U8296 (N_8296,N_7907,N_7987);
xnor U8297 (N_8297,N_7897,N_7944);
nand U8298 (N_8298,N_7849,N_7810);
xor U8299 (N_8299,N_7814,N_7948);
nor U8300 (N_8300,N_7940,N_7987);
or U8301 (N_8301,N_7829,N_8094);
xor U8302 (N_8302,N_7835,N_7902);
and U8303 (N_8303,N_7999,N_7813);
nor U8304 (N_8304,N_7879,N_8054);
and U8305 (N_8305,N_7991,N_8017);
or U8306 (N_8306,N_7848,N_7866);
and U8307 (N_8307,N_7803,N_7934);
or U8308 (N_8308,N_8033,N_8096);
or U8309 (N_8309,N_7889,N_7835);
nand U8310 (N_8310,N_7829,N_7953);
nor U8311 (N_8311,N_8082,N_7807);
nor U8312 (N_8312,N_7975,N_7904);
or U8313 (N_8313,N_7937,N_7906);
or U8314 (N_8314,N_7860,N_8069);
nor U8315 (N_8315,N_8026,N_8001);
nand U8316 (N_8316,N_7879,N_7848);
or U8317 (N_8317,N_7845,N_7884);
nand U8318 (N_8318,N_8068,N_7972);
nand U8319 (N_8319,N_7915,N_8083);
or U8320 (N_8320,N_8099,N_8028);
nand U8321 (N_8321,N_7809,N_7855);
xnor U8322 (N_8322,N_7911,N_8034);
and U8323 (N_8323,N_7836,N_8001);
nor U8324 (N_8324,N_8070,N_7970);
and U8325 (N_8325,N_7824,N_7992);
nand U8326 (N_8326,N_7812,N_8051);
nand U8327 (N_8327,N_8047,N_8007);
and U8328 (N_8328,N_7890,N_7947);
and U8329 (N_8329,N_7960,N_8022);
or U8330 (N_8330,N_8063,N_8043);
xnor U8331 (N_8331,N_7991,N_7856);
nor U8332 (N_8332,N_7886,N_7933);
nand U8333 (N_8333,N_7844,N_8012);
nor U8334 (N_8334,N_7933,N_7956);
and U8335 (N_8335,N_8011,N_8036);
nand U8336 (N_8336,N_8045,N_8063);
nand U8337 (N_8337,N_8034,N_7820);
xnor U8338 (N_8338,N_8058,N_8081);
xnor U8339 (N_8339,N_7830,N_8064);
and U8340 (N_8340,N_8040,N_7948);
xnor U8341 (N_8341,N_7859,N_7909);
or U8342 (N_8342,N_7800,N_8094);
nand U8343 (N_8343,N_8001,N_8062);
nor U8344 (N_8344,N_7906,N_8029);
nand U8345 (N_8345,N_7823,N_7924);
and U8346 (N_8346,N_7824,N_7967);
nor U8347 (N_8347,N_8055,N_7838);
nand U8348 (N_8348,N_7896,N_7932);
nor U8349 (N_8349,N_8028,N_7901);
or U8350 (N_8350,N_8018,N_8075);
xnor U8351 (N_8351,N_8014,N_7840);
and U8352 (N_8352,N_7873,N_8006);
nor U8353 (N_8353,N_8018,N_7852);
or U8354 (N_8354,N_7964,N_7944);
nand U8355 (N_8355,N_8053,N_7836);
xor U8356 (N_8356,N_8089,N_7820);
and U8357 (N_8357,N_7877,N_7851);
or U8358 (N_8358,N_7879,N_7973);
xnor U8359 (N_8359,N_7878,N_7997);
nor U8360 (N_8360,N_7918,N_7978);
xnor U8361 (N_8361,N_7898,N_7893);
or U8362 (N_8362,N_8084,N_7990);
or U8363 (N_8363,N_7928,N_8055);
or U8364 (N_8364,N_8026,N_7826);
nand U8365 (N_8365,N_7828,N_7863);
nor U8366 (N_8366,N_7875,N_7834);
and U8367 (N_8367,N_7998,N_8052);
xnor U8368 (N_8368,N_8065,N_8082);
xnor U8369 (N_8369,N_8042,N_7880);
nand U8370 (N_8370,N_8064,N_7963);
nor U8371 (N_8371,N_7935,N_7833);
and U8372 (N_8372,N_7913,N_8048);
nand U8373 (N_8373,N_7817,N_7927);
xnor U8374 (N_8374,N_7942,N_7936);
nor U8375 (N_8375,N_7809,N_7915);
xor U8376 (N_8376,N_7802,N_7989);
nand U8377 (N_8377,N_7926,N_7995);
nor U8378 (N_8378,N_7949,N_8043);
or U8379 (N_8379,N_7806,N_7844);
nor U8380 (N_8380,N_7883,N_7963);
or U8381 (N_8381,N_8076,N_8032);
and U8382 (N_8382,N_7836,N_7801);
nand U8383 (N_8383,N_7898,N_7947);
or U8384 (N_8384,N_7908,N_7858);
and U8385 (N_8385,N_7935,N_8070);
xor U8386 (N_8386,N_7872,N_7807);
and U8387 (N_8387,N_7818,N_7865);
and U8388 (N_8388,N_8091,N_7819);
and U8389 (N_8389,N_7937,N_8081);
and U8390 (N_8390,N_8039,N_8013);
or U8391 (N_8391,N_7901,N_8097);
or U8392 (N_8392,N_8041,N_7999);
xor U8393 (N_8393,N_7954,N_8060);
nand U8394 (N_8394,N_8084,N_7818);
and U8395 (N_8395,N_7824,N_8090);
nand U8396 (N_8396,N_7902,N_8005);
and U8397 (N_8397,N_7980,N_8019);
xor U8398 (N_8398,N_7869,N_8017);
or U8399 (N_8399,N_8044,N_7878);
nor U8400 (N_8400,N_8301,N_8156);
nand U8401 (N_8401,N_8363,N_8125);
or U8402 (N_8402,N_8333,N_8190);
nor U8403 (N_8403,N_8145,N_8211);
or U8404 (N_8404,N_8329,N_8216);
nor U8405 (N_8405,N_8326,N_8116);
nand U8406 (N_8406,N_8210,N_8318);
xor U8407 (N_8407,N_8105,N_8205);
nor U8408 (N_8408,N_8246,N_8235);
nor U8409 (N_8409,N_8231,N_8163);
nand U8410 (N_8410,N_8239,N_8154);
nand U8411 (N_8411,N_8153,N_8300);
or U8412 (N_8412,N_8142,N_8180);
xor U8413 (N_8413,N_8152,N_8327);
xnor U8414 (N_8414,N_8330,N_8174);
or U8415 (N_8415,N_8214,N_8126);
and U8416 (N_8416,N_8387,N_8218);
xor U8417 (N_8417,N_8147,N_8386);
nand U8418 (N_8418,N_8309,N_8134);
or U8419 (N_8419,N_8340,N_8259);
nor U8420 (N_8420,N_8306,N_8117);
nand U8421 (N_8421,N_8391,N_8290);
xnor U8422 (N_8422,N_8398,N_8118);
or U8423 (N_8423,N_8222,N_8230);
nor U8424 (N_8424,N_8279,N_8351);
xor U8425 (N_8425,N_8352,N_8191);
xnor U8426 (N_8426,N_8269,N_8292);
xnor U8427 (N_8427,N_8106,N_8114);
xor U8428 (N_8428,N_8171,N_8139);
and U8429 (N_8429,N_8347,N_8354);
and U8430 (N_8430,N_8291,N_8141);
nor U8431 (N_8431,N_8220,N_8249);
nor U8432 (N_8432,N_8315,N_8332);
or U8433 (N_8433,N_8227,N_8388);
and U8434 (N_8434,N_8295,N_8375);
or U8435 (N_8435,N_8189,N_8202);
nand U8436 (N_8436,N_8208,N_8353);
nand U8437 (N_8437,N_8167,N_8224);
nand U8438 (N_8438,N_8390,N_8150);
nand U8439 (N_8439,N_8339,N_8135);
or U8440 (N_8440,N_8314,N_8286);
xnor U8441 (N_8441,N_8376,N_8273);
nor U8442 (N_8442,N_8251,N_8337);
or U8443 (N_8443,N_8252,N_8275);
nand U8444 (N_8444,N_8313,N_8158);
xor U8445 (N_8445,N_8360,N_8317);
nor U8446 (N_8446,N_8304,N_8209);
nand U8447 (N_8447,N_8311,N_8155);
or U8448 (N_8448,N_8392,N_8272);
or U8449 (N_8449,N_8103,N_8120);
nand U8450 (N_8450,N_8395,N_8350);
and U8451 (N_8451,N_8284,N_8133);
nor U8452 (N_8452,N_8123,N_8294);
or U8453 (N_8453,N_8336,N_8207);
or U8454 (N_8454,N_8299,N_8308);
nand U8455 (N_8455,N_8271,N_8267);
nor U8456 (N_8456,N_8138,N_8128);
nor U8457 (N_8457,N_8185,N_8377);
nor U8458 (N_8458,N_8338,N_8260);
nor U8459 (N_8459,N_8248,N_8172);
xnor U8460 (N_8460,N_8215,N_8140);
and U8461 (N_8461,N_8255,N_8241);
nor U8462 (N_8462,N_8240,N_8162);
or U8463 (N_8463,N_8266,N_8320);
xor U8464 (N_8464,N_8293,N_8369);
xnor U8465 (N_8465,N_8157,N_8285);
or U8466 (N_8466,N_8362,N_8223);
or U8467 (N_8467,N_8345,N_8198);
nand U8468 (N_8468,N_8217,N_8161);
nand U8469 (N_8469,N_8199,N_8335);
nor U8470 (N_8470,N_8371,N_8358);
or U8471 (N_8471,N_8316,N_8264);
xor U8472 (N_8472,N_8160,N_8121);
nand U8473 (N_8473,N_8247,N_8281);
or U8474 (N_8474,N_8130,N_8393);
and U8475 (N_8475,N_8184,N_8280);
nand U8476 (N_8476,N_8288,N_8378);
and U8477 (N_8477,N_8245,N_8151);
and U8478 (N_8478,N_8197,N_8310);
xor U8479 (N_8479,N_8312,N_8107);
nor U8480 (N_8480,N_8263,N_8226);
nand U8481 (N_8481,N_8177,N_8319);
or U8482 (N_8482,N_8183,N_8349);
and U8483 (N_8483,N_8144,N_8195);
xor U8484 (N_8484,N_8364,N_8397);
and U8485 (N_8485,N_8149,N_8385);
nor U8486 (N_8486,N_8127,N_8297);
or U8487 (N_8487,N_8256,N_8379);
nand U8488 (N_8488,N_8146,N_8348);
nand U8489 (N_8489,N_8307,N_8206);
nand U8490 (N_8490,N_8282,N_8303);
xor U8491 (N_8491,N_8182,N_8221);
and U8492 (N_8492,N_8186,N_8173);
or U8493 (N_8493,N_8170,N_8178);
or U8494 (N_8494,N_8359,N_8112);
or U8495 (N_8495,N_8165,N_8334);
xnor U8496 (N_8496,N_8225,N_8396);
nor U8497 (N_8497,N_8324,N_8229);
or U8498 (N_8498,N_8296,N_8305);
or U8499 (N_8499,N_8110,N_8361);
xor U8500 (N_8500,N_8382,N_8356);
nand U8501 (N_8501,N_8113,N_8366);
and U8502 (N_8502,N_8270,N_8200);
or U8503 (N_8503,N_8373,N_8322);
xnor U8504 (N_8504,N_8115,N_8236);
nand U8505 (N_8505,N_8384,N_8261);
nand U8506 (N_8506,N_8268,N_8302);
nor U8507 (N_8507,N_8129,N_8283);
xnor U8508 (N_8508,N_8242,N_8323);
or U8509 (N_8509,N_8321,N_8325);
nor U8510 (N_8510,N_8394,N_8254);
nand U8511 (N_8511,N_8109,N_8357);
and U8512 (N_8512,N_8342,N_8212);
and U8513 (N_8513,N_8346,N_8381);
and U8514 (N_8514,N_8343,N_8237);
xor U8515 (N_8515,N_8399,N_8278);
xnor U8516 (N_8516,N_8374,N_8257);
nand U8517 (N_8517,N_8213,N_8370);
xor U8518 (N_8518,N_8159,N_8203);
and U8519 (N_8519,N_8101,N_8287);
xor U8520 (N_8520,N_8262,N_8367);
nand U8521 (N_8521,N_8274,N_8244);
nand U8522 (N_8522,N_8250,N_8298);
xnor U8523 (N_8523,N_8131,N_8119);
nand U8524 (N_8524,N_8108,N_8124);
or U8525 (N_8525,N_8233,N_8258);
xor U8526 (N_8526,N_8100,N_8276);
xor U8527 (N_8527,N_8234,N_8368);
nor U8528 (N_8528,N_8204,N_8164);
and U8529 (N_8529,N_8389,N_8232);
or U8530 (N_8530,N_8136,N_8277);
or U8531 (N_8531,N_8201,N_8102);
nand U8532 (N_8532,N_8265,N_8194);
nand U8533 (N_8533,N_8181,N_8228);
xor U8534 (N_8534,N_8253,N_8365);
xnor U8535 (N_8535,N_8380,N_8192);
and U8536 (N_8536,N_8289,N_8179);
nor U8537 (N_8537,N_8193,N_8176);
xor U8538 (N_8538,N_8169,N_8328);
and U8539 (N_8539,N_8383,N_8187);
nand U8540 (N_8540,N_8196,N_8122);
or U8541 (N_8541,N_8104,N_8166);
xor U8542 (N_8542,N_8148,N_8219);
and U8543 (N_8543,N_8143,N_8344);
nor U8544 (N_8544,N_8331,N_8137);
nand U8545 (N_8545,N_8238,N_8243);
xor U8546 (N_8546,N_8341,N_8372);
or U8547 (N_8547,N_8168,N_8355);
xor U8548 (N_8548,N_8188,N_8111);
xnor U8549 (N_8549,N_8132,N_8175);
or U8550 (N_8550,N_8374,N_8242);
and U8551 (N_8551,N_8103,N_8399);
or U8552 (N_8552,N_8274,N_8278);
and U8553 (N_8553,N_8263,N_8385);
xnor U8554 (N_8554,N_8302,N_8181);
nand U8555 (N_8555,N_8305,N_8249);
or U8556 (N_8556,N_8247,N_8334);
or U8557 (N_8557,N_8114,N_8377);
nand U8558 (N_8558,N_8308,N_8358);
nor U8559 (N_8559,N_8160,N_8347);
or U8560 (N_8560,N_8250,N_8312);
xor U8561 (N_8561,N_8112,N_8279);
xor U8562 (N_8562,N_8251,N_8196);
or U8563 (N_8563,N_8291,N_8353);
and U8564 (N_8564,N_8185,N_8128);
nor U8565 (N_8565,N_8256,N_8153);
xor U8566 (N_8566,N_8277,N_8261);
nor U8567 (N_8567,N_8212,N_8263);
nand U8568 (N_8568,N_8391,N_8352);
nor U8569 (N_8569,N_8210,N_8150);
nand U8570 (N_8570,N_8362,N_8194);
nor U8571 (N_8571,N_8348,N_8382);
xnor U8572 (N_8572,N_8212,N_8275);
nand U8573 (N_8573,N_8328,N_8299);
nand U8574 (N_8574,N_8219,N_8127);
nor U8575 (N_8575,N_8203,N_8346);
or U8576 (N_8576,N_8170,N_8163);
and U8577 (N_8577,N_8390,N_8356);
or U8578 (N_8578,N_8138,N_8347);
nand U8579 (N_8579,N_8388,N_8291);
xor U8580 (N_8580,N_8135,N_8371);
or U8581 (N_8581,N_8379,N_8174);
or U8582 (N_8582,N_8319,N_8145);
or U8583 (N_8583,N_8197,N_8114);
nor U8584 (N_8584,N_8157,N_8284);
xor U8585 (N_8585,N_8191,N_8139);
and U8586 (N_8586,N_8353,N_8121);
and U8587 (N_8587,N_8154,N_8257);
nand U8588 (N_8588,N_8126,N_8299);
xnor U8589 (N_8589,N_8396,N_8117);
or U8590 (N_8590,N_8201,N_8374);
xnor U8591 (N_8591,N_8365,N_8313);
or U8592 (N_8592,N_8238,N_8242);
xnor U8593 (N_8593,N_8237,N_8259);
and U8594 (N_8594,N_8106,N_8179);
and U8595 (N_8595,N_8257,N_8148);
xnor U8596 (N_8596,N_8156,N_8129);
nand U8597 (N_8597,N_8149,N_8314);
or U8598 (N_8598,N_8219,N_8381);
xor U8599 (N_8599,N_8202,N_8201);
nor U8600 (N_8600,N_8323,N_8298);
nor U8601 (N_8601,N_8368,N_8320);
nand U8602 (N_8602,N_8294,N_8391);
nor U8603 (N_8603,N_8372,N_8242);
and U8604 (N_8604,N_8102,N_8198);
or U8605 (N_8605,N_8141,N_8399);
xnor U8606 (N_8606,N_8222,N_8134);
xnor U8607 (N_8607,N_8297,N_8136);
or U8608 (N_8608,N_8120,N_8109);
nand U8609 (N_8609,N_8202,N_8215);
nor U8610 (N_8610,N_8200,N_8286);
and U8611 (N_8611,N_8389,N_8204);
or U8612 (N_8612,N_8345,N_8202);
nand U8613 (N_8613,N_8270,N_8396);
or U8614 (N_8614,N_8163,N_8237);
nor U8615 (N_8615,N_8155,N_8333);
xor U8616 (N_8616,N_8388,N_8349);
nand U8617 (N_8617,N_8196,N_8181);
or U8618 (N_8618,N_8206,N_8163);
or U8619 (N_8619,N_8338,N_8393);
nand U8620 (N_8620,N_8271,N_8187);
xnor U8621 (N_8621,N_8284,N_8392);
nor U8622 (N_8622,N_8329,N_8101);
xnor U8623 (N_8623,N_8205,N_8243);
nand U8624 (N_8624,N_8244,N_8352);
xnor U8625 (N_8625,N_8248,N_8273);
nor U8626 (N_8626,N_8394,N_8311);
and U8627 (N_8627,N_8354,N_8209);
nor U8628 (N_8628,N_8108,N_8174);
or U8629 (N_8629,N_8271,N_8239);
nor U8630 (N_8630,N_8259,N_8248);
nand U8631 (N_8631,N_8313,N_8251);
nor U8632 (N_8632,N_8127,N_8269);
nor U8633 (N_8633,N_8194,N_8179);
nor U8634 (N_8634,N_8172,N_8263);
or U8635 (N_8635,N_8232,N_8295);
and U8636 (N_8636,N_8380,N_8120);
nand U8637 (N_8637,N_8147,N_8312);
and U8638 (N_8638,N_8272,N_8247);
xnor U8639 (N_8639,N_8192,N_8315);
xnor U8640 (N_8640,N_8347,N_8151);
or U8641 (N_8641,N_8230,N_8172);
or U8642 (N_8642,N_8160,N_8337);
or U8643 (N_8643,N_8336,N_8111);
or U8644 (N_8644,N_8386,N_8330);
nand U8645 (N_8645,N_8149,N_8292);
nand U8646 (N_8646,N_8276,N_8333);
nand U8647 (N_8647,N_8190,N_8313);
nor U8648 (N_8648,N_8127,N_8133);
nand U8649 (N_8649,N_8142,N_8114);
xnor U8650 (N_8650,N_8398,N_8302);
or U8651 (N_8651,N_8297,N_8261);
nand U8652 (N_8652,N_8386,N_8117);
nand U8653 (N_8653,N_8310,N_8303);
or U8654 (N_8654,N_8357,N_8284);
xor U8655 (N_8655,N_8114,N_8214);
xor U8656 (N_8656,N_8310,N_8123);
or U8657 (N_8657,N_8134,N_8109);
nand U8658 (N_8658,N_8387,N_8132);
nand U8659 (N_8659,N_8139,N_8162);
nand U8660 (N_8660,N_8339,N_8197);
or U8661 (N_8661,N_8291,N_8185);
xor U8662 (N_8662,N_8239,N_8135);
xnor U8663 (N_8663,N_8389,N_8193);
xor U8664 (N_8664,N_8268,N_8158);
xnor U8665 (N_8665,N_8182,N_8200);
and U8666 (N_8666,N_8337,N_8138);
and U8667 (N_8667,N_8173,N_8288);
or U8668 (N_8668,N_8338,N_8109);
nor U8669 (N_8669,N_8201,N_8289);
xor U8670 (N_8670,N_8383,N_8132);
or U8671 (N_8671,N_8200,N_8394);
or U8672 (N_8672,N_8240,N_8307);
nand U8673 (N_8673,N_8369,N_8200);
nor U8674 (N_8674,N_8205,N_8208);
or U8675 (N_8675,N_8229,N_8119);
and U8676 (N_8676,N_8293,N_8150);
or U8677 (N_8677,N_8221,N_8303);
nor U8678 (N_8678,N_8283,N_8209);
nor U8679 (N_8679,N_8111,N_8253);
nand U8680 (N_8680,N_8331,N_8158);
xnor U8681 (N_8681,N_8249,N_8300);
or U8682 (N_8682,N_8282,N_8317);
nand U8683 (N_8683,N_8192,N_8143);
xnor U8684 (N_8684,N_8103,N_8342);
and U8685 (N_8685,N_8296,N_8185);
and U8686 (N_8686,N_8193,N_8217);
nand U8687 (N_8687,N_8175,N_8167);
nor U8688 (N_8688,N_8287,N_8244);
nand U8689 (N_8689,N_8182,N_8191);
and U8690 (N_8690,N_8282,N_8245);
and U8691 (N_8691,N_8342,N_8277);
nand U8692 (N_8692,N_8315,N_8239);
nor U8693 (N_8693,N_8106,N_8305);
and U8694 (N_8694,N_8217,N_8206);
xor U8695 (N_8695,N_8258,N_8238);
xor U8696 (N_8696,N_8214,N_8346);
nand U8697 (N_8697,N_8363,N_8293);
and U8698 (N_8698,N_8130,N_8321);
xnor U8699 (N_8699,N_8383,N_8391);
nand U8700 (N_8700,N_8472,N_8619);
nor U8701 (N_8701,N_8586,N_8560);
nor U8702 (N_8702,N_8431,N_8682);
and U8703 (N_8703,N_8425,N_8649);
nand U8704 (N_8704,N_8426,N_8508);
nand U8705 (N_8705,N_8666,N_8630);
and U8706 (N_8706,N_8443,N_8541);
xnor U8707 (N_8707,N_8640,N_8579);
or U8708 (N_8708,N_8684,N_8459);
or U8709 (N_8709,N_8435,N_8688);
nor U8710 (N_8710,N_8632,N_8520);
nand U8711 (N_8711,N_8618,N_8698);
or U8712 (N_8712,N_8559,N_8518);
and U8713 (N_8713,N_8599,N_8625);
nand U8714 (N_8714,N_8552,N_8661);
nor U8715 (N_8715,N_8416,N_8571);
or U8716 (N_8716,N_8486,N_8617);
nor U8717 (N_8717,N_8580,N_8608);
and U8718 (N_8718,N_8536,N_8500);
nor U8719 (N_8719,N_8653,N_8525);
xor U8720 (N_8720,N_8457,N_8427);
nor U8721 (N_8721,N_8480,N_8503);
and U8722 (N_8722,N_8411,N_8695);
nor U8723 (N_8723,N_8643,N_8658);
and U8724 (N_8724,N_8495,N_8657);
or U8725 (N_8725,N_8476,N_8590);
nand U8726 (N_8726,N_8672,N_8542);
nand U8727 (N_8727,N_8696,N_8568);
nand U8728 (N_8728,N_8497,N_8417);
nor U8729 (N_8729,N_8422,N_8401);
or U8730 (N_8730,N_8467,N_8504);
or U8731 (N_8731,N_8488,N_8523);
xnor U8732 (N_8732,N_8670,N_8479);
or U8733 (N_8733,N_8626,N_8623);
xnor U8734 (N_8734,N_8487,N_8515);
xor U8735 (N_8735,N_8470,N_8464);
xor U8736 (N_8736,N_8562,N_8613);
and U8737 (N_8737,N_8578,N_8421);
nand U8738 (N_8738,N_8535,N_8496);
xor U8739 (N_8739,N_8585,N_8573);
and U8740 (N_8740,N_8668,N_8442);
xnor U8741 (N_8741,N_8642,N_8544);
nand U8742 (N_8742,N_8566,N_8655);
nand U8743 (N_8743,N_8533,N_8483);
or U8744 (N_8744,N_8597,N_8678);
xor U8745 (N_8745,N_8663,N_8538);
or U8746 (N_8746,N_8424,N_8452);
and U8747 (N_8747,N_8635,N_8582);
and U8748 (N_8748,N_8673,N_8647);
nor U8749 (N_8749,N_8412,N_8569);
and U8750 (N_8750,N_8434,N_8689);
nor U8751 (N_8751,N_8546,N_8437);
xor U8752 (N_8752,N_8505,N_8662);
and U8753 (N_8753,N_8502,N_8664);
xnor U8754 (N_8754,N_8484,N_8547);
xnor U8755 (N_8755,N_8624,N_8561);
and U8756 (N_8756,N_8641,N_8529);
or U8757 (N_8757,N_8448,N_8687);
or U8758 (N_8758,N_8444,N_8469);
and U8759 (N_8759,N_8592,N_8446);
xor U8760 (N_8760,N_8419,N_8473);
xor U8761 (N_8761,N_8548,N_8636);
nor U8762 (N_8762,N_8414,N_8492);
nor U8763 (N_8763,N_8438,N_8455);
nor U8764 (N_8764,N_8622,N_8449);
xnor U8765 (N_8765,N_8587,N_8506);
xor U8766 (N_8766,N_8601,N_8403);
and U8767 (N_8767,N_8517,N_8602);
and U8768 (N_8768,N_8699,N_8621);
nor U8769 (N_8769,N_8482,N_8441);
nand U8770 (N_8770,N_8490,N_8567);
nand U8771 (N_8771,N_8491,N_8671);
or U8772 (N_8772,N_8454,N_8501);
nand U8773 (N_8773,N_8596,N_8588);
or U8774 (N_8774,N_8679,N_8609);
nand U8775 (N_8775,N_8514,N_8477);
nor U8776 (N_8776,N_8408,N_8516);
or U8777 (N_8777,N_8659,N_8453);
and U8778 (N_8778,N_8557,N_8512);
xnor U8779 (N_8779,N_8634,N_8558);
nand U8780 (N_8780,N_8526,N_8674);
xnor U8781 (N_8781,N_8451,N_8584);
xor U8782 (N_8782,N_8598,N_8400);
or U8783 (N_8783,N_8406,N_8466);
and U8784 (N_8784,N_8474,N_8428);
nand U8785 (N_8785,N_8697,N_8583);
nand U8786 (N_8786,N_8494,N_8651);
and U8787 (N_8787,N_8550,N_8530);
nand U8788 (N_8788,N_8534,N_8549);
and U8789 (N_8789,N_8461,N_8681);
and U8790 (N_8790,N_8633,N_8439);
and U8791 (N_8791,N_8574,N_8648);
or U8792 (N_8792,N_8519,N_8570);
nor U8793 (N_8793,N_8652,N_8691);
or U8794 (N_8794,N_8465,N_8595);
nor U8795 (N_8795,N_8460,N_8611);
and U8796 (N_8796,N_8540,N_8654);
nor U8797 (N_8797,N_8436,N_8450);
and U8798 (N_8798,N_8667,N_8620);
nor U8799 (N_8799,N_8565,N_8686);
nand U8800 (N_8800,N_8509,N_8627);
or U8801 (N_8801,N_8410,N_8458);
nand U8802 (N_8802,N_8615,N_8507);
and U8803 (N_8803,N_8591,N_8471);
nor U8804 (N_8804,N_8528,N_8554);
nor U8805 (N_8805,N_8575,N_8527);
or U8806 (N_8806,N_8481,N_8612);
nor U8807 (N_8807,N_8493,N_8551);
or U8808 (N_8808,N_8628,N_8631);
nand U8809 (N_8809,N_8489,N_8485);
and U8810 (N_8810,N_8430,N_8420);
and U8811 (N_8811,N_8407,N_8593);
or U8812 (N_8812,N_8676,N_8532);
nor U8813 (N_8813,N_8610,N_8510);
nor U8814 (N_8814,N_8603,N_8607);
or U8815 (N_8815,N_8462,N_8616);
or U8816 (N_8816,N_8475,N_8604);
nor U8817 (N_8817,N_8629,N_8415);
xnor U8818 (N_8818,N_8677,N_8440);
xor U8819 (N_8819,N_8429,N_8650);
or U8820 (N_8820,N_8638,N_8690);
nor U8821 (N_8821,N_8683,N_8445);
and U8822 (N_8822,N_8577,N_8433);
nand U8823 (N_8823,N_8555,N_8511);
xor U8824 (N_8824,N_8564,N_8675);
and U8825 (N_8825,N_8693,N_8637);
and U8826 (N_8826,N_8669,N_8543);
xnor U8827 (N_8827,N_8513,N_8539);
nor U8828 (N_8828,N_8614,N_8645);
and U8829 (N_8829,N_8685,N_8537);
nand U8830 (N_8830,N_8522,N_8594);
and U8831 (N_8831,N_8589,N_8524);
and U8832 (N_8832,N_8456,N_8463);
nand U8833 (N_8833,N_8639,N_8405);
and U8834 (N_8834,N_8423,N_8665);
nand U8835 (N_8835,N_8531,N_8498);
or U8836 (N_8836,N_8556,N_8600);
nand U8837 (N_8837,N_8478,N_8646);
and U8838 (N_8838,N_8660,N_8432);
nand U8839 (N_8839,N_8499,N_8581);
nor U8840 (N_8840,N_8545,N_8680);
nand U8841 (N_8841,N_8656,N_8553);
nand U8842 (N_8842,N_8605,N_8521);
or U8843 (N_8843,N_8644,N_8576);
xnor U8844 (N_8844,N_8694,N_8563);
and U8845 (N_8845,N_8606,N_8409);
xnor U8846 (N_8846,N_8468,N_8404);
nand U8847 (N_8847,N_8692,N_8572);
and U8848 (N_8848,N_8413,N_8447);
and U8849 (N_8849,N_8402,N_8418);
xor U8850 (N_8850,N_8530,N_8617);
xor U8851 (N_8851,N_8599,N_8450);
xor U8852 (N_8852,N_8532,N_8529);
xor U8853 (N_8853,N_8679,N_8506);
and U8854 (N_8854,N_8490,N_8613);
xnor U8855 (N_8855,N_8433,N_8601);
nand U8856 (N_8856,N_8424,N_8685);
nand U8857 (N_8857,N_8432,N_8618);
and U8858 (N_8858,N_8570,N_8448);
nand U8859 (N_8859,N_8502,N_8643);
nand U8860 (N_8860,N_8411,N_8697);
nor U8861 (N_8861,N_8585,N_8555);
nand U8862 (N_8862,N_8609,N_8684);
and U8863 (N_8863,N_8408,N_8698);
nor U8864 (N_8864,N_8518,N_8614);
nand U8865 (N_8865,N_8547,N_8608);
nand U8866 (N_8866,N_8630,N_8675);
nor U8867 (N_8867,N_8614,N_8556);
nand U8868 (N_8868,N_8499,N_8544);
or U8869 (N_8869,N_8528,N_8473);
nor U8870 (N_8870,N_8527,N_8510);
nand U8871 (N_8871,N_8543,N_8503);
and U8872 (N_8872,N_8498,N_8678);
xnor U8873 (N_8873,N_8650,N_8472);
and U8874 (N_8874,N_8615,N_8551);
nor U8875 (N_8875,N_8544,N_8480);
xor U8876 (N_8876,N_8450,N_8533);
nor U8877 (N_8877,N_8403,N_8612);
nand U8878 (N_8878,N_8663,N_8457);
or U8879 (N_8879,N_8624,N_8438);
nor U8880 (N_8880,N_8461,N_8459);
nand U8881 (N_8881,N_8657,N_8650);
nand U8882 (N_8882,N_8635,N_8521);
xor U8883 (N_8883,N_8467,N_8670);
nor U8884 (N_8884,N_8663,N_8523);
and U8885 (N_8885,N_8548,N_8506);
and U8886 (N_8886,N_8617,N_8642);
nand U8887 (N_8887,N_8427,N_8669);
nand U8888 (N_8888,N_8658,N_8582);
and U8889 (N_8889,N_8508,N_8685);
nand U8890 (N_8890,N_8504,N_8495);
nand U8891 (N_8891,N_8493,N_8627);
or U8892 (N_8892,N_8602,N_8453);
or U8893 (N_8893,N_8633,N_8478);
xor U8894 (N_8894,N_8665,N_8474);
xnor U8895 (N_8895,N_8405,N_8603);
nor U8896 (N_8896,N_8591,N_8667);
xor U8897 (N_8897,N_8482,N_8501);
or U8898 (N_8898,N_8501,N_8505);
and U8899 (N_8899,N_8423,N_8543);
and U8900 (N_8900,N_8445,N_8414);
xnor U8901 (N_8901,N_8618,N_8616);
nor U8902 (N_8902,N_8522,N_8695);
or U8903 (N_8903,N_8648,N_8577);
nor U8904 (N_8904,N_8477,N_8620);
or U8905 (N_8905,N_8407,N_8495);
or U8906 (N_8906,N_8539,N_8508);
xor U8907 (N_8907,N_8439,N_8572);
xnor U8908 (N_8908,N_8541,N_8625);
xnor U8909 (N_8909,N_8429,N_8432);
nor U8910 (N_8910,N_8402,N_8614);
nand U8911 (N_8911,N_8474,N_8669);
and U8912 (N_8912,N_8528,N_8603);
or U8913 (N_8913,N_8618,N_8534);
nand U8914 (N_8914,N_8581,N_8684);
or U8915 (N_8915,N_8689,N_8606);
xnor U8916 (N_8916,N_8501,N_8537);
nor U8917 (N_8917,N_8452,N_8563);
and U8918 (N_8918,N_8644,N_8476);
or U8919 (N_8919,N_8669,N_8688);
nor U8920 (N_8920,N_8528,N_8520);
and U8921 (N_8921,N_8534,N_8691);
nand U8922 (N_8922,N_8615,N_8594);
or U8923 (N_8923,N_8552,N_8437);
or U8924 (N_8924,N_8459,N_8421);
xor U8925 (N_8925,N_8459,N_8538);
nor U8926 (N_8926,N_8405,N_8453);
nor U8927 (N_8927,N_8463,N_8659);
or U8928 (N_8928,N_8668,N_8459);
xnor U8929 (N_8929,N_8548,N_8557);
or U8930 (N_8930,N_8437,N_8637);
or U8931 (N_8931,N_8592,N_8467);
nand U8932 (N_8932,N_8402,N_8470);
or U8933 (N_8933,N_8604,N_8544);
and U8934 (N_8934,N_8423,N_8529);
xnor U8935 (N_8935,N_8550,N_8613);
or U8936 (N_8936,N_8674,N_8549);
nor U8937 (N_8937,N_8437,N_8525);
nor U8938 (N_8938,N_8408,N_8586);
nor U8939 (N_8939,N_8489,N_8651);
or U8940 (N_8940,N_8443,N_8680);
and U8941 (N_8941,N_8435,N_8670);
nor U8942 (N_8942,N_8478,N_8569);
nand U8943 (N_8943,N_8524,N_8421);
nor U8944 (N_8944,N_8423,N_8556);
nand U8945 (N_8945,N_8545,N_8607);
nor U8946 (N_8946,N_8511,N_8452);
or U8947 (N_8947,N_8633,N_8518);
xor U8948 (N_8948,N_8404,N_8623);
nand U8949 (N_8949,N_8550,N_8465);
or U8950 (N_8950,N_8600,N_8441);
nand U8951 (N_8951,N_8475,N_8483);
and U8952 (N_8952,N_8435,N_8522);
nor U8953 (N_8953,N_8509,N_8673);
nor U8954 (N_8954,N_8696,N_8461);
nand U8955 (N_8955,N_8472,N_8629);
and U8956 (N_8956,N_8477,N_8518);
and U8957 (N_8957,N_8603,N_8667);
nor U8958 (N_8958,N_8499,N_8663);
nand U8959 (N_8959,N_8605,N_8691);
or U8960 (N_8960,N_8512,N_8589);
xnor U8961 (N_8961,N_8452,N_8481);
and U8962 (N_8962,N_8679,N_8690);
or U8963 (N_8963,N_8629,N_8438);
nor U8964 (N_8964,N_8621,N_8546);
and U8965 (N_8965,N_8472,N_8568);
nand U8966 (N_8966,N_8567,N_8515);
and U8967 (N_8967,N_8523,N_8582);
and U8968 (N_8968,N_8429,N_8420);
xor U8969 (N_8969,N_8662,N_8441);
nand U8970 (N_8970,N_8573,N_8681);
xnor U8971 (N_8971,N_8570,N_8496);
nor U8972 (N_8972,N_8574,N_8441);
xor U8973 (N_8973,N_8433,N_8643);
and U8974 (N_8974,N_8518,N_8500);
and U8975 (N_8975,N_8697,N_8582);
xnor U8976 (N_8976,N_8553,N_8630);
or U8977 (N_8977,N_8549,N_8615);
nand U8978 (N_8978,N_8564,N_8663);
and U8979 (N_8979,N_8493,N_8682);
nand U8980 (N_8980,N_8605,N_8506);
and U8981 (N_8981,N_8543,N_8656);
nand U8982 (N_8982,N_8512,N_8657);
nor U8983 (N_8983,N_8426,N_8674);
xnor U8984 (N_8984,N_8427,N_8482);
xnor U8985 (N_8985,N_8633,N_8442);
nor U8986 (N_8986,N_8696,N_8508);
and U8987 (N_8987,N_8524,N_8557);
nand U8988 (N_8988,N_8572,N_8407);
or U8989 (N_8989,N_8544,N_8492);
xnor U8990 (N_8990,N_8525,N_8666);
xor U8991 (N_8991,N_8685,N_8487);
nand U8992 (N_8992,N_8433,N_8644);
xor U8993 (N_8993,N_8456,N_8623);
nand U8994 (N_8994,N_8461,N_8575);
xnor U8995 (N_8995,N_8455,N_8434);
nand U8996 (N_8996,N_8623,N_8643);
nand U8997 (N_8997,N_8534,N_8679);
nor U8998 (N_8998,N_8666,N_8437);
or U8999 (N_8999,N_8411,N_8424);
nand U9000 (N_9000,N_8979,N_8921);
nor U9001 (N_9001,N_8822,N_8932);
nor U9002 (N_9002,N_8842,N_8915);
nand U9003 (N_9003,N_8759,N_8919);
nor U9004 (N_9004,N_8729,N_8821);
or U9005 (N_9005,N_8862,N_8866);
and U9006 (N_9006,N_8793,N_8951);
nor U9007 (N_9007,N_8788,N_8723);
nand U9008 (N_9008,N_8733,N_8929);
nand U9009 (N_9009,N_8827,N_8888);
nand U9010 (N_9010,N_8976,N_8839);
or U9011 (N_9011,N_8844,N_8909);
or U9012 (N_9012,N_8837,N_8703);
nor U9013 (N_9013,N_8900,N_8934);
nor U9014 (N_9014,N_8717,N_8949);
nand U9015 (N_9015,N_8722,N_8969);
and U9016 (N_9016,N_8987,N_8700);
or U9017 (N_9017,N_8803,N_8898);
xor U9018 (N_9018,N_8805,N_8928);
nor U9019 (N_9019,N_8778,N_8876);
nand U9020 (N_9020,N_8799,N_8754);
nand U9021 (N_9021,N_8871,N_8953);
or U9022 (N_9022,N_8978,N_8774);
nor U9023 (N_9023,N_8742,N_8920);
and U9024 (N_9024,N_8877,N_8975);
nor U9025 (N_9025,N_8814,N_8972);
or U9026 (N_9026,N_8776,N_8791);
nor U9027 (N_9027,N_8829,N_8771);
or U9028 (N_9028,N_8835,N_8780);
nor U9029 (N_9029,N_8712,N_8811);
or U9030 (N_9030,N_8935,N_8859);
and U9031 (N_9031,N_8707,N_8738);
and U9032 (N_9032,N_8881,N_8817);
nand U9033 (N_9033,N_8708,N_8794);
nor U9034 (N_9034,N_8907,N_8954);
or U9035 (N_9035,N_8850,N_8983);
or U9036 (N_9036,N_8783,N_8970);
and U9037 (N_9037,N_8767,N_8965);
xnor U9038 (N_9038,N_8816,N_8856);
or U9039 (N_9039,N_8705,N_8853);
nor U9040 (N_9040,N_8779,N_8724);
nand U9041 (N_9041,N_8746,N_8751);
nand U9042 (N_9042,N_8899,N_8818);
and U9043 (N_9043,N_8875,N_8865);
nand U9044 (N_9044,N_8873,N_8796);
and U9045 (N_9045,N_8937,N_8882);
and U9046 (N_9046,N_8913,N_8889);
nand U9047 (N_9047,N_8710,N_8996);
or U9048 (N_9048,N_8823,N_8936);
and U9049 (N_9049,N_8988,N_8752);
xor U9050 (N_9050,N_8906,N_8874);
and U9051 (N_9051,N_8897,N_8930);
or U9052 (N_9052,N_8880,N_8769);
nor U9053 (N_9053,N_8702,N_8834);
nor U9054 (N_9054,N_8838,N_8728);
xnor U9055 (N_9055,N_8739,N_8787);
nor U9056 (N_9056,N_8857,N_8872);
or U9057 (N_9057,N_8706,N_8721);
nand U9058 (N_9058,N_8768,N_8843);
nand U9059 (N_9059,N_8910,N_8826);
and U9060 (N_9060,N_8962,N_8786);
nand U9061 (N_9061,N_8955,N_8845);
nor U9062 (N_9062,N_8895,N_8918);
and U9063 (N_9063,N_8950,N_8775);
nor U9064 (N_9064,N_8961,N_8830);
nor U9065 (N_9065,N_8758,N_8896);
or U9066 (N_9066,N_8824,N_8938);
xor U9067 (N_9067,N_8958,N_8741);
and U9068 (N_9068,N_8841,N_8784);
and U9069 (N_9069,N_8781,N_8812);
and U9070 (N_9070,N_8851,N_8798);
xor U9071 (N_9071,N_8765,N_8763);
nand U9072 (N_9072,N_8736,N_8947);
and U9073 (N_9073,N_8870,N_8734);
nand U9074 (N_9074,N_8886,N_8737);
or U9075 (N_9075,N_8730,N_8815);
and U9076 (N_9076,N_8790,N_8755);
nor U9077 (N_9077,N_8740,N_8802);
nor U9078 (N_9078,N_8985,N_8840);
nor U9079 (N_9079,N_8847,N_8832);
nor U9080 (N_9080,N_8854,N_8861);
nor U9081 (N_9081,N_8743,N_8714);
xnor U9082 (N_9082,N_8891,N_8848);
or U9083 (N_9083,N_8719,N_8745);
nor U9084 (N_9084,N_8989,N_8789);
or U9085 (N_9085,N_8998,N_8809);
or U9086 (N_9086,N_8810,N_8792);
and U9087 (N_9087,N_8952,N_8849);
nor U9088 (N_9088,N_8960,N_8997);
and U9089 (N_9089,N_8766,N_8863);
nand U9090 (N_9090,N_8903,N_8933);
or U9091 (N_9091,N_8963,N_8939);
nor U9092 (N_9092,N_8764,N_8797);
or U9093 (N_9093,N_8864,N_8761);
and U9094 (N_9094,N_8868,N_8867);
nor U9095 (N_9095,N_8828,N_8749);
nor U9096 (N_9096,N_8804,N_8912);
or U9097 (N_9097,N_8924,N_8777);
xnor U9098 (N_9098,N_8760,N_8831);
nand U9099 (N_9099,N_8931,N_8825);
nor U9100 (N_9100,N_8990,N_8750);
xnor U9101 (N_9101,N_8715,N_8801);
xor U9102 (N_9102,N_8701,N_8991);
or U9103 (N_9103,N_8785,N_8883);
xor U9104 (N_9104,N_8852,N_8995);
and U9105 (N_9105,N_8981,N_8946);
or U9106 (N_9106,N_8709,N_8977);
and U9107 (N_9107,N_8948,N_8885);
or U9108 (N_9108,N_8968,N_8894);
or U9109 (N_9109,N_8993,N_8984);
or U9110 (N_9110,N_8860,N_8732);
nor U9111 (N_9111,N_8800,N_8902);
nor U9112 (N_9112,N_8711,N_8762);
nor U9113 (N_9113,N_8770,N_8893);
nor U9114 (N_9114,N_8942,N_8973);
and U9115 (N_9115,N_8846,N_8757);
xnor U9116 (N_9116,N_8748,N_8753);
and U9117 (N_9117,N_8772,N_8966);
and U9118 (N_9118,N_8994,N_8756);
nand U9119 (N_9119,N_8808,N_8904);
and U9120 (N_9120,N_8713,N_8806);
and U9121 (N_9121,N_8959,N_8890);
nor U9122 (N_9122,N_8858,N_8901);
and U9123 (N_9123,N_8726,N_8916);
and U9124 (N_9124,N_8725,N_8922);
nor U9125 (N_9125,N_8884,N_8944);
and U9126 (N_9126,N_8869,N_8911);
nor U9127 (N_9127,N_8782,N_8704);
nand U9128 (N_9128,N_8819,N_8999);
xor U9129 (N_9129,N_8744,N_8878);
nand U9130 (N_9130,N_8923,N_8855);
nor U9131 (N_9131,N_8720,N_8917);
nor U9132 (N_9132,N_8914,N_8887);
xor U9133 (N_9133,N_8982,N_8964);
nand U9134 (N_9134,N_8836,N_8892);
or U9135 (N_9135,N_8773,N_8956);
or U9136 (N_9136,N_8731,N_8820);
and U9137 (N_9137,N_8974,N_8747);
or U9138 (N_9138,N_8967,N_8833);
nor U9139 (N_9139,N_8905,N_8927);
nor U9140 (N_9140,N_8813,N_8971);
or U9141 (N_9141,N_8926,N_8727);
nor U9142 (N_9142,N_8718,N_8735);
xnor U9143 (N_9143,N_8908,N_8943);
and U9144 (N_9144,N_8992,N_8807);
nand U9145 (N_9145,N_8795,N_8716);
nand U9146 (N_9146,N_8879,N_8957);
xor U9147 (N_9147,N_8941,N_8945);
and U9148 (N_9148,N_8940,N_8986);
or U9149 (N_9149,N_8980,N_8925);
or U9150 (N_9150,N_8726,N_8875);
and U9151 (N_9151,N_8743,N_8703);
or U9152 (N_9152,N_8937,N_8729);
nand U9153 (N_9153,N_8845,N_8773);
xnor U9154 (N_9154,N_8862,N_8721);
nor U9155 (N_9155,N_8981,N_8976);
xor U9156 (N_9156,N_8899,N_8734);
nand U9157 (N_9157,N_8858,N_8804);
nor U9158 (N_9158,N_8885,N_8756);
nor U9159 (N_9159,N_8733,N_8911);
nor U9160 (N_9160,N_8711,N_8752);
nor U9161 (N_9161,N_8898,N_8820);
and U9162 (N_9162,N_8743,N_8983);
xor U9163 (N_9163,N_8931,N_8864);
and U9164 (N_9164,N_8852,N_8915);
nor U9165 (N_9165,N_8704,N_8913);
nand U9166 (N_9166,N_8898,N_8789);
or U9167 (N_9167,N_8789,N_8976);
or U9168 (N_9168,N_8901,N_8798);
nand U9169 (N_9169,N_8800,N_8944);
and U9170 (N_9170,N_8953,N_8779);
xor U9171 (N_9171,N_8797,N_8971);
and U9172 (N_9172,N_8973,N_8844);
nor U9173 (N_9173,N_8709,N_8733);
and U9174 (N_9174,N_8982,N_8981);
xor U9175 (N_9175,N_8834,N_8970);
nand U9176 (N_9176,N_8733,N_8792);
nand U9177 (N_9177,N_8812,N_8733);
and U9178 (N_9178,N_8726,N_8841);
nand U9179 (N_9179,N_8732,N_8769);
and U9180 (N_9180,N_8779,N_8944);
and U9181 (N_9181,N_8938,N_8819);
or U9182 (N_9182,N_8792,N_8885);
xor U9183 (N_9183,N_8788,N_8935);
xnor U9184 (N_9184,N_8810,N_8719);
xor U9185 (N_9185,N_8848,N_8958);
xor U9186 (N_9186,N_8834,N_8868);
nor U9187 (N_9187,N_8796,N_8710);
xnor U9188 (N_9188,N_8853,N_8943);
and U9189 (N_9189,N_8837,N_8896);
nor U9190 (N_9190,N_8876,N_8716);
nor U9191 (N_9191,N_8989,N_8838);
xor U9192 (N_9192,N_8979,N_8792);
and U9193 (N_9193,N_8847,N_8841);
nor U9194 (N_9194,N_8926,N_8811);
and U9195 (N_9195,N_8939,N_8949);
xor U9196 (N_9196,N_8987,N_8954);
nand U9197 (N_9197,N_8959,N_8834);
and U9198 (N_9198,N_8846,N_8909);
nor U9199 (N_9199,N_8859,N_8778);
nand U9200 (N_9200,N_8900,N_8702);
and U9201 (N_9201,N_8902,N_8903);
or U9202 (N_9202,N_8963,N_8744);
xor U9203 (N_9203,N_8994,N_8774);
and U9204 (N_9204,N_8902,N_8904);
nand U9205 (N_9205,N_8892,N_8765);
nor U9206 (N_9206,N_8811,N_8767);
nand U9207 (N_9207,N_8889,N_8928);
or U9208 (N_9208,N_8866,N_8826);
or U9209 (N_9209,N_8855,N_8942);
xor U9210 (N_9210,N_8903,N_8953);
nor U9211 (N_9211,N_8858,N_8956);
xor U9212 (N_9212,N_8912,N_8840);
and U9213 (N_9213,N_8729,N_8924);
or U9214 (N_9214,N_8761,N_8935);
or U9215 (N_9215,N_8912,N_8814);
nor U9216 (N_9216,N_8708,N_8922);
nand U9217 (N_9217,N_8988,N_8817);
nor U9218 (N_9218,N_8862,N_8820);
nand U9219 (N_9219,N_8808,N_8761);
or U9220 (N_9220,N_8762,N_8845);
nor U9221 (N_9221,N_8771,N_8785);
xor U9222 (N_9222,N_8901,N_8803);
and U9223 (N_9223,N_8853,N_8909);
nor U9224 (N_9224,N_8850,N_8999);
xor U9225 (N_9225,N_8856,N_8961);
xor U9226 (N_9226,N_8724,N_8700);
nor U9227 (N_9227,N_8955,N_8827);
or U9228 (N_9228,N_8994,N_8903);
and U9229 (N_9229,N_8887,N_8874);
xor U9230 (N_9230,N_8789,N_8722);
or U9231 (N_9231,N_8856,N_8781);
xnor U9232 (N_9232,N_8812,N_8805);
nor U9233 (N_9233,N_8893,N_8762);
xnor U9234 (N_9234,N_8837,N_8724);
nor U9235 (N_9235,N_8709,N_8904);
xnor U9236 (N_9236,N_8961,N_8892);
and U9237 (N_9237,N_8720,N_8703);
nand U9238 (N_9238,N_8968,N_8807);
or U9239 (N_9239,N_8736,N_8957);
nand U9240 (N_9240,N_8888,N_8904);
and U9241 (N_9241,N_8736,N_8929);
xnor U9242 (N_9242,N_8923,N_8762);
nand U9243 (N_9243,N_8849,N_8742);
nor U9244 (N_9244,N_8791,N_8834);
and U9245 (N_9245,N_8976,N_8809);
nand U9246 (N_9246,N_8829,N_8772);
nor U9247 (N_9247,N_8741,N_8831);
and U9248 (N_9248,N_8987,N_8885);
nor U9249 (N_9249,N_8885,N_8830);
nand U9250 (N_9250,N_8932,N_8710);
xnor U9251 (N_9251,N_8847,N_8949);
and U9252 (N_9252,N_8987,N_8875);
or U9253 (N_9253,N_8814,N_8932);
nor U9254 (N_9254,N_8887,N_8832);
xor U9255 (N_9255,N_8757,N_8976);
nor U9256 (N_9256,N_8998,N_8878);
and U9257 (N_9257,N_8776,N_8789);
nand U9258 (N_9258,N_8955,N_8860);
nand U9259 (N_9259,N_8701,N_8915);
or U9260 (N_9260,N_8753,N_8766);
nor U9261 (N_9261,N_8990,N_8948);
and U9262 (N_9262,N_8831,N_8930);
xor U9263 (N_9263,N_8956,N_8804);
or U9264 (N_9264,N_8952,N_8973);
and U9265 (N_9265,N_8964,N_8730);
or U9266 (N_9266,N_8786,N_8806);
nand U9267 (N_9267,N_8958,N_8824);
and U9268 (N_9268,N_8956,N_8946);
nand U9269 (N_9269,N_8956,N_8799);
and U9270 (N_9270,N_8937,N_8913);
xor U9271 (N_9271,N_8979,N_8761);
nand U9272 (N_9272,N_8920,N_8843);
and U9273 (N_9273,N_8881,N_8913);
xnor U9274 (N_9274,N_8952,N_8954);
or U9275 (N_9275,N_8874,N_8712);
and U9276 (N_9276,N_8937,N_8820);
nand U9277 (N_9277,N_8793,N_8769);
or U9278 (N_9278,N_8939,N_8874);
nand U9279 (N_9279,N_8964,N_8991);
or U9280 (N_9280,N_8706,N_8923);
nor U9281 (N_9281,N_8813,N_8958);
or U9282 (N_9282,N_8937,N_8877);
xor U9283 (N_9283,N_8781,N_8971);
nor U9284 (N_9284,N_8765,N_8994);
and U9285 (N_9285,N_8902,N_8752);
and U9286 (N_9286,N_8710,N_8889);
nand U9287 (N_9287,N_8946,N_8735);
nor U9288 (N_9288,N_8961,N_8945);
nand U9289 (N_9289,N_8904,N_8984);
and U9290 (N_9290,N_8741,N_8987);
nand U9291 (N_9291,N_8905,N_8901);
and U9292 (N_9292,N_8780,N_8880);
xnor U9293 (N_9293,N_8942,N_8716);
and U9294 (N_9294,N_8743,N_8960);
and U9295 (N_9295,N_8778,N_8909);
or U9296 (N_9296,N_8891,N_8724);
nand U9297 (N_9297,N_8737,N_8821);
nand U9298 (N_9298,N_8846,N_8774);
and U9299 (N_9299,N_8991,N_8742);
nor U9300 (N_9300,N_9286,N_9077);
xnor U9301 (N_9301,N_9215,N_9064);
nand U9302 (N_9302,N_9070,N_9166);
nor U9303 (N_9303,N_9183,N_9116);
nand U9304 (N_9304,N_9225,N_9269);
and U9305 (N_9305,N_9181,N_9178);
or U9306 (N_9306,N_9283,N_9232);
nor U9307 (N_9307,N_9069,N_9289);
or U9308 (N_9308,N_9271,N_9090);
nor U9309 (N_9309,N_9270,N_9009);
nor U9310 (N_9310,N_9012,N_9109);
nor U9311 (N_9311,N_9204,N_9282);
nand U9312 (N_9312,N_9210,N_9035);
xnor U9313 (N_9313,N_9057,N_9044);
nand U9314 (N_9314,N_9056,N_9139);
nand U9315 (N_9315,N_9160,N_9081);
nor U9316 (N_9316,N_9261,N_9117);
or U9317 (N_9317,N_9138,N_9144);
nand U9318 (N_9318,N_9120,N_9074);
or U9319 (N_9319,N_9112,N_9260);
nor U9320 (N_9320,N_9280,N_9172);
or U9321 (N_9321,N_9072,N_9294);
and U9322 (N_9322,N_9218,N_9195);
or U9323 (N_9323,N_9060,N_9005);
or U9324 (N_9324,N_9121,N_9251);
xnor U9325 (N_9325,N_9094,N_9292);
nor U9326 (N_9326,N_9023,N_9141);
nand U9327 (N_9327,N_9084,N_9017);
nand U9328 (N_9328,N_9149,N_9290);
and U9329 (N_9329,N_9004,N_9246);
or U9330 (N_9330,N_9046,N_9273);
and U9331 (N_9331,N_9257,N_9266);
nand U9332 (N_9332,N_9182,N_9051);
or U9333 (N_9333,N_9102,N_9100);
and U9334 (N_9334,N_9157,N_9095);
or U9335 (N_9335,N_9099,N_9132);
xnor U9336 (N_9336,N_9186,N_9253);
nand U9337 (N_9337,N_9002,N_9192);
and U9338 (N_9338,N_9152,N_9043);
or U9339 (N_9339,N_9163,N_9140);
and U9340 (N_9340,N_9103,N_9089);
xor U9341 (N_9341,N_9206,N_9168);
nand U9342 (N_9342,N_9025,N_9231);
xor U9343 (N_9343,N_9174,N_9092);
nand U9344 (N_9344,N_9086,N_9021);
or U9345 (N_9345,N_9156,N_9104);
and U9346 (N_9346,N_9297,N_9027);
nand U9347 (N_9347,N_9287,N_9202);
or U9348 (N_9348,N_9101,N_9063);
or U9349 (N_9349,N_9284,N_9265);
nor U9350 (N_9350,N_9019,N_9001);
and U9351 (N_9351,N_9032,N_9125);
nor U9352 (N_9352,N_9217,N_9123);
or U9353 (N_9353,N_9224,N_9212);
or U9354 (N_9354,N_9041,N_9244);
xor U9355 (N_9355,N_9039,N_9226);
nand U9356 (N_9356,N_9298,N_9184);
nand U9357 (N_9357,N_9016,N_9259);
nor U9358 (N_9358,N_9096,N_9110);
nor U9359 (N_9359,N_9071,N_9201);
nand U9360 (N_9360,N_9198,N_9010);
nand U9361 (N_9361,N_9158,N_9208);
nand U9362 (N_9362,N_9136,N_9119);
or U9363 (N_9363,N_9254,N_9033);
and U9364 (N_9364,N_9008,N_9238);
and U9365 (N_9365,N_9180,N_9024);
nor U9366 (N_9366,N_9219,N_9170);
nand U9367 (N_9367,N_9030,N_9250);
nor U9368 (N_9368,N_9278,N_9179);
xnor U9369 (N_9369,N_9291,N_9142);
and U9370 (N_9370,N_9239,N_9194);
and U9371 (N_9371,N_9240,N_9167);
or U9372 (N_9372,N_9088,N_9153);
xor U9373 (N_9373,N_9113,N_9122);
nor U9374 (N_9374,N_9093,N_9052);
and U9375 (N_9375,N_9078,N_9288);
xor U9376 (N_9376,N_9247,N_9196);
nand U9377 (N_9377,N_9227,N_9191);
nor U9378 (N_9378,N_9159,N_9143);
and U9379 (N_9379,N_9193,N_9176);
nand U9380 (N_9380,N_9135,N_9020);
and U9381 (N_9381,N_9091,N_9105);
and U9382 (N_9382,N_9299,N_9130);
and U9383 (N_9383,N_9114,N_9209);
xor U9384 (N_9384,N_9173,N_9047);
xor U9385 (N_9385,N_9131,N_9028);
xor U9386 (N_9386,N_9235,N_9067);
xnor U9387 (N_9387,N_9128,N_9042);
or U9388 (N_9388,N_9048,N_9248);
or U9389 (N_9389,N_9211,N_9061);
nor U9390 (N_9390,N_9222,N_9034);
or U9391 (N_9391,N_9189,N_9029);
nor U9392 (N_9392,N_9296,N_9097);
nand U9393 (N_9393,N_9169,N_9245);
xor U9394 (N_9394,N_9111,N_9221);
or U9395 (N_9395,N_9080,N_9126);
xnor U9396 (N_9396,N_9068,N_9236);
or U9397 (N_9397,N_9188,N_9082);
and U9398 (N_9398,N_9038,N_9161);
xnor U9399 (N_9399,N_9274,N_9106);
or U9400 (N_9400,N_9147,N_9098);
or U9401 (N_9401,N_9264,N_9268);
or U9402 (N_9402,N_9045,N_9079);
nor U9403 (N_9403,N_9285,N_9205);
nand U9404 (N_9404,N_9148,N_9199);
xor U9405 (N_9405,N_9256,N_9137);
and U9406 (N_9406,N_9272,N_9151);
nor U9407 (N_9407,N_9065,N_9175);
or U9408 (N_9408,N_9076,N_9243);
and U9409 (N_9409,N_9000,N_9073);
or U9410 (N_9410,N_9293,N_9133);
or U9411 (N_9411,N_9150,N_9177);
or U9412 (N_9412,N_9200,N_9127);
nand U9413 (N_9413,N_9164,N_9059);
nor U9414 (N_9414,N_9262,N_9134);
or U9415 (N_9415,N_9162,N_9154);
or U9416 (N_9416,N_9187,N_9066);
and U9417 (N_9417,N_9075,N_9049);
nand U9418 (N_9418,N_9234,N_9129);
nor U9419 (N_9419,N_9015,N_9108);
nor U9420 (N_9420,N_9267,N_9022);
nand U9421 (N_9421,N_9083,N_9255);
xor U9422 (N_9422,N_9054,N_9007);
or U9423 (N_9423,N_9155,N_9295);
or U9424 (N_9424,N_9146,N_9279);
xor U9425 (N_9425,N_9118,N_9115);
nand U9426 (N_9426,N_9145,N_9036);
nand U9427 (N_9427,N_9124,N_9228);
and U9428 (N_9428,N_9275,N_9190);
xor U9429 (N_9429,N_9214,N_9087);
nor U9430 (N_9430,N_9062,N_9252);
nand U9431 (N_9431,N_9230,N_9249);
nand U9432 (N_9432,N_9011,N_9223);
nand U9433 (N_9433,N_9220,N_9207);
nor U9434 (N_9434,N_9003,N_9058);
nor U9435 (N_9435,N_9031,N_9263);
nor U9436 (N_9436,N_9050,N_9277);
or U9437 (N_9437,N_9006,N_9107);
and U9438 (N_9438,N_9013,N_9026);
and U9439 (N_9439,N_9037,N_9165);
and U9440 (N_9440,N_9242,N_9014);
and U9441 (N_9441,N_9055,N_9040);
xor U9442 (N_9442,N_9185,N_9258);
nand U9443 (N_9443,N_9197,N_9085);
xor U9444 (N_9444,N_9229,N_9171);
or U9445 (N_9445,N_9233,N_9213);
nor U9446 (N_9446,N_9237,N_9018);
nor U9447 (N_9447,N_9053,N_9241);
xnor U9448 (N_9448,N_9281,N_9203);
xnor U9449 (N_9449,N_9276,N_9216);
nor U9450 (N_9450,N_9232,N_9049);
xor U9451 (N_9451,N_9215,N_9143);
nand U9452 (N_9452,N_9068,N_9160);
and U9453 (N_9453,N_9174,N_9031);
xor U9454 (N_9454,N_9095,N_9114);
xor U9455 (N_9455,N_9267,N_9259);
nand U9456 (N_9456,N_9225,N_9274);
or U9457 (N_9457,N_9165,N_9298);
or U9458 (N_9458,N_9039,N_9250);
and U9459 (N_9459,N_9165,N_9250);
xor U9460 (N_9460,N_9024,N_9158);
xor U9461 (N_9461,N_9270,N_9259);
nor U9462 (N_9462,N_9184,N_9241);
and U9463 (N_9463,N_9157,N_9190);
or U9464 (N_9464,N_9079,N_9247);
or U9465 (N_9465,N_9030,N_9285);
or U9466 (N_9466,N_9113,N_9252);
nor U9467 (N_9467,N_9226,N_9284);
and U9468 (N_9468,N_9214,N_9118);
nand U9469 (N_9469,N_9043,N_9134);
and U9470 (N_9470,N_9270,N_9119);
or U9471 (N_9471,N_9229,N_9255);
and U9472 (N_9472,N_9106,N_9116);
or U9473 (N_9473,N_9018,N_9145);
or U9474 (N_9474,N_9004,N_9115);
or U9475 (N_9475,N_9170,N_9083);
xnor U9476 (N_9476,N_9002,N_9050);
xor U9477 (N_9477,N_9132,N_9225);
nor U9478 (N_9478,N_9013,N_9102);
nand U9479 (N_9479,N_9153,N_9253);
and U9480 (N_9480,N_9063,N_9185);
nor U9481 (N_9481,N_9024,N_9080);
and U9482 (N_9482,N_9239,N_9034);
or U9483 (N_9483,N_9202,N_9219);
and U9484 (N_9484,N_9002,N_9158);
and U9485 (N_9485,N_9043,N_9205);
and U9486 (N_9486,N_9110,N_9014);
nor U9487 (N_9487,N_9132,N_9291);
nor U9488 (N_9488,N_9043,N_9229);
or U9489 (N_9489,N_9103,N_9144);
or U9490 (N_9490,N_9025,N_9032);
nand U9491 (N_9491,N_9237,N_9251);
or U9492 (N_9492,N_9105,N_9266);
xor U9493 (N_9493,N_9283,N_9264);
nor U9494 (N_9494,N_9125,N_9129);
and U9495 (N_9495,N_9143,N_9029);
xnor U9496 (N_9496,N_9201,N_9245);
and U9497 (N_9497,N_9179,N_9068);
xor U9498 (N_9498,N_9199,N_9076);
nor U9499 (N_9499,N_9150,N_9270);
xnor U9500 (N_9500,N_9234,N_9028);
xor U9501 (N_9501,N_9093,N_9291);
and U9502 (N_9502,N_9140,N_9276);
nand U9503 (N_9503,N_9207,N_9016);
and U9504 (N_9504,N_9081,N_9112);
and U9505 (N_9505,N_9101,N_9241);
xor U9506 (N_9506,N_9255,N_9181);
nor U9507 (N_9507,N_9005,N_9011);
and U9508 (N_9508,N_9192,N_9262);
or U9509 (N_9509,N_9214,N_9180);
and U9510 (N_9510,N_9053,N_9281);
or U9511 (N_9511,N_9162,N_9231);
nor U9512 (N_9512,N_9216,N_9050);
nor U9513 (N_9513,N_9094,N_9139);
xnor U9514 (N_9514,N_9252,N_9022);
or U9515 (N_9515,N_9136,N_9010);
nand U9516 (N_9516,N_9104,N_9123);
or U9517 (N_9517,N_9073,N_9289);
nand U9518 (N_9518,N_9111,N_9286);
xor U9519 (N_9519,N_9061,N_9009);
xnor U9520 (N_9520,N_9212,N_9246);
nor U9521 (N_9521,N_9259,N_9024);
nor U9522 (N_9522,N_9160,N_9097);
nor U9523 (N_9523,N_9277,N_9048);
and U9524 (N_9524,N_9092,N_9080);
xor U9525 (N_9525,N_9080,N_9012);
nand U9526 (N_9526,N_9264,N_9191);
nand U9527 (N_9527,N_9147,N_9141);
and U9528 (N_9528,N_9199,N_9112);
xor U9529 (N_9529,N_9022,N_9221);
or U9530 (N_9530,N_9171,N_9262);
xnor U9531 (N_9531,N_9239,N_9024);
nand U9532 (N_9532,N_9238,N_9024);
nand U9533 (N_9533,N_9048,N_9085);
xnor U9534 (N_9534,N_9131,N_9158);
xor U9535 (N_9535,N_9059,N_9267);
and U9536 (N_9536,N_9064,N_9166);
nand U9537 (N_9537,N_9284,N_9257);
nand U9538 (N_9538,N_9178,N_9280);
xor U9539 (N_9539,N_9003,N_9271);
or U9540 (N_9540,N_9016,N_9007);
or U9541 (N_9541,N_9184,N_9105);
nor U9542 (N_9542,N_9278,N_9158);
and U9543 (N_9543,N_9129,N_9093);
xor U9544 (N_9544,N_9142,N_9194);
and U9545 (N_9545,N_9055,N_9269);
xnor U9546 (N_9546,N_9148,N_9012);
xnor U9547 (N_9547,N_9159,N_9144);
nand U9548 (N_9548,N_9216,N_9042);
xor U9549 (N_9549,N_9035,N_9283);
nand U9550 (N_9550,N_9070,N_9122);
xnor U9551 (N_9551,N_9119,N_9123);
nand U9552 (N_9552,N_9209,N_9264);
and U9553 (N_9553,N_9049,N_9219);
nor U9554 (N_9554,N_9013,N_9129);
and U9555 (N_9555,N_9081,N_9146);
or U9556 (N_9556,N_9044,N_9193);
nand U9557 (N_9557,N_9174,N_9246);
nand U9558 (N_9558,N_9079,N_9017);
or U9559 (N_9559,N_9296,N_9271);
xor U9560 (N_9560,N_9290,N_9224);
nor U9561 (N_9561,N_9062,N_9297);
or U9562 (N_9562,N_9294,N_9132);
and U9563 (N_9563,N_9273,N_9259);
xor U9564 (N_9564,N_9273,N_9097);
and U9565 (N_9565,N_9291,N_9278);
nor U9566 (N_9566,N_9108,N_9214);
nor U9567 (N_9567,N_9046,N_9017);
and U9568 (N_9568,N_9231,N_9131);
and U9569 (N_9569,N_9162,N_9145);
xor U9570 (N_9570,N_9071,N_9127);
nor U9571 (N_9571,N_9171,N_9092);
and U9572 (N_9572,N_9174,N_9164);
or U9573 (N_9573,N_9184,N_9257);
nand U9574 (N_9574,N_9031,N_9264);
nor U9575 (N_9575,N_9175,N_9246);
and U9576 (N_9576,N_9154,N_9098);
xor U9577 (N_9577,N_9163,N_9166);
nor U9578 (N_9578,N_9018,N_9094);
xnor U9579 (N_9579,N_9136,N_9191);
or U9580 (N_9580,N_9195,N_9258);
nor U9581 (N_9581,N_9110,N_9129);
nand U9582 (N_9582,N_9096,N_9099);
nor U9583 (N_9583,N_9214,N_9159);
xnor U9584 (N_9584,N_9103,N_9234);
and U9585 (N_9585,N_9298,N_9213);
xnor U9586 (N_9586,N_9033,N_9259);
or U9587 (N_9587,N_9205,N_9200);
xnor U9588 (N_9588,N_9198,N_9050);
nand U9589 (N_9589,N_9245,N_9284);
or U9590 (N_9590,N_9168,N_9090);
or U9591 (N_9591,N_9137,N_9121);
or U9592 (N_9592,N_9189,N_9156);
xor U9593 (N_9593,N_9169,N_9099);
nor U9594 (N_9594,N_9035,N_9183);
nand U9595 (N_9595,N_9142,N_9038);
or U9596 (N_9596,N_9157,N_9155);
nor U9597 (N_9597,N_9136,N_9153);
and U9598 (N_9598,N_9187,N_9168);
nor U9599 (N_9599,N_9029,N_9021);
xor U9600 (N_9600,N_9559,N_9549);
or U9601 (N_9601,N_9435,N_9486);
xnor U9602 (N_9602,N_9517,N_9510);
and U9603 (N_9603,N_9531,N_9467);
xor U9604 (N_9604,N_9375,N_9525);
nand U9605 (N_9605,N_9381,N_9518);
nor U9606 (N_9606,N_9479,N_9499);
or U9607 (N_9607,N_9573,N_9300);
or U9608 (N_9608,N_9461,N_9474);
or U9609 (N_9609,N_9352,N_9506);
nor U9610 (N_9610,N_9521,N_9459);
or U9611 (N_9611,N_9338,N_9555);
xnor U9612 (N_9612,N_9571,N_9445);
nor U9613 (N_9613,N_9313,N_9356);
and U9614 (N_9614,N_9504,N_9449);
or U9615 (N_9615,N_9568,N_9582);
xnor U9616 (N_9616,N_9359,N_9316);
and U9617 (N_9617,N_9505,N_9481);
or U9618 (N_9618,N_9351,N_9304);
xnor U9619 (N_9619,N_9419,N_9306);
nand U9620 (N_9620,N_9524,N_9401);
or U9621 (N_9621,N_9452,N_9410);
or U9622 (N_9622,N_9578,N_9430);
xor U9623 (N_9623,N_9412,N_9466);
xor U9624 (N_9624,N_9345,N_9454);
xor U9625 (N_9625,N_9404,N_9364);
and U9626 (N_9626,N_9408,N_9339);
xor U9627 (N_9627,N_9317,N_9436);
nand U9628 (N_9628,N_9538,N_9589);
nand U9629 (N_9629,N_9355,N_9353);
or U9630 (N_9630,N_9534,N_9315);
xnor U9631 (N_9631,N_9455,N_9354);
nor U9632 (N_9632,N_9584,N_9453);
xor U9633 (N_9633,N_9565,N_9309);
xnor U9634 (N_9634,N_9580,N_9411);
nor U9635 (N_9635,N_9484,N_9558);
and U9636 (N_9636,N_9554,N_9488);
nand U9637 (N_9637,N_9368,N_9407);
nor U9638 (N_9638,N_9437,N_9386);
nand U9639 (N_9639,N_9475,N_9468);
or U9640 (N_9640,N_9331,N_9358);
xnor U9641 (N_9641,N_9507,N_9539);
or U9642 (N_9642,N_9397,N_9402);
nand U9643 (N_9643,N_9428,N_9492);
nand U9644 (N_9644,N_9370,N_9464);
or U9645 (N_9645,N_9463,N_9372);
nand U9646 (N_9646,N_9320,N_9363);
and U9647 (N_9647,N_9596,N_9348);
or U9648 (N_9648,N_9442,N_9482);
or U9649 (N_9649,N_9498,N_9491);
or U9650 (N_9650,N_9540,N_9593);
nor U9651 (N_9651,N_9567,N_9414);
and U9652 (N_9652,N_9350,N_9537);
or U9653 (N_9653,N_9590,N_9421);
and U9654 (N_9654,N_9599,N_9462);
and U9655 (N_9655,N_9377,N_9399);
nor U9656 (N_9656,N_9497,N_9328);
nand U9657 (N_9657,N_9438,N_9325);
nor U9658 (N_9658,N_9519,N_9418);
or U9659 (N_9659,N_9321,N_9529);
xnor U9660 (N_9660,N_9423,N_9542);
or U9661 (N_9661,N_9457,N_9420);
or U9662 (N_9662,N_9406,N_9574);
nor U9663 (N_9663,N_9324,N_9380);
xnor U9664 (N_9664,N_9456,N_9310);
xnor U9665 (N_9665,N_9367,N_9340);
xor U9666 (N_9666,N_9560,N_9583);
or U9667 (N_9667,N_9302,N_9523);
and U9668 (N_9668,N_9308,N_9458);
and U9669 (N_9669,N_9569,N_9556);
or U9670 (N_9670,N_9417,N_9485);
and U9671 (N_9671,N_9480,N_9342);
or U9672 (N_9672,N_9303,N_9477);
xor U9673 (N_9673,N_9346,N_9581);
nor U9674 (N_9674,N_9541,N_9373);
or U9675 (N_9675,N_9398,N_9545);
or U9676 (N_9676,N_9566,N_9512);
or U9677 (N_9677,N_9326,N_9471);
or U9678 (N_9678,N_9347,N_9576);
nand U9679 (N_9679,N_9337,N_9476);
xor U9680 (N_9680,N_9444,N_9335);
or U9681 (N_9681,N_9385,N_9330);
and U9682 (N_9682,N_9334,N_9514);
nand U9683 (N_9683,N_9392,N_9557);
nand U9684 (N_9684,N_9450,N_9509);
nor U9685 (N_9685,N_9371,N_9516);
or U9686 (N_9686,N_9594,N_9305);
xor U9687 (N_9687,N_9333,N_9429);
or U9688 (N_9688,N_9301,N_9446);
and U9689 (N_9689,N_9469,N_9434);
nand U9690 (N_9690,N_9487,N_9522);
or U9691 (N_9691,N_9447,N_9595);
nor U9692 (N_9692,N_9562,N_9588);
nand U9693 (N_9693,N_9426,N_9473);
nand U9694 (N_9694,N_9443,N_9493);
nor U9695 (N_9695,N_9451,N_9388);
nand U9696 (N_9696,N_9563,N_9470);
nor U9697 (N_9697,N_9403,N_9378);
xnor U9698 (N_9698,N_9585,N_9513);
nor U9699 (N_9699,N_9322,N_9472);
and U9700 (N_9700,N_9441,N_9547);
and U9701 (N_9701,N_9478,N_9495);
and U9702 (N_9702,N_9366,N_9400);
and U9703 (N_9703,N_9344,N_9508);
and U9704 (N_9704,N_9391,N_9527);
xnor U9705 (N_9705,N_9553,N_9361);
or U9706 (N_9706,N_9327,N_9496);
and U9707 (N_9707,N_9369,N_9307);
xnor U9708 (N_9708,N_9544,N_9416);
or U9709 (N_9709,N_9376,N_9405);
nand U9710 (N_9710,N_9393,N_9439);
and U9711 (N_9711,N_9501,N_9389);
xor U9712 (N_9712,N_9341,N_9343);
and U9713 (N_9713,N_9586,N_9379);
xor U9714 (N_9714,N_9536,N_9413);
xor U9715 (N_9715,N_9548,N_9490);
or U9716 (N_9716,N_9329,N_9424);
and U9717 (N_9717,N_9591,N_9311);
nor U9718 (N_9718,N_9415,N_9323);
nand U9719 (N_9719,N_9579,N_9374);
or U9720 (N_9720,N_9395,N_9460);
or U9721 (N_9721,N_9382,N_9448);
xnor U9722 (N_9722,N_9390,N_9530);
xnor U9723 (N_9723,N_9465,N_9592);
and U9724 (N_9724,N_9365,N_9483);
nand U9725 (N_9725,N_9432,N_9387);
nand U9726 (N_9726,N_9561,N_9520);
and U9727 (N_9727,N_9500,N_9362);
nand U9728 (N_9728,N_9577,N_9551);
or U9729 (N_9729,N_9564,N_9427);
or U9730 (N_9730,N_9336,N_9394);
or U9731 (N_9731,N_9312,N_9433);
xor U9732 (N_9732,N_9528,N_9384);
nand U9733 (N_9733,N_9332,N_9526);
nor U9734 (N_9734,N_9535,N_9409);
nand U9735 (N_9735,N_9587,N_9572);
nor U9736 (N_9736,N_9597,N_9546);
nand U9737 (N_9737,N_9383,N_9533);
or U9738 (N_9738,N_9440,N_9314);
xor U9739 (N_9739,N_9502,N_9511);
nand U9740 (N_9740,N_9431,N_9349);
xnor U9741 (N_9741,N_9494,N_9357);
nor U9742 (N_9742,N_9318,N_9570);
nor U9743 (N_9743,N_9503,N_9532);
and U9744 (N_9744,N_9319,N_9396);
nand U9745 (N_9745,N_9422,N_9552);
and U9746 (N_9746,N_9550,N_9360);
or U9747 (N_9747,N_9515,N_9543);
nor U9748 (N_9748,N_9598,N_9489);
or U9749 (N_9749,N_9575,N_9425);
xor U9750 (N_9750,N_9343,N_9460);
and U9751 (N_9751,N_9458,N_9340);
xor U9752 (N_9752,N_9591,N_9561);
and U9753 (N_9753,N_9499,N_9576);
nor U9754 (N_9754,N_9419,N_9470);
nand U9755 (N_9755,N_9486,N_9428);
nand U9756 (N_9756,N_9447,N_9534);
nor U9757 (N_9757,N_9487,N_9593);
or U9758 (N_9758,N_9593,N_9477);
xnor U9759 (N_9759,N_9560,N_9439);
nand U9760 (N_9760,N_9575,N_9473);
and U9761 (N_9761,N_9307,N_9453);
xnor U9762 (N_9762,N_9513,N_9427);
xnor U9763 (N_9763,N_9304,N_9416);
xnor U9764 (N_9764,N_9565,N_9485);
or U9765 (N_9765,N_9510,N_9528);
or U9766 (N_9766,N_9503,N_9571);
nor U9767 (N_9767,N_9501,N_9356);
xnor U9768 (N_9768,N_9353,N_9567);
or U9769 (N_9769,N_9489,N_9338);
and U9770 (N_9770,N_9428,N_9515);
and U9771 (N_9771,N_9316,N_9393);
nand U9772 (N_9772,N_9502,N_9429);
and U9773 (N_9773,N_9529,N_9403);
and U9774 (N_9774,N_9385,N_9313);
nor U9775 (N_9775,N_9557,N_9408);
nor U9776 (N_9776,N_9534,N_9375);
nor U9777 (N_9777,N_9515,N_9400);
or U9778 (N_9778,N_9322,N_9434);
nor U9779 (N_9779,N_9580,N_9501);
and U9780 (N_9780,N_9428,N_9440);
xnor U9781 (N_9781,N_9321,N_9547);
nor U9782 (N_9782,N_9539,N_9542);
nor U9783 (N_9783,N_9334,N_9419);
and U9784 (N_9784,N_9477,N_9355);
nand U9785 (N_9785,N_9384,N_9479);
nand U9786 (N_9786,N_9532,N_9544);
nor U9787 (N_9787,N_9552,N_9318);
and U9788 (N_9788,N_9431,N_9336);
nor U9789 (N_9789,N_9597,N_9439);
and U9790 (N_9790,N_9539,N_9317);
nand U9791 (N_9791,N_9492,N_9514);
and U9792 (N_9792,N_9509,N_9533);
and U9793 (N_9793,N_9386,N_9480);
nand U9794 (N_9794,N_9403,N_9497);
and U9795 (N_9795,N_9478,N_9514);
xnor U9796 (N_9796,N_9303,N_9511);
or U9797 (N_9797,N_9532,N_9380);
nand U9798 (N_9798,N_9492,N_9487);
or U9799 (N_9799,N_9437,N_9466);
nand U9800 (N_9800,N_9353,N_9422);
xor U9801 (N_9801,N_9317,N_9441);
nor U9802 (N_9802,N_9381,N_9355);
and U9803 (N_9803,N_9559,N_9349);
or U9804 (N_9804,N_9375,N_9454);
or U9805 (N_9805,N_9516,N_9534);
nor U9806 (N_9806,N_9333,N_9482);
nand U9807 (N_9807,N_9519,N_9499);
nor U9808 (N_9808,N_9322,N_9568);
nor U9809 (N_9809,N_9448,N_9431);
xor U9810 (N_9810,N_9441,N_9501);
and U9811 (N_9811,N_9587,N_9579);
nand U9812 (N_9812,N_9592,N_9419);
nand U9813 (N_9813,N_9322,N_9431);
or U9814 (N_9814,N_9482,N_9308);
or U9815 (N_9815,N_9464,N_9428);
or U9816 (N_9816,N_9457,N_9314);
nor U9817 (N_9817,N_9428,N_9327);
xor U9818 (N_9818,N_9445,N_9407);
or U9819 (N_9819,N_9448,N_9401);
and U9820 (N_9820,N_9582,N_9326);
and U9821 (N_9821,N_9461,N_9369);
nand U9822 (N_9822,N_9587,N_9483);
and U9823 (N_9823,N_9448,N_9527);
or U9824 (N_9824,N_9481,N_9366);
xor U9825 (N_9825,N_9350,N_9556);
or U9826 (N_9826,N_9300,N_9533);
xnor U9827 (N_9827,N_9330,N_9594);
or U9828 (N_9828,N_9518,N_9368);
nor U9829 (N_9829,N_9472,N_9378);
nor U9830 (N_9830,N_9320,N_9369);
nand U9831 (N_9831,N_9405,N_9366);
nor U9832 (N_9832,N_9352,N_9573);
nor U9833 (N_9833,N_9303,N_9342);
and U9834 (N_9834,N_9550,N_9310);
nor U9835 (N_9835,N_9302,N_9578);
nor U9836 (N_9836,N_9461,N_9386);
nand U9837 (N_9837,N_9569,N_9403);
xnor U9838 (N_9838,N_9532,N_9586);
xnor U9839 (N_9839,N_9376,N_9509);
or U9840 (N_9840,N_9563,N_9386);
nand U9841 (N_9841,N_9469,N_9304);
and U9842 (N_9842,N_9512,N_9563);
and U9843 (N_9843,N_9416,N_9316);
xor U9844 (N_9844,N_9464,N_9480);
nor U9845 (N_9845,N_9571,N_9424);
nand U9846 (N_9846,N_9542,N_9348);
xnor U9847 (N_9847,N_9376,N_9514);
nor U9848 (N_9848,N_9421,N_9409);
nor U9849 (N_9849,N_9585,N_9503);
nor U9850 (N_9850,N_9495,N_9343);
xnor U9851 (N_9851,N_9382,N_9510);
or U9852 (N_9852,N_9499,N_9547);
and U9853 (N_9853,N_9475,N_9529);
or U9854 (N_9854,N_9436,N_9397);
nor U9855 (N_9855,N_9456,N_9304);
nand U9856 (N_9856,N_9428,N_9396);
xor U9857 (N_9857,N_9403,N_9355);
nor U9858 (N_9858,N_9513,N_9524);
nor U9859 (N_9859,N_9527,N_9586);
xor U9860 (N_9860,N_9519,N_9594);
and U9861 (N_9861,N_9563,N_9589);
nand U9862 (N_9862,N_9595,N_9317);
nand U9863 (N_9863,N_9555,N_9578);
nand U9864 (N_9864,N_9514,N_9581);
xnor U9865 (N_9865,N_9309,N_9535);
nor U9866 (N_9866,N_9318,N_9449);
nor U9867 (N_9867,N_9317,N_9582);
nor U9868 (N_9868,N_9528,N_9308);
xor U9869 (N_9869,N_9584,N_9432);
or U9870 (N_9870,N_9490,N_9373);
nand U9871 (N_9871,N_9452,N_9493);
or U9872 (N_9872,N_9433,N_9557);
nor U9873 (N_9873,N_9417,N_9528);
or U9874 (N_9874,N_9385,N_9300);
nor U9875 (N_9875,N_9453,N_9579);
xnor U9876 (N_9876,N_9321,N_9425);
nor U9877 (N_9877,N_9587,N_9404);
or U9878 (N_9878,N_9500,N_9401);
and U9879 (N_9879,N_9418,N_9599);
xnor U9880 (N_9880,N_9332,N_9387);
nand U9881 (N_9881,N_9419,N_9481);
nand U9882 (N_9882,N_9458,N_9420);
nor U9883 (N_9883,N_9574,N_9517);
nand U9884 (N_9884,N_9482,N_9454);
nand U9885 (N_9885,N_9368,N_9376);
or U9886 (N_9886,N_9460,N_9513);
xnor U9887 (N_9887,N_9435,N_9335);
and U9888 (N_9888,N_9477,N_9351);
or U9889 (N_9889,N_9411,N_9395);
xnor U9890 (N_9890,N_9304,N_9418);
or U9891 (N_9891,N_9439,N_9465);
nand U9892 (N_9892,N_9303,N_9498);
xor U9893 (N_9893,N_9348,N_9445);
nor U9894 (N_9894,N_9380,N_9426);
nand U9895 (N_9895,N_9363,N_9555);
and U9896 (N_9896,N_9335,N_9402);
and U9897 (N_9897,N_9555,N_9531);
nor U9898 (N_9898,N_9546,N_9347);
xor U9899 (N_9899,N_9331,N_9502);
or U9900 (N_9900,N_9784,N_9675);
or U9901 (N_9901,N_9621,N_9674);
nor U9902 (N_9902,N_9861,N_9803);
xor U9903 (N_9903,N_9759,N_9658);
and U9904 (N_9904,N_9827,N_9722);
or U9905 (N_9905,N_9677,N_9726);
or U9906 (N_9906,N_9643,N_9685);
nand U9907 (N_9907,N_9758,N_9737);
xor U9908 (N_9908,N_9801,N_9734);
xnor U9909 (N_9909,N_9633,N_9662);
nand U9910 (N_9910,N_9775,N_9707);
and U9911 (N_9911,N_9738,N_9661);
xor U9912 (N_9912,N_9770,N_9657);
xnor U9913 (N_9913,N_9636,N_9787);
xor U9914 (N_9914,N_9730,N_9620);
nand U9915 (N_9915,N_9741,N_9755);
and U9916 (N_9916,N_9644,N_9849);
and U9917 (N_9917,N_9890,N_9720);
nor U9918 (N_9918,N_9867,N_9795);
and U9919 (N_9919,N_9863,N_9690);
or U9920 (N_9920,N_9860,N_9842);
xnor U9921 (N_9921,N_9871,N_9857);
xor U9922 (N_9922,N_9805,N_9696);
or U9923 (N_9923,N_9650,N_9873);
xnor U9924 (N_9924,N_9659,N_9774);
or U9925 (N_9925,N_9750,N_9893);
nand U9926 (N_9926,N_9879,N_9616);
nor U9927 (N_9927,N_9828,N_9664);
and U9928 (N_9928,N_9679,N_9723);
or U9929 (N_9929,N_9660,N_9671);
or U9930 (N_9930,N_9818,N_9804);
and U9931 (N_9931,N_9872,N_9712);
or U9932 (N_9932,N_9794,N_9646);
nand U9933 (N_9933,N_9825,N_9702);
or U9934 (N_9934,N_9883,N_9673);
nand U9935 (N_9935,N_9683,N_9859);
xnor U9936 (N_9936,N_9791,N_9826);
and U9937 (N_9937,N_9709,N_9779);
or U9938 (N_9938,N_9830,N_9780);
nand U9939 (N_9939,N_9713,N_9672);
nor U9940 (N_9940,N_9769,N_9700);
nand U9941 (N_9941,N_9699,N_9776);
nor U9942 (N_9942,N_9808,N_9733);
nor U9943 (N_9943,N_9751,N_9884);
or U9944 (N_9944,N_9718,N_9724);
and U9945 (N_9945,N_9687,N_9817);
xnor U9946 (N_9946,N_9831,N_9792);
and U9947 (N_9947,N_9630,N_9611);
or U9948 (N_9948,N_9823,N_9848);
nor U9949 (N_9949,N_9645,N_9868);
and U9950 (N_9950,N_9766,N_9882);
and U9951 (N_9951,N_9614,N_9815);
and U9952 (N_9952,N_9874,N_9742);
xor U9953 (N_9953,N_9889,N_9802);
nand U9954 (N_9954,N_9878,N_9880);
or U9955 (N_9955,N_9789,N_9788);
nand U9956 (N_9956,N_9866,N_9606);
and U9957 (N_9957,N_9684,N_9813);
nor U9958 (N_9958,N_9716,N_9695);
or U9959 (N_9959,N_9881,N_9745);
nor U9960 (N_9960,N_9717,N_9739);
nand U9961 (N_9961,N_9666,N_9607);
or U9962 (N_9962,N_9631,N_9894);
or U9963 (N_9963,N_9604,N_9731);
or U9964 (N_9964,N_9875,N_9809);
xor U9965 (N_9965,N_9897,N_9855);
and U9966 (N_9966,N_9782,N_9836);
and U9967 (N_9967,N_9710,N_9747);
nor U9968 (N_9968,N_9693,N_9654);
or U9969 (N_9969,N_9697,N_9752);
and U9970 (N_9970,N_9760,N_9834);
xnor U9971 (N_9971,N_9680,N_9768);
nor U9972 (N_9972,N_9870,N_9609);
or U9973 (N_9973,N_9719,N_9886);
nand U9974 (N_9974,N_9892,N_9708);
nand U9975 (N_9975,N_9885,N_9624);
nand U9976 (N_9976,N_9623,N_9856);
and U9977 (N_9977,N_9656,N_9891);
or U9978 (N_9978,N_9898,N_9667);
xor U9979 (N_9979,N_9689,N_9844);
nand U9980 (N_9980,N_9668,N_9688);
and U9981 (N_9981,N_9772,N_9835);
and U9982 (N_9982,N_9841,N_9704);
or U9983 (N_9983,N_9613,N_9816);
and U9984 (N_9984,N_9676,N_9845);
xor U9985 (N_9985,N_9729,N_9744);
xor U9986 (N_9986,N_9773,N_9698);
nand U9987 (N_9987,N_9832,N_9888);
and U9988 (N_9988,N_9852,N_9819);
and U9989 (N_9989,N_9781,N_9627);
nand U9990 (N_9990,N_9612,N_9632);
nor U9991 (N_9991,N_9833,N_9850);
and U9992 (N_9992,N_9601,N_9798);
nor U9993 (N_9993,N_9846,N_9663);
xor U9994 (N_9994,N_9896,N_9701);
or U9995 (N_9995,N_9865,N_9838);
xnor U9996 (N_9996,N_9858,N_9767);
nand U9997 (N_9997,N_9635,N_9622);
xor U9998 (N_9998,N_9869,N_9610);
and U9999 (N_9999,N_9692,N_9652);
nand U10000 (N_10000,N_9640,N_9847);
nand U10001 (N_10001,N_9619,N_9777);
nor U10002 (N_10002,N_9732,N_9761);
nand U10003 (N_10003,N_9763,N_9617);
and U10004 (N_10004,N_9853,N_9754);
nor U10005 (N_10005,N_9655,N_9820);
nor U10006 (N_10006,N_9649,N_9615);
or U10007 (N_10007,N_9669,N_9839);
and U10008 (N_10008,N_9771,N_9851);
nand U10009 (N_10009,N_9691,N_9665);
xnor U10010 (N_10010,N_9641,N_9748);
and U10011 (N_10011,N_9806,N_9715);
and U10012 (N_10012,N_9637,N_9783);
nand U10013 (N_10013,N_9786,N_9647);
and U10014 (N_10014,N_9799,N_9762);
and U10015 (N_10015,N_9682,N_9686);
xnor U10016 (N_10016,N_9837,N_9887);
xor U10017 (N_10017,N_9600,N_9814);
and U10018 (N_10018,N_9793,N_9796);
nor U10019 (N_10019,N_9822,N_9812);
xnor U10020 (N_10020,N_9678,N_9876);
nor U10021 (N_10021,N_9648,N_9602);
and U10022 (N_10022,N_9714,N_9603);
xnor U10023 (N_10023,N_9629,N_9743);
or U10024 (N_10024,N_9736,N_9810);
nand U10025 (N_10025,N_9778,N_9625);
and U10026 (N_10026,N_9811,N_9639);
xnor U10027 (N_10027,N_9728,N_9725);
nand U10028 (N_10028,N_9864,N_9829);
or U10029 (N_10029,N_9608,N_9757);
nor U10030 (N_10030,N_9605,N_9653);
or U10031 (N_10031,N_9764,N_9628);
nor U10032 (N_10032,N_9854,N_9765);
or U10033 (N_10033,N_9626,N_9749);
xnor U10034 (N_10034,N_9681,N_9727);
nand U10035 (N_10035,N_9895,N_9824);
or U10036 (N_10036,N_9899,N_9746);
and U10037 (N_10037,N_9862,N_9807);
nor U10038 (N_10038,N_9840,N_9618);
nor U10039 (N_10039,N_9740,N_9651);
xor U10040 (N_10040,N_9711,N_9721);
and U10041 (N_10041,N_9821,N_9638);
or U10042 (N_10042,N_9800,N_9756);
and U10043 (N_10043,N_9705,N_9735);
nand U10044 (N_10044,N_9843,N_9694);
and U10045 (N_10045,N_9785,N_9634);
and U10046 (N_10046,N_9642,N_9670);
or U10047 (N_10047,N_9753,N_9703);
or U10048 (N_10048,N_9706,N_9877);
nor U10049 (N_10049,N_9797,N_9790);
and U10050 (N_10050,N_9640,N_9714);
nand U10051 (N_10051,N_9630,N_9898);
and U10052 (N_10052,N_9859,N_9813);
nor U10053 (N_10053,N_9632,N_9733);
and U10054 (N_10054,N_9833,N_9607);
nor U10055 (N_10055,N_9863,N_9795);
xnor U10056 (N_10056,N_9710,N_9618);
and U10057 (N_10057,N_9610,N_9676);
nor U10058 (N_10058,N_9882,N_9845);
or U10059 (N_10059,N_9876,N_9853);
and U10060 (N_10060,N_9736,N_9680);
or U10061 (N_10061,N_9828,N_9851);
nor U10062 (N_10062,N_9677,N_9806);
nand U10063 (N_10063,N_9795,N_9673);
nand U10064 (N_10064,N_9774,N_9694);
nor U10065 (N_10065,N_9828,N_9753);
or U10066 (N_10066,N_9791,N_9885);
nand U10067 (N_10067,N_9600,N_9649);
nor U10068 (N_10068,N_9824,N_9783);
nor U10069 (N_10069,N_9864,N_9730);
xor U10070 (N_10070,N_9654,N_9721);
or U10071 (N_10071,N_9800,N_9843);
or U10072 (N_10072,N_9606,N_9832);
xor U10073 (N_10073,N_9639,N_9861);
xnor U10074 (N_10074,N_9702,N_9896);
or U10075 (N_10075,N_9699,N_9682);
and U10076 (N_10076,N_9653,N_9728);
nor U10077 (N_10077,N_9798,N_9774);
and U10078 (N_10078,N_9642,N_9652);
nor U10079 (N_10079,N_9778,N_9861);
nand U10080 (N_10080,N_9812,N_9632);
nor U10081 (N_10081,N_9715,N_9611);
nor U10082 (N_10082,N_9601,N_9742);
nor U10083 (N_10083,N_9623,N_9637);
nor U10084 (N_10084,N_9640,N_9860);
or U10085 (N_10085,N_9713,N_9626);
and U10086 (N_10086,N_9789,N_9751);
or U10087 (N_10087,N_9668,N_9876);
nor U10088 (N_10088,N_9858,N_9654);
nor U10089 (N_10089,N_9840,N_9694);
nand U10090 (N_10090,N_9740,N_9762);
and U10091 (N_10091,N_9774,N_9758);
xor U10092 (N_10092,N_9645,N_9854);
nor U10093 (N_10093,N_9661,N_9724);
and U10094 (N_10094,N_9615,N_9768);
nor U10095 (N_10095,N_9809,N_9710);
xnor U10096 (N_10096,N_9762,N_9776);
and U10097 (N_10097,N_9648,N_9719);
and U10098 (N_10098,N_9736,N_9671);
nand U10099 (N_10099,N_9612,N_9864);
nand U10100 (N_10100,N_9772,N_9776);
or U10101 (N_10101,N_9840,N_9664);
nor U10102 (N_10102,N_9891,N_9717);
xor U10103 (N_10103,N_9885,N_9851);
or U10104 (N_10104,N_9827,N_9771);
or U10105 (N_10105,N_9776,N_9774);
or U10106 (N_10106,N_9822,N_9773);
nand U10107 (N_10107,N_9815,N_9813);
and U10108 (N_10108,N_9661,N_9896);
xnor U10109 (N_10109,N_9647,N_9698);
xor U10110 (N_10110,N_9659,N_9703);
nand U10111 (N_10111,N_9695,N_9737);
nor U10112 (N_10112,N_9871,N_9658);
xor U10113 (N_10113,N_9860,N_9675);
nor U10114 (N_10114,N_9888,N_9646);
nand U10115 (N_10115,N_9613,N_9773);
nor U10116 (N_10116,N_9798,N_9789);
nor U10117 (N_10117,N_9646,N_9710);
and U10118 (N_10118,N_9648,N_9876);
and U10119 (N_10119,N_9635,N_9796);
and U10120 (N_10120,N_9753,N_9899);
nor U10121 (N_10121,N_9757,N_9862);
or U10122 (N_10122,N_9881,N_9894);
and U10123 (N_10123,N_9741,N_9896);
xor U10124 (N_10124,N_9747,N_9611);
nand U10125 (N_10125,N_9694,N_9870);
and U10126 (N_10126,N_9840,N_9739);
nor U10127 (N_10127,N_9869,N_9750);
and U10128 (N_10128,N_9687,N_9630);
or U10129 (N_10129,N_9836,N_9683);
and U10130 (N_10130,N_9714,N_9686);
nor U10131 (N_10131,N_9702,N_9809);
nor U10132 (N_10132,N_9749,N_9799);
xnor U10133 (N_10133,N_9799,N_9880);
xor U10134 (N_10134,N_9782,N_9826);
nand U10135 (N_10135,N_9829,N_9891);
xnor U10136 (N_10136,N_9651,N_9732);
nor U10137 (N_10137,N_9699,N_9619);
and U10138 (N_10138,N_9647,N_9654);
xor U10139 (N_10139,N_9732,N_9625);
nor U10140 (N_10140,N_9682,N_9781);
nor U10141 (N_10141,N_9679,N_9883);
nor U10142 (N_10142,N_9647,N_9615);
xnor U10143 (N_10143,N_9852,N_9830);
nor U10144 (N_10144,N_9723,N_9600);
or U10145 (N_10145,N_9658,N_9790);
nor U10146 (N_10146,N_9886,N_9616);
nand U10147 (N_10147,N_9756,N_9683);
nor U10148 (N_10148,N_9670,N_9683);
nor U10149 (N_10149,N_9843,N_9728);
nor U10150 (N_10150,N_9646,N_9740);
or U10151 (N_10151,N_9750,N_9600);
and U10152 (N_10152,N_9719,N_9711);
and U10153 (N_10153,N_9647,N_9878);
and U10154 (N_10154,N_9709,N_9641);
nand U10155 (N_10155,N_9678,N_9852);
and U10156 (N_10156,N_9615,N_9618);
and U10157 (N_10157,N_9787,N_9866);
and U10158 (N_10158,N_9710,N_9640);
or U10159 (N_10159,N_9617,N_9700);
and U10160 (N_10160,N_9755,N_9602);
nor U10161 (N_10161,N_9644,N_9638);
xor U10162 (N_10162,N_9777,N_9881);
and U10163 (N_10163,N_9855,N_9671);
nor U10164 (N_10164,N_9737,N_9657);
nor U10165 (N_10165,N_9638,N_9773);
nor U10166 (N_10166,N_9796,N_9624);
nand U10167 (N_10167,N_9619,N_9877);
or U10168 (N_10168,N_9867,N_9684);
nor U10169 (N_10169,N_9821,N_9825);
nor U10170 (N_10170,N_9652,N_9747);
or U10171 (N_10171,N_9715,N_9829);
nand U10172 (N_10172,N_9826,N_9836);
nor U10173 (N_10173,N_9759,N_9894);
nor U10174 (N_10174,N_9819,N_9620);
nor U10175 (N_10175,N_9745,N_9711);
xor U10176 (N_10176,N_9872,N_9676);
or U10177 (N_10177,N_9714,N_9820);
and U10178 (N_10178,N_9878,N_9683);
nor U10179 (N_10179,N_9738,N_9800);
nor U10180 (N_10180,N_9791,N_9713);
xnor U10181 (N_10181,N_9724,N_9867);
nand U10182 (N_10182,N_9656,N_9677);
nand U10183 (N_10183,N_9646,N_9667);
nor U10184 (N_10184,N_9863,N_9603);
xor U10185 (N_10185,N_9622,N_9673);
xor U10186 (N_10186,N_9668,N_9773);
or U10187 (N_10187,N_9743,N_9650);
xor U10188 (N_10188,N_9836,N_9878);
or U10189 (N_10189,N_9712,N_9647);
or U10190 (N_10190,N_9899,N_9718);
nor U10191 (N_10191,N_9610,N_9782);
nor U10192 (N_10192,N_9615,N_9670);
xor U10193 (N_10193,N_9835,N_9626);
nand U10194 (N_10194,N_9843,N_9872);
or U10195 (N_10195,N_9878,N_9633);
and U10196 (N_10196,N_9635,N_9629);
nand U10197 (N_10197,N_9740,N_9788);
xor U10198 (N_10198,N_9769,N_9794);
and U10199 (N_10199,N_9752,N_9684);
nor U10200 (N_10200,N_9962,N_10088);
and U10201 (N_10201,N_9909,N_10184);
or U10202 (N_10202,N_9934,N_10045);
xnor U10203 (N_10203,N_10108,N_10195);
nor U10204 (N_10204,N_9963,N_10020);
xnor U10205 (N_10205,N_9967,N_9924);
xnor U10206 (N_10206,N_9933,N_10018);
or U10207 (N_10207,N_10077,N_10130);
nand U10208 (N_10208,N_10192,N_10090);
nor U10209 (N_10209,N_10132,N_9911);
or U10210 (N_10210,N_9970,N_9942);
nand U10211 (N_10211,N_9913,N_10063);
xnor U10212 (N_10212,N_10099,N_10006);
xnor U10213 (N_10213,N_10129,N_10101);
nand U10214 (N_10214,N_9938,N_10084);
nor U10215 (N_10215,N_10120,N_10128);
or U10216 (N_10216,N_10068,N_9925);
nand U10217 (N_10217,N_9984,N_10143);
or U10218 (N_10218,N_10150,N_10087);
or U10219 (N_10219,N_10017,N_10049);
nor U10220 (N_10220,N_9990,N_10030);
nor U10221 (N_10221,N_10188,N_10034);
and U10222 (N_10222,N_10069,N_10076);
nor U10223 (N_10223,N_9906,N_10151);
nor U10224 (N_10224,N_10021,N_9921);
nand U10225 (N_10225,N_10080,N_10111);
or U10226 (N_10226,N_10031,N_10038);
nor U10227 (N_10227,N_10062,N_10089);
nand U10228 (N_10228,N_10092,N_10053);
nor U10229 (N_10229,N_10160,N_10023);
nand U10230 (N_10230,N_10078,N_10010);
or U10231 (N_10231,N_10060,N_10033);
xor U10232 (N_10232,N_10012,N_9964);
xor U10233 (N_10233,N_9972,N_10171);
and U10234 (N_10234,N_10015,N_10165);
or U10235 (N_10235,N_10114,N_9959);
nor U10236 (N_10236,N_10048,N_9904);
nor U10237 (N_10237,N_10110,N_10113);
nor U10238 (N_10238,N_10106,N_9987);
xor U10239 (N_10239,N_10029,N_10152);
and U10240 (N_10240,N_10169,N_10140);
xnor U10241 (N_10241,N_10144,N_10066);
xor U10242 (N_10242,N_9993,N_10139);
nand U10243 (N_10243,N_9928,N_9955);
nor U10244 (N_10244,N_9992,N_10162);
xnor U10245 (N_10245,N_10134,N_9902);
nor U10246 (N_10246,N_10157,N_9979);
nor U10247 (N_10247,N_9939,N_9919);
or U10248 (N_10248,N_10054,N_10124);
nor U10249 (N_10249,N_10005,N_10001);
xnor U10250 (N_10250,N_9903,N_9931);
nand U10251 (N_10251,N_10127,N_9944);
nor U10252 (N_10252,N_9985,N_10137);
nand U10253 (N_10253,N_9943,N_10047);
nor U10254 (N_10254,N_10148,N_10037);
and U10255 (N_10255,N_10187,N_9976);
nor U10256 (N_10256,N_10107,N_9941);
nor U10257 (N_10257,N_10071,N_10098);
and U10258 (N_10258,N_9956,N_9920);
nand U10259 (N_10259,N_9929,N_10198);
or U10260 (N_10260,N_10170,N_10135);
and U10261 (N_10261,N_10147,N_9936);
or U10262 (N_10262,N_9994,N_10154);
xor U10263 (N_10263,N_10167,N_9997);
nor U10264 (N_10264,N_10052,N_10178);
xnor U10265 (N_10265,N_10081,N_10191);
nand U10266 (N_10266,N_9914,N_9969);
nor U10267 (N_10267,N_10168,N_10174);
or U10268 (N_10268,N_9980,N_10011);
nand U10269 (N_10269,N_9968,N_9958);
nor U10270 (N_10270,N_9901,N_10036);
xnor U10271 (N_10271,N_9986,N_9926);
or U10272 (N_10272,N_10105,N_10014);
xnor U10273 (N_10273,N_9960,N_10093);
or U10274 (N_10274,N_10112,N_10126);
or U10275 (N_10275,N_9927,N_10156);
nor U10276 (N_10276,N_10193,N_9910);
nor U10277 (N_10277,N_10176,N_10196);
and U10278 (N_10278,N_10158,N_9991);
and U10279 (N_10279,N_10159,N_10166);
or U10280 (N_10280,N_10040,N_9988);
nor U10281 (N_10281,N_10061,N_9947);
nand U10282 (N_10282,N_10046,N_10003);
xor U10283 (N_10283,N_10185,N_10027);
nor U10284 (N_10284,N_10073,N_10032);
nor U10285 (N_10285,N_9952,N_10199);
xor U10286 (N_10286,N_10025,N_10072);
or U10287 (N_10287,N_9917,N_9954);
and U10288 (N_10288,N_10115,N_10097);
nor U10289 (N_10289,N_10022,N_9999);
and U10290 (N_10290,N_10117,N_9918);
or U10291 (N_10291,N_10104,N_9945);
xnor U10292 (N_10292,N_9923,N_10056);
nor U10293 (N_10293,N_10197,N_9957);
nor U10294 (N_10294,N_10125,N_10136);
nand U10295 (N_10295,N_10075,N_9978);
and U10296 (N_10296,N_10179,N_10059);
nor U10297 (N_10297,N_10164,N_9922);
nor U10298 (N_10298,N_9915,N_10024);
nand U10299 (N_10299,N_10064,N_10183);
xor U10300 (N_10300,N_10175,N_10067);
nand U10301 (N_10301,N_9974,N_9983);
nand U10302 (N_10302,N_10058,N_10163);
nor U10303 (N_10303,N_9982,N_9966);
and U10304 (N_10304,N_10122,N_9908);
nor U10305 (N_10305,N_10116,N_9940);
or U10306 (N_10306,N_10055,N_10103);
and U10307 (N_10307,N_10177,N_10182);
nor U10308 (N_10308,N_10041,N_9946);
nor U10309 (N_10309,N_9948,N_10035);
xor U10310 (N_10310,N_10057,N_10082);
and U10311 (N_10311,N_10086,N_10149);
nor U10312 (N_10312,N_10119,N_10118);
xnor U10313 (N_10313,N_10002,N_9950);
and U10314 (N_10314,N_9937,N_9975);
nand U10315 (N_10315,N_10096,N_10100);
and U10316 (N_10316,N_10007,N_9935);
nand U10317 (N_10317,N_10173,N_10181);
and U10318 (N_10318,N_9951,N_10095);
xnor U10319 (N_10319,N_9953,N_10094);
or U10320 (N_10320,N_10145,N_10186);
or U10321 (N_10321,N_10013,N_9973);
xor U10322 (N_10322,N_10004,N_9995);
nand U10323 (N_10323,N_10091,N_10050);
or U10324 (N_10324,N_10180,N_10043);
nor U10325 (N_10325,N_10146,N_9905);
nor U10326 (N_10326,N_10009,N_9930);
or U10327 (N_10327,N_9916,N_10123);
xor U10328 (N_10328,N_9998,N_10083);
nand U10329 (N_10329,N_9981,N_9977);
xnor U10330 (N_10330,N_10142,N_10051);
nor U10331 (N_10331,N_10016,N_10155);
nand U10332 (N_10332,N_9996,N_10102);
xnor U10333 (N_10333,N_10085,N_10028);
xor U10334 (N_10334,N_10039,N_10044);
xor U10335 (N_10335,N_10121,N_10000);
nor U10336 (N_10336,N_10161,N_9971);
or U10337 (N_10337,N_10109,N_10074);
or U10338 (N_10338,N_9949,N_10026);
or U10339 (N_10339,N_10138,N_10042);
or U10340 (N_10340,N_9932,N_9900);
nor U10341 (N_10341,N_10133,N_10019);
xor U10342 (N_10342,N_9961,N_10065);
xor U10343 (N_10343,N_10008,N_10131);
or U10344 (N_10344,N_10194,N_9965);
or U10345 (N_10345,N_10190,N_9912);
or U10346 (N_10346,N_10079,N_10141);
nand U10347 (N_10347,N_9989,N_10172);
or U10348 (N_10348,N_10189,N_10153);
nand U10349 (N_10349,N_9907,N_10070);
nor U10350 (N_10350,N_10119,N_10108);
nand U10351 (N_10351,N_10048,N_9969);
nor U10352 (N_10352,N_10103,N_10013);
and U10353 (N_10353,N_10035,N_9915);
xor U10354 (N_10354,N_10064,N_9970);
or U10355 (N_10355,N_9916,N_10053);
nand U10356 (N_10356,N_9938,N_10177);
and U10357 (N_10357,N_10001,N_10196);
xnor U10358 (N_10358,N_10047,N_9958);
nor U10359 (N_10359,N_9918,N_10061);
and U10360 (N_10360,N_10183,N_9904);
xnor U10361 (N_10361,N_9948,N_9909);
nand U10362 (N_10362,N_10117,N_10056);
or U10363 (N_10363,N_9966,N_10046);
and U10364 (N_10364,N_10044,N_10041);
or U10365 (N_10365,N_9918,N_10121);
nand U10366 (N_10366,N_10118,N_10111);
or U10367 (N_10367,N_9910,N_10042);
nand U10368 (N_10368,N_9961,N_9989);
nand U10369 (N_10369,N_10100,N_9954);
and U10370 (N_10370,N_9965,N_10108);
nand U10371 (N_10371,N_10169,N_9938);
nor U10372 (N_10372,N_10133,N_9935);
or U10373 (N_10373,N_10167,N_10148);
nand U10374 (N_10374,N_10023,N_9933);
xnor U10375 (N_10375,N_10180,N_10173);
or U10376 (N_10376,N_10133,N_10053);
and U10377 (N_10377,N_9952,N_9970);
nor U10378 (N_10378,N_10135,N_9906);
nand U10379 (N_10379,N_10072,N_9937);
xor U10380 (N_10380,N_9935,N_9968);
xor U10381 (N_10381,N_10167,N_10062);
or U10382 (N_10382,N_10059,N_9918);
or U10383 (N_10383,N_10056,N_10100);
nor U10384 (N_10384,N_10086,N_9914);
or U10385 (N_10385,N_9990,N_10136);
nor U10386 (N_10386,N_10180,N_10019);
nand U10387 (N_10387,N_9975,N_10146);
nor U10388 (N_10388,N_10035,N_10033);
nor U10389 (N_10389,N_10085,N_10128);
and U10390 (N_10390,N_9902,N_9942);
or U10391 (N_10391,N_9929,N_10147);
or U10392 (N_10392,N_10183,N_10068);
xnor U10393 (N_10393,N_9955,N_9915);
nand U10394 (N_10394,N_10105,N_10083);
nor U10395 (N_10395,N_9990,N_10134);
nor U10396 (N_10396,N_10162,N_9940);
and U10397 (N_10397,N_10154,N_10028);
or U10398 (N_10398,N_10131,N_10105);
xor U10399 (N_10399,N_9963,N_9901);
or U10400 (N_10400,N_9965,N_9923);
nor U10401 (N_10401,N_10181,N_10073);
nor U10402 (N_10402,N_9943,N_9903);
nor U10403 (N_10403,N_10139,N_9900);
nand U10404 (N_10404,N_10157,N_9959);
nor U10405 (N_10405,N_10081,N_10109);
nor U10406 (N_10406,N_10197,N_10134);
or U10407 (N_10407,N_9915,N_10009);
and U10408 (N_10408,N_10149,N_10099);
xnor U10409 (N_10409,N_9956,N_10135);
nand U10410 (N_10410,N_10096,N_10109);
nor U10411 (N_10411,N_10135,N_10104);
or U10412 (N_10412,N_10044,N_10070);
and U10413 (N_10413,N_9915,N_10196);
xnor U10414 (N_10414,N_10131,N_10180);
nor U10415 (N_10415,N_10022,N_10084);
or U10416 (N_10416,N_10110,N_10177);
nor U10417 (N_10417,N_9984,N_9956);
or U10418 (N_10418,N_9965,N_9911);
nand U10419 (N_10419,N_10150,N_10164);
nor U10420 (N_10420,N_10170,N_9991);
and U10421 (N_10421,N_10063,N_10105);
nor U10422 (N_10422,N_10065,N_10036);
nor U10423 (N_10423,N_10076,N_9909);
nor U10424 (N_10424,N_10179,N_10138);
xnor U10425 (N_10425,N_10011,N_10188);
or U10426 (N_10426,N_10090,N_10187);
nand U10427 (N_10427,N_9904,N_10000);
nor U10428 (N_10428,N_9956,N_10118);
or U10429 (N_10429,N_9961,N_9964);
nor U10430 (N_10430,N_9949,N_10143);
nor U10431 (N_10431,N_10108,N_10139);
and U10432 (N_10432,N_10144,N_10188);
nor U10433 (N_10433,N_10145,N_9903);
xnor U10434 (N_10434,N_10182,N_10122);
xor U10435 (N_10435,N_9971,N_10115);
nor U10436 (N_10436,N_10171,N_10034);
nor U10437 (N_10437,N_9929,N_10003);
and U10438 (N_10438,N_10126,N_10001);
xnor U10439 (N_10439,N_10119,N_10092);
nor U10440 (N_10440,N_10077,N_10197);
nand U10441 (N_10441,N_10186,N_9978);
or U10442 (N_10442,N_10131,N_9952);
nor U10443 (N_10443,N_10187,N_9999);
nor U10444 (N_10444,N_9971,N_9941);
xnor U10445 (N_10445,N_10029,N_10190);
nor U10446 (N_10446,N_9916,N_10115);
xor U10447 (N_10447,N_10124,N_10043);
nand U10448 (N_10448,N_10086,N_9956);
xnor U10449 (N_10449,N_10060,N_9999);
nor U10450 (N_10450,N_10147,N_9970);
nor U10451 (N_10451,N_9995,N_10097);
nand U10452 (N_10452,N_10039,N_10075);
or U10453 (N_10453,N_9973,N_10105);
nor U10454 (N_10454,N_9990,N_10148);
nand U10455 (N_10455,N_9943,N_10078);
nand U10456 (N_10456,N_10090,N_10131);
xnor U10457 (N_10457,N_10179,N_10046);
and U10458 (N_10458,N_10014,N_10135);
nand U10459 (N_10459,N_10048,N_10053);
and U10460 (N_10460,N_10073,N_9957);
xnor U10461 (N_10461,N_9916,N_10126);
xnor U10462 (N_10462,N_10123,N_9918);
nand U10463 (N_10463,N_9921,N_10197);
nand U10464 (N_10464,N_9909,N_9969);
xnor U10465 (N_10465,N_9931,N_10116);
or U10466 (N_10466,N_9904,N_10139);
or U10467 (N_10467,N_10138,N_10169);
and U10468 (N_10468,N_9907,N_10164);
nor U10469 (N_10469,N_10130,N_9955);
nand U10470 (N_10470,N_9923,N_10001);
nor U10471 (N_10471,N_10030,N_9952);
nand U10472 (N_10472,N_10185,N_9908);
nand U10473 (N_10473,N_10124,N_10142);
and U10474 (N_10474,N_10133,N_9930);
nand U10475 (N_10475,N_9934,N_9952);
or U10476 (N_10476,N_9964,N_10157);
or U10477 (N_10477,N_10121,N_10008);
nand U10478 (N_10478,N_10018,N_10105);
and U10479 (N_10479,N_10157,N_10058);
nor U10480 (N_10480,N_9945,N_9921);
and U10481 (N_10481,N_10037,N_10125);
xor U10482 (N_10482,N_9993,N_9981);
and U10483 (N_10483,N_10079,N_10125);
and U10484 (N_10484,N_10142,N_9992);
or U10485 (N_10485,N_10186,N_10128);
xnor U10486 (N_10486,N_10192,N_9994);
nand U10487 (N_10487,N_10038,N_10017);
and U10488 (N_10488,N_10099,N_9901);
xnor U10489 (N_10489,N_10127,N_9961);
nor U10490 (N_10490,N_10043,N_10115);
and U10491 (N_10491,N_10010,N_10006);
xor U10492 (N_10492,N_10047,N_9997);
and U10493 (N_10493,N_10135,N_10131);
nor U10494 (N_10494,N_10149,N_10049);
or U10495 (N_10495,N_9970,N_9945);
xnor U10496 (N_10496,N_10123,N_10096);
and U10497 (N_10497,N_9971,N_9949);
and U10498 (N_10498,N_10038,N_9985);
nand U10499 (N_10499,N_10141,N_10108);
nor U10500 (N_10500,N_10283,N_10495);
or U10501 (N_10501,N_10437,N_10232);
or U10502 (N_10502,N_10366,N_10406);
nand U10503 (N_10503,N_10315,N_10256);
or U10504 (N_10504,N_10409,N_10439);
or U10505 (N_10505,N_10402,N_10261);
nor U10506 (N_10506,N_10248,N_10350);
and U10507 (N_10507,N_10246,N_10419);
and U10508 (N_10508,N_10314,N_10247);
or U10509 (N_10509,N_10210,N_10252);
nor U10510 (N_10510,N_10223,N_10368);
xnor U10511 (N_10511,N_10490,N_10454);
or U10512 (N_10512,N_10474,N_10408);
xnor U10513 (N_10513,N_10341,N_10268);
xor U10514 (N_10514,N_10317,N_10231);
or U10515 (N_10515,N_10237,N_10332);
and U10516 (N_10516,N_10357,N_10399);
nand U10517 (N_10517,N_10496,N_10438);
or U10518 (N_10518,N_10395,N_10219);
nand U10519 (N_10519,N_10420,N_10461);
nor U10520 (N_10520,N_10291,N_10220);
nor U10521 (N_10521,N_10456,N_10309);
nor U10522 (N_10522,N_10352,N_10233);
nor U10523 (N_10523,N_10325,N_10426);
nand U10524 (N_10524,N_10326,N_10388);
nor U10525 (N_10525,N_10398,N_10462);
or U10526 (N_10526,N_10303,N_10282);
nor U10527 (N_10527,N_10382,N_10413);
and U10528 (N_10528,N_10458,N_10414);
nand U10529 (N_10529,N_10227,N_10381);
nand U10530 (N_10530,N_10400,N_10370);
and U10531 (N_10531,N_10239,N_10385);
and U10532 (N_10532,N_10287,N_10344);
and U10533 (N_10533,N_10207,N_10307);
xnor U10534 (N_10534,N_10353,N_10410);
xnor U10535 (N_10535,N_10243,N_10453);
nand U10536 (N_10536,N_10355,N_10215);
or U10537 (N_10537,N_10432,N_10304);
nor U10538 (N_10538,N_10488,N_10298);
nand U10539 (N_10539,N_10440,N_10201);
nor U10540 (N_10540,N_10306,N_10205);
xnor U10541 (N_10541,N_10292,N_10258);
nor U10542 (N_10542,N_10242,N_10333);
xor U10543 (N_10543,N_10296,N_10280);
nor U10544 (N_10544,N_10305,N_10200);
nor U10545 (N_10545,N_10289,N_10202);
or U10546 (N_10546,N_10324,N_10444);
or U10547 (N_10547,N_10466,N_10312);
nor U10548 (N_10548,N_10442,N_10234);
xor U10549 (N_10549,N_10241,N_10340);
xnor U10550 (N_10550,N_10404,N_10469);
nor U10551 (N_10551,N_10269,N_10313);
xor U10552 (N_10552,N_10473,N_10389);
nor U10553 (N_10553,N_10323,N_10288);
nand U10554 (N_10554,N_10417,N_10468);
and U10555 (N_10555,N_10351,N_10491);
nand U10556 (N_10556,N_10452,N_10411);
and U10557 (N_10557,N_10475,N_10228);
and U10558 (N_10558,N_10331,N_10446);
nor U10559 (N_10559,N_10492,N_10369);
xor U10560 (N_10560,N_10266,N_10421);
nand U10561 (N_10561,N_10362,N_10273);
nand U10562 (N_10562,N_10345,N_10270);
xor U10563 (N_10563,N_10321,N_10229);
nand U10564 (N_10564,N_10257,N_10250);
xnor U10565 (N_10565,N_10396,N_10300);
or U10566 (N_10566,N_10482,N_10459);
nand U10567 (N_10567,N_10218,N_10375);
nand U10568 (N_10568,N_10271,N_10483);
xnor U10569 (N_10569,N_10486,N_10221);
nor U10570 (N_10570,N_10477,N_10240);
nand U10571 (N_10571,N_10464,N_10476);
xor U10572 (N_10572,N_10371,N_10293);
xnor U10573 (N_10573,N_10425,N_10481);
xor U10574 (N_10574,N_10278,N_10479);
xnor U10575 (N_10575,N_10367,N_10485);
and U10576 (N_10576,N_10415,N_10275);
xor U10577 (N_10577,N_10354,N_10412);
and U10578 (N_10578,N_10390,N_10214);
nand U10579 (N_10579,N_10467,N_10329);
nor U10580 (N_10580,N_10254,N_10272);
or U10581 (N_10581,N_10379,N_10360);
or U10582 (N_10582,N_10251,N_10445);
or U10583 (N_10583,N_10363,N_10392);
or U10584 (N_10584,N_10443,N_10471);
nand U10585 (N_10585,N_10397,N_10489);
or U10586 (N_10586,N_10203,N_10498);
nor U10587 (N_10587,N_10424,N_10327);
and U10588 (N_10588,N_10384,N_10224);
xor U10589 (N_10589,N_10487,N_10274);
or U10590 (N_10590,N_10322,N_10276);
xor U10591 (N_10591,N_10295,N_10418);
and U10592 (N_10592,N_10428,N_10302);
nor U10593 (N_10593,N_10290,N_10301);
nor U10594 (N_10594,N_10284,N_10431);
or U10595 (N_10595,N_10376,N_10334);
nor U10596 (N_10596,N_10441,N_10447);
or U10597 (N_10597,N_10436,N_10416);
nor U10598 (N_10598,N_10267,N_10364);
nand U10599 (N_10599,N_10222,N_10225);
xor U10600 (N_10600,N_10245,N_10338);
xor U10601 (N_10601,N_10238,N_10429);
and U10602 (N_10602,N_10457,N_10244);
nor U10603 (N_10603,N_10451,N_10497);
xnor U10604 (N_10604,N_10335,N_10455);
or U10605 (N_10605,N_10320,N_10212);
xnor U10606 (N_10606,N_10365,N_10405);
and U10607 (N_10607,N_10263,N_10356);
nand U10608 (N_10608,N_10211,N_10401);
xor U10609 (N_10609,N_10226,N_10387);
or U10610 (N_10610,N_10260,N_10294);
and U10611 (N_10611,N_10349,N_10297);
and U10612 (N_10612,N_10372,N_10430);
or U10613 (N_10613,N_10435,N_10448);
or U10614 (N_10614,N_10336,N_10374);
nor U10615 (N_10615,N_10433,N_10391);
and U10616 (N_10616,N_10262,N_10265);
and U10617 (N_10617,N_10348,N_10358);
xnor U10618 (N_10618,N_10299,N_10472);
or U10619 (N_10619,N_10434,N_10423);
or U10620 (N_10620,N_10380,N_10318);
nor U10621 (N_10621,N_10480,N_10383);
xnor U10622 (N_10622,N_10499,N_10230);
nand U10623 (N_10623,N_10264,N_10337);
or U10624 (N_10624,N_10393,N_10470);
and U10625 (N_10625,N_10449,N_10361);
and U10626 (N_10626,N_10216,N_10259);
nand U10627 (N_10627,N_10378,N_10460);
nand U10628 (N_10628,N_10281,N_10373);
nor U10629 (N_10629,N_10394,N_10494);
and U10630 (N_10630,N_10347,N_10316);
nand U10631 (N_10631,N_10463,N_10310);
nor U10632 (N_10632,N_10285,N_10213);
nor U10633 (N_10633,N_10204,N_10328);
or U10634 (N_10634,N_10255,N_10403);
xnor U10635 (N_10635,N_10279,N_10478);
and U10636 (N_10636,N_10450,N_10277);
xor U10637 (N_10637,N_10217,N_10236);
or U10638 (N_10638,N_10308,N_10339);
nand U10639 (N_10639,N_10342,N_10493);
or U10640 (N_10640,N_10319,N_10206);
or U10641 (N_10641,N_10235,N_10343);
and U10642 (N_10642,N_10209,N_10427);
or U10643 (N_10643,N_10286,N_10359);
or U10644 (N_10644,N_10407,N_10377);
and U10645 (N_10645,N_10249,N_10346);
nor U10646 (N_10646,N_10253,N_10311);
xor U10647 (N_10647,N_10386,N_10208);
xor U10648 (N_10648,N_10484,N_10422);
nand U10649 (N_10649,N_10465,N_10330);
or U10650 (N_10650,N_10402,N_10309);
and U10651 (N_10651,N_10342,N_10412);
nor U10652 (N_10652,N_10242,N_10463);
or U10653 (N_10653,N_10325,N_10241);
nor U10654 (N_10654,N_10271,N_10227);
and U10655 (N_10655,N_10390,N_10405);
nand U10656 (N_10656,N_10418,N_10238);
nor U10657 (N_10657,N_10344,N_10341);
and U10658 (N_10658,N_10372,N_10423);
or U10659 (N_10659,N_10441,N_10342);
xor U10660 (N_10660,N_10274,N_10319);
nor U10661 (N_10661,N_10427,N_10392);
or U10662 (N_10662,N_10219,N_10259);
xor U10663 (N_10663,N_10411,N_10288);
and U10664 (N_10664,N_10241,N_10392);
and U10665 (N_10665,N_10366,N_10210);
nand U10666 (N_10666,N_10430,N_10269);
and U10667 (N_10667,N_10410,N_10456);
nor U10668 (N_10668,N_10405,N_10452);
nor U10669 (N_10669,N_10218,N_10406);
or U10670 (N_10670,N_10374,N_10426);
or U10671 (N_10671,N_10226,N_10242);
and U10672 (N_10672,N_10224,N_10329);
nand U10673 (N_10673,N_10338,N_10369);
nor U10674 (N_10674,N_10352,N_10256);
nand U10675 (N_10675,N_10356,N_10334);
and U10676 (N_10676,N_10394,N_10349);
nor U10677 (N_10677,N_10454,N_10324);
nor U10678 (N_10678,N_10364,N_10424);
and U10679 (N_10679,N_10305,N_10489);
or U10680 (N_10680,N_10311,N_10258);
nand U10681 (N_10681,N_10459,N_10280);
or U10682 (N_10682,N_10349,N_10290);
or U10683 (N_10683,N_10439,N_10454);
nor U10684 (N_10684,N_10256,N_10433);
nand U10685 (N_10685,N_10332,N_10287);
or U10686 (N_10686,N_10327,N_10427);
or U10687 (N_10687,N_10451,N_10201);
or U10688 (N_10688,N_10477,N_10347);
or U10689 (N_10689,N_10299,N_10317);
nand U10690 (N_10690,N_10299,N_10297);
nor U10691 (N_10691,N_10472,N_10326);
or U10692 (N_10692,N_10265,N_10315);
or U10693 (N_10693,N_10433,N_10298);
nand U10694 (N_10694,N_10200,N_10323);
or U10695 (N_10695,N_10316,N_10214);
xor U10696 (N_10696,N_10381,N_10323);
nor U10697 (N_10697,N_10342,N_10218);
and U10698 (N_10698,N_10234,N_10402);
nor U10699 (N_10699,N_10356,N_10228);
nor U10700 (N_10700,N_10337,N_10338);
nor U10701 (N_10701,N_10466,N_10393);
nor U10702 (N_10702,N_10219,N_10315);
xnor U10703 (N_10703,N_10339,N_10454);
xor U10704 (N_10704,N_10228,N_10297);
nand U10705 (N_10705,N_10350,N_10389);
nand U10706 (N_10706,N_10438,N_10291);
or U10707 (N_10707,N_10427,N_10479);
xnor U10708 (N_10708,N_10306,N_10254);
xor U10709 (N_10709,N_10246,N_10433);
nand U10710 (N_10710,N_10220,N_10451);
nand U10711 (N_10711,N_10359,N_10229);
nand U10712 (N_10712,N_10320,N_10262);
nor U10713 (N_10713,N_10415,N_10351);
nor U10714 (N_10714,N_10407,N_10205);
nand U10715 (N_10715,N_10428,N_10219);
nand U10716 (N_10716,N_10445,N_10465);
nand U10717 (N_10717,N_10319,N_10352);
xor U10718 (N_10718,N_10388,N_10227);
nand U10719 (N_10719,N_10347,N_10496);
or U10720 (N_10720,N_10325,N_10339);
nor U10721 (N_10721,N_10290,N_10417);
nand U10722 (N_10722,N_10274,N_10286);
nor U10723 (N_10723,N_10457,N_10245);
and U10724 (N_10724,N_10327,N_10361);
xor U10725 (N_10725,N_10369,N_10404);
or U10726 (N_10726,N_10474,N_10345);
xnor U10727 (N_10727,N_10285,N_10358);
xor U10728 (N_10728,N_10291,N_10388);
and U10729 (N_10729,N_10287,N_10210);
nor U10730 (N_10730,N_10254,N_10250);
or U10731 (N_10731,N_10232,N_10486);
nand U10732 (N_10732,N_10359,N_10203);
or U10733 (N_10733,N_10314,N_10285);
or U10734 (N_10734,N_10269,N_10349);
or U10735 (N_10735,N_10271,N_10298);
nand U10736 (N_10736,N_10315,N_10399);
or U10737 (N_10737,N_10211,N_10391);
nand U10738 (N_10738,N_10243,N_10469);
or U10739 (N_10739,N_10489,N_10258);
nor U10740 (N_10740,N_10461,N_10438);
nand U10741 (N_10741,N_10454,N_10411);
or U10742 (N_10742,N_10411,N_10282);
xnor U10743 (N_10743,N_10360,N_10470);
nand U10744 (N_10744,N_10434,N_10346);
and U10745 (N_10745,N_10204,N_10337);
and U10746 (N_10746,N_10244,N_10479);
nand U10747 (N_10747,N_10290,N_10239);
and U10748 (N_10748,N_10276,N_10258);
or U10749 (N_10749,N_10295,N_10356);
nor U10750 (N_10750,N_10375,N_10431);
xnor U10751 (N_10751,N_10401,N_10312);
or U10752 (N_10752,N_10311,N_10448);
nand U10753 (N_10753,N_10379,N_10234);
and U10754 (N_10754,N_10361,N_10475);
xnor U10755 (N_10755,N_10270,N_10265);
xor U10756 (N_10756,N_10498,N_10366);
xnor U10757 (N_10757,N_10345,N_10444);
xnor U10758 (N_10758,N_10282,N_10300);
nor U10759 (N_10759,N_10226,N_10205);
and U10760 (N_10760,N_10376,N_10229);
nor U10761 (N_10761,N_10408,N_10244);
xor U10762 (N_10762,N_10304,N_10412);
or U10763 (N_10763,N_10257,N_10251);
and U10764 (N_10764,N_10287,N_10451);
nand U10765 (N_10765,N_10277,N_10231);
or U10766 (N_10766,N_10402,N_10492);
and U10767 (N_10767,N_10456,N_10273);
xor U10768 (N_10768,N_10256,N_10324);
nand U10769 (N_10769,N_10430,N_10381);
or U10770 (N_10770,N_10486,N_10283);
or U10771 (N_10771,N_10336,N_10221);
xor U10772 (N_10772,N_10354,N_10430);
and U10773 (N_10773,N_10477,N_10248);
nand U10774 (N_10774,N_10444,N_10301);
nand U10775 (N_10775,N_10385,N_10488);
and U10776 (N_10776,N_10245,N_10206);
or U10777 (N_10777,N_10341,N_10478);
nand U10778 (N_10778,N_10409,N_10378);
xor U10779 (N_10779,N_10419,N_10310);
xnor U10780 (N_10780,N_10386,N_10394);
nor U10781 (N_10781,N_10261,N_10464);
nand U10782 (N_10782,N_10314,N_10202);
nand U10783 (N_10783,N_10320,N_10217);
xor U10784 (N_10784,N_10353,N_10473);
or U10785 (N_10785,N_10359,N_10450);
and U10786 (N_10786,N_10401,N_10405);
or U10787 (N_10787,N_10420,N_10439);
xnor U10788 (N_10788,N_10438,N_10231);
nor U10789 (N_10789,N_10368,N_10398);
xnor U10790 (N_10790,N_10229,N_10353);
nor U10791 (N_10791,N_10238,N_10405);
or U10792 (N_10792,N_10311,N_10340);
xnor U10793 (N_10793,N_10216,N_10372);
xor U10794 (N_10794,N_10291,N_10422);
nand U10795 (N_10795,N_10327,N_10204);
xnor U10796 (N_10796,N_10355,N_10352);
xor U10797 (N_10797,N_10481,N_10373);
nor U10798 (N_10798,N_10494,N_10387);
nand U10799 (N_10799,N_10222,N_10452);
nor U10800 (N_10800,N_10638,N_10764);
xnor U10801 (N_10801,N_10711,N_10729);
nor U10802 (N_10802,N_10613,N_10581);
nand U10803 (N_10803,N_10626,N_10589);
xnor U10804 (N_10804,N_10639,N_10798);
nor U10805 (N_10805,N_10701,N_10509);
nand U10806 (N_10806,N_10650,N_10541);
nand U10807 (N_10807,N_10681,N_10607);
or U10808 (N_10808,N_10679,N_10722);
nor U10809 (N_10809,N_10591,N_10765);
nor U10810 (N_10810,N_10732,N_10597);
or U10811 (N_10811,N_10572,N_10715);
and U10812 (N_10812,N_10636,N_10538);
nor U10813 (N_10813,N_10696,N_10789);
or U10814 (N_10814,N_10657,N_10579);
and U10815 (N_10815,N_10551,N_10601);
or U10816 (N_10816,N_10616,N_10698);
or U10817 (N_10817,N_10796,N_10521);
xor U10818 (N_10818,N_10506,N_10659);
xnor U10819 (N_10819,N_10625,N_10645);
nand U10820 (N_10820,N_10554,N_10710);
nor U10821 (N_10821,N_10767,N_10622);
nor U10822 (N_10822,N_10550,N_10629);
or U10823 (N_10823,N_10564,N_10654);
xor U10824 (N_10824,N_10708,N_10669);
nand U10825 (N_10825,N_10682,N_10713);
and U10826 (N_10826,N_10632,N_10548);
and U10827 (N_10827,N_10678,N_10686);
nor U10828 (N_10828,N_10621,N_10615);
xor U10829 (N_10829,N_10664,N_10536);
nor U10830 (N_10830,N_10772,N_10658);
nor U10831 (N_10831,N_10515,N_10552);
xnor U10832 (N_10832,N_10748,N_10555);
and U10833 (N_10833,N_10504,N_10533);
and U10834 (N_10834,N_10699,N_10665);
nand U10835 (N_10835,N_10736,N_10777);
or U10836 (N_10836,N_10633,N_10714);
or U10837 (N_10837,N_10751,N_10797);
and U10838 (N_10838,N_10584,N_10576);
nand U10839 (N_10839,N_10680,N_10582);
nand U10840 (N_10840,N_10532,N_10624);
or U10841 (N_10841,N_10676,N_10531);
nand U10842 (N_10842,N_10547,N_10518);
xor U10843 (N_10843,N_10525,N_10718);
or U10844 (N_10844,N_10743,N_10562);
and U10845 (N_10845,N_10724,N_10642);
and U10846 (N_10846,N_10760,N_10725);
nand U10847 (N_10847,N_10747,N_10731);
or U10848 (N_10848,N_10691,N_10675);
nand U10849 (N_10849,N_10684,N_10575);
or U10850 (N_10850,N_10662,N_10566);
nand U10851 (N_10851,N_10542,N_10598);
xnor U10852 (N_10852,N_10539,N_10794);
or U10853 (N_10853,N_10644,N_10631);
nor U10854 (N_10854,N_10513,N_10526);
nand U10855 (N_10855,N_10685,N_10611);
xor U10856 (N_10856,N_10688,N_10744);
xnor U10857 (N_10857,N_10619,N_10653);
or U10858 (N_10858,N_10578,N_10635);
and U10859 (N_10859,N_10740,N_10630);
nand U10860 (N_10860,N_10719,N_10690);
xnor U10861 (N_10861,N_10637,N_10648);
nor U10862 (N_10862,N_10553,N_10647);
xnor U10863 (N_10863,N_10683,N_10565);
xnor U10864 (N_10864,N_10706,N_10671);
nor U10865 (N_10865,N_10754,N_10573);
nor U10866 (N_10866,N_10757,N_10508);
nor U10867 (N_10867,N_10500,N_10605);
xnor U10868 (N_10868,N_10783,N_10762);
nor U10869 (N_10869,N_10778,N_10721);
and U10870 (N_10870,N_10663,N_10733);
xor U10871 (N_10871,N_10535,N_10528);
xor U10872 (N_10872,N_10559,N_10694);
nand U10873 (N_10873,N_10689,N_10609);
or U10874 (N_10874,N_10560,N_10503);
or U10875 (N_10875,N_10524,N_10599);
nor U10876 (N_10876,N_10695,N_10792);
or U10877 (N_10877,N_10540,N_10668);
and U10878 (N_10878,N_10771,N_10571);
xnor U10879 (N_10879,N_10577,N_10716);
and U10880 (N_10880,N_10614,N_10612);
xnor U10881 (N_10881,N_10738,N_10580);
xor U10882 (N_10882,N_10501,N_10784);
xnor U10883 (N_10883,N_10769,N_10750);
nand U10884 (N_10884,N_10779,N_10793);
nor U10885 (N_10885,N_10723,N_10652);
and U10886 (N_10886,N_10594,N_10569);
nor U10887 (N_10887,N_10693,N_10752);
xor U10888 (N_10888,N_10727,N_10561);
nand U10889 (N_10889,N_10546,N_10790);
or U10890 (N_10890,N_10737,N_10726);
xnor U10891 (N_10891,N_10585,N_10623);
nor U10892 (N_10892,N_10795,N_10505);
and U10893 (N_10893,N_10590,N_10558);
and U10894 (N_10894,N_10742,N_10735);
xor U10895 (N_10895,N_10655,N_10507);
or U10896 (N_10896,N_10527,N_10774);
xnor U10897 (N_10897,N_10730,N_10502);
nor U10898 (N_10898,N_10746,N_10570);
and U10899 (N_10899,N_10717,N_10606);
xor U10900 (N_10900,N_10745,N_10557);
or U10901 (N_10901,N_10586,N_10641);
nor U10902 (N_10902,N_10620,N_10768);
nor U10903 (N_10903,N_10643,N_10704);
xnor U10904 (N_10904,N_10781,N_10608);
nor U10905 (N_10905,N_10567,N_10734);
and U10906 (N_10906,N_10692,N_10697);
nor U10907 (N_10907,N_10511,N_10780);
nor U10908 (N_10908,N_10674,N_10703);
nand U10909 (N_10909,N_10753,N_10687);
nor U10910 (N_10910,N_10770,N_10728);
nand U10911 (N_10911,N_10785,N_10593);
xnor U10912 (N_10912,N_10596,N_10755);
or U10913 (N_10913,N_10523,N_10628);
and U10914 (N_10914,N_10782,N_10574);
and U10915 (N_10915,N_10617,N_10700);
nor U10916 (N_10916,N_10766,N_10707);
and U10917 (N_10917,N_10512,N_10775);
and U10918 (N_10918,N_10763,N_10530);
nor U10919 (N_10919,N_10670,N_10739);
and U10920 (N_10920,N_10634,N_10741);
or U10921 (N_10921,N_10517,N_10712);
xnor U10922 (N_10922,N_10514,N_10758);
nor U10923 (N_10923,N_10543,N_10588);
nor U10924 (N_10924,N_10661,N_10651);
nor U10925 (N_10925,N_10602,N_10660);
and U10926 (N_10926,N_10720,N_10672);
and U10927 (N_10927,N_10510,N_10595);
or U10928 (N_10928,N_10537,N_10583);
xor U10929 (N_10929,N_10759,N_10756);
nor U10930 (N_10930,N_10556,N_10786);
nand U10931 (N_10931,N_10519,N_10568);
xor U10932 (N_10932,N_10603,N_10749);
nor U10933 (N_10933,N_10544,N_10761);
or U10934 (N_10934,N_10618,N_10627);
or U10935 (N_10935,N_10705,N_10667);
or U10936 (N_10936,N_10520,N_10549);
and U10937 (N_10937,N_10646,N_10773);
xor U10938 (N_10938,N_10677,N_10791);
nor U10939 (N_10939,N_10788,N_10534);
nor U10940 (N_10940,N_10563,N_10529);
xor U10941 (N_10941,N_10640,N_10522);
and U10942 (N_10942,N_10610,N_10587);
or U10943 (N_10943,N_10799,N_10545);
and U10944 (N_10944,N_10649,N_10600);
nor U10945 (N_10945,N_10666,N_10516);
nand U10946 (N_10946,N_10709,N_10604);
nor U10947 (N_10947,N_10787,N_10702);
and U10948 (N_10948,N_10656,N_10592);
nor U10949 (N_10949,N_10673,N_10776);
xnor U10950 (N_10950,N_10646,N_10584);
and U10951 (N_10951,N_10616,N_10786);
xor U10952 (N_10952,N_10734,N_10508);
xnor U10953 (N_10953,N_10619,N_10550);
nor U10954 (N_10954,N_10676,N_10553);
or U10955 (N_10955,N_10790,N_10618);
and U10956 (N_10956,N_10570,N_10634);
xor U10957 (N_10957,N_10601,N_10759);
xor U10958 (N_10958,N_10799,N_10726);
nand U10959 (N_10959,N_10737,N_10531);
nand U10960 (N_10960,N_10705,N_10790);
or U10961 (N_10961,N_10749,N_10755);
nand U10962 (N_10962,N_10542,N_10618);
and U10963 (N_10963,N_10508,N_10738);
and U10964 (N_10964,N_10784,N_10704);
nor U10965 (N_10965,N_10513,N_10598);
and U10966 (N_10966,N_10517,N_10683);
nand U10967 (N_10967,N_10748,N_10764);
nand U10968 (N_10968,N_10503,N_10535);
xnor U10969 (N_10969,N_10560,N_10519);
or U10970 (N_10970,N_10715,N_10738);
and U10971 (N_10971,N_10640,N_10703);
xnor U10972 (N_10972,N_10569,N_10564);
nor U10973 (N_10973,N_10544,N_10670);
or U10974 (N_10974,N_10721,N_10658);
or U10975 (N_10975,N_10742,N_10508);
nor U10976 (N_10976,N_10783,N_10791);
or U10977 (N_10977,N_10762,N_10639);
or U10978 (N_10978,N_10753,N_10764);
or U10979 (N_10979,N_10751,N_10790);
or U10980 (N_10980,N_10619,N_10567);
xnor U10981 (N_10981,N_10626,N_10728);
xor U10982 (N_10982,N_10722,N_10760);
nand U10983 (N_10983,N_10749,N_10744);
nand U10984 (N_10984,N_10584,N_10667);
nand U10985 (N_10985,N_10767,N_10707);
nand U10986 (N_10986,N_10644,N_10581);
and U10987 (N_10987,N_10647,N_10752);
xor U10988 (N_10988,N_10719,N_10642);
nand U10989 (N_10989,N_10580,N_10610);
nor U10990 (N_10990,N_10526,N_10542);
xnor U10991 (N_10991,N_10504,N_10651);
or U10992 (N_10992,N_10768,N_10512);
or U10993 (N_10993,N_10686,N_10512);
nand U10994 (N_10994,N_10565,N_10590);
and U10995 (N_10995,N_10562,N_10718);
nand U10996 (N_10996,N_10557,N_10572);
and U10997 (N_10997,N_10579,N_10540);
xor U10998 (N_10998,N_10799,N_10665);
xor U10999 (N_10999,N_10715,N_10671);
and U11000 (N_11000,N_10736,N_10786);
nand U11001 (N_11001,N_10697,N_10766);
and U11002 (N_11002,N_10663,N_10615);
nor U11003 (N_11003,N_10795,N_10756);
xor U11004 (N_11004,N_10603,N_10771);
or U11005 (N_11005,N_10580,N_10636);
or U11006 (N_11006,N_10501,N_10610);
and U11007 (N_11007,N_10686,N_10500);
and U11008 (N_11008,N_10625,N_10562);
nand U11009 (N_11009,N_10550,N_10728);
nand U11010 (N_11010,N_10643,N_10507);
nor U11011 (N_11011,N_10538,N_10539);
nand U11012 (N_11012,N_10743,N_10571);
xor U11013 (N_11013,N_10649,N_10565);
xor U11014 (N_11014,N_10742,N_10658);
or U11015 (N_11015,N_10675,N_10596);
xnor U11016 (N_11016,N_10798,N_10727);
or U11017 (N_11017,N_10696,N_10763);
nor U11018 (N_11018,N_10704,N_10515);
or U11019 (N_11019,N_10529,N_10791);
nand U11020 (N_11020,N_10515,N_10669);
or U11021 (N_11021,N_10606,N_10691);
xor U11022 (N_11022,N_10524,N_10759);
or U11023 (N_11023,N_10688,N_10592);
nor U11024 (N_11024,N_10535,N_10674);
or U11025 (N_11025,N_10691,N_10750);
or U11026 (N_11026,N_10518,N_10773);
or U11027 (N_11027,N_10504,N_10634);
or U11028 (N_11028,N_10590,N_10638);
xnor U11029 (N_11029,N_10742,N_10669);
nand U11030 (N_11030,N_10558,N_10577);
xor U11031 (N_11031,N_10652,N_10799);
and U11032 (N_11032,N_10597,N_10734);
or U11033 (N_11033,N_10603,N_10701);
nand U11034 (N_11034,N_10608,N_10634);
xor U11035 (N_11035,N_10677,N_10649);
or U11036 (N_11036,N_10557,N_10789);
nand U11037 (N_11037,N_10758,N_10750);
nor U11038 (N_11038,N_10762,N_10509);
nand U11039 (N_11039,N_10716,N_10644);
xnor U11040 (N_11040,N_10614,N_10587);
or U11041 (N_11041,N_10689,N_10524);
nand U11042 (N_11042,N_10522,N_10586);
nand U11043 (N_11043,N_10724,N_10605);
or U11044 (N_11044,N_10718,N_10734);
or U11045 (N_11045,N_10593,N_10641);
or U11046 (N_11046,N_10559,N_10712);
and U11047 (N_11047,N_10524,N_10540);
nand U11048 (N_11048,N_10690,N_10736);
or U11049 (N_11049,N_10707,N_10697);
nor U11050 (N_11050,N_10666,N_10508);
and U11051 (N_11051,N_10604,N_10631);
nand U11052 (N_11052,N_10544,N_10595);
and U11053 (N_11053,N_10728,N_10531);
xnor U11054 (N_11054,N_10551,N_10681);
nand U11055 (N_11055,N_10551,N_10782);
and U11056 (N_11056,N_10593,N_10649);
and U11057 (N_11057,N_10564,N_10656);
and U11058 (N_11058,N_10704,N_10577);
or U11059 (N_11059,N_10755,N_10675);
or U11060 (N_11060,N_10541,N_10759);
nand U11061 (N_11061,N_10578,N_10514);
xor U11062 (N_11062,N_10631,N_10503);
nor U11063 (N_11063,N_10757,N_10510);
or U11064 (N_11064,N_10745,N_10520);
or U11065 (N_11065,N_10774,N_10775);
xnor U11066 (N_11066,N_10775,N_10651);
or U11067 (N_11067,N_10637,N_10548);
nor U11068 (N_11068,N_10525,N_10532);
and U11069 (N_11069,N_10756,N_10783);
and U11070 (N_11070,N_10635,N_10642);
nand U11071 (N_11071,N_10682,N_10650);
and U11072 (N_11072,N_10785,N_10770);
or U11073 (N_11073,N_10741,N_10700);
nor U11074 (N_11074,N_10767,N_10615);
nand U11075 (N_11075,N_10632,N_10789);
nand U11076 (N_11076,N_10628,N_10771);
xnor U11077 (N_11077,N_10692,N_10667);
xor U11078 (N_11078,N_10637,N_10703);
and U11079 (N_11079,N_10758,N_10751);
nor U11080 (N_11080,N_10713,N_10522);
nand U11081 (N_11081,N_10739,N_10611);
nand U11082 (N_11082,N_10668,N_10655);
nand U11083 (N_11083,N_10568,N_10508);
nand U11084 (N_11084,N_10580,N_10581);
xnor U11085 (N_11085,N_10738,N_10643);
or U11086 (N_11086,N_10593,N_10768);
nor U11087 (N_11087,N_10601,N_10663);
xnor U11088 (N_11088,N_10588,N_10511);
xor U11089 (N_11089,N_10528,N_10720);
and U11090 (N_11090,N_10670,N_10606);
or U11091 (N_11091,N_10781,N_10742);
or U11092 (N_11092,N_10569,N_10528);
nor U11093 (N_11093,N_10731,N_10703);
and U11094 (N_11094,N_10769,N_10505);
xor U11095 (N_11095,N_10602,N_10753);
or U11096 (N_11096,N_10555,N_10529);
xor U11097 (N_11097,N_10704,N_10520);
nor U11098 (N_11098,N_10533,N_10717);
or U11099 (N_11099,N_10726,N_10592);
and U11100 (N_11100,N_11032,N_10984);
nand U11101 (N_11101,N_11006,N_10894);
and U11102 (N_11102,N_11094,N_11075);
or U11103 (N_11103,N_11027,N_10864);
or U11104 (N_11104,N_11051,N_11034);
nand U11105 (N_11105,N_10877,N_10952);
nand U11106 (N_11106,N_10902,N_10897);
nand U11107 (N_11107,N_10932,N_11039);
nor U11108 (N_11108,N_10987,N_11057);
or U11109 (N_11109,N_10971,N_10816);
or U11110 (N_11110,N_10921,N_10994);
and U11111 (N_11111,N_11055,N_11058);
and U11112 (N_11112,N_11007,N_10918);
and U11113 (N_11113,N_10859,N_10800);
and U11114 (N_11114,N_11059,N_11091);
or U11115 (N_11115,N_11013,N_10972);
xnor U11116 (N_11116,N_10953,N_10978);
nor U11117 (N_11117,N_11000,N_11012);
or U11118 (N_11118,N_10882,N_11070);
and U11119 (N_11119,N_10834,N_10819);
or U11120 (N_11120,N_10803,N_10881);
or U11121 (N_11121,N_10958,N_10880);
nor U11122 (N_11122,N_11081,N_10846);
nor U11123 (N_11123,N_11066,N_10874);
nor U11124 (N_11124,N_11011,N_10906);
or U11125 (N_11125,N_10948,N_11024);
and U11126 (N_11126,N_11088,N_10910);
nand U11127 (N_11127,N_11092,N_10837);
nand U11128 (N_11128,N_10830,N_11043);
and U11129 (N_11129,N_10946,N_10878);
nand U11130 (N_11130,N_10991,N_11082);
and U11131 (N_11131,N_10852,N_10916);
and U11132 (N_11132,N_10925,N_10802);
and U11133 (N_11133,N_11080,N_10839);
or U11134 (N_11134,N_10934,N_10960);
xor U11135 (N_11135,N_10854,N_10823);
xor U11136 (N_11136,N_10895,N_10967);
nand U11137 (N_11137,N_10840,N_10871);
xnor U11138 (N_11138,N_11033,N_10982);
and U11139 (N_11139,N_11040,N_10838);
xnor U11140 (N_11140,N_10810,N_11064);
xor U11141 (N_11141,N_10937,N_11009);
xor U11142 (N_11142,N_10997,N_10806);
xnor U11143 (N_11143,N_11016,N_10957);
nand U11144 (N_11144,N_10805,N_10985);
xor U11145 (N_11145,N_11093,N_10930);
nor U11146 (N_11146,N_11071,N_11085);
nor U11147 (N_11147,N_11079,N_10890);
or U11148 (N_11148,N_10924,N_10841);
and U11149 (N_11149,N_10817,N_10973);
xor U11150 (N_11150,N_10965,N_10945);
nor U11151 (N_11151,N_10913,N_10992);
nor U11152 (N_11152,N_11045,N_10980);
xnor U11153 (N_11153,N_10820,N_11077);
or U11154 (N_11154,N_10824,N_11083);
xnor U11155 (N_11155,N_10942,N_11074);
or U11156 (N_11156,N_11019,N_11004);
nor U11157 (N_11157,N_11061,N_10876);
nor U11158 (N_11158,N_11098,N_11029);
nand U11159 (N_11159,N_11008,N_10833);
or U11160 (N_11160,N_10848,N_11072);
and U11161 (N_11161,N_11044,N_10993);
or U11162 (N_11162,N_11028,N_10861);
or U11163 (N_11163,N_11048,N_10964);
or U11164 (N_11164,N_11015,N_10939);
nor U11165 (N_11165,N_11047,N_10844);
nand U11166 (N_11166,N_10917,N_10961);
and U11167 (N_11167,N_10983,N_10856);
or U11168 (N_11168,N_10832,N_10996);
and U11169 (N_11169,N_10970,N_10893);
nand U11170 (N_11170,N_10842,N_10995);
nor U11171 (N_11171,N_10979,N_11096);
nand U11172 (N_11172,N_10849,N_10908);
and U11173 (N_11173,N_10875,N_10883);
xnor U11174 (N_11174,N_10956,N_10828);
nand U11175 (N_11175,N_10821,N_10929);
nor U11176 (N_11176,N_11046,N_11017);
or U11177 (N_11177,N_10857,N_10866);
and U11178 (N_11178,N_10903,N_10969);
nand U11179 (N_11179,N_10826,N_10868);
xor U11180 (N_11180,N_10928,N_10815);
nand U11181 (N_11181,N_10990,N_11020);
and U11182 (N_11182,N_10814,N_10845);
or U11183 (N_11183,N_11089,N_10981);
xor U11184 (N_11184,N_10988,N_11026);
xnor U11185 (N_11185,N_11062,N_10954);
and U11186 (N_11186,N_10940,N_10850);
or U11187 (N_11187,N_10963,N_10922);
or U11188 (N_11188,N_10827,N_10955);
and U11189 (N_11189,N_10879,N_10872);
or U11190 (N_11190,N_10949,N_10809);
xnor U11191 (N_11191,N_10891,N_11097);
or U11192 (N_11192,N_10889,N_11095);
and U11193 (N_11193,N_10905,N_10920);
nand U11194 (N_11194,N_10843,N_10862);
xnor U11195 (N_11195,N_10836,N_10888);
and U11196 (N_11196,N_10904,N_11054);
or U11197 (N_11197,N_10898,N_11023);
nand U11198 (N_11198,N_11041,N_11035);
xnor U11199 (N_11199,N_11099,N_11002);
nand U11200 (N_11200,N_10936,N_11087);
or U11201 (N_11201,N_11069,N_10915);
nand U11202 (N_11202,N_11068,N_10977);
xor U11203 (N_11203,N_11090,N_10907);
xor U11204 (N_11204,N_10912,N_11021);
or U11205 (N_11205,N_11031,N_10813);
xnor U11206 (N_11206,N_11001,N_10974);
xnor U11207 (N_11207,N_10886,N_11076);
and U11208 (N_11208,N_10825,N_10927);
nor U11209 (N_11209,N_10919,N_11042);
nand U11210 (N_11210,N_11065,N_10976);
or U11211 (N_11211,N_10938,N_10944);
xnor U11212 (N_11212,N_10892,N_10801);
nor U11213 (N_11213,N_10887,N_11003);
nand U11214 (N_11214,N_10867,N_10818);
nor U11215 (N_11215,N_10858,N_11060);
or U11216 (N_11216,N_11014,N_10822);
xor U11217 (N_11217,N_10962,N_10926);
nand U11218 (N_11218,N_10998,N_10986);
and U11219 (N_11219,N_10851,N_11022);
and U11220 (N_11220,N_10811,N_10950);
nand U11221 (N_11221,N_10935,N_11050);
nor U11222 (N_11222,N_10873,N_10808);
and U11223 (N_11223,N_11084,N_10968);
nor U11224 (N_11224,N_10899,N_10829);
xnor U11225 (N_11225,N_10966,N_11005);
nor U11226 (N_11226,N_10911,N_11038);
and U11227 (N_11227,N_10900,N_11018);
nand U11228 (N_11228,N_11025,N_10923);
xor U11229 (N_11229,N_11063,N_10933);
nor U11230 (N_11230,N_10865,N_10853);
nor U11231 (N_11231,N_10931,N_10835);
nor U11232 (N_11232,N_10999,N_11086);
or U11233 (N_11233,N_10804,N_11036);
xnor U11234 (N_11234,N_10884,N_10812);
nand U11235 (N_11235,N_11067,N_10951);
nand U11236 (N_11236,N_11052,N_10914);
or U11237 (N_11237,N_11010,N_10885);
and U11238 (N_11238,N_10807,N_10847);
or U11239 (N_11239,N_11078,N_10860);
or U11240 (N_11240,N_10947,N_10855);
xor U11241 (N_11241,N_11037,N_10975);
nor U11242 (N_11242,N_10941,N_10869);
nor U11243 (N_11243,N_10870,N_10896);
and U11244 (N_11244,N_11073,N_11056);
or U11245 (N_11245,N_11030,N_10909);
xor U11246 (N_11246,N_11053,N_10943);
or U11247 (N_11247,N_11049,N_10831);
xor U11248 (N_11248,N_10901,N_10863);
or U11249 (N_11249,N_10989,N_10959);
nor U11250 (N_11250,N_11039,N_11068);
nor U11251 (N_11251,N_10954,N_10999);
xor U11252 (N_11252,N_10964,N_10800);
xnor U11253 (N_11253,N_10910,N_10868);
nor U11254 (N_11254,N_10921,N_10811);
xor U11255 (N_11255,N_10912,N_10996);
and U11256 (N_11256,N_10917,N_10835);
nand U11257 (N_11257,N_10815,N_10997);
or U11258 (N_11258,N_10888,N_10926);
and U11259 (N_11259,N_10884,N_10801);
nand U11260 (N_11260,N_11082,N_10808);
xnor U11261 (N_11261,N_10959,N_10914);
nor U11262 (N_11262,N_11052,N_10897);
nand U11263 (N_11263,N_11088,N_11010);
and U11264 (N_11264,N_10949,N_10846);
nand U11265 (N_11265,N_11047,N_11005);
nand U11266 (N_11266,N_11006,N_11059);
and U11267 (N_11267,N_10819,N_11066);
or U11268 (N_11268,N_10953,N_10996);
and U11269 (N_11269,N_10920,N_10953);
or U11270 (N_11270,N_11010,N_10946);
nand U11271 (N_11271,N_10895,N_10801);
or U11272 (N_11272,N_11004,N_10944);
and U11273 (N_11273,N_11074,N_11035);
and U11274 (N_11274,N_11056,N_10909);
xnor U11275 (N_11275,N_10899,N_10977);
xor U11276 (N_11276,N_11073,N_10846);
nand U11277 (N_11277,N_10848,N_10928);
xor U11278 (N_11278,N_11099,N_10929);
xnor U11279 (N_11279,N_10931,N_10836);
or U11280 (N_11280,N_10979,N_10821);
and U11281 (N_11281,N_10819,N_10883);
and U11282 (N_11282,N_10883,N_10822);
xnor U11283 (N_11283,N_10899,N_10803);
and U11284 (N_11284,N_10844,N_10914);
and U11285 (N_11285,N_10866,N_10985);
or U11286 (N_11286,N_11083,N_11078);
nor U11287 (N_11287,N_10844,N_11084);
nand U11288 (N_11288,N_10933,N_11079);
and U11289 (N_11289,N_11075,N_11085);
nor U11290 (N_11290,N_10882,N_11008);
and U11291 (N_11291,N_11022,N_11085);
xnor U11292 (N_11292,N_10839,N_10885);
and U11293 (N_11293,N_11070,N_11055);
xor U11294 (N_11294,N_10843,N_10808);
nand U11295 (N_11295,N_10997,N_10891);
and U11296 (N_11296,N_11006,N_11087);
or U11297 (N_11297,N_11000,N_10957);
and U11298 (N_11298,N_10808,N_11036);
or U11299 (N_11299,N_11009,N_10945);
xor U11300 (N_11300,N_10887,N_10895);
and U11301 (N_11301,N_10954,N_10995);
or U11302 (N_11302,N_10912,N_10935);
or U11303 (N_11303,N_10814,N_11030);
nand U11304 (N_11304,N_10806,N_10864);
and U11305 (N_11305,N_10936,N_10935);
or U11306 (N_11306,N_10863,N_10837);
nor U11307 (N_11307,N_11049,N_11075);
xnor U11308 (N_11308,N_10971,N_10914);
or U11309 (N_11309,N_10876,N_10829);
nor U11310 (N_11310,N_10887,N_10983);
nand U11311 (N_11311,N_11076,N_11050);
or U11312 (N_11312,N_11035,N_10812);
and U11313 (N_11313,N_10823,N_10803);
nor U11314 (N_11314,N_11024,N_10827);
or U11315 (N_11315,N_10815,N_11022);
xnor U11316 (N_11316,N_10909,N_11021);
and U11317 (N_11317,N_11044,N_10860);
nand U11318 (N_11318,N_10955,N_11042);
and U11319 (N_11319,N_10832,N_10849);
xor U11320 (N_11320,N_11094,N_11015);
and U11321 (N_11321,N_10978,N_11077);
nand U11322 (N_11322,N_10913,N_10850);
or U11323 (N_11323,N_10809,N_11035);
nand U11324 (N_11324,N_10905,N_11074);
xnor U11325 (N_11325,N_10977,N_10863);
nand U11326 (N_11326,N_10855,N_10944);
xnor U11327 (N_11327,N_10855,N_10960);
or U11328 (N_11328,N_10984,N_10868);
xnor U11329 (N_11329,N_10954,N_10894);
nor U11330 (N_11330,N_10977,N_11048);
nand U11331 (N_11331,N_10884,N_11052);
nand U11332 (N_11332,N_10902,N_10924);
and U11333 (N_11333,N_11054,N_11097);
nor U11334 (N_11334,N_11028,N_10804);
and U11335 (N_11335,N_10986,N_10800);
and U11336 (N_11336,N_11034,N_11040);
nand U11337 (N_11337,N_10822,N_11058);
nor U11338 (N_11338,N_11067,N_10837);
or U11339 (N_11339,N_10880,N_11001);
xnor U11340 (N_11340,N_11015,N_11064);
xor U11341 (N_11341,N_10800,N_10831);
nand U11342 (N_11342,N_10988,N_10979);
nand U11343 (N_11343,N_11044,N_10845);
xor U11344 (N_11344,N_10978,N_10813);
nand U11345 (N_11345,N_10918,N_10804);
and U11346 (N_11346,N_11015,N_10816);
or U11347 (N_11347,N_10832,N_10926);
nor U11348 (N_11348,N_10936,N_10863);
and U11349 (N_11349,N_10976,N_10870);
or U11350 (N_11350,N_10934,N_10989);
and U11351 (N_11351,N_10953,N_10884);
and U11352 (N_11352,N_10898,N_11007);
or U11353 (N_11353,N_10990,N_10873);
xor U11354 (N_11354,N_10868,N_10985);
nor U11355 (N_11355,N_10852,N_11023);
nand U11356 (N_11356,N_10957,N_10838);
nor U11357 (N_11357,N_10824,N_11087);
and U11358 (N_11358,N_10814,N_11068);
or U11359 (N_11359,N_10852,N_10860);
xor U11360 (N_11360,N_10911,N_11035);
nor U11361 (N_11361,N_11055,N_11007);
nand U11362 (N_11362,N_10988,N_11005);
or U11363 (N_11363,N_10880,N_10944);
xor U11364 (N_11364,N_10975,N_11071);
xor U11365 (N_11365,N_11092,N_11070);
nor U11366 (N_11366,N_10943,N_11066);
or U11367 (N_11367,N_10913,N_10902);
xor U11368 (N_11368,N_10803,N_10956);
xnor U11369 (N_11369,N_11090,N_11036);
nor U11370 (N_11370,N_10927,N_11072);
xnor U11371 (N_11371,N_11063,N_10985);
and U11372 (N_11372,N_11013,N_11071);
nand U11373 (N_11373,N_10890,N_10920);
nor U11374 (N_11374,N_11001,N_10847);
or U11375 (N_11375,N_10919,N_10853);
or U11376 (N_11376,N_10804,N_11009);
nand U11377 (N_11377,N_11057,N_10832);
xor U11378 (N_11378,N_11045,N_11029);
nand U11379 (N_11379,N_10873,N_10968);
xor U11380 (N_11380,N_10942,N_10886);
nor U11381 (N_11381,N_11072,N_10923);
xor U11382 (N_11382,N_10975,N_11017);
xor U11383 (N_11383,N_10811,N_10869);
nor U11384 (N_11384,N_11058,N_10900);
xor U11385 (N_11385,N_11077,N_10824);
nand U11386 (N_11386,N_10808,N_10917);
or U11387 (N_11387,N_11013,N_10811);
and U11388 (N_11388,N_10921,N_10825);
nor U11389 (N_11389,N_10876,N_10961);
and U11390 (N_11390,N_11091,N_11017);
xor U11391 (N_11391,N_10839,N_10935);
nor U11392 (N_11392,N_11030,N_10981);
nand U11393 (N_11393,N_10931,N_11094);
and U11394 (N_11394,N_10802,N_10856);
nor U11395 (N_11395,N_10950,N_10951);
nor U11396 (N_11396,N_10833,N_11082);
and U11397 (N_11397,N_11005,N_11084);
nor U11398 (N_11398,N_11039,N_10980);
or U11399 (N_11399,N_10979,N_10802);
nor U11400 (N_11400,N_11223,N_11390);
or U11401 (N_11401,N_11160,N_11343);
or U11402 (N_11402,N_11161,N_11113);
or U11403 (N_11403,N_11370,N_11145);
nand U11404 (N_11404,N_11338,N_11101);
or U11405 (N_11405,N_11240,N_11248);
nor U11406 (N_11406,N_11300,N_11244);
nor U11407 (N_11407,N_11380,N_11295);
nor U11408 (N_11408,N_11126,N_11329);
or U11409 (N_11409,N_11315,N_11335);
and U11410 (N_11410,N_11368,N_11144);
nand U11411 (N_11411,N_11388,N_11189);
nor U11412 (N_11412,N_11112,N_11167);
nor U11413 (N_11413,N_11103,N_11301);
and U11414 (N_11414,N_11379,N_11376);
xnor U11415 (N_11415,N_11243,N_11196);
nor U11416 (N_11416,N_11206,N_11361);
and U11417 (N_11417,N_11362,N_11195);
nor U11418 (N_11418,N_11305,N_11227);
or U11419 (N_11419,N_11217,N_11228);
nand U11420 (N_11420,N_11247,N_11266);
nor U11421 (N_11421,N_11194,N_11313);
xor U11422 (N_11422,N_11364,N_11131);
and U11423 (N_11423,N_11245,N_11324);
or U11424 (N_11424,N_11234,N_11382);
or U11425 (N_11425,N_11287,N_11381);
nor U11426 (N_11426,N_11229,N_11304);
or U11427 (N_11427,N_11232,N_11186);
and U11428 (N_11428,N_11250,N_11256);
nor U11429 (N_11429,N_11321,N_11188);
xor U11430 (N_11430,N_11175,N_11262);
xor U11431 (N_11431,N_11200,N_11233);
or U11432 (N_11432,N_11166,N_11298);
xnor U11433 (N_11433,N_11183,N_11235);
and U11434 (N_11434,N_11385,N_11163);
nand U11435 (N_11435,N_11237,N_11303);
or U11436 (N_11436,N_11312,N_11215);
or U11437 (N_11437,N_11387,N_11174);
nor U11438 (N_11438,N_11374,N_11274);
or U11439 (N_11439,N_11273,N_11155);
nand U11440 (N_11440,N_11171,N_11164);
xnor U11441 (N_11441,N_11299,N_11213);
or U11442 (N_11442,N_11284,N_11185);
nand U11443 (N_11443,N_11261,N_11346);
and U11444 (N_11444,N_11187,N_11204);
nor U11445 (N_11445,N_11396,N_11136);
xnor U11446 (N_11446,N_11283,N_11139);
nor U11447 (N_11447,N_11292,N_11178);
nand U11448 (N_11448,N_11259,N_11358);
xor U11449 (N_11449,N_11123,N_11306);
nor U11450 (N_11450,N_11307,N_11340);
nor U11451 (N_11451,N_11350,N_11330);
nand U11452 (N_11452,N_11326,N_11116);
xor U11453 (N_11453,N_11179,N_11129);
or U11454 (N_11454,N_11115,N_11114);
nor U11455 (N_11455,N_11279,N_11354);
xnor U11456 (N_11456,N_11201,N_11149);
nand U11457 (N_11457,N_11272,N_11141);
or U11458 (N_11458,N_11276,N_11208);
or U11459 (N_11459,N_11357,N_11102);
nand U11460 (N_11460,N_11260,N_11318);
nand U11461 (N_11461,N_11207,N_11137);
or U11462 (N_11462,N_11110,N_11369);
and U11463 (N_11463,N_11107,N_11105);
xor U11464 (N_11464,N_11323,N_11290);
or U11465 (N_11465,N_11325,N_11127);
or U11466 (N_11466,N_11220,N_11359);
nand U11467 (N_11467,N_11302,N_11109);
xnor U11468 (N_11468,N_11265,N_11372);
and U11469 (N_11469,N_11333,N_11365);
nor U11470 (N_11470,N_11367,N_11199);
nor U11471 (N_11471,N_11211,N_11192);
nor U11472 (N_11472,N_11389,N_11218);
xnor U11473 (N_11473,N_11399,N_11366);
and U11474 (N_11474,N_11216,N_11239);
or U11475 (N_11475,N_11226,N_11135);
nor U11476 (N_11476,N_11236,N_11339);
nor U11477 (N_11477,N_11251,N_11269);
or U11478 (N_11478,N_11319,N_11397);
and U11479 (N_11479,N_11225,N_11386);
nor U11480 (N_11480,N_11162,N_11132);
and U11481 (N_11481,N_11373,N_11224);
xnor U11482 (N_11482,N_11184,N_11134);
and U11483 (N_11483,N_11352,N_11125);
nand U11484 (N_11484,N_11173,N_11106);
and U11485 (N_11485,N_11275,N_11331);
nor U11486 (N_11486,N_11271,N_11242);
nor U11487 (N_11487,N_11308,N_11176);
xnor U11488 (N_11488,N_11241,N_11210);
and U11489 (N_11489,N_11316,N_11293);
nand U11490 (N_11490,N_11314,N_11375);
xor U11491 (N_11491,N_11360,N_11157);
xor U11492 (N_11492,N_11311,N_11363);
nand U11493 (N_11493,N_11347,N_11336);
nor U11494 (N_11494,N_11289,N_11278);
xor U11495 (N_11495,N_11221,N_11341);
xor U11496 (N_11496,N_11356,N_11252);
and U11497 (N_11497,N_11190,N_11191);
and U11498 (N_11498,N_11180,N_11230);
nor U11499 (N_11499,N_11282,N_11142);
xnor U11500 (N_11500,N_11124,N_11197);
and U11501 (N_11501,N_11222,N_11398);
xor U11502 (N_11502,N_11263,N_11281);
and U11503 (N_11503,N_11320,N_11392);
or U11504 (N_11504,N_11296,N_11118);
nand U11505 (N_11505,N_11165,N_11146);
xor U11506 (N_11506,N_11377,N_11253);
nor U11507 (N_11507,N_11153,N_11143);
and U11508 (N_11508,N_11344,N_11159);
xor U11509 (N_11509,N_11177,N_11152);
nor U11510 (N_11510,N_11342,N_11169);
xor U11511 (N_11511,N_11255,N_11355);
and U11512 (N_11512,N_11291,N_11310);
and U11513 (N_11513,N_11257,N_11212);
nor U11514 (N_11514,N_11328,N_11268);
nor U11515 (N_11515,N_11384,N_11285);
nor U11516 (N_11516,N_11351,N_11147);
nor U11517 (N_11517,N_11383,N_11108);
nor U11518 (N_11518,N_11203,N_11202);
xnor U11519 (N_11519,N_11117,N_11294);
nor U11520 (N_11520,N_11394,N_11286);
and U11521 (N_11521,N_11317,N_11297);
nand U11522 (N_11522,N_11395,N_11121);
or U11523 (N_11523,N_11205,N_11120);
nand U11524 (N_11524,N_11104,N_11172);
and U11525 (N_11525,N_11264,N_11198);
or U11526 (N_11526,N_11182,N_11332);
nor U11527 (N_11527,N_11193,N_11214);
or U11528 (N_11528,N_11231,N_11209);
and U11529 (N_11529,N_11219,N_11334);
and U11530 (N_11530,N_11122,N_11154);
and U11531 (N_11531,N_11249,N_11270);
xnor U11532 (N_11532,N_11158,N_11378);
nand U11533 (N_11533,N_11156,N_11181);
nand U11534 (N_11534,N_11337,N_11258);
or U11535 (N_11535,N_11238,N_11111);
or U11536 (N_11536,N_11371,N_11119);
or U11537 (N_11537,N_11130,N_11267);
xnor U11538 (N_11538,N_11100,N_11288);
and U11539 (N_11539,N_11345,N_11246);
nor U11540 (N_11540,N_11150,N_11309);
or U11541 (N_11541,N_11277,N_11393);
xor U11542 (N_11542,N_11280,N_11140);
or U11543 (N_11543,N_11353,N_11348);
xor U11544 (N_11544,N_11391,N_11170);
xor U11545 (N_11545,N_11254,N_11128);
xor U11546 (N_11546,N_11138,N_11322);
or U11547 (N_11547,N_11148,N_11349);
and U11548 (N_11548,N_11327,N_11168);
or U11549 (N_11549,N_11133,N_11151);
nand U11550 (N_11550,N_11176,N_11246);
or U11551 (N_11551,N_11171,N_11251);
nor U11552 (N_11552,N_11244,N_11365);
nor U11553 (N_11553,N_11390,N_11198);
and U11554 (N_11554,N_11256,N_11367);
nand U11555 (N_11555,N_11321,N_11314);
or U11556 (N_11556,N_11333,N_11378);
nor U11557 (N_11557,N_11325,N_11293);
or U11558 (N_11558,N_11377,N_11249);
xnor U11559 (N_11559,N_11230,N_11359);
or U11560 (N_11560,N_11106,N_11245);
xor U11561 (N_11561,N_11111,N_11323);
and U11562 (N_11562,N_11355,N_11163);
and U11563 (N_11563,N_11349,N_11176);
or U11564 (N_11564,N_11266,N_11347);
and U11565 (N_11565,N_11120,N_11334);
nor U11566 (N_11566,N_11211,N_11251);
nor U11567 (N_11567,N_11198,N_11227);
nor U11568 (N_11568,N_11161,N_11309);
and U11569 (N_11569,N_11141,N_11383);
xor U11570 (N_11570,N_11270,N_11136);
and U11571 (N_11571,N_11392,N_11283);
or U11572 (N_11572,N_11191,N_11280);
nor U11573 (N_11573,N_11365,N_11378);
and U11574 (N_11574,N_11399,N_11205);
nor U11575 (N_11575,N_11157,N_11102);
or U11576 (N_11576,N_11199,N_11118);
or U11577 (N_11577,N_11200,N_11192);
xor U11578 (N_11578,N_11320,N_11339);
nor U11579 (N_11579,N_11304,N_11122);
and U11580 (N_11580,N_11304,N_11205);
nor U11581 (N_11581,N_11222,N_11283);
and U11582 (N_11582,N_11398,N_11261);
nor U11583 (N_11583,N_11356,N_11346);
or U11584 (N_11584,N_11377,N_11284);
or U11585 (N_11585,N_11293,N_11150);
or U11586 (N_11586,N_11144,N_11259);
nor U11587 (N_11587,N_11292,N_11346);
nand U11588 (N_11588,N_11217,N_11225);
or U11589 (N_11589,N_11379,N_11277);
or U11590 (N_11590,N_11231,N_11136);
nand U11591 (N_11591,N_11201,N_11127);
and U11592 (N_11592,N_11366,N_11303);
nand U11593 (N_11593,N_11280,N_11250);
and U11594 (N_11594,N_11121,N_11205);
nor U11595 (N_11595,N_11372,N_11153);
or U11596 (N_11596,N_11270,N_11301);
nand U11597 (N_11597,N_11311,N_11270);
and U11598 (N_11598,N_11335,N_11351);
and U11599 (N_11599,N_11287,N_11266);
or U11600 (N_11600,N_11301,N_11224);
and U11601 (N_11601,N_11391,N_11148);
and U11602 (N_11602,N_11365,N_11189);
nor U11603 (N_11603,N_11282,N_11292);
xnor U11604 (N_11604,N_11160,N_11341);
or U11605 (N_11605,N_11160,N_11197);
or U11606 (N_11606,N_11118,N_11121);
or U11607 (N_11607,N_11229,N_11204);
and U11608 (N_11608,N_11286,N_11106);
or U11609 (N_11609,N_11199,N_11293);
nor U11610 (N_11610,N_11367,N_11308);
and U11611 (N_11611,N_11212,N_11244);
nor U11612 (N_11612,N_11126,N_11171);
nor U11613 (N_11613,N_11209,N_11230);
or U11614 (N_11614,N_11336,N_11224);
nand U11615 (N_11615,N_11171,N_11362);
nor U11616 (N_11616,N_11164,N_11279);
xor U11617 (N_11617,N_11103,N_11199);
nand U11618 (N_11618,N_11209,N_11111);
and U11619 (N_11619,N_11267,N_11133);
and U11620 (N_11620,N_11288,N_11345);
nand U11621 (N_11621,N_11307,N_11265);
and U11622 (N_11622,N_11119,N_11351);
xor U11623 (N_11623,N_11118,N_11104);
nor U11624 (N_11624,N_11271,N_11331);
or U11625 (N_11625,N_11268,N_11245);
and U11626 (N_11626,N_11259,N_11227);
and U11627 (N_11627,N_11211,N_11254);
nor U11628 (N_11628,N_11114,N_11324);
nor U11629 (N_11629,N_11248,N_11291);
and U11630 (N_11630,N_11339,N_11310);
xor U11631 (N_11631,N_11395,N_11292);
nor U11632 (N_11632,N_11225,N_11154);
or U11633 (N_11633,N_11238,N_11380);
xor U11634 (N_11634,N_11215,N_11372);
xor U11635 (N_11635,N_11377,N_11306);
and U11636 (N_11636,N_11338,N_11158);
and U11637 (N_11637,N_11393,N_11289);
xnor U11638 (N_11638,N_11255,N_11236);
xor U11639 (N_11639,N_11107,N_11109);
nand U11640 (N_11640,N_11311,N_11151);
and U11641 (N_11641,N_11343,N_11291);
xor U11642 (N_11642,N_11346,N_11265);
xnor U11643 (N_11643,N_11376,N_11337);
nor U11644 (N_11644,N_11307,N_11287);
nor U11645 (N_11645,N_11366,N_11214);
xor U11646 (N_11646,N_11111,N_11219);
or U11647 (N_11647,N_11290,N_11398);
xor U11648 (N_11648,N_11202,N_11256);
and U11649 (N_11649,N_11318,N_11240);
and U11650 (N_11650,N_11335,N_11269);
and U11651 (N_11651,N_11322,N_11394);
nand U11652 (N_11652,N_11261,N_11275);
and U11653 (N_11653,N_11192,N_11216);
nand U11654 (N_11654,N_11273,N_11278);
or U11655 (N_11655,N_11393,N_11274);
nand U11656 (N_11656,N_11100,N_11266);
and U11657 (N_11657,N_11157,N_11114);
nand U11658 (N_11658,N_11392,N_11256);
nand U11659 (N_11659,N_11398,N_11220);
and U11660 (N_11660,N_11256,N_11237);
or U11661 (N_11661,N_11358,N_11364);
nand U11662 (N_11662,N_11111,N_11374);
nand U11663 (N_11663,N_11111,N_11366);
nand U11664 (N_11664,N_11114,N_11354);
nor U11665 (N_11665,N_11352,N_11276);
or U11666 (N_11666,N_11280,N_11256);
or U11667 (N_11667,N_11205,N_11236);
nor U11668 (N_11668,N_11300,N_11230);
and U11669 (N_11669,N_11196,N_11207);
nor U11670 (N_11670,N_11182,N_11222);
xor U11671 (N_11671,N_11343,N_11104);
nor U11672 (N_11672,N_11351,N_11155);
or U11673 (N_11673,N_11162,N_11219);
nor U11674 (N_11674,N_11168,N_11334);
nor U11675 (N_11675,N_11170,N_11354);
or U11676 (N_11676,N_11314,N_11104);
xnor U11677 (N_11677,N_11291,N_11372);
nor U11678 (N_11678,N_11255,N_11175);
and U11679 (N_11679,N_11285,N_11263);
nor U11680 (N_11680,N_11114,N_11203);
nor U11681 (N_11681,N_11362,N_11222);
xor U11682 (N_11682,N_11169,N_11334);
nor U11683 (N_11683,N_11142,N_11196);
or U11684 (N_11684,N_11318,N_11284);
xor U11685 (N_11685,N_11323,N_11221);
xor U11686 (N_11686,N_11343,N_11121);
or U11687 (N_11687,N_11301,N_11140);
nand U11688 (N_11688,N_11135,N_11301);
or U11689 (N_11689,N_11297,N_11227);
nand U11690 (N_11690,N_11322,N_11176);
xor U11691 (N_11691,N_11337,N_11102);
nand U11692 (N_11692,N_11283,N_11279);
and U11693 (N_11693,N_11266,N_11357);
nor U11694 (N_11694,N_11124,N_11121);
nor U11695 (N_11695,N_11374,N_11129);
nand U11696 (N_11696,N_11139,N_11184);
or U11697 (N_11697,N_11323,N_11225);
xnor U11698 (N_11698,N_11199,N_11331);
nand U11699 (N_11699,N_11148,N_11104);
xor U11700 (N_11700,N_11621,N_11451);
nor U11701 (N_11701,N_11671,N_11416);
nor U11702 (N_11702,N_11571,N_11646);
and U11703 (N_11703,N_11524,N_11594);
nor U11704 (N_11704,N_11670,N_11475);
nor U11705 (N_11705,N_11543,N_11401);
or U11706 (N_11706,N_11420,N_11580);
nand U11707 (N_11707,N_11688,N_11417);
and U11708 (N_11708,N_11477,N_11677);
and U11709 (N_11709,N_11648,N_11427);
xor U11710 (N_11710,N_11406,N_11601);
or U11711 (N_11711,N_11561,N_11687);
xor U11712 (N_11712,N_11668,N_11483);
and U11713 (N_11713,N_11603,N_11513);
or U11714 (N_11714,N_11560,N_11473);
xnor U11715 (N_11715,N_11622,N_11500);
nor U11716 (N_11716,N_11564,N_11482);
nand U11717 (N_11717,N_11472,N_11486);
xor U11718 (N_11718,N_11557,N_11529);
nor U11719 (N_11719,N_11534,N_11609);
and U11720 (N_11720,N_11680,N_11569);
nor U11721 (N_11721,N_11628,N_11585);
or U11722 (N_11722,N_11428,N_11515);
or U11723 (N_11723,N_11501,N_11685);
xor U11724 (N_11724,N_11471,N_11597);
and U11725 (N_11725,N_11422,N_11662);
and U11726 (N_11726,N_11689,N_11568);
nor U11727 (N_11727,N_11694,N_11492);
and U11728 (N_11728,N_11613,N_11429);
xor U11729 (N_11729,N_11699,N_11460);
nor U11730 (N_11730,N_11653,N_11425);
nand U11731 (N_11731,N_11474,N_11542);
and U11732 (N_11732,N_11638,N_11457);
and U11733 (N_11733,N_11587,N_11517);
xnor U11734 (N_11734,N_11645,N_11678);
nor U11735 (N_11735,N_11600,N_11518);
nor U11736 (N_11736,N_11658,N_11440);
xnor U11737 (N_11737,N_11665,N_11540);
nor U11738 (N_11738,N_11554,N_11562);
or U11739 (N_11739,N_11655,N_11511);
or U11740 (N_11740,N_11606,N_11552);
nand U11741 (N_11741,N_11498,N_11442);
nand U11742 (N_11742,N_11528,N_11634);
or U11743 (N_11743,N_11667,N_11488);
nand U11744 (N_11744,N_11481,N_11546);
or U11745 (N_11745,N_11445,N_11432);
nor U11746 (N_11746,N_11467,N_11647);
and U11747 (N_11747,N_11499,N_11454);
and U11748 (N_11748,N_11510,N_11676);
and U11749 (N_11749,N_11490,N_11408);
nor U11750 (N_11750,N_11559,N_11531);
xor U11751 (N_11751,N_11526,N_11436);
and U11752 (N_11752,N_11595,N_11636);
nor U11753 (N_11753,N_11404,N_11593);
nor U11754 (N_11754,N_11579,N_11468);
and U11755 (N_11755,N_11502,N_11565);
nand U11756 (N_11756,N_11405,N_11679);
nor U11757 (N_11757,N_11589,N_11489);
or U11758 (N_11758,N_11447,N_11469);
nor U11759 (N_11759,N_11617,N_11435);
nand U11760 (N_11760,N_11566,N_11459);
and U11761 (N_11761,N_11410,N_11413);
nor U11762 (N_11762,N_11553,N_11484);
nor U11763 (N_11763,N_11444,N_11683);
nor U11764 (N_11764,N_11642,N_11581);
and U11765 (N_11765,N_11627,N_11591);
nand U11766 (N_11766,N_11575,N_11519);
nor U11767 (N_11767,N_11539,N_11558);
xnor U11768 (N_11768,N_11615,N_11663);
xnor U11769 (N_11769,N_11551,N_11675);
nor U11770 (N_11770,N_11686,N_11614);
nand U11771 (N_11771,N_11437,N_11415);
or U11772 (N_11772,N_11516,N_11697);
xnor U11773 (N_11773,N_11548,N_11497);
nor U11774 (N_11774,N_11430,N_11682);
nor U11775 (N_11775,N_11637,N_11434);
and U11776 (N_11776,N_11547,N_11657);
nor U11777 (N_11777,N_11419,N_11470);
nand U11778 (N_11778,N_11629,N_11448);
xor U11779 (N_11779,N_11660,N_11403);
nor U11780 (N_11780,N_11431,N_11608);
nand U11781 (N_11781,N_11590,N_11583);
or U11782 (N_11782,N_11476,N_11643);
and U11783 (N_11783,N_11669,N_11570);
and U11784 (N_11784,N_11535,N_11479);
xnor U11785 (N_11785,N_11414,N_11426);
or U11786 (N_11786,N_11478,N_11423);
and U11787 (N_11787,N_11521,N_11620);
nand U11788 (N_11788,N_11659,N_11684);
nor U11789 (N_11789,N_11592,N_11654);
nor U11790 (N_11790,N_11544,N_11549);
nor U11791 (N_11791,N_11598,N_11433);
xnor U11792 (N_11792,N_11602,N_11690);
and U11793 (N_11793,N_11466,N_11503);
nand U11794 (N_11794,N_11495,N_11418);
nor U11795 (N_11795,N_11672,N_11443);
nand U11796 (N_11796,N_11578,N_11650);
and U11797 (N_11797,N_11572,N_11584);
nand U11798 (N_11798,N_11661,N_11604);
or U11799 (N_11799,N_11596,N_11691);
and U11800 (N_11800,N_11487,N_11441);
and U11801 (N_11801,N_11631,N_11599);
xnor U11802 (N_11802,N_11449,N_11520);
nand U11803 (N_11803,N_11639,N_11563);
nor U11804 (N_11804,N_11402,N_11541);
or U11805 (N_11805,N_11491,N_11652);
nor U11806 (N_11806,N_11530,N_11463);
or U11807 (N_11807,N_11522,N_11681);
and U11808 (N_11808,N_11623,N_11506);
nor U11809 (N_11809,N_11494,N_11605);
and U11810 (N_11810,N_11574,N_11616);
xor U11811 (N_11811,N_11532,N_11509);
xor U11812 (N_11812,N_11656,N_11525);
xor U11813 (N_11813,N_11446,N_11412);
xor U11814 (N_11814,N_11512,N_11538);
nor U11815 (N_11815,N_11633,N_11577);
or U11816 (N_11816,N_11695,N_11456);
nor U11817 (N_11817,N_11644,N_11619);
and U11818 (N_11818,N_11651,N_11458);
and U11819 (N_11819,N_11480,N_11462);
nor U11820 (N_11820,N_11640,N_11400);
nor U11821 (N_11821,N_11626,N_11523);
and U11822 (N_11822,N_11625,N_11555);
and U11823 (N_11823,N_11545,N_11438);
nor U11824 (N_11824,N_11421,N_11537);
or U11825 (N_11825,N_11607,N_11586);
or U11826 (N_11826,N_11666,N_11464);
nand U11827 (N_11827,N_11641,N_11618);
nand U11828 (N_11828,N_11576,N_11696);
nand U11829 (N_11829,N_11493,N_11664);
or U11830 (N_11830,N_11635,N_11649);
nand U11831 (N_11831,N_11461,N_11411);
nand U11832 (N_11832,N_11692,N_11504);
nand U11833 (N_11833,N_11556,N_11698);
nor U11834 (N_11834,N_11674,N_11582);
nand U11835 (N_11835,N_11505,N_11624);
or U11836 (N_11836,N_11507,N_11527);
or U11837 (N_11837,N_11508,N_11439);
and U11838 (N_11838,N_11536,N_11407);
and U11839 (N_11839,N_11632,N_11514);
xnor U11840 (N_11840,N_11409,N_11673);
and U11841 (N_11841,N_11424,N_11450);
nand U11842 (N_11842,N_11452,N_11588);
nand U11843 (N_11843,N_11453,N_11610);
xnor U11844 (N_11844,N_11612,N_11630);
or U11845 (N_11845,N_11496,N_11573);
nand U11846 (N_11846,N_11533,N_11567);
xnor U11847 (N_11847,N_11550,N_11465);
nand U11848 (N_11848,N_11485,N_11611);
and U11849 (N_11849,N_11693,N_11455);
or U11850 (N_11850,N_11584,N_11622);
and U11851 (N_11851,N_11574,N_11656);
xnor U11852 (N_11852,N_11519,N_11671);
xnor U11853 (N_11853,N_11534,N_11422);
and U11854 (N_11854,N_11503,N_11607);
and U11855 (N_11855,N_11401,N_11564);
xnor U11856 (N_11856,N_11488,N_11436);
nor U11857 (N_11857,N_11690,N_11693);
nor U11858 (N_11858,N_11688,N_11580);
nand U11859 (N_11859,N_11506,N_11552);
nand U11860 (N_11860,N_11638,N_11543);
and U11861 (N_11861,N_11620,N_11602);
and U11862 (N_11862,N_11633,N_11533);
xnor U11863 (N_11863,N_11437,N_11543);
and U11864 (N_11864,N_11418,N_11486);
nand U11865 (N_11865,N_11503,N_11455);
xor U11866 (N_11866,N_11669,N_11499);
or U11867 (N_11867,N_11684,N_11638);
and U11868 (N_11868,N_11541,N_11572);
or U11869 (N_11869,N_11432,N_11558);
or U11870 (N_11870,N_11590,N_11401);
and U11871 (N_11871,N_11673,N_11435);
or U11872 (N_11872,N_11657,N_11619);
nor U11873 (N_11873,N_11632,N_11429);
nand U11874 (N_11874,N_11422,N_11553);
nand U11875 (N_11875,N_11427,N_11428);
and U11876 (N_11876,N_11456,N_11443);
nand U11877 (N_11877,N_11634,N_11517);
and U11878 (N_11878,N_11658,N_11400);
nor U11879 (N_11879,N_11455,N_11409);
nand U11880 (N_11880,N_11425,N_11424);
nor U11881 (N_11881,N_11419,N_11525);
or U11882 (N_11882,N_11463,N_11448);
or U11883 (N_11883,N_11626,N_11682);
or U11884 (N_11884,N_11679,N_11448);
and U11885 (N_11885,N_11605,N_11552);
nand U11886 (N_11886,N_11422,N_11679);
or U11887 (N_11887,N_11402,N_11442);
nor U11888 (N_11888,N_11626,N_11583);
and U11889 (N_11889,N_11487,N_11468);
nand U11890 (N_11890,N_11596,N_11432);
xnor U11891 (N_11891,N_11452,N_11445);
xor U11892 (N_11892,N_11564,N_11470);
or U11893 (N_11893,N_11459,N_11509);
nor U11894 (N_11894,N_11468,N_11433);
and U11895 (N_11895,N_11565,N_11509);
and U11896 (N_11896,N_11552,N_11594);
nand U11897 (N_11897,N_11564,N_11645);
nand U11898 (N_11898,N_11673,N_11629);
and U11899 (N_11899,N_11520,N_11672);
or U11900 (N_11900,N_11672,N_11593);
xnor U11901 (N_11901,N_11464,N_11550);
xor U11902 (N_11902,N_11419,N_11456);
nand U11903 (N_11903,N_11629,N_11644);
or U11904 (N_11904,N_11584,N_11440);
nand U11905 (N_11905,N_11620,N_11678);
or U11906 (N_11906,N_11473,N_11419);
or U11907 (N_11907,N_11516,N_11563);
xor U11908 (N_11908,N_11660,N_11699);
xnor U11909 (N_11909,N_11618,N_11576);
xnor U11910 (N_11910,N_11470,N_11554);
or U11911 (N_11911,N_11596,N_11468);
nor U11912 (N_11912,N_11663,N_11625);
xnor U11913 (N_11913,N_11480,N_11606);
xnor U11914 (N_11914,N_11627,N_11617);
nor U11915 (N_11915,N_11650,N_11565);
or U11916 (N_11916,N_11444,N_11532);
or U11917 (N_11917,N_11430,N_11575);
nor U11918 (N_11918,N_11467,N_11422);
or U11919 (N_11919,N_11424,N_11498);
xor U11920 (N_11920,N_11589,N_11487);
nand U11921 (N_11921,N_11650,N_11640);
nand U11922 (N_11922,N_11496,N_11582);
xor U11923 (N_11923,N_11449,N_11516);
and U11924 (N_11924,N_11437,N_11624);
and U11925 (N_11925,N_11489,N_11469);
nand U11926 (N_11926,N_11678,N_11409);
nor U11927 (N_11927,N_11657,N_11521);
xnor U11928 (N_11928,N_11643,N_11523);
nand U11929 (N_11929,N_11675,N_11533);
nand U11930 (N_11930,N_11653,N_11461);
nor U11931 (N_11931,N_11679,N_11578);
or U11932 (N_11932,N_11491,N_11661);
and U11933 (N_11933,N_11570,N_11578);
or U11934 (N_11934,N_11646,N_11671);
nand U11935 (N_11935,N_11545,N_11479);
nor U11936 (N_11936,N_11429,N_11554);
xor U11937 (N_11937,N_11538,N_11683);
and U11938 (N_11938,N_11694,N_11423);
nor U11939 (N_11939,N_11669,N_11534);
or U11940 (N_11940,N_11624,N_11493);
and U11941 (N_11941,N_11563,N_11519);
xnor U11942 (N_11942,N_11407,N_11573);
and U11943 (N_11943,N_11613,N_11660);
or U11944 (N_11944,N_11518,N_11422);
or U11945 (N_11945,N_11540,N_11680);
nand U11946 (N_11946,N_11494,N_11529);
or U11947 (N_11947,N_11442,N_11573);
nand U11948 (N_11948,N_11690,N_11467);
nand U11949 (N_11949,N_11407,N_11688);
nand U11950 (N_11950,N_11699,N_11403);
or U11951 (N_11951,N_11608,N_11471);
or U11952 (N_11952,N_11683,N_11670);
and U11953 (N_11953,N_11565,N_11685);
or U11954 (N_11954,N_11638,N_11554);
nor U11955 (N_11955,N_11674,N_11437);
nor U11956 (N_11956,N_11472,N_11446);
nor U11957 (N_11957,N_11648,N_11599);
and U11958 (N_11958,N_11682,N_11665);
and U11959 (N_11959,N_11401,N_11526);
xor U11960 (N_11960,N_11583,N_11451);
or U11961 (N_11961,N_11664,N_11535);
nor U11962 (N_11962,N_11685,N_11632);
nand U11963 (N_11963,N_11525,N_11593);
xor U11964 (N_11964,N_11673,N_11619);
nor U11965 (N_11965,N_11480,N_11559);
nand U11966 (N_11966,N_11636,N_11456);
or U11967 (N_11967,N_11492,N_11584);
xor U11968 (N_11968,N_11619,N_11648);
xor U11969 (N_11969,N_11455,N_11430);
xnor U11970 (N_11970,N_11528,N_11536);
and U11971 (N_11971,N_11400,N_11420);
and U11972 (N_11972,N_11507,N_11549);
and U11973 (N_11973,N_11667,N_11569);
xnor U11974 (N_11974,N_11479,N_11632);
xor U11975 (N_11975,N_11502,N_11524);
or U11976 (N_11976,N_11653,N_11599);
or U11977 (N_11977,N_11672,N_11558);
or U11978 (N_11978,N_11557,N_11463);
nor U11979 (N_11979,N_11541,N_11434);
or U11980 (N_11980,N_11695,N_11415);
xnor U11981 (N_11981,N_11406,N_11531);
and U11982 (N_11982,N_11553,N_11459);
or U11983 (N_11983,N_11693,N_11515);
xnor U11984 (N_11984,N_11458,N_11508);
nor U11985 (N_11985,N_11474,N_11691);
or U11986 (N_11986,N_11662,N_11617);
or U11987 (N_11987,N_11434,N_11657);
nand U11988 (N_11988,N_11640,N_11673);
or U11989 (N_11989,N_11473,N_11602);
nor U11990 (N_11990,N_11632,N_11445);
nor U11991 (N_11991,N_11615,N_11607);
nand U11992 (N_11992,N_11412,N_11414);
nor U11993 (N_11993,N_11411,N_11655);
nand U11994 (N_11994,N_11537,N_11534);
nor U11995 (N_11995,N_11631,N_11591);
nor U11996 (N_11996,N_11612,N_11444);
or U11997 (N_11997,N_11476,N_11673);
xor U11998 (N_11998,N_11636,N_11659);
and U11999 (N_11999,N_11446,N_11582);
xor U12000 (N_12000,N_11712,N_11821);
and U12001 (N_12001,N_11895,N_11874);
nor U12002 (N_12002,N_11826,N_11870);
or U12003 (N_12003,N_11805,N_11950);
and U12004 (N_12004,N_11735,N_11803);
xnor U12005 (N_12005,N_11916,N_11938);
and U12006 (N_12006,N_11811,N_11965);
nand U12007 (N_12007,N_11867,N_11937);
nor U12008 (N_12008,N_11987,N_11845);
and U12009 (N_12009,N_11892,N_11922);
and U12010 (N_12010,N_11994,N_11762);
nor U12011 (N_12011,N_11843,N_11827);
and U12012 (N_12012,N_11800,N_11801);
nand U12013 (N_12013,N_11782,N_11723);
or U12014 (N_12014,N_11775,N_11879);
nand U12015 (N_12015,N_11856,N_11751);
and U12016 (N_12016,N_11972,N_11899);
or U12017 (N_12017,N_11898,N_11716);
or U12018 (N_12018,N_11809,N_11822);
nor U12019 (N_12019,N_11816,N_11711);
nor U12020 (N_12020,N_11906,N_11846);
xnor U12021 (N_12021,N_11731,N_11862);
nand U12022 (N_12022,N_11741,N_11812);
and U12023 (N_12023,N_11941,N_11842);
or U12024 (N_12024,N_11838,N_11761);
and U12025 (N_12025,N_11981,N_11768);
or U12026 (N_12026,N_11792,N_11980);
xnor U12027 (N_12027,N_11736,N_11900);
nand U12028 (N_12028,N_11959,N_11920);
xor U12029 (N_12029,N_11714,N_11902);
nor U12030 (N_12030,N_11832,N_11844);
or U12031 (N_12031,N_11992,N_11797);
and U12032 (N_12032,N_11753,N_11763);
nor U12033 (N_12033,N_11884,N_11880);
nor U12034 (N_12034,N_11923,N_11943);
and U12035 (N_12035,N_11745,N_11926);
or U12036 (N_12036,N_11836,N_11869);
or U12037 (N_12037,N_11705,N_11828);
nand U12038 (N_12038,N_11726,N_11969);
or U12039 (N_12039,N_11730,N_11947);
nand U12040 (N_12040,N_11991,N_11964);
or U12041 (N_12041,N_11982,N_11848);
or U12042 (N_12042,N_11772,N_11977);
xor U12043 (N_12043,N_11984,N_11993);
nand U12044 (N_12044,N_11917,N_11910);
and U12045 (N_12045,N_11933,N_11894);
nand U12046 (N_12046,N_11824,N_11791);
nor U12047 (N_12047,N_11854,N_11949);
and U12048 (N_12048,N_11935,N_11976);
and U12049 (N_12049,N_11721,N_11960);
and U12050 (N_12050,N_11742,N_11759);
nor U12051 (N_12051,N_11882,N_11789);
and U12052 (N_12052,N_11897,N_11860);
nand U12053 (N_12053,N_11784,N_11804);
and U12054 (N_12054,N_11810,N_11718);
nand U12055 (N_12055,N_11924,N_11795);
nor U12056 (N_12056,N_11866,N_11806);
nor U12057 (N_12057,N_11825,N_11889);
nand U12058 (N_12058,N_11748,N_11975);
nor U12059 (N_12059,N_11749,N_11750);
and U12060 (N_12060,N_11781,N_11799);
nand U12061 (N_12061,N_11814,N_11903);
nor U12062 (N_12062,N_11754,N_11934);
and U12063 (N_12063,N_11946,N_11872);
nor U12064 (N_12064,N_11757,N_11953);
or U12065 (N_12065,N_11907,N_11998);
nor U12066 (N_12066,N_11706,N_11853);
nand U12067 (N_12067,N_11807,N_11888);
nand U12068 (N_12068,N_11700,N_11715);
nor U12069 (N_12069,N_11904,N_11999);
xor U12070 (N_12070,N_11883,N_11841);
nand U12071 (N_12071,N_11720,N_11722);
nand U12072 (N_12072,N_11908,N_11771);
xnor U12073 (N_12073,N_11985,N_11927);
xnor U12074 (N_12074,N_11817,N_11939);
xor U12075 (N_12075,N_11905,N_11914);
or U12076 (N_12076,N_11861,N_11776);
nor U12077 (N_12077,N_11778,N_11855);
and U12078 (N_12078,N_11983,N_11995);
nand U12079 (N_12079,N_11990,N_11833);
xnor U12080 (N_12080,N_11743,N_11859);
or U12081 (N_12081,N_11793,N_11737);
nand U12082 (N_12082,N_11978,N_11858);
nor U12083 (N_12083,N_11948,N_11760);
or U12084 (N_12084,N_11819,N_11729);
nand U12085 (N_12085,N_11878,N_11971);
and U12086 (N_12086,N_11864,N_11790);
or U12087 (N_12087,N_11871,N_11945);
or U12088 (N_12088,N_11961,N_11918);
nor U12089 (N_12089,N_11876,N_11967);
xor U12090 (N_12090,N_11837,N_11732);
or U12091 (N_12091,N_11932,N_11930);
or U12092 (N_12092,N_11875,N_11955);
and U12093 (N_12093,N_11713,N_11952);
nor U12094 (N_12094,N_11777,N_11830);
nor U12095 (N_12095,N_11786,N_11909);
and U12096 (N_12096,N_11849,N_11954);
xnor U12097 (N_12097,N_11708,N_11988);
xnor U12098 (N_12098,N_11709,N_11840);
or U12099 (N_12099,N_11766,N_11733);
nor U12100 (N_12100,N_11752,N_11957);
and U12101 (N_12101,N_11783,N_11746);
and U12102 (N_12102,N_11813,N_11802);
or U12103 (N_12103,N_11857,N_11765);
and U12104 (N_12104,N_11928,N_11758);
nor U12105 (N_12105,N_11796,N_11767);
nor U12106 (N_12106,N_11850,N_11929);
and U12107 (N_12107,N_11808,N_11703);
nor U12108 (N_12108,N_11891,N_11707);
nand U12109 (N_12109,N_11823,N_11986);
xnor U12110 (N_12110,N_11893,N_11925);
or U12111 (N_12111,N_11764,N_11996);
nor U12112 (N_12112,N_11734,N_11829);
xnor U12113 (N_12113,N_11719,N_11873);
nor U12114 (N_12114,N_11727,N_11728);
nor U12115 (N_12115,N_11725,N_11785);
nand U12116 (N_12116,N_11755,N_11962);
nand U12117 (N_12117,N_11968,N_11798);
xnor U12118 (N_12118,N_11717,N_11944);
and U12119 (N_12119,N_11912,N_11958);
nor U12120 (N_12120,N_11970,N_11877);
nor U12121 (N_12121,N_11911,N_11747);
xnor U12122 (N_12122,N_11710,N_11702);
or U12123 (N_12123,N_11973,N_11921);
nor U12124 (N_12124,N_11834,N_11966);
nor U12125 (N_12125,N_11738,N_11890);
nor U12126 (N_12126,N_11963,N_11769);
and U12127 (N_12127,N_11724,N_11989);
xor U12128 (N_12128,N_11704,N_11779);
nor U12129 (N_12129,N_11770,N_11831);
nor U12130 (N_12130,N_11868,N_11865);
xor U12131 (N_12131,N_11852,N_11896);
or U12132 (N_12132,N_11787,N_11919);
nand U12133 (N_12133,N_11997,N_11940);
xnor U12134 (N_12134,N_11820,N_11835);
xnor U12135 (N_12135,N_11887,N_11851);
nand U12136 (N_12136,N_11774,N_11913);
and U12137 (N_12137,N_11839,N_11773);
nand U12138 (N_12138,N_11815,N_11788);
or U12139 (N_12139,N_11956,N_11744);
or U12140 (N_12140,N_11756,N_11740);
xor U12141 (N_12141,N_11863,N_11979);
nor U12142 (N_12142,N_11739,N_11885);
or U12143 (N_12143,N_11915,N_11974);
nand U12144 (N_12144,N_11942,N_11818);
xnor U12145 (N_12145,N_11936,N_11847);
nand U12146 (N_12146,N_11931,N_11701);
nand U12147 (N_12147,N_11951,N_11794);
nand U12148 (N_12148,N_11780,N_11901);
nor U12149 (N_12149,N_11881,N_11886);
or U12150 (N_12150,N_11945,N_11749);
xnor U12151 (N_12151,N_11919,N_11894);
xnor U12152 (N_12152,N_11978,N_11779);
nor U12153 (N_12153,N_11867,N_11739);
nand U12154 (N_12154,N_11831,N_11709);
nand U12155 (N_12155,N_11873,N_11794);
nor U12156 (N_12156,N_11747,N_11910);
xor U12157 (N_12157,N_11748,N_11769);
nor U12158 (N_12158,N_11801,N_11886);
nor U12159 (N_12159,N_11722,N_11706);
and U12160 (N_12160,N_11971,N_11937);
nand U12161 (N_12161,N_11831,N_11718);
nor U12162 (N_12162,N_11716,N_11979);
and U12163 (N_12163,N_11772,N_11842);
xor U12164 (N_12164,N_11768,N_11893);
and U12165 (N_12165,N_11896,N_11816);
nand U12166 (N_12166,N_11798,N_11728);
or U12167 (N_12167,N_11737,N_11988);
xnor U12168 (N_12168,N_11927,N_11728);
and U12169 (N_12169,N_11871,N_11843);
xnor U12170 (N_12170,N_11864,N_11865);
nor U12171 (N_12171,N_11764,N_11815);
nor U12172 (N_12172,N_11977,N_11838);
nand U12173 (N_12173,N_11707,N_11807);
xnor U12174 (N_12174,N_11972,N_11933);
and U12175 (N_12175,N_11879,N_11901);
nor U12176 (N_12176,N_11868,N_11846);
xnor U12177 (N_12177,N_11788,N_11811);
xor U12178 (N_12178,N_11983,N_11973);
and U12179 (N_12179,N_11986,N_11774);
xor U12180 (N_12180,N_11982,N_11811);
and U12181 (N_12181,N_11769,N_11713);
xnor U12182 (N_12182,N_11935,N_11980);
or U12183 (N_12183,N_11920,N_11966);
nor U12184 (N_12184,N_11789,N_11919);
nor U12185 (N_12185,N_11923,N_11908);
nor U12186 (N_12186,N_11955,N_11896);
and U12187 (N_12187,N_11756,N_11967);
nor U12188 (N_12188,N_11846,N_11749);
nand U12189 (N_12189,N_11985,N_11789);
nand U12190 (N_12190,N_11784,N_11742);
or U12191 (N_12191,N_11874,N_11865);
nand U12192 (N_12192,N_11887,N_11987);
or U12193 (N_12193,N_11873,N_11764);
or U12194 (N_12194,N_11759,N_11960);
xnor U12195 (N_12195,N_11817,N_11742);
xnor U12196 (N_12196,N_11828,N_11826);
or U12197 (N_12197,N_11950,N_11791);
xor U12198 (N_12198,N_11797,N_11749);
nor U12199 (N_12199,N_11781,N_11971);
nor U12200 (N_12200,N_11783,N_11972);
or U12201 (N_12201,N_11795,N_11849);
and U12202 (N_12202,N_11978,N_11748);
or U12203 (N_12203,N_11903,N_11785);
and U12204 (N_12204,N_11726,N_11705);
nand U12205 (N_12205,N_11798,N_11780);
xnor U12206 (N_12206,N_11895,N_11906);
and U12207 (N_12207,N_11882,N_11874);
or U12208 (N_12208,N_11727,N_11873);
nand U12209 (N_12209,N_11989,N_11967);
nor U12210 (N_12210,N_11700,N_11982);
and U12211 (N_12211,N_11798,N_11768);
xor U12212 (N_12212,N_11707,N_11991);
or U12213 (N_12213,N_11880,N_11809);
nor U12214 (N_12214,N_11827,N_11936);
or U12215 (N_12215,N_11804,N_11708);
or U12216 (N_12216,N_11954,N_11837);
or U12217 (N_12217,N_11775,N_11906);
nor U12218 (N_12218,N_11971,N_11714);
nand U12219 (N_12219,N_11930,N_11913);
nor U12220 (N_12220,N_11866,N_11960);
nand U12221 (N_12221,N_11862,N_11705);
nand U12222 (N_12222,N_11848,N_11935);
or U12223 (N_12223,N_11985,N_11802);
nand U12224 (N_12224,N_11723,N_11938);
or U12225 (N_12225,N_11787,N_11821);
and U12226 (N_12226,N_11739,N_11702);
and U12227 (N_12227,N_11739,N_11711);
and U12228 (N_12228,N_11935,N_11939);
nor U12229 (N_12229,N_11764,N_11875);
and U12230 (N_12230,N_11715,N_11939);
nor U12231 (N_12231,N_11955,N_11704);
nand U12232 (N_12232,N_11771,N_11888);
xnor U12233 (N_12233,N_11866,N_11872);
and U12234 (N_12234,N_11858,N_11907);
nor U12235 (N_12235,N_11951,N_11709);
nor U12236 (N_12236,N_11971,N_11818);
nor U12237 (N_12237,N_11719,N_11952);
xnor U12238 (N_12238,N_11830,N_11764);
and U12239 (N_12239,N_11701,N_11898);
nand U12240 (N_12240,N_11765,N_11981);
nor U12241 (N_12241,N_11817,N_11920);
xor U12242 (N_12242,N_11907,N_11875);
nor U12243 (N_12243,N_11907,N_11911);
or U12244 (N_12244,N_11946,N_11911);
or U12245 (N_12245,N_11942,N_11859);
and U12246 (N_12246,N_11843,N_11938);
nand U12247 (N_12247,N_11989,N_11754);
nor U12248 (N_12248,N_11927,N_11802);
and U12249 (N_12249,N_11992,N_11796);
xor U12250 (N_12250,N_11754,N_11761);
nand U12251 (N_12251,N_11813,N_11812);
nand U12252 (N_12252,N_11869,N_11802);
nand U12253 (N_12253,N_11810,N_11878);
or U12254 (N_12254,N_11714,N_11910);
or U12255 (N_12255,N_11981,N_11887);
or U12256 (N_12256,N_11728,N_11932);
xnor U12257 (N_12257,N_11897,N_11847);
nand U12258 (N_12258,N_11715,N_11851);
xor U12259 (N_12259,N_11952,N_11765);
nand U12260 (N_12260,N_11918,N_11766);
nand U12261 (N_12261,N_11931,N_11954);
or U12262 (N_12262,N_11884,N_11775);
and U12263 (N_12263,N_11705,N_11964);
xnor U12264 (N_12264,N_11867,N_11836);
xor U12265 (N_12265,N_11910,N_11956);
nor U12266 (N_12266,N_11972,N_11893);
and U12267 (N_12267,N_11720,N_11947);
and U12268 (N_12268,N_11901,N_11762);
and U12269 (N_12269,N_11775,N_11799);
or U12270 (N_12270,N_11858,N_11712);
and U12271 (N_12271,N_11899,N_11770);
and U12272 (N_12272,N_11771,N_11854);
nand U12273 (N_12273,N_11920,N_11822);
and U12274 (N_12274,N_11712,N_11781);
xor U12275 (N_12275,N_11925,N_11815);
or U12276 (N_12276,N_11999,N_11719);
or U12277 (N_12277,N_11976,N_11842);
xnor U12278 (N_12278,N_11940,N_11908);
nand U12279 (N_12279,N_11817,N_11883);
and U12280 (N_12280,N_11862,N_11769);
and U12281 (N_12281,N_11959,N_11845);
nor U12282 (N_12282,N_11964,N_11930);
nor U12283 (N_12283,N_11890,N_11772);
nor U12284 (N_12284,N_11737,N_11893);
or U12285 (N_12285,N_11921,N_11892);
nor U12286 (N_12286,N_11902,N_11827);
nor U12287 (N_12287,N_11853,N_11971);
xnor U12288 (N_12288,N_11869,N_11873);
or U12289 (N_12289,N_11795,N_11952);
xor U12290 (N_12290,N_11816,N_11860);
nor U12291 (N_12291,N_11827,N_11900);
and U12292 (N_12292,N_11965,N_11938);
nor U12293 (N_12293,N_11856,N_11992);
xor U12294 (N_12294,N_11787,N_11827);
nand U12295 (N_12295,N_11753,N_11943);
nand U12296 (N_12296,N_11705,N_11710);
and U12297 (N_12297,N_11772,N_11862);
nand U12298 (N_12298,N_11840,N_11784);
xnor U12299 (N_12299,N_11894,N_11963);
or U12300 (N_12300,N_12019,N_12174);
nand U12301 (N_12301,N_12245,N_12214);
nand U12302 (N_12302,N_12079,N_12118);
nor U12303 (N_12303,N_12018,N_12142);
or U12304 (N_12304,N_12060,N_12171);
or U12305 (N_12305,N_12216,N_12059);
or U12306 (N_12306,N_12194,N_12246);
xor U12307 (N_12307,N_12011,N_12092);
and U12308 (N_12308,N_12058,N_12145);
nor U12309 (N_12309,N_12232,N_12243);
xor U12310 (N_12310,N_12144,N_12131);
nor U12311 (N_12311,N_12101,N_12028);
and U12312 (N_12312,N_12136,N_12147);
xor U12313 (N_12313,N_12062,N_12017);
nor U12314 (N_12314,N_12172,N_12029);
xor U12315 (N_12315,N_12100,N_12225);
nor U12316 (N_12316,N_12219,N_12054);
xnor U12317 (N_12317,N_12117,N_12266);
nand U12318 (N_12318,N_12251,N_12258);
nand U12319 (N_12319,N_12153,N_12031);
xor U12320 (N_12320,N_12154,N_12016);
xor U12321 (N_12321,N_12257,N_12247);
or U12322 (N_12322,N_12264,N_12066);
xor U12323 (N_12323,N_12170,N_12040);
nor U12324 (N_12324,N_12033,N_12067);
or U12325 (N_12325,N_12150,N_12269);
or U12326 (N_12326,N_12037,N_12053);
nand U12327 (N_12327,N_12096,N_12263);
and U12328 (N_12328,N_12122,N_12157);
nand U12329 (N_12329,N_12270,N_12267);
xnor U12330 (N_12330,N_12006,N_12215);
or U12331 (N_12331,N_12143,N_12176);
xnor U12332 (N_12332,N_12293,N_12074);
and U12333 (N_12333,N_12152,N_12111);
xnor U12334 (N_12334,N_12272,N_12201);
and U12335 (N_12335,N_12109,N_12296);
or U12336 (N_12336,N_12119,N_12043);
xor U12337 (N_12337,N_12129,N_12090);
nand U12338 (N_12338,N_12095,N_12127);
nor U12339 (N_12339,N_12038,N_12291);
or U12340 (N_12340,N_12072,N_12009);
nor U12341 (N_12341,N_12022,N_12000);
and U12342 (N_12342,N_12250,N_12180);
xnor U12343 (N_12343,N_12107,N_12056);
nor U12344 (N_12344,N_12173,N_12024);
and U12345 (N_12345,N_12212,N_12160);
xor U12346 (N_12346,N_12290,N_12032);
nand U12347 (N_12347,N_12244,N_12004);
nand U12348 (N_12348,N_12086,N_12146);
nor U12349 (N_12349,N_12030,N_12242);
xnor U12350 (N_12350,N_12276,N_12190);
nand U12351 (N_12351,N_12260,N_12163);
and U12352 (N_12352,N_12284,N_12078);
nand U12353 (N_12353,N_12139,N_12188);
or U12354 (N_12354,N_12230,N_12262);
and U12355 (N_12355,N_12076,N_12121);
or U12356 (N_12356,N_12034,N_12192);
or U12357 (N_12357,N_12141,N_12283);
xor U12358 (N_12358,N_12233,N_12197);
or U12359 (N_12359,N_12104,N_12097);
or U12360 (N_12360,N_12140,N_12281);
nand U12361 (N_12361,N_12259,N_12158);
and U12362 (N_12362,N_12252,N_12110);
and U12363 (N_12363,N_12021,N_12186);
nor U12364 (N_12364,N_12205,N_12108);
xor U12365 (N_12365,N_12049,N_12134);
and U12366 (N_12366,N_12130,N_12268);
xor U12367 (N_12367,N_12105,N_12255);
nand U12368 (N_12368,N_12013,N_12206);
nand U12369 (N_12369,N_12189,N_12112);
and U12370 (N_12370,N_12099,N_12210);
xor U12371 (N_12371,N_12120,N_12159);
or U12372 (N_12372,N_12227,N_12229);
or U12373 (N_12373,N_12115,N_12015);
nor U12374 (N_12374,N_12231,N_12014);
nand U12375 (N_12375,N_12133,N_12277);
nand U12376 (N_12376,N_12077,N_12237);
xor U12377 (N_12377,N_12084,N_12080);
or U12378 (N_12378,N_12203,N_12199);
and U12379 (N_12379,N_12063,N_12007);
nor U12380 (N_12380,N_12012,N_12036);
and U12381 (N_12381,N_12087,N_12178);
nor U12382 (N_12382,N_12195,N_12184);
xnor U12383 (N_12383,N_12202,N_12102);
nor U12384 (N_12384,N_12116,N_12200);
nand U12385 (N_12385,N_12208,N_12274);
nand U12386 (N_12386,N_12070,N_12135);
or U12387 (N_12387,N_12023,N_12295);
nand U12388 (N_12388,N_12299,N_12224);
or U12389 (N_12389,N_12048,N_12287);
xnor U12390 (N_12390,N_12228,N_12236);
nand U12391 (N_12391,N_12156,N_12113);
nand U12392 (N_12392,N_12273,N_12137);
nor U12393 (N_12393,N_12183,N_12047);
nand U12394 (N_12394,N_12285,N_12039);
xnor U12395 (N_12395,N_12106,N_12148);
and U12396 (N_12396,N_12292,N_12114);
and U12397 (N_12397,N_12179,N_12051);
nand U12398 (N_12398,N_12068,N_12223);
xor U12399 (N_12399,N_12278,N_12123);
and U12400 (N_12400,N_12003,N_12149);
or U12401 (N_12401,N_12249,N_12041);
nor U12402 (N_12402,N_12089,N_12103);
nand U12403 (N_12403,N_12220,N_12005);
xnor U12404 (N_12404,N_12128,N_12085);
xor U12405 (N_12405,N_12168,N_12052);
or U12406 (N_12406,N_12193,N_12044);
xnor U12407 (N_12407,N_12280,N_12075);
or U12408 (N_12408,N_12254,N_12177);
xnor U12409 (N_12409,N_12198,N_12234);
nor U12410 (N_12410,N_12046,N_12162);
and U12411 (N_12411,N_12167,N_12235);
and U12412 (N_12412,N_12161,N_12204);
xor U12413 (N_12413,N_12238,N_12138);
nand U12414 (N_12414,N_12045,N_12191);
nand U12415 (N_12415,N_12221,N_12185);
nor U12416 (N_12416,N_12265,N_12166);
or U12417 (N_12417,N_12207,N_12226);
nand U12418 (N_12418,N_12002,N_12298);
nor U12419 (N_12419,N_12001,N_12010);
and U12420 (N_12420,N_12248,N_12271);
nor U12421 (N_12421,N_12042,N_12294);
and U12422 (N_12422,N_12050,N_12061);
or U12423 (N_12423,N_12125,N_12094);
xor U12424 (N_12424,N_12241,N_12217);
or U12425 (N_12425,N_12196,N_12124);
nand U12426 (N_12426,N_12169,N_12093);
nor U12427 (N_12427,N_12151,N_12261);
and U12428 (N_12428,N_12279,N_12155);
nand U12429 (N_12429,N_12182,N_12091);
xnor U12430 (N_12430,N_12175,N_12055);
nor U12431 (N_12431,N_12098,N_12057);
or U12432 (N_12432,N_12289,N_12081);
nor U12433 (N_12433,N_12073,N_12027);
nand U12434 (N_12434,N_12126,N_12211);
nand U12435 (N_12435,N_12297,N_12240);
or U12436 (N_12436,N_12218,N_12187);
or U12437 (N_12437,N_12165,N_12035);
and U12438 (N_12438,N_12020,N_12222);
or U12439 (N_12439,N_12071,N_12069);
and U12440 (N_12440,N_12282,N_12275);
or U12441 (N_12441,N_12164,N_12082);
xnor U12442 (N_12442,N_12088,N_12256);
xnor U12443 (N_12443,N_12025,N_12083);
xnor U12444 (N_12444,N_12213,N_12065);
and U12445 (N_12445,N_12132,N_12181);
nand U12446 (N_12446,N_12064,N_12026);
and U12447 (N_12447,N_12286,N_12253);
nand U12448 (N_12448,N_12209,N_12008);
or U12449 (N_12449,N_12239,N_12288);
nand U12450 (N_12450,N_12297,N_12077);
and U12451 (N_12451,N_12212,N_12237);
or U12452 (N_12452,N_12289,N_12067);
nor U12453 (N_12453,N_12079,N_12158);
and U12454 (N_12454,N_12163,N_12247);
xnor U12455 (N_12455,N_12052,N_12192);
or U12456 (N_12456,N_12157,N_12260);
nor U12457 (N_12457,N_12160,N_12193);
xnor U12458 (N_12458,N_12239,N_12065);
nand U12459 (N_12459,N_12044,N_12177);
nand U12460 (N_12460,N_12103,N_12102);
xor U12461 (N_12461,N_12037,N_12060);
and U12462 (N_12462,N_12041,N_12063);
xor U12463 (N_12463,N_12276,N_12128);
nor U12464 (N_12464,N_12184,N_12215);
nand U12465 (N_12465,N_12127,N_12251);
and U12466 (N_12466,N_12135,N_12174);
or U12467 (N_12467,N_12158,N_12032);
nand U12468 (N_12468,N_12038,N_12262);
and U12469 (N_12469,N_12214,N_12278);
nand U12470 (N_12470,N_12244,N_12299);
or U12471 (N_12471,N_12025,N_12116);
nand U12472 (N_12472,N_12198,N_12169);
xor U12473 (N_12473,N_12286,N_12093);
xnor U12474 (N_12474,N_12139,N_12017);
xor U12475 (N_12475,N_12050,N_12101);
and U12476 (N_12476,N_12274,N_12275);
nor U12477 (N_12477,N_12057,N_12020);
or U12478 (N_12478,N_12265,N_12003);
nor U12479 (N_12479,N_12061,N_12053);
and U12480 (N_12480,N_12279,N_12223);
xnor U12481 (N_12481,N_12001,N_12255);
nand U12482 (N_12482,N_12283,N_12041);
nor U12483 (N_12483,N_12274,N_12025);
or U12484 (N_12484,N_12122,N_12193);
or U12485 (N_12485,N_12075,N_12178);
and U12486 (N_12486,N_12157,N_12027);
and U12487 (N_12487,N_12280,N_12010);
and U12488 (N_12488,N_12190,N_12208);
nor U12489 (N_12489,N_12081,N_12038);
and U12490 (N_12490,N_12048,N_12262);
and U12491 (N_12491,N_12246,N_12180);
and U12492 (N_12492,N_12050,N_12001);
or U12493 (N_12493,N_12286,N_12205);
nor U12494 (N_12494,N_12072,N_12083);
and U12495 (N_12495,N_12196,N_12085);
xor U12496 (N_12496,N_12264,N_12036);
or U12497 (N_12497,N_12218,N_12152);
nor U12498 (N_12498,N_12023,N_12125);
or U12499 (N_12499,N_12025,N_12250);
xor U12500 (N_12500,N_12022,N_12252);
or U12501 (N_12501,N_12088,N_12027);
and U12502 (N_12502,N_12054,N_12162);
nand U12503 (N_12503,N_12159,N_12292);
and U12504 (N_12504,N_12294,N_12153);
nor U12505 (N_12505,N_12062,N_12080);
or U12506 (N_12506,N_12238,N_12069);
nor U12507 (N_12507,N_12242,N_12150);
nand U12508 (N_12508,N_12016,N_12155);
and U12509 (N_12509,N_12178,N_12006);
or U12510 (N_12510,N_12186,N_12191);
xnor U12511 (N_12511,N_12014,N_12065);
xor U12512 (N_12512,N_12276,N_12193);
nand U12513 (N_12513,N_12195,N_12063);
nand U12514 (N_12514,N_12238,N_12167);
nand U12515 (N_12515,N_12141,N_12290);
and U12516 (N_12516,N_12190,N_12139);
nand U12517 (N_12517,N_12145,N_12287);
nor U12518 (N_12518,N_12023,N_12081);
xnor U12519 (N_12519,N_12280,N_12063);
nor U12520 (N_12520,N_12228,N_12255);
xnor U12521 (N_12521,N_12152,N_12011);
or U12522 (N_12522,N_12014,N_12132);
xnor U12523 (N_12523,N_12113,N_12124);
or U12524 (N_12524,N_12046,N_12084);
and U12525 (N_12525,N_12094,N_12193);
and U12526 (N_12526,N_12110,N_12112);
and U12527 (N_12527,N_12038,N_12234);
or U12528 (N_12528,N_12035,N_12186);
nor U12529 (N_12529,N_12011,N_12164);
nor U12530 (N_12530,N_12128,N_12157);
and U12531 (N_12531,N_12196,N_12037);
xnor U12532 (N_12532,N_12172,N_12263);
nand U12533 (N_12533,N_12140,N_12257);
xnor U12534 (N_12534,N_12239,N_12045);
nor U12535 (N_12535,N_12060,N_12109);
and U12536 (N_12536,N_12186,N_12193);
or U12537 (N_12537,N_12041,N_12048);
nor U12538 (N_12538,N_12182,N_12043);
nand U12539 (N_12539,N_12287,N_12245);
and U12540 (N_12540,N_12219,N_12107);
nand U12541 (N_12541,N_12277,N_12000);
xor U12542 (N_12542,N_12142,N_12003);
or U12543 (N_12543,N_12274,N_12195);
nor U12544 (N_12544,N_12241,N_12094);
or U12545 (N_12545,N_12281,N_12283);
nand U12546 (N_12546,N_12095,N_12159);
nor U12547 (N_12547,N_12280,N_12241);
or U12548 (N_12548,N_12268,N_12234);
nand U12549 (N_12549,N_12177,N_12211);
nor U12550 (N_12550,N_12036,N_12196);
or U12551 (N_12551,N_12092,N_12166);
xnor U12552 (N_12552,N_12048,N_12198);
or U12553 (N_12553,N_12184,N_12136);
nor U12554 (N_12554,N_12199,N_12064);
xnor U12555 (N_12555,N_12046,N_12276);
and U12556 (N_12556,N_12286,N_12262);
or U12557 (N_12557,N_12100,N_12217);
and U12558 (N_12558,N_12181,N_12080);
nand U12559 (N_12559,N_12210,N_12024);
and U12560 (N_12560,N_12049,N_12243);
xor U12561 (N_12561,N_12235,N_12146);
and U12562 (N_12562,N_12245,N_12209);
nand U12563 (N_12563,N_12002,N_12293);
nor U12564 (N_12564,N_12197,N_12107);
and U12565 (N_12565,N_12240,N_12065);
xnor U12566 (N_12566,N_12070,N_12210);
and U12567 (N_12567,N_12115,N_12155);
xor U12568 (N_12568,N_12281,N_12099);
xor U12569 (N_12569,N_12127,N_12258);
xor U12570 (N_12570,N_12228,N_12080);
and U12571 (N_12571,N_12152,N_12220);
and U12572 (N_12572,N_12055,N_12285);
and U12573 (N_12573,N_12139,N_12216);
and U12574 (N_12574,N_12096,N_12213);
or U12575 (N_12575,N_12084,N_12088);
nand U12576 (N_12576,N_12144,N_12235);
xor U12577 (N_12577,N_12225,N_12057);
nand U12578 (N_12578,N_12246,N_12149);
or U12579 (N_12579,N_12007,N_12003);
nor U12580 (N_12580,N_12274,N_12104);
and U12581 (N_12581,N_12029,N_12167);
or U12582 (N_12582,N_12038,N_12226);
nand U12583 (N_12583,N_12015,N_12253);
nand U12584 (N_12584,N_12077,N_12013);
nand U12585 (N_12585,N_12176,N_12139);
nor U12586 (N_12586,N_12264,N_12175);
nor U12587 (N_12587,N_12174,N_12028);
xor U12588 (N_12588,N_12085,N_12059);
or U12589 (N_12589,N_12096,N_12024);
and U12590 (N_12590,N_12078,N_12174);
nand U12591 (N_12591,N_12096,N_12265);
nor U12592 (N_12592,N_12002,N_12223);
xnor U12593 (N_12593,N_12064,N_12269);
or U12594 (N_12594,N_12043,N_12003);
nor U12595 (N_12595,N_12169,N_12050);
or U12596 (N_12596,N_12164,N_12117);
nand U12597 (N_12597,N_12206,N_12184);
xor U12598 (N_12598,N_12010,N_12296);
or U12599 (N_12599,N_12231,N_12102);
and U12600 (N_12600,N_12461,N_12393);
nand U12601 (N_12601,N_12401,N_12412);
and U12602 (N_12602,N_12356,N_12431);
xor U12603 (N_12603,N_12436,N_12538);
nand U12604 (N_12604,N_12333,N_12512);
xor U12605 (N_12605,N_12334,N_12561);
and U12606 (N_12606,N_12300,N_12419);
nand U12607 (N_12607,N_12439,N_12345);
nor U12608 (N_12608,N_12408,N_12591);
xnor U12609 (N_12609,N_12448,N_12596);
and U12610 (N_12610,N_12368,N_12315);
xnor U12611 (N_12611,N_12380,N_12305);
nor U12612 (N_12612,N_12579,N_12492);
or U12613 (N_12613,N_12336,N_12599);
nor U12614 (N_12614,N_12468,N_12396);
nor U12615 (N_12615,N_12351,N_12577);
nand U12616 (N_12616,N_12500,N_12574);
xnor U12617 (N_12617,N_12306,N_12455);
nor U12618 (N_12618,N_12411,N_12421);
xnor U12619 (N_12619,N_12328,N_12312);
nand U12620 (N_12620,N_12390,N_12330);
xor U12621 (N_12621,N_12331,N_12418);
or U12622 (N_12622,N_12363,N_12435);
and U12623 (N_12623,N_12589,N_12536);
and U12624 (N_12624,N_12511,N_12495);
nor U12625 (N_12625,N_12433,N_12598);
or U12626 (N_12626,N_12490,N_12587);
nand U12627 (N_12627,N_12365,N_12434);
and U12628 (N_12628,N_12357,N_12387);
xor U12629 (N_12629,N_12469,N_12338);
xor U12630 (N_12630,N_12335,N_12402);
nand U12631 (N_12631,N_12485,N_12568);
xnor U12632 (N_12632,N_12530,N_12456);
nand U12633 (N_12633,N_12354,N_12420);
or U12634 (N_12634,N_12593,N_12339);
and U12635 (N_12635,N_12491,N_12590);
or U12636 (N_12636,N_12484,N_12551);
xnor U12637 (N_12637,N_12503,N_12454);
xor U12638 (N_12638,N_12376,N_12509);
nor U12639 (N_12639,N_12447,N_12475);
nand U12640 (N_12640,N_12580,N_12319);
nand U12641 (N_12641,N_12426,N_12374);
and U12642 (N_12642,N_12405,N_12377);
xnor U12643 (N_12643,N_12443,N_12440);
nor U12644 (N_12644,N_12459,N_12321);
nor U12645 (N_12645,N_12373,N_12352);
nand U12646 (N_12646,N_12597,N_12566);
and U12647 (N_12647,N_12432,N_12358);
xor U12648 (N_12648,N_12323,N_12449);
nor U12649 (N_12649,N_12350,N_12310);
nor U12650 (N_12650,N_12472,N_12481);
and U12651 (N_12651,N_12592,N_12437);
nand U12652 (N_12652,N_12406,N_12410);
and U12653 (N_12653,N_12366,N_12375);
nand U12654 (N_12654,N_12582,N_12462);
nor U12655 (N_12655,N_12570,N_12471);
or U12656 (N_12656,N_12559,N_12325);
and U12657 (N_12657,N_12514,N_12362);
and U12658 (N_12658,N_12516,N_12318);
and U12659 (N_12659,N_12554,N_12422);
and U12660 (N_12660,N_12483,N_12413);
xor U12661 (N_12661,N_12513,N_12557);
and U12662 (N_12662,N_12427,N_12348);
xnor U12663 (N_12663,N_12531,N_12391);
nand U12664 (N_12664,N_12314,N_12409);
nand U12665 (N_12665,N_12476,N_12301);
or U12666 (N_12666,N_12463,N_12478);
and U12667 (N_12667,N_12424,N_12322);
nand U12668 (N_12668,N_12520,N_12320);
nor U12669 (N_12669,N_12558,N_12403);
or U12670 (N_12670,N_12453,N_12488);
and U12671 (N_12671,N_12355,N_12415);
or U12672 (N_12672,N_12372,N_12458);
or U12673 (N_12673,N_12517,N_12581);
nor U12674 (N_12674,N_12304,N_12311);
nor U12675 (N_12675,N_12585,N_12508);
nand U12676 (N_12676,N_12444,N_12552);
or U12677 (N_12677,N_12389,N_12539);
xnor U12678 (N_12678,N_12360,N_12571);
and U12679 (N_12679,N_12445,N_12398);
nand U12680 (N_12680,N_12425,N_12546);
nor U12681 (N_12681,N_12502,N_12553);
nor U12682 (N_12682,N_12400,N_12370);
nand U12683 (N_12683,N_12479,N_12569);
nor U12684 (N_12684,N_12493,N_12567);
nand U12685 (N_12685,N_12303,N_12562);
or U12686 (N_12686,N_12515,N_12510);
and U12687 (N_12687,N_12450,N_12429);
nand U12688 (N_12688,N_12340,N_12525);
nand U12689 (N_12689,N_12353,N_12364);
nand U12690 (N_12690,N_12466,N_12535);
or U12691 (N_12691,N_12317,N_12576);
xnor U12692 (N_12692,N_12361,N_12498);
or U12693 (N_12693,N_12385,N_12344);
nand U12694 (N_12694,N_12473,N_12359);
or U12695 (N_12695,N_12392,N_12543);
nor U12696 (N_12696,N_12383,N_12595);
nor U12697 (N_12697,N_12332,N_12457);
or U12698 (N_12698,N_12451,N_12480);
or U12699 (N_12699,N_12524,N_12346);
or U12700 (N_12700,N_12417,N_12326);
xor U12701 (N_12701,N_12347,N_12464);
nor U12702 (N_12702,N_12441,N_12528);
and U12703 (N_12703,N_12465,N_12533);
nand U12704 (N_12704,N_12486,N_12341);
and U12705 (N_12705,N_12518,N_12474);
nor U12706 (N_12706,N_12423,N_12494);
nand U12707 (N_12707,N_12397,N_12499);
xnor U12708 (N_12708,N_12501,N_12371);
or U12709 (N_12709,N_12522,N_12523);
or U12710 (N_12710,N_12428,N_12532);
or U12711 (N_12711,N_12594,N_12544);
or U12712 (N_12712,N_12438,N_12382);
or U12713 (N_12713,N_12404,N_12540);
nand U12714 (N_12714,N_12496,N_12343);
or U12715 (N_12715,N_12487,N_12497);
nand U12716 (N_12716,N_12329,N_12395);
or U12717 (N_12717,N_12505,N_12414);
xor U12718 (N_12718,N_12572,N_12555);
nor U12719 (N_12719,N_12342,N_12313);
or U12720 (N_12720,N_12407,N_12583);
or U12721 (N_12721,N_12477,N_12563);
or U12722 (N_12722,N_12316,N_12337);
nand U12723 (N_12723,N_12542,N_12534);
and U12724 (N_12724,N_12399,N_12526);
nor U12725 (N_12725,N_12386,N_12349);
nand U12726 (N_12726,N_12573,N_12564);
or U12727 (N_12727,N_12489,N_12504);
nand U12728 (N_12728,N_12452,N_12327);
and U12729 (N_12729,N_12384,N_12367);
or U12730 (N_12730,N_12560,N_12548);
nor U12731 (N_12731,N_12586,N_12545);
xor U12732 (N_12732,N_12467,N_12541);
nor U12733 (N_12733,N_12588,N_12521);
xnor U12734 (N_12734,N_12460,N_12394);
and U12735 (N_12735,N_12507,N_12527);
xnor U12736 (N_12736,N_12308,N_12416);
nor U12737 (N_12737,N_12584,N_12578);
nor U12738 (N_12738,N_12379,N_12549);
or U12739 (N_12739,N_12470,N_12430);
nand U12740 (N_12740,N_12482,N_12381);
xor U12741 (N_12741,N_12537,N_12575);
nand U12742 (N_12742,N_12506,N_12388);
and U12743 (N_12743,N_12565,N_12378);
xnor U12744 (N_12744,N_12309,N_12446);
xor U12745 (N_12745,N_12442,N_12324);
and U12746 (N_12746,N_12550,N_12369);
or U12747 (N_12747,N_12519,N_12556);
or U12748 (N_12748,N_12307,N_12529);
nand U12749 (N_12749,N_12302,N_12547);
nand U12750 (N_12750,N_12440,N_12304);
nand U12751 (N_12751,N_12395,N_12310);
nor U12752 (N_12752,N_12511,N_12322);
or U12753 (N_12753,N_12323,N_12331);
nand U12754 (N_12754,N_12413,N_12336);
nand U12755 (N_12755,N_12565,N_12431);
nor U12756 (N_12756,N_12408,N_12526);
nand U12757 (N_12757,N_12391,N_12339);
and U12758 (N_12758,N_12315,N_12591);
nor U12759 (N_12759,N_12407,N_12420);
and U12760 (N_12760,N_12395,N_12505);
nor U12761 (N_12761,N_12439,N_12519);
nor U12762 (N_12762,N_12572,N_12403);
or U12763 (N_12763,N_12599,N_12452);
nand U12764 (N_12764,N_12597,N_12385);
nor U12765 (N_12765,N_12419,N_12347);
nor U12766 (N_12766,N_12531,N_12517);
nor U12767 (N_12767,N_12411,N_12358);
nand U12768 (N_12768,N_12511,N_12429);
xnor U12769 (N_12769,N_12413,N_12572);
or U12770 (N_12770,N_12428,N_12517);
nor U12771 (N_12771,N_12507,N_12373);
and U12772 (N_12772,N_12320,N_12586);
nor U12773 (N_12773,N_12589,N_12597);
nor U12774 (N_12774,N_12576,N_12556);
or U12775 (N_12775,N_12317,N_12343);
nor U12776 (N_12776,N_12431,N_12328);
or U12777 (N_12777,N_12509,N_12549);
nor U12778 (N_12778,N_12345,N_12450);
or U12779 (N_12779,N_12311,N_12393);
and U12780 (N_12780,N_12565,N_12596);
or U12781 (N_12781,N_12536,N_12592);
nor U12782 (N_12782,N_12457,N_12543);
and U12783 (N_12783,N_12567,N_12432);
nand U12784 (N_12784,N_12584,N_12573);
xor U12785 (N_12785,N_12477,N_12486);
and U12786 (N_12786,N_12533,N_12436);
nor U12787 (N_12787,N_12414,N_12534);
or U12788 (N_12788,N_12363,N_12485);
or U12789 (N_12789,N_12415,N_12495);
and U12790 (N_12790,N_12446,N_12556);
or U12791 (N_12791,N_12464,N_12337);
or U12792 (N_12792,N_12531,N_12456);
xor U12793 (N_12793,N_12587,N_12318);
nand U12794 (N_12794,N_12458,N_12302);
or U12795 (N_12795,N_12341,N_12378);
nor U12796 (N_12796,N_12581,N_12552);
or U12797 (N_12797,N_12407,N_12502);
or U12798 (N_12798,N_12450,N_12549);
and U12799 (N_12799,N_12444,N_12467);
nor U12800 (N_12800,N_12599,N_12304);
nor U12801 (N_12801,N_12369,N_12405);
nor U12802 (N_12802,N_12331,N_12450);
and U12803 (N_12803,N_12350,N_12345);
nand U12804 (N_12804,N_12582,N_12449);
and U12805 (N_12805,N_12458,N_12571);
or U12806 (N_12806,N_12471,N_12361);
xor U12807 (N_12807,N_12542,N_12363);
xnor U12808 (N_12808,N_12477,N_12420);
or U12809 (N_12809,N_12505,N_12478);
or U12810 (N_12810,N_12561,N_12505);
and U12811 (N_12811,N_12531,N_12523);
nand U12812 (N_12812,N_12447,N_12592);
or U12813 (N_12813,N_12335,N_12553);
nor U12814 (N_12814,N_12530,N_12571);
xnor U12815 (N_12815,N_12412,N_12311);
nand U12816 (N_12816,N_12465,N_12392);
xor U12817 (N_12817,N_12325,N_12493);
xnor U12818 (N_12818,N_12588,N_12412);
nand U12819 (N_12819,N_12534,N_12334);
xnor U12820 (N_12820,N_12415,N_12340);
and U12821 (N_12821,N_12317,N_12592);
and U12822 (N_12822,N_12476,N_12354);
nor U12823 (N_12823,N_12414,N_12427);
and U12824 (N_12824,N_12497,N_12594);
and U12825 (N_12825,N_12496,N_12428);
and U12826 (N_12826,N_12343,N_12351);
nand U12827 (N_12827,N_12473,N_12385);
xor U12828 (N_12828,N_12452,N_12415);
xnor U12829 (N_12829,N_12569,N_12598);
or U12830 (N_12830,N_12515,N_12411);
and U12831 (N_12831,N_12571,N_12341);
and U12832 (N_12832,N_12354,N_12358);
and U12833 (N_12833,N_12430,N_12332);
nand U12834 (N_12834,N_12329,N_12422);
nand U12835 (N_12835,N_12561,N_12410);
nor U12836 (N_12836,N_12488,N_12423);
or U12837 (N_12837,N_12576,N_12488);
and U12838 (N_12838,N_12453,N_12317);
and U12839 (N_12839,N_12575,N_12579);
or U12840 (N_12840,N_12404,N_12432);
xor U12841 (N_12841,N_12556,N_12590);
nor U12842 (N_12842,N_12546,N_12585);
xnor U12843 (N_12843,N_12593,N_12511);
or U12844 (N_12844,N_12566,N_12364);
and U12845 (N_12845,N_12491,N_12489);
xor U12846 (N_12846,N_12394,N_12504);
and U12847 (N_12847,N_12501,N_12411);
and U12848 (N_12848,N_12452,N_12331);
nand U12849 (N_12849,N_12375,N_12518);
nand U12850 (N_12850,N_12491,N_12487);
xnor U12851 (N_12851,N_12556,N_12326);
or U12852 (N_12852,N_12402,N_12397);
and U12853 (N_12853,N_12392,N_12405);
nor U12854 (N_12854,N_12425,N_12426);
or U12855 (N_12855,N_12524,N_12443);
xnor U12856 (N_12856,N_12440,N_12540);
or U12857 (N_12857,N_12406,N_12523);
or U12858 (N_12858,N_12328,N_12376);
and U12859 (N_12859,N_12339,N_12346);
or U12860 (N_12860,N_12395,N_12581);
or U12861 (N_12861,N_12328,N_12521);
nand U12862 (N_12862,N_12320,N_12527);
nand U12863 (N_12863,N_12589,N_12451);
or U12864 (N_12864,N_12521,N_12575);
nor U12865 (N_12865,N_12476,N_12496);
nor U12866 (N_12866,N_12472,N_12401);
xor U12867 (N_12867,N_12570,N_12367);
nand U12868 (N_12868,N_12334,N_12462);
or U12869 (N_12869,N_12382,N_12450);
nor U12870 (N_12870,N_12522,N_12419);
nand U12871 (N_12871,N_12469,N_12558);
nand U12872 (N_12872,N_12580,N_12484);
or U12873 (N_12873,N_12310,N_12387);
xnor U12874 (N_12874,N_12316,N_12572);
and U12875 (N_12875,N_12372,N_12349);
or U12876 (N_12876,N_12426,N_12508);
nand U12877 (N_12877,N_12340,N_12428);
nand U12878 (N_12878,N_12393,N_12580);
and U12879 (N_12879,N_12382,N_12491);
nor U12880 (N_12880,N_12560,N_12484);
nand U12881 (N_12881,N_12401,N_12544);
or U12882 (N_12882,N_12375,N_12587);
xnor U12883 (N_12883,N_12303,N_12505);
and U12884 (N_12884,N_12533,N_12405);
and U12885 (N_12885,N_12369,N_12501);
or U12886 (N_12886,N_12559,N_12427);
xnor U12887 (N_12887,N_12406,N_12390);
nor U12888 (N_12888,N_12374,N_12457);
nor U12889 (N_12889,N_12316,N_12595);
and U12890 (N_12890,N_12425,N_12564);
xor U12891 (N_12891,N_12546,N_12593);
nor U12892 (N_12892,N_12515,N_12520);
xor U12893 (N_12893,N_12405,N_12326);
xor U12894 (N_12894,N_12586,N_12531);
xnor U12895 (N_12895,N_12364,N_12571);
nor U12896 (N_12896,N_12548,N_12572);
and U12897 (N_12897,N_12337,N_12422);
and U12898 (N_12898,N_12549,N_12503);
nor U12899 (N_12899,N_12551,N_12562);
nand U12900 (N_12900,N_12845,N_12709);
or U12901 (N_12901,N_12753,N_12648);
xor U12902 (N_12902,N_12713,N_12768);
and U12903 (N_12903,N_12803,N_12838);
xnor U12904 (N_12904,N_12862,N_12836);
xnor U12905 (N_12905,N_12815,N_12766);
and U12906 (N_12906,N_12634,N_12851);
and U12907 (N_12907,N_12623,N_12647);
and U12908 (N_12908,N_12805,N_12692);
and U12909 (N_12909,N_12624,N_12777);
nor U12910 (N_12910,N_12716,N_12835);
xor U12911 (N_12911,N_12846,N_12849);
and U12912 (N_12912,N_12797,N_12744);
nor U12913 (N_12913,N_12730,N_12725);
and U12914 (N_12914,N_12787,N_12733);
nor U12915 (N_12915,N_12834,N_12617);
nand U12916 (N_12916,N_12873,N_12652);
or U12917 (N_12917,N_12664,N_12636);
nor U12918 (N_12918,N_12656,N_12706);
and U12919 (N_12919,N_12635,N_12813);
nor U12920 (N_12920,N_12864,N_12653);
and U12921 (N_12921,N_12602,N_12764);
or U12922 (N_12922,N_12823,N_12639);
nand U12923 (N_12923,N_12893,N_12760);
and U12924 (N_12924,N_12681,N_12609);
nand U12925 (N_12925,N_12798,N_12612);
or U12926 (N_12926,N_12689,N_12734);
nor U12927 (N_12927,N_12640,N_12847);
nor U12928 (N_12928,N_12743,N_12742);
xnor U12929 (N_12929,N_12718,N_12699);
xnor U12930 (N_12930,N_12691,N_12765);
nand U12931 (N_12931,N_12898,N_12857);
nor U12932 (N_12932,N_12806,N_12606);
xor U12933 (N_12933,N_12605,N_12723);
nor U12934 (N_12934,N_12858,N_12831);
or U12935 (N_12935,N_12795,N_12601);
and U12936 (N_12936,N_12745,N_12661);
nor U12937 (N_12937,N_12790,N_12679);
or U12938 (N_12938,N_12626,N_12702);
and U12939 (N_12939,N_12868,N_12613);
or U12940 (N_12940,N_12735,N_12822);
or U12941 (N_12941,N_12750,N_12856);
nand U12942 (N_12942,N_12839,N_12881);
nand U12943 (N_12943,N_12837,N_12774);
nor U12944 (N_12944,N_12708,N_12872);
and U12945 (N_12945,N_12791,N_12841);
nand U12946 (N_12946,N_12759,N_12801);
or U12947 (N_12947,N_12603,N_12625);
nor U12948 (N_12948,N_12853,N_12789);
nand U12949 (N_12949,N_12818,N_12794);
and U12950 (N_12950,N_12659,N_12869);
nor U12951 (N_12951,N_12894,N_12642);
xor U12952 (N_12952,N_12690,N_12761);
xnor U12953 (N_12953,N_12863,N_12663);
or U12954 (N_12954,N_12871,N_12649);
nor U12955 (N_12955,N_12855,N_12678);
nor U12956 (N_12956,N_12781,N_12804);
or U12957 (N_12957,N_12828,N_12891);
or U12958 (N_12958,N_12703,N_12695);
xor U12959 (N_12959,N_12683,N_12719);
nand U12960 (N_12960,N_12641,N_12687);
and U12961 (N_12961,N_12820,N_12756);
and U12962 (N_12962,N_12680,N_12608);
and U12963 (N_12963,N_12704,N_12650);
or U12964 (N_12964,N_12767,N_12645);
nand U12965 (N_12965,N_12827,N_12840);
nor U12966 (N_12966,N_12693,N_12694);
or U12967 (N_12967,N_12769,N_12630);
xor U12968 (N_12968,N_12685,N_12620);
and U12969 (N_12969,N_12728,N_12779);
xnor U12970 (N_12970,N_12877,N_12727);
nand U12971 (N_12971,N_12722,N_12721);
or U12972 (N_12972,N_12758,N_12772);
xor U12973 (N_12973,N_12657,N_12705);
nand U12974 (N_12974,N_12684,N_12665);
or U12975 (N_12975,N_12622,N_12786);
and U12976 (N_12976,N_12701,N_12780);
and U12977 (N_12977,N_12671,N_12668);
nand U12978 (N_12978,N_12829,N_12682);
nor U12979 (N_12979,N_12778,N_12658);
and U12980 (N_12980,N_12763,N_12866);
nor U12981 (N_12981,N_12771,N_12707);
xor U12982 (N_12982,N_12850,N_12631);
xor U12983 (N_12983,N_12646,N_12710);
nor U12984 (N_12984,N_12875,N_12809);
or U12985 (N_12985,N_12812,N_12627);
or U12986 (N_12986,N_12654,N_12715);
nor U12987 (N_12987,N_12825,N_12770);
nor U12988 (N_12988,N_12852,N_12662);
xnor U12989 (N_12989,N_12886,N_12824);
nand U12990 (N_12990,N_12633,N_12861);
or U12991 (N_12991,N_12638,N_12666);
nor U12992 (N_12992,N_12669,N_12629);
nand U12993 (N_12993,N_12783,N_12688);
or U12994 (N_12994,N_12667,N_12832);
and U12995 (N_12995,N_12843,N_12773);
or U12996 (N_12996,N_12746,N_12878);
nand U12997 (N_12997,N_12632,N_12614);
and U12998 (N_12998,N_12738,N_12736);
nor U12999 (N_12999,N_12802,N_12740);
nor U13000 (N_13000,N_12616,N_12782);
nand U13001 (N_13001,N_12888,N_12628);
nand U13002 (N_13002,N_12830,N_12672);
nand U13003 (N_13003,N_12890,N_12615);
and U13004 (N_13004,N_12749,N_12887);
xnor U13005 (N_13005,N_12810,N_12848);
nand U13006 (N_13006,N_12676,N_12660);
nor U13007 (N_13007,N_12619,N_12885);
and U13008 (N_13008,N_12607,N_12842);
nand U13009 (N_13009,N_12816,N_12747);
or U13010 (N_13010,N_12686,N_12826);
nor U13011 (N_13011,N_12754,N_12712);
nand U13012 (N_13012,N_12817,N_12610);
and U13013 (N_13013,N_12819,N_12844);
nand U13014 (N_13014,N_12739,N_12698);
or U13015 (N_13015,N_12882,N_12755);
or U13016 (N_13016,N_12611,N_12618);
xnor U13017 (N_13017,N_12697,N_12673);
nor U13018 (N_13018,N_12892,N_12860);
nand U13019 (N_13019,N_12762,N_12800);
nand U13020 (N_13020,N_12883,N_12833);
xor U13021 (N_13021,N_12784,N_12600);
and U13022 (N_13022,N_12811,N_12876);
or U13023 (N_13023,N_12896,N_12859);
nor U13024 (N_13024,N_12732,N_12655);
xor U13025 (N_13025,N_12788,N_12821);
nor U13026 (N_13026,N_12895,N_12731);
and U13027 (N_13027,N_12865,N_12899);
and U13028 (N_13028,N_12696,N_12889);
nand U13029 (N_13029,N_12670,N_12621);
nor U13030 (N_13030,N_12677,N_12751);
nor U13031 (N_13031,N_12752,N_12793);
xnor U13032 (N_13032,N_12757,N_12748);
nor U13033 (N_13033,N_12729,N_12674);
and U13034 (N_13034,N_12741,N_12799);
xor U13035 (N_13035,N_12808,N_12796);
and U13036 (N_13036,N_12714,N_12637);
nor U13037 (N_13037,N_12700,N_12724);
nand U13038 (N_13038,N_12737,N_12814);
nand U13039 (N_13039,N_12792,N_12776);
nand U13040 (N_13040,N_12854,N_12807);
and U13041 (N_13041,N_12874,N_12651);
or U13042 (N_13042,N_12897,N_12775);
xor U13043 (N_13043,N_12720,N_12879);
or U13044 (N_13044,N_12717,N_12726);
xnor U13045 (N_13045,N_12644,N_12884);
nand U13046 (N_13046,N_12711,N_12867);
and U13047 (N_13047,N_12604,N_12870);
or U13048 (N_13048,N_12675,N_12643);
or U13049 (N_13049,N_12880,N_12785);
nor U13050 (N_13050,N_12784,N_12783);
nor U13051 (N_13051,N_12615,N_12878);
xnor U13052 (N_13052,N_12723,N_12766);
and U13053 (N_13053,N_12611,N_12638);
and U13054 (N_13054,N_12653,N_12710);
or U13055 (N_13055,N_12871,N_12633);
nand U13056 (N_13056,N_12704,N_12608);
or U13057 (N_13057,N_12767,N_12656);
and U13058 (N_13058,N_12812,N_12879);
and U13059 (N_13059,N_12843,N_12814);
nand U13060 (N_13060,N_12616,N_12676);
and U13061 (N_13061,N_12620,N_12659);
and U13062 (N_13062,N_12659,N_12653);
and U13063 (N_13063,N_12715,N_12712);
or U13064 (N_13064,N_12867,N_12797);
xnor U13065 (N_13065,N_12865,N_12673);
and U13066 (N_13066,N_12768,N_12731);
xor U13067 (N_13067,N_12604,N_12790);
nor U13068 (N_13068,N_12799,N_12899);
nor U13069 (N_13069,N_12898,N_12770);
nand U13070 (N_13070,N_12882,N_12634);
and U13071 (N_13071,N_12842,N_12828);
and U13072 (N_13072,N_12826,N_12873);
xor U13073 (N_13073,N_12636,N_12852);
nor U13074 (N_13074,N_12626,N_12745);
and U13075 (N_13075,N_12635,N_12702);
or U13076 (N_13076,N_12875,N_12651);
nor U13077 (N_13077,N_12753,N_12625);
xnor U13078 (N_13078,N_12837,N_12714);
nand U13079 (N_13079,N_12804,N_12611);
nor U13080 (N_13080,N_12621,N_12742);
and U13081 (N_13081,N_12680,N_12652);
and U13082 (N_13082,N_12725,N_12629);
nor U13083 (N_13083,N_12735,N_12763);
nand U13084 (N_13084,N_12760,N_12701);
nand U13085 (N_13085,N_12888,N_12854);
and U13086 (N_13086,N_12629,N_12859);
and U13087 (N_13087,N_12791,N_12834);
nand U13088 (N_13088,N_12812,N_12632);
or U13089 (N_13089,N_12822,N_12824);
nand U13090 (N_13090,N_12634,N_12798);
and U13091 (N_13091,N_12713,N_12813);
nor U13092 (N_13092,N_12669,N_12603);
nand U13093 (N_13093,N_12718,N_12655);
nand U13094 (N_13094,N_12869,N_12890);
nor U13095 (N_13095,N_12832,N_12807);
nor U13096 (N_13096,N_12777,N_12674);
nor U13097 (N_13097,N_12759,N_12677);
or U13098 (N_13098,N_12775,N_12623);
nor U13099 (N_13099,N_12898,N_12859);
or U13100 (N_13100,N_12689,N_12853);
xnor U13101 (N_13101,N_12601,N_12605);
and U13102 (N_13102,N_12627,N_12806);
nor U13103 (N_13103,N_12791,N_12764);
and U13104 (N_13104,N_12660,N_12847);
or U13105 (N_13105,N_12703,N_12762);
nor U13106 (N_13106,N_12750,N_12731);
nor U13107 (N_13107,N_12689,N_12825);
nor U13108 (N_13108,N_12677,N_12778);
or U13109 (N_13109,N_12682,N_12723);
xor U13110 (N_13110,N_12722,N_12671);
nand U13111 (N_13111,N_12655,N_12700);
and U13112 (N_13112,N_12762,N_12645);
nor U13113 (N_13113,N_12749,N_12837);
or U13114 (N_13114,N_12739,N_12747);
nand U13115 (N_13115,N_12851,N_12826);
xnor U13116 (N_13116,N_12847,N_12727);
and U13117 (N_13117,N_12724,N_12832);
and U13118 (N_13118,N_12673,N_12758);
nor U13119 (N_13119,N_12816,N_12661);
nor U13120 (N_13120,N_12632,N_12854);
nand U13121 (N_13121,N_12876,N_12707);
nand U13122 (N_13122,N_12757,N_12775);
nand U13123 (N_13123,N_12827,N_12717);
nand U13124 (N_13124,N_12645,N_12674);
xor U13125 (N_13125,N_12881,N_12669);
nand U13126 (N_13126,N_12805,N_12887);
xnor U13127 (N_13127,N_12897,N_12729);
nor U13128 (N_13128,N_12879,N_12896);
nor U13129 (N_13129,N_12672,N_12625);
or U13130 (N_13130,N_12797,N_12782);
or U13131 (N_13131,N_12672,N_12693);
xor U13132 (N_13132,N_12620,N_12693);
xnor U13133 (N_13133,N_12663,N_12783);
nor U13134 (N_13134,N_12711,N_12694);
and U13135 (N_13135,N_12785,N_12772);
and U13136 (N_13136,N_12607,N_12663);
nand U13137 (N_13137,N_12714,N_12720);
xnor U13138 (N_13138,N_12826,N_12892);
or U13139 (N_13139,N_12607,N_12669);
and U13140 (N_13140,N_12656,N_12822);
and U13141 (N_13141,N_12663,N_12626);
nor U13142 (N_13142,N_12838,N_12852);
nor U13143 (N_13143,N_12801,N_12683);
nor U13144 (N_13144,N_12717,N_12852);
nand U13145 (N_13145,N_12619,N_12817);
nor U13146 (N_13146,N_12852,N_12837);
nand U13147 (N_13147,N_12687,N_12703);
nor U13148 (N_13148,N_12610,N_12864);
nand U13149 (N_13149,N_12675,N_12647);
or U13150 (N_13150,N_12633,N_12660);
and U13151 (N_13151,N_12897,N_12618);
nand U13152 (N_13152,N_12615,N_12832);
or U13153 (N_13153,N_12678,N_12872);
and U13154 (N_13154,N_12705,N_12881);
nand U13155 (N_13155,N_12806,N_12717);
or U13156 (N_13156,N_12807,N_12611);
or U13157 (N_13157,N_12732,N_12666);
nand U13158 (N_13158,N_12771,N_12690);
and U13159 (N_13159,N_12813,N_12731);
nor U13160 (N_13160,N_12849,N_12894);
and U13161 (N_13161,N_12762,N_12712);
nand U13162 (N_13162,N_12681,N_12871);
or U13163 (N_13163,N_12696,N_12603);
or U13164 (N_13164,N_12660,N_12850);
or U13165 (N_13165,N_12831,N_12739);
and U13166 (N_13166,N_12655,N_12806);
or U13167 (N_13167,N_12791,N_12895);
nand U13168 (N_13168,N_12665,N_12657);
and U13169 (N_13169,N_12895,N_12693);
and U13170 (N_13170,N_12820,N_12784);
xnor U13171 (N_13171,N_12813,N_12788);
xnor U13172 (N_13172,N_12848,N_12786);
xnor U13173 (N_13173,N_12828,N_12884);
nor U13174 (N_13174,N_12721,N_12803);
and U13175 (N_13175,N_12739,N_12736);
nand U13176 (N_13176,N_12815,N_12639);
xnor U13177 (N_13177,N_12840,N_12752);
and U13178 (N_13178,N_12768,N_12892);
nand U13179 (N_13179,N_12825,N_12659);
and U13180 (N_13180,N_12743,N_12753);
xnor U13181 (N_13181,N_12850,N_12855);
xor U13182 (N_13182,N_12819,N_12899);
nand U13183 (N_13183,N_12735,N_12740);
and U13184 (N_13184,N_12621,N_12760);
or U13185 (N_13185,N_12679,N_12773);
nor U13186 (N_13186,N_12815,N_12855);
nand U13187 (N_13187,N_12643,N_12703);
and U13188 (N_13188,N_12789,N_12762);
or U13189 (N_13189,N_12725,N_12862);
nand U13190 (N_13190,N_12655,N_12640);
nor U13191 (N_13191,N_12844,N_12733);
nor U13192 (N_13192,N_12842,N_12884);
or U13193 (N_13193,N_12659,N_12602);
xnor U13194 (N_13194,N_12833,N_12832);
nand U13195 (N_13195,N_12707,N_12693);
or U13196 (N_13196,N_12739,N_12682);
or U13197 (N_13197,N_12884,N_12862);
or U13198 (N_13198,N_12860,N_12778);
nor U13199 (N_13199,N_12628,N_12690);
nand U13200 (N_13200,N_13095,N_12902);
and U13201 (N_13201,N_12900,N_13103);
nor U13202 (N_13202,N_13014,N_13017);
and U13203 (N_13203,N_13078,N_13054);
and U13204 (N_13204,N_13036,N_12981);
and U13205 (N_13205,N_13172,N_13148);
nor U13206 (N_13206,N_12976,N_13004);
or U13207 (N_13207,N_13030,N_13191);
and U13208 (N_13208,N_13114,N_12954);
xnor U13209 (N_13209,N_13021,N_13136);
nand U13210 (N_13210,N_12987,N_12946);
and U13211 (N_13211,N_13049,N_13129);
xor U13212 (N_13212,N_13174,N_13074);
nor U13213 (N_13213,N_13016,N_13052);
xnor U13214 (N_13214,N_12940,N_12982);
nor U13215 (N_13215,N_13150,N_13183);
xnor U13216 (N_13216,N_13090,N_13112);
and U13217 (N_13217,N_12989,N_13110);
nor U13218 (N_13218,N_13029,N_13080);
nand U13219 (N_13219,N_12991,N_13087);
nor U13220 (N_13220,N_13138,N_13184);
or U13221 (N_13221,N_13012,N_13135);
or U13222 (N_13222,N_13157,N_12959);
or U13223 (N_13223,N_13194,N_12917);
or U13224 (N_13224,N_13193,N_13145);
xnor U13225 (N_13225,N_13189,N_13108);
nand U13226 (N_13226,N_13062,N_12951);
or U13227 (N_13227,N_13180,N_13038);
nand U13228 (N_13228,N_12903,N_13133);
and U13229 (N_13229,N_12968,N_12980);
xor U13230 (N_13230,N_13175,N_13072);
nor U13231 (N_13231,N_12908,N_12979);
or U13232 (N_13232,N_12935,N_13130);
nor U13233 (N_13233,N_13040,N_13031);
or U13234 (N_13234,N_13067,N_13056);
and U13235 (N_13235,N_13020,N_12911);
nor U13236 (N_13236,N_13161,N_13117);
or U13237 (N_13237,N_12969,N_12945);
xor U13238 (N_13238,N_13064,N_13026);
or U13239 (N_13239,N_12921,N_13005);
and U13240 (N_13240,N_12997,N_12985);
and U13241 (N_13241,N_13053,N_12922);
and U13242 (N_13242,N_13085,N_12933);
or U13243 (N_13243,N_13088,N_13164);
or U13244 (N_13244,N_13034,N_12942);
xnor U13245 (N_13245,N_12961,N_13097);
and U13246 (N_13246,N_13007,N_12978);
or U13247 (N_13247,N_13028,N_13094);
nor U13248 (N_13248,N_12960,N_13156);
or U13249 (N_13249,N_12926,N_13141);
xnor U13250 (N_13250,N_12970,N_13107);
nand U13251 (N_13251,N_13185,N_12994);
xnor U13252 (N_13252,N_13155,N_13122);
xnor U13253 (N_13253,N_13023,N_13058);
xnor U13254 (N_13254,N_12918,N_13163);
xnor U13255 (N_13255,N_12962,N_13001);
xor U13256 (N_13256,N_13153,N_13105);
or U13257 (N_13257,N_13169,N_13042);
or U13258 (N_13258,N_13027,N_12986);
and U13259 (N_13259,N_13000,N_13082);
xnor U13260 (N_13260,N_12957,N_12958);
and U13261 (N_13261,N_13166,N_13162);
xor U13262 (N_13262,N_13176,N_12913);
nand U13263 (N_13263,N_13069,N_13048);
or U13264 (N_13264,N_13178,N_13143);
nand U13265 (N_13265,N_13009,N_13065);
nor U13266 (N_13266,N_13102,N_12936);
nor U13267 (N_13267,N_13081,N_13154);
nand U13268 (N_13268,N_12906,N_13137);
nand U13269 (N_13269,N_13010,N_12929);
and U13270 (N_13270,N_12924,N_13181);
xor U13271 (N_13271,N_13131,N_12905);
or U13272 (N_13272,N_12931,N_13177);
nor U13273 (N_13273,N_13077,N_13170);
and U13274 (N_13274,N_13047,N_13092);
nand U13275 (N_13275,N_13116,N_13091);
xor U13276 (N_13276,N_13195,N_13199);
or U13277 (N_13277,N_12938,N_12914);
xor U13278 (N_13278,N_13043,N_13096);
nand U13279 (N_13279,N_12920,N_13147);
xor U13280 (N_13280,N_12919,N_12955);
or U13281 (N_13281,N_12965,N_13139);
nand U13282 (N_13282,N_13119,N_12901);
or U13283 (N_13283,N_13011,N_13025);
nor U13284 (N_13284,N_12993,N_12996);
or U13285 (N_13285,N_13120,N_13035);
xnor U13286 (N_13286,N_12964,N_13073);
and U13287 (N_13287,N_12998,N_13186);
nand U13288 (N_13288,N_13152,N_13046);
and U13289 (N_13289,N_13086,N_12925);
nor U13290 (N_13290,N_13093,N_12948);
or U13291 (N_13291,N_13041,N_12947);
nand U13292 (N_13292,N_13167,N_13075);
nor U13293 (N_13293,N_13124,N_12930);
xor U13294 (N_13294,N_13101,N_13179);
nand U13295 (N_13295,N_12963,N_13061);
and U13296 (N_13296,N_12988,N_13063);
or U13297 (N_13297,N_13019,N_13160);
nor U13298 (N_13298,N_13018,N_13118);
nor U13299 (N_13299,N_12973,N_13050);
xnor U13300 (N_13300,N_13057,N_13008);
xnor U13301 (N_13301,N_13151,N_12952);
and U13302 (N_13302,N_13100,N_13099);
and U13303 (N_13303,N_13198,N_13127);
and U13304 (N_13304,N_13128,N_12923);
or U13305 (N_13305,N_13089,N_12916);
nor U13306 (N_13306,N_12912,N_13168);
and U13307 (N_13307,N_12977,N_13051);
nor U13308 (N_13308,N_13071,N_13146);
xor U13309 (N_13309,N_12944,N_12984);
nand U13310 (N_13310,N_12995,N_13002);
nor U13311 (N_13311,N_12967,N_13190);
and U13312 (N_13312,N_13188,N_13076);
or U13313 (N_13313,N_13192,N_13125);
xnor U13314 (N_13314,N_13165,N_13111);
xnor U13315 (N_13315,N_12974,N_13032);
and U13316 (N_13316,N_13144,N_13134);
nand U13317 (N_13317,N_12943,N_13171);
nand U13318 (N_13318,N_13113,N_12904);
nor U13319 (N_13319,N_13003,N_13055);
xor U13320 (N_13320,N_13182,N_12950);
xnor U13321 (N_13321,N_12907,N_13060);
or U13322 (N_13322,N_13142,N_12999);
nand U13323 (N_13323,N_12915,N_13013);
or U13324 (N_13324,N_12975,N_12990);
nor U13325 (N_13325,N_12953,N_13037);
and U13326 (N_13326,N_13098,N_13132);
nor U13327 (N_13327,N_13115,N_13196);
xor U13328 (N_13328,N_13158,N_13173);
or U13329 (N_13329,N_12966,N_13044);
or U13330 (N_13330,N_12971,N_13084);
and U13331 (N_13331,N_12927,N_12910);
nor U13332 (N_13332,N_13033,N_13159);
xnor U13333 (N_13333,N_13022,N_12941);
nor U13334 (N_13334,N_12949,N_13121);
nand U13335 (N_13335,N_13083,N_13070);
nand U13336 (N_13336,N_13079,N_12992);
or U13337 (N_13337,N_12909,N_13104);
xor U13338 (N_13338,N_13123,N_13126);
or U13339 (N_13339,N_13015,N_13024);
nor U13340 (N_13340,N_13045,N_13066);
and U13341 (N_13341,N_12932,N_13140);
xor U13342 (N_13342,N_12934,N_12928);
nor U13343 (N_13343,N_12939,N_13109);
nand U13344 (N_13344,N_13106,N_12983);
nor U13345 (N_13345,N_13068,N_12956);
or U13346 (N_13346,N_13006,N_13197);
and U13347 (N_13347,N_13149,N_12937);
nand U13348 (N_13348,N_13039,N_12972);
and U13349 (N_13349,N_13059,N_13187);
or U13350 (N_13350,N_13050,N_13021);
xor U13351 (N_13351,N_13058,N_12905);
nor U13352 (N_13352,N_12944,N_12965);
nor U13353 (N_13353,N_12907,N_12920);
nand U13354 (N_13354,N_13023,N_12903);
and U13355 (N_13355,N_13165,N_13010);
nand U13356 (N_13356,N_13136,N_13197);
and U13357 (N_13357,N_13157,N_12937);
nor U13358 (N_13358,N_13001,N_12988);
xor U13359 (N_13359,N_13090,N_13022);
nand U13360 (N_13360,N_12956,N_13043);
or U13361 (N_13361,N_13149,N_12956);
or U13362 (N_13362,N_13069,N_13193);
xor U13363 (N_13363,N_13155,N_13046);
xor U13364 (N_13364,N_12955,N_13044);
and U13365 (N_13365,N_12939,N_12906);
and U13366 (N_13366,N_12915,N_13071);
xor U13367 (N_13367,N_12950,N_13156);
xnor U13368 (N_13368,N_12983,N_13090);
or U13369 (N_13369,N_13177,N_13131);
or U13370 (N_13370,N_13053,N_13026);
or U13371 (N_13371,N_13024,N_13034);
and U13372 (N_13372,N_13087,N_12915);
nor U13373 (N_13373,N_13178,N_13006);
and U13374 (N_13374,N_12937,N_12967);
and U13375 (N_13375,N_12913,N_13197);
xnor U13376 (N_13376,N_13125,N_12900);
xor U13377 (N_13377,N_13111,N_13099);
or U13378 (N_13378,N_12981,N_13048);
xor U13379 (N_13379,N_12954,N_12904);
and U13380 (N_13380,N_13114,N_12958);
or U13381 (N_13381,N_13111,N_12947);
or U13382 (N_13382,N_13096,N_13081);
nand U13383 (N_13383,N_13105,N_13022);
and U13384 (N_13384,N_12944,N_13143);
or U13385 (N_13385,N_13142,N_13158);
nand U13386 (N_13386,N_12974,N_12945);
nor U13387 (N_13387,N_13004,N_12971);
or U13388 (N_13388,N_12960,N_13132);
or U13389 (N_13389,N_13111,N_13072);
and U13390 (N_13390,N_13178,N_13024);
and U13391 (N_13391,N_13169,N_13013);
xor U13392 (N_13392,N_12977,N_12948);
and U13393 (N_13393,N_12983,N_12950);
xnor U13394 (N_13394,N_13052,N_13108);
xor U13395 (N_13395,N_13001,N_13137);
nor U13396 (N_13396,N_13152,N_13049);
and U13397 (N_13397,N_13077,N_13067);
xnor U13398 (N_13398,N_12967,N_12951);
nor U13399 (N_13399,N_12961,N_13024);
and U13400 (N_13400,N_12957,N_13106);
or U13401 (N_13401,N_12983,N_12912);
nor U13402 (N_13402,N_12908,N_12914);
or U13403 (N_13403,N_13191,N_13101);
or U13404 (N_13404,N_13108,N_13011);
nand U13405 (N_13405,N_13185,N_13044);
and U13406 (N_13406,N_13068,N_12995);
or U13407 (N_13407,N_13005,N_12965);
xor U13408 (N_13408,N_12955,N_13002);
xor U13409 (N_13409,N_12947,N_13059);
nor U13410 (N_13410,N_13174,N_12990);
and U13411 (N_13411,N_12996,N_13057);
nor U13412 (N_13412,N_13118,N_13003);
and U13413 (N_13413,N_13053,N_13014);
and U13414 (N_13414,N_13157,N_13094);
or U13415 (N_13415,N_13040,N_12989);
nand U13416 (N_13416,N_12991,N_12951);
nand U13417 (N_13417,N_12983,N_13148);
nor U13418 (N_13418,N_12993,N_12901);
and U13419 (N_13419,N_13132,N_13052);
xor U13420 (N_13420,N_13186,N_12980);
xor U13421 (N_13421,N_12951,N_13030);
or U13422 (N_13422,N_13193,N_13132);
nand U13423 (N_13423,N_13196,N_13022);
or U13424 (N_13424,N_12951,N_13071);
and U13425 (N_13425,N_13110,N_13050);
xor U13426 (N_13426,N_12974,N_13002);
xnor U13427 (N_13427,N_13189,N_13133);
and U13428 (N_13428,N_13081,N_13159);
or U13429 (N_13429,N_13122,N_12963);
or U13430 (N_13430,N_12926,N_13015);
or U13431 (N_13431,N_13156,N_13093);
nand U13432 (N_13432,N_12947,N_12932);
nor U13433 (N_13433,N_12924,N_13071);
or U13434 (N_13434,N_13071,N_12988);
xnor U13435 (N_13435,N_12947,N_13104);
and U13436 (N_13436,N_13125,N_13013);
or U13437 (N_13437,N_13002,N_13015);
or U13438 (N_13438,N_13073,N_13187);
nor U13439 (N_13439,N_13103,N_13013);
or U13440 (N_13440,N_12961,N_13148);
or U13441 (N_13441,N_12976,N_13013);
nor U13442 (N_13442,N_12999,N_13073);
and U13443 (N_13443,N_13127,N_13159);
nor U13444 (N_13444,N_13106,N_13091);
and U13445 (N_13445,N_13039,N_13007);
nor U13446 (N_13446,N_13015,N_13165);
nor U13447 (N_13447,N_12928,N_13106);
or U13448 (N_13448,N_12938,N_13023);
xor U13449 (N_13449,N_13160,N_13045);
or U13450 (N_13450,N_13028,N_12988);
nand U13451 (N_13451,N_13003,N_13004);
and U13452 (N_13452,N_12985,N_13008);
and U13453 (N_13453,N_13176,N_13192);
nor U13454 (N_13454,N_12954,N_13148);
or U13455 (N_13455,N_12963,N_13062);
and U13456 (N_13456,N_13050,N_13152);
or U13457 (N_13457,N_13010,N_13036);
and U13458 (N_13458,N_13029,N_13091);
nor U13459 (N_13459,N_12964,N_12918);
xor U13460 (N_13460,N_12993,N_13198);
and U13461 (N_13461,N_13119,N_12986);
xor U13462 (N_13462,N_12971,N_12915);
xnor U13463 (N_13463,N_13159,N_12940);
or U13464 (N_13464,N_13080,N_13163);
nand U13465 (N_13465,N_13095,N_12982);
xor U13466 (N_13466,N_12900,N_13041);
nand U13467 (N_13467,N_13035,N_13034);
and U13468 (N_13468,N_13149,N_13092);
xor U13469 (N_13469,N_12965,N_13140);
nor U13470 (N_13470,N_13143,N_13164);
xnor U13471 (N_13471,N_13052,N_13063);
nand U13472 (N_13472,N_13080,N_12941);
nand U13473 (N_13473,N_13122,N_13038);
xor U13474 (N_13474,N_13004,N_13070);
nand U13475 (N_13475,N_13141,N_13180);
nand U13476 (N_13476,N_13020,N_13180);
or U13477 (N_13477,N_12965,N_13145);
xor U13478 (N_13478,N_12945,N_13177);
nand U13479 (N_13479,N_13171,N_13120);
nor U13480 (N_13480,N_13015,N_12919);
nor U13481 (N_13481,N_12965,N_12922);
nand U13482 (N_13482,N_13073,N_12907);
xnor U13483 (N_13483,N_13090,N_12901);
xnor U13484 (N_13484,N_12908,N_12938);
nor U13485 (N_13485,N_13008,N_12930);
nor U13486 (N_13486,N_13118,N_12940);
xor U13487 (N_13487,N_13131,N_13102);
nor U13488 (N_13488,N_13042,N_13069);
or U13489 (N_13489,N_13046,N_13019);
nand U13490 (N_13490,N_13152,N_13154);
nor U13491 (N_13491,N_13079,N_12962);
nand U13492 (N_13492,N_13145,N_13061);
xnor U13493 (N_13493,N_13158,N_12937);
xnor U13494 (N_13494,N_13118,N_12952);
xnor U13495 (N_13495,N_13168,N_12989);
nand U13496 (N_13496,N_13134,N_12901);
or U13497 (N_13497,N_13103,N_12912);
or U13498 (N_13498,N_12926,N_13023);
or U13499 (N_13499,N_13109,N_13073);
xor U13500 (N_13500,N_13296,N_13465);
nand U13501 (N_13501,N_13409,N_13406);
or U13502 (N_13502,N_13416,N_13272);
xnor U13503 (N_13503,N_13372,N_13303);
and U13504 (N_13504,N_13264,N_13466);
and U13505 (N_13505,N_13291,N_13282);
or U13506 (N_13506,N_13387,N_13359);
and U13507 (N_13507,N_13366,N_13382);
nand U13508 (N_13508,N_13398,N_13358);
or U13509 (N_13509,N_13364,N_13220);
nand U13510 (N_13510,N_13227,N_13297);
or U13511 (N_13511,N_13413,N_13311);
xor U13512 (N_13512,N_13336,N_13400);
or U13513 (N_13513,N_13208,N_13280);
nand U13514 (N_13514,N_13232,N_13434);
or U13515 (N_13515,N_13223,N_13460);
or U13516 (N_13516,N_13402,N_13392);
xor U13517 (N_13517,N_13329,N_13249);
nor U13518 (N_13518,N_13214,N_13486);
nor U13519 (N_13519,N_13447,N_13260);
nand U13520 (N_13520,N_13467,N_13342);
or U13521 (N_13521,N_13229,N_13320);
nand U13522 (N_13522,N_13271,N_13234);
xor U13523 (N_13523,N_13217,N_13201);
nor U13524 (N_13524,N_13492,N_13339);
nand U13525 (N_13525,N_13381,N_13301);
nand U13526 (N_13526,N_13463,N_13491);
nand U13527 (N_13527,N_13474,N_13228);
xnor U13528 (N_13528,N_13482,N_13425);
nand U13529 (N_13529,N_13391,N_13457);
nand U13530 (N_13530,N_13389,N_13266);
nand U13531 (N_13531,N_13315,N_13341);
xnor U13532 (N_13532,N_13484,N_13485);
and U13533 (N_13533,N_13452,N_13489);
nand U13534 (N_13534,N_13356,N_13243);
nand U13535 (N_13535,N_13397,N_13313);
xor U13536 (N_13536,N_13377,N_13351);
xor U13537 (N_13537,N_13479,N_13395);
or U13538 (N_13538,N_13327,N_13308);
xor U13539 (N_13539,N_13470,N_13407);
xor U13540 (N_13540,N_13499,N_13498);
nor U13541 (N_13541,N_13293,N_13419);
nor U13542 (N_13542,N_13240,N_13455);
nand U13543 (N_13543,N_13362,N_13403);
or U13544 (N_13544,N_13317,N_13261);
nor U13545 (N_13545,N_13378,N_13340);
xor U13546 (N_13546,N_13429,N_13443);
xnor U13547 (N_13547,N_13284,N_13335);
xnor U13548 (N_13548,N_13442,N_13276);
xnor U13549 (N_13549,N_13314,N_13269);
nor U13550 (N_13550,N_13350,N_13411);
nor U13551 (N_13551,N_13368,N_13490);
nand U13552 (N_13552,N_13242,N_13399);
and U13553 (N_13553,N_13424,N_13253);
and U13554 (N_13554,N_13423,N_13393);
and U13555 (N_13555,N_13202,N_13417);
xnor U13556 (N_13556,N_13312,N_13277);
nand U13557 (N_13557,N_13451,N_13306);
nand U13558 (N_13558,N_13450,N_13255);
and U13559 (N_13559,N_13493,N_13204);
xor U13560 (N_13560,N_13440,N_13310);
nor U13561 (N_13561,N_13379,N_13241);
xnor U13562 (N_13562,N_13328,N_13436);
and U13563 (N_13563,N_13290,N_13412);
nand U13564 (N_13564,N_13322,N_13363);
nand U13565 (N_13565,N_13278,N_13346);
or U13566 (N_13566,N_13235,N_13371);
nand U13567 (N_13567,N_13349,N_13325);
nor U13568 (N_13568,N_13388,N_13401);
and U13569 (N_13569,N_13225,N_13219);
nand U13570 (N_13570,N_13332,N_13333);
nand U13571 (N_13571,N_13321,N_13287);
nand U13572 (N_13572,N_13275,N_13439);
xnor U13573 (N_13573,N_13238,N_13244);
nand U13574 (N_13574,N_13268,N_13343);
nor U13575 (N_13575,N_13274,N_13211);
or U13576 (N_13576,N_13469,N_13471);
nand U13577 (N_13577,N_13319,N_13352);
and U13578 (N_13578,N_13257,N_13464);
nand U13579 (N_13579,N_13222,N_13385);
and U13580 (N_13580,N_13298,N_13408);
nor U13581 (N_13581,N_13360,N_13294);
nand U13582 (N_13582,N_13203,N_13250);
nand U13583 (N_13583,N_13483,N_13421);
or U13584 (N_13584,N_13444,N_13207);
nor U13585 (N_13585,N_13273,N_13441);
nand U13586 (N_13586,N_13410,N_13295);
or U13587 (N_13587,N_13258,N_13449);
and U13588 (N_13588,N_13422,N_13361);
or U13589 (N_13589,N_13376,N_13259);
nor U13590 (N_13590,N_13231,N_13236);
and U13591 (N_13591,N_13344,N_13237);
or U13592 (N_13592,N_13367,N_13330);
xor U13593 (N_13593,N_13307,N_13200);
nor U13594 (N_13594,N_13221,N_13256);
and U13595 (N_13595,N_13283,N_13326);
nand U13596 (N_13596,N_13438,N_13292);
and U13597 (N_13597,N_13472,N_13209);
nand U13598 (N_13598,N_13248,N_13286);
xor U13599 (N_13599,N_13337,N_13239);
nor U13600 (N_13600,N_13458,N_13288);
or U13601 (N_13601,N_13216,N_13380);
and U13602 (N_13602,N_13354,N_13475);
or U13603 (N_13603,N_13233,N_13430);
and U13604 (N_13604,N_13299,N_13494);
nand U13605 (N_13605,N_13246,N_13418);
or U13606 (N_13606,N_13390,N_13496);
or U13607 (N_13607,N_13215,N_13396);
or U13608 (N_13608,N_13427,N_13426);
and U13609 (N_13609,N_13446,N_13263);
nor U13610 (N_13610,N_13477,N_13357);
nor U13611 (N_13611,N_13267,N_13394);
xor U13612 (N_13612,N_13384,N_13247);
or U13613 (N_13613,N_13369,N_13495);
nor U13614 (N_13614,N_13448,N_13254);
xnor U13615 (N_13615,N_13270,N_13281);
xor U13616 (N_13616,N_13213,N_13468);
xnor U13617 (N_13617,N_13245,N_13375);
and U13618 (N_13618,N_13265,N_13334);
xnor U13619 (N_13619,N_13252,N_13461);
nor U13620 (N_13620,N_13355,N_13453);
or U13621 (N_13621,N_13476,N_13353);
nand U13622 (N_13622,N_13230,N_13210);
or U13623 (N_13623,N_13437,N_13414);
xnor U13624 (N_13624,N_13383,N_13365);
or U13625 (N_13625,N_13279,N_13487);
nand U13626 (N_13626,N_13445,N_13224);
xnor U13627 (N_13627,N_13323,N_13212);
nand U13628 (N_13628,N_13318,N_13488);
xor U13629 (N_13629,N_13462,N_13420);
or U13630 (N_13630,N_13473,N_13302);
nor U13631 (N_13631,N_13497,N_13348);
nor U13632 (N_13632,N_13316,N_13226);
or U13633 (N_13633,N_13262,N_13218);
xor U13634 (N_13634,N_13480,N_13370);
or U13635 (N_13635,N_13324,N_13338);
and U13636 (N_13636,N_13374,N_13456);
or U13637 (N_13637,N_13206,N_13481);
or U13638 (N_13638,N_13205,N_13300);
and U13639 (N_13639,N_13331,N_13304);
nor U13640 (N_13640,N_13251,N_13435);
xnor U13641 (N_13641,N_13347,N_13405);
xor U13642 (N_13642,N_13404,N_13478);
nand U13643 (N_13643,N_13454,N_13345);
xnor U13644 (N_13644,N_13428,N_13373);
nor U13645 (N_13645,N_13386,N_13433);
or U13646 (N_13646,N_13431,N_13309);
xnor U13647 (N_13647,N_13285,N_13415);
xnor U13648 (N_13648,N_13432,N_13289);
and U13649 (N_13649,N_13305,N_13459);
nand U13650 (N_13650,N_13268,N_13244);
nand U13651 (N_13651,N_13345,N_13349);
nand U13652 (N_13652,N_13457,N_13282);
or U13653 (N_13653,N_13436,N_13319);
xnor U13654 (N_13654,N_13449,N_13220);
nor U13655 (N_13655,N_13484,N_13284);
or U13656 (N_13656,N_13255,N_13281);
or U13657 (N_13657,N_13469,N_13381);
xnor U13658 (N_13658,N_13391,N_13468);
and U13659 (N_13659,N_13253,N_13314);
or U13660 (N_13660,N_13317,N_13418);
nor U13661 (N_13661,N_13405,N_13304);
xor U13662 (N_13662,N_13476,N_13438);
nor U13663 (N_13663,N_13229,N_13474);
xnor U13664 (N_13664,N_13253,N_13298);
and U13665 (N_13665,N_13449,N_13447);
xnor U13666 (N_13666,N_13391,N_13285);
nor U13667 (N_13667,N_13492,N_13421);
or U13668 (N_13668,N_13302,N_13462);
xor U13669 (N_13669,N_13256,N_13330);
nor U13670 (N_13670,N_13351,N_13210);
nand U13671 (N_13671,N_13227,N_13238);
xor U13672 (N_13672,N_13297,N_13375);
nand U13673 (N_13673,N_13211,N_13470);
xnor U13674 (N_13674,N_13286,N_13457);
and U13675 (N_13675,N_13244,N_13463);
and U13676 (N_13676,N_13457,N_13447);
nand U13677 (N_13677,N_13210,N_13200);
and U13678 (N_13678,N_13362,N_13258);
and U13679 (N_13679,N_13285,N_13315);
nor U13680 (N_13680,N_13440,N_13418);
and U13681 (N_13681,N_13215,N_13302);
nand U13682 (N_13682,N_13450,N_13442);
xor U13683 (N_13683,N_13234,N_13238);
or U13684 (N_13684,N_13230,N_13357);
xor U13685 (N_13685,N_13397,N_13228);
and U13686 (N_13686,N_13375,N_13266);
and U13687 (N_13687,N_13487,N_13481);
and U13688 (N_13688,N_13325,N_13471);
and U13689 (N_13689,N_13252,N_13458);
nor U13690 (N_13690,N_13449,N_13210);
nor U13691 (N_13691,N_13379,N_13268);
nand U13692 (N_13692,N_13426,N_13482);
nand U13693 (N_13693,N_13388,N_13202);
nand U13694 (N_13694,N_13382,N_13397);
and U13695 (N_13695,N_13213,N_13300);
xnor U13696 (N_13696,N_13280,N_13268);
nand U13697 (N_13697,N_13384,N_13263);
nand U13698 (N_13698,N_13271,N_13405);
nand U13699 (N_13699,N_13233,N_13404);
xor U13700 (N_13700,N_13240,N_13200);
or U13701 (N_13701,N_13418,N_13456);
xor U13702 (N_13702,N_13413,N_13213);
and U13703 (N_13703,N_13287,N_13391);
nand U13704 (N_13704,N_13318,N_13249);
and U13705 (N_13705,N_13301,N_13413);
nor U13706 (N_13706,N_13308,N_13357);
or U13707 (N_13707,N_13339,N_13366);
nor U13708 (N_13708,N_13317,N_13379);
xnor U13709 (N_13709,N_13202,N_13376);
and U13710 (N_13710,N_13248,N_13461);
xor U13711 (N_13711,N_13467,N_13358);
xnor U13712 (N_13712,N_13488,N_13423);
nor U13713 (N_13713,N_13373,N_13238);
xnor U13714 (N_13714,N_13240,N_13335);
nor U13715 (N_13715,N_13473,N_13312);
nand U13716 (N_13716,N_13283,N_13363);
or U13717 (N_13717,N_13215,N_13311);
nand U13718 (N_13718,N_13412,N_13207);
xor U13719 (N_13719,N_13488,N_13305);
nor U13720 (N_13720,N_13414,N_13296);
nand U13721 (N_13721,N_13484,N_13226);
or U13722 (N_13722,N_13266,N_13221);
xor U13723 (N_13723,N_13373,N_13426);
nand U13724 (N_13724,N_13413,N_13225);
nand U13725 (N_13725,N_13304,N_13217);
nor U13726 (N_13726,N_13271,N_13291);
or U13727 (N_13727,N_13236,N_13440);
nor U13728 (N_13728,N_13485,N_13306);
and U13729 (N_13729,N_13365,N_13309);
nor U13730 (N_13730,N_13399,N_13465);
nor U13731 (N_13731,N_13297,N_13270);
xnor U13732 (N_13732,N_13401,N_13394);
nand U13733 (N_13733,N_13425,N_13330);
nand U13734 (N_13734,N_13317,N_13280);
xnor U13735 (N_13735,N_13391,N_13482);
or U13736 (N_13736,N_13449,N_13313);
and U13737 (N_13737,N_13468,N_13220);
nand U13738 (N_13738,N_13395,N_13262);
nand U13739 (N_13739,N_13359,N_13301);
nor U13740 (N_13740,N_13494,N_13202);
nor U13741 (N_13741,N_13397,N_13487);
and U13742 (N_13742,N_13362,N_13324);
nand U13743 (N_13743,N_13295,N_13204);
nand U13744 (N_13744,N_13372,N_13241);
nand U13745 (N_13745,N_13291,N_13210);
nand U13746 (N_13746,N_13339,N_13252);
xor U13747 (N_13747,N_13289,N_13459);
nor U13748 (N_13748,N_13359,N_13416);
and U13749 (N_13749,N_13230,N_13331);
nor U13750 (N_13750,N_13334,N_13346);
xor U13751 (N_13751,N_13428,N_13361);
nand U13752 (N_13752,N_13300,N_13466);
and U13753 (N_13753,N_13344,N_13387);
nand U13754 (N_13754,N_13260,N_13388);
nand U13755 (N_13755,N_13271,N_13269);
or U13756 (N_13756,N_13464,N_13485);
nor U13757 (N_13757,N_13422,N_13433);
nor U13758 (N_13758,N_13331,N_13226);
and U13759 (N_13759,N_13444,N_13351);
or U13760 (N_13760,N_13205,N_13375);
or U13761 (N_13761,N_13432,N_13321);
or U13762 (N_13762,N_13460,N_13444);
nor U13763 (N_13763,N_13383,N_13319);
and U13764 (N_13764,N_13317,N_13202);
nand U13765 (N_13765,N_13361,N_13267);
nand U13766 (N_13766,N_13361,N_13247);
or U13767 (N_13767,N_13409,N_13431);
xor U13768 (N_13768,N_13374,N_13471);
or U13769 (N_13769,N_13435,N_13422);
and U13770 (N_13770,N_13484,N_13462);
xnor U13771 (N_13771,N_13457,N_13222);
nor U13772 (N_13772,N_13235,N_13454);
nor U13773 (N_13773,N_13377,N_13463);
nor U13774 (N_13774,N_13258,N_13271);
nand U13775 (N_13775,N_13282,N_13218);
nand U13776 (N_13776,N_13217,N_13470);
nor U13777 (N_13777,N_13445,N_13286);
xor U13778 (N_13778,N_13385,N_13459);
nand U13779 (N_13779,N_13441,N_13462);
nand U13780 (N_13780,N_13288,N_13462);
xor U13781 (N_13781,N_13368,N_13264);
nor U13782 (N_13782,N_13473,N_13332);
and U13783 (N_13783,N_13410,N_13489);
nand U13784 (N_13784,N_13400,N_13232);
nand U13785 (N_13785,N_13215,N_13418);
and U13786 (N_13786,N_13365,N_13205);
nor U13787 (N_13787,N_13497,N_13317);
and U13788 (N_13788,N_13234,N_13339);
xor U13789 (N_13789,N_13342,N_13473);
or U13790 (N_13790,N_13364,N_13267);
xor U13791 (N_13791,N_13243,N_13292);
xnor U13792 (N_13792,N_13316,N_13351);
or U13793 (N_13793,N_13469,N_13379);
nand U13794 (N_13794,N_13463,N_13324);
or U13795 (N_13795,N_13246,N_13460);
or U13796 (N_13796,N_13276,N_13367);
xor U13797 (N_13797,N_13376,N_13499);
and U13798 (N_13798,N_13225,N_13468);
nand U13799 (N_13799,N_13280,N_13241);
nand U13800 (N_13800,N_13655,N_13561);
xor U13801 (N_13801,N_13538,N_13694);
and U13802 (N_13802,N_13589,N_13748);
nor U13803 (N_13803,N_13560,N_13578);
nand U13804 (N_13804,N_13516,N_13558);
or U13805 (N_13805,N_13547,N_13763);
or U13806 (N_13806,N_13778,N_13752);
xor U13807 (N_13807,N_13537,N_13684);
nand U13808 (N_13808,N_13587,N_13786);
or U13809 (N_13809,N_13795,N_13730);
nand U13810 (N_13810,N_13588,N_13500);
or U13811 (N_13811,N_13712,N_13606);
xnor U13812 (N_13812,N_13534,N_13768);
nand U13813 (N_13813,N_13650,N_13724);
nand U13814 (N_13814,N_13671,N_13703);
and U13815 (N_13815,N_13636,N_13743);
or U13816 (N_13816,N_13581,N_13766);
or U13817 (N_13817,N_13510,N_13754);
and U13818 (N_13818,N_13612,N_13523);
or U13819 (N_13819,N_13770,N_13539);
or U13820 (N_13820,N_13758,N_13676);
nand U13821 (N_13821,N_13624,N_13511);
nor U13822 (N_13822,N_13557,N_13501);
or U13823 (N_13823,N_13717,N_13701);
nor U13824 (N_13824,N_13663,N_13540);
and U13825 (N_13825,N_13673,N_13771);
nand U13826 (N_13826,N_13633,N_13692);
nand U13827 (N_13827,N_13575,N_13610);
nand U13828 (N_13828,N_13562,N_13652);
and U13829 (N_13829,N_13546,N_13729);
nor U13830 (N_13830,N_13735,N_13648);
or U13831 (N_13831,N_13765,N_13661);
and U13832 (N_13832,N_13611,N_13638);
and U13833 (N_13833,N_13660,N_13642);
nand U13834 (N_13834,N_13598,N_13625);
or U13835 (N_13835,N_13622,N_13618);
xor U13836 (N_13836,N_13640,N_13721);
xor U13837 (N_13837,N_13720,N_13797);
or U13838 (N_13838,N_13619,N_13744);
xor U13839 (N_13839,N_13616,N_13774);
xor U13840 (N_13840,N_13653,N_13704);
or U13841 (N_13841,N_13631,N_13769);
or U13842 (N_13842,N_13722,N_13686);
xnor U13843 (N_13843,N_13544,N_13515);
nand U13844 (N_13844,N_13741,N_13759);
or U13845 (N_13845,N_13691,N_13506);
or U13846 (N_13846,N_13723,N_13607);
nand U13847 (N_13847,N_13714,N_13702);
or U13848 (N_13848,N_13545,N_13525);
nor U13849 (N_13849,N_13597,N_13678);
or U13850 (N_13850,N_13502,N_13629);
and U13851 (N_13851,N_13617,N_13666);
or U13852 (N_13852,N_13750,N_13570);
nor U13853 (N_13853,N_13621,N_13669);
nand U13854 (N_13854,N_13541,N_13643);
xor U13855 (N_13855,N_13708,N_13637);
xnor U13856 (N_13856,N_13667,N_13608);
nor U13857 (N_13857,N_13605,N_13734);
or U13858 (N_13858,N_13591,N_13577);
and U13859 (N_13859,N_13664,N_13792);
or U13860 (N_13860,N_13665,N_13559);
xnor U13861 (N_13861,N_13739,N_13555);
xor U13862 (N_13862,N_13767,N_13609);
nand U13863 (N_13863,N_13527,N_13590);
or U13864 (N_13864,N_13674,N_13695);
and U13865 (N_13865,N_13747,N_13614);
xnor U13866 (N_13866,N_13505,N_13715);
xor U13867 (N_13867,N_13646,N_13514);
nand U13868 (N_13868,N_13751,N_13794);
nor U13869 (N_13869,N_13574,N_13680);
and U13870 (N_13870,N_13566,N_13572);
nor U13871 (N_13871,N_13519,N_13716);
or U13872 (N_13872,N_13738,N_13543);
nand U13873 (N_13873,N_13718,N_13594);
nand U13874 (N_13874,N_13761,N_13745);
or U13875 (N_13875,N_13571,N_13756);
nor U13876 (N_13876,N_13528,N_13706);
nor U13877 (N_13877,N_13634,N_13728);
xnor U13878 (N_13878,N_13707,N_13705);
xnor U13879 (N_13879,N_13777,N_13697);
xor U13880 (N_13880,N_13567,N_13710);
xor U13881 (N_13881,N_13579,N_13632);
and U13882 (N_13882,N_13799,N_13656);
nor U13883 (N_13883,N_13682,N_13757);
xor U13884 (N_13884,N_13796,N_13635);
nor U13885 (N_13885,N_13583,N_13709);
nand U13886 (N_13886,N_13564,N_13530);
and U13887 (N_13887,N_13503,N_13569);
nand U13888 (N_13888,N_13736,N_13781);
nand U13889 (N_13889,N_13762,N_13615);
xor U13890 (N_13890,N_13689,N_13536);
nand U13891 (N_13891,N_13764,N_13776);
and U13892 (N_13892,N_13737,N_13772);
and U13893 (N_13893,N_13782,N_13732);
xor U13894 (N_13894,N_13688,N_13753);
and U13895 (N_13895,N_13602,N_13662);
nand U13896 (N_13896,N_13604,N_13654);
nor U13897 (N_13897,N_13725,N_13649);
and U13898 (N_13898,N_13627,N_13672);
nor U13899 (N_13899,N_13513,N_13585);
xor U13900 (N_13900,N_13563,N_13573);
and U13901 (N_13901,N_13698,N_13613);
or U13902 (N_13902,N_13524,N_13526);
and U13903 (N_13903,N_13601,N_13670);
nor U13904 (N_13904,N_13647,N_13532);
xor U13905 (N_13905,N_13584,N_13517);
and U13906 (N_13906,N_13711,N_13639);
xor U13907 (N_13907,N_13580,N_13785);
nor U13908 (N_13908,N_13760,N_13749);
xnor U13909 (N_13909,N_13586,N_13508);
and U13910 (N_13910,N_13790,N_13623);
and U13911 (N_13911,N_13630,N_13641);
or U13912 (N_13912,N_13690,N_13521);
xor U13913 (N_13913,N_13775,N_13683);
and U13914 (N_13914,N_13783,N_13522);
and U13915 (N_13915,N_13582,N_13626);
or U13916 (N_13916,N_13719,N_13620);
nand U13917 (N_13917,N_13507,N_13677);
nor U13918 (N_13918,N_13727,N_13657);
nor U13919 (N_13919,N_13509,N_13791);
nor U13920 (N_13920,N_13518,N_13568);
nand U13921 (N_13921,N_13595,N_13787);
xor U13922 (N_13922,N_13600,N_13713);
nand U13923 (N_13923,N_13779,N_13645);
xor U13924 (N_13924,N_13789,N_13599);
and U13925 (N_13925,N_13529,N_13512);
or U13926 (N_13926,N_13780,N_13554);
and U13927 (N_13927,N_13726,N_13504);
xor U13928 (N_13928,N_13651,N_13733);
nor U13929 (N_13929,N_13731,N_13693);
or U13930 (N_13930,N_13548,N_13593);
nand U13931 (N_13931,N_13784,N_13742);
nor U13932 (N_13932,N_13793,N_13556);
nand U13933 (N_13933,N_13531,N_13746);
xor U13934 (N_13934,N_13542,N_13668);
nand U13935 (N_13935,N_13679,N_13681);
and U13936 (N_13936,N_13687,N_13565);
nor U13937 (N_13937,N_13788,N_13535);
or U13938 (N_13938,N_13685,N_13550);
and U13939 (N_13939,N_13700,N_13551);
nand U13940 (N_13940,N_13773,N_13596);
nand U13941 (N_13941,N_13603,N_13576);
and U13942 (N_13942,N_13552,N_13755);
nand U13943 (N_13943,N_13628,N_13658);
and U13944 (N_13944,N_13699,N_13644);
nand U13945 (N_13945,N_13740,N_13696);
nand U13946 (N_13946,N_13659,N_13549);
nor U13947 (N_13947,N_13520,N_13798);
xor U13948 (N_13948,N_13675,N_13592);
nand U13949 (N_13949,N_13553,N_13533);
nor U13950 (N_13950,N_13728,N_13525);
and U13951 (N_13951,N_13799,N_13695);
nand U13952 (N_13952,N_13544,N_13599);
and U13953 (N_13953,N_13621,N_13629);
xor U13954 (N_13954,N_13652,N_13601);
nor U13955 (N_13955,N_13564,N_13528);
or U13956 (N_13956,N_13666,N_13651);
nand U13957 (N_13957,N_13579,N_13669);
and U13958 (N_13958,N_13744,N_13623);
and U13959 (N_13959,N_13623,N_13562);
xnor U13960 (N_13960,N_13570,N_13794);
and U13961 (N_13961,N_13607,N_13660);
nor U13962 (N_13962,N_13768,N_13679);
nand U13963 (N_13963,N_13548,N_13539);
nor U13964 (N_13964,N_13603,N_13584);
nor U13965 (N_13965,N_13673,N_13621);
xnor U13966 (N_13966,N_13714,N_13741);
nand U13967 (N_13967,N_13565,N_13691);
xnor U13968 (N_13968,N_13613,N_13562);
nor U13969 (N_13969,N_13531,N_13748);
nor U13970 (N_13970,N_13611,N_13626);
nand U13971 (N_13971,N_13712,N_13647);
or U13972 (N_13972,N_13504,N_13655);
nand U13973 (N_13973,N_13520,N_13690);
nand U13974 (N_13974,N_13767,N_13769);
and U13975 (N_13975,N_13687,N_13667);
or U13976 (N_13976,N_13754,N_13607);
or U13977 (N_13977,N_13583,N_13724);
and U13978 (N_13978,N_13614,N_13787);
nand U13979 (N_13979,N_13691,N_13713);
xnor U13980 (N_13980,N_13766,N_13700);
and U13981 (N_13981,N_13665,N_13542);
and U13982 (N_13982,N_13769,N_13575);
xor U13983 (N_13983,N_13625,N_13767);
or U13984 (N_13984,N_13631,N_13603);
and U13985 (N_13985,N_13641,N_13532);
xnor U13986 (N_13986,N_13680,N_13522);
and U13987 (N_13987,N_13693,N_13567);
and U13988 (N_13988,N_13710,N_13636);
or U13989 (N_13989,N_13523,N_13515);
nand U13990 (N_13990,N_13757,N_13798);
nand U13991 (N_13991,N_13598,N_13540);
nor U13992 (N_13992,N_13655,N_13625);
or U13993 (N_13993,N_13676,N_13725);
or U13994 (N_13994,N_13627,N_13655);
or U13995 (N_13995,N_13649,N_13595);
nand U13996 (N_13996,N_13687,N_13535);
xnor U13997 (N_13997,N_13707,N_13504);
nand U13998 (N_13998,N_13753,N_13777);
nand U13999 (N_13999,N_13558,N_13721);
xnor U14000 (N_14000,N_13796,N_13702);
or U14001 (N_14001,N_13697,N_13546);
xnor U14002 (N_14002,N_13651,N_13569);
nand U14003 (N_14003,N_13693,N_13598);
and U14004 (N_14004,N_13616,N_13729);
and U14005 (N_14005,N_13780,N_13722);
and U14006 (N_14006,N_13743,N_13666);
and U14007 (N_14007,N_13636,N_13701);
nor U14008 (N_14008,N_13666,N_13662);
nor U14009 (N_14009,N_13701,N_13542);
and U14010 (N_14010,N_13723,N_13706);
and U14011 (N_14011,N_13776,N_13571);
nand U14012 (N_14012,N_13619,N_13787);
or U14013 (N_14013,N_13533,N_13785);
or U14014 (N_14014,N_13564,N_13793);
xor U14015 (N_14015,N_13514,N_13766);
nand U14016 (N_14016,N_13658,N_13587);
xnor U14017 (N_14017,N_13705,N_13562);
xnor U14018 (N_14018,N_13783,N_13563);
nor U14019 (N_14019,N_13720,N_13609);
or U14020 (N_14020,N_13712,N_13572);
xor U14021 (N_14021,N_13558,N_13663);
and U14022 (N_14022,N_13679,N_13719);
nand U14023 (N_14023,N_13600,N_13749);
and U14024 (N_14024,N_13755,N_13640);
nand U14025 (N_14025,N_13657,N_13768);
and U14026 (N_14026,N_13781,N_13741);
or U14027 (N_14027,N_13705,N_13554);
nand U14028 (N_14028,N_13748,N_13516);
and U14029 (N_14029,N_13739,N_13594);
nand U14030 (N_14030,N_13542,N_13601);
nand U14031 (N_14031,N_13769,N_13514);
nor U14032 (N_14032,N_13628,N_13635);
or U14033 (N_14033,N_13641,N_13751);
nand U14034 (N_14034,N_13569,N_13693);
nand U14035 (N_14035,N_13542,N_13719);
nor U14036 (N_14036,N_13524,N_13585);
nor U14037 (N_14037,N_13750,N_13653);
nand U14038 (N_14038,N_13631,N_13741);
xnor U14039 (N_14039,N_13633,N_13653);
nor U14040 (N_14040,N_13614,N_13558);
nand U14041 (N_14041,N_13723,N_13585);
xor U14042 (N_14042,N_13794,N_13612);
nor U14043 (N_14043,N_13664,N_13696);
or U14044 (N_14044,N_13630,N_13505);
or U14045 (N_14045,N_13651,N_13661);
and U14046 (N_14046,N_13513,N_13598);
and U14047 (N_14047,N_13657,N_13702);
xnor U14048 (N_14048,N_13781,N_13547);
nand U14049 (N_14049,N_13690,N_13604);
xnor U14050 (N_14050,N_13688,N_13668);
and U14051 (N_14051,N_13764,N_13788);
and U14052 (N_14052,N_13538,N_13570);
or U14053 (N_14053,N_13618,N_13552);
or U14054 (N_14054,N_13680,N_13780);
or U14055 (N_14055,N_13718,N_13510);
nand U14056 (N_14056,N_13682,N_13693);
nand U14057 (N_14057,N_13722,N_13533);
or U14058 (N_14058,N_13653,N_13536);
xor U14059 (N_14059,N_13595,N_13538);
xor U14060 (N_14060,N_13625,N_13523);
and U14061 (N_14061,N_13530,N_13720);
and U14062 (N_14062,N_13570,N_13636);
nand U14063 (N_14063,N_13538,N_13795);
or U14064 (N_14064,N_13719,N_13640);
or U14065 (N_14065,N_13547,N_13659);
nor U14066 (N_14066,N_13584,N_13688);
nor U14067 (N_14067,N_13579,N_13591);
nand U14068 (N_14068,N_13523,N_13560);
nor U14069 (N_14069,N_13720,N_13648);
nand U14070 (N_14070,N_13720,N_13675);
nor U14071 (N_14071,N_13700,N_13651);
or U14072 (N_14072,N_13648,N_13667);
nand U14073 (N_14073,N_13514,N_13792);
nand U14074 (N_14074,N_13757,N_13668);
nand U14075 (N_14075,N_13541,N_13748);
or U14076 (N_14076,N_13631,N_13734);
or U14077 (N_14077,N_13666,N_13785);
nand U14078 (N_14078,N_13683,N_13579);
nand U14079 (N_14079,N_13575,N_13624);
nor U14080 (N_14080,N_13563,N_13636);
nor U14081 (N_14081,N_13787,N_13649);
or U14082 (N_14082,N_13662,N_13581);
nand U14083 (N_14083,N_13718,N_13780);
or U14084 (N_14084,N_13717,N_13770);
and U14085 (N_14085,N_13735,N_13746);
xor U14086 (N_14086,N_13510,N_13559);
and U14087 (N_14087,N_13731,N_13560);
and U14088 (N_14088,N_13644,N_13629);
nand U14089 (N_14089,N_13502,N_13518);
and U14090 (N_14090,N_13542,N_13505);
xnor U14091 (N_14091,N_13732,N_13555);
or U14092 (N_14092,N_13658,N_13674);
nand U14093 (N_14093,N_13505,N_13585);
or U14094 (N_14094,N_13759,N_13782);
nand U14095 (N_14095,N_13524,N_13606);
or U14096 (N_14096,N_13677,N_13792);
xnor U14097 (N_14097,N_13659,N_13749);
or U14098 (N_14098,N_13664,N_13629);
xor U14099 (N_14099,N_13615,N_13797);
nor U14100 (N_14100,N_13818,N_13834);
or U14101 (N_14101,N_13901,N_13972);
nand U14102 (N_14102,N_13918,N_13993);
or U14103 (N_14103,N_14089,N_13952);
and U14104 (N_14104,N_13998,N_14044);
or U14105 (N_14105,N_14010,N_14052);
nor U14106 (N_14106,N_14032,N_13904);
and U14107 (N_14107,N_14008,N_13829);
or U14108 (N_14108,N_14023,N_13898);
nor U14109 (N_14109,N_13843,N_13945);
nor U14110 (N_14110,N_13827,N_14054);
nand U14111 (N_14111,N_13932,N_13988);
or U14112 (N_14112,N_13963,N_13833);
or U14113 (N_14113,N_13846,N_13985);
nor U14114 (N_14114,N_13810,N_13971);
or U14115 (N_14115,N_13978,N_13936);
and U14116 (N_14116,N_13990,N_13970);
xor U14117 (N_14117,N_14070,N_13864);
xnor U14118 (N_14118,N_14088,N_13938);
nor U14119 (N_14119,N_14085,N_14056);
and U14120 (N_14120,N_14005,N_13876);
or U14121 (N_14121,N_14021,N_13844);
nand U14122 (N_14122,N_14087,N_13995);
and U14123 (N_14123,N_13841,N_13839);
xor U14124 (N_14124,N_14000,N_14038);
and U14125 (N_14125,N_14036,N_13861);
and U14126 (N_14126,N_13836,N_13911);
nand U14127 (N_14127,N_13812,N_14048);
or U14128 (N_14128,N_13958,N_13851);
nor U14129 (N_14129,N_13916,N_13959);
nand U14130 (N_14130,N_14068,N_13824);
xnor U14131 (N_14131,N_13814,N_13821);
xor U14132 (N_14132,N_14096,N_13919);
or U14133 (N_14133,N_13875,N_13879);
xor U14134 (N_14134,N_13892,N_13878);
and U14135 (N_14135,N_13953,N_13873);
nand U14136 (N_14136,N_13913,N_13884);
nor U14137 (N_14137,N_13940,N_13874);
xnor U14138 (N_14138,N_13908,N_13928);
xor U14139 (N_14139,N_13862,N_13950);
nand U14140 (N_14140,N_14003,N_14067);
or U14141 (N_14141,N_13969,N_14018);
xor U14142 (N_14142,N_13866,N_14016);
xor U14143 (N_14143,N_13830,N_13820);
nand U14144 (N_14144,N_13897,N_13962);
or U14145 (N_14145,N_13907,N_13973);
xnor U14146 (N_14146,N_14046,N_14086);
or U14147 (N_14147,N_13832,N_13996);
xnor U14148 (N_14148,N_13927,N_14027);
nor U14149 (N_14149,N_13934,N_13822);
and U14150 (N_14150,N_13885,N_13888);
or U14151 (N_14151,N_13980,N_14053);
and U14152 (N_14152,N_13823,N_13889);
nor U14153 (N_14153,N_14039,N_13886);
and U14154 (N_14154,N_14082,N_14051);
nor U14155 (N_14155,N_13867,N_13806);
xor U14156 (N_14156,N_13912,N_13997);
and U14157 (N_14157,N_13893,N_14094);
nand U14158 (N_14158,N_13850,N_13986);
nor U14159 (N_14159,N_14061,N_13840);
nand U14160 (N_14160,N_13966,N_13808);
nand U14161 (N_14161,N_13807,N_14079);
or U14162 (N_14162,N_13903,N_13948);
and U14163 (N_14163,N_13954,N_13992);
nand U14164 (N_14164,N_14097,N_13925);
xor U14165 (N_14165,N_13856,N_14066);
or U14166 (N_14166,N_13848,N_13802);
nor U14167 (N_14167,N_13955,N_13964);
nor U14168 (N_14168,N_14047,N_13880);
nand U14169 (N_14169,N_14099,N_13917);
and U14170 (N_14170,N_14095,N_13989);
or U14171 (N_14171,N_14081,N_13883);
or U14172 (N_14172,N_14040,N_13894);
nand U14173 (N_14173,N_13881,N_13984);
nor U14174 (N_14174,N_14071,N_13852);
and U14175 (N_14175,N_13842,N_13943);
and U14176 (N_14176,N_13965,N_13860);
nor U14177 (N_14177,N_14043,N_13976);
nand U14178 (N_14178,N_13803,N_13982);
or U14179 (N_14179,N_14031,N_14057);
or U14180 (N_14180,N_13923,N_13921);
or U14181 (N_14181,N_14029,N_13933);
nand U14182 (N_14182,N_13999,N_13809);
or U14183 (N_14183,N_13828,N_14030);
xnor U14184 (N_14184,N_13960,N_14041);
nor U14185 (N_14185,N_14074,N_13899);
or U14186 (N_14186,N_13882,N_13871);
or U14187 (N_14187,N_13855,N_14078);
nor U14188 (N_14188,N_14092,N_13974);
xnor U14189 (N_14189,N_14072,N_14022);
and U14190 (N_14190,N_13804,N_13957);
nor U14191 (N_14191,N_13922,N_14014);
and U14192 (N_14192,N_13831,N_14049);
nand U14193 (N_14193,N_13951,N_13854);
nand U14194 (N_14194,N_14028,N_13914);
and U14195 (N_14195,N_14059,N_14050);
xnor U14196 (N_14196,N_14062,N_14025);
nor U14197 (N_14197,N_14055,N_13944);
nand U14198 (N_14198,N_14090,N_13956);
and U14199 (N_14199,N_13935,N_14083);
and U14200 (N_14200,N_13967,N_13910);
nor U14201 (N_14201,N_13939,N_13915);
xnor U14202 (N_14202,N_13946,N_14093);
nand U14203 (N_14203,N_13929,N_14013);
or U14204 (N_14204,N_14017,N_13896);
nand U14205 (N_14205,N_13994,N_13931);
nor U14206 (N_14206,N_14033,N_13975);
nor U14207 (N_14207,N_13863,N_13890);
and U14208 (N_14208,N_13909,N_13847);
xnor U14209 (N_14209,N_13845,N_14058);
or U14210 (N_14210,N_13817,N_13869);
and U14211 (N_14211,N_13977,N_14075);
and U14212 (N_14212,N_14073,N_14015);
xor U14213 (N_14213,N_13865,N_13811);
nor U14214 (N_14214,N_13905,N_13941);
xnor U14215 (N_14215,N_13983,N_13981);
nand U14216 (N_14216,N_14019,N_13877);
or U14217 (N_14217,N_14064,N_13801);
nor U14218 (N_14218,N_13900,N_13968);
xnor U14219 (N_14219,N_13895,N_13924);
xor U14220 (N_14220,N_14026,N_14076);
nand U14221 (N_14221,N_13835,N_13849);
or U14222 (N_14222,N_13815,N_13870);
xnor U14223 (N_14223,N_13805,N_13937);
xor U14224 (N_14224,N_14060,N_14077);
and U14225 (N_14225,N_14065,N_14004);
xnor U14226 (N_14226,N_14009,N_14012);
and U14227 (N_14227,N_13891,N_13868);
nand U14228 (N_14228,N_13819,N_13902);
xor U14229 (N_14229,N_13991,N_14024);
nor U14230 (N_14230,N_13930,N_14063);
and U14231 (N_14231,N_14002,N_13853);
xor U14232 (N_14232,N_14098,N_14080);
and U14233 (N_14233,N_14035,N_13961);
nand U14234 (N_14234,N_13857,N_13947);
nand U14235 (N_14235,N_14069,N_13979);
or U14236 (N_14236,N_13825,N_13858);
or U14237 (N_14237,N_13837,N_14020);
nand U14238 (N_14238,N_13920,N_13859);
and U14239 (N_14239,N_14011,N_14042);
and U14240 (N_14240,N_13826,N_13838);
nand U14241 (N_14241,N_13872,N_14006);
nand U14242 (N_14242,N_14037,N_14007);
or U14243 (N_14243,N_13926,N_13816);
xor U14244 (N_14244,N_14091,N_13887);
nor U14245 (N_14245,N_13949,N_14034);
xnor U14246 (N_14246,N_13942,N_13813);
nand U14247 (N_14247,N_13800,N_13906);
nor U14248 (N_14248,N_14045,N_14001);
nor U14249 (N_14249,N_13987,N_14084);
nand U14250 (N_14250,N_13859,N_14054);
nor U14251 (N_14251,N_13841,N_14057);
xnor U14252 (N_14252,N_14038,N_13977);
or U14253 (N_14253,N_13955,N_13942);
nor U14254 (N_14254,N_13946,N_14023);
xor U14255 (N_14255,N_13803,N_13856);
nand U14256 (N_14256,N_13893,N_13819);
or U14257 (N_14257,N_14039,N_13815);
nor U14258 (N_14258,N_13931,N_13949);
or U14259 (N_14259,N_13822,N_14039);
nor U14260 (N_14260,N_13932,N_13953);
and U14261 (N_14261,N_13886,N_14080);
xor U14262 (N_14262,N_14035,N_13842);
nand U14263 (N_14263,N_14052,N_14004);
or U14264 (N_14264,N_14070,N_13997);
and U14265 (N_14265,N_14009,N_14007);
nand U14266 (N_14266,N_13838,N_13957);
or U14267 (N_14267,N_14016,N_14031);
or U14268 (N_14268,N_13959,N_14050);
and U14269 (N_14269,N_13967,N_13880);
nor U14270 (N_14270,N_13984,N_13902);
xor U14271 (N_14271,N_14025,N_13897);
or U14272 (N_14272,N_13893,N_14056);
or U14273 (N_14273,N_13879,N_13968);
nor U14274 (N_14274,N_13808,N_13827);
or U14275 (N_14275,N_13985,N_13940);
or U14276 (N_14276,N_14040,N_13915);
xnor U14277 (N_14277,N_13829,N_13969);
nor U14278 (N_14278,N_13832,N_14081);
nand U14279 (N_14279,N_14081,N_13914);
and U14280 (N_14280,N_14058,N_14009);
nor U14281 (N_14281,N_14068,N_13837);
nand U14282 (N_14282,N_13932,N_14014);
nor U14283 (N_14283,N_14043,N_13967);
or U14284 (N_14284,N_13809,N_14096);
xnor U14285 (N_14285,N_13999,N_13996);
or U14286 (N_14286,N_13956,N_13971);
xnor U14287 (N_14287,N_14037,N_14000);
nand U14288 (N_14288,N_14063,N_13836);
and U14289 (N_14289,N_14095,N_14021);
xnor U14290 (N_14290,N_14042,N_13932);
or U14291 (N_14291,N_13824,N_13978);
xor U14292 (N_14292,N_13997,N_14074);
and U14293 (N_14293,N_13852,N_13981);
and U14294 (N_14294,N_13819,N_13978);
nor U14295 (N_14295,N_13853,N_13829);
or U14296 (N_14296,N_13867,N_13952);
xor U14297 (N_14297,N_13979,N_13977);
nor U14298 (N_14298,N_13885,N_14056);
or U14299 (N_14299,N_14076,N_13973);
or U14300 (N_14300,N_13866,N_13964);
xor U14301 (N_14301,N_14015,N_13856);
xor U14302 (N_14302,N_14009,N_14020);
nor U14303 (N_14303,N_13912,N_14069);
xor U14304 (N_14304,N_14029,N_14071);
nand U14305 (N_14305,N_13801,N_14023);
nor U14306 (N_14306,N_14091,N_13802);
xor U14307 (N_14307,N_13968,N_13931);
xor U14308 (N_14308,N_13968,N_14018);
nor U14309 (N_14309,N_13866,N_13926);
xor U14310 (N_14310,N_13858,N_13962);
or U14311 (N_14311,N_13958,N_13944);
nand U14312 (N_14312,N_13931,N_13899);
nand U14313 (N_14313,N_13851,N_13895);
nor U14314 (N_14314,N_13847,N_14062);
or U14315 (N_14315,N_14006,N_14017);
nand U14316 (N_14316,N_13858,N_14095);
and U14317 (N_14317,N_13818,N_13837);
nand U14318 (N_14318,N_14051,N_13800);
and U14319 (N_14319,N_14022,N_14050);
nor U14320 (N_14320,N_13876,N_13989);
nand U14321 (N_14321,N_14081,N_13907);
xor U14322 (N_14322,N_13935,N_13898);
xnor U14323 (N_14323,N_13820,N_13934);
or U14324 (N_14324,N_13982,N_13977);
and U14325 (N_14325,N_13867,N_14037);
nor U14326 (N_14326,N_13808,N_14000);
nand U14327 (N_14327,N_13901,N_13815);
and U14328 (N_14328,N_13847,N_13921);
or U14329 (N_14329,N_13923,N_13962);
xor U14330 (N_14330,N_14019,N_13939);
nand U14331 (N_14331,N_13917,N_13860);
nand U14332 (N_14332,N_13938,N_14062);
nand U14333 (N_14333,N_13819,N_14029);
xnor U14334 (N_14334,N_13813,N_14021);
xor U14335 (N_14335,N_14027,N_13940);
nand U14336 (N_14336,N_13825,N_14002);
or U14337 (N_14337,N_13900,N_13989);
xnor U14338 (N_14338,N_14015,N_13942);
nor U14339 (N_14339,N_14028,N_14015);
and U14340 (N_14340,N_14051,N_13932);
nand U14341 (N_14341,N_14089,N_14034);
or U14342 (N_14342,N_13926,N_13800);
xnor U14343 (N_14343,N_13881,N_13833);
nand U14344 (N_14344,N_13876,N_13985);
or U14345 (N_14345,N_14026,N_13929);
and U14346 (N_14346,N_13883,N_13966);
or U14347 (N_14347,N_13960,N_13867);
and U14348 (N_14348,N_13912,N_13810);
and U14349 (N_14349,N_13892,N_13929);
xnor U14350 (N_14350,N_13867,N_14004);
nand U14351 (N_14351,N_13888,N_14008);
xnor U14352 (N_14352,N_14039,N_14034);
xnor U14353 (N_14353,N_13899,N_14044);
and U14354 (N_14354,N_13855,N_13877);
nor U14355 (N_14355,N_14020,N_13936);
nor U14356 (N_14356,N_13921,N_13932);
xnor U14357 (N_14357,N_14051,N_13811);
nor U14358 (N_14358,N_14043,N_13972);
xor U14359 (N_14359,N_13906,N_13905);
nor U14360 (N_14360,N_13830,N_13855);
or U14361 (N_14361,N_13834,N_13856);
and U14362 (N_14362,N_13988,N_13852);
nand U14363 (N_14363,N_13917,N_13828);
or U14364 (N_14364,N_13908,N_13874);
or U14365 (N_14365,N_13916,N_14044);
or U14366 (N_14366,N_13879,N_14018);
or U14367 (N_14367,N_13826,N_13904);
and U14368 (N_14368,N_13952,N_14003);
nor U14369 (N_14369,N_13806,N_13934);
xnor U14370 (N_14370,N_13874,N_13860);
nor U14371 (N_14371,N_13820,N_14093);
and U14372 (N_14372,N_13893,N_14031);
xnor U14373 (N_14373,N_13980,N_13861);
or U14374 (N_14374,N_13869,N_13984);
xnor U14375 (N_14375,N_13886,N_13878);
and U14376 (N_14376,N_13918,N_13826);
nand U14377 (N_14377,N_13808,N_13866);
and U14378 (N_14378,N_14080,N_14081);
nand U14379 (N_14379,N_13852,N_14084);
or U14380 (N_14380,N_14077,N_13851);
nand U14381 (N_14381,N_13838,N_13846);
nor U14382 (N_14382,N_14053,N_14093);
nor U14383 (N_14383,N_13938,N_14043);
nand U14384 (N_14384,N_14000,N_13934);
xor U14385 (N_14385,N_13936,N_13897);
and U14386 (N_14386,N_13830,N_13961);
and U14387 (N_14387,N_13906,N_13862);
nor U14388 (N_14388,N_13809,N_13860);
or U14389 (N_14389,N_13939,N_13894);
and U14390 (N_14390,N_14010,N_14018);
and U14391 (N_14391,N_13871,N_13941);
and U14392 (N_14392,N_13864,N_13950);
xnor U14393 (N_14393,N_14029,N_14030);
and U14394 (N_14394,N_14007,N_13823);
xnor U14395 (N_14395,N_13978,N_13901);
or U14396 (N_14396,N_14076,N_13855);
nand U14397 (N_14397,N_13944,N_14057);
nand U14398 (N_14398,N_14013,N_13955);
nor U14399 (N_14399,N_13878,N_13807);
nand U14400 (N_14400,N_14232,N_14160);
and U14401 (N_14401,N_14381,N_14121);
nand U14402 (N_14402,N_14233,N_14378);
or U14403 (N_14403,N_14146,N_14132);
or U14404 (N_14404,N_14138,N_14155);
xnor U14405 (N_14405,N_14323,N_14330);
xnor U14406 (N_14406,N_14311,N_14398);
nand U14407 (N_14407,N_14290,N_14310);
xor U14408 (N_14408,N_14273,N_14343);
xnor U14409 (N_14409,N_14141,N_14136);
or U14410 (N_14410,N_14271,N_14113);
and U14411 (N_14411,N_14102,N_14105);
and U14412 (N_14412,N_14336,N_14352);
nor U14413 (N_14413,N_14103,N_14151);
xor U14414 (N_14414,N_14143,N_14298);
and U14415 (N_14415,N_14209,N_14110);
nand U14416 (N_14416,N_14388,N_14373);
nand U14417 (N_14417,N_14314,N_14159);
nor U14418 (N_14418,N_14197,N_14237);
and U14419 (N_14419,N_14297,N_14302);
nor U14420 (N_14420,N_14194,N_14335);
or U14421 (N_14421,N_14384,N_14184);
xor U14422 (N_14422,N_14111,N_14235);
nor U14423 (N_14423,N_14361,N_14285);
and U14424 (N_14424,N_14345,N_14312);
xor U14425 (N_14425,N_14327,N_14210);
nor U14426 (N_14426,N_14245,N_14180);
nand U14427 (N_14427,N_14203,N_14274);
or U14428 (N_14428,N_14291,N_14251);
xnor U14429 (N_14429,N_14179,N_14288);
or U14430 (N_14430,N_14128,N_14137);
nand U14431 (N_14431,N_14346,N_14217);
nor U14432 (N_14432,N_14223,N_14258);
nand U14433 (N_14433,N_14222,N_14161);
nand U14434 (N_14434,N_14351,N_14199);
nor U14435 (N_14435,N_14394,N_14305);
nor U14436 (N_14436,N_14348,N_14249);
nand U14437 (N_14437,N_14148,N_14192);
nand U14438 (N_14438,N_14124,N_14317);
xor U14439 (N_14439,N_14172,N_14269);
xor U14440 (N_14440,N_14322,N_14218);
nand U14441 (N_14441,N_14153,N_14385);
and U14442 (N_14442,N_14278,N_14375);
nor U14443 (N_14443,N_14100,N_14119);
and U14444 (N_14444,N_14123,N_14283);
xor U14445 (N_14445,N_14115,N_14204);
or U14446 (N_14446,N_14248,N_14207);
nand U14447 (N_14447,N_14307,N_14337);
nand U14448 (N_14448,N_14157,N_14185);
and U14449 (N_14449,N_14170,N_14377);
or U14450 (N_14450,N_14272,N_14395);
and U14451 (N_14451,N_14347,N_14397);
and U14452 (N_14452,N_14193,N_14396);
nor U14453 (N_14453,N_14147,N_14133);
and U14454 (N_14454,N_14301,N_14380);
xor U14455 (N_14455,N_14164,N_14112);
xor U14456 (N_14456,N_14122,N_14333);
nand U14457 (N_14457,N_14247,N_14349);
or U14458 (N_14458,N_14230,N_14226);
nand U14459 (N_14459,N_14229,N_14366);
nor U14460 (N_14460,N_14324,N_14162);
and U14461 (N_14461,N_14332,N_14340);
xor U14462 (N_14462,N_14279,N_14399);
xor U14463 (N_14463,N_14221,N_14383);
nor U14464 (N_14464,N_14236,N_14242);
nor U14465 (N_14465,N_14254,N_14107);
and U14466 (N_14466,N_14265,N_14227);
xor U14467 (N_14467,N_14319,N_14326);
nor U14468 (N_14468,N_14144,N_14268);
nor U14469 (N_14469,N_14156,N_14244);
or U14470 (N_14470,N_14356,N_14270);
or U14471 (N_14471,N_14306,N_14320);
xnor U14472 (N_14472,N_14211,N_14339);
and U14473 (N_14473,N_14262,N_14140);
and U14474 (N_14474,N_14364,N_14292);
xnor U14475 (N_14475,N_14101,N_14154);
xnor U14476 (N_14476,N_14240,N_14300);
and U14477 (N_14477,N_14304,N_14241);
xor U14478 (N_14478,N_14321,N_14250);
xor U14479 (N_14479,N_14167,N_14176);
nand U14480 (N_14480,N_14374,N_14390);
and U14481 (N_14481,N_14116,N_14277);
xnor U14482 (N_14482,N_14369,N_14256);
or U14483 (N_14483,N_14208,N_14216);
nor U14484 (N_14484,N_14393,N_14360);
or U14485 (N_14485,N_14252,N_14253);
nand U14486 (N_14486,N_14299,N_14125);
nand U14487 (N_14487,N_14341,N_14282);
and U14488 (N_14488,N_14120,N_14201);
or U14489 (N_14489,N_14165,N_14359);
nor U14490 (N_14490,N_14135,N_14225);
nor U14491 (N_14491,N_14382,N_14246);
xor U14492 (N_14492,N_14353,N_14309);
and U14493 (N_14493,N_14266,N_14202);
or U14494 (N_14494,N_14189,N_14200);
xor U14495 (N_14495,N_14114,N_14354);
or U14496 (N_14496,N_14130,N_14166);
nor U14497 (N_14497,N_14280,N_14183);
and U14498 (N_14498,N_14386,N_14328);
or U14499 (N_14499,N_14308,N_14205);
and U14500 (N_14500,N_14220,N_14379);
nor U14501 (N_14501,N_14387,N_14342);
xor U14502 (N_14502,N_14257,N_14368);
xnor U14503 (N_14503,N_14198,N_14255);
or U14504 (N_14504,N_14303,N_14267);
or U14505 (N_14505,N_14287,N_14163);
nand U14506 (N_14506,N_14259,N_14158);
nor U14507 (N_14507,N_14372,N_14129);
nor U14508 (N_14508,N_14392,N_14171);
or U14509 (N_14509,N_14338,N_14215);
nor U14510 (N_14510,N_14108,N_14178);
and U14511 (N_14511,N_14318,N_14173);
nor U14512 (N_14512,N_14296,N_14334);
and U14513 (N_14513,N_14175,N_14182);
nand U14514 (N_14514,N_14239,N_14294);
xnor U14515 (N_14515,N_14325,N_14362);
nor U14516 (N_14516,N_14391,N_14186);
nor U14517 (N_14517,N_14231,N_14264);
nand U14518 (N_14518,N_14367,N_14219);
or U14519 (N_14519,N_14109,N_14126);
nor U14520 (N_14520,N_14181,N_14260);
xor U14521 (N_14521,N_14196,N_14224);
xnor U14522 (N_14522,N_14243,N_14263);
xor U14523 (N_14523,N_14376,N_14131);
or U14524 (N_14524,N_14295,N_14355);
nand U14525 (N_14525,N_14127,N_14261);
nor U14526 (N_14526,N_14139,N_14149);
xor U14527 (N_14527,N_14358,N_14316);
or U14528 (N_14528,N_14195,N_14191);
or U14529 (N_14529,N_14371,N_14187);
nand U14530 (N_14530,N_14365,N_14214);
xnor U14531 (N_14531,N_14281,N_14118);
nor U14532 (N_14532,N_14117,N_14106);
nand U14533 (N_14533,N_14363,N_14152);
and U14534 (N_14534,N_14228,N_14357);
xnor U14535 (N_14535,N_14344,N_14350);
xnor U14536 (N_14536,N_14313,N_14212);
nor U14537 (N_14537,N_14168,N_14331);
and U14538 (N_14538,N_14169,N_14150);
and U14539 (N_14539,N_14104,N_14275);
or U14540 (N_14540,N_14284,N_14293);
xor U14541 (N_14541,N_14206,N_14134);
nand U14542 (N_14542,N_14174,N_14370);
nor U14543 (N_14543,N_14188,N_14190);
and U14544 (N_14544,N_14213,N_14142);
xnor U14545 (N_14545,N_14238,N_14315);
nor U14546 (N_14546,N_14234,N_14329);
nor U14547 (N_14547,N_14286,N_14276);
nand U14548 (N_14548,N_14145,N_14289);
or U14549 (N_14549,N_14389,N_14177);
nand U14550 (N_14550,N_14361,N_14279);
nand U14551 (N_14551,N_14113,N_14128);
and U14552 (N_14552,N_14359,N_14147);
nand U14553 (N_14553,N_14173,N_14186);
xor U14554 (N_14554,N_14386,N_14225);
xnor U14555 (N_14555,N_14236,N_14133);
and U14556 (N_14556,N_14268,N_14353);
xnor U14557 (N_14557,N_14376,N_14240);
xnor U14558 (N_14558,N_14267,N_14308);
nor U14559 (N_14559,N_14146,N_14381);
nor U14560 (N_14560,N_14325,N_14184);
or U14561 (N_14561,N_14228,N_14379);
nand U14562 (N_14562,N_14334,N_14161);
or U14563 (N_14563,N_14250,N_14331);
xnor U14564 (N_14564,N_14106,N_14197);
nor U14565 (N_14565,N_14138,N_14229);
and U14566 (N_14566,N_14211,N_14120);
nor U14567 (N_14567,N_14323,N_14146);
xnor U14568 (N_14568,N_14115,N_14267);
or U14569 (N_14569,N_14262,N_14151);
xor U14570 (N_14570,N_14389,N_14143);
and U14571 (N_14571,N_14121,N_14183);
or U14572 (N_14572,N_14130,N_14144);
and U14573 (N_14573,N_14396,N_14300);
nor U14574 (N_14574,N_14274,N_14211);
and U14575 (N_14575,N_14289,N_14228);
nor U14576 (N_14576,N_14140,N_14355);
nor U14577 (N_14577,N_14263,N_14274);
nand U14578 (N_14578,N_14365,N_14107);
or U14579 (N_14579,N_14319,N_14100);
or U14580 (N_14580,N_14351,N_14158);
xor U14581 (N_14581,N_14383,N_14369);
nor U14582 (N_14582,N_14211,N_14121);
or U14583 (N_14583,N_14311,N_14241);
xnor U14584 (N_14584,N_14342,N_14225);
nand U14585 (N_14585,N_14314,N_14149);
nor U14586 (N_14586,N_14147,N_14343);
nand U14587 (N_14587,N_14234,N_14162);
nor U14588 (N_14588,N_14115,N_14105);
or U14589 (N_14589,N_14297,N_14151);
xnor U14590 (N_14590,N_14387,N_14213);
and U14591 (N_14591,N_14392,N_14380);
nor U14592 (N_14592,N_14274,N_14236);
nor U14593 (N_14593,N_14362,N_14104);
and U14594 (N_14594,N_14178,N_14169);
or U14595 (N_14595,N_14160,N_14133);
nor U14596 (N_14596,N_14360,N_14250);
nor U14597 (N_14597,N_14332,N_14148);
nor U14598 (N_14598,N_14198,N_14241);
nand U14599 (N_14599,N_14262,N_14193);
xor U14600 (N_14600,N_14355,N_14352);
nor U14601 (N_14601,N_14155,N_14264);
nor U14602 (N_14602,N_14274,N_14111);
xor U14603 (N_14603,N_14363,N_14389);
xor U14604 (N_14604,N_14247,N_14194);
xor U14605 (N_14605,N_14210,N_14161);
nand U14606 (N_14606,N_14390,N_14137);
and U14607 (N_14607,N_14273,N_14146);
or U14608 (N_14608,N_14222,N_14359);
nand U14609 (N_14609,N_14142,N_14334);
nor U14610 (N_14610,N_14131,N_14168);
xnor U14611 (N_14611,N_14130,N_14373);
or U14612 (N_14612,N_14143,N_14399);
nand U14613 (N_14613,N_14364,N_14357);
or U14614 (N_14614,N_14139,N_14331);
and U14615 (N_14615,N_14104,N_14246);
nor U14616 (N_14616,N_14254,N_14262);
and U14617 (N_14617,N_14318,N_14153);
nor U14618 (N_14618,N_14128,N_14114);
xor U14619 (N_14619,N_14238,N_14193);
or U14620 (N_14620,N_14341,N_14238);
or U14621 (N_14621,N_14109,N_14240);
or U14622 (N_14622,N_14138,N_14390);
or U14623 (N_14623,N_14275,N_14174);
nor U14624 (N_14624,N_14303,N_14114);
nand U14625 (N_14625,N_14181,N_14224);
or U14626 (N_14626,N_14129,N_14289);
nand U14627 (N_14627,N_14117,N_14344);
nor U14628 (N_14628,N_14196,N_14100);
xor U14629 (N_14629,N_14387,N_14334);
nand U14630 (N_14630,N_14212,N_14336);
or U14631 (N_14631,N_14347,N_14286);
or U14632 (N_14632,N_14120,N_14182);
and U14633 (N_14633,N_14230,N_14358);
nor U14634 (N_14634,N_14385,N_14292);
xor U14635 (N_14635,N_14139,N_14304);
nor U14636 (N_14636,N_14282,N_14213);
or U14637 (N_14637,N_14362,N_14259);
nand U14638 (N_14638,N_14178,N_14141);
nor U14639 (N_14639,N_14140,N_14129);
nor U14640 (N_14640,N_14323,N_14189);
or U14641 (N_14641,N_14231,N_14259);
xor U14642 (N_14642,N_14297,N_14288);
and U14643 (N_14643,N_14119,N_14317);
xor U14644 (N_14644,N_14136,N_14244);
or U14645 (N_14645,N_14337,N_14341);
nand U14646 (N_14646,N_14216,N_14127);
and U14647 (N_14647,N_14344,N_14125);
or U14648 (N_14648,N_14169,N_14319);
nand U14649 (N_14649,N_14109,N_14102);
or U14650 (N_14650,N_14397,N_14287);
xnor U14651 (N_14651,N_14148,N_14234);
nand U14652 (N_14652,N_14141,N_14308);
nand U14653 (N_14653,N_14294,N_14103);
nand U14654 (N_14654,N_14141,N_14343);
nand U14655 (N_14655,N_14331,N_14323);
nor U14656 (N_14656,N_14171,N_14265);
nor U14657 (N_14657,N_14326,N_14179);
nand U14658 (N_14658,N_14302,N_14272);
and U14659 (N_14659,N_14340,N_14375);
nand U14660 (N_14660,N_14161,N_14269);
xnor U14661 (N_14661,N_14198,N_14376);
xor U14662 (N_14662,N_14288,N_14358);
xnor U14663 (N_14663,N_14383,N_14100);
xnor U14664 (N_14664,N_14105,N_14101);
xnor U14665 (N_14665,N_14302,N_14239);
xor U14666 (N_14666,N_14357,N_14353);
nand U14667 (N_14667,N_14238,N_14240);
and U14668 (N_14668,N_14168,N_14343);
or U14669 (N_14669,N_14327,N_14270);
nor U14670 (N_14670,N_14117,N_14147);
xnor U14671 (N_14671,N_14213,N_14139);
or U14672 (N_14672,N_14319,N_14261);
nand U14673 (N_14673,N_14300,N_14110);
nor U14674 (N_14674,N_14275,N_14207);
and U14675 (N_14675,N_14121,N_14331);
or U14676 (N_14676,N_14341,N_14145);
or U14677 (N_14677,N_14254,N_14127);
nand U14678 (N_14678,N_14219,N_14188);
and U14679 (N_14679,N_14201,N_14233);
and U14680 (N_14680,N_14287,N_14124);
nand U14681 (N_14681,N_14359,N_14283);
or U14682 (N_14682,N_14138,N_14226);
nor U14683 (N_14683,N_14362,N_14183);
nand U14684 (N_14684,N_14232,N_14365);
nor U14685 (N_14685,N_14338,N_14184);
and U14686 (N_14686,N_14165,N_14373);
or U14687 (N_14687,N_14264,N_14164);
or U14688 (N_14688,N_14382,N_14369);
or U14689 (N_14689,N_14393,N_14308);
nor U14690 (N_14690,N_14165,N_14306);
and U14691 (N_14691,N_14180,N_14386);
nand U14692 (N_14692,N_14254,N_14362);
or U14693 (N_14693,N_14123,N_14175);
and U14694 (N_14694,N_14171,N_14276);
and U14695 (N_14695,N_14294,N_14358);
nand U14696 (N_14696,N_14275,N_14183);
nor U14697 (N_14697,N_14397,N_14293);
or U14698 (N_14698,N_14309,N_14119);
or U14699 (N_14699,N_14109,N_14360);
or U14700 (N_14700,N_14610,N_14426);
xor U14701 (N_14701,N_14415,N_14460);
nor U14702 (N_14702,N_14541,N_14492);
nor U14703 (N_14703,N_14548,N_14424);
and U14704 (N_14704,N_14425,N_14502);
or U14705 (N_14705,N_14442,N_14446);
and U14706 (N_14706,N_14454,N_14698);
nand U14707 (N_14707,N_14571,N_14532);
xnor U14708 (N_14708,N_14633,N_14579);
nand U14709 (N_14709,N_14540,N_14597);
or U14710 (N_14710,N_14476,N_14543);
xor U14711 (N_14711,N_14521,N_14598);
nand U14712 (N_14712,N_14483,N_14494);
and U14713 (N_14713,N_14674,N_14662);
nand U14714 (N_14714,N_14650,N_14625);
nand U14715 (N_14715,N_14689,N_14513);
xor U14716 (N_14716,N_14501,N_14453);
or U14717 (N_14717,N_14622,N_14599);
xor U14718 (N_14718,N_14652,N_14692);
and U14719 (N_14719,N_14518,N_14410);
xnor U14720 (N_14720,N_14470,N_14581);
and U14721 (N_14721,N_14432,N_14455);
xnor U14722 (N_14722,N_14627,N_14639);
nand U14723 (N_14723,N_14606,N_14507);
and U14724 (N_14724,N_14462,N_14451);
xnor U14725 (N_14725,N_14527,N_14684);
nand U14726 (N_14726,N_14616,N_14665);
xnor U14727 (N_14727,N_14550,N_14576);
nand U14728 (N_14728,N_14509,N_14551);
or U14729 (N_14729,N_14456,N_14634);
xnor U14730 (N_14730,N_14419,N_14624);
and U14731 (N_14731,N_14528,N_14457);
and U14732 (N_14732,N_14587,N_14436);
and U14733 (N_14733,N_14429,N_14525);
xor U14734 (N_14734,N_14495,N_14638);
or U14735 (N_14735,N_14407,N_14575);
and U14736 (N_14736,N_14626,N_14516);
nand U14737 (N_14737,N_14449,N_14542);
and U14738 (N_14738,N_14416,N_14601);
and U14739 (N_14739,N_14435,N_14549);
nand U14740 (N_14740,N_14623,N_14517);
nand U14741 (N_14741,N_14481,N_14589);
or U14742 (N_14742,N_14668,N_14572);
nand U14743 (N_14743,N_14594,N_14673);
xnor U14744 (N_14744,N_14503,N_14539);
nor U14745 (N_14745,N_14484,N_14422);
or U14746 (N_14746,N_14679,N_14580);
xnor U14747 (N_14747,N_14605,N_14535);
nand U14748 (N_14748,N_14568,N_14671);
xnor U14749 (N_14749,N_14508,N_14531);
and U14750 (N_14750,N_14615,N_14467);
xnor U14751 (N_14751,N_14590,N_14440);
nor U14752 (N_14752,N_14413,N_14649);
nor U14753 (N_14753,N_14602,N_14524);
xor U14754 (N_14754,N_14658,N_14408);
xor U14755 (N_14755,N_14497,N_14667);
xor U14756 (N_14756,N_14574,N_14584);
nand U14757 (N_14757,N_14617,N_14653);
xnor U14758 (N_14758,N_14683,N_14657);
nor U14759 (N_14759,N_14678,N_14491);
and U14760 (N_14760,N_14635,N_14669);
or U14761 (N_14761,N_14444,N_14629);
or U14762 (N_14762,N_14465,N_14439);
or U14763 (N_14763,N_14695,N_14666);
and U14764 (N_14764,N_14418,N_14428);
nor U14765 (N_14765,N_14447,N_14489);
xnor U14766 (N_14766,N_14564,N_14619);
and U14767 (N_14767,N_14438,N_14530);
and U14768 (N_14768,N_14560,N_14488);
xor U14769 (N_14769,N_14504,N_14402);
xnor U14770 (N_14770,N_14515,N_14559);
nor U14771 (N_14771,N_14686,N_14696);
nor U14772 (N_14772,N_14681,N_14500);
nor U14773 (N_14773,N_14620,N_14687);
nor U14774 (N_14774,N_14582,N_14643);
xnor U14775 (N_14775,N_14557,N_14421);
nand U14776 (N_14776,N_14526,N_14403);
nor U14777 (N_14777,N_14431,N_14443);
nor U14778 (N_14778,N_14642,N_14406);
or U14779 (N_14779,N_14573,N_14563);
nor U14780 (N_14780,N_14663,N_14472);
xnor U14781 (N_14781,N_14511,N_14609);
and U14782 (N_14782,N_14697,N_14570);
nand U14783 (N_14783,N_14473,N_14485);
and U14784 (N_14784,N_14591,N_14478);
or U14785 (N_14785,N_14621,N_14654);
nand U14786 (N_14786,N_14676,N_14423);
nor U14787 (N_14787,N_14506,N_14401);
nand U14788 (N_14788,N_14510,N_14505);
and U14789 (N_14789,N_14538,N_14523);
xor U14790 (N_14790,N_14644,N_14434);
nand U14791 (N_14791,N_14534,N_14637);
nor U14792 (N_14792,N_14595,N_14417);
nor U14793 (N_14793,N_14566,N_14612);
and U14794 (N_14794,N_14533,N_14567);
or U14795 (N_14795,N_14630,N_14400);
nand U14796 (N_14796,N_14675,N_14420);
or U14797 (N_14797,N_14477,N_14588);
and U14798 (N_14798,N_14690,N_14618);
xnor U14799 (N_14799,N_14682,N_14544);
nand U14800 (N_14800,N_14520,N_14640);
and U14801 (N_14801,N_14655,N_14466);
xor U14802 (N_14802,N_14512,N_14448);
nand U14803 (N_14803,N_14433,N_14585);
xnor U14804 (N_14804,N_14441,N_14546);
xnor U14805 (N_14805,N_14558,N_14445);
and U14806 (N_14806,N_14479,N_14450);
and U14807 (N_14807,N_14583,N_14593);
nand U14808 (N_14808,N_14699,N_14604);
xnor U14809 (N_14809,N_14554,N_14656);
or U14810 (N_14810,N_14519,N_14670);
nor U14811 (N_14811,N_14645,N_14586);
nor U14812 (N_14812,N_14592,N_14646);
xor U14813 (N_14813,N_14536,N_14493);
or U14814 (N_14814,N_14636,N_14468);
nor U14815 (N_14815,N_14556,N_14562);
xor U14816 (N_14816,N_14461,N_14458);
or U14817 (N_14817,N_14685,N_14691);
and U14818 (N_14818,N_14555,N_14614);
nand U14819 (N_14819,N_14409,N_14659);
or U14820 (N_14820,N_14482,N_14514);
nand U14821 (N_14821,N_14577,N_14430);
nand U14822 (N_14822,N_14596,N_14628);
nand U14823 (N_14823,N_14641,N_14463);
nor U14824 (N_14824,N_14561,N_14688);
nor U14825 (N_14825,N_14693,N_14651);
xnor U14826 (N_14826,N_14677,N_14487);
or U14827 (N_14827,N_14661,N_14537);
nor U14828 (N_14828,N_14469,N_14427);
xnor U14829 (N_14829,N_14452,N_14600);
nand U14830 (N_14830,N_14664,N_14498);
nor U14831 (N_14831,N_14607,N_14608);
xor U14832 (N_14832,N_14480,N_14411);
nand U14833 (N_14833,N_14522,N_14648);
xnor U14834 (N_14834,N_14631,N_14545);
nor U14835 (N_14835,N_14404,N_14459);
or U14836 (N_14836,N_14553,N_14499);
or U14837 (N_14837,N_14552,N_14490);
or U14838 (N_14838,N_14613,N_14694);
xor U14839 (N_14839,N_14437,N_14647);
or U14840 (N_14840,N_14496,N_14565);
nor U14841 (N_14841,N_14412,N_14611);
nand U14842 (N_14842,N_14464,N_14569);
xor U14843 (N_14843,N_14578,N_14547);
nand U14844 (N_14844,N_14660,N_14414);
and U14845 (N_14845,N_14486,N_14474);
and U14846 (N_14846,N_14529,N_14475);
nand U14847 (N_14847,N_14672,N_14632);
or U14848 (N_14848,N_14680,N_14603);
or U14849 (N_14849,N_14471,N_14405);
nand U14850 (N_14850,N_14589,N_14534);
xor U14851 (N_14851,N_14565,N_14651);
nor U14852 (N_14852,N_14624,N_14417);
nand U14853 (N_14853,N_14699,N_14616);
or U14854 (N_14854,N_14582,N_14591);
or U14855 (N_14855,N_14537,N_14548);
or U14856 (N_14856,N_14615,N_14528);
or U14857 (N_14857,N_14539,N_14406);
xnor U14858 (N_14858,N_14485,N_14628);
and U14859 (N_14859,N_14633,N_14603);
and U14860 (N_14860,N_14581,N_14495);
nand U14861 (N_14861,N_14699,N_14608);
and U14862 (N_14862,N_14649,N_14559);
and U14863 (N_14863,N_14684,N_14507);
or U14864 (N_14864,N_14640,N_14653);
nor U14865 (N_14865,N_14673,N_14600);
nand U14866 (N_14866,N_14425,N_14520);
or U14867 (N_14867,N_14652,N_14429);
nand U14868 (N_14868,N_14438,N_14649);
xor U14869 (N_14869,N_14509,N_14552);
nand U14870 (N_14870,N_14510,N_14427);
or U14871 (N_14871,N_14666,N_14418);
nand U14872 (N_14872,N_14657,N_14675);
and U14873 (N_14873,N_14691,N_14564);
xor U14874 (N_14874,N_14434,N_14532);
xor U14875 (N_14875,N_14466,N_14638);
nor U14876 (N_14876,N_14500,N_14443);
nor U14877 (N_14877,N_14584,N_14510);
nor U14878 (N_14878,N_14478,N_14420);
or U14879 (N_14879,N_14434,N_14542);
nand U14880 (N_14880,N_14671,N_14529);
and U14881 (N_14881,N_14405,N_14589);
and U14882 (N_14882,N_14689,N_14683);
nand U14883 (N_14883,N_14467,N_14442);
or U14884 (N_14884,N_14421,N_14612);
nor U14885 (N_14885,N_14502,N_14506);
nor U14886 (N_14886,N_14689,N_14662);
xor U14887 (N_14887,N_14533,N_14457);
nor U14888 (N_14888,N_14628,N_14431);
nand U14889 (N_14889,N_14641,N_14584);
and U14890 (N_14890,N_14691,N_14533);
nor U14891 (N_14891,N_14457,N_14456);
and U14892 (N_14892,N_14678,N_14535);
nand U14893 (N_14893,N_14483,N_14436);
and U14894 (N_14894,N_14650,N_14498);
nand U14895 (N_14895,N_14560,N_14503);
or U14896 (N_14896,N_14690,N_14459);
nand U14897 (N_14897,N_14581,N_14591);
nor U14898 (N_14898,N_14600,N_14544);
xnor U14899 (N_14899,N_14644,N_14440);
nor U14900 (N_14900,N_14698,N_14531);
nor U14901 (N_14901,N_14532,N_14527);
or U14902 (N_14902,N_14640,N_14541);
or U14903 (N_14903,N_14690,N_14539);
and U14904 (N_14904,N_14485,N_14463);
nand U14905 (N_14905,N_14536,N_14610);
nand U14906 (N_14906,N_14482,N_14683);
xnor U14907 (N_14907,N_14499,N_14485);
or U14908 (N_14908,N_14465,N_14610);
nor U14909 (N_14909,N_14555,N_14682);
or U14910 (N_14910,N_14530,N_14636);
nand U14911 (N_14911,N_14494,N_14508);
nor U14912 (N_14912,N_14668,N_14691);
nand U14913 (N_14913,N_14543,N_14676);
nor U14914 (N_14914,N_14585,N_14566);
xor U14915 (N_14915,N_14513,N_14583);
nor U14916 (N_14916,N_14652,N_14615);
nor U14917 (N_14917,N_14424,N_14689);
or U14918 (N_14918,N_14585,N_14554);
nor U14919 (N_14919,N_14556,N_14458);
nor U14920 (N_14920,N_14500,N_14496);
and U14921 (N_14921,N_14574,N_14549);
nor U14922 (N_14922,N_14513,N_14438);
nand U14923 (N_14923,N_14509,N_14433);
nor U14924 (N_14924,N_14465,N_14584);
or U14925 (N_14925,N_14688,N_14527);
or U14926 (N_14926,N_14611,N_14463);
or U14927 (N_14927,N_14576,N_14667);
and U14928 (N_14928,N_14596,N_14561);
xor U14929 (N_14929,N_14656,N_14508);
and U14930 (N_14930,N_14500,N_14592);
nand U14931 (N_14931,N_14508,N_14642);
nand U14932 (N_14932,N_14644,N_14485);
nand U14933 (N_14933,N_14438,N_14610);
or U14934 (N_14934,N_14523,N_14413);
nor U14935 (N_14935,N_14651,N_14654);
and U14936 (N_14936,N_14683,N_14445);
or U14937 (N_14937,N_14657,N_14536);
or U14938 (N_14938,N_14494,N_14604);
or U14939 (N_14939,N_14426,N_14429);
nor U14940 (N_14940,N_14520,N_14611);
and U14941 (N_14941,N_14626,N_14688);
nor U14942 (N_14942,N_14502,N_14620);
and U14943 (N_14943,N_14522,N_14414);
xor U14944 (N_14944,N_14591,N_14614);
or U14945 (N_14945,N_14699,N_14670);
and U14946 (N_14946,N_14554,N_14506);
nand U14947 (N_14947,N_14403,N_14553);
xnor U14948 (N_14948,N_14666,N_14419);
nor U14949 (N_14949,N_14660,N_14542);
or U14950 (N_14950,N_14677,N_14468);
and U14951 (N_14951,N_14627,N_14458);
and U14952 (N_14952,N_14544,N_14474);
and U14953 (N_14953,N_14647,N_14483);
and U14954 (N_14954,N_14451,N_14621);
nor U14955 (N_14955,N_14527,N_14622);
and U14956 (N_14956,N_14526,N_14663);
nand U14957 (N_14957,N_14580,N_14641);
xor U14958 (N_14958,N_14668,N_14596);
nand U14959 (N_14959,N_14523,N_14567);
xnor U14960 (N_14960,N_14452,N_14408);
nand U14961 (N_14961,N_14565,N_14481);
nor U14962 (N_14962,N_14473,N_14679);
or U14963 (N_14963,N_14458,N_14678);
and U14964 (N_14964,N_14679,N_14437);
nor U14965 (N_14965,N_14655,N_14491);
xor U14966 (N_14966,N_14630,N_14421);
and U14967 (N_14967,N_14419,N_14539);
xor U14968 (N_14968,N_14408,N_14558);
nand U14969 (N_14969,N_14679,N_14648);
xnor U14970 (N_14970,N_14508,N_14635);
or U14971 (N_14971,N_14688,N_14643);
nand U14972 (N_14972,N_14644,N_14667);
and U14973 (N_14973,N_14536,N_14484);
and U14974 (N_14974,N_14543,N_14649);
nor U14975 (N_14975,N_14692,N_14673);
nand U14976 (N_14976,N_14639,N_14469);
nor U14977 (N_14977,N_14591,N_14510);
xnor U14978 (N_14978,N_14594,N_14606);
nor U14979 (N_14979,N_14667,N_14627);
or U14980 (N_14980,N_14596,N_14469);
nand U14981 (N_14981,N_14689,N_14459);
nor U14982 (N_14982,N_14570,N_14615);
xor U14983 (N_14983,N_14517,N_14427);
nor U14984 (N_14984,N_14596,N_14486);
or U14985 (N_14985,N_14678,N_14453);
or U14986 (N_14986,N_14680,N_14696);
nand U14987 (N_14987,N_14513,N_14564);
nor U14988 (N_14988,N_14502,N_14405);
nand U14989 (N_14989,N_14444,N_14520);
nor U14990 (N_14990,N_14645,N_14494);
xnor U14991 (N_14991,N_14582,N_14430);
and U14992 (N_14992,N_14498,N_14545);
or U14993 (N_14993,N_14565,N_14650);
and U14994 (N_14994,N_14564,N_14697);
nor U14995 (N_14995,N_14488,N_14688);
xnor U14996 (N_14996,N_14644,N_14632);
nand U14997 (N_14997,N_14446,N_14580);
nor U14998 (N_14998,N_14484,N_14472);
or U14999 (N_14999,N_14458,N_14614);
and UO_0 (O_0,N_14954,N_14710);
nor UO_1 (O_1,N_14856,N_14817);
and UO_2 (O_2,N_14712,N_14792);
and UO_3 (O_3,N_14744,N_14759);
xnor UO_4 (O_4,N_14861,N_14715);
xnor UO_5 (O_5,N_14998,N_14776);
nor UO_6 (O_6,N_14769,N_14795);
or UO_7 (O_7,N_14873,N_14900);
or UO_8 (O_8,N_14868,N_14944);
xnor UO_9 (O_9,N_14791,N_14870);
xnor UO_10 (O_10,N_14849,N_14837);
and UO_11 (O_11,N_14888,N_14717);
nand UO_12 (O_12,N_14863,N_14765);
or UO_13 (O_13,N_14726,N_14799);
xnor UO_14 (O_14,N_14818,N_14939);
nor UO_15 (O_15,N_14931,N_14794);
xnor UO_16 (O_16,N_14806,N_14842);
xnor UO_17 (O_17,N_14737,N_14831);
xor UO_18 (O_18,N_14902,N_14993);
or UO_19 (O_19,N_14956,N_14908);
and UO_20 (O_20,N_14760,N_14735);
xnor UO_21 (O_21,N_14946,N_14814);
nand UO_22 (O_22,N_14730,N_14921);
xor UO_23 (O_23,N_14770,N_14941);
xor UO_24 (O_24,N_14723,N_14816);
nand UO_25 (O_25,N_14811,N_14906);
and UO_26 (O_26,N_14968,N_14739);
nand UO_27 (O_27,N_14777,N_14729);
and UO_28 (O_28,N_14854,N_14898);
and UO_29 (O_29,N_14766,N_14706);
and UO_30 (O_30,N_14901,N_14882);
xnor UO_31 (O_31,N_14787,N_14962);
xnor UO_32 (O_32,N_14820,N_14878);
xnor UO_33 (O_33,N_14858,N_14793);
nor UO_34 (O_34,N_14782,N_14978);
xor UO_35 (O_35,N_14815,N_14952);
and UO_36 (O_36,N_14913,N_14757);
or UO_37 (O_37,N_14753,N_14788);
xnor UO_38 (O_38,N_14992,N_14751);
or UO_39 (O_39,N_14948,N_14876);
nand UO_40 (O_40,N_14745,N_14994);
or UO_41 (O_41,N_14862,N_14713);
or UO_42 (O_42,N_14724,N_14988);
nand UO_43 (O_43,N_14722,N_14890);
nand UO_44 (O_44,N_14918,N_14860);
nor UO_45 (O_45,N_14971,N_14927);
and UO_46 (O_46,N_14880,N_14865);
nand UO_47 (O_47,N_14775,N_14986);
and UO_48 (O_48,N_14917,N_14938);
or UO_49 (O_49,N_14984,N_14711);
or UO_50 (O_50,N_14910,N_14989);
nor UO_51 (O_51,N_14852,N_14881);
and UO_52 (O_52,N_14889,N_14884);
xor UO_53 (O_53,N_14920,N_14975);
and UO_54 (O_54,N_14802,N_14924);
nor UO_55 (O_55,N_14701,N_14841);
nand UO_56 (O_56,N_14976,N_14705);
xnor UO_57 (O_57,N_14801,N_14909);
or UO_58 (O_58,N_14828,N_14821);
nor UO_59 (O_59,N_14797,N_14812);
or UO_60 (O_60,N_14961,N_14869);
or UO_61 (O_61,N_14859,N_14747);
nor UO_62 (O_62,N_14982,N_14707);
and UO_63 (O_63,N_14825,N_14926);
and UO_64 (O_64,N_14995,N_14919);
nand UO_65 (O_65,N_14768,N_14979);
or UO_66 (O_66,N_14779,N_14819);
nor UO_67 (O_67,N_14830,N_14848);
nor UO_68 (O_68,N_14959,N_14991);
nand UO_69 (O_69,N_14762,N_14877);
nor UO_70 (O_70,N_14960,N_14704);
or UO_71 (O_71,N_14951,N_14923);
and UO_72 (O_72,N_14969,N_14839);
nand UO_73 (O_73,N_14866,N_14864);
nand UO_74 (O_74,N_14851,N_14936);
or UO_75 (O_75,N_14955,N_14703);
and UO_76 (O_76,N_14754,N_14785);
xor UO_77 (O_77,N_14824,N_14702);
and UO_78 (O_78,N_14823,N_14846);
nand UO_79 (O_79,N_14734,N_14980);
nand UO_80 (O_80,N_14829,N_14727);
nand UO_81 (O_81,N_14749,N_14790);
or UO_82 (O_82,N_14891,N_14965);
and UO_83 (O_83,N_14832,N_14725);
and UO_84 (O_84,N_14748,N_14855);
or UO_85 (O_85,N_14853,N_14700);
nor UO_86 (O_86,N_14930,N_14763);
nand UO_87 (O_87,N_14983,N_14987);
or UO_88 (O_88,N_14718,N_14732);
or UO_89 (O_89,N_14928,N_14741);
nor UO_90 (O_90,N_14997,N_14772);
and UO_91 (O_91,N_14714,N_14963);
and UO_92 (O_92,N_14774,N_14733);
xor UO_93 (O_93,N_14874,N_14835);
xor UO_94 (O_94,N_14771,N_14950);
xnor UO_95 (O_95,N_14742,N_14778);
and UO_96 (O_96,N_14721,N_14808);
or UO_97 (O_97,N_14949,N_14847);
or UO_98 (O_98,N_14905,N_14767);
nor UO_99 (O_99,N_14780,N_14844);
xnor UO_100 (O_100,N_14999,N_14807);
or UO_101 (O_101,N_14892,N_14916);
and UO_102 (O_102,N_14789,N_14897);
nand UO_103 (O_103,N_14929,N_14894);
nand UO_104 (O_104,N_14758,N_14940);
nor UO_105 (O_105,N_14904,N_14925);
nor UO_106 (O_106,N_14893,N_14738);
nor UO_107 (O_107,N_14945,N_14843);
xnor UO_108 (O_108,N_14761,N_14899);
nor UO_109 (O_109,N_14895,N_14716);
and UO_110 (O_110,N_14784,N_14903);
nand UO_111 (O_111,N_14964,N_14786);
or UO_112 (O_112,N_14834,N_14755);
xor UO_113 (O_113,N_14883,N_14708);
or UO_114 (O_114,N_14958,N_14875);
xnor UO_115 (O_115,N_14990,N_14886);
xnor UO_116 (O_116,N_14957,N_14934);
nand UO_117 (O_117,N_14709,N_14872);
nor UO_118 (O_118,N_14798,N_14809);
nor UO_119 (O_119,N_14915,N_14827);
nand UO_120 (O_120,N_14731,N_14887);
or UO_121 (O_121,N_14996,N_14836);
and UO_122 (O_122,N_14935,N_14746);
or UO_123 (O_123,N_14740,N_14728);
xnor UO_124 (O_124,N_14750,N_14764);
and UO_125 (O_125,N_14850,N_14783);
or UO_126 (O_126,N_14867,N_14833);
nand UO_127 (O_127,N_14879,N_14813);
nand UO_128 (O_128,N_14736,N_14911);
nand UO_129 (O_129,N_14985,N_14810);
or UO_130 (O_130,N_14773,N_14974);
nor UO_131 (O_131,N_14932,N_14967);
nand UO_132 (O_132,N_14973,N_14896);
nor UO_133 (O_133,N_14752,N_14803);
xor UO_134 (O_134,N_14838,N_14937);
and UO_135 (O_135,N_14720,N_14977);
nor UO_136 (O_136,N_14943,N_14719);
nand UO_137 (O_137,N_14914,N_14781);
nor UO_138 (O_138,N_14743,N_14826);
or UO_139 (O_139,N_14966,N_14907);
xnor UO_140 (O_140,N_14845,N_14942);
nor UO_141 (O_141,N_14981,N_14871);
and UO_142 (O_142,N_14972,N_14857);
xnor UO_143 (O_143,N_14756,N_14922);
and UO_144 (O_144,N_14947,N_14885);
xnor UO_145 (O_145,N_14953,N_14804);
or UO_146 (O_146,N_14933,N_14800);
or UO_147 (O_147,N_14796,N_14912);
or UO_148 (O_148,N_14822,N_14840);
nand UO_149 (O_149,N_14805,N_14970);
xor UO_150 (O_150,N_14884,N_14833);
and UO_151 (O_151,N_14870,N_14731);
and UO_152 (O_152,N_14788,N_14930);
xnor UO_153 (O_153,N_14804,N_14770);
and UO_154 (O_154,N_14931,N_14985);
and UO_155 (O_155,N_14823,N_14866);
xnor UO_156 (O_156,N_14765,N_14917);
nand UO_157 (O_157,N_14789,N_14975);
nand UO_158 (O_158,N_14957,N_14791);
and UO_159 (O_159,N_14943,N_14775);
nor UO_160 (O_160,N_14927,N_14929);
xnor UO_161 (O_161,N_14758,N_14871);
xnor UO_162 (O_162,N_14944,N_14927);
xnor UO_163 (O_163,N_14925,N_14724);
and UO_164 (O_164,N_14768,N_14706);
xor UO_165 (O_165,N_14732,N_14727);
xnor UO_166 (O_166,N_14767,N_14966);
and UO_167 (O_167,N_14854,N_14822);
xor UO_168 (O_168,N_14739,N_14916);
nand UO_169 (O_169,N_14768,N_14960);
nor UO_170 (O_170,N_14884,N_14735);
xor UO_171 (O_171,N_14819,N_14776);
xor UO_172 (O_172,N_14727,N_14823);
nand UO_173 (O_173,N_14839,N_14707);
nor UO_174 (O_174,N_14998,N_14804);
nor UO_175 (O_175,N_14730,N_14968);
nor UO_176 (O_176,N_14766,N_14713);
or UO_177 (O_177,N_14869,N_14933);
or UO_178 (O_178,N_14949,N_14857);
and UO_179 (O_179,N_14723,N_14796);
or UO_180 (O_180,N_14789,N_14925);
and UO_181 (O_181,N_14971,N_14930);
and UO_182 (O_182,N_14986,N_14818);
nand UO_183 (O_183,N_14810,N_14823);
and UO_184 (O_184,N_14918,N_14781);
nor UO_185 (O_185,N_14751,N_14885);
or UO_186 (O_186,N_14776,N_14772);
and UO_187 (O_187,N_14748,N_14981);
nand UO_188 (O_188,N_14810,N_14908);
or UO_189 (O_189,N_14879,N_14886);
or UO_190 (O_190,N_14863,N_14984);
nand UO_191 (O_191,N_14868,N_14863);
nand UO_192 (O_192,N_14757,N_14751);
xor UO_193 (O_193,N_14920,N_14870);
nor UO_194 (O_194,N_14887,N_14875);
and UO_195 (O_195,N_14845,N_14755);
nor UO_196 (O_196,N_14981,N_14815);
nor UO_197 (O_197,N_14868,N_14949);
and UO_198 (O_198,N_14860,N_14839);
xor UO_199 (O_199,N_14776,N_14798);
xnor UO_200 (O_200,N_14891,N_14909);
nor UO_201 (O_201,N_14851,N_14764);
and UO_202 (O_202,N_14890,N_14811);
or UO_203 (O_203,N_14954,N_14828);
and UO_204 (O_204,N_14751,N_14977);
xnor UO_205 (O_205,N_14922,N_14774);
xor UO_206 (O_206,N_14866,N_14970);
and UO_207 (O_207,N_14715,N_14964);
nand UO_208 (O_208,N_14833,N_14958);
nor UO_209 (O_209,N_14801,N_14835);
xnor UO_210 (O_210,N_14823,N_14773);
nor UO_211 (O_211,N_14776,N_14978);
nor UO_212 (O_212,N_14917,N_14968);
xor UO_213 (O_213,N_14886,N_14758);
nor UO_214 (O_214,N_14858,N_14788);
or UO_215 (O_215,N_14886,N_14882);
and UO_216 (O_216,N_14762,N_14934);
xnor UO_217 (O_217,N_14879,N_14745);
and UO_218 (O_218,N_14836,N_14861);
nor UO_219 (O_219,N_14881,N_14912);
nand UO_220 (O_220,N_14845,N_14876);
nand UO_221 (O_221,N_14906,N_14872);
nor UO_222 (O_222,N_14825,N_14921);
or UO_223 (O_223,N_14986,N_14910);
xor UO_224 (O_224,N_14949,N_14928);
or UO_225 (O_225,N_14970,N_14916);
or UO_226 (O_226,N_14949,N_14782);
nand UO_227 (O_227,N_14819,N_14932);
and UO_228 (O_228,N_14834,N_14941);
xor UO_229 (O_229,N_14978,N_14991);
or UO_230 (O_230,N_14816,N_14764);
nor UO_231 (O_231,N_14971,N_14777);
or UO_232 (O_232,N_14913,N_14812);
nor UO_233 (O_233,N_14796,N_14704);
and UO_234 (O_234,N_14880,N_14748);
or UO_235 (O_235,N_14793,N_14832);
and UO_236 (O_236,N_14899,N_14938);
and UO_237 (O_237,N_14911,N_14830);
xnor UO_238 (O_238,N_14738,N_14751);
and UO_239 (O_239,N_14878,N_14838);
nand UO_240 (O_240,N_14878,N_14711);
nor UO_241 (O_241,N_14703,N_14726);
nand UO_242 (O_242,N_14824,N_14783);
and UO_243 (O_243,N_14962,N_14952);
and UO_244 (O_244,N_14998,N_14722);
or UO_245 (O_245,N_14795,N_14808);
nor UO_246 (O_246,N_14845,N_14861);
and UO_247 (O_247,N_14743,N_14926);
and UO_248 (O_248,N_14990,N_14859);
nor UO_249 (O_249,N_14831,N_14912);
and UO_250 (O_250,N_14788,N_14834);
xnor UO_251 (O_251,N_14919,N_14747);
or UO_252 (O_252,N_14718,N_14986);
xnor UO_253 (O_253,N_14914,N_14721);
and UO_254 (O_254,N_14712,N_14829);
xnor UO_255 (O_255,N_14853,N_14945);
and UO_256 (O_256,N_14999,N_14991);
or UO_257 (O_257,N_14865,N_14748);
xnor UO_258 (O_258,N_14847,N_14990);
nand UO_259 (O_259,N_14973,N_14986);
and UO_260 (O_260,N_14921,N_14799);
nor UO_261 (O_261,N_14882,N_14954);
or UO_262 (O_262,N_14951,N_14998);
nand UO_263 (O_263,N_14952,N_14987);
nand UO_264 (O_264,N_14908,N_14928);
nor UO_265 (O_265,N_14996,N_14892);
nor UO_266 (O_266,N_14778,N_14704);
nor UO_267 (O_267,N_14867,N_14946);
nor UO_268 (O_268,N_14832,N_14701);
nor UO_269 (O_269,N_14747,N_14865);
or UO_270 (O_270,N_14899,N_14742);
xor UO_271 (O_271,N_14803,N_14866);
xnor UO_272 (O_272,N_14982,N_14774);
nor UO_273 (O_273,N_14752,N_14819);
xor UO_274 (O_274,N_14976,N_14791);
nor UO_275 (O_275,N_14862,N_14895);
and UO_276 (O_276,N_14923,N_14881);
and UO_277 (O_277,N_14894,N_14716);
xor UO_278 (O_278,N_14777,N_14722);
nand UO_279 (O_279,N_14894,N_14877);
and UO_280 (O_280,N_14918,N_14811);
nand UO_281 (O_281,N_14931,N_14875);
or UO_282 (O_282,N_14949,N_14824);
nand UO_283 (O_283,N_14851,N_14813);
or UO_284 (O_284,N_14903,N_14778);
xor UO_285 (O_285,N_14751,N_14998);
or UO_286 (O_286,N_14871,N_14817);
and UO_287 (O_287,N_14889,N_14851);
nor UO_288 (O_288,N_14946,N_14968);
or UO_289 (O_289,N_14933,N_14718);
nand UO_290 (O_290,N_14927,N_14785);
nor UO_291 (O_291,N_14992,N_14748);
or UO_292 (O_292,N_14994,N_14883);
or UO_293 (O_293,N_14798,N_14911);
nor UO_294 (O_294,N_14723,N_14785);
or UO_295 (O_295,N_14950,N_14936);
xor UO_296 (O_296,N_14801,N_14953);
nand UO_297 (O_297,N_14921,N_14781);
xnor UO_298 (O_298,N_14749,N_14890);
nand UO_299 (O_299,N_14839,N_14943);
and UO_300 (O_300,N_14886,N_14747);
nor UO_301 (O_301,N_14828,N_14912);
nor UO_302 (O_302,N_14857,N_14999);
nor UO_303 (O_303,N_14844,N_14786);
and UO_304 (O_304,N_14752,N_14756);
nand UO_305 (O_305,N_14907,N_14854);
and UO_306 (O_306,N_14732,N_14853);
and UO_307 (O_307,N_14934,N_14757);
nand UO_308 (O_308,N_14828,N_14745);
or UO_309 (O_309,N_14960,N_14743);
nand UO_310 (O_310,N_14972,N_14899);
nand UO_311 (O_311,N_14709,N_14988);
and UO_312 (O_312,N_14728,N_14787);
nand UO_313 (O_313,N_14834,N_14935);
nor UO_314 (O_314,N_14904,N_14713);
xor UO_315 (O_315,N_14995,N_14894);
or UO_316 (O_316,N_14796,N_14863);
nor UO_317 (O_317,N_14786,N_14960);
nand UO_318 (O_318,N_14768,N_14875);
nor UO_319 (O_319,N_14729,N_14956);
nor UO_320 (O_320,N_14900,N_14757);
nor UO_321 (O_321,N_14966,N_14935);
nand UO_322 (O_322,N_14714,N_14929);
nand UO_323 (O_323,N_14865,N_14716);
nor UO_324 (O_324,N_14725,N_14871);
xnor UO_325 (O_325,N_14972,N_14725);
and UO_326 (O_326,N_14905,N_14881);
xnor UO_327 (O_327,N_14943,N_14737);
nand UO_328 (O_328,N_14952,N_14766);
nand UO_329 (O_329,N_14900,N_14722);
nand UO_330 (O_330,N_14802,N_14704);
or UO_331 (O_331,N_14991,N_14976);
nand UO_332 (O_332,N_14916,N_14846);
and UO_333 (O_333,N_14778,N_14799);
xor UO_334 (O_334,N_14789,N_14862);
xnor UO_335 (O_335,N_14994,N_14869);
or UO_336 (O_336,N_14774,N_14889);
nand UO_337 (O_337,N_14774,N_14744);
nor UO_338 (O_338,N_14835,N_14717);
nand UO_339 (O_339,N_14922,N_14853);
and UO_340 (O_340,N_14835,N_14962);
or UO_341 (O_341,N_14759,N_14785);
or UO_342 (O_342,N_14964,N_14710);
or UO_343 (O_343,N_14742,N_14736);
and UO_344 (O_344,N_14738,N_14736);
xor UO_345 (O_345,N_14866,N_14778);
and UO_346 (O_346,N_14980,N_14908);
or UO_347 (O_347,N_14738,N_14968);
nand UO_348 (O_348,N_14938,N_14742);
and UO_349 (O_349,N_14993,N_14839);
or UO_350 (O_350,N_14873,N_14937);
xnor UO_351 (O_351,N_14861,N_14868);
xor UO_352 (O_352,N_14895,N_14999);
nand UO_353 (O_353,N_14707,N_14916);
nor UO_354 (O_354,N_14975,N_14964);
and UO_355 (O_355,N_14741,N_14745);
nand UO_356 (O_356,N_14783,N_14956);
xor UO_357 (O_357,N_14913,N_14713);
and UO_358 (O_358,N_14817,N_14727);
or UO_359 (O_359,N_14860,N_14768);
xor UO_360 (O_360,N_14762,N_14907);
nor UO_361 (O_361,N_14742,N_14963);
xnor UO_362 (O_362,N_14824,N_14933);
and UO_363 (O_363,N_14975,N_14738);
nor UO_364 (O_364,N_14997,N_14967);
xor UO_365 (O_365,N_14752,N_14839);
and UO_366 (O_366,N_14785,N_14813);
nor UO_367 (O_367,N_14849,N_14909);
and UO_368 (O_368,N_14968,N_14808);
xor UO_369 (O_369,N_14857,N_14983);
nand UO_370 (O_370,N_14756,N_14936);
xnor UO_371 (O_371,N_14892,N_14733);
or UO_372 (O_372,N_14887,N_14914);
xnor UO_373 (O_373,N_14961,N_14995);
xnor UO_374 (O_374,N_14945,N_14993);
nor UO_375 (O_375,N_14954,N_14984);
nand UO_376 (O_376,N_14734,N_14700);
or UO_377 (O_377,N_14759,N_14732);
xor UO_378 (O_378,N_14789,N_14710);
nand UO_379 (O_379,N_14737,N_14847);
or UO_380 (O_380,N_14952,N_14830);
nand UO_381 (O_381,N_14823,N_14887);
and UO_382 (O_382,N_14933,N_14924);
and UO_383 (O_383,N_14741,N_14926);
and UO_384 (O_384,N_14866,N_14755);
nand UO_385 (O_385,N_14973,N_14868);
or UO_386 (O_386,N_14872,N_14949);
nor UO_387 (O_387,N_14839,N_14956);
nor UO_388 (O_388,N_14762,N_14983);
and UO_389 (O_389,N_14743,N_14787);
nand UO_390 (O_390,N_14721,N_14990);
nor UO_391 (O_391,N_14781,N_14730);
nor UO_392 (O_392,N_14791,N_14919);
nand UO_393 (O_393,N_14908,N_14945);
nor UO_394 (O_394,N_14980,N_14827);
and UO_395 (O_395,N_14783,N_14740);
xnor UO_396 (O_396,N_14792,N_14803);
nor UO_397 (O_397,N_14998,N_14948);
nor UO_398 (O_398,N_14968,N_14799);
nand UO_399 (O_399,N_14935,N_14921);
and UO_400 (O_400,N_14978,N_14912);
nand UO_401 (O_401,N_14915,N_14843);
xnor UO_402 (O_402,N_14950,N_14720);
nand UO_403 (O_403,N_14972,N_14911);
or UO_404 (O_404,N_14817,N_14818);
nand UO_405 (O_405,N_14930,N_14982);
nand UO_406 (O_406,N_14782,N_14952);
and UO_407 (O_407,N_14884,N_14725);
or UO_408 (O_408,N_14999,N_14773);
xor UO_409 (O_409,N_14779,N_14828);
nand UO_410 (O_410,N_14709,N_14738);
and UO_411 (O_411,N_14709,N_14776);
or UO_412 (O_412,N_14959,N_14876);
nand UO_413 (O_413,N_14884,N_14771);
nand UO_414 (O_414,N_14834,N_14801);
or UO_415 (O_415,N_14755,N_14736);
and UO_416 (O_416,N_14766,N_14712);
nand UO_417 (O_417,N_14880,N_14964);
nor UO_418 (O_418,N_14860,N_14794);
nor UO_419 (O_419,N_14720,N_14703);
xor UO_420 (O_420,N_14709,N_14735);
nor UO_421 (O_421,N_14957,N_14762);
xor UO_422 (O_422,N_14726,N_14915);
xnor UO_423 (O_423,N_14826,N_14907);
nor UO_424 (O_424,N_14848,N_14798);
and UO_425 (O_425,N_14858,N_14893);
and UO_426 (O_426,N_14742,N_14861);
or UO_427 (O_427,N_14701,N_14970);
xnor UO_428 (O_428,N_14743,N_14812);
nand UO_429 (O_429,N_14716,N_14977);
and UO_430 (O_430,N_14773,N_14879);
nand UO_431 (O_431,N_14829,N_14797);
or UO_432 (O_432,N_14855,N_14793);
nor UO_433 (O_433,N_14987,N_14891);
xor UO_434 (O_434,N_14959,N_14750);
nor UO_435 (O_435,N_14756,N_14820);
xnor UO_436 (O_436,N_14996,N_14735);
nand UO_437 (O_437,N_14841,N_14822);
nand UO_438 (O_438,N_14937,N_14821);
xor UO_439 (O_439,N_14730,N_14995);
and UO_440 (O_440,N_14953,N_14731);
and UO_441 (O_441,N_14911,N_14809);
nor UO_442 (O_442,N_14718,N_14970);
or UO_443 (O_443,N_14736,N_14760);
xor UO_444 (O_444,N_14852,N_14865);
nand UO_445 (O_445,N_14902,N_14937);
nor UO_446 (O_446,N_14800,N_14766);
and UO_447 (O_447,N_14881,N_14756);
xor UO_448 (O_448,N_14802,N_14831);
and UO_449 (O_449,N_14766,N_14703);
xnor UO_450 (O_450,N_14769,N_14721);
nand UO_451 (O_451,N_14849,N_14861);
nor UO_452 (O_452,N_14995,N_14832);
and UO_453 (O_453,N_14890,N_14888);
nor UO_454 (O_454,N_14737,N_14983);
nand UO_455 (O_455,N_14985,N_14803);
nand UO_456 (O_456,N_14768,N_14799);
xor UO_457 (O_457,N_14938,N_14738);
xor UO_458 (O_458,N_14715,N_14959);
xnor UO_459 (O_459,N_14981,N_14781);
nand UO_460 (O_460,N_14736,N_14794);
nor UO_461 (O_461,N_14909,N_14866);
or UO_462 (O_462,N_14828,N_14713);
or UO_463 (O_463,N_14916,N_14871);
xnor UO_464 (O_464,N_14730,N_14793);
nand UO_465 (O_465,N_14934,N_14996);
nand UO_466 (O_466,N_14865,N_14972);
nor UO_467 (O_467,N_14975,N_14870);
nor UO_468 (O_468,N_14921,N_14803);
nor UO_469 (O_469,N_14857,N_14882);
nor UO_470 (O_470,N_14864,N_14739);
nor UO_471 (O_471,N_14865,N_14841);
or UO_472 (O_472,N_14955,N_14929);
or UO_473 (O_473,N_14884,N_14830);
nand UO_474 (O_474,N_14868,N_14947);
and UO_475 (O_475,N_14936,N_14967);
nor UO_476 (O_476,N_14899,N_14753);
nand UO_477 (O_477,N_14801,N_14969);
nand UO_478 (O_478,N_14972,N_14738);
nand UO_479 (O_479,N_14975,N_14865);
nand UO_480 (O_480,N_14904,N_14707);
or UO_481 (O_481,N_14734,N_14787);
or UO_482 (O_482,N_14965,N_14883);
or UO_483 (O_483,N_14756,N_14773);
nand UO_484 (O_484,N_14973,N_14920);
or UO_485 (O_485,N_14865,N_14809);
or UO_486 (O_486,N_14711,N_14954);
nor UO_487 (O_487,N_14860,N_14837);
and UO_488 (O_488,N_14882,N_14759);
nand UO_489 (O_489,N_14906,N_14764);
nor UO_490 (O_490,N_14826,N_14723);
or UO_491 (O_491,N_14912,N_14920);
or UO_492 (O_492,N_14722,N_14992);
xor UO_493 (O_493,N_14884,N_14834);
or UO_494 (O_494,N_14974,N_14931);
xnor UO_495 (O_495,N_14828,N_14965);
or UO_496 (O_496,N_14732,N_14719);
xnor UO_497 (O_497,N_14881,N_14806);
or UO_498 (O_498,N_14849,N_14811);
and UO_499 (O_499,N_14756,N_14728);
nor UO_500 (O_500,N_14761,N_14923);
and UO_501 (O_501,N_14802,N_14970);
nand UO_502 (O_502,N_14858,N_14927);
nand UO_503 (O_503,N_14931,N_14978);
nor UO_504 (O_504,N_14843,N_14802);
nand UO_505 (O_505,N_14734,N_14753);
nor UO_506 (O_506,N_14790,N_14827);
nor UO_507 (O_507,N_14737,N_14900);
or UO_508 (O_508,N_14961,N_14724);
xnor UO_509 (O_509,N_14728,N_14749);
and UO_510 (O_510,N_14978,N_14775);
and UO_511 (O_511,N_14743,N_14871);
nand UO_512 (O_512,N_14938,N_14724);
xnor UO_513 (O_513,N_14754,N_14903);
or UO_514 (O_514,N_14867,N_14737);
nor UO_515 (O_515,N_14745,N_14742);
nor UO_516 (O_516,N_14940,N_14767);
xnor UO_517 (O_517,N_14791,N_14814);
nand UO_518 (O_518,N_14943,N_14832);
nand UO_519 (O_519,N_14920,N_14710);
and UO_520 (O_520,N_14888,N_14991);
xnor UO_521 (O_521,N_14940,N_14746);
nor UO_522 (O_522,N_14761,N_14910);
or UO_523 (O_523,N_14878,N_14813);
and UO_524 (O_524,N_14738,N_14943);
nor UO_525 (O_525,N_14874,N_14893);
nand UO_526 (O_526,N_14848,N_14847);
nor UO_527 (O_527,N_14896,N_14800);
nand UO_528 (O_528,N_14776,N_14823);
or UO_529 (O_529,N_14962,N_14939);
xor UO_530 (O_530,N_14798,N_14910);
and UO_531 (O_531,N_14770,N_14975);
nand UO_532 (O_532,N_14915,N_14861);
or UO_533 (O_533,N_14790,N_14802);
nand UO_534 (O_534,N_14772,N_14875);
nor UO_535 (O_535,N_14751,N_14821);
and UO_536 (O_536,N_14999,N_14741);
xnor UO_537 (O_537,N_14719,N_14842);
xor UO_538 (O_538,N_14774,N_14800);
nand UO_539 (O_539,N_14739,N_14841);
nor UO_540 (O_540,N_14865,N_14794);
nor UO_541 (O_541,N_14935,N_14854);
or UO_542 (O_542,N_14903,N_14915);
nand UO_543 (O_543,N_14882,N_14736);
xor UO_544 (O_544,N_14812,N_14833);
or UO_545 (O_545,N_14995,N_14801);
and UO_546 (O_546,N_14973,N_14795);
nor UO_547 (O_547,N_14906,N_14776);
or UO_548 (O_548,N_14956,N_14955);
xnor UO_549 (O_549,N_14939,N_14716);
nand UO_550 (O_550,N_14703,N_14735);
nor UO_551 (O_551,N_14881,N_14848);
xnor UO_552 (O_552,N_14861,N_14816);
xnor UO_553 (O_553,N_14808,N_14987);
xnor UO_554 (O_554,N_14802,N_14731);
nor UO_555 (O_555,N_14763,N_14700);
and UO_556 (O_556,N_14747,N_14843);
nand UO_557 (O_557,N_14787,N_14871);
xnor UO_558 (O_558,N_14954,N_14919);
nor UO_559 (O_559,N_14718,N_14798);
xor UO_560 (O_560,N_14737,N_14888);
nor UO_561 (O_561,N_14929,N_14756);
xor UO_562 (O_562,N_14974,N_14711);
and UO_563 (O_563,N_14829,N_14981);
nand UO_564 (O_564,N_14965,N_14925);
nor UO_565 (O_565,N_14767,N_14867);
nor UO_566 (O_566,N_14905,N_14863);
or UO_567 (O_567,N_14820,N_14984);
xor UO_568 (O_568,N_14881,N_14924);
nor UO_569 (O_569,N_14987,N_14855);
xnor UO_570 (O_570,N_14785,N_14828);
nor UO_571 (O_571,N_14926,N_14748);
nand UO_572 (O_572,N_14799,N_14874);
nor UO_573 (O_573,N_14974,N_14941);
nor UO_574 (O_574,N_14707,N_14716);
nand UO_575 (O_575,N_14723,N_14954);
nor UO_576 (O_576,N_14709,N_14783);
nand UO_577 (O_577,N_14765,N_14795);
or UO_578 (O_578,N_14853,N_14718);
and UO_579 (O_579,N_14800,N_14703);
nor UO_580 (O_580,N_14819,N_14802);
or UO_581 (O_581,N_14775,N_14767);
xnor UO_582 (O_582,N_14794,N_14753);
nor UO_583 (O_583,N_14782,N_14870);
nand UO_584 (O_584,N_14967,N_14957);
and UO_585 (O_585,N_14843,N_14738);
nor UO_586 (O_586,N_14739,N_14854);
xor UO_587 (O_587,N_14767,N_14740);
nor UO_588 (O_588,N_14719,N_14749);
or UO_589 (O_589,N_14800,N_14968);
or UO_590 (O_590,N_14815,N_14848);
and UO_591 (O_591,N_14836,N_14909);
and UO_592 (O_592,N_14965,N_14932);
nor UO_593 (O_593,N_14808,N_14851);
or UO_594 (O_594,N_14742,N_14868);
and UO_595 (O_595,N_14890,N_14785);
and UO_596 (O_596,N_14954,N_14945);
and UO_597 (O_597,N_14925,N_14720);
or UO_598 (O_598,N_14791,N_14780);
xor UO_599 (O_599,N_14797,N_14966);
xor UO_600 (O_600,N_14884,N_14899);
or UO_601 (O_601,N_14859,N_14845);
xor UO_602 (O_602,N_14716,N_14813);
and UO_603 (O_603,N_14744,N_14987);
nor UO_604 (O_604,N_14752,N_14816);
nor UO_605 (O_605,N_14889,N_14902);
or UO_606 (O_606,N_14823,N_14721);
xnor UO_607 (O_607,N_14938,N_14739);
and UO_608 (O_608,N_14844,N_14879);
nand UO_609 (O_609,N_14989,N_14919);
nor UO_610 (O_610,N_14934,N_14715);
xor UO_611 (O_611,N_14838,N_14886);
nand UO_612 (O_612,N_14791,N_14705);
nand UO_613 (O_613,N_14883,N_14957);
nand UO_614 (O_614,N_14726,N_14713);
and UO_615 (O_615,N_14744,N_14898);
nor UO_616 (O_616,N_14947,N_14895);
nand UO_617 (O_617,N_14959,N_14882);
nor UO_618 (O_618,N_14997,N_14881);
xnor UO_619 (O_619,N_14871,N_14731);
xor UO_620 (O_620,N_14946,N_14857);
nor UO_621 (O_621,N_14910,N_14930);
nor UO_622 (O_622,N_14979,N_14739);
nand UO_623 (O_623,N_14825,N_14973);
xnor UO_624 (O_624,N_14949,N_14916);
nand UO_625 (O_625,N_14877,N_14976);
xor UO_626 (O_626,N_14953,N_14863);
xnor UO_627 (O_627,N_14740,N_14969);
or UO_628 (O_628,N_14955,N_14845);
nand UO_629 (O_629,N_14788,N_14963);
nor UO_630 (O_630,N_14968,N_14802);
and UO_631 (O_631,N_14772,N_14762);
nor UO_632 (O_632,N_14922,N_14948);
xor UO_633 (O_633,N_14848,N_14700);
or UO_634 (O_634,N_14802,N_14906);
xnor UO_635 (O_635,N_14812,N_14958);
xor UO_636 (O_636,N_14907,N_14733);
xnor UO_637 (O_637,N_14943,N_14932);
nor UO_638 (O_638,N_14883,N_14838);
and UO_639 (O_639,N_14985,N_14700);
nand UO_640 (O_640,N_14983,N_14799);
nor UO_641 (O_641,N_14797,N_14950);
xnor UO_642 (O_642,N_14922,N_14828);
nor UO_643 (O_643,N_14975,N_14904);
nand UO_644 (O_644,N_14981,N_14893);
xor UO_645 (O_645,N_14740,N_14737);
or UO_646 (O_646,N_14943,N_14853);
and UO_647 (O_647,N_14895,N_14968);
nand UO_648 (O_648,N_14834,N_14953);
nand UO_649 (O_649,N_14744,N_14864);
nand UO_650 (O_650,N_14781,N_14785);
nor UO_651 (O_651,N_14940,N_14712);
nor UO_652 (O_652,N_14995,N_14896);
nor UO_653 (O_653,N_14823,N_14770);
nor UO_654 (O_654,N_14825,N_14782);
nand UO_655 (O_655,N_14806,N_14747);
or UO_656 (O_656,N_14852,N_14850);
and UO_657 (O_657,N_14811,N_14838);
and UO_658 (O_658,N_14803,N_14970);
nand UO_659 (O_659,N_14903,N_14900);
xor UO_660 (O_660,N_14771,N_14762);
nor UO_661 (O_661,N_14960,N_14718);
nand UO_662 (O_662,N_14703,N_14914);
nor UO_663 (O_663,N_14888,N_14881);
xnor UO_664 (O_664,N_14979,N_14807);
nand UO_665 (O_665,N_14956,N_14916);
and UO_666 (O_666,N_14877,N_14787);
xnor UO_667 (O_667,N_14739,N_14830);
or UO_668 (O_668,N_14754,N_14879);
xor UO_669 (O_669,N_14818,N_14815);
xnor UO_670 (O_670,N_14754,N_14791);
nor UO_671 (O_671,N_14938,N_14942);
nor UO_672 (O_672,N_14832,N_14717);
nor UO_673 (O_673,N_14885,N_14981);
nand UO_674 (O_674,N_14980,N_14715);
nor UO_675 (O_675,N_14731,N_14728);
nand UO_676 (O_676,N_14819,N_14861);
xor UO_677 (O_677,N_14759,N_14860);
nand UO_678 (O_678,N_14937,N_14732);
xor UO_679 (O_679,N_14730,N_14889);
or UO_680 (O_680,N_14803,N_14788);
nor UO_681 (O_681,N_14813,N_14993);
nor UO_682 (O_682,N_14876,N_14723);
and UO_683 (O_683,N_14800,N_14918);
and UO_684 (O_684,N_14799,N_14739);
nor UO_685 (O_685,N_14919,N_14942);
or UO_686 (O_686,N_14848,N_14917);
nand UO_687 (O_687,N_14792,N_14736);
and UO_688 (O_688,N_14963,N_14808);
nand UO_689 (O_689,N_14844,N_14775);
nand UO_690 (O_690,N_14701,N_14982);
or UO_691 (O_691,N_14751,N_14818);
nand UO_692 (O_692,N_14719,N_14993);
nor UO_693 (O_693,N_14744,N_14982);
and UO_694 (O_694,N_14839,N_14758);
and UO_695 (O_695,N_14807,N_14992);
and UO_696 (O_696,N_14898,N_14821);
xor UO_697 (O_697,N_14940,N_14938);
xor UO_698 (O_698,N_14934,N_14818);
and UO_699 (O_699,N_14799,N_14814);
xor UO_700 (O_700,N_14894,N_14831);
nor UO_701 (O_701,N_14978,N_14956);
nor UO_702 (O_702,N_14704,N_14887);
nor UO_703 (O_703,N_14861,N_14859);
nand UO_704 (O_704,N_14847,N_14989);
and UO_705 (O_705,N_14837,N_14771);
or UO_706 (O_706,N_14815,N_14719);
nand UO_707 (O_707,N_14708,N_14730);
xor UO_708 (O_708,N_14801,N_14760);
nor UO_709 (O_709,N_14992,N_14768);
nor UO_710 (O_710,N_14858,N_14772);
nor UO_711 (O_711,N_14812,N_14712);
xor UO_712 (O_712,N_14724,N_14853);
xnor UO_713 (O_713,N_14992,N_14818);
nor UO_714 (O_714,N_14986,N_14942);
or UO_715 (O_715,N_14792,N_14819);
or UO_716 (O_716,N_14872,N_14924);
or UO_717 (O_717,N_14926,N_14948);
and UO_718 (O_718,N_14892,N_14727);
nor UO_719 (O_719,N_14989,N_14773);
or UO_720 (O_720,N_14763,N_14871);
nand UO_721 (O_721,N_14745,N_14732);
nor UO_722 (O_722,N_14918,N_14717);
or UO_723 (O_723,N_14859,N_14904);
or UO_724 (O_724,N_14833,N_14957);
nor UO_725 (O_725,N_14921,N_14960);
nand UO_726 (O_726,N_14823,N_14828);
nand UO_727 (O_727,N_14961,N_14959);
and UO_728 (O_728,N_14987,N_14772);
nor UO_729 (O_729,N_14914,N_14785);
or UO_730 (O_730,N_14782,N_14986);
nand UO_731 (O_731,N_14793,N_14869);
and UO_732 (O_732,N_14973,N_14964);
and UO_733 (O_733,N_14744,N_14972);
and UO_734 (O_734,N_14977,N_14707);
or UO_735 (O_735,N_14760,N_14875);
or UO_736 (O_736,N_14774,N_14807);
nor UO_737 (O_737,N_14933,N_14716);
xor UO_738 (O_738,N_14807,N_14867);
and UO_739 (O_739,N_14851,N_14976);
nor UO_740 (O_740,N_14880,N_14900);
or UO_741 (O_741,N_14759,N_14795);
nor UO_742 (O_742,N_14883,N_14826);
or UO_743 (O_743,N_14916,N_14824);
xnor UO_744 (O_744,N_14881,N_14856);
nand UO_745 (O_745,N_14772,N_14712);
nor UO_746 (O_746,N_14740,N_14807);
nand UO_747 (O_747,N_14906,N_14772);
or UO_748 (O_748,N_14993,N_14842);
nand UO_749 (O_749,N_14976,N_14706);
and UO_750 (O_750,N_14939,N_14781);
or UO_751 (O_751,N_14922,N_14902);
nand UO_752 (O_752,N_14960,N_14802);
and UO_753 (O_753,N_14955,N_14788);
nor UO_754 (O_754,N_14768,N_14790);
xor UO_755 (O_755,N_14853,N_14918);
or UO_756 (O_756,N_14875,N_14832);
and UO_757 (O_757,N_14975,N_14756);
or UO_758 (O_758,N_14809,N_14789);
nor UO_759 (O_759,N_14712,N_14895);
nand UO_760 (O_760,N_14866,N_14734);
or UO_761 (O_761,N_14723,N_14867);
nand UO_762 (O_762,N_14902,N_14761);
nand UO_763 (O_763,N_14932,N_14837);
xnor UO_764 (O_764,N_14881,N_14793);
xor UO_765 (O_765,N_14824,N_14780);
and UO_766 (O_766,N_14911,N_14894);
and UO_767 (O_767,N_14745,N_14752);
nor UO_768 (O_768,N_14971,N_14727);
xor UO_769 (O_769,N_14978,N_14846);
nor UO_770 (O_770,N_14730,N_14914);
nor UO_771 (O_771,N_14883,N_14860);
and UO_772 (O_772,N_14828,N_14920);
nor UO_773 (O_773,N_14816,N_14724);
or UO_774 (O_774,N_14872,N_14819);
and UO_775 (O_775,N_14829,N_14782);
xor UO_776 (O_776,N_14999,N_14792);
nor UO_777 (O_777,N_14722,N_14896);
and UO_778 (O_778,N_14907,N_14901);
xor UO_779 (O_779,N_14915,N_14763);
or UO_780 (O_780,N_14842,N_14897);
nor UO_781 (O_781,N_14909,N_14933);
nor UO_782 (O_782,N_14960,N_14710);
nor UO_783 (O_783,N_14760,N_14798);
nand UO_784 (O_784,N_14945,N_14999);
nand UO_785 (O_785,N_14713,N_14826);
nor UO_786 (O_786,N_14741,N_14882);
and UO_787 (O_787,N_14931,N_14702);
xnor UO_788 (O_788,N_14782,N_14886);
or UO_789 (O_789,N_14704,N_14864);
xor UO_790 (O_790,N_14798,N_14756);
and UO_791 (O_791,N_14990,N_14727);
nand UO_792 (O_792,N_14975,N_14868);
nand UO_793 (O_793,N_14700,N_14806);
and UO_794 (O_794,N_14862,N_14785);
or UO_795 (O_795,N_14769,N_14947);
nor UO_796 (O_796,N_14932,N_14926);
nand UO_797 (O_797,N_14788,N_14838);
or UO_798 (O_798,N_14967,N_14968);
nor UO_799 (O_799,N_14954,N_14939);
xor UO_800 (O_800,N_14894,N_14782);
or UO_801 (O_801,N_14882,N_14878);
or UO_802 (O_802,N_14953,N_14789);
or UO_803 (O_803,N_14895,N_14978);
and UO_804 (O_804,N_14709,N_14863);
xnor UO_805 (O_805,N_14736,N_14916);
or UO_806 (O_806,N_14956,N_14782);
and UO_807 (O_807,N_14928,N_14721);
xnor UO_808 (O_808,N_14976,N_14715);
or UO_809 (O_809,N_14904,N_14748);
nor UO_810 (O_810,N_14721,N_14988);
xnor UO_811 (O_811,N_14702,N_14876);
nor UO_812 (O_812,N_14901,N_14707);
xor UO_813 (O_813,N_14875,N_14759);
nand UO_814 (O_814,N_14879,N_14740);
xor UO_815 (O_815,N_14817,N_14821);
nor UO_816 (O_816,N_14707,N_14866);
nor UO_817 (O_817,N_14997,N_14718);
nor UO_818 (O_818,N_14787,N_14718);
nor UO_819 (O_819,N_14863,N_14721);
or UO_820 (O_820,N_14950,N_14708);
xor UO_821 (O_821,N_14767,N_14790);
nor UO_822 (O_822,N_14871,N_14892);
xor UO_823 (O_823,N_14793,N_14866);
nor UO_824 (O_824,N_14987,N_14945);
nor UO_825 (O_825,N_14886,N_14799);
nand UO_826 (O_826,N_14767,N_14999);
nand UO_827 (O_827,N_14980,N_14767);
nor UO_828 (O_828,N_14749,N_14722);
nand UO_829 (O_829,N_14881,N_14959);
xnor UO_830 (O_830,N_14720,N_14815);
or UO_831 (O_831,N_14887,N_14955);
or UO_832 (O_832,N_14874,N_14763);
xor UO_833 (O_833,N_14746,N_14711);
nor UO_834 (O_834,N_14822,N_14772);
nor UO_835 (O_835,N_14839,N_14853);
nor UO_836 (O_836,N_14931,N_14879);
nor UO_837 (O_837,N_14836,N_14704);
nand UO_838 (O_838,N_14800,N_14847);
nand UO_839 (O_839,N_14943,N_14896);
xnor UO_840 (O_840,N_14865,N_14767);
or UO_841 (O_841,N_14841,N_14710);
xnor UO_842 (O_842,N_14773,N_14968);
nand UO_843 (O_843,N_14720,N_14730);
nand UO_844 (O_844,N_14967,N_14747);
xor UO_845 (O_845,N_14756,N_14946);
nand UO_846 (O_846,N_14775,N_14859);
nor UO_847 (O_847,N_14816,N_14887);
nand UO_848 (O_848,N_14853,N_14880);
and UO_849 (O_849,N_14993,N_14891);
xnor UO_850 (O_850,N_14710,N_14740);
and UO_851 (O_851,N_14872,N_14770);
or UO_852 (O_852,N_14938,N_14961);
nor UO_853 (O_853,N_14885,N_14839);
and UO_854 (O_854,N_14979,N_14901);
nor UO_855 (O_855,N_14729,N_14927);
or UO_856 (O_856,N_14888,N_14754);
nor UO_857 (O_857,N_14928,N_14901);
or UO_858 (O_858,N_14714,N_14925);
and UO_859 (O_859,N_14920,N_14924);
nor UO_860 (O_860,N_14867,N_14987);
xor UO_861 (O_861,N_14772,N_14803);
and UO_862 (O_862,N_14848,N_14913);
xor UO_863 (O_863,N_14924,N_14989);
or UO_864 (O_864,N_14989,N_14854);
or UO_865 (O_865,N_14878,N_14713);
and UO_866 (O_866,N_14937,N_14776);
or UO_867 (O_867,N_14920,N_14835);
nand UO_868 (O_868,N_14865,N_14932);
nand UO_869 (O_869,N_14979,N_14858);
nor UO_870 (O_870,N_14850,N_14943);
or UO_871 (O_871,N_14789,N_14806);
or UO_872 (O_872,N_14980,N_14876);
and UO_873 (O_873,N_14817,N_14897);
or UO_874 (O_874,N_14716,N_14856);
nor UO_875 (O_875,N_14737,N_14988);
xor UO_876 (O_876,N_14715,N_14922);
and UO_877 (O_877,N_14812,N_14782);
xnor UO_878 (O_878,N_14746,N_14808);
nor UO_879 (O_879,N_14884,N_14870);
xnor UO_880 (O_880,N_14990,N_14946);
and UO_881 (O_881,N_14997,N_14965);
nor UO_882 (O_882,N_14827,N_14811);
nor UO_883 (O_883,N_14792,N_14795);
or UO_884 (O_884,N_14797,N_14890);
xor UO_885 (O_885,N_14993,N_14732);
nor UO_886 (O_886,N_14731,N_14740);
xnor UO_887 (O_887,N_14898,N_14952);
and UO_888 (O_888,N_14927,N_14784);
nor UO_889 (O_889,N_14780,N_14832);
nor UO_890 (O_890,N_14966,N_14892);
nand UO_891 (O_891,N_14980,N_14959);
nor UO_892 (O_892,N_14846,N_14825);
nor UO_893 (O_893,N_14951,N_14713);
and UO_894 (O_894,N_14919,N_14793);
nor UO_895 (O_895,N_14745,N_14810);
and UO_896 (O_896,N_14884,N_14897);
or UO_897 (O_897,N_14754,N_14819);
and UO_898 (O_898,N_14766,N_14799);
nand UO_899 (O_899,N_14977,N_14802);
xnor UO_900 (O_900,N_14869,N_14969);
xnor UO_901 (O_901,N_14867,N_14942);
nand UO_902 (O_902,N_14979,N_14833);
and UO_903 (O_903,N_14866,N_14986);
and UO_904 (O_904,N_14902,N_14753);
and UO_905 (O_905,N_14776,N_14815);
xnor UO_906 (O_906,N_14972,N_14853);
or UO_907 (O_907,N_14837,N_14894);
or UO_908 (O_908,N_14932,N_14966);
xor UO_909 (O_909,N_14988,N_14743);
and UO_910 (O_910,N_14928,N_14703);
nor UO_911 (O_911,N_14741,N_14764);
and UO_912 (O_912,N_14951,N_14761);
xnor UO_913 (O_913,N_14832,N_14774);
xnor UO_914 (O_914,N_14752,N_14754);
or UO_915 (O_915,N_14766,N_14955);
and UO_916 (O_916,N_14900,N_14749);
nor UO_917 (O_917,N_14834,N_14734);
and UO_918 (O_918,N_14710,N_14947);
nand UO_919 (O_919,N_14904,N_14732);
nor UO_920 (O_920,N_14708,N_14897);
nor UO_921 (O_921,N_14917,N_14862);
or UO_922 (O_922,N_14843,N_14800);
xor UO_923 (O_923,N_14874,N_14864);
xor UO_924 (O_924,N_14978,N_14848);
xor UO_925 (O_925,N_14933,N_14935);
xnor UO_926 (O_926,N_14751,N_14731);
and UO_927 (O_927,N_14901,N_14899);
and UO_928 (O_928,N_14952,N_14891);
or UO_929 (O_929,N_14740,N_14988);
xnor UO_930 (O_930,N_14794,N_14858);
or UO_931 (O_931,N_14961,N_14772);
xor UO_932 (O_932,N_14801,N_14754);
and UO_933 (O_933,N_14931,N_14754);
nand UO_934 (O_934,N_14837,N_14920);
xor UO_935 (O_935,N_14833,N_14796);
and UO_936 (O_936,N_14833,N_14962);
or UO_937 (O_937,N_14737,N_14809);
and UO_938 (O_938,N_14816,N_14967);
or UO_939 (O_939,N_14780,N_14911);
and UO_940 (O_940,N_14887,N_14981);
and UO_941 (O_941,N_14702,N_14877);
xor UO_942 (O_942,N_14840,N_14701);
nor UO_943 (O_943,N_14800,N_14863);
xor UO_944 (O_944,N_14967,N_14761);
and UO_945 (O_945,N_14937,N_14816);
nand UO_946 (O_946,N_14877,N_14880);
and UO_947 (O_947,N_14897,N_14763);
or UO_948 (O_948,N_14757,N_14942);
nand UO_949 (O_949,N_14764,N_14726);
or UO_950 (O_950,N_14881,N_14704);
or UO_951 (O_951,N_14780,N_14808);
or UO_952 (O_952,N_14954,N_14702);
nor UO_953 (O_953,N_14783,N_14869);
nand UO_954 (O_954,N_14752,N_14895);
nand UO_955 (O_955,N_14905,N_14735);
xor UO_956 (O_956,N_14833,N_14757);
and UO_957 (O_957,N_14840,N_14843);
and UO_958 (O_958,N_14940,N_14831);
xor UO_959 (O_959,N_14762,N_14719);
or UO_960 (O_960,N_14796,N_14793);
or UO_961 (O_961,N_14894,N_14873);
and UO_962 (O_962,N_14942,N_14805);
nand UO_963 (O_963,N_14957,N_14778);
xor UO_964 (O_964,N_14783,N_14734);
xor UO_965 (O_965,N_14856,N_14762);
and UO_966 (O_966,N_14777,N_14954);
nor UO_967 (O_967,N_14832,N_14910);
nor UO_968 (O_968,N_14749,N_14725);
nor UO_969 (O_969,N_14700,N_14714);
or UO_970 (O_970,N_14981,N_14940);
nor UO_971 (O_971,N_14954,N_14904);
xor UO_972 (O_972,N_14821,N_14886);
xor UO_973 (O_973,N_14869,N_14720);
or UO_974 (O_974,N_14962,N_14753);
or UO_975 (O_975,N_14970,N_14955);
nand UO_976 (O_976,N_14872,N_14882);
nor UO_977 (O_977,N_14788,N_14978);
and UO_978 (O_978,N_14875,N_14748);
nor UO_979 (O_979,N_14795,N_14772);
and UO_980 (O_980,N_14995,N_14718);
or UO_981 (O_981,N_14847,N_14811);
xor UO_982 (O_982,N_14861,N_14840);
nand UO_983 (O_983,N_14862,N_14747);
and UO_984 (O_984,N_14817,N_14815);
xor UO_985 (O_985,N_14908,N_14967);
and UO_986 (O_986,N_14912,N_14801);
or UO_987 (O_987,N_14885,N_14975);
nor UO_988 (O_988,N_14896,N_14827);
nor UO_989 (O_989,N_14856,N_14889);
or UO_990 (O_990,N_14952,N_14994);
or UO_991 (O_991,N_14943,N_14902);
nor UO_992 (O_992,N_14952,N_14978);
nand UO_993 (O_993,N_14801,N_14887);
xnor UO_994 (O_994,N_14849,N_14853);
or UO_995 (O_995,N_14719,N_14922);
nor UO_996 (O_996,N_14784,N_14707);
xnor UO_997 (O_997,N_14889,N_14780);
or UO_998 (O_998,N_14767,N_14771);
xnor UO_999 (O_999,N_14925,N_14977);
and UO_1000 (O_1000,N_14973,N_14906);
or UO_1001 (O_1001,N_14914,N_14992);
or UO_1002 (O_1002,N_14866,N_14979);
xor UO_1003 (O_1003,N_14703,N_14806);
nand UO_1004 (O_1004,N_14982,N_14715);
and UO_1005 (O_1005,N_14764,N_14878);
nor UO_1006 (O_1006,N_14791,N_14808);
nand UO_1007 (O_1007,N_14741,N_14802);
nand UO_1008 (O_1008,N_14945,N_14725);
xnor UO_1009 (O_1009,N_14713,N_14778);
nand UO_1010 (O_1010,N_14815,N_14963);
nand UO_1011 (O_1011,N_14783,N_14787);
nor UO_1012 (O_1012,N_14821,N_14787);
and UO_1013 (O_1013,N_14907,N_14783);
xor UO_1014 (O_1014,N_14783,N_14922);
nor UO_1015 (O_1015,N_14905,N_14707);
xnor UO_1016 (O_1016,N_14768,N_14964);
xnor UO_1017 (O_1017,N_14765,N_14981);
nand UO_1018 (O_1018,N_14962,N_14888);
nand UO_1019 (O_1019,N_14869,N_14952);
nor UO_1020 (O_1020,N_14814,N_14779);
xor UO_1021 (O_1021,N_14857,N_14953);
nand UO_1022 (O_1022,N_14980,N_14780);
nor UO_1023 (O_1023,N_14879,N_14910);
nand UO_1024 (O_1024,N_14920,N_14905);
or UO_1025 (O_1025,N_14945,N_14704);
or UO_1026 (O_1026,N_14944,N_14960);
and UO_1027 (O_1027,N_14756,N_14830);
xnor UO_1028 (O_1028,N_14990,N_14705);
nand UO_1029 (O_1029,N_14977,N_14748);
xnor UO_1030 (O_1030,N_14946,N_14971);
and UO_1031 (O_1031,N_14745,N_14702);
nand UO_1032 (O_1032,N_14792,N_14740);
nand UO_1033 (O_1033,N_14976,N_14794);
nand UO_1034 (O_1034,N_14945,N_14774);
xor UO_1035 (O_1035,N_14872,N_14808);
nand UO_1036 (O_1036,N_14849,N_14992);
nand UO_1037 (O_1037,N_14800,N_14886);
xor UO_1038 (O_1038,N_14981,N_14870);
nor UO_1039 (O_1039,N_14917,N_14726);
nand UO_1040 (O_1040,N_14822,N_14944);
nor UO_1041 (O_1041,N_14987,N_14714);
xnor UO_1042 (O_1042,N_14715,N_14775);
or UO_1043 (O_1043,N_14873,N_14982);
xor UO_1044 (O_1044,N_14953,N_14785);
nor UO_1045 (O_1045,N_14927,N_14931);
nor UO_1046 (O_1046,N_14725,N_14835);
nand UO_1047 (O_1047,N_14783,N_14724);
and UO_1048 (O_1048,N_14975,N_14778);
nor UO_1049 (O_1049,N_14736,N_14988);
nand UO_1050 (O_1050,N_14907,N_14888);
nand UO_1051 (O_1051,N_14736,N_14996);
nor UO_1052 (O_1052,N_14953,N_14865);
nor UO_1053 (O_1053,N_14759,N_14995);
nand UO_1054 (O_1054,N_14783,N_14949);
or UO_1055 (O_1055,N_14750,N_14711);
nor UO_1056 (O_1056,N_14708,N_14853);
or UO_1057 (O_1057,N_14956,N_14792);
or UO_1058 (O_1058,N_14875,N_14915);
xnor UO_1059 (O_1059,N_14845,N_14983);
nand UO_1060 (O_1060,N_14946,N_14824);
or UO_1061 (O_1061,N_14961,N_14825);
nand UO_1062 (O_1062,N_14817,N_14729);
or UO_1063 (O_1063,N_14829,N_14886);
xnor UO_1064 (O_1064,N_14861,N_14880);
nand UO_1065 (O_1065,N_14811,N_14810);
and UO_1066 (O_1066,N_14931,N_14815);
nor UO_1067 (O_1067,N_14994,N_14872);
and UO_1068 (O_1068,N_14812,N_14747);
and UO_1069 (O_1069,N_14891,N_14940);
and UO_1070 (O_1070,N_14996,N_14779);
nand UO_1071 (O_1071,N_14971,N_14761);
nor UO_1072 (O_1072,N_14799,N_14839);
xor UO_1073 (O_1073,N_14860,N_14833);
xnor UO_1074 (O_1074,N_14930,N_14970);
nor UO_1075 (O_1075,N_14704,N_14920);
nand UO_1076 (O_1076,N_14879,N_14744);
nand UO_1077 (O_1077,N_14997,N_14763);
nand UO_1078 (O_1078,N_14906,N_14704);
nor UO_1079 (O_1079,N_14991,N_14768);
or UO_1080 (O_1080,N_14882,N_14731);
nor UO_1081 (O_1081,N_14757,N_14907);
xnor UO_1082 (O_1082,N_14754,N_14742);
and UO_1083 (O_1083,N_14935,N_14750);
nor UO_1084 (O_1084,N_14920,N_14857);
xor UO_1085 (O_1085,N_14791,N_14735);
and UO_1086 (O_1086,N_14936,N_14872);
nor UO_1087 (O_1087,N_14825,N_14873);
nor UO_1088 (O_1088,N_14843,N_14841);
xor UO_1089 (O_1089,N_14944,N_14888);
and UO_1090 (O_1090,N_14819,N_14830);
or UO_1091 (O_1091,N_14704,N_14852);
or UO_1092 (O_1092,N_14988,N_14809);
and UO_1093 (O_1093,N_14929,N_14890);
and UO_1094 (O_1094,N_14796,N_14960);
nor UO_1095 (O_1095,N_14964,N_14994);
nand UO_1096 (O_1096,N_14914,N_14836);
and UO_1097 (O_1097,N_14723,N_14974);
nand UO_1098 (O_1098,N_14972,N_14932);
nor UO_1099 (O_1099,N_14775,N_14759);
nor UO_1100 (O_1100,N_14926,N_14772);
xor UO_1101 (O_1101,N_14925,N_14872);
or UO_1102 (O_1102,N_14905,N_14981);
xor UO_1103 (O_1103,N_14981,N_14840);
nand UO_1104 (O_1104,N_14984,N_14712);
xnor UO_1105 (O_1105,N_14825,N_14736);
nor UO_1106 (O_1106,N_14902,N_14769);
or UO_1107 (O_1107,N_14813,N_14859);
or UO_1108 (O_1108,N_14876,N_14904);
and UO_1109 (O_1109,N_14890,N_14979);
xnor UO_1110 (O_1110,N_14873,N_14754);
or UO_1111 (O_1111,N_14902,N_14813);
and UO_1112 (O_1112,N_14771,N_14860);
xnor UO_1113 (O_1113,N_14744,N_14772);
nor UO_1114 (O_1114,N_14915,N_14964);
nand UO_1115 (O_1115,N_14855,N_14878);
nand UO_1116 (O_1116,N_14745,N_14701);
and UO_1117 (O_1117,N_14792,N_14830);
and UO_1118 (O_1118,N_14881,N_14721);
nor UO_1119 (O_1119,N_14983,N_14975);
and UO_1120 (O_1120,N_14972,N_14747);
and UO_1121 (O_1121,N_14872,N_14835);
or UO_1122 (O_1122,N_14816,N_14933);
xor UO_1123 (O_1123,N_14729,N_14761);
and UO_1124 (O_1124,N_14900,N_14901);
or UO_1125 (O_1125,N_14711,N_14892);
nand UO_1126 (O_1126,N_14989,N_14828);
nand UO_1127 (O_1127,N_14940,N_14925);
and UO_1128 (O_1128,N_14855,N_14956);
nor UO_1129 (O_1129,N_14732,N_14962);
xnor UO_1130 (O_1130,N_14728,N_14980);
xor UO_1131 (O_1131,N_14947,N_14915);
and UO_1132 (O_1132,N_14949,N_14984);
nand UO_1133 (O_1133,N_14702,N_14871);
and UO_1134 (O_1134,N_14709,N_14837);
nor UO_1135 (O_1135,N_14726,N_14727);
or UO_1136 (O_1136,N_14913,N_14755);
nor UO_1137 (O_1137,N_14889,N_14762);
or UO_1138 (O_1138,N_14839,N_14745);
and UO_1139 (O_1139,N_14955,N_14995);
and UO_1140 (O_1140,N_14950,N_14826);
and UO_1141 (O_1141,N_14797,N_14767);
or UO_1142 (O_1142,N_14786,N_14832);
and UO_1143 (O_1143,N_14865,N_14778);
and UO_1144 (O_1144,N_14769,N_14925);
and UO_1145 (O_1145,N_14974,N_14938);
xor UO_1146 (O_1146,N_14844,N_14983);
and UO_1147 (O_1147,N_14785,N_14942);
and UO_1148 (O_1148,N_14844,N_14785);
or UO_1149 (O_1149,N_14818,N_14771);
and UO_1150 (O_1150,N_14804,N_14967);
nor UO_1151 (O_1151,N_14750,N_14819);
xnor UO_1152 (O_1152,N_14793,N_14781);
or UO_1153 (O_1153,N_14771,N_14774);
and UO_1154 (O_1154,N_14797,N_14735);
or UO_1155 (O_1155,N_14856,N_14938);
or UO_1156 (O_1156,N_14738,N_14724);
or UO_1157 (O_1157,N_14811,N_14988);
nand UO_1158 (O_1158,N_14968,N_14716);
and UO_1159 (O_1159,N_14735,N_14969);
nand UO_1160 (O_1160,N_14737,N_14755);
and UO_1161 (O_1161,N_14929,N_14786);
nand UO_1162 (O_1162,N_14914,N_14896);
or UO_1163 (O_1163,N_14889,N_14969);
or UO_1164 (O_1164,N_14774,N_14853);
and UO_1165 (O_1165,N_14748,N_14874);
and UO_1166 (O_1166,N_14799,N_14767);
or UO_1167 (O_1167,N_14886,N_14852);
or UO_1168 (O_1168,N_14819,N_14864);
xnor UO_1169 (O_1169,N_14730,N_14944);
or UO_1170 (O_1170,N_14988,N_14875);
and UO_1171 (O_1171,N_14794,N_14977);
or UO_1172 (O_1172,N_14879,N_14898);
or UO_1173 (O_1173,N_14942,N_14999);
or UO_1174 (O_1174,N_14825,N_14844);
xnor UO_1175 (O_1175,N_14944,N_14748);
or UO_1176 (O_1176,N_14747,N_14816);
nor UO_1177 (O_1177,N_14914,N_14899);
xor UO_1178 (O_1178,N_14816,N_14913);
nand UO_1179 (O_1179,N_14982,N_14894);
and UO_1180 (O_1180,N_14851,N_14750);
or UO_1181 (O_1181,N_14767,N_14753);
nand UO_1182 (O_1182,N_14900,N_14803);
or UO_1183 (O_1183,N_14912,N_14986);
nor UO_1184 (O_1184,N_14720,N_14973);
nor UO_1185 (O_1185,N_14984,N_14827);
and UO_1186 (O_1186,N_14773,N_14784);
nand UO_1187 (O_1187,N_14797,N_14763);
xnor UO_1188 (O_1188,N_14923,N_14738);
nor UO_1189 (O_1189,N_14981,N_14777);
and UO_1190 (O_1190,N_14718,N_14868);
and UO_1191 (O_1191,N_14944,N_14851);
nor UO_1192 (O_1192,N_14901,N_14896);
nor UO_1193 (O_1193,N_14925,N_14756);
or UO_1194 (O_1194,N_14983,N_14810);
nand UO_1195 (O_1195,N_14999,N_14843);
and UO_1196 (O_1196,N_14968,N_14820);
xnor UO_1197 (O_1197,N_14791,N_14777);
nand UO_1198 (O_1198,N_14943,N_14926);
and UO_1199 (O_1199,N_14898,N_14977);
or UO_1200 (O_1200,N_14995,N_14833);
nand UO_1201 (O_1201,N_14771,N_14775);
xor UO_1202 (O_1202,N_14949,N_14938);
nor UO_1203 (O_1203,N_14754,N_14965);
nand UO_1204 (O_1204,N_14993,N_14703);
nand UO_1205 (O_1205,N_14919,N_14719);
xor UO_1206 (O_1206,N_14829,N_14806);
xnor UO_1207 (O_1207,N_14818,N_14983);
xor UO_1208 (O_1208,N_14983,N_14715);
nand UO_1209 (O_1209,N_14893,N_14785);
or UO_1210 (O_1210,N_14836,N_14932);
xnor UO_1211 (O_1211,N_14829,N_14916);
nor UO_1212 (O_1212,N_14921,N_14955);
or UO_1213 (O_1213,N_14857,N_14935);
and UO_1214 (O_1214,N_14724,N_14992);
or UO_1215 (O_1215,N_14910,N_14963);
and UO_1216 (O_1216,N_14934,N_14748);
nor UO_1217 (O_1217,N_14975,N_14727);
xnor UO_1218 (O_1218,N_14886,N_14956);
and UO_1219 (O_1219,N_14812,N_14790);
and UO_1220 (O_1220,N_14764,N_14783);
xnor UO_1221 (O_1221,N_14724,N_14732);
nand UO_1222 (O_1222,N_14819,N_14842);
and UO_1223 (O_1223,N_14715,N_14741);
and UO_1224 (O_1224,N_14863,N_14816);
and UO_1225 (O_1225,N_14880,N_14731);
nor UO_1226 (O_1226,N_14986,N_14981);
nor UO_1227 (O_1227,N_14897,N_14971);
nor UO_1228 (O_1228,N_14914,N_14772);
and UO_1229 (O_1229,N_14987,N_14838);
xnor UO_1230 (O_1230,N_14813,N_14847);
nand UO_1231 (O_1231,N_14930,N_14963);
xnor UO_1232 (O_1232,N_14765,N_14735);
or UO_1233 (O_1233,N_14754,N_14794);
nor UO_1234 (O_1234,N_14964,N_14764);
xnor UO_1235 (O_1235,N_14880,N_14967);
xnor UO_1236 (O_1236,N_14936,N_14834);
nand UO_1237 (O_1237,N_14801,N_14945);
nand UO_1238 (O_1238,N_14831,N_14986);
and UO_1239 (O_1239,N_14975,N_14906);
and UO_1240 (O_1240,N_14838,N_14704);
or UO_1241 (O_1241,N_14867,N_14764);
and UO_1242 (O_1242,N_14754,N_14833);
or UO_1243 (O_1243,N_14782,N_14765);
or UO_1244 (O_1244,N_14882,N_14907);
or UO_1245 (O_1245,N_14911,N_14801);
and UO_1246 (O_1246,N_14738,N_14834);
xor UO_1247 (O_1247,N_14781,N_14985);
and UO_1248 (O_1248,N_14864,N_14761);
or UO_1249 (O_1249,N_14707,N_14984);
or UO_1250 (O_1250,N_14716,N_14760);
nor UO_1251 (O_1251,N_14961,N_14929);
nand UO_1252 (O_1252,N_14972,N_14769);
or UO_1253 (O_1253,N_14781,N_14849);
nor UO_1254 (O_1254,N_14939,N_14805);
or UO_1255 (O_1255,N_14942,N_14853);
or UO_1256 (O_1256,N_14831,N_14702);
nand UO_1257 (O_1257,N_14910,N_14891);
or UO_1258 (O_1258,N_14999,N_14929);
nor UO_1259 (O_1259,N_14745,N_14990);
nor UO_1260 (O_1260,N_14886,N_14993);
nand UO_1261 (O_1261,N_14969,N_14895);
nand UO_1262 (O_1262,N_14971,N_14832);
xor UO_1263 (O_1263,N_14921,N_14867);
and UO_1264 (O_1264,N_14706,N_14777);
or UO_1265 (O_1265,N_14764,N_14713);
xnor UO_1266 (O_1266,N_14935,N_14812);
nor UO_1267 (O_1267,N_14816,N_14728);
nor UO_1268 (O_1268,N_14838,N_14834);
xor UO_1269 (O_1269,N_14729,N_14967);
xor UO_1270 (O_1270,N_14721,N_14931);
nor UO_1271 (O_1271,N_14932,N_14984);
or UO_1272 (O_1272,N_14732,N_14780);
xnor UO_1273 (O_1273,N_14737,N_14712);
and UO_1274 (O_1274,N_14725,N_14731);
nand UO_1275 (O_1275,N_14724,N_14763);
nand UO_1276 (O_1276,N_14921,N_14861);
nand UO_1277 (O_1277,N_14756,N_14742);
and UO_1278 (O_1278,N_14917,N_14999);
nand UO_1279 (O_1279,N_14874,N_14980);
nor UO_1280 (O_1280,N_14902,N_14780);
or UO_1281 (O_1281,N_14729,N_14930);
nor UO_1282 (O_1282,N_14786,N_14748);
nand UO_1283 (O_1283,N_14810,N_14975);
nand UO_1284 (O_1284,N_14769,N_14747);
nor UO_1285 (O_1285,N_14819,N_14886);
xnor UO_1286 (O_1286,N_14707,N_14942);
or UO_1287 (O_1287,N_14890,N_14908);
xor UO_1288 (O_1288,N_14727,N_14766);
and UO_1289 (O_1289,N_14838,N_14763);
nand UO_1290 (O_1290,N_14737,N_14919);
xor UO_1291 (O_1291,N_14851,N_14735);
nand UO_1292 (O_1292,N_14919,N_14863);
nor UO_1293 (O_1293,N_14920,N_14998);
nand UO_1294 (O_1294,N_14922,N_14812);
nand UO_1295 (O_1295,N_14982,N_14903);
nand UO_1296 (O_1296,N_14930,N_14810);
nor UO_1297 (O_1297,N_14899,N_14925);
nor UO_1298 (O_1298,N_14856,N_14876);
or UO_1299 (O_1299,N_14951,N_14769);
nor UO_1300 (O_1300,N_14903,N_14955);
or UO_1301 (O_1301,N_14703,N_14712);
and UO_1302 (O_1302,N_14966,N_14974);
or UO_1303 (O_1303,N_14995,N_14900);
nand UO_1304 (O_1304,N_14990,N_14749);
or UO_1305 (O_1305,N_14883,N_14785);
nor UO_1306 (O_1306,N_14707,N_14963);
nand UO_1307 (O_1307,N_14992,N_14721);
nand UO_1308 (O_1308,N_14904,N_14882);
nand UO_1309 (O_1309,N_14961,N_14985);
xor UO_1310 (O_1310,N_14782,N_14999);
nand UO_1311 (O_1311,N_14776,N_14729);
nor UO_1312 (O_1312,N_14883,N_14808);
and UO_1313 (O_1313,N_14735,N_14815);
nor UO_1314 (O_1314,N_14839,N_14944);
or UO_1315 (O_1315,N_14712,N_14866);
nor UO_1316 (O_1316,N_14948,N_14786);
nand UO_1317 (O_1317,N_14943,N_14835);
xor UO_1318 (O_1318,N_14983,N_14837);
xor UO_1319 (O_1319,N_14939,N_14908);
or UO_1320 (O_1320,N_14753,N_14805);
xnor UO_1321 (O_1321,N_14706,N_14912);
xor UO_1322 (O_1322,N_14961,N_14839);
nor UO_1323 (O_1323,N_14741,N_14997);
nor UO_1324 (O_1324,N_14783,N_14861);
xor UO_1325 (O_1325,N_14810,N_14734);
nor UO_1326 (O_1326,N_14834,N_14985);
and UO_1327 (O_1327,N_14805,N_14754);
xnor UO_1328 (O_1328,N_14836,N_14899);
xnor UO_1329 (O_1329,N_14832,N_14925);
nor UO_1330 (O_1330,N_14754,N_14995);
nand UO_1331 (O_1331,N_14846,N_14873);
and UO_1332 (O_1332,N_14787,N_14794);
nand UO_1333 (O_1333,N_14705,N_14818);
xor UO_1334 (O_1334,N_14702,N_14874);
xnor UO_1335 (O_1335,N_14837,N_14976);
xor UO_1336 (O_1336,N_14929,N_14996);
nor UO_1337 (O_1337,N_14922,N_14966);
nor UO_1338 (O_1338,N_14821,N_14921);
or UO_1339 (O_1339,N_14906,N_14741);
and UO_1340 (O_1340,N_14947,N_14949);
xor UO_1341 (O_1341,N_14826,N_14781);
xnor UO_1342 (O_1342,N_14740,N_14837);
nor UO_1343 (O_1343,N_14731,N_14859);
xor UO_1344 (O_1344,N_14873,N_14958);
or UO_1345 (O_1345,N_14879,N_14796);
or UO_1346 (O_1346,N_14924,N_14832);
nand UO_1347 (O_1347,N_14994,N_14734);
or UO_1348 (O_1348,N_14931,N_14742);
nor UO_1349 (O_1349,N_14777,N_14863);
nand UO_1350 (O_1350,N_14884,N_14864);
and UO_1351 (O_1351,N_14888,N_14719);
nor UO_1352 (O_1352,N_14717,N_14901);
and UO_1353 (O_1353,N_14982,N_14935);
nand UO_1354 (O_1354,N_14937,N_14965);
xor UO_1355 (O_1355,N_14737,N_14746);
and UO_1356 (O_1356,N_14980,N_14787);
or UO_1357 (O_1357,N_14785,N_14700);
or UO_1358 (O_1358,N_14957,N_14852);
or UO_1359 (O_1359,N_14901,N_14933);
or UO_1360 (O_1360,N_14754,N_14964);
nand UO_1361 (O_1361,N_14766,N_14837);
xor UO_1362 (O_1362,N_14950,N_14897);
nand UO_1363 (O_1363,N_14996,N_14986);
and UO_1364 (O_1364,N_14826,N_14844);
xnor UO_1365 (O_1365,N_14841,N_14823);
or UO_1366 (O_1366,N_14760,N_14804);
nor UO_1367 (O_1367,N_14785,N_14808);
or UO_1368 (O_1368,N_14828,N_14882);
and UO_1369 (O_1369,N_14835,N_14854);
xor UO_1370 (O_1370,N_14749,N_14791);
xnor UO_1371 (O_1371,N_14858,N_14768);
and UO_1372 (O_1372,N_14970,N_14876);
and UO_1373 (O_1373,N_14786,N_14926);
nand UO_1374 (O_1374,N_14899,N_14713);
and UO_1375 (O_1375,N_14828,N_14826);
and UO_1376 (O_1376,N_14937,N_14948);
nor UO_1377 (O_1377,N_14784,N_14788);
and UO_1378 (O_1378,N_14803,N_14895);
or UO_1379 (O_1379,N_14830,N_14738);
or UO_1380 (O_1380,N_14825,N_14900);
nand UO_1381 (O_1381,N_14857,N_14883);
or UO_1382 (O_1382,N_14965,N_14954);
nand UO_1383 (O_1383,N_14709,N_14933);
and UO_1384 (O_1384,N_14977,N_14994);
nor UO_1385 (O_1385,N_14922,N_14850);
xor UO_1386 (O_1386,N_14938,N_14803);
xnor UO_1387 (O_1387,N_14899,N_14875);
nor UO_1388 (O_1388,N_14709,N_14854);
or UO_1389 (O_1389,N_14782,N_14929);
nor UO_1390 (O_1390,N_14824,N_14762);
or UO_1391 (O_1391,N_14980,N_14955);
xor UO_1392 (O_1392,N_14791,N_14903);
nand UO_1393 (O_1393,N_14921,N_14997);
nand UO_1394 (O_1394,N_14845,N_14915);
xnor UO_1395 (O_1395,N_14734,N_14818);
nand UO_1396 (O_1396,N_14808,N_14752);
nor UO_1397 (O_1397,N_14934,N_14842);
or UO_1398 (O_1398,N_14971,N_14938);
and UO_1399 (O_1399,N_14881,N_14948);
and UO_1400 (O_1400,N_14811,N_14750);
and UO_1401 (O_1401,N_14706,N_14701);
and UO_1402 (O_1402,N_14952,N_14903);
and UO_1403 (O_1403,N_14887,N_14939);
nand UO_1404 (O_1404,N_14851,N_14998);
xnor UO_1405 (O_1405,N_14990,N_14719);
nand UO_1406 (O_1406,N_14808,N_14948);
nor UO_1407 (O_1407,N_14732,N_14842);
or UO_1408 (O_1408,N_14744,N_14938);
or UO_1409 (O_1409,N_14965,N_14818);
or UO_1410 (O_1410,N_14858,N_14785);
xor UO_1411 (O_1411,N_14864,N_14875);
xnor UO_1412 (O_1412,N_14759,N_14888);
nor UO_1413 (O_1413,N_14856,N_14840);
or UO_1414 (O_1414,N_14886,N_14830);
xor UO_1415 (O_1415,N_14802,N_14915);
and UO_1416 (O_1416,N_14751,N_14764);
or UO_1417 (O_1417,N_14856,N_14917);
nor UO_1418 (O_1418,N_14847,N_14826);
and UO_1419 (O_1419,N_14893,N_14911);
xor UO_1420 (O_1420,N_14994,N_14887);
or UO_1421 (O_1421,N_14996,N_14982);
xor UO_1422 (O_1422,N_14793,N_14911);
nand UO_1423 (O_1423,N_14725,N_14822);
and UO_1424 (O_1424,N_14773,N_14752);
xnor UO_1425 (O_1425,N_14902,N_14701);
and UO_1426 (O_1426,N_14724,N_14962);
xnor UO_1427 (O_1427,N_14739,N_14750);
and UO_1428 (O_1428,N_14753,N_14998);
xor UO_1429 (O_1429,N_14863,N_14793);
nand UO_1430 (O_1430,N_14777,N_14715);
nand UO_1431 (O_1431,N_14912,N_14872);
nand UO_1432 (O_1432,N_14961,N_14897);
nand UO_1433 (O_1433,N_14923,N_14981);
nor UO_1434 (O_1434,N_14926,N_14702);
and UO_1435 (O_1435,N_14937,N_14985);
and UO_1436 (O_1436,N_14966,N_14857);
xnor UO_1437 (O_1437,N_14898,N_14811);
nor UO_1438 (O_1438,N_14877,N_14747);
and UO_1439 (O_1439,N_14999,N_14886);
xor UO_1440 (O_1440,N_14814,N_14798);
nand UO_1441 (O_1441,N_14749,N_14777);
nor UO_1442 (O_1442,N_14926,N_14904);
nand UO_1443 (O_1443,N_14707,N_14753);
nor UO_1444 (O_1444,N_14842,N_14977);
or UO_1445 (O_1445,N_14819,N_14763);
or UO_1446 (O_1446,N_14771,N_14876);
or UO_1447 (O_1447,N_14779,N_14893);
xnor UO_1448 (O_1448,N_14893,N_14832);
or UO_1449 (O_1449,N_14968,N_14852);
nor UO_1450 (O_1450,N_14700,N_14962);
and UO_1451 (O_1451,N_14987,N_14900);
nor UO_1452 (O_1452,N_14927,N_14923);
or UO_1453 (O_1453,N_14777,N_14922);
and UO_1454 (O_1454,N_14873,N_14780);
nand UO_1455 (O_1455,N_14817,N_14981);
nor UO_1456 (O_1456,N_14744,N_14845);
and UO_1457 (O_1457,N_14809,N_14869);
nand UO_1458 (O_1458,N_14917,N_14769);
nand UO_1459 (O_1459,N_14972,N_14745);
nor UO_1460 (O_1460,N_14713,N_14870);
or UO_1461 (O_1461,N_14771,N_14786);
or UO_1462 (O_1462,N_14762,N_14916);
nor UO_1463 (O_1463,N_14783,N_14811);
or UO_1464 (O_1464,N_14984,N_14920);
xor UO_1465 (O_1465,N_14742,N_14734);
xor UO_1466 (O_1466,N_14917,N_14704);
and UO_1467 (O_1467,N_14751,N_14928);
nand UO_1468 (O_1468,N_14767,N_14735);
nand UO_1469 (O_1469,N_14919,N_14996);
or UO_1470 (O_1470,N_14966,N_14752);
nand UO_1471 (O_1471,N_14724,N_14984);
and UO_1472 (O_1472,N_14967,N_14948);
nand UO_1473 (O_1473,N_14944,N_14793);
xnor UO_1474 (O_1474,N_14834,N_14809);
and UO_1475 (O_1475,N_14937,N_14857);
and UO_1476 (O_1476,N_14780,N_14939);
xor UO_1477 (O_1477,N_14850,N_14830);
and UO_1478 (O_1478,N_14949,N_14835);
and UO_1479 (O_1479,N_14885,N_14716);
and UO_1480 (O_1480,N_14783,N_14969);
or UO_1481 (O_1481,N_14916,N_14752);
and UO_1482 (O_1482,N_14841,N_14859);
nand UO_1483 (O_1483,N_14814,N_14998);
nor UO_1484 (O_1484,N_14811,N_14891);
nor UO_1485 (O_1485,N_14705,N_14756);
nand UO_1486 (O_1486,N_14905,N_14829);
or UO_1487 (O_1487,N_14759,N_14820);
nor UO_1488 (O_1488,N_14858,N_14861);
nor UO_1489 (O_1489,N_14799,N_14998);
nand UO_1490 (O_1490,N_14734,N_14931);
and UO_1491 (O_1491,N_14703,N_14777);
nand UO_1492 (O_1492,N_14748,N_14828);
nor UO_1493 (O_1493,N_14737,N_14921);
xor UO_1494 (O_1494,N_14876,N_14767);
or UO_1495 (O_1495,N_14795,N_14713);
or UO_1496 (O_1496,N_14849,N_14703);
and UO_1497 (O_1497,N_14945,N_14920);
nand UO_1498 (O_1498,N_14702,N_14819);
or UO_1499 (O_1499,N_14774,N_14745);
xnor UO_1500 (O_1500,N_14856,N_14833);
or UO_1501 (O_1501,N_14858,N_14899);
nand UO_1502 (O_1502,N_14793,N_14808);
and UO_1503 (O_1503,N_14721,N_14930);
nand UO_1504 (O_1504,N_14705,N_14715);
nor UO_1505 (O_1505,N_14744,N_14788);
xnor UO_1506 (O_1506,N_14885,N_14829);
and UO_1507 (O_1507,N_14724,N_14894);
nor UO_1508 (O_1508,N_14910,N_14950);
nor UO_1509 (O_1509,N_14831,N_14936);
or UO_1510 (O_1510,N_14841,N_14777);
nor UO_1511 (O_1511,N_14827,N_14707);
nand UO_1512 (O_1512,N_14892,N_14717);
nand UO_1513 (O_1513,N_14882,N_14798);
nand UO_1514 (O_1514,N_14920,N_14971);
nor UO_1515 (O_1515,N_14978,N_14799);
xor UO_1516 (O_1516,N_14714,N_14782);
nor UO_1517 (O_1517,N_14704,N_14840);
and UO_1518 (O_1518,N_14742,N_14977);
nand UO_1519 (O_1519,N_14959,N_14723);
and UO_1520 (O_1520,N_14897,N_14891);
nor UO_1521 (O_1521,N_14904,N_14938);
nor UO_1522 (O_1522,N_14762,N_14898);
nand UO_1523 (O_1523,N_14988,N_14869);
xnor UO_1524 (O_1524,N_14799,N_14885);
and UO_1525 (O_1525,N_14881,N_14985);
xor UO_1526 (O_1526,N_14885,N_14925);
xor UO_1527 (O_1527,N_14992,N_14763);
xor UO_1528 (O_1528,N_14774,N_14760);
nand UO_1529 (O_1529,N_14948,N_14746);
and UO_1530 (O_1530,N_14957,N_14802);
and UO_1531 (O_1531,N_14844,N_14981);
xor UO_1532 (O_1532,N_14872,N_14714);
xor UO_1533 (O_1533,N_14993,N_14875);
or UO_1534 (O_1534,N_14779,N_14783);
and UO_1535 (O_1535,N_14866,N_14869);
xnor UO_1536 (O_1536,N_14987,N_14871);
or UO_1537 (O_1537,N_14730,N_14812);
and UO_1538 (O_1538,N_14728,N_14755);
nor UO_1539 (O_1539,N_14814,N_14909);
xnor UO_1540 (O_1540,N_14826,N_14843);
and UO_1541 (O_1541,N_14763,N_14824);
or UO_1542 (O_1542,N_14792,N_14908);
nor UO_1543 (O_1543,N_14999,N_14738);
and UO_1544 (O_1544,N_14777,N_14892);
nor UO_1545 (O_1545,N_14766,N_14827);
nor UO_1546 (O_1546,N_14727,N_14910);
xor UO_1547 (O_1547,N_14760,N_14983);
or UO_1548 (O_1548,N_14829,N_14892);
nand UO_1549 (O_1549,N_14887,N_14744);
xor UO_1550 (O_1550,N_14995,N_14923);
and UO_1551 (O_1551,N_14754,N_14734);
and UO_1552 (O_1552,N_14963,N_14891);
nor UO_1553 (O_1553,N_14924,N_14860);
nor UO_1554 (O_1554,N_14867,N_14820);
nor UO_1555 (O_1555,N_14841,N_14704);
nor UO_1556 (O_1556,N_14995,N_14866);
nand UO_1557 (O_1557,N_14906,N_14855);
nor UO_1558 (O_1558,N_14741,N_14784);
xnor UO_1559 (O_1559,N_14909,N_14991);
nor UO_1560 (O_1560,N_14974,N_14759);
or UO_1561 (O_1561,N_14736,N_14857);
or UO_1562 (O_1562,N_14703,N_14793);
or UO_1563 (O_1563,N_14918,N_14748);
and UO_1564 (O_1564,N_14763,N_14991);
nand UO_1565 (O_1565,N_14848,N_14814);
and UO_1566 (O_1566,N_14889,N_14753);
xnor UO_1567 (O_1567,N_14849,N_14821);
xnor UO_1568 (O_1568,N_14846,N_14864);
nor UO_1569 (O_1569,N_14740,N_14749);
or UO_1570 (O_1570,N_14923,N_14860);
or UO_1571 (O_1571,N_14986,N_14949);
xor UO_1572 (O_1572,N_14888,N_14927);
or UO_1573 (O_1573,N_14740,N_14893);
or UO_1574 (O_1574,N_14754,N_14823);
xnor UO_1575 (O_1575,N_14992,N_14738);
nor UO_1576 (O_1576,N_14808,N_14926);
xor UO_1577 (O_1577,N_14977,N_14827);
xnor UO_1578 (O_1578,N_14788,N_14738);
or UO_1579 (O_1579,N_14944,N_14940);
or UO_1580 (O_1580,N_14986,N_14740);
nor UO_1581 (O_1581,N_14763,N_14813);
nand UO_1582 (O_1582,N_14970,N_14784);
and UO_1583 (O_1583,N_14932,N_14935);
or UO_1584 (O_1584,N_14822,N_14861);
nand UO_1585 (O_1585,N_14726,N_14725);
or UO_1586 (O_1586,N_14845,N_14793);
nand UO_1587 (O_1587,N_14968,N_14944);
xnor UO_1588 (O_1588,N_14814,N_14928);
nand UO_1589 (O_1589,N_14880,N_14891);
nor UO_1590 (O_1590,N_14975,N_14842);
nand UO_1591 (O_1591,N_14808,N_14972);
nand UO_1592 (O_1592,N_14714,N_14994);
or UO_1593 (O_1593,N_14951,N_14890);
or UO_1594 (O_1594,N_14913,N_14834);
and UO_1595 (O_1595,N_14861,N_14871);
nor UO_1596 (O_1596,N_14941,N_14870);
xor UO_1597 (O_1597,N_14892,N_14895);
or UO_1598 (O_1598,N_14789,N_14765);
xor UO_1599 (O_1599,N_14782,N_14732);
or UO_1600 (O_1600,N_14742,N_14772);
or UO_1601 (O_1601,N_14990,N_14802);
xnor UO_1602 (O_1602,N_14877,N_14808);
and UO_1603 (O_1603,N_14944,N_14769);
and UO_1604 (O_1604,N_14740,N_14863);
nor UO_1605 (O_1605,N_14790,N_14872);
nor UO_1606 (O_1606,N_14743,N_14869);
xnor UO_1607 (O_1607,N_14829,N_14861);
and UO_1608 (O_1608,N_14742,N_14829);
nand UO_1609 (O_1609,N_14979,N_14811);
or UO_1610 (O_1610,N_14979,N_14931);
or UO_1611 (O_1611,N_14990,N_14959);
nand UO_1612 (O_1612,N_14854,N_14759);
and UO_1613 (O_1613,N_14961,N_14810);
nand UO_1614 (O_1614,N_14825,N_14910);
xor UO_1615 (O_1615,N_14946,N_14987);
nand UO_1616 (O_1616,N_14860,N_14876);
or UO_1617 (O_1617,N_14963,N_14980);
nand UO_1618 (O_1618,N_14828,N_14799);
and UO_1619 (O_1619,N_14866,N_14725);
nand UO_1620 (O_1620,N_14711,N_14931);
nand UO_1621 (O_1621,N_14948,N_14777);
and UO_1622 (O_1622,N_14904,N_14958);
nor UO_1623 (O_1623,N_14958,N_14798);
nand UO_1624 (O_1624,N_14894,N_14725);
xor UO_1625 (O_1625,N_14984,N_14860);
nor UO_1626 (O_1626,N_14847,N_14839);
and UO_1627 (O_1627,N_14926,N_14938);
nor UO_1628 (O_1628,N_14909,N_14784);
or UO_1629 (O_1629,N_14880,N_14941);
xor UO_1630 (O_1630,N_14933,N_14905);
nand UO_1631 (O_1631,N_14919,N_14855);
nand UO_1632 (O_1632,N_14740,N_14982);
xor UO_1633 (O_1633,N_14989,N_14955);
nand UO_1634 (O_1634,N_14732,N_14945);
xnor UO_1635 (O_1635,N_14927,N_14974);
nor UO_1636 (O_1636,N_14787,N_14789);
or UO_1637 (O_1637,N_14925,N_14921);
xnor UO_1638 (O_1638,N_14877,N_14751);
xnor UO_1639 (O_1639,N_14945,N_14867);
nor UO_1640 (O_1640,N_14714,N_14736);
xnor UO_1641 (O_1641,N_14950,N_14750);
xnor UO_1642 (O_1642,N_14986,N_14733);
nand UO_1643 (O_1643,N_14931,N_14908);
and UO_1644 (O_1644,N_14982,N_14844);
xor UO_1645 (O_1645,N_14847,N_14770);
xor UO_1646 (O_1646,N_14949,N_14746);
nand UO_1647 (O_1647,N_14926,N_14705);
nand UO_1648 (O_1648,N_14824,N_14984);
xnor UO_1649 (O_1649,N_14965,N_14777);
nor UO_1650 (O_1650,N_14909,N_14797);
and UO_1651 (O_1651,N_14902,N_14771);
nand UO_1652 (O_1652,N_14884,N_14744);
xor UO_1653 (O_1653,N_14961,N_14967);
nor UO_1654 (O_1654,N_14771,N_14850);
nor UO_1655 (O_1655,N_14896,N_14867);
xor UO_1656 (O_1656,N_14845,N_14718);
xnor UO_1657 (O_1657,N_14902,N_14914);
nand UO_1658 (O_1658,N_14735,N_14999);
nor UO_1659 (O_1659,N_14925,N_14791);
or UO_1660 (O_1660,N_14759,N_14874);
and UO_1661 (O_1661,N_14862,N_14736);
and UO_1662 (O_1662,N_14960,N_14758);
or UO_1663 (O_1663,N_14912,N_14953);
nor UO_1664 (O_1664,N_14803,N_14960);
or UO_1665 (O_1665,N_14926,N_14947);
and UO_1666 (O_1666,N_14877,N_14785);
or UO_1667 (O_1667,N_14856,N_14703);
or UO_1668 (O_1668,N_14858,N_14977);
xor UO_1669 (O_1669,N_14843,N_14906);
or UO_1670 (O_1670,N_14886,N_14921);
xnor UO_1671 (O_1671,N_14894,N_14850);
or UO_1672 (O_1672,N_14839,N_14933);
and UO_1673 (O_1673,N_14972,N_14815);
xnor UO_1674 (O_1674,N_14950,N_14916);
nand UO_1675 (O_1675,N_14709,N_14998);
nor UO_1676 (O_1676,N_14772,N_14749);
nor UO_1677 (O_1677,N_14750,N_14883);
nand UO_1678 (O_1678,N_14788,N_14767);
and UO_1679 (O_1679,N_14924,N_14772);
nand UO_1680 (O_1680,N_14911,N_14993);
nor UO_1681 (O_1681,N_14747,N_14908);
nor UO_1682 (O_1682,N_14772,N_14710);
nor UO_1683 (O_1683,N_14881,N_14845);
xnor UO_1684 (O_1684,N_14921,N_14856);
nand UO_1685 (O_1685,N_14855,N_14916);
or UO_1686 (O_1686,N_14739,N_14704);
nor UO_1687 (O_1687,N_14819,N_14964);
or UO_1688 (O_1688,N_14892,N_14989);
xnor UO_1689 (O_1689,N_14848,N_14802);
and UO_1690 (O_1690,N_14941,N_14797);
nand UO_1691 (O_1691,N_14831,N_14923);
nand UO_1692 (O_1692,N_14940,N_14818);
nor UO_1693 (O_1693,N_14700,N_14910);
nor UO_1694 (O_1694,N_14839,N_14869);
and UO_1695 (O_1695,N_14748,N_14702);
nand UO_1696 (O_1696,N_14948,N_14725);
xor UO_1697 (O_1697,N_14762,N_14962);
and UO_1698 (O_1698,N_14887,N_14817);
nor UO_1699 (O_1699,N_14937,N_14938);
and UO_1700 (O_1700,N_14930,N_14724);
nand UO_1701 (O_1701,N_14741,N_14936);
or UO_1702 (O_1702,N_14828,N_14832);
nand UO_1703 (O_1703,N_14784,N_14912);
nand UO_1704 (O_1704,N_14835,N_14777);
or UO_1705 (O_1705,N_14898,N_14880);
nand UO_1706 (O_1706,N_14745,N_14865);
nand UO_1707 (O_1707,N_14891,N_14972);
nor UO_1708 (O_1708,N_14717,N_14843);
nand UO_1709 (O_1709,N_14866,N_14714);
and UO_1710 (O_1710,N_14826,N_14900);
or UO_1711 (O_1711,N_14851,N_14973);
nand UO_1712 (O_1712,N_14720,N_14763);
nor UO_1713 (O_1713,N_14978,N_14713);
nand UO_1714 (O_1714,N_14939,N_14881);
or UO_1715 (O_1715,N_14880,N_14818);
nor UO_1716 (O_1716,N_14991,N_14742);
nor UO_1717 (O_1717,N_14914,N_14947);
xnor UO_1718 (O_1718,N_14867,N_14995);
xor UO_1719 (O_1719,N_14879,N_14761);
and UO_1720 (O_1720,N_14768,N_14941);
and UO_1721 (O_1721,N_14862,N_14837);
xor UO_1722 (O_1722,N_14893,N_14706);
nor UO_1723 (O_1723,N_14837,N_14767);
nor UO_1724 (O_1724,N_14913,N_14734);
and UO_1725 (O_1725,N_14772,N_14996);
nor UO_1726 (O_1726,N_14931,N_14801);
nor UO_1727 (O_1727,N_14994,N_14871);
nand UO_1728 (O_1728,N_14928,N_14757);
and UO_1729 (O_1729,N_14812,N_14883);
nor UO_1730 (O_1730,N_14905,N_14984);
or UO_1731 (O_1731,N_14788,N_14837);
and UO_1732 (O_1732,N_14756,N_14815);
or UO_1733 (O_1733,N_14891,N_14955);
nand UO_1734 (O_1734,N_14805,N_14787);
nand UO_1735 (O_1735,N_14709,N_14888);
and UO_1736 (O_1736,N_14783,N_14752);
or UO_1737 (O_1737,N_14714,N_14986);
nor UO_1738 (O_1738,N_14841,N_14909);
nor UO_1739 (O_1739,N_14901,N_14721);
or UO_1740 (O_1740,N_14703,N_14821);
and UO_1741 (O_1741,N_14750,N_14875);
or UO_1742 (O_1742,N_14925,N_14999);
nand UO_1743 (O_1743,N_14951,N_14956);
nor UO_1744 (O_1744,N_14950,N_14971);
xor UO_1745 (O_1745,N_14719,N_14989);
nand UO_1746 (O_1746,N_14712,N_14727);
xor UO_1747 (O_1747,N_14791,N_14834);
nand UO_1748 (O_1748,N_14970,N_14985);
or UO_1749 (O_1749,N_14808,N_14983);
xor UO_1750 (O_1750,N_14803,N_14919);
and UO_1751 (O_1751,N_14950,N_14787);
and UO_1752 (O_1752,N_14727,N_14878);
and UO_1753 (O_1753,N_14896,N_14793);
nand UO_1754 (O_1754,N_14942,N_14992);
or UO_1755 (O_1755,N_14914,N_14823);
nor UO_1756 (O_1756,N_14851,N_14877);
xnor UO_1757 (O_1757,N_14857,N_14951);
nand UO_1758 (O_1758,N_14980,N_14831);
or UO_1759 (O_1759,N_14946,N_14760);
and UO_1760 (O_1760,N_14776,N_14740);
or UO_1761 (O_1761,N_14942,N_14937);
nand UO_1762 (O_1762,N_14943,N_14725);
and UO_1763 (O_1763,N_14919,N_14839);
nand UO_1764 (O_1764,N_14789,N_14879);
xnor UO_1765 (O_1765,N_14718,N_14987);
nor UO_1766 (O_1766,N_14752,N_14720);
and UO_1767 (O_1767,N_14986,N_14762);
nand UO_1768 (O_1768,N_14839,N_14733);
or UO_1769 (O_1769,N_14881,N_14732);
nor UO_1770 (O_1770,N_14762,N_14766);
nand UO_1771 (O_1771,N_14750,N_14976);
and UO_1772 (O_1772,N_14708,N_14815);
nand UO_1773 (O_1773,N_14820,N_14778);
nand UO_1774 (O_1774,N_14859,N_14914);
xnor UO_1775 (O_1775,N_14984,N_14987);
and UO_1776 (O_1776,N_14885,N_14813);
and UO_1777 (O_1777,N_14928,N_14877);
nand UO_1778 (O_1778,N_14952,N_14966);
and UO_1779 (O_1779,N_14813,N_14982);
or UO_1780 (O_1780,N_14927,N_14843);
or UO_1781 (O_1781,N_14963,N_14918);
or UO_1782 (O_1782,N_14766,N_14925);
nor UO_1783 (O_1783,N_14772,N_14718);
xnor UO_1784 (O_1784,N_14885,N_14904);
nor UO_1785 (O_1785,N_14845,N_14740);
or UO_1786 (O_1786,N_14923,N_14890);
xor UO_1787 (O_1787,N_14994,N_14839);
xnor UO_1788 (O_1788,N_14900,N_14814);
nor UO_1789 (O_1789,N_14704,N_14915);
nand UO_1790 (O_1790,N_14880,N_14767);
nor UO_1791 (O_1791,N_14836,N_14777);
or UO_1792 (O_1792,N_14963,N_14894);
nand UO_1793 (O_1793,N_14802,N_14725);
or UO_1794 (O_1794,N_14888,N_14851);
nor UO_1795 (O_1795,N_14724,N_14946);
and UO_1796 (O_1796,N_14737,N_14895);
xor UO_1797 (O_1797,N_14726,N_14782);
xor UO_1798 (O_1798,N_14967,N_14783);
or UO_1799 (O_1799,N_14812,N_14998);
and UO_1800 (O_1800,N_14992,N_14798);
nand UO_1801 (O_1801,N_14920,N_14784);
xnor UO_1802 (O_1802,N_14820,N_14728);
nand UO_1803 (O_1803,N_14742,N_14946);
xnor UO_1804 (O_1804,N_14821,N_14820);
nor UO_1805 (O_1805,N_14735,N_14972);
or UO_1806 (O_1806,N_14900,N_14889);
xor UO_1807 (O_1807,N_14924,N_14747);
nand UO_1808 (O_1808,N_14965,N_14752);
or UO_1809 (O_1809,N_14946,N_14722);
nand UO_1810 (O_1810,N_14775,N_14702);
or UO_1811 (O_1811,N_14765,N_14984);
nand UO_1812 (O_1812,N_14990,N_14814);
nor UO_1813 (O_1813,N_14806,N_14814);
or UO_1814 (O_1814,N_14821,N_14993);
xnor UO_1815 (O_1815,N_14905,N_14787);
nor UO_1816 (O_1816,N_14793,N_14731);
or UO_1817 (O_1817,N_14714,N_14870);
and UO_1818 (O_1818,N_14929,N_14793);
and UO_1819 (O_1819,N_14823,N_14767);
nand UO_1820 (O_1820,N_14840,N_14867);
xor UO_1821 (O_1821,N_14982,N_14967);
xor UO_1822 (O_1822,N_14771,N_14969);
nand UO_1823 (O_1823,N_14958,N_14707);
or UO_1824 (O_1824,N_14834,N_14757);
nor UO_1825 (O_1825,N_14931,N_14915);
and UO_1826 (O_1826,N_14813,N_14883);
nand UO_1827 (O_1827,N_14988,N_14960);
xnor UO_1828 (O_1828,N_14999,N_14815);
and UO_1829 (O_1829,N_14814,N_14861);
nor UO_1830 (O_1830,N_14794,N_14823);
nor UO_1831 (O_1831,N_14994,N_14707);
nor UO_1832 (O_1832,N_14946,N_14949);
nand UO_1833 (O_1833,N_14831,N_14846);
and UO_1834 (O_1834,N_14986,N_14980);
nand UO_1835 (O_1835,N_14956,N_14748);
nand UO_1836 (O_1836,N_14915,N_14901);
xnor UO_1837 (O_1837,N_14820,N_14793);
nor UO_1838 (O_1838,N_14863,N_14986);
xnor UO_1839 (O_1839,N_14787,N_14811);
nand UO_1840 (O_1840,N_14833,N_14828);
xor UO_1841 (O_1841,N_14788,N_14769);
nor UO_1842 (O_1842,N_14731,N_14927);
nor UO_1843 (O_1843,N_14962,N_14823);
xor UO_1844 (O_1844,N_14761,N_14839);
nand UO_1845 (O_1845,N_14805,N_14902);
nand UO_1846 (O_1846,N_14824,N_14813);
xnor UO_1847 (O_1847,N_14706,N_14770);
nor UO_1848 (O_1848,N_14929,N_14770);
xnor UO_1849 (O_1849,N_14966,N_14707);
or UO_1850 (O_1850,N_14795,N_14911);
nor UO_1851 (O_1851,N_14951,N_14839);
nand UO_1852 (O_1852,N_14824,N_14874);
nand UO_1853 (O_1853,N_14883,N_14931);
xor UO_1854 (O_1854,N_14880,N_14885);
nor UO_1855 (O_1855,N_14789,N_14847);
and UO_1856 (O_1856,N_14819,N_14983);
or UO_1857 (O_1857,N_14717,N_14737);
xor UO_1858 (O_1858,N_14889,N_14943);
nand UO_1859 (O_1859,N_14936,N_14954);
and UO_1860 (O_1860,N_14967,N_14811);
xor UO_1861 (O_1861,N_14968,N_14842);
nand UO_1862 (O_1862,N_14947,N_14925);
nor UO_1863 (O_1863,N_14961,N_14735);
and UO_1864 (O_1864,N_14921,N_14884);
and UO_1865 (O_1865,N_14927,N_14871);
nor UO_1866 (O_1866,N_14839,N_14779);
nor UO_1867 (O_1867,N_14766,N_14949);
xnor UO_1868 (O_1868,N_14710,N_14978);
nor UO_1869 (O_1869,N_14840,N_14868);
or UO_1870 (O_1870,N_14741,N_14896);
nand UO_1871 (O_1871,N_14907,N_14728);
or UO_1872 (O_1872,N_14777,N_14839);
or UO_1873 (O_1873,N_14969,N_14759);
or UO_1874 (O_1874,N_14934,N_14737);
xnor UO_1875 (O_1875,N_14917,N_14900);
nor UO_1876 (O_1876,N_14920,N_14886);
and UO_1877 (O_1877,N_14791,N_14733);
nor UO_1878 (O_1878,N_14742,N_14799);
nor UO_1879 (O_1879,N_14943,N_14952);
nand UO_1880 (O_1880,N_14860,N_14972);
and UO_1881 (O_1881,N_14783,N_14852);
nor UO_1882 (O_1882,N_14856,N_14781);
or UO_1883 (O_1883,N_14713,N_14831);
nand UO_1884 (O_1884,N_14796,N_14783);
xor UO_1885 (O_1885,N_14818,N_14931);
and UO_1886 (O_1886,N_14747,N_14941);
and UO_1887 (O_1887,N_14964,N_14728);
nand UO_1888 (O_1888,N_14721,N_14730);
nand UO_1889 (O_1889,N_14999,N_14899);
and UO_1890 (O_1890,N_14727,N_14769);
nor UO_1891 (O_1891,N_14892,N_14967);
nor UO_1892 (O_1892,N_14903,N_14740);
and UO_1893 (O_1893,N_14726,N_14759);
or UO_1894 (O_1894,N_14720,N_14937);
nand UO_1895 (O_1895,N_14967,N_14814);
and UO_1896 (O_1896,N_14809,N_14778);
xnor UO_1897 (O_1897,N_14771,N_14755);
nor UO_1898 (O_1898,N_14910,N_14735);
and UO_1899 (O_1899,N_14959,N_14707);
nand UO_1900 (O_1900,N_14897,N_14870);
xnor UO_1901 (O_1901,N_14793,N_14921);
or UO_1902 (O_1902,N_14725,N_14938);
and UO_1903 (O_1903,N_14845,N_14830);
nand UO_1904 (O_1904,N_14971,N_14909);
nor UO_1905 (O_1905,N_14969,N_14757);
nor UO_1906 (O_1906,N_14922,N_14872);
nor UO_1907 (O_1907,N_14920,N_14801);
or UO_1908 (O_1908,N_14709,N_14951);
nor UO_1909 (O_1909,N_14967,N_14862);
xor UO_1910 (O_1910,N_14763,N_14868);
xor UO_1911 (O_1911,N_14758,N_14870);
xnor UO_1912 (O_1912,N_14829,N_14977);
xor UO_1913 (O_1913,N_14915,N_14764);
nand UO_1914 (O_1914,N_14918,N_14900);
nand UO_1915 (O_1915,N_14745,N_14944);
nor UO_1916 (O_1916,N_14847,N_14857);
and UO_1917 (O_1917,N_14956,N_14785);
nor UO_1918 (O_1918,N_14882,N_14910);
nor UO_1919 (O_1919,N_14799,N_14705);
nor UO_1920 (O_1920,N_14835,N_14783);
or UO_1921 (O_1921,N_14890,N_14968);
xor UO_1922 (O_1922,N_14974,N_14749);
nand UO_1923 (O_1923,N_14829,N_14725);
or UO_1924 (O_1924,N_14728,N_14864);
xnor UO_1925 (O_1925,N_14905,N_14824);
or UO_1926 (O_1926,N_14996,N_14744);
and UO_1927 (O_1927,N_14708,N_14740);
nand UO_1928 (O_1928,N_14743,N_14934);
nand UO_1929 (O_1929,N_14963,N_14890);
and UO_1930 (O_1930,N_14989,N_14787);
xor UO_1931 (O_1931,N_14847,N_14971);
or UO_1932 (O_1932,N_14832,N_14856);
xnor UO_1933 (O_1933,N_14983,N_14719);
nor UO_1934 (O_1934,N_14775,N_14925);
nand UO_1935 (O_1935,N_14721,N_14945);
or UO_1936 (O_1936,N_14896,N_14763);
xnor UO_1937 (O_1937,N_14783,N_14866);
xor UO_1938 (O_1938,N_14744,N_14723);
and UO_1939 (O_1939,N_14731,N_14919);
or UO_1940 (O_1940,N_14875,N_14738);
and UO_1941 (O_1941,N_14983,N_14754);
nor UO_1942 (O_1942,N_14836,N_14838);
and UO_1943 (O_1943,N_14923,N_14944);
or UO_1944 (O_1944,N_14859,N_14958);
xor UO_1945 (O_1945,N_14863,N_14840);
nor UO_1946 (O_1946,N_14727,N_14721);
nand UO_1947 (O_1947,N_14705,N_14803);
nand UO_1948 (O_1948,N_14779,N_14895);
nand UO_1949 (O_1949,N_14928,N_14943);
xnor UO_1950 (O_1950,N_14994,N_14841);
or UO_1951 (O_1951,N_14766,N_14906);
nand UO_1952 (O_1952,N_14968,N_14753);
nand UO_1953 (O_1953,N_14924,N_14713);
and UO_1954 (O_1954,N_14906,N_14983);
nand UO_1955 (O_1955,N_14869,N_14800);
xnor UO_1956 (O_1956,N_14820,N_14861);
or UO_1957 (O_1957,N_14823,N_14947);
nand UO_1958 (O_1958,N_14895,N_14863);
xor UO_1959 (O_1959,N_14764,N_14857);
or UO_1960 (O_1960,N_14911,N_14927);
xor UO_1961 (O_1961,N_14958,N_14783);
xor UO_1962 (O_1962,N_14742,N_14794);
nand UO_1963 (O_1963,N_14945,N_14829);
xor UO_1964 (O_1964,N_14942,N_14751);
nor UO_1965 (O_1965,N_14841,N_14900);
nand UO_1966 (O_1966,N_14715,N_14766);
nor UO_1967 (O_1967,N_14756,N_14879);
xnor UO_1968 (O_1968,N_14839,N_14754);
xnor UO_1969 (O_1969,N_14789,N_14904);
nand UO_1970 (O_1970,N_14731,N_14929);
and UO_1971 (O_1971,N_14876,N_14775);
or UO_1972 (O_1972,N_14874,N_14722);
xor UO_1973 (O_1973,N_14885,N_14711);
and UO_1974 (O_1974,N_14860,N_14847);
nand UO_1975 (O_1975,N_14964,N_14909);
nor UO_1976 (O_1976,N_14710,N_14851);
nor UO_1977 (O_1977,N_14970,N_14780);
or UO_1978 (O_1978,N_14745,N_14868);
xor UO_1979 (O_1979,N_14949,N_14748);
nand UO_1980 (O_1980,N_14864,N_14965);
and UO_1981 (O_1981,N_14897,N_14892);
xnor UO_1982 (O_1982,N_14723,N_14894);
xnor UO_1983 (O_1983,N_14706,N_14992);
nand UO_1984 (O_1984,N_14841,N_14824);
and UO_1985 (O_1985,N_14838,N_14721);
nand UO_1986 (O_1986,N_14741,N_14721);
and UO_1987 (O_1987,N_14906,N_14861);
nand UO_1988 (O_1988,N_14917,N_14826);
nor UO_1989 (O_1989,N_14902,N_14924);
or UO_1990 (O_1990,N_14909,N_14713);
and UO_1991 (O_1991,N_14895,N_14880);
and UO_1992 (O_1992,N_14969,N_14884);
and UO_1993 (O_1993,N_14940,N_14703);
nand UO_1994 (O_1994,N_14703,N_14862);
nand UO_1995 (O_1995,N_14794,N_14986);
or UO_1996 (O_1996,N_14735,N_14732);
nor UO_1997 (O_1997,N_14834,N_14907);
and UO_1998 (O_1998,N_14741,N_14894);
nand UO_1999 (O_1999,N_14917,N_14823);
endmodule