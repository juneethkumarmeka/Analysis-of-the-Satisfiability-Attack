module basic_2500_25000_3000_4_levels_5xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19025,N_19026,N_19027,N_19028,N_19029,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19186,N_19187,N_19188,N_19189,N_19190,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19253,N_19254,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19325,N_19326,N_19327,N_19328,N_19329,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19400,N_19401,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19464,N_19465,N_19466,N_19467,N_19469,N_19470,N_19471,N_19472,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19533,N_19534,N_19535,N_19536,N_19537,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19871,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19978,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19996,N_19997,N_19999,N_20000,N_20001,N_20002,N_20003,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20206,N_20207,N_20209,N_20210,N_20211,N_20212,N_20213,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20230,N_20231,N_20232,N_20234,N_20235,N_20236,N_20237,N_20238,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20363,N_20364,N_20365,N_20367,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20413,N_20414,N_20415,N_20416,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20458,N_20459,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20533,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_21000,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21376,N_21378,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21635,N_21636,N_21637,N_21638,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21736,N_21737,N_21738,N_21739,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22038,N_22039,N_22040,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22320,N_22321,N_22322,N_22323,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22839,N_22840,N_22841,N_22842,N_22844,N_22845,N_22846,N_22847,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22859,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22935,N_22936,N_22937,N_22938,N_22939,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23168,N_23169,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23561,N_23562,N_23563,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23732,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23872,N_23873,N_23874,N_23875,N_23876,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24066,N_24067,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24087,N_24089,N_24090,N_24091,N_24092,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24266,N_24267,N_24269,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24302,N_24303,N_24304,N_24305,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24488,N_24490,N_24491,N_24492,N_24493,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24521,N_24522,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24709,N_24710,N_24711,N_24712,N_24713,N_24715,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
or U0 (N_0,In_1337,In_101);
or U1 (N_1,In_246,In_77);
or U2 (N_2,In_334,In_1866);
and U3 (N_3,In_1184,In_2006);
nor U4 (N_4,In_1531,In_1366);
nor U5 (N_5,In_769,In_1657);
nor U6 (N_6,In_451,In_907);
nand U7 (N_7,In_1164,In_1524);
or U8 (N_8,In_641,In_2329);
nor U9 (N_9,In_2115,In_1559);
nor U10 (N_10,In_706,In_1112);
or U11 (N_11,In_532,In_885);
xor U12 (N_12,In_762,In_2281);
nor U13 (N_13,In_1514,In_1260);
nand U14 (N_14,In_845,In_2240);
nand U15 (N_15,In_2407,In_1257);
or U16 (N_16,In_349,In_1359);
and U17 (N_17,In_617,In_1379);
and U18 (N_18,In_1212,In_414);
nor U19 (N_19,In_312,In_1046);
nor U20 (N_20,In_2125,In_1110);
or U21 (N_21,In_780,In_1326);
or U22 (N_22,In_1828,In_2122);
and U23 (N_23,In_758,In_1729);
or U24 (N_24,In_289,In_87);
nand U25 (N_25,In_2018,In_757);
nor U26 (N_26,In_1087,In_2064);
nand U27 (N_27,In_1061,In_765);
nand U28 (N_28,In_2076,In_789);
and U29 (N_29,In_2192,In_1352);
and U30 (N_30,In_692,In_803);
nand U31 (N_31,In_248,In_1801);
nand U32 (N_32,In_2382,In_2171);
xnor U33 (N_33,In_2313,In_2442);
or U34 (N_34,In_1758,In_1195);
nand U35 (N_35,In_2424,In_1188);
nand U36 (N_36,In_936,In_1655);
or U37 (N_37,In_2188,In_1426);
xor U38 (N_38,In_982,In_639);
nor U39 (N_39,In_139,In_57);
and U40 (N_40,In_1398,In_2189);
nand U41 (N_41,In_2210,In_445);
nor U42 (N_42,In_1367,In_8);
or U43 (N_43,In_314,In_1011);
xor U44 (N_44,In_1249,In_1896);
and U45 (N_45,In_1662,In_2293);
nor U46 (N_46,In_150,In_350);
nand U47 (N_47,In_1295,In_1093);
or U48 (N_48,In_908,In_1939);
nand U49 (N_49,In_1837,In_2054);
nand U50 (N_50,In_914,In_1769);
nor U51 (N_51,In_1375,In_375);
xnor U52 (N_52,In_2147,In_186);
and U53 (N_53,In_183,In_233);
or U54 (N_54,In_657,In_2430);
and U55 (N_55,In_1245,In_524);
or U56 (N_56,In_1323,In_1667);
xor U57 (N_57,In_776,In_2203);
xor U58 (N_58,In_2426,In_1085);
nor U59 (N_59,In_2050,In_81);
or U60 (N_60,In_2110,In_2066);
nand U61 (N_61,In_748,In_1728);
nand U62 (N_62,In_2355,In_1401);
nor U63 (N_63,In_992,In_670);
or U64 (N_64,In_1380,In_1369);
nand U65 (N_65,In_1481,In_178);
xor U66 (N_66,In_1575,In_1621);
and U67 (N_67,In_1283,In_837);
xor U68 (N_68,In_1428,In_593);
nor U69 (N_69,In_841,In_2463);
and U70 (N_70,In_1607,In_550);
nor U71 (N_71,In_1176,In_2004);
nand U72 (N_72,In_1020,In_2146);
or U73 (N_73,In_2255,In_1127);
and U74 (N_74,In_2184,In_1392);
nor U75 (N_75,In_569,In_494);
or U76 (N_76,In_1450,In_1754);
xnor U77 (N_77,In_2428,In_440);
and U78 (N_78,In_1892,In_31);
nor U79 (N_79,In_1183,In_168);
nand U80 (N_80,In_2395,In_2116);
nand U81 (N_81,In_33,In_1010);
or U82 (N_82,In_927,In_324);
or U83 (N_83,In_26,In_2071);
and U84 (N_84,In_2303,In_516);
nor U85 (N_85,In_2237,In_731);
and U86 (N_86,In_2141,In_2261);
nand U87 (N_87,In_2423,In_277);
and U88 (N_88,In_503,In_1965);
and U89 (N_89,In_1564,In_408);
or U90 (N_90,In_22,In_2457);
nand U91 (N_91,In_1686,In_2316);
nand U92 (N_92,In_1290,In_467);
nor U93 (N_93,In_1731,In_1854);
xor U94 (N_94,In_1306,In_1605);
xor U95 (N_95,In_2140,In_1119);
nor U96 (N_96,In_1756,In_1037);
nand U97 (N_97,In_1318,In_106);
and U98 (N_98,In_1313,In_985);
nand U99 (N_99,In_1641,In_1882);
and U100 (N_100,In_2021,In_986);
nand U101 (N_101,In_2246,In_1623);
nand U102 (N_102,In_1272,In_1515);
nand U103 (N_103,In_2485,In_1873);
nor U104 (N_104,In_1252,In_736);
and U105 (N_105,In_142,In_1000);
nor U106 (N_106,In_1957,In_751);
and U107 (N_107,In_1064,In_1682);
and U108 (N_108,In_935,In_1904);
and U109 (N_109,In_423,In_589);
xor U110 (N_110,In_1142,In_2175);
or U111 (N_111,In_665,In_660);
or U112 (N_112,In_327,In_2222);
xor U113 (N_113,In_1973,In_942);
nand U114 (N_114,In_2165,In_1421);
or U115 (N_115,In_357,In_416);
or U116 (N_116,In_259,In_1441);
nand U117 (N_117,In_1884,In_2160);
xor U118 (N_118,In_717,In_664);
nor U119 (N_119,In_505,In_2086);
and U120 (N_120,In_1237,In_869);
or U121 (N_121,In_216,In_1031);
or U122 (N_122,In_1130,In_12);
nand U123 (N_123,In_1557,In_632);
nand U124 (N_124,In_1258,In_1716);
and U125 (N_125,In_431,In_1143);
and U126 (N_126,In_2164,In_1541);
nand U127 (N_127,In_439,In_2363);
nand U128 (N_128,In_2392,In_1717);
or U129 (N_129,In_622,In_586);
nand U130 (N_130,In_604,In_669);
nand U131 (N_131,In_1256,In_2080);
or U132 (N_132,In_2072,In_1674);
nand U133 (N_133,In_1096,In_1362);
xor U134 (N_134,In_1349,In_605);
and U135 (N_135,In_412,In_954);
xnor U136 (N_136,In_1587,In_2221);
nor U137 (N_137,In_556,In_1689);
nor U138 (N_138,In_95,In_1972);
xnor U139 (N_139,In_1203,In_1156);
and U140 (N_140,In_1343,In_1786);
or U141 (N_141,In_298,In_797);
or U142 (N_142,In_760,In_1592);
and U143 (N_143,In_976,In_678);
nand U144 (N_144,In_2475,In_1415);
nand U145 (N_145,In_2204,In_268);
or U146 (N_146,In_1719,In_1453);
nand U147 (N_147,In_1849,In_666);
or U148 (N_148,In_1660,In_192);
and U149 (N_149,In_46,In_689);
xnor U150 (N_150,In_112,In_5);
nand U151 (N_151,In_235,In_2254);
or U152 (N_152,In_1395,In_2307);
or U153 (N_153,In_577,In_1498);
nor U154 (N_154,In_1806,In_1937);
or U155 (N_155,In_713,In_174);
or U156 (N_156,In_307,In_273);
or U157 (N_157,In_1800,In_902);
and U158 (N_158,In_286,In_482);
or U159 (N_159,In_1779,In_293);
and U160 (N_160,In_13,In_103);
nor U161 (N_161,In_828,In_1547);
nor U162 (N_162,In_1831,In_2301);
nand U163 (N_163,In_170,In_462);
xnor U164 (N_164,In_2036,In_86);
xnor U165 (N_165,In_671,In_1981);
nor U166 (N_166,In_1799,In_177);
or U167 (N_167,In_1693,In_283);
or U168 (N_168,In_994,In_965);
and U169 (N_169,In_650,In_924);
and U170 (N_170,In_2191,In_2119);
or U171 (N_171,In_1763,In_1107);
and U172 (N_172,In_1467,In_455);
nor U173 (N_173,In_2262,In_1646);
or U174 (N_174,In_1906,In_1386);
nor U175 (N_175,In_2497,In_2335);
or U176 (N_176,In_1797,In_160);
and U177 (N_177,In_1509,In_137);
nand U178 (N_178,In_30,In_661);
and U179 (N_179,In_529,In_1566);
nor U180 (N_180,In_2354,In_2443);
nor U181 (N_181,In_834,In_971);
or U182 (N_182,In_1676,In_164);
nand U183 (N_183,In_683,In_1893);
and U184 (N_184,In_2317,In_242);
nand U185 (N_185,In_1132,In_2067);
nor U186 (N_186,In_539,In_1824);
or U187 (N_187,In_860,In_970);
or U188 (N_188,In_1919,In_620);
and U189 (N_189,In_2228,In_1472);
nand U190 (N_190,In_2142,In_2233);
and U191 (N_191,In_2121,In_1014);
nand U192 (N_192,In_1140,In_1712);
xnor U193 (N_193,In_899,In_1139);
and U194 (N_194,In_694,In_93);
or U195 (N_195,In_321,In_502);
and U196 (N_196,In_1992,In_397);
nor U197 (N_197,In_351,In_1118);
or U198 (N_198,In_999,In_117);
or U199 (N_199,In_880,In_972);
nand U200 (N_200,In_1852,In_996);
or U201 (N_201,In_598,In_311);
or U202 (N_202,In_1659,In_688);
and U203 (N_203,In_2253,In_1840);
and U204 (N_204,In_681,In_2450);
or U205 (N_205,In_1262,In_1340);
or U206 (N_206,In_1320,In_481);
xnor U207 (N_207,In_572,In_1865);
nand U208 (N_208,In_113,In_1294);
and U209 (N_209,In_1781,In_738);
and U210 (N_210,In_1200,In_1572);
and U211 (N_211,In_690,In_1325);
xnor U212 (N_212,In_804,In_1608);
and U213 (N_213,In_1982,In_1846);
nor U214 (N_214,In_1264,In_1382);
and U215 (N_215,In_411,In_236);
xnor U216 (N_216,In_1739,In_2098);
or U217 (N_217,In_2062,In_166);
or U218 (N_218,In_2389,In_879);
or U219 (N_219,In_653,In_1815);
or U220 (N_220,In_119,In_1791);
nand U221 (N_221,In_1850,In_1927);
nand U222 (N_222,In_1796,In_1813);
nand U223 (N_223,In_2367,In_1172);
and U224 (N_224,In_1247,In_1170);
nor U225 (N_225,In_612,In_1309);
or U226 (N_226,In_17,In_1400);
nand U227 (N_227,In_2042,In_2492);
nand U228 (N_228,In_14,In_450);
and U229 (N_229,In_2084,In_781);
and U230 (N_230,In_1568,In_234);
and U231 (N_231,In_2238,In_1098);
or U232 (N_232,In_1502,In_1049);
nand U233 (N_233,In_517,In_2333);
xnor U234 (N_234,In_858,In_1876);
or U235 (N_235,In_2352,In_1335);
or U236 (N_236,In_2077,In_1371);
and U237 (N_237,In_92,In_1926);
nand U238 (N_238,In_303,In_365);
and U239 (N_239,In_2490,In_2386);
or U240 (N_240,In_2187,In_1416);
nor U241 (N_241,In_470,In_11);
nor U242 (N_242,In_562,In_558);
and U243 (N_243,In_2200,In_266);
nand U244 (N_244,In_2266,In_1825);
nor U245 (N_245,In_1629,In_721);
and U246 (N_246,In_1021,In_764);
nand U247 (N_247,In_332,In_114);
nor U248 (N_248,In_2208,In_2153);
and U249 (N_249,In_2046,In_722);
nor U250 (N_250,In_1522,In_606);
and U251 (N_251,In_1534,In_1696);
nand U252 (N_252,In_306,In_1417);
or U253 (N_253,In_295,In_1947);
nand U254 (N_254,In_1289,In_1962);
nor U255 (N_255,In_857,In_2069);
xnor U256 (N_256,In_1631,In_495);
xor U257 (N_257,In_1388,In_730);
xnor U258 (N_258,In_1241,In_2111);
or U259 (N_259,In_1339,In_2414);
or U260 (N_260,In_1776,In_1069);
and U261 (N_261,In_488,In_405);
nor U262 (N_262,In_1594,In_537);
nand U263 (N_263,In_648,In_1553);
nor U264 (N_264,In_15,In_1869);
and U265 (N_265,In_1802,In_1617);
xor U266 (N_266,In_1701,In_2406);
and U267 (N_267,In_342,In_275);
nor U268 (N_268,In_91,In_566);
nor U269 (N_269,In_1868,In_1597);
and U270 (N_270,In_1685,In_1698);
and U271 (N_271,In_313,In_424);
nand U272 (N_272,In_527,In_2251);
or U273 (N_273,In_2309,In_461);
xnor U274 (N_274,In_1993,In_1749);
nand U275 (N_275,In_403,In_2195);
and U276 (N_276,In_1787,In_887);
nor U277 (N_277,In_1711,In_1439);
and U278 (N_278,In_1527,In_1651);
or U279 (N_279,In_479,In_1333);
or U280 (N_280,In_1554,In_1591);
and U281 (N_281,In_132,In_1720);
nand U282 (N_282,In_833,In_2059);
nor U283 (N_283,In_382,In_1773);
nor U284 (N_284,In_107,In_711);
xnor U285 (N_285,In_1723,In_1954);
xor U286 (N_286,In_2305,In_1206);
or U287 (N_287,In_652,In_919);
nand U288 (N_288,In_476,In_2132);
and U289 (N_289,In_794,In_1533);
nand U290 (N_290,In_1016,In_2483);
and U291 (N_291,In_131,In_2390);
nand U292 (N_292,In_581,In_767);
nand U293 (N_293,In_2136,In_76);
nor U294 (N_294,In_2431,In_2090);
nor U295 (N_295,In_1956,In_436);
nor U296 (N_296,In_120,In_507);
nor U297 (N_297,In_2365,In_1671);
or U298 (N_298,In_55,In_161);
and U299 (N_299,In_154,In_2462);
nand U300 (N_300,In_2276,In_1518);
and U301 (N_301,In_1028,In_2044);
nor U302 (N_302,In_251,In_1297);
or U303 (N_303,In_1454,In_2405);
and U304 (N_304,In_715,In_2338);
nor U305 (N_305,In_469,In_1963);
or U306 (N_306,In_883,In_1690);
xor U307 (N_307,In_946,In_1826);
nand U308 (N_308,In_1878,In_1032);
nor U309 (N_309,In_1035,In_2170);
or U310 (N_310,In_2214,In_2114);
and U311 (N_311,In_2473,In_460);
or U312 (N_312,In_214,In_844);
nor U313 (N_313,In_873,In_963);
and U314 (N_314,In_948,In_1268);
nand U315 (N_315,In_145,In_535);
nand U316 (N_316,In_1699,In_2020);
and U317 (N_317,In_1473,In_536);
or U318 (N_318,In_2011,In_1480);
nand U319 (N_319,In_1510,In_404);
and U320 (N_320,In_143,In_2229);
nor U321 (N_321,In_2271,In_2138);
or U322 (N_322,In_512,In_1210);
or U323 (N_323,In_1665,In_1910);
or U324 (N_324,In_2244,In_68);
xor U325 (N_325,In_1034,In_2133);
nor U326 (N_326,In_185,In_737);
nand U327 (N_327,In_1603,In_1135);
nor U328 (N_328,In_975,In_1948);
nand U329 (N_329,In_741,In_2026);
or U330 (N_330,In_1742,In_2479);
xnor U331 (N_331,In_1780,In_1635);
and U332 (N_332,In_381,In_1669);
xnor U333 (N_333,In_1025,In_1538);
and U334 (N_334,In_753,In_50);
nor U335 (N_335,In_474,In_1908);
or U336 (N_336,In_1223,In_1209);
nor U337 (N_337,In_2369,In_1990);
nand U338 (N_338,In_1161,In_1979);
nor U339 (N_339,In_441,In_2033);
nand U340 (N_340,In_2498,In_659);
nand U341 (N_341,In_220,In_618);
nor U342 (N_342,In_1331,In_83);
nand U343 (N_343,In_2014,In_795);
nand U344 (N_344,In_2101,In_38);
and U345 (N_345,In_1714,In_705);
or U346 (N_346,In_60,In_247);
nand U347 (N_347,In_1038,In_2275);
or U348 (N_348,In_2408,In_1471);
or U349 (N_349,In_41,In_600);
or U350 (N_350,In_637,In_124);
and U351 (N_351,In_1404,In_1234);
nand U352 (N_352,In_1765,In_513);
xor U353 (N_353,In_232,In_563);
nor U354 (N_354,In_1961,In_54);
and U355 (N_355,In_169,In_1839);
nor U356 (N_356,In_1059,In_1879);
or U357 (N_357,In_511,In_1785);
or U358 (N_358,In_1269,In_878);
nor U359 (N_359,In_1497,In_1341);
nand U360 (N_360,In_2264,In_2433);
nand U361 (N_361,In_1120,In_1909);
and U362 (N_362,In_1980,In_2263);
or U363 (N_363,In_2093,In_1073);
or U364 (N_364,In_1642,In_1013);
and U365 (N_365,In_2081,In_830);
nand U366 (N_366,In_2087,In_1935);
or U367 (N_367,In_379,In_1610);
or U368 (N_368,In_1647,In_2061);
or U369 (N_369,In_135,In_65);
nor U370 (N_370,In_1108,In_1745);
xor U371 (N_371,In_1726,In_853);
nand U372 (N_372,In_2332,In_783);
nand U373 (N_373,In_759,In_231);
nor U374 (N_374,In_1520,In_920);
nor U375 (N_375,In_2057,In_2350);
and U376 (N_376,In_595,In_94);
and U377 (N_377,In_1949,In_2009);
or U378 (N_378,In_2190,In_2124);
and U379 (N_379,In_2104,In_554);
nor U380 (N_380,In_1503,In_667);
nand U381 (N_381,In_480,In_262);
nand U382 (N_382,In_1158,In_928);
nor U383 (N_383,In_2480,In_702);
nand U384 (N_384,In_1040,In_2312);
nand U385 (N_385,In_2465,In_1571);
and U386 (N_386,In_634,In_2477);
nor U387 (N_387,In_1478,In_2144);
nand U388 (N_388,In_2314,In_1602);
nand U389 (N_389,In_1422,In_2274);
nand U390 (N_390,In_2048,In_1934);
nand U391 (N_391,In_892,In_709);
nor U392 (N_392,In_1946,In_320);
and U393 (N_393,In_2419,In_208);
and U394 (N_394,In_2489,In_1823);
nor U395 (N_395,In_73,In_257);
nor U396 (N_396,In_2447,In_193);
xnor U397 (N_397,In_952,In_2356);
nor U398 (N_398,In_1296,In_209);
nand U399 (N_399,In_888,In_1736);
or U400 (N_400,In_1880,In_360);
or U401 (N_401,In_1584,In_319);
xor U402 (N_402,In_1162,In_1638);
nand U403 (N_403,In_1407,In_725);
nand U404 (N_404,In_299,In_1881);
nand U405 (N_405,In_933,In_84);
or U406 (N_406,In_2280,In_1902);
or U407 (N_407,In_1163,In_561);
nand U408 (N_408,In_36,In_410);
nand U409 (N_409,In_2211,In_1793);
and U410 (N_410,In_1692,In_823);
and U411 (N_411,In_1001,In_548);
nor U412 (N_412,In_1221,In_1084);
nor U413 (N_413,In_1194,In_1319);
and U414 (N_414,In_1871,In_1875);
nor U415 (N_415,In_701,In_1540);
nand U416 (N_416,In_1966,In_2085);
nand U417 (N_417,In_2055,In_2045);
xor U418 (N_418,In_194,In_1895);
xor U419 (N_419,In_624,In_1899);
xnor U420 (N_420,In_227,In_149);
nor U421 (N_421,In_2287,In_932);
xor U422 (N_422,In_1933,In_323);
nor U423 (N_423,In_1894,In_1886);
nor U424 (N_424,In_698,In_1004);
and U425 (N_425,In_656,In_1921);
nor U426 (N_426,In_2396,In_627);
or U427 (N_427,In_2242,In_3);
and U428 (N_428,In_2092,In_80);
or U429 (N_429,In_1137,In_574);
or U430 (N_430,In_1991,In_237);
nor U431 (N_431,In_1431,In_534);
and U432 (N_432,In_465,In_2385);
or U433 (N_433,In_1370,In_1457);
nand U434 (N_434,In_1435,In_1207);
nand U435 (N_435,In_1298,In_1039);
and U436 (N_436,In_1490,In_364);
nand U437 (N_437,In_422,In_1687);
nand U438 (N_438,In_1500,In_255);
and U439 (N_439,In_1626,In_300);
xnor U440 (N_440,In_1704,In_1483);
or U441 (N_441,In_1350,In_1412);
nand U442 (N_442,In_1075,In_1746);
or U443 (N_443,In_1233,In_318);
or U444 (N_444,In_2278,In_2182);
or U445 (N_445,In_2288,In_180);
and U446 (N_446,In_425,In_891);
nand U447 (N_447,In_1987,In_339);
and U448 (N_448,In_2401,In_1694);
nor U449 (N_449,In_129,In_40);
xnor U450 (N_450,In_1389,In_2464);
and U451 (N_451,In_294,In_1009);
nand U452 (N_452,In_865,In_2323);
or U453 (N_453,In_925,In_1443);
and U454 (N_454,In_889,In_1002);
or U455 (N_455,In_1271,In_584);
or U456 (N_456,In_1440,In_374);
and U457 (N_457,In_2375,In_361);
nand U458 (N_458,In_281,In_1134);
and U459 (N_459,In_1618,In_1938);
or U460 (N_460,In_2118,In_2260);
nand U461 (N_461,In_551,In_1627);
or U462 (N_462,In_787,In_733);
nand U463 (N_463,In_1166,In_1253);
nor U464 (N_464,In_337,In_610);
or U465 (N_465,In_2285,In_48);
nand U466 (N_466,In_520,In_1474);
or U467 (N_467,In_1589,In_815);
or U468 (N_468,In_34,In_1818);
nand U469 (N_469,In_1705,In_2013);
or U470 (N_470,In_2102,In_181);
and U471 (N_471,In_1236,In_591);
nand U472 (N_472,In_1266,In_10);
nand U473 (N_473,In_402,In_1585);
or U474 (N_474,In_1606,In_203);
or U475 (N_475,In_642,In_419);
nor U476 (N_476,In_2010,In_2035);
nor U477 (N_477,In_1387,In_2100);
and U478 (N_478,In_1710,In_2482);
or U479 (N_479,In_1914,In_1857);
and U480 (N_480,In_571,In_955);
nor U481 (N_481,In_140,In_2034);
xor U482 (N_482,In_317,In_1616);
nor U483 (N_483,In_842,In_1688);
and U484 (N_484,In_1707,In_2345);
nand U485 (N_485,In_583,In_2448);
nor U486 (N_486,In_1214,In_1402);
nand U487 (N_487,In_1461,In_243);
and U488 (N_488,In_1622,In_1361);
and U489 (N_489,In_2008,In_2);
nand U490 (N_490,In_1877,In_1812);
or U491 (N_491,In_2403,In_358);
and U492 (N_492,In_1066,In_974);
nor U493 (N_493,In_2041,In_373);
nand U494 (N_494,In_213,In_2223);
and U495 (N_495,In_839,In_212);
or U496 (N_496,In_1834,In_813);
nand U497 (N_497,In_1955,In_1446);
and U498 (N_498,In_1177,In_2476);
nor U499 (N_499,In_173,In_1887);
nand U500 (N_500,In_1543,In_1654);
nor U501 (N_501,In_1764,In_827);
nand U502 (N_502,In_260,In_2272);
xor U503 (N_503,In_1775,In_1102);
nor U504 (N_504,In_744,In_2232);
and U505 (N_505,In_1625,In_1770);
nand U506 (N_506,In_644,In_1488);
nand U507 (N_507,In_745,In_2353);
nor U508 (N_508,In_1639,In_9);
nor U509 (N_509,In_742,In_2466);
nand U510 (N_510,In_1327,In_63);
xor U511 (N_511,In_1144,In_1519);
or U512 (N_512,In_2012,In_676);
or U513 (N_513,In_949,In_1310);
nor U514 (N_514,In_542,In_207);
and U515 (N_515,In_388,In_1218);
or U516 (N_516,In_1250,In_872);
nand U517 (N_517,In_710,In_956);
nand U518 (N_518,In_728,In_2319);
xnor U519 (N_519,In_1077,In_1109);
or U520 (N_520,In_2331,In_1810);
and U521 (N_521,In_906,In_1023);
nor U522 (N_522,In_1805,In_239);
or U523 (N_523,In_1501,In_575);
or U524 (N_524,In_472,In_110);
nor U525 (N_525,In_1019,In_1464);
nor U526 (N_526,In_704,In_2056);
and U527 (N_527,In_1024,In_343);
or U528 (N_528,In_2183,In_219);
and U529 (N_529,In_631,In_662);
nor U530 (N_530,In_1232,In_1795);
nand U531 (N_531,In_1358,In_750);
and U532 (N_532,In_1442,In_102);
or U533 (N_533,In_724,In_2032);
and U534 (N_534,In_2197,In_1489);
xnor U535 (N_535,In_398,In_1219);
nand U536 (N_536,In_2371,In_2306);
xnor U537 (N_537,In_1578,In_1149);
and U538 (N_538,In_1652,In_981);
or U539 (N_539,In_400,In_2181);
nand U540 (N_540,In_541,In_1215);
nor U541 (N_541,In_1315,In_2145);
nand U542 (N_542,In_1867,In_740);
nand U543 (N_543,In_1640,In_967);
nor U544 (N_544,In_921,In_2341);
nand U545 (N_545,In_39,In_2364);
and U546 (N_546,In_824,In_2163);
and U547 (N_547,In_1596,In_1111);
nor U548 (N_548,In_775,In_134);
nand U549 (N_549,In_1858,In_296);
nor U550 (N_550,In_2030,In_226);
nand U551 (N_551,In_2470,In_1737);
or U552 (N_552,In_947,In_1141);
nand U553 (N_553,In_401,In_732);
or U554 (N_554,In_1190,In_1372);
nor U555 (N_555,In_2215,In_943);
nor U556 (N_556,In_1433,In_2284);
nor U557 (N_557,In_1008,In_1827);
nand U558 (N_558,In_1978,In_254);
nor U559 (N_559,In_1374,In_2446);
nor U560 (N_560,In_614,In_396);
nor U561 (N_561,In_893,In_1964);
and U562 (N_562,In_377,In_362);
or U563 (N_563,In_1276,In_2366);
and U564 (N_564,In_961,In_1280);
nand U565 (N_565,In_1322,In_1573);
and U566 (N_566,In_67,In_636);
xor U567 (N_567,In_2294,In_1491);
xnor U568 (N_568,In_697,In_1094);
nor U569 (N_569,In_2321,In_2231);
or U570 (N_570,In_153,In_2220);
nand U571 (N_571,In_1700,In_210);
nand U572 (N_572,In_52,In_66);
nand U573 (N_573,In_2436,In_1917);
xor U574 (N_574,In_719,In_2474);
and U575 (N_575,In_1357,In_1444);
nand U576 (N_576,In_779,In_1124);
or U577 (N_577,In_2455,In_2001);
and U578 (N_578,In_746,In_2089);
xor U579 (N_579,In_126,In_1383);
or U580 (N_580,In_1479,In_1609);
nand U581 (N_581,In_387,In_2201);
and U582 (N_582,In_348,In_23);
and U583 (N_583,In_1345,In_2387);
nor U584 (N_584,In_2007,In_2016);
and U585 (N_585,In_696,In_1168);
and U586 (N_586,In_1732,In_851);
nor U587 (N_587,In_2429,In_301);
nor U588 (N_588,In_1410,In_1356);
xnor U589 (N_589,In_700,In_456);
and U590 (N_590,In_1076,In_1542);
nor U591 (N_591,In_58,In_2308);
or U592 (N_592,In_1044,In_687);
xnor U593 (N_593,In_647,In_2368);
nand U594 (N_594,In_1462,In_684);
nand U595 (N_595,In_786,In_386);
nor U596 (N_596,In_2486,In_1673);
nor U597 (N_597,In_1872,In_1018);
xnor U598 (N_598,In_2162,In_1959);
or U599 (N_599,In_1281,In_1808);
xnor U600 (N_600,In_1744,In_47);
and U601 (N_601,In_1804,In_1248);
nand U602 (N_602,In_71,In_1274);
nand U603 (N_603,In_61,In_1516);
or U604 (N_604,In_272,In_1208);
and U605 (N_605,In_1300,In_2344);
xnor U606 (N_606,In_877,In_1278);
nor U607 (N_607,In_1027,In_1684);
or U608 (N_608,In_2005,In_88);
nand U609 (N_609,In_6,In_2298);
and U610 (N_610,In_1136,In_394);
nand U611 (N_611,In_1944,In_831);
xnor U612 (N_612,In_874,In_432);
or U613 (N_613,In_2091,In_2402);
and U614 (N_614,In_448,In_621);
or U615 (N_615,In_1539,In_2258);
and U616 (N_616,In_2252,In_543);
nand U617 (N_617,In_1299,In_304);
nor U618 (N_618,In_1664,In_2404);
nand U619 (N_619,In_1782,In_1907);
nor U620 (N_620,In_1513,In_847);
or U621 (N_621,In_329,In_987);
nor U622 (N_622,In_1492,In_1675);
and U623 (N_623,In_1121,In_1153);
and U624 (N_624,In_151,In_1619);
xnor U625 (N_625,In_1586,In_1321);
and U626 (N_626,In_167,In_1192);
nand U627 (N_627,In_1169,In_1324);
and U628 (N_628,In_2340,In_2444);
nand U629 (N_629,In_818,In_1943);
nand U630 (N_630,In_1661,In_2247);
nand U631 (N_631,In_1653,In_2299);
nor U632 (N_632,In_1403,In_1809);
and U633 (N_633,In_325,In_2234);
nand U634 (N_634,In_1680,In_2441);
and U635 (N_635,In_1870,In_1983);
nor U636 (N_636,In_1406,In_2346);
nor U637 (N_637,In_1958,In_1182);
nand U638 (N_638,In_1259,In_680);
or U639 (N_639,In_2279,In_1465);
xnor U640 (N_640,In_245,In_1279);
or U641 (N_641,In_587,In_1434);
nand U642 (N_642,In_130,In_1942);
nor U643 (N_643,In_718,In_894);
and U644 (N_644,In_770,In_163);
and U645 (N_645,In_1565,In_1506);
and U646 (N_646,In_478,In_2304);
nor U647 (N_647,In_1856,In_1555);
or U648 (N_648,In_1495,In_1523);
and U649 (N_649,In_1173,In_1579);
or U650 (N_650,In_2172,In_1752);
xor U651 (N_651,In_1614,In_56);
and U652 (N_652,In_898,In_434);
and U653 (N_653,In_2206,In_2213);
nand U654 (N_654,In_1577,In_991);
nor U655 (N_655,In_316,In_922);
and U656 (N_656,In_70,In_547);
nor U657 (N_657,In_1792,In_805);
and U658 (N_658,In_72,In_1042);
or U659 (N_659,In_2399,In_582);
nor U660 (N_660,In_930,In_1329);
and U661 (N_661,In_1448,In_2265);
or U662 (N_662,In_1985,In_2174);
nor U663 (N_663,In_1063,In_1929);
and U664 (N_664,In_2282,In_2360);
and U665 (N_665,In_870,In_2472);
and U666 (N_666,In_1159,In_2028);
and U667 (N_667,In_148,In_1974);
and U668 (N_668,In_1836,In_983);
nand U669 (N_669,In_2158,In_1548);
nor U670 (N_670,In_515,In_2449);
nand U671 (N_671,In_2166,In_1054);
nand U672 (N_672,In_1521,In_1157);
xor U673 (N_673,In_2373,In_206);
nand U674 (N_674,In_549,In_2380);
nand U675 (N_675,In_1537,In_1832);
and U676 (N_676,In_1022,In_335);
and U677 (N_677,In_2453,In_336);
and U678 (N_678,In_929,In_729);
and U679 (N_679,In_640,In_265);
nand U680 (N_680,In_123,In_290);
nand U681 (N_681,In_2393,In_881);
or U682 (N_682,In_2216,In_1709);
nand U683 (N_683,In_1181,In_2015);
nor U684 (N_684,In_544,In_1855);
nor U685 (N_685,In_2148,In_308);
nand U686 (N_686,In_217,In_490);
xnor U687 (N_687,In_2416,In_1911);
xor U688 (N_688,In_579,In_35);
or U689 (N_689,In_1423,In_2194);
nor U690 (N_690,In_133,In_2250);
nor U691 (N_691,In_1468,In_1224);
and U692 (N_692,In_1859,In_1405);
nand U693 (N_693,In_668,In_1251);
nand U694 (N_694,In_2243,In_1811);
and U695 (N_695,In_1220,In_1185);
and U696 (N_696,In_1302,In_802);
nor U697 (N_697,In_2039,In_1486);
and U698 (N_698,In_172,In_829);
or U699 (N_699,In_900,In_1360);
and U700 (N_700,In_1819,In_449);
or U701 (N_701,In_1466,In_1920);
and U702 (N_702,In_2461,In_663);
or U703 (N_703,In_2378,In_2432);
nand U704 (N_704,In_944,In_221);
and U705 (N_705,In_816,In_1117);
and U706 (N_706,In_1790,In_1385);
nand U707 (N_707,In_1438,In_200);
nor U708 (N_708,In_785,In_1202);
and U709 (N_709,In_121,In_32);
or U710 (N_710,In_1377,In_810);
nand U711 (N_711,In_1560,In_2002);
nand U712 (N_712,In_2219,In_848);
nor U713 (N_713,In_1390,In_596);
and U714 (N_714,In_1384,In_1003);
nand U715 (N_715,In_225,In_1912);
or U716 (N_716,In_1235,In_2196);
xnor U717 (N_717,In_2257,In_526);
and U718 (N_718,In_836,In_2040);
and U719 (N_719,In_493,In_1766);
nor U720 (N_720,In_162,In_2202);
or U721 (N_721,In_1767,In_1007);
and U722 (N_722,In_1864,In_726);
and U723 (N_723,In_825,In_2178);
nand U724 (N_724,In_958,In_471);
xor U725 (N_725,In_310,In_658);
or U726 (N_726,In_1267,In_176);
xor U727 (N_727,In_2047,In_1725);
nor U728 (N_728,In_2337,In_792);
or U729 (N_729,In_165,In_2289);
and U730 (N_730,In_2412,In_158);
nor U731 (N_731,In_1291,In_2273);
or U732 (N_732,In_2325,In_1860);
and U733 (N_733,In_1941,In_409);
nor U734 (N_734,In_264,In_2079);
nor U735 (N_735,In_691,In_159);
nor U736 (N_736,In_1097,In_2411);
nand U737 (N_737,In_1658,In_292);
nor U738 (N_738,In_1691,In_2459);
nand U739 (N_739,In_261,In_2456);
nor U740 (N_740,In_806,In_649);
nor U741 (N_741,In_1905,In_438);
nor U742 (N_742,In_2239,In_754);
nor U743 (N_743,In_814,In_1637);
nor U744 (N_744,In_1351,In_1487);
nand U745 (N_745,In_1050,In_2458);
nand U746 (N_746,In_105,In_979);
nor U747 (N_747,In_2088,In_1068);
xor U748 (N_748,In_1342,In_997);
or U749 (N_749,In_832,In_2417);
and U750 (N_750,In_1888,In_2126);
and U751 (N_751,In_279,In_393);
xor U752 (N_752,In_2043,In_501);
nand U753 (N_753,In_980,In_1128);
and U754 (N_754,In_720,In_1649);
nor U755 (N_755,In_399,In_138);
or U756 (N_756,In_1734,In_2495);
nor U757 (N_757,In_1317,In_1580);
nor U758 (N_758,In_735,In_1048);
and U759 (N_759,In_1216,In_196);
nor U760 (N_760,In_2290,In_1822);
and U761 (N_761,In_1043,In_1969);
nand U762 (N_762,In_1078,In_1970);
or U763 (N_763,In_707,In_2400);
nand U764 (N_764,In_2025,In_288);
nor U765 (N_765,In_1505,In_1175);
and U766 (N_766,In_1463,In_1430);
xor U767 (N_767,In_428,In_1079);
and U768 (N_768,In_1930,In_568);
and U769 (N_769,In_791,In_1475);
nand U770 (N_770,In_915,In_1449);
or U771 (N_771,In_695,In_886);
and U772 (N_772,In_1951,In_884);
and U773 (N_773,In_187,In_1612);
or U774 (N_774,In_1240,In_2075);
xor U775 (N_775,In_826,In_2139);
nor U776 (N_776,In_1774,In_2017);
nor U777 (N_777,In_2438,In_2128);
nand U778 (N_778,In_1601,In_1683);
or U779 (N_779,In_1238,In_1074);
nand U780 (N_780,In_497,In_1469);
nand U781 (N_781,In_1145,In_1115);
nor U782 (N_782,In_1552,In_2471);
nor U783 (N_783,In_1376,In_2027);
or U784 (N_784,In_1088,In_1845);
xor U785 (N_785,In_2179,In_2248);
or U786 (N_786,In_1645,In_190);
nor U787 (N_787,In_457,In_385);
nand U788 (N_788,In_2023,In_468);
nor U789 (N_789,In_2421,In_1425);
and U790 (N_790,In_1945,In_241);
nand U791 (N_791,In_2381,In_433);
and U792 (N_792,In_859,In_484);
nor U793 (N_793,In_309,In_1485);
and U794 (N_794,In_356,In_1517);
nor U795 (N_795,In_28,In_1604);
xor U796 (N_796,In_466,In_1844);
and U797 (N_797,In_53,In_699);
nor U798 (N_798,In_1217,In_18);
xnor U799 (N_799,In_2113,In_799);
nand U800 (N_800,In_601,In_2349);
or U801 (N_801,In_2060,In_228);
nand U802 (N_802,In_1628,In_147);
and U803 (N_803,In_2209,In_1198);
nand U804 (N_804,In_1570,In_1613);
nor U805 (N_805,In_523,In_951);
nor U806 (N_806,In_2488,In_615);
nor U807 (N_807,In_1330,In_452);
nor U808 (N_808,In_2391,In_1814);
or U809 (N_809,In_485,In_2058);
or U810 (N_810,In_1663,In_1995);
nor U811 (N_811,In_995,In_21);
nand U812 (N_812,In_1432,In_723);
or U813 (N_813,In_2224,In_1151);
and U814 (N_814,In_2478,In_2499);
and U815 (N_815,In_359,In_1051);
nand U816 (N_816,In_766,In_1529);
or U817 (N_817,In_1397,In_808);
nor U818 (N_818,In_96,In_2420);
or U819 (N_819,In_1470,In_2112);
nor U820 (N_820,In_1284,In_911);
xnor U821 (N_821,In_1060,In_863);
nor U822 (N_822,In_609,In_2445);
nand U823 (N_823,In_1741,In_843);
nor U824 (N_824,In_654,In_1355);
and U825 (N_825,In_90,In_1740);
or U826 (N_826,In_49,In_2347);
and U827 (N_827,In_1666,In_2131);
nor U828 (N_828,In_1225,In_2484);
or U829 (N_829,In_182,In_1065);
nor U830 (N_830,In_2063,In_918);
nor U831 (N_831,In_2302,In_1830);
or U832 (N_832,In_2177,In_623);
and U833 (N_833,In_1842,In_44);
nand U834 (N_834,In_1748,In_1615);
nor U835 (N_835,In_852,In_2370);
and U836 (N_836,In_2397,In_218);
nand U837 (N_837,In_1598,In_1885);
nand U838 (N_838,In_491,In_1286);
and U839 (N_839,In_2460,In_2109);
nor U840 (N_840,In_1057,In_146);
and U841 (N_841,In_777,In_1082);
xor U842 (N_842,In_968,In_413);
xor U843 (N_843,In_817,In_2467);
or U844 (N_844,In_1952,In_1545);
or U845 (N_845,In_1147,In_2398);
and U846 (N_846,In_2096,In_672);
or U847 (N_847,In_679,In_1817);
or U848 (N_848,In_7,In_1427);
nor U849 (N_849,In_580,In_64);
nand U850 (N_850,In_525,In_2388);
and U851 (N_851,In_1316,In_1301);
and U852 (N_852,In_1724,In_2343);
nor U853 (N_853,In_444,In_1146);
or U854 (N_854,In_1644,In_2134);
nand U855 (N_855,In_2051,In_1624);
nor U856 (N_856,In_1455,In_1532);
or U857 (N_857,In_1925,In_1750);
and U858 (N_858,In_291,In_2225);
and U859 (N_859,In_1530,In_655);
or U860 (N_860,In_1496,In_2049);
nand U861 (N_861,In_2031,In_1988);
nor U862 (N_862,In_778,In_211);
nand U863 (N_863,In_189,In_1999);
xnor U864 (N_864,In_633,In_16);
nor U865 (N_865,In_2270,In_1936);
nand U866 (N_866,In_1986,In_1556);
nor U867 (N_867,In_59,In_1191);
or U868 (N_868,In_2019,In_1263);
nor U869 (N_869,In_1678,In_2212);
and U870 (N_870,In_1015,In_2103);
nor U871 (N_871,In_761,In_1620);
xnor U872 (N_872,In_2318,In_2073);
and U873 (N_873,In_1436,In_1155);
nand U874 (N_874,In_1650,In_1582);
xor U875 (N_875,In_1989,In_973);
and U876 (N_876,In_1563,In_945);
or U877 (N_877,In_686,In_240);
nand U878 (N_878,In_198,In_521);
nor U879 (N_879,In_415,In_2259);
and U880 (N_880,In_270,In_1931);
nor U881 (N_881,In_258,In_406);
or U882 (N_882,In_628,In_854);
or U883 (N_883,In_1308,In_518);
nand U884 (N_884,In_2469,In_984);
or U885 (N_885,In_504,In_821);
and U886 (N_886,In_99,In_1794);
or U887 (N_887,In_939,In_1747);
and U888 (N_888,In_2143,In_1347);
or U889 (N_889,In_597,In_1771);
nor U890 (N_890,In_1484,In_1975);
nor U891 (N_891,In_1095,In_1451);
and U892 (N_892,In_788,In_499);
or U893 (N_893,In_1903,In_2351);
and U894 (N_894,In_346,In_909);
or U895 (N_895,In_1273,In_1006);
and U896 (N_896,In_703,In_1196);
and U897 (N_897,In_913,In_395);
and U898 (N_898,In_341,In_2267);
and U899 (N_899,In_199,In_1730);
and U900 (N_900,In_1820,In_1525);
and U901 (N_901,In_376,In_533);
xor U902 (N_902,In_1239,In_682);
nor U903 (N_903,In_905,In_1544);
and U904 (N_904,In_1072,In_553);
and U905 (N_905,In_1030,In_1364);
xor U906 (N_906,In_1636,In_613);
nand U907 (N_907,In_122,In_1713);
and U908 (N_908,In_371,In_1230);
and U909 (N_909,In_1368,In_2358);
and U910 (N_910,In_937,In_1677);
or U911 (N_911,In_2117,In_838);
nor U912 (N_912,In_1706,In_1968);
nand U913 (N_913,In_510,In_1967);
xor U914 (N_914,In_673,In_1045);
nand U915 (N_915,In_1311,In_1226);
xor U916 (N_916,In_1131,In_1265);
nor U917 (N_917,In_202,In_2159);
and U918 (N_918,In_1197,In_1447);
and U919 (N_919,In_1148,In_1456);
nor U920 (N_920,In_876,In_800);
or U921 (N_921,In_1154,In_1976);
xor U922 (N_922,In_819,In_391);
or U923 (N_923,In_1703,In_368);
nor U924 (N_924,In_903,In_530);
nor U925 (N_925,In_1549,In_136);
nor U926 (N_926,In_1922,In_1199);
xor U927 (N_927,In_1898,In_1254);
or U928 (N_928,In_2230,In_616);
and U929 (N_929,In_1399,In_2468);
or U930 (N_930,In_565,In_674);
and U931 (N_931,In_1588,In_1816);
nor U932 (N_932,In_380,In_849);
or U933 (N_933,In_2422,In_1751);
or U934 (N_934,In_384,In_1721);
or U935 (N_935,In_223,In_473);
or U936 (N_936,In_2434,In_37);
and U937 (N_937,In_287,In_638);
nor U938 (N_938,In_302,In_1104);
or U939 (N_939,In_1648,In_85);
nand U940 (N_940,In_1755,In_1971);
nor U941 (N_941,In_2120,In_2029);
nor U942 (N_942,In_2249,In_152);
xnor U943 (N_943,In_1213,In_812);
nor U944 (N_944,In_2135,In_835);
and U945 (N_945,In_1753,In_347);
nor U946 (N_946,In_2130,In_2106);
and U947 (N_947,In_2161,In_184);
nand U948 (N_948,In_901,In_2193);
nand U949 (N_949,In_1546,In_2186);
xor U950 (N_950,In_693,In_0);
nor U951 (N_951,In_486,In_1874);
xnor U952 (N_952,In_755,In_2286);
xnor U953 (N_953,In_1477,In_1821);
nand U954 (N_954,In_426,In_1656);
xor U955 (N_955,In_442,In_2137);
nor U956 (N_956,In_2435,In_2291);
or U957 (N_957,In_1508,In_383);
nor U958 (N_958,In_1843,In_1798);
or U959 (N_959,In_1735,In_2095);
and U960 (N_960,In_2328,In_1285);
xnor U961 (N_961,In_1915,In_1883);
or U962 (N_962,In_1344,In_895);
nand U963 (N_963,In_500,In_603);
xnor U964 (N_964,In_1070,In_390);
nand U965 (N_965,In_278,In_1697);
nand U966 (N_966,In_369,In_840);
nor U967 (N_967,In_602,In_1348);
and U968 (N_968,In_352,In_904);
or U969 (N_969,In_111,In_1996);
or U970 (N_970,In_2327,In_2082);
nand U971 (N_971,In_1924,In_1160);
or U972 (N_972,In_864,In_2384);
nor U973 (N_973,In_716,In_1633);
and U974 (N_974,In_338,In_483);
nor U975 (N_975,In_978,In_127);
and U976 (N_976,In_782,In_1055);
or U977 (N_977,In_345,In_626);
nor U978 (N_978,In_538,In_2123);
and U979 (N_979,In_630,In_1133);
or U980 (N_980,In_1630,In_29);
xnor U981 (N_981,In_98,In_1353);
or U982 (N_982,In_608,In_2496);
nand U983 (N_983,In_2339,In_1420);
nor U984 (N_984,In_1103,In_2074);
nand U985 (N_985,In_2207,In_197);
nor U986 (N_986,In_1762,In_97);
and U987 (N_987,In_222,In_590);
or U988 (N_988,In_1228,In_790);
nand U989 (N_989,In_2491,In_2198);
nand U990 (N_990,In_2334,In_1833);
nor U991 (N_991,In_370,In_1336);
nor U992 (N_992,In_389,In_454);
xnor U993 (N_993,In_45,In_798);
nor U994 (N_994,In_2357,In_1174);
xor U995 (N_995,In_89,In_429);
and U996 (N_996,In_1179,In_714);
or U997 (N_997,In_25,In_867);
nor U998 (N_998,In_959,In_645);
and U999 (N_999,In_2394,In_1599);
and U1000 (N_1000,In_447,In_1760);
nor U1001 (N_1001,In_940,In_407);
and U1002 (N_1002,In_2283,In_1314);
nand U1003 (N_1003,In_2277,In_2413);
xor U1004 (N_1004,In_917,In_328);
or U1005 (N_1005,In_896,In_1058);
nand U1006 (N_1006,In_1201,In_578);
xnor U1007 (N_1007,In_923,In_2493);
nand U1008 (N_1008,In_1994,In_1092);
nand U1009 (N_1009,In_1152,In_1026);
nor U1010 (N_1010,In_82,In_191);
and U1011 (N_1011,In_1838,In_871);
and U1012 (N_1012,In_331,In_2383);
or U1013 (N_1013,In_24,In_1114);
or U1014 (N_1014,In_363,In_969);
and U1015 (N_1015,In_756,In_496);
and U1016 (N_1016,In_856,In_875);
xor U1017 (N_1017,In_2454,In_1312);
and U1018 (N_1018,In_2199,In_2218);
or U1019 (N_1019,In_475,In_2362);
or U1020 (N_1020,In_2226,In_560);
or U1021 (N_1021,In_557,In_2149);
and U1022 (N_1022,In_1738,In_576);
nand U1023 (N_1023,In_367,In_1901);
nand U1024 (N_1024,In_1890,In_477);
xor U1025 (N_1025,In_2361,In_509);
or U1026 (N_1026,In_912,In_1950);
nor U1027 (N_1027,In_1365,In_646);
and U1028 (N_1028,In_1180,In_253);
or U1029 (N_1029,In_1891,In_238);
and U1030 (N_1030,In_2176,In_2418);
and U1031 (N_1031,In_2205,In_1100);
nand U1032 (N_1032,In_204,In_2326);
nand U1033 (N_1033,In_774,In_446);
nor U1034 (N_1034,In_1581,In_1918);
nor U1035 (N_1035,In_1129,In_2235);
nand U1036 (N_1036,In_950,In_811);
nor U1037 (N_1037,In_1551,In_1727);
nor U1038 (N_1038,In_230,In_205);
nor U1039 (N_1039,In_459,In_807);
nor U1040 (N_1040,In_1733,In_966);
or U1041 (N_1041,In_685,In_531);
or U1042 (N_1042,In_1244,In_19);
nand U1043 (N_1043,In_1507,In_179);
nor U1044 (N_1044,In_1101,In_100);
nor U1045 (N_1045,In_1122,In_267);
or U1046 (N_1046,In_625,In_1086);
or U1047 (N_1047,In_1851,In_555);
nand U1048 (N_1048,In_1071,In_594);
xnor U1049 (N_1049,In_1165,In_1561);
nand U1050 (N_1050,In_573,In_2003);
nand U1051 (N_1051,In_1668,In_1445);
nand U1052 (N_1052,In_464,In_69);
or U1053 (N_1053,In_1632,In_1080);
xnor U1054 (N_1054,In_74,In_2024);
nand U1055 (N_1055,In_1067,In_938);
nor U1056 (N_1056,In_675,In_392);
and U1057 (N_1057,In_417,In_749);
and U1058 (N_1058,In_366,In_1702);
and U1059 (N_1059,In_570,In_1772);
or U1060 (N_1060,In_340,In_2425);
and U1061 (N_1061,In_868,In_599);
xor U1062 (N_1062,In_1229,In_1287);
nand U1063 (N_1063,In_1504,In_1718);
nor U1064 (N_1064,In_326,In_1913);
and U1065 (N_1065,In_2150,In_2156);
nand U1066 (N_1066,In_353,In_1848);
nand U1067 (N_1067,In_1062,In_1611);
nor U1068 (N_1068,In_1670,In_1036);
nand U1069 (N_1069,In_1106,In_1222);
nand U1070 (N_1070,In_201,In_78);
and U1071 (N_1071,In_964,In_1381);
nor U1072 (N_1072,In_1275,In_1123);
nor U1073 (N_1073,In_2376,In_1408);
nor U1074 (N_1074,In_977,In_771);
nor U1075 (N_1075,In_1889,In_1803);
xnor U1076 (N_1076,In_619,In_1807);
and U1077 (N_1077,In_4,In_1960);
nand U1078 (N_1078,In_354,In_1783);
xnor U1079 (N_1079,In_1334,In_27);
and U1080 (N_1080,In_1715,In_784);
nand U1081 (N_1081,In_75,In_188);
and U1082 (N_1082,In_993,In_1012);
nor U1083 (N_1083,In_1460,In_1338);
nand U1084 (N_1084,In_1411,In_1424);
xor U1085 (N_1085,In_1923,In_712);
and U1086 (N_1086,In_2439,In_344);
nor U1087 (N_1087,In_1998,In_1307);
or U1088 (N_1088,In_1784,In_250);
or U1089 (N_1089,In_2105,In_1997);
and U1090 (N_1090,In_1029,In_1105);
xor U1091 (N_1091,In_229,In_651);
nand U1092 (N_1092,In_2037,In_611);
nand U1093 (N_1093,In_355,In_271);
nand U1094 (N_1094,In_941,In_1761);
nand U1095 (N_1095,In_916,In_1778);
nor U1096 (N_1096,In_1550,In_171);
nand U1097 (N_1097,In_269,In_1354);
and U1098 (N_1098,In_453,In_1681);
nand U1099 (N_1099,In_2000,In_1759);
nor U1100 (N_1100,In_1459,In_1743);
nor U1101 (N_1101,In_42,In_2359);
nor U1102 (N_1102,In_2129,In_1757);
or U1103 (N_1103,In_1396,In_378);
nand U1104 (N_1104,In_1041,In_2481);
xnor U1105 (N_1105,In_2241,In_1005);
and U1106 (N_1106,In_1288,In_282);
nor U1107 (N_1107,In_1113,In_1270);
nand U1108 (N_1108,In_20,In_708);
and U1109 (N_1109,In_796,In_458);
or U1110 (N_1110,In_2097,In_989);
and U1111 (N_1111,In_2151,In_773);
nor U1112 (N_1112,In_244,In_2256);
nor U1113 (N_1113,In_435,In_988);
and U1114 (N_1114,In_1231,In_104);
nand U1115 (N_1115,In_421,In_1414);
or U1116 (N_1116,In_1413,In_1595);
nand U1117 (N_1117,In_157,In_333);
and U1118 (N_1118,In_155,In_546);
nor U1119 (N_1119,In_498,In_2295);
or U1120 (N_1120,In_1116,In_215);
xor U1121 (N_1121,In_990,In_276);
nor U1122 (N_1122,In_2322,In_1567);
and U1123 (N_1123,In_2167,In_1788);
nor U1124 (N_1124,In_1282,In_1409);
nor U1125 (N_1125,In_592,In_1841);
xor U1126 (N_1126,In_763,In_2168);
or U1127 (N_1127,In_252,In_2038);
xor U1128 (N_1128,In_528,In_1277);
nand U1129 (N_1129,In_2296,In_1476);
nor U1130 (N_1130,In_1862,In_156);
and U1131 (N_1131,In_2127,In_855);
and U1132 (N_1132,In_2180,In_1391);
nor U1133 (N_1133,In_809,In_585);
nand U1134 (N_1134,In_897,In_1722);
nand U1135 (N_1135,In_2494,In_2108);
or U1136 (N_1136,In_2083,In_2227);
and U1137 (N_1137,In_727,In_2094);
nor U1138 (N_1138,In_882,In_1017);
nand U1139 (N_1139,In_118,In_2315);
nand U1140 (N_1140,In_1847,In_1033);
or U1141 (N_1141,In_108,In_1512);
and U1142 (N_1142,In_1305,In_2269);
nand U1143 (N_1143,In_1499,In_1695);
or U1144 (N_1144,In_443,In_1511);
and U1145 (N_1145,In_2336,In_1091);
nand U1146 (N_1146,In_734,In_747);
xnor U1147 (N_1147,In_420,In_2022);
nor U1148 (N_1148,In_305,In_801);
or U1149 (N_1149,In_1292,In_1679);
or U1150 (N_1150,In_1193,In_1363);
nor U1151 (N_1151,In_1056,In_1242);
or U1152 (N_1152,In_2374,In_1634);
or U1153 (N_1153,In_567,In_1293);
nor U1154 (N_1154,In_629,In_2173);
nor U1155 (N_1155,In_559,In_1977);
and U1156 (N_1156,In_1829,In_1576);
nor U1157 (N_1157,In_2330,In_1227);
nor U1158 (N_1158,In_1777,In_2245);
or U1159 (N_1159,In_1255,In_427);
xnor U1160 (N_1160,In_1394,In_1768);
nand U1161 (N_1161,In_926,In_2155);
nand U1162 (N_1162,In_489,In_522);
nand U1163 (N_1163,In_79,In_1);
or U1164 (N_1164,In_820,In_1090);
and U1165 (N_1165,In_545,In_862);
nor U1166 (N_1166,In_1126,In_953);
xor U1167 (N_1167,In_910,In_1643);
or U1168 (N_1168,In_1482,In_1171);
nand U1169 (N_1169,In_1261,In_1535);
nand U1170 (N_1170,In_2440,In_866);
xnor U1171 (N_1171,In_1150,In_2451);
nor U1172 (N_1172,In_772,In_934);
nor U1173 (N_1173,In_284,In_1187);
and U1174 (N_1174,In_1167,In_144);
or U1175 (N_1175,In_846,In_2070);
nand U1176 (N_1176,In_957,In_2310);
and U1177 (N_1177,In_2415,In_1081);
nor U1178 (N_1178,In_2410,In_768);
or U1179 (N_1179,In_1863,In_2379);
or U1180 (N_1180,In_1897,In_1528);
or U1181 (N_1181,In_2342,In_2437);
nor U1182 (N_1182,In_2372,In_175);
and U1183 (N_1183,In_1672,In_1419);
or U1184 (N_1184,In_1204,In_822);
xnor U1185 (N_1185,In_962,In_1178);
nor U1186 (N_1186,In_2292,In_280);
and U1187 (N_1187,In_315,In_2099);
and U1188 (N_1188,In_1429,In_793);
nand U1189 (N_1189,In_297,In_1099);
nand U1190 (N_1190,In_372,In_109);
and U1191 (N_1191,In_1452,In_2068);
and U1192 (N_1192,In_1304,In_677);
nor U1193 (N_1193,In_1047,In_540);
and U1194 (N_1194,In_125,In_1189);
nor U1195 (N_1195,In_263,In_1984);
nand U1196 (N_1196,In_2154,In_1600);
nor U1197 (N_1197,In_195,In_1853);
xnor U1198 (N_1198,In_463,In_1493);
or U1199 (N_1199,In_1494,In_2297);
and U1200 (N_1200,In_2377,In_931);
or U1201 (N_1201,In_1089,In_51);
and U1202 (N_1202,In_2324,In_861);
nand U1203 (N_1203,In_1569,In_2217);
and U1204 (N_1204,In_2107,In_2078);
nor U1205 (N_1205,In_1186,In_1583);
nand U1206 (N_1206,In_1458,In_1940);
or U1207 (N_1207,In_2065,In_1861);
nand U1208 (N_1208,In_2320,In_128);
xnor U1209 (N_1209,In_1835,In_998);
or U1210 (N_1210,In_635,In_2052);
nand U1211 (N_1211,In_1053,In_552);
nor U1212 (N_1212,In_1789,In_1211);
nor U1213 (N_1213,In_1437,In_2157);
nand U1214 (N_1214,In_514,In_1373);
and U1215 (N_1215,In_437,In_752);
and U1216 (N_1216,In_1590,In_1558);
and U1217 (N_1217,In_1303,In_274);
nand U1218 (N_1218,In_1243,In_2409);
or U1219 (N_1219,In_1953,In_322);
nand U1220 (N_1220,In_430,In_1346);
and U1221 (N_1221,In_1246,In_1418);
or U1222 (N_1222,In_224,In_487);
or U1223 (N_1223,In_2236,In_2268);
nor U1224 (N_1224,In_960,In_418);
xnor U1225 (N_1225,In_2169,In_2152);
xnor U1226 (N_1226,In_1932,In_2300);
nor U1227 (N_1227,In_1328,In_607);
or U1228 (N_1228,In_643,In_1332);
nor U1229 (N_1229,In_739,In_1536);
nor U1230 (N_1230,In_2487,In_330);
or U1231 (N_1231,In_1378,In_1708);
nor U1232 (N_1232,In_2311,In_1526);
nor U1233 (N_1233,In_1562,In_2427);
and U1234 (N_1234,In_850,In_249);
nor U1235 (N_1235,In_1574,In_508);
or U1236 (N_1236,In_1205,In_116);
or U1237 (N_1237,In_1138,In_1393);
and U1238 (N_1238,In_2185,In_1916);
xor U1239 (N_1239,In_492,In_1593);
and U1240 (N_1240,In_519,In_62);
xnor U1241 (N_1241,In_890,In_1125);
and U1242 (N_1242,In_2452,In_2053);
or U1243 (N_1243,In_115,In_1928);
or U1244 (N_1244,In_1083,In_43);
and U1245 (N_1245,In_743,In_1900);
nand U1246 (N_1246,In_2348,In_588);
nand U1247 (N_1247,In_506,In_285);
nand U1248 (N_1248,In_256,In_1052);
nor U1249 (N_1249,In_564,In_141);
and U1250 (N_1250,In_82,In_197);
nand U1251 (N_1251,In_693,In_2368);
nand U1252 (N_1252,In_885,In_1952);
nor U1253 (N_1253,In_359,In_1867);
nor U1254 (N_1254,In_1642,In_2072);
and U1255 (N_1255,In_1085,In_2180);
or U1256 (N_1256,In_1615,In_2497);
nand U1257 (N_1257,In_1631,In_146);
and U1258 (N_1258,In_608,In_2001);
or U1259 (N_1259,In_1647,In_32);
or U1260 (N_1260,In_2065,In_160);
or U1261 (N_1261,In_431,In_1436);
or U1262 (N_1262,In_84,In_1539);
nand U1263 (N_1263,In_116,In_1823);
and U1264 (N_1264,In_1037,In_1417);
and U1265 (N_1265,In_2005,In_265);
nor U1266 (N_1266,In_1086,In_182);
nor U1267 (N_1267,In_575,In_2058);
xnor U1268 (N_1268,In_2394,In_1029);
or U1269 (N_1269,In_1265,In_1671);
nor U1270 (N_1270,In_231,In_2004);
and U1271 (N_1271,In_1004,In_2246);
and U1272 (N_1272,In_880,In_202);
xnor U1273 (N_1273,In_403,In_954);
xnor U1274 (N_1274,In_1109,In_1433);
xor U1275 (N_1275,In_18,In_68);
nand U1276 (N_1276,In_1078,In_1648);
nand U1277 (N_1277,In_1903,In_1403);
xnor U1278 (N_1278,In_1428,In_2191);
and U1279 (N_1279,In_1308,In_2490);
and U1280 (N_1280,In_809,In_616);
nor U1281 (N_1281,In_783,In_1231);
nor U1282 (N_1282,In_1968,In_699);
or U1283 (N_1283,In_971,In_1245);
and U1284 (N_1284,In_80,In_472);
nor U1285 (N_1285,In_484,In_1473);
and U1286 (N_1286,In_1976,In_1113);
and U1287 (N_1287,In_348,In_37);
nand U1288 (N_1288,In_681,In_2471);
nand U1289 (N_1289,In_2113,In_1054);
nor U1290 (N_1290,In_2306,In_1625);
and U1291 (N_1291,In_836,In_1742);
and U1292 (N_1292,In_1060,In_2237);
xnor U1293 (N_1293,In_624,In_5);
or U1294 (N_1294,In_834,In_2113);
xnor U1295 (N_1295,In_219,In_1856);
or U1296 (N_1296,In_494,In_2032);
nor U1297 (N_1297,In_1866,In_939);
nor U1298 (N_1298,In_2035,In_675);
nor U1299 (N_1299,In_1687,In_1882);
or U1300 (N_1300,In_1276,In_2457);
nand U1301 (N_1301,In_509,In_1879);
xnor U1302 (N_1302,In_2374,In_774);
xnor U1303 (N_1303,In_1758,In_1346);
and U1304 (N_1304,In_2097,In_1070);
nand U1305 (N_1305,In_2378,In_1875);
nor U1306 (N_1306,In_1760,In_1071);
xor U1307 (N_1307,In_1396,In_884);
xnor U1308 (N_1308,In_1104,In_2017);
nor U1309 (N_1309,In_1382,In_404);
or U1310 (N_1310,In_775,In_847);
or U1311 (N_1311,In_2438,In_2032);
nor U1312 (N_1312,In_1293,In_903);
nor U1313 (N_1313,In_684,In_198);
xnor U1314 (N_1314,In_2042,In_2208);
and U1315 (N_1315,In_2433,In_1991);
and U1316 (N_1316,In_1337,In_2247);
and U1317 (N_1317,In_2297,In_2163);
nand U1318 (N_1318,In_648,In_1118);
or U1319 (N_1319,In_2067,In_747);
nor U1320 (N_1320,In_1323,In_1854);
nand U1321 (N_1321,In_1591,In_601);
nor U1322 (N_1322,In_1215,In_246);
nand U1323 (N_1323,In_1690,In_660);
and U1324 (N_1324,In_1131,In_2160);
nand U1325 (N_1325,In_41,In_2122);
xor U1326 (N_1326,In_925,In_623);
or U1327 (N_1327,In_1519,In_98);
xor U1328 (N_1328,In_298,In_764);
nand U1329 (N_1329,In_1184,In_1519);
and U1330 (N_1330,In_1506,In_927);
and U1331 (N_1331,In_568,In_980);
nand U1332 (N_1332,In_1226,In_1748);
and U1333 (N_1333,In_2496,In_1075);
or U1334 (N_1334,In_1425,In_1747);
and U1335 (N_1335,In_566,In_2353);
nand U1336 (N_1336,In_1635,In_1303);
xnor U1337 (N_1337,In_1767,In_2300);
and U1338 (N_1338,In_1830,In_1229);
and U1339 (N_1339,In_1827,In_1723);
or U1340 (N_1340,In_1608,In_1718);
nand U1341 (N_1341,In_39,In_1653);
nor U1342 (N_1342,In_2291,In_313);
xor U1343 (N_1343,In_2109,In_1916);
nand U1344 (N_1344,In_651,In_1585);
nand U1345 (N_1345,In_790,In_2135);
and U1346 (N_1346,In_2145,In_66);
or U1347 (N_1347,In_765,In_2297);
nor U1348 (N_1348,In_839,In_2094);
nand U1349 (N_1349,In_1968,In_605);
nand U1350 (N_1350,In_944,In_807);
and U1351 (N_1351,In_264,In_1754);
nor U1352 (N_1352,In_1189,In_2375);
or U1353 (N_1353,In_2359,In_626);
nand U1354 (N_1354,In_1957,In_502);
nor U1355 (N_1355,In_1334,In_1137);
nor U1356 (N_1356,In_810,In_1434);
or U1357 (N_1357,In_1085,In_571);
or U1358 (N_1358,In_1615,In_1629);
nor U1359 (N_1359,In_1596,In_365);
nor U1360 (N_1360,In_2290,In_122);
nor U1361 (N_1361,In_2148,In_471);
and U1362 (N_1362,In_1987,In_144);
or U1363 (N_1363,In_1356,In_1812);
nand U1364 (N_1364,In_24,In_189);
nand U1365 (N_1365,In_2104,In_1137);
nor U1366 (N_1366,In_81,In_157);
or U1367 (N_1367,In_1555,In_810);
nor U1368 (N_1368,In_1630,In_685);
xnor U1369 (N_1369,In_665,In_1264);
nand U1370 (N_1370,In_878,In_2159);
or U1371 (N_1371,In_1590,In_2342);
nor U1372 (N_1372,In_1350,In_1677);
nand U1373 (N_1373,In_1777,In_3);
or U1374 (N_1374,In_195,In_483);
and U1375 (N_1375,In_2486,In_289);
and U1376 (N_1376,In_2364,In_2436);
nor U1377 (N_1377,In_2368,In_616);
nand U1378 (N_1378,In_1060,In_2117);
nor U1379 (N_1379,In_1000,In_1748);
nand U1380 (N_1380,In_2070,In_1280);
nand U1381 (N_1381,In_29,In_1636);
nor U1382 (N_1382,In_1221,In_176);
nand U1383 (N_1383,In_959,In_2134);
nand U1384 (N_1384,In_328,In_37);
and U1385 (N_1385,In_1151,In_1932);
nor U1386 (N_1386,In_2481,In_2011);
xnor U1387 (N_1387,In_1412,In_1162);
or U1388 (N_1388,In_2360,In_505);
xor U1389 (N_1389,In_2066,In_371);
or U1390 (N_1390,In_658,In_1497);
and U1391 (N_1391,In_43,In_1351);
nand U1392 (N_1392,In_1125,In_1151);
or U1393 (N_1393,In_425,In_1562);
and U1394 (N_1394,In_2283,In_88);
xor U1395 (N_1395,In_1075,In_39);
xor U1396 (N_1396,In_2361,In_215);
nand U1397 (N_1397,In_1321,In_1275);
and U1398 (N_1398,In_2054,In_2222);
and U1399 (N_1399,In_1792,In_1727);
nand U1400 (N_1400,In_1754,In_801);
or U1401 (N_1401,In_1747,In_1216);
nand U1402 (N_1402,In_242,In_237);
or U1403 (N_1403,In_981,In_2252);
xor U1404 (N_1404,In_1182,In_1262);
xor U1405 (N_1405,In_1290,In_500);
or U1406 (N_1406,In_1587,In_1442);
or U1407 (N_1407,In_2306,In_1165);
nor U1408 (N_1408,In_2079,In_2032);
nor U1409 (N_1409,In_1982,In_1416);
or U1410 (N_1410,In_592,In_2420);
nand U1411 (N_1411,In_1578,In_1277);
or U1412 (N_1412,In_595,In_171);
nand U1413 (N_1413,In_2313,In_1231);
or U1414 (N_1414,In_1130,In_210);
and U1415 (N_1415,In_740,In_420);
and U1416 (N_1416,In_811,In_1264);
and U1417 (N_1417,In_2384,In_89);
xnor U1418 (N_1418,In_108,In_2000);
nor U1419 (N_1419,In_1483,In_817);
nand U1420 (N_1420,In_1859,In_2286);
nor U1421 (N_1421,In_2319,In_1635);
or U1422 (N_1422,In_775,In_2025);
nand U1423 (N_1423,In_2425,In_1351);
or U1424 (N_1424,In_979,In_1025);
nand U1425 (N_1425,In_946,In_1577);
nand U1426 (N_1426,In_2444,In_1108);
nand U1427 (N_1427,In_869,In_173);
xnor U1428 (N_1428,In_2250,In_456);
and U1429 (N_1429,In_1161,In_37);
and U1430 (N_1430,In_1563,In_1772);
nand U1431 (N_1431,In_1587,In_186);
nor U1432 (N_1432,In_230,In_203);
nor U1433 (N_1433,In_1007,In_2398);
nor U1434 (N_1434,In_1448,In_2461);
xnor U1435 (N_1435,In_1752,In_1826);
xnor U1436 (N_1436,In_720,In_626);
and U1437 (N_1437,In_2173,In_2257);
xnor U1438 (N_1438,In_911,In_2200);
nor U1439 (N_1439,In_1909,In_853);
or U1440 (N_1440,In_2347,In_566);
nor U1441 (N_1441,In_291,In_924);
and U1442 (N_1442,In_368,In_738);
nand U1443 (N_1443,In_2026,In_1399);
and U1444 (N_1444,In_110,In_1619);
and U1445 (N_1445,In_1962,In_2192);
or U1446 (N_1446,In_1505,In_1537);
xor U1447 (N_1447,In_921,In_528);
nand U1448 (N_1448,In_1471,In_1792);
xor U1449 (N_1449,In_1577,In_888);
or U1450 (N_1450,In_1393,In_136);
nand U1451 (N_1451,In_2319,In_944);
nand U1452 (N_1452,In_835,In_1548);
nand U1453 (N_1453,In_847,In_2327);
and U1454 (N_1454,In_1341,In_376);
or U1455 (N_1455,In_1806,In_106);
nor U1456 (N_1456,In_753,In_520);
nand U1457 (N_1457,In_1370,In_135);
xnor U1458 (N_1458,In_148,In_646);
nor U1459 (N_1459,In_2153,In_2172);
nand U1460 (N_1460,In_106,In_1556);
and U1461 (N_1461,In_1787,In_1717);
and U1462 (N_1462,In_1158,In_927);
nor U1463 (N_1463,In_644,In_389);
nor U1464 (N_1464,In_211,In_1991);
xnor U1465 (N_1465,In_674,In_1025);
nor U1466 (N_1466,In_1945,In_2401);
and U1467 (N_1467,In_601,In_2287);
nand U1468 (N_1468,In_448,In_979);
and U1469 (N_1469,In_292,In_715);
xnor U1470 (N_1470,In_2344,In_814);
and U1471 (N_1471,In_445,In_43);
or U1472 (N_1472,In_760,In_1038);
and U1473 (N_1473,In_1299,In_1418);
and U1474 (N_1474,In_723,In_1903);
nor U1475 (N_1475,In_2407,In_582);
or U1476 (N_1476,In_437,In_533);
nor U1477 (N_1477,In_518,In_752);
nor U1478 (N_1478,In_1520,In_657);
or U1479 (N_1479,In_1692,In_1789);
nand U1480 (N_1480,In_2375,In_1496);
nand U1481 (N_1481,In_888,In_1273);
nand U1482 (N_1482,In_1240,In_1664);
or U1483 (N_1483,In_1354,In_42);
nor U1484 (N_1484,In_1299,In_1536);
nor U1485 (N_1485,In_1241,In_1366);
nand U1486 (N_1486,In_1599,In_2194);
nor U1487 (N_1487,In_1053,In_2027);
nor U1488 (N_1488,In_1919,In_2148);
nand U1489 (N_1489,In_2373,In_683);
nand U1490 (N_1490,In_221,In_1069);
or U1491 (N_1491,In_1874,In_120);
nand U1492 (N_1492,In_1288,In_489);
or U1493 (N_1493,In_1312,In_1477);
or U1494 (N_1494,In_905,In_2327);
and U1495 (N_1495,In_105,In_284);
and U1496 (N_1496,In_1732,In_2302);
nor U1497 (N_1497,In_1836,In_2);
nor U1498 (N_1498,In_2006,In_37);
nand U1499 (N_1499,In_387,In_2106);
nor U1500 (N_1500,In_1158,In_1076);
nand U1501 (N_1501,In_2001,In_1901);
nand U1502 (N_1502,In_890,In_449);
nor U1503 (N_1503,In_257,In_1785);
and U1504 (N_1504,In_2062,In_228);
or U1505 (N_1505,In_2290,In_2029);
and U1506 (N_1506,In_807,In_2478);
or U1507 (N_1507,In_1224,In_484);
and U1508 (N_1508,In_827,In_1800);
or U1509 (N_1509,In_378,In_802);
xor U1510 (N_1510,In_2199,In_1863);
nor U1511 (N_1511,In_2462,In_449);
and U1512 (N_1512,In_2471,In_2315);
nor U1513 (N_1513,In_498,In_14);
or U1514 (N_1514,In_1140,In_558);
nand U1515 (N_1515,In_1058,In_296);
nand U1516 (N_1516,In_845,In_250);
and U1517 (N_1517,In_1436,In_2429);
nand U1518 (N_1518,In_1472,In_655);
nand U1519 (N_1519,In_827,In_1633);
xor U1520 (N_1520,In_191,In_1407);
nand U1521 (N_1521,In_1810,In_1732);
nor U1522 (N_1522,In_2096,In_748);
nor U1523 (N_1523,In_1413,In_1672);
or U1524 (N_1524,In_2102,In_1067);
xor U1525 (N_1525,In_1322,In_808);
and U1526 (N_1526,In_1596,In_2379);
and U1527 (N_1527,In_240,In_574);
and U1528 (N_1528,In_1741,In_129);
and U1529 (N_1529,In_973,In_18);
or U1530 (N_1530,In_543,In_526);
nand U1531 (N_1531,In_468,In_1336);
and U1532 (N_1532,In_998,In_2256);
or U1533 (N_1533,In_1230,In_1587);
or U1534 (N_1534,In_1459,In_1880);
xor U1535 (N_1535,In_736,In_1633);
nor U1536 (N_1536,In_1981,In_2467);
xor U1537 (N_1537,In_858,In_1986);
and U1538 (N_1538,In_692,In_136);
or U1539 (N_1539,In_26,In_1914);
xor U1540 (N_1540,In_1917,In_1436);
nand U1541 (N_1541,In_146,In_735);
nand U1542 (N_1542,In_837,In_162);
or U1543 (N_1543,In_163,In_2137);
nor U1544 (N_1544,In_891,In_441);
nor U1545 (N_1545,In_1248,In_2402);
and U1546 (N_1546,In_2439,In_1234);
nand U1547 (N_1547,In_1088,In_1493);
nand U1548 (N_1548,In_2108,In_1989);
and U1549 (N_1549,In_2031,In_500);
nand U1550 (N_1550,In_612,In_1835);
nand U1551 (N_1551,In_801,In_2141);
nand U1552 (N_1552,In_1816,In_2095);
nand U1553 (N_1553,In_1962,In_44);
and U1554 (N_1554,In_78,In_2467);
and U1555 (N_1555,In_1750,In_2234);
and U1556 (N_1556,In_1469,In_1263);
or U1557 (N_1557,In_2053,In_1416);
nand U1558 (N_1558,In_310,In_781);
xnor U1559 (N_1559,In_888,In_347);
and U1560 (N_1560,In_83,In_2213);
nand U1561 (N_1561,In_1120,In_1365);
and U1562 (N_1562,In_485,In_1309);
nand U1563 (N_1563,In_183,In_1836);
or U1564 (N_1564,In_388,In_904);
or U1565 (N_1565,In_1434,In_779);
nand U1566 (N_1566,In_1406,In_1850);
nor U1567 (N_1567,In_533,In_416);
or U1568 (N_1568,In_985,In_975);
nand U1569 (N_1569,In_614,In_98);
nor U1570 (N_1570,In_222,In_2034);
and U1571 (N_1571,In_1407,In_2396);
nor U1572 (N_1572,In_755,In_194);
and U1573 (N_1573,In_399,In_431);
and U1574 (N_1574,In_963,In_646);
and U1575 (N_1575,In_1213,In_1083);
xnor U1576 (N_1576,In_449,In_755);
and U1577 (N_1577,In_1696,In_447);
nand U1578 (N_1578,In_2096,In_435);
and U1579 (N_1579,In_1095,In_788);
nand U1580 (N_1580,In_160,In_243);
nor U1581 (N_1581,In_2201,In_2184);
nor U1582 (N_1582,In_859,In_2216);
and U1583 (N_1583,In_763,In_1083);
or U1584 (N_1584,In_2049,In_1338);
xor U1585 (N_1585,In_2049,In_1160);
xnor U1586 (N_1586,In_963,In_2486);
nor U1587 (N_1587,In_93,In_1718);
or U1588 (N_1588,In_301,In_1903);
nand U1589 (N_1589,In_192,In_1486);
nor U1590 (N_1590,In_745,In_2211);
and U1591 (N_1591,In_290,In_132);
and U1592 (N_1592,In_366,In_2072);
xor U1593 (N_1593,In_396,In_31);
and U1594 (N_1594,In_1175,In_551);
nand U1595 (N_1595,In_1896,In_1957);
or U1596 (N_1596,In_1935,In_619);
and U1597 (N_1597,In_1012,In_508);
xor U1598 (N_1598,In_2237,In_1541);
and U1599 (N_1599,In_799,In_743);
nand U1600 (N_1600,In_253,In_523);
or U1601 (N_1601,In_1302,In_410);
and U1602 (N_1602,In_2069,In_1931);
nor U1603 (N_1603,In_2291,In_1620);
nor U1604 (N_1604,In_927,In_967);
xor U1605 (N_1605,In_1504,In_415);
or U1606 (N_1606,In_407,In_686);
nand U1607 (N_1607,In_1103,In_1912);
and U1608 (N_1608,In_1020,In_644);
and U1609 (N_1609,In_2481,In_2369);
nor U1610 (N_1610,In_740,In_2254);
or U1611 (N_1611,In_1689,In_2380);
or U1612 (N_1612,In_2437,In_832);
nand U1613 (N_1613,In_2132,In_2024);
and U1614 (N_1614,In_456,In_1124);
and U1615 (N_1615,In_1436,In_260);
nand U1616 (N_1616,In_375,In_1505);
xor U1617 (N_1617,In_1258,In_2384);
and U1618 (N_1618,In_2282,In_524);
nor U1619 (N_1619,In_1418,In_2374);
nand U1620 (N_1620,In_80,In_1473);
and U1621 (N_1621,In_1361,In_2399);
or U1622 (N_1622,In_1949,In_557);
nor U1623 (N_1623,In_1691,In_1156);
nor U1624 (N_1624,In_920,In_1004);
nor U1625 (N_1625,In_1970,In_765);
and U1626 (N_1626,In_54,In_1604);
and U1627 (N_1627,In_795,In_72);
or U1628 (N_1628,In_570,In_1646);
xnor U1629 (N_1629,In_602,In_2018);
or U1630 (N_1630,In_2218,In_1376);
or U1631 (N_1631,In_1777,In_1337);
or U1632 (N_1632,In_1413,In_2086);
and U1633 (N_1633,In_1749,In_2200);
nand U1634 (N_1634,In_2055,In_183);
nor U1635 (N_1635,In_1123,In_1988);
xnor U1636 (N_1636,In_1075,In_1747);
or U1637 (N_1637,In_709,In_1240);
nand U1638 (N_1638,In_1247,In_746);
nor U1639 (N_1639,In_2360,In_2402);
nor U1640 (N_1640,In_2104,In_450);
or U1641 (N_1641,In_349,In_1712);
nand U1642 (N_1642,In_1403,In_1221);
or U1643 (N_1643,In_313,In_1290);
nand U1644 (N_1644,In_1503,In_1283);
or U1645 (N_1645,In_854,In_1055);
or U1646 (N_1646,In_1939,In_537);
nor U1647 (N_1647,In_573,In_2399);
nor U1648 (N_1648,In_1186,In_1765);
nor U1649 (N_1649,In_696,In_802);
and U1650 (N_1650,In_1970,In_521);
nand U1651 (N_1651,In_516,In_1158);
and U1652 (N_1652,In_2008,In_1364);
or U1653 (N_1653,In_2304,In_2391);
or U1654 (N_1654,In_366,In_1281);
nor U1655 (N_1655,In_2120,In_460);
nor U1656 (N_1656,In_1376,In_885);
or U1657 (N_1657,In_1548,In_670);
and U1658 (N_1658,In_1463,In_356);
and U1659 (N_1659,In_998,In_2481);
or U1660 (N_1660,In_2244,In_994);
or U1661 (N_1661,In_1883,In_372);
and U1662 (N_1662,In_1664,In_2420);
and U1663 (N_1663,In_504,In_2411);
xor U1664 (N_1664,In_670,In_880);
nand U1665 (N_1665,In_2462,In_1635);
nor U1666 (N_1666,In_1637,In_1890);
nor U1667 (N_1667,In_1712,In_601);
and U1668 (N_1668,In_1864,In_203);
nand U1669 (N_1669,In_323,In_1543);
nor U1670 (N_1670,In_1868,In_1466);
nand U1671 (N_1671,In_2039,In_795);
nor U1672 (N_1672,In_2346,In_466);
nand U1673 (N_1673,In_2138,In_1110);
xor U1674 (N_1674,In_1268,In_255);
and U1675 (N_1675,In_335,In_1568);
and U1676 (N_1676,In_511,In_1954);
or U1677 (N_1677,In_2239,In_467);
and U1678 (N_1678,In_1890,In_995);
nand U1679 (N_1679,In_1269,In_1688);
nand U1680 (N_1680,In_662,In_2035);
xnor U1681 (N_1681,In_1177,In_1092);
xnor U1682 (N_1682,In_191,In_1003);
nand U1683 (N_1683,In_2007,In_769);
nand U1684 (N_1684,In_1802,In_402);
nor U1685 (N_1685,In_2018,In_1934);
xor U1686 (N_1686,In_2410,In_898);
nor U1687 (N_1687,In_592,In_1763);
nor U1688 (N_1688,In_2408,In_1915);
nor U1689 (N_1689,In_2479,In_1661);
nand U1690 (N_1690,In_721,In_2066);
xor U1691 (N_1691,In_1375,In_419);
and U1692 (N_1692,In_870,In_1170);
and U1693 (N_1693,In_719,In_1403);
nor U1694 (N_1694,In_543,In_1397);
nor U1695 (N_1695,In_4,In_983);
and U1696 (N_1696,In_2038,In_790);
and U1697 (N_1697,In_1850,In_411);
nor U1698 (N_1698,In_2107,In_634);
nand U1699 (N_1699,In_130,In_1427);
nand U1700 (N_1700,In_1644,In_1670);
xor U1701 (N_1701,In_1066,In_1205);
or U1702 (N_1702,In_866,In_926);
or U1703 (N_1703,In_1563,In_2484);
nor U1704 (N_1704,In_2177,In_117);
xnor U1705 (N_1705,In_2180,In_422);
nand U1706 (N_1706,In_1618,In_316);
nor U1707 (N_1707,In_893,In_1195);
or U1708 (N_1708,In_938,In_2129);
and U1709 (N_1709,In_1368,In_1740);
nand U1710 (N_1710,In_1740,In_1658);
xnor U1711 (N_1711,In_857,In_361);
nand U1712 (N_1712,In_1652,In_2351);
or U1713 (N_1713,In_174,In_25);
nor U1714 (N_1714,In_200,In_141);
xor U1715 (N_1715,In_2368,In_1076);
nand U1716 (N_1716,In_781,In_1533);
and U1717 (N_1717,In_2098,In_414);
nand U1718 (N_1718,In_1122,In_2157);
nand U1719 (N_1719,In_1382,In_1756);
and U1720 (N_1720,In_2369,In_566);
nor U1721 (N_1721,In_390,In_1660);
nand U1722 (N_1722,In_2007,In_1525);
nand U1723 (N_1723,In_1271,In_806);
and U1724 (N_1724,In_1316,In_1870);
nand U1725 (N_1725,In_916,In_1260);
and U1726 (N_1726,In_2410,In_126);
nand U1727 (N_1727,In_827,In_346);
nand U1728 (N_1728,In_2135,In_2086);
or U1729 (N_1729,In_8,In_565);
or U1730 (N_1730,In_2388,In_2406);
nor U1731 (N_1731,In_2083,In_515);
xor U1732 (N_1732,In_1297,In_1823);
nand U1733 (N_1733,In_636,In_1119);
nand U1734 (N_1734,In_1,In_1672);
nand U1735 (N_1735,In_2100,In_444);
nor U1736 (N_1736,In_1356,In_396);
or U1737 (N_1737,In_2489,In_2285);
or U1738 (N_1738,In_1370,In_632);
or U1739 (N_1739,In_1284,In_2169);
and U1740 (N_1740,In_1560,In_1449);
nor U1741 (N_1741,In_890,In_405);
xnor U1742 (N_1742,In_25,In_1036);
and U1743 (N_1743,In_733,In_1820);
nand U1744 (N_1744,In_1,In_843);
nand U1745 (N_1745,In_1222,In_117);
nand U1746 (N_1746,In_869,In_499);
nand U1747 (N_1747,In_44,In_1856);
nand U1748 (N_1748,In_238,In_2107);
nor U1749 (N_1749,In_2240,In_1290);
xnor U1750 (N_1750,In_511,In_184);
xnor U1751 (N_1751,In_612,In_2320);
or U1752 (N_1752,In_988,In_253);
nand U1753 (N_1753,In_1490,In_2246);
nand U1754 (N_1754,In_2206,In_2225);
and U1755 (N_1755,In_818,In_696);
nand U1756 (N_1756,In_1315,In_2014);
nor U1757 (N_1757,In_1427,In_533);
nand U1758 (N_1758,In_239,In_2138);
nor U1759 (N_1759,In_1235,In_350);
nand U1760 (N_1760,In_1410,In_579);
nor U1761 (N_1761,In_1939,In_612);
or U1762 (N_1762,In_2483,In_1638);
nand U1763 (N_1763,In_1588,In_1607);
xnor U1764 (N_1764,In_2217,In_2001);
nor U1765 (N_1765,In_911,In_348);
and U1766 (N_1766,In_217,In_2041);
or U1767 (N_1767,In_282,In_2061);
nor U1768 (N_1768,In_569,In_2370);
or U1769 (N_1769,In_654,In_1074);
nand U1770 (N_1770,In_2244,In_1815);
nor U1771 (N_1771,In_48,In_310);
and U1772 (N_1772,In_1304,In_1002);
and U1773 (N_1773,In_797,In_1515);
or U1774 (N_1774,In_2125,In_723);
nor U1775 (N_1775,In_889,In_734);
or U1776 (N_1776,In_2441,In_2309);
and U1777 (N_1777,In_1834,In_1350);
nor U1778 (N_1778,In_1112,In_1820);
nor U1779 (N_1779,In_1372,In_2071);
and U1780 (N_1780,In_1905,In_1425);
and U1781 (N_1781,In_2196,In_1733);
and U1782 (N_1782,In_376,In_679);
nand U1783 (N_1783,In_2023,In_1084);
nand U1784 (N_1784,In_45,In_448);
nor U1785 (N_1785,In_1047,In_428);
nand U1786 (N_1786,In_1046,In_712);
or U1787 (N_1787,In_1901,In_69);
and U1788 (N_1788,In_1016,In_929);
nor U1789 (N_1789,In_987,In_749);
nor U1790 (N_1790,In_1092,In_1002);
nor U1791 (N_1791,In_1119,In_908);
and U1792 (N_1792,In_1003,In_1267);
nor U1793 (N_1793,In_1135,In_301);
and U1794 (N_1794,In_113,In_2088);
nor U1795 (N_1795,In_9,In_2220);
and U1796 (N_1796,In_1133,In_2197);
nor U1797 (N_1797,In_1604,In_1730);
or U1798 (N_1798,In_1108,In_1061);
nor U1799 (N_1799,In_2175,In_1454);
nand U1800 (N_1800,In_2239,In_420);
nor U1801 (N_1801,In_1421,In_259);
or U1802 (N_1802,In_17,In_140);
xnor U1803 (N_1803,In_1803,In_1904);
nor U1804 (N_1804,In_1262,In_1796);
nand U1805 (N_1805,In_568,In_493);
and U1806 (N_1806,In_1882,In_701);
nor U1807 (N_1807,In_1927,In_2462);
or U1808 (N_1808,In_1747,In_652);
xnor U1809 (N_1809,In_194,In_589);
nand U1810 (N_1810,In_1962,In_573);
nand U1811 (N_1811,In_1254,In_876);
or U1812 (N_1812,In_2270,In_1862);
and U1813 (N_1813,In_2467,In_2303);
and U1814 (N_1814,In_2221,In_376);
and U1815 (N_1815,In_501,In_991);
or U1816 (N_1816,In_1105,In_350);
nand U1817 (N_1817,In_1578,In_1777);
nor U1818 (N_1818,In_541,In_439);
or U1819 (N_1819,In_143,In_2047);
nor U1820 (N_1820,In_1655,In_1063);
nor U1821 (N_1821,In_123,In_2087);
or U1822 (N_1822,In_1907,In_2359);
and U1823 (N_1823,In_372,In_194);
nor U1824 (N_1824,In_194,In_1577);
nor U1825 (N_1825,In_1909,In_1860);
and U1826 (N_1826,In_1681,In_1247);
and U1827 (N_1827,In_312,In_439);
and U1828 (N_1828,In_2010,In_1461);
nand U1829 (N_1829,In_2321,In_1251);
xor U1830 (N_1830,In_929,In_2123);
nand U1831 (N_1831,In_120,In_525);
xor U1832 (N_1832,In_254,In_1980);
or U1833 (N_1833,In_626,In_1932);
nand U1834 (N_1834,In_1095,In_1805);
nand U1835 (N_1835,In_1295,In_301);
nor U1836 (N_1836,In_763,In_1901);
nor U1837 (N_1837,In_1431,In_1079);
xor U1838 (N_1838,In_1701,In_2239);
nand U1839 (N_1839,In_2333,In_1271);
xor U1840 (N_1840,In_1099,In_653);
nor U1841 (N_1841,In_1561,In_1302);
and U1842 (N_1842,In_1726,In_542);
or U1843 (N_1843,In_1870,In_1830);
nand U1844 (N_1844,In_2490,In_304);
and U1845 (N_1845,In_2235,In_1396);
nand U1846 (N_1846,In_1277,In_1427);
nand U1847 (N_1847,In_1469,In_381);
and U1848 (N_1848,In_353,In_2242);
nand U1849 (N_1849,In_1880,In_77);
xnor U1850 (N_1850,In_2145,In_1559);
nand U1851 (N_1851,In_1114,In_435);
nor U1852 (N_1852,In_2383,In_1635);
nand U1853 (N_1853,In_1178,In_2090);
or U1854 (N_1854,In_1786,In_396);
and U1855 (N_1855,In_1932,In_2329);
and U1856 (N_1856,In_925,In_997);
nor U1857 (N_1857,In_1076,In_2405);
nand U1858 (N_1858,In_435,In_426);
nor U1859 (N_1859,In_1716,In_2209);
nand U1860 (N_1860,In_1788,In_725);
nand U1861 (N_1861,In_2277,In_1338);
nand U1862 (N_1862,In_101,In_2025);
or U1863 (N_1863,In_531,In_2100);
and U1864 (N_1864,In_834,In_1037);
xnor U1865 (N_1865,In_391,In_932);
or U1866 (N_1866,In_157,In_1224);
nor U1867 (N_1867,In_1529,In_2464);
nand U1868 (N_1868,In_86,In_1312);
or U1869 (N_1869,In_423,In_382);
and U1870 (N_1870,In_1090,In_1086);
nand U1871 (N_1871,In_1361,In_1938);
nor U1872 (N_1872,In_1252,In_613);
nand U1873 (N_1873,In_1465,In_1862);
nor U1874 (N_1874,In_1926,In_2288);
nor U1875 (N_1875,In_1778,In_249);
and U1876 (N_1876,In_307,In_143);
nand U1877 (N_1877,In_2496,In_211);
and U1878 (N_1878,In_2334,In_2127);
xnor U1879 (N_1879,In_1801,In_2189);
or U1880 (N_1880,In_275,In_648);
and U1881 (N_1881,In_1882,In_1588);
or U1882 (N_1882,In_343,In_1857);
xor U1883 (N_1883,In_1264,In_853);
and U1884 (N_1884,In_1136,In_518);
xor U1885 (N_1885,In_2342,In_978);
or U1886 (N_1886,In_2241,In_883);
nand U1887 (N_1887,In_2483,In_1105);
and U1888 (N_1888,In_1447,In_2470);
xor U1889 (N_1889,In_1057,In_1717);
nand U1890 (N_1890,In_1494,In_1539);
or U1891 (N_1891,In_1954,In_2088);
nand U1892 (N_1892,In_1629,In_1467);
nand U1893 (N_1893,In_959,In_2393);
and U1894 (N_1894,In_2150,In_254);
and U1895 (N_1895,In_55,In_530);
nand U1896 (N_1896,In_1215,In_1921);
or U1897 (N_1897,In_1541,In_455);
or U1898 (N_1898,In_335,In_1649);
nor U1899 (N_1899,In_703,In_610);
and U1900 (N_1900,In_2332,In_523);
and U1901 (N_1901,In_1695,In_1001);
or U1902 (N_1902,In_244,In_2094);
or U1903 (N_1903,In_88,In_1112);
and U1904 (N_1904,In_2493,In_1995);
or U1905 (N_1905,In_1483,In_334);
nand U1906 (N_1906,In_329,In_2272);
nand U1907 (N_1907,In_1126,In_241);
or U1908 (N_1908,In_274,In_2209);
nand U1909 (N_1909,In_1025,In_684);
xor U1910 (N_1910,In_2366,In_1003);
and U1911 (N_1911,In_1142,In_1052);
or U1912 (N_1912,In_1993,In_2008);
nand U1913 (N_1913,In_933,In_864);
nand U1914 (N_1914,In_2031,In_1049);
nor U1915 (N_1915,In_572,In_1186);
and U1916 (N_1916,In_1433,In_1531);
and U1917 (N_1917,In_726,In_1596);
and U1918 (N_1918,In_1133,In_1041);
and U1919 (N_1919,In_1954,In_605);
or U1920 (N_1920,In_599,In_2062);
and U1921 (N_1921,In_1605,In_1478);
nor U1922 (N_1922,In_1070,In_2320);
nand U1923 (N_1923,In_1948,In_633);
nor U1924 (N_1924,In_1139,In_1928);
and U1925 (N_1925,In_1733,In_2042);
xnor U1926 (N_1926,In_1424,In_1601);
nand U1927 (N_1927,In_924,In_1751);
xnor U1928 (N_1928,In_1338,In_118);
or U1929 (N_1929,In_1167,In_2003);
nor U1930 (N_1930,In_1121,In_782);
nor U1931 (N_1931,In_1862,In_2103);
nor U1932 (N_1932,In_896,In_155);
or U1933 (N_1933,In_892,In_661);
nor U1934 (N_1934,In_1395,In_881);
nor U1935 (N_1935,In_2396,In_1726);
xnor U1936 (N_1936,In_2299,In_652);
nor U1937 (N_1937,In_382,In_2385);
nand U1938 (N_1938,In_795,In_364);
nor U1939 (N_1939,In_2243,In_1711);
and U1940 (N_1940,In_1327,In_168);
or U1941 (N_1941,In_1838,In_1962);
xnor U1942 (N_1942,In_2050,In_822);
and U1943 (N_1943,In_325,In_1756);
and U1944 (N_1944,In_840,In_1721);
or U1945 (N_1945,In_2441,In_132);
and U1946 (N_1946,In_676,In_2276);
and U1947 (N_1947,In_1243,In_1889);
nor U1948 (N_1948,In_1352,In_1579);
xnor U1949 (N_1949,In_1755,In_118);
and U1950 (N_1950,In_2391,In_2009);
nor U1951 (N_1951,In_1526,In_1135);
and U1952 (N_1952,In_17,In_161);
and U1953 (N_1953,In_1463,In_1312);
nor U1954 (N_1954,In_1879,In_2114);
nor U1955 (N_1955,In_974,In_1913);
or U1956 (N_1956,In_1875,In_830);
nor U1957 (N_1957,In_1956,In_2220);
and U1958 (N_1958,In_2011,In_2136);
nor U1959 (N_1959,In_138,In_2086);
nand U1960 (N_1960,In_2400,In_216);
or U1961 (N_1961,In_1789,In_2236);
nor U1962 (N_1962,In_1771,In_2401);
and U1963 (N_1963,In_1432,In_404);
and U1964 (N_1964,In_1416,In_1721);
nor U1965 (N_1965,In_1314,In_1801);
nand U1966 (N_1966,In_1470,In_1762);
xnor U1967 (N_1967,In_2206,In_2253);
nand U1968 (N_1968,In_736,In_1890);
and U1969 (N_1969,In_1105,In_774);
or U1970 (N_1970,In_51,In_2029);
or U1971 (N_1971,In_1200,In_1523);
nor U1972 (N_1972,In_631,In_1140);
nor U1973 (N_1973,In_636,In_147);
and U1974 (N_1974,In_96,In_1028);
and U1975 (N_1975,In_34,In_1440);
and U1976 (N_1976,In_174,In_1952);
and U1977 (N_1977,In_2094,In_1525);
or U1978 (N_1978,In_1833,In_846);
nand U1979 (N_1979,In_527,In_1738);
and U1980 (N_1980,In_163,In_959);
nand U1981 (N_1981,In_1482,In_343);
or U1982 (N_1982,In_835,In_1913);
nor U1983 (N_1983,In_1544,In_1664);
nor U1984 (N_1984,In_876,In_1545);
nor U1985 (N_1985,In_1924,In_558);
and U1986 (N_1986,In_550,In_967);
and U1987 (N_1987,In_185,In_752);
nand U1988 (N_1988,In_1386,In_2020);
nand U1989 (N_1989,In_767,In_1700);
and U1990 (N_1990,In_2143,In_2346);
nand U1991 (N_1991,In_1431,In_382);
nand U1992 (N_1992,In_890,In_91);
nand U1993 (N_1993,In_406,In_2437);
nor U1994 (N_1994,In_1358,In_754);
nor U1995 (N_1995,In_1789,In_467);
nand U1996 (N_1996,In_125,In_2271);
nor U1997 (N_1997,In_2028,In_1872);
nand U1998 (N_1998,In_1149,In_2136);
or U1999 (N_1999,In_912,In_383);
and U2000 (N_2000,In_411,In_1701);
and U2001 (N_2001,In_1105,In_1289);
nand U2002 (N_2002,In_1536,In_2283);
and U2003 (N_2003,In_1373,In_2060);
or U2004 (N_2004,In_1643,In_1986);
and U2005 (N_2005,In_1633,In_777);
nand U2006 (N_2006,In_1836,In_1882);
or U2007 (N_2007,In_1823,In_1397);
or U2008 (N_2008,In_2104,In_2178);
nand U2009 (N_2009,In_1362,In_858);
and U2010 (N_2010,In_1341,In_2226);
nand U2011 (N_2011,In_2410,In_1069);
and U2012 (N_2012,In_757,In_137);
or U2013 (N_2013,In_1557,In_680);
or U2014 (N_2014,In_1488,In_595);
nand U2015 (N_2015,In_1876,In_380);
nand U2016 (N_2016,In_1751,In_1516);
nor U2017 (N_2017,In_305,In_1257);
nand U2018 (N_2018,In_569,In_926);
and U2019 (N_2019,In_887,In_2018);
or U2020 (N_2020,In_1647,In_288);
xor U2021 (N_2021,In_1541,In_1666);
nor U2022 (N_2022,In_1078,In_95);
nand U2023 (N_2023,In_2122,In_2316);
or U2024 (N_2024,In_920,In_1435);
nand U2025 (N_2025,In_1849,In_1487);
and U2026 (N_2026,In_2194,In_2011);
nor U2027 (N_2027,In_946,In_641);
nand U2028 (N_2028,In_1534,In_580);
or U2029 (N_2029,In_2091,In_1905);
or U2030 (N_2030,In_838,In_800);
nor U2031 (N_2031,In_1496,In_5);
or U2032 (N_2032,In_981,In_192);
and U2033 (N_2033,In_296,In_1001);
xnor U2034 (N_2034,In_2096,In_145);
xnor U2035 (N_2035,In_1679,In_1837);
or U2036 (N_2036,In_2414,In_1123);
and U2037 (N_2037,In_232,In_1887);
nand U2038 (N_2038,In_1502,In_218);
or U2039 (N_2039,In_77,In_1038);
nand U2040 (N_2040,In_110,In_1457);
nor U2041 (N_2041,In_1603,In_857);
nand U2042 (N_2042,In_1747,In_8);
and U2043 (N_2043,In_317,In_2495);
xnor U2044 (N_2044,In_281,In_1565);
and U2045 (N_2045,In_1607,In_527);
nor U2046 (N_2046,In_1795,In_2434);
or U2047 (N_2047,In_1885,In_1786);
or U2048 (N_2048,In_1368,In_1545);
or U2049 (N_2049,In_344,In_2161);
nand U2050 (N_2050,In_305,In_1420);
and U2051 (N_2051,In_81,In_1635);
and U2052 (N_2052,In_1600,In_2169);
or U2053 (N_2053,In_696,In_224);
and U2054 (N_2054,In_184,In_832);
nor U2055 (N_2055,In_365,In_1007);
and U2056 (N_2056,In_1972,In_1449);
nor U2057 (N_2057,In_1297,In_964);
and U2058 (N_2058,In_184,In_166);
and U2059 (N_2059,In_824,In_387);
nand U2060 (N_2060,In_567,In_1494);
nand U2061 (N_2061,In_2205,In_2387);
or U2062 (N_2062,In_1371,In_1299);
and U2063 (N_2063,In_1794,In_1488);
nor U2064 (N_2064,In_2046,In_2431);
nand U2065 (N_2065,In_801,In_1302);
nor U2066 (N_2066,In_244,In_2434);
and U2067 (N_2067,In_1134,In_1970);
or U2068 (N_2068,In_280,In_1846);
or U2069 (N_2069,In_1835,In_453);
nand U2070 (N_2070,In_1610,In_258);
and U2071 (N_2071,In_31,In_2165);
and U2072 (N_2072,In_1109,In_1104);
and U2073 (N_2073,In_949,In_1608);
and U2074 (N_2074,In_1383,In_2063);
nor U2075 (N_2075,In_1481,In_1791);
and U2076 (N_2076,In_1679,In_934);
nand U2077 (N_2077,In_1023,In_2349);
and U2078 (N_2078,In_1539,In_483);
and U2079 (N_2079,In_878,In_1220);
nand U2080 (N_2080,In_242,In_1230);
and U2081 (N_2081,In_507,In_1817);
nand U2082 (N_2082,In_1522,In_257);
nor U2083 (N_2083,In_5,In_1889);
or U2084 (N_2084,In_385,In_1521);
and U2085 (N_2085,In_1936,In_1946);
xor U2086 (N_2086,In_140,In_861);
and U2087 (N_2087,In_1526,In_898);
nor U2088 (N_2088,In_1585,In_601);
nor U2089 (N_2089,In_1506,In_1414);
nor U2090 (N_2090,In_1964,In_1413);
or U2091 (N_2091,In_1149,In_146);
nand U2092 (N_2092,In_1164,In_1484);
and U2093 (N_2093,In_1258,In_2106);
and U2094 (N_2094,In_1954,In_779);
xnor U2095 (N_2095,In_2490,In_548);
nand U2096 (N_2096,In_1248,In_70);
nor U2097 (N_2097,In_2007,In_835);
or U2098 (N_2098,In_245,In_1623);
or U2099 (N_2099,In_1865,In_1650);
or U2100 (N_2100,In_1550,In_1631);
and U2101 (N_2101,In_214,In_1645);
and U2102 (N_2102,In_923,In_1447);
nor U2103 (N_2103,In_130,In_839);
nand U2104 (N_2104,In_33,In_1992);
nor U2105 (N_2105,In_2386,In_2025);
nand U2106 (N_2106,In_1052,In_136);
xnor U2107 (N_2107,In_2043,In_878);
or U2108 (N_2108,In_732,In_503);
or U2109 (N_2109,In_1632,In_1285);
nand U2110 (N_2110,In_1713,In_2118);
xor U2111 (N_2111,In_276,In_23);
nand U2112 (N_2112,In_1791,In_2402);
and U2113 (N_2113,In_412,In_2053);
nand U2114 (N_2114,In_2353,In_2378);
nand U2115 (N_2115,In_2139,In_1828);
or U2116 (N_2116,In_188,In_645);
and U2117 (N_2117,In_2005,In_2122);
nand U2118 (N_2118,In_1972,In_993);
and U2119 (N_2119,In_1809,In_1210);
nand U2120 (N_2120,In_299,In_1654);
nor U2121 (N_2121,In_2150,In_1234);
nand U2122 (N_2122,In_786,In_2325);
nand U2123 (N_2123,In_29,In_997);
or U2124 (N_2124,In_561,In_495);
nor U2125 (N_2125,In_2258,In_621);
and U2126 (N_2126,In_1651,In_2005);
and U2127 (N_2127,In_451,In_2495);
nor U2128 (N_2128,In_381,In_872);
nand U2129 (N_2129,In_1766,In_1745);
or U2130 (N_2130,In_1385,In_2088);
nand U2131 (N_2131,In_229,In_1053);
nor U2132 (N_2132,In_166,In_2339);
xor U2133 (N_2133,In_1558,In_267);
nor U2134 (N_2134,In_2416,In_1585);
nor U2135 (N_2135,In_945,In_2364);
nand U2136 (N_2136,In_2332,In_1251);
or U2137 (N_2137,In_1542,In_2228);
or U2138 (N_2138,In_691,In_670);
nor U2139 (N_2139,In_87,In_2418);
and U2140 (N_2140,In_299,In_2442);
and U2141 (N_2141,In_383,In_1220);
nand U2142 (N_2142,In_1941,In_173);
nor U2143 (N_2143,In_444,In_2249);
or U2144 (N_2144,In_12,In_1149);
nand U2145 (N_2145,In_2035,In_1232);
and U2146 (N_2146,In_2153,In_1174);
or U2147 (N_2147,In_1368,In_1748);
or U2148 (N_2148,In_1101,In_1163);
and U2149 (N_2149,In_105,In_1307);
or U2150 (N_2150,In_2493,In_2047);
or U2151 (N_2151,In_237,In_72);
nor U2152 (N_2152,In_1889,In_2436);
or U2153 (N_2153,In_1650,In_1205);
nand U2154 (N_2154,In_2315,In_1333);
nand U2155 (N_2155,In_1217,In_1493);
and U2156 (N_2156,In_823,In_1145);
and U2157 (N_2157,In_570,In_500);
and U2158 (N_2158,In_2474,In_162);
nor U2159 (N_2159,In_101,In_2080);
nor U2160 (N_2160,In_2139,In_2121);
and U2161 (N_2161,In_2325,In_263);
nand U2162 (N_2162,In_1868,In_808);
or U2163 (N_2163,In_1397,In_1000);
nand U2164 (N_2164,In_2418,In_1356);
and U2165 (N_2165,In_2438,In_320);
and U2166 (N_2166,In_656,In_793);
nor U2167 (N_2167,In_1050,In_2169);
or U2168 (N_2168,In_373,In_1236);
and U2169 (N_2169,In_2292,In_1771);
or U2170 (N_2170,In_2188,In_2168);
xnor U2171 (N_2171,In_101,In_852);
nor U2172 (N_2172,In_942,In_392);
nand U2173 (N_2173,In_415,In_558);
and U2174 (N_2174,In_1521,In_1143);
or U2175 (N_2175,In_2262,In_1725);
nand U2176 (N_2176,In_333,In_450);
nand U2177 (N_2177,In_1829,In_645);
nand U2178 (N_2178,In_7,In_1199);
and U2179 (N_2179,In_2417,In_503);
and U2180 (N_2180,In_1749,In_1476);
and U2181 (N_2181,In_780,In_1304);
and U2182 (N_2182,In_1688,In_2185);
nand U2183 (N_2183,In_1139,In_1681);
and U2184 (N_2184,In_684,In_110);
xor U2185 (N_2185,In_1852,In_972);
nor U2186 (N_2186,In_978,In_1824);
or U2187 (N_2187,In_663,In_1547);
nor U2188 (N_2188,In_348,In_2254);
nor U2189 (N_2189,In_2328,In_1860);
nor U2190 (N_2190,In_925,In_1550);
and U2191 (N_2191,In_2123,In_1773);
or U2192 (N_2192,In_1426,In_1345);
or U2193 (N_2193,In_560,In_1130);
xor U2194 (N_2194,In_1994,In_2336);
xor U2195 (N_2195,In_230,In_1109);
and U2196 (N_2196,In_1661,In_733);
or U2197 (N_2197,In_285,In_189);
or U2198 (N_2198,In_130,In_1796);
nor U2199 (N_2199,In_720,In_136);
and U2200 (N_2200,In_2443,In_943);
and U2201 (N_2201,In_580,In_1332);
or U2202 (N_2202,In_856,In_909);
nor U2203 (N_2203,In_965,In_730);
nand U2204 (N_2204,In_130,In_1269);
and U2205 (N_2205,In_1581,In_1434);
and U2206 (N_2206,In_538,In_2011);
nor U2207 (N_2207,In_2468,In_2186);
or U2208 (N_2208,In_1415,In_2112);
and U2209 (N_2209,In_1327,In_1747);
and U2210 (N_2210,In_1507,In_1116);
nor U2211 (N_2211,In_840,In_2199);
nor U2212 (N_2212,In_2184,In_2175);
or U2213 (N_2213,In_1657,In_31);
xnor U2214 (N_2214,In_964,In_722);
nand U2215 (N_2215,In_1467,In_2383);
nor U2216 (N_2216,In_1395,In_993);
and U2217 (N_2217,In_1118,In_2143);
nor U2218 (N_2218,In_2087,In_1507);
nor U2219 (N_2219,In_2107,In_1116);
nand U2220 (N_2220,In_1549,In_1199);
and U2221 (N_2221,In_2044,In_2485);
nor U2222 (N_2222,In_424,In_206);
or U2223 (N_2223,In_662,In_793);
or U2224 (N_2224,In_497,In_1562);
and U2225 (N_2225,In_1614,In_938);
nand U2226 (N_2226,In_1439,In_90);
and U2227 (N_2227,In_353,In_1251);
nand U2228 (N_2228,In_1406,In_1158);
and U2229 (N_2229,In_1333,In_996);
nand U2230 (N_2230,In_1468,In_719);
nor U2231 (N_2231,In_729,In_1131);
or U2232 (N_2232,In_180,In_778);
and U2233 (N_2233,In_1221,In_1607);
or U2234 (N_2234,In_2431,In_710);
and U2235 (N_2235,In_1499,In_1823);
xor U2236 (N_2236,In_1153,In_389);
and U2237 (N_2237,In_1328,In_1271);
and U2238 (N_2238,In_2283,In_192);
nand U2239 (N_2239,In_2434,In_939);
nor U2240 (N_2240,In_1306,In_660);
nor U2241 (N_2241,In_2292,In_585);
nand U2242 (N_2242,In_1866,In_367);
or U2243 (N_2243,In_479,In_725);
nand U2244 (N_2244,In_535,In_1131);
nor U2245 (N_2245,In_704,In_2001);
xnor U2246 (N_2246,In_2224,In_25);
or U2247 (N_2247,In_541,In_837);
and U2248 (N_2248,In_146,In_1549);
nand U2249 (N_2249,In_1954,In_1216);
nor U2250 (N_2250,In_659,In_1577);
nor U2251 (N_2251,In_1088,In_1026);
nand U2252 (N_2252,In_987,In_1960);
nor U2253 (N_2253,In_16,In_1138);
or U2254 (N_2254,In_2481,In_1168);
or U2255 (N_2255,In_290,In_239);
nor U2256 (N_2256,In_963,In_1795);
nor U2257 (N_2257,In_515,In_1507);
xor U2258 (N_2258,In_2349,In_839);
and U2259 (N_2259,In_374,In_2187);
and U2260 (N_2260,In_1661,In_209);
nand U2261 (N_2261,In_2472,In_2006);
and U2262 (N_2262,In_23,In_1264);
or U2263 (N_2263,In_2214,In_693);
or U2264 (N_2264,In_113,In_1293);
xnor U2265 (N_2265,In_190,In_983);
nand U2266 (N_2266,In_1831,In_494);
nor U2267 (N_2267,In_1717,In_51);
nor U2268 (N_2268,In_1929,In_1143);
and U2269 (N_2269,In_2091,In_1583);
nor U2270 (N_2270,In_75,In_2423);
and U2271 (N_2271,In_2135,In_1843);
nand U2272 (N_2272,In_2073,In_529);
and U2273 (N_2273,In_569,In_1434);
and U2274 (N_2274,In_791,In_1667);
and U2275 (N_2275,In_1616,In_1378);
and U2276 (N_2276,In_2151,In_1435);
nor U2277 (N_2277,In_1761,In_2460);
nor U2278 (N_2278,In_769,In_1599);
nand U2279 (N_2279,In_667,In_190);
nor U2280 (N_2280,In_1524,In_1925);
nor U2281 (N_2281,In_2061,In_1497);
xor U2282 (N_2282,In_657,In_1962);
or U2283 (N_2283,In_702,In_589);
nand U2284 (N_2284,In_2238,In_555);
nand U2285 (N_2285,In_877,In_153);
nor U2286 (N_2286,In_1076,In_800);
or U2287 (N_2287,In_1550,In_1947);
nor U2288 (N_2288,In_1060,In_780);
or U2289 (N_2289,In_2183,In_1348);
and U2290 (N_2290,In_405,In_1943);
and U2291 (N_2291,In_1040,In_2368);
and U2292 (N_2292,In_271,In_2393);
and U2293 (N_2293,In_1733,In_2396);
and U2294 (N_2294,In_1992,In_2370);
xnor U2295 (N_2295,In_1973,In_1280);
and U2296 (N_2296,In_582,In_1661);
xor U2297 (N_2297,In_54,In_1003);
and U2298 (N_2298,In_236,In_1695);
or U2299 (N_2299,In_1292,In_2077);
nor U2300 (N_2300,In_2254,In_1174);
or U2301 (N_2301,In_1642,In_2174);
and U2302 (N_2302,In_2480,In_1572);
nor U2303 (N_2303,In_1390,In_363);
and U2304 (N_2304,In_760,In_2017);
or U2305 (N_2305,In_1122,In_115);
nor U2306 (N_2306,In_676,In_2056);
nor U2307 (N_2307,In_1967,In_795);
nor U2308 (N_2308,In_2331,In_1339);
or U2309 (N_2309,In_1861,In_2388);
and U2310 (N_2310,In_888,In_1338);
nand U2311 (N_2311,In_2246,In_740);
and U2312 (N_2312,In_1167,In_294);
xnor U2313 (N_2313,In_477,In_2267);
and U2314 (N_2314,In_1462,In_2442);
and U2315 (N_2315,In_1450,In_1935);
or U2316 (N_2316,In_2389,In_1724);
nor U2317 (N_2317,In_1789,In_1276);
nand U2318 (N_2318,In_1750,In_1667);
nor U2319 (N_2319,In_1472,In_561);
nand U2320 (N_2320,In_686,In_896);
or U2321 (N_2321,In_296,In_1410);
nand U2322 (N_2322,In_1197,In_426);
nor U2323 (N_2323,In_1928,In_1002);
or U2324 (N_2324,In_2294,In_1801);
nand U2325 (N_2325,In_2356,In_197);
nand U2326 (N_2326,In_652,In_995);
or U2327 (N_2327,In_778,In_1997);
nand U2328 (N_2328,In_144,In_81);
nand U2329 (N_2329,In_1045,In_101);
nand U2330 (N_2330,In_5,In_1489);
xor U2331 (N_2331,In_2453,In_2008);
nand U2332 (N_2332,In_2299,In_687);
nor U2333 (N_2333,In_1047,In_8);
nand U2334 (N_2334,In_2321,In_2243);
nor U2335 (N_2335,In_72,In_177);
nor U2336 (N_2336,In_218,In_2160);
nor U2337 (N_2337,In_1261,In_1338);
or U2338 (N_2338,In_1633,In_1616);
nor U2339 (N_2339,In_1610,In_987);
xnor U2340 (N_2340,In_1678,In_1500);
xor U2341 (N_2341,In_614,In_353);
xnor U2342 (N_2342,In_823,In_2039);
and U2343 (N_2343,In_501,In_1271);
or U2344 (N_2344,In_661,In_60);
nand U2345 (N_2345,In_429,In_640);
nand U2346 (N_2346,In_1866,In_17);
nor U2347 (N_2347,In_2201,In_474);
xor U2348 (N_2348,In_405,In_647);
and U2349 (N_2349,In_326,In_1416);
nand U2350 (N_2350,In_2008,In_1599);
xor U2351 (N_2351,In_1676,In_1967);
nand U2352 (N_2352,In_1531,In_1684);
nor U2353 (N_2353,In_2062,In_2438);
nand U2354 (N_2354,In_1624,In_442);
nand U2355 (N_2355,In_1840,In_1172);
and U2356 (N_2356,In_2115,In_367);
or U2357 (N_2357,In_189,In_125);
nand U2358 (N_2358,In_1517,In_351);
and U2359 (N_2359,In_1140,In_2405);
or U2360 (N_2360,In_1987,In_1500);
or U2361 (N_2361,In_182,In_2069);
or U2362 (N_2362,In_942,In_2144);
nor U2363 (N_2363,In_691,In_2252);
or U2364 (N_2364,In_1538,In_731);
xor U2365 (N_2365,In_1487,In_1452);
xor U2366 (N_2366,In_763,In_2016);
nand U2367 (N_2367,In_394,In_404);
and U2368 (N_2368,In_303,In_176);
xnor U2369 (N_2369,In_1063,In_1016);
or U2370 (N_2370,In_2498,In_617);
xnor U2371 (N_2371,In_1777,In_2016);
nor U2372 (N_2372,In_1870,In_220);
nand U2373 (N_2373,In_1975,In_660);
nor U2374 (N_2374,In_743,In_366);
nand U2375 (N_2375,In_1427,In_1721);
nand U2376 (N_2376,In_1259,In_2082);
and U2377 (N_2377,In_707,In_2269);
nand U2378 (N_2378,In_2345,In_1102);
and U2379 (N_2379,In_2157,In_1168);
and U2380 (N_2380,In_708,In_1149);
or U2381 (N_2381,In_929,In_1561);
or U2382 (N_2382,In_1781,In_666);
nand U2383 (N_2383,In_1001,In_1598);
nand U2384 (N_2384,In_1122,In_1496);
or U2385 (N_2385,In_1943,In_559);
nor U2386 (N_2386,In_1854,In_2258);
nor U2387 (N_2387,In_723,In_449);
xnor U2388 (N_2388,In_722,In_1468);
nor U2389 (N_2389,In_2422,In_1222);
nand U2390 (N_2390,In_87,In_2102);
nor U2391 (N_2391,In_2434,In_2333);
xnor U2392 (N_2392,In_1352,In_760);
nand U2393 (N_2393,In_53,In_1826);
and U2394 (N_2394,In_1959,In_2242);
and U2395 (N_2395,In_296,In_856);
nand U2396 (N_2396,In_1713,In_1500);
and U2397 (N_2397,In_2205,In_1498);
nor U2398 (N_2398,In_2272,In_1571);
and U2399 (N_2399,In_552,In_1003);
nand U2400 (N_2400,In_1848,In_2433);
or U2401 (N_2401,In_330,In_1903);
and U2402 (N_2402,In_1506,In_1613);
or U2403 (N_2403,In_1191,In_1575);
and U2404 (N_2404,In_1476,In_298);
or U2405 (N_2405,In_1932,In_1486);
nor U2406 (N_2406,In_853,In_1724);
and U2407 (N_2407,In_210,In_2105);
nor U2408 (N_2408,In_1747,In_199);
or U2409 (N_2409,In_1074,In_1888);
and U2410 (N_2410,In_1908,In_150);
nand U2411 (N_2411,In_836,In_754);
nand U2412 (N_2412,In_217,In_478);
or U2413 (N_2413,In_459,In_1480);
and U2414 (N_2414,In_2218,In_1789);
nor U2415 (N_2415,In_1378,In_2283);
nor U2416 (N_2416,In_602,In_316);
and U2417 (N_2417,In_778,In_2287);
or U2418 (N_2418,In_1460,In_631);
xor U2419 (N_2419,In_38,In_453);
or U2420 (N_2420,In_1621,In_1470);
or U2421 (N_2421,In_1239,In_1535);
and U2422 (N_2422,In_570,In_1442);
or U2423 (N_2423,In_516,In_2138);
nand U2424 (N_2424,In_1861,In_1958);
and U2425 (N_2425,In_1733,In_1613);
and U2426 (N_2426,In_917,In_1822);
nand U2427 (N_2427,In_352,In_272);
nor U2428 (N_2428,In_819,In_49);
and U2429 (N_2429,In_1385,In_1873);
xnor U2430 (N_2430,In_392,In_1854);
nor U2431 (N_2431,In_2065,In_1271);
and U2432 (N_2432,In_1846,In_1685);
nand U2433 (N_2433,In_2015,In_572);
nor U2434 (N_2434,In_2123,In_1779);
or U2435 (N_2435,In_1274,In_2075);
nor U2436 (N_2436,In_1498,In_2398);
nand U2437 (N_2437,In_1074,In_650);
or U2438 (N_2438,In_1722,In_2107);
or U2439 (N_2439,In_326,In_595);
nand U2440 (N_2440,In_2173,In_1985);
nand U2441 (N_2441,In_2323,In_493);
or U2442 (N_2442,In_827,In_1901);
nand U2443 (N_2443,In_2033,In_133);
or U2444 (N_2444,In_476,In_1268);
nand U2445 (N_2445,In_830,In_157);
nand U2446 (N_2446,In_8,In_1056);
nand U2447 (N_2447,In_1962,In_159);
nor U2448 (N_2448,In_1992,In_1328);
nand U2449 (N_2449,In_1554,In_2213);
or U2450 (N_2450,In_359,In_1368);
nor U2451 (N_2451,In_944,In_2435);
xnor U2452 (N_2452,In_574,In_1747);
or U2453 (N_2453,In_1229,In_2432);
nor U2454 (N_2454,In_1114,In_1945);
and U2455 (N_2455,In_1352,In_1416);
and U2456 (N_2456,In_1945,In_100);
or U2457 (N_2457,In_1525,In_449);
and U2458 (N_2458,In_310,In_1251);
nand U2459 (N_2459,In_1815,In_1488);
and U2460 (N_2460,In_519,In_1983);
nor U2461 (N_2461,In_1447,In_684);
nor U2462 (N_2462,In_145,In_2269);
or U2463 (N_2463,In_1783,In_19);
and U2464 (N_2464,In_1245,In_837);
nand U2465 (N_2465,In_2111,In_2190);
or U2466 (N_2466,In_2374,In_1162);
and U2467 (N_2467,In_2440,In_411);
nor U2468 (N_2468,In_1405,In_1827);
nor U2469 (N_2469,In_1654,In_1509);
nor U2470 (N_2470,In_1353,In_1037);
nor U2471 (N_2471,In_563,In_2288);
nor U2472 (N_2472,In_879,In_803);
xor U2473 (N_2473,In_2374,In_1293);
xnor U2474 (N_2474,In_1020,In_1598);
nor U2475 (N_2475,In_621,In_2193);
xor U2476 (N_2476,In_64,In_1452);
xor U2477 (N_2477,In_137,In_1813);
xor U2478 (N_2478,In_1699,In_548);
nor U2479 (N_2479,In_593,In_1359);
and U2480 (N_2480,In_1616,In_562);
nor U2481 (N_2481,In_1709,In_2068);
or U2482 (N_2482,In_2007,In_70);
nand U2483 (N_2483,In_2051,In_1809);
or U2484 (N_2484,In_2179,In_1855);
nand U2485 (N_2485,In_2141,In_2002);
xnor U2486 (N_2486,In_256,In_1615);
and U2487 (N_2487,In_328,In_1415);
and U2488 (N_2488,In_1102,In_1724);
and U2489 (N_2489,In_2218,In_1279);
xor U2490 (N_2490,In_664,In_158);
and U2491 (N_2491,In_2218,In_110);
and U2492 (N_2492,In_1829,In_1434);
and U2493 (N_2493,In_2379,In_559);
or U2494 (N_2494,In_982,In_82);
nand U2495 (N_2495,In_1073,In_1175);
nor U2496 (N_2496,In_1110,In_756);
xor U2497 (N_2497,In_493,In_1287);
nand U2498 (N_2498,In_1132,In_414);
nor U2499 (N_2499,In_1822,In_1492);
nor U2500 (N_2500,In_1299,In_270);
or U2501 (N_2501,In_2154,In_2187);
nor U2502 (N_2502,In_1024,In_244);
nand U2503 (N_2503,In_2013,In_2169);
and U2504 (N_2504,In_668,In_418);
nand U2505 (N_2505,In_586,In_690);
and U2506 (N_2506,In_103,In_1254);
or U2507 (N_2507,In_1001,In_569);
nor U2508 (N_2508,In_1439,In_2422);
nand U2509 (N_2509,In_465,In_1947);
nand U2510 (N_2510,In_1608,In_2138);
nand U2511 (N_2511,In_2154,In_1055);
or U2512 (N_2512,In_1980,In_729);
nand U2513 (N_2513,In_374,In_4);
and U2514 (N_2514,In_566,In_876);
nor U2515 (N_2515,In_1251,In_2171);
or U2516 (N_2516,In_2467,In_315);
and U2517 (N_2517,In_554,In_157);
nor U2518 (N_2518,In_2200,In_199);
or U2519 (N_2519,In_994,In_2343);
nor U2520 (N_2520,In_606,In_1935);
nand U2521 (N_2521,In_312,In_2429);
xor U2522 (N_2522,In_949,In_916);
or U2523 (N_2523,In_490,In_1189);
or U2524 (N_2524,In_1832,In_2237);
and U2525 (N_2525,In_758,In_2166);
and U2526 (N_2526,In_1022,In_31);
or U2527 (N_2527,In_2192,In_536);
nor U2528 (N_2528,In_680,In_2134);
or U2529 (N_2529,In_1502,In_2230);
nand U2530 (N_2530,In_1211,In_1212);
or U2531 (N_2531,In_1491,In_924);
xnor U2532 (N_2532,In_1968,In_1932);
nor U2533 (N_2533,In_92,In_1945);
and U2534 (N_2534,In_1359,In_119);
or U2535 (N_2535,In_985,In_2150);
nand U2536 (N_2536,In_179,In_1913);
xnor U2537 (N_2537,In_98,In_1514);
or U2538 (N_2538,In_1135,In_757);
and U2539 (N_2539,In_857,In_2139);
or U2540 (N_2540,In_128,In_402);
nor U2541 (N_2541,In_512,In_189);
nand U2542 (N_2542,In_909,In_135);
and U2543 (N_2543,In_759,In_1301);
or U2544 (N_2544,In_2127,In_890);
nand U2545 (N_2545,In_1705,In_1816);
and U2546 (N_2546,In_1090,In_1412);
nand U2547 (N_2547,In_2238,In_2214);
nand U2548 (N_2548,In_433,In_1313);
and U2549 (N_2549,In_1025,In_1218);
or U2550 (N_2550,In_111,In_1389);
nand U2551 (N_2551,In_1466,In_1688);
nor U2552 (N_2552,In_805,In_1003);
or U2553 (N_2553,In_2141,In_503);
and U2554 (N_2554,In_931,In_2257);
and U2555 (N_2555,In_1930,In_114);
nand U2556 (N_2556,In_1397,In_1063);
or U2557 (N_2557,In_2109,In_1401);
or U2558 (N_2558,In_976,In_2037);
nor U2559 (N_2559,In_28,In_2465);
nor U2560 (N_2560,In_1475,In_1785);
and U2561 (N_2561,In_2294,In_2034);
nand U2562 (N_2562,In_960,In_373);
or U2563 (N_2563,In_2070,In_1670);
and U2564 (N_2564,In_146,In_162);
nand U2565 (N_2565,In_565,In_2257);
or U2566 (N_2566,In_2066,In_627);
or U2567 (N_2567,In_2400,In_1545);
nor U2568 (N_2568,In_1329,In_776);
nand U2569 (N_2569,In_760,In_693);
and U2570 (N_2570,In_361,In_667);
nand U2571 (N_2571,In_528,In_289);
nor U2572 (N_2572,In_2251,In_2461);
xor U2573 (N_2573,In_2219,In_1723);
nor U2574 (N_2574,In_1661,In_2264);
nand U2575 (N_2575,In_1454,In_540);
or U2576 (N_2576,In_1062,In_2221);
nand U2577 (N_2577,In_2429,In_2456);
and U2578 (N_2578,In_770,In_229);
and U2579 (N_2579,In_9,In_2308);
or U2580 (N_2580,In_159,In_994);
and U2581 (N_2581,In_1602,In_2340);
and U2582 (N_2582,In_460,In_1216);
nor U2583 (N_2583,In_485,In_351);
nand U2584 (N_2584,In_1011,In_1939);
and U2585 (N_2585,In_1538,In_2167);
nand U2586 (N_2586,In_2414,In_1434);
and U2587 (N_2587,In_996,In_2234);
xnor U2588 (N_2588,In_423,In_2052);
or U2589 (N_2589,In_1458,In_1768);
nor U2590 (N_2590,In_1357,In_2241);
xnor U2591 (N_2591,In_431,In_984);
or U2592 (N_2592,In_470,In_1304);
and U2593 (N_2593,In_702,In_902);
nand U2594 (N_2594,In_2363,In_1231);
or U2595 (N_2595,In_180,In_1461);
xor U2596 (N_2596,In_1140,In_43);
nor U2597 (N_2597,In_812,In_2323);
and U2598 (N_2598,In_1689,In_841);
or U2599 (N_2599,In_1410,In_2073);
nand U2600 (N_2600,In_1899,In_2485);
and U2601 (N_2601,In_1031,In_1849);
and U2602 (N_2602,In_1503,In_494);
and U2603 (N_2603,In_941,In_621);
nand U2604 (N_2604,In_1102,In_375);
and U2605 (N_2605,In_1876,In_252);
or U2606 (N_2606,In_470,In_2421);
or U2607 (N_2607,In_822,In_88);
nand U2608 (N_2608,In_2219,In_871);
nand U2609 (N_2609,In_1496,In_547);
or U2610 (N_2610,In_712,In_1163);
or U2611 (N_2611,In_2253,In_1908);
nand U2612 (N_2612,In_1445,In_2439);
xor U2613 (N_2613,In_1274,In_1696);
nand U2614 (N_2614,In_2281,In_964);
or U2615 (N_2615,In_47,In_2233);
and U2616 (N_2616,In_655,In_967);
nand U2617 (N_2617,In_742,In_1905);
nand U2618 (N_2618,In_2003,In_808);
or U2619 (N_2619,In_486,In_336);
nand U2620 (N_2620,In_1689,In_2142);
or U2621 (N_2621,In_208,In_1812);
nor U2622 (N_2622,In_1369,In_1337);
nand U2623 (N_2623,In_1332,In_608);
nor U2624 (N_2624,In_711,In_246);
xor U2625 (N_2625,In_472,In_614);
nor U2626 (N_2626,In_1336,In_460);
nor U2627 (N_2627,In_1266,In_871);
or U2628 (N_2628,In_2160,In_635);
xnor U2629 (N_2629,In_2336,In_791);
or U2630 (N_2630,In_579,In_672);
nor U2631 (N_2631,In_2331,In_1302);
and U2632 (N_2632,In_1713,In_843);
xnor U2633 (N_2633,In_928,In_1656);
and U2634 (N_2634,In_1987,In_45);
and U2635 (N_2635,In_2364,In_1474);
nand U2636 (N_2636,In_2302,In_10);
nand U2637 (N_2637,In_1681,In_1223);
and U2638 (N_2638,In_1273,In_1194);
and U2639 (N_2639,In_504,In_2450);
nor U2640 (N_2640,In_585,In_1159);
nor U2641 (N_2641,In_2384,In_2359);
nand U2642 (N_2642,In_2229,In_1243);
or U2643 (N_2643,In_845,In_1789);
nand U2644 (N_2644,In_1360,In_1138);
and U2645 (N_2645,In_980,In_1162);
or U2646 (N_2646,In_945,In_1147);
and U2647 (N_2647,In_591,In_2109);
or U2648 (N_2648,In_1058,In_1851);
and U2649 (N_2649,In_2408,In_1597);
and U2650 (N_2650,In_1825,In_1806);
or U2651 (N_2651,In_149,In_2104);
and U2652 (N_2652,In_1337,In_1108);
or U2653 (N_2653,In_553,In_68);
and U2654 (N_2654,In_2029,In_1251);
and U2655 (N_2655,In_1991,In_1111);
xor U2656 (N_2656,In_1084,In_1211);
nor U2657 (N_2657,In_1472,In_1941);
or U2658 (N_2658,In_878,In_1496);
and U2659 (N_2659,In_2415,In_1663);
and U2660 (N_2660,In_109,In_752);
xnor U2661 (N_2661,In_1959,In_1680);
nor U2662 (N_2662,In_1869,In_1774);
or U2663 (N_2663,In_1290,In_831);
nand U2664 (N_2664,In_2020,In_1241);
nor U2665 (N_2665,In_763,In_2298);
and U2666 (N_2666,In_2448,In_2439);
and U2667 (N_2667,In_831,In_1436);
or U2668 (N_2668,In_903,In_794);
nor U2669 (N_2669,In_708,In_1303);
and U2670 (N_2670,In_793,In_83);
xnor U2671 (N_2671,In_910,In_374);
and U2672 (N_2672,In_1273,In_375);
and U2673 (N_2673,In_1292,In_956);
nand U2674 (N_2674,In_879,In_511);
nor U2675 (N_2675,In_1454,In_106);
nand U2676 (N_2676,In_1247,In_1978);
or U2677 (N_2677,In_964,In_1628);
nor U2678 (N_2678,In_189,In_736);
nand U2679 (N_2679,In_435,In_1801);
nand U2680 (N_2680,In_200,In_954);
or U2681 (N_2681,In_1342,In_2467);
and U2682 (N_2682,In_1164,In_1396);
nor U2683 (N_2683,In_328,In_1759);
nand U2684 (N_2684,In_1321,In_1965);
xnor U2685 (N_2685,In_92,In_544);
nor U2686 (N_2686,In_1651,In_2348);
nand U2687 (N_2687,In_1387,In_107);
and U2688 (N_2688,In_408,In_677);
nand U2689 (N_2689,In_1046,In_1582);
nand U2690 (N_2690,In_1172,In_991);
or U2691 (N_2691,In_2198,In_1230);
xor U2692 (N_2692,In_528,In_1659);
and U2693 (N_2693,In_804,In_1103);
nor U2694 (N_2694,In_2043,In_926);
nand U2695 (N_2695,In_165,In_534);
and U2696 (N_2696,In_315,In_1494);
or U2697 (N_2697,In_1945,In_714);
or U2698 (N_2698,In_2354,In_568);
and U2699 (N_2699,In_2301,In_1980);
nor U2700 (N_2700,In_766,In_1612);
or U2701 (N_2701,In_280,In_1155);
and U2702 (N_2702,In_2121,In_2002);
and U2703 (N_2703,In_777,In_595);
xnor U2704 (N_2704,In_1730,In_1921);
nor U2705 (N_2705,In_650,In_2283);
nand U2706 (N_2706,In_1453,In_119);
nand U2707 (N_2707,In_9,In_1649);
or U2708 (N_2708,In_2156,In_1202);
nand U2709 (N_2709,In_1636,In_1558);
and U2710 (N_2710,In_2206,In_1849);
and U2711 (N_2711,In_551,In_2336);
nand U2712 (N_2712,In_1765,In_1580);
or U2713 (N_2713,In_1596,In_623);
or U2714 (N_2714,In_45,In_1662);
and U2715 (N_2715,In_1369,In_1088);
nor U2716 (N_2716,In_1105,In_1283);
or U2717 (N_2717,In_495,In_365);
nand U2718 (N_2718,In_260,In_971);
nor U2719 (N_2719,In_591,In_980);
nor U2720 (N_2720,In_1109,In_668);
or U2721 (N_2721,In_786,In_1282);
and U2722 (N_2722,In_1866,In_2432);
xor U2723 (N_2723,In_1782,In_1054);
or U2724 (N_2724,In_1233,In_125);
and U2725 (N_2725,In_863,In_1855);
and U2726 (N_2726,In_2010,In_1802);
or U2727 (N_2727,In_400,In_2119);
nand U2728 (N_2728,In_1566,In_2002);
or U2729 (N_2729,In_451,In_633);
or U2730 (N_2730,In_1841,In_1445);
xor U2731 (N_2731,In_1269,In_1656);
and U2732 (N_2732,In_2157,In_1977);
nor U2733 (N_2733,In_936,In_1044);
and U2734 (N_2734,In_2358,In_121);
or U2735 (N_2735,In_783,In_1719);
or U2736 (N_2736,In_635,In_1969);
and U2737 (N_2737,In_329,In_746);
nand U2738 (N_2738,In_1577,In_2243);
nor U2739 (N_2739,In_1017,In_982);
or U2740 (N_2740,In_573,In_2107);
nand U2741 (N_2741,In_1223,In_1064);
nor U2742 (N_2742,In_332,In_268);
or U2743 (N_2743,In_700,In_1559);
nor U2744 (N_2744,In_256,In_1015);
and U2745 (N_2745,In_1716,In_1852);
nor U2746 (N_2746,In_1628,In_220);
nor U2747 (N_2747,In_1183,In_1398);
xnor U2748 (N_2748,In_52,In_76);
nor U2749 (N_2749,In_1396,In_998);
nor U2750 (N_2750,In_829,In_1293);
xnor U2751 (N_2751,In_1862,In_2046);
or U2752 (N_2752,In_384,In_1886);
nand U2753 (N_2753,In_1258,In_2303);
and U2754 (N_2754,In_1492,In_1100);
and U2755 (N_2755,In_2187,In_1837);
and U2756 (N_2756,In_968,In_2087);
nor U2757 (N_2757,In_1007,In_2430);
and U2758 (N_2758,In_1906,In_1339);
or U2759 (N_2759,In_1884,In_2410);
or U2760 (N_2760,In_2215,In_1282);
nand U2761 (N_2761,In_252,In_1607);
and U2762 (N_2762,In_710,In_2082);
nand U2763 (N_2763,In_1887,In_2439);
xor U2764 (N_2764,In_102,In_2002);
nor U2765 (N_2765,In_2244,In_1921);
or U2766 (N_2766,In_648,In_2125);
nand U2767 (N_2767,In_230,In_334);
nor U2768 (N_2768,In_2408,In_2454);
and U2769 (N_2769,In_2019,In_1003);
nand U2770 (N_2770,In_727,In_1329);
xor U2771 (N_2771,In_1440,In_1745);
nand U2772 (N_2772,In_1636,In_2098);
nand U2773 (N_2773,In_1486,In_1109);
xnor U2774 (N_2774,In_2087,In_317);
and U2775 (N_2775,In_1201,In_984);
and U2776 (N_2776,In_660,In_360);
xor U2777 (N_2777,In_1578,In_1668);
or U2778 (N_2778,In_661,In_1283);
or U2779 (N_2779,In_2306,In_1815);
nand U2780 (N_2780,In_367,In_797);
or U2781 (N_2781,In_1919,In_127);
nor U2782 (N_2782,In_1420,In_2283);
and U2783 (N_2783,In_2301,In_198);
or U2784 (N_2784,In_746,In_776);
and U2785 (N_2785,In_996,In_1589);
or U2786 (N_2786,In_2160,In_799);
or U2787 (N_2787,In_2018,In_1705);
xnor U2788 (N_2788,In_556,In_1926);
nand U2789 (N_2789,In_335,In_1677);
nand U2790 (N_2790,In_630,In_539);
nor U2791 (N_2791,In_805,In_930);
nand U2792 (N_2792,In_2073,In_1503);
and U2793 (N_2793,In_1557,In_2479);
nor U2794 (N_2794,In_576,In_908);
nand U2795 (N_2795,In_1039,In_1966);
and U2796 (N_2796,In_735,In_361);
and U2797 (N_2797,In_0,In_2121);
nand U2798 (N_2798,In_446,In_1539);
nand U2799 (N_2799,In_627,In_2469);
xor U2800 (N_2800,In_628,In_2131);
xor U2801 (N_2801,In_773,In_411);
or U2802 (N_2802,In_75,In_178);
nand U2803 (N_2803,In_402,In_285);
nand U2804 (N_2804,In_1919,In_310);
nand U2805 (N_2805,In_728,In_571);
nand U2806 (N_2806,In_1873,In_610);
or U2807 (N_2807,In_999,In_789);
nand U2808 (N_2808,In_1538,In_1118);
nand U2809 (N_2809,In_754,In_1185);
xor U2810 (N_2810,In_1651,In_570);
and U2811 (N_2811,In_962,In_1376);
nand U2812 (N_2812,In_97,In_2007);
nor U2813 (N_2813,In_2156,In_2037);
and U2814 (N_2814,In_582,In_2173);
nor U2815 (N_2815,In_69,In_2057);
or U2816 (N_2816,In_151,In_2240);
xnor U2817 (N_2817,In_327,In_2395);
nand U2818 (N_2818,In_1909,In_666);
and U2819 (N_2819,In_152,In_2389);
nor U2820 (N_2820,In_1583,In_1591);
nand U2821 (N_2821,In_1586,In_1710);
nor U2822 (N_2822,In_2045,In_2025);
or U2823 (N_2823,In_1509,In_1042);
and U2824 (N_2824,In_2151,In_712);
xor U2825 (N_2825,In_1716,In_661);
nor U2826 (N_2826,In_1200,In_70);
nor U2827 (N_2827,In_680,In_1090);
or U2828 (N_2828,In_728,In_333);
or U2829 (N_2829,In_519,In_228);
and U2830 (N_2830,In_56,In_2418);
xor U2831 (N_2831,In_1481,In_853);
or U2832 (N_2832,In_1352,In_2252);
nor U2833 (N_2833,In_228,In_650);
and U2834 (N_2834,In_1213,In_1474);
and U2835 (N_2835,In_736,In_90);
and U2836 (N_2836,In_416,In_1786);
nand U2837 (N_2837,In_457,In_1301);
and U2838 (N_2838,In_880,In_1177);
xnor U2839 (N_2839,In_975,In_2234);
xor U2840 (N_2840,In_2383,In_978);
or U2841 (N_2841,In_336,In_286);
and U2842 (N_2842,In_1876,In_2141);
or U2843 (N_2843,In_393,In_878);
or U2844 (N_2844,In_334,In_1315);
or U2845 (N_2845,In_1493,In_1896);
or U2846 (N_2846,In_2279,In_1096);
and U2847 (N_2847,In_1061,In_1897);
or U2848 (N_2848,In_586,In_2211);
nor U2849 (N_2849,In_404,In_1764);
or U2850 (N_2850,In_630,In_1219);
nor U2851 (N_2851,In_341,In_1003);
and U2852 (N_2852,In_981,In_2207);
nor U2853 (N_2853,In_2097,In_1275);
or U2854 (N_2854,In_1047,In_1622);
nor U2855 (N_2855,In_483,In_926);
and U2856 (N_2856,In_97,In_2253);
xor U2857 (N_2857,In_1653,In_175);
or U2858 (N_2858,In_1933,In_1214);
nand U2859 (N_2859,In_2382,In_342);
or U2860 (N_2860,In_397,In_468);
or U2861 (N_2861,In_762,In_1442);
or U2862 (N_2862,In_139,In_1052);
nand U2863 (N_2863,In_1579,In_231);
and U2864 (N_2864,In_1655,In_2002);
or U2865 (N_2865,In_2362,In_234);
nand U2866 (N_2866,In_1720,In_1716);
xnor U2867 (N_2867,In_1808,In_2074);
nand U2868 (N_2868,In_1767,In_925);
or U2869 (N_2869,In_2398,In_489);
nand U2870 (N_2870,In_2449,In_1289);
and U2871 (N_2871,In_374,In_1017);
or U2872 (N_2872,In_1500,In_1946);
nand U2873 (N_2873,In_2162,In_1401);
or U2874 (N_2874,In_200,In_889);
nor U2875 (N_2875,In_1752,In_2423);
and U2876 (N_2876,In_1631,In_1297);
nor U2877 (N_2877,In_106,In_2042);
nand U2878 (N_2878,In_1641,In_278);
nor U2879 (N_2879,In_897,In_644);
and U2880 (N_2880,In_1705,In_1379);
nor U2881 (N_2881,In_1485,In_2250);
or U2882 (N_2882,In_1945,In_348);
nand U2883 (N_2883,In_507,In_139);
and U2884 (N_2884,In_2144,In_1721);
or U2885 (N_2885,In_2080,In_284);
and U2886 (N_2886,In_1450,In_1050);
or U2887 (N_2887,In_1937,In_904);
nand U2888 (N_2888,In_1780,In_2303);
and U2889 (N_2889,In_946,In_589);
nand U2890 (N_2890,In_181,In_1178);
and U2891 (N_2891,In_2199,In_1237);
nand U2892 (N_2892,In_987,In_1959);
nand U2893 (N_2893,In_2125,In_1908);
nand U2894 (N_2894,In_468,In_626);
and U2895 (N_2895,In_2293,In_1433);
xnor U2896 (N_2896,In_288,In_404);
xnor U2897 (N_2897,In_1702,In_159);
nand U2898 (N_2898,In_1254,In_1505);
nor U2899 (N_2899,In_200,In_1923);
nand U2900 (N_2900,In_753,In_984);
nor U2901 (N_2901,In_722,In_1428);
xnor U2902 (N_2902,In_55,In_1489);
or U2903 (N_2903,In_2323,In_1332);
and U2904 (N_2904,In_311,In_1143);
and U2905 (N_2905,In_2270,In_2054);
nor U2906 (N_2906,In_917,In_2140);
xor U2907 (N_2907,In_1734,In_1433);
nand U2908 (N_2908,In_2259,In_345);
or U2909 (N_2909,In_280,In_1395);
nand U2910 (N_2910,In_18,In_496);
nor U2911 (N_2911,In_2084,In_2170);
or U2912 (N_2912,In_1437,In_2350);
nand U2913 (N_2913,In_2118,In_229);
or U2914 (N_2914,In_2006,In_1017);
nand U2915 (N_2915,In_2462,In_865);
nor U2916 (N_2916,In_2130,In_1870);
nand U2917 (N_2917,In_240,In_624);
and U2918 (N_2918,In_2316,In_232);
and U2919 (N_2919,In_108,In_737);
or U2920 (N_2920,In_2148,In_118);
xnor U2921 (N_2921,In_1367,In_2377);
nand U2922 (N_2922,In_2410,In_861);
and U2923 (N_2923,In_770,In_1337);
nand U2924 (N_2924,In_1210,In_1137);
nor U2925 (N_2925,In_1758,In_2156);
nand U2926 (N_2926,In_2337,In_2311);
nand U2927 (N_2927,In_1433,In_351);
nand U2928 (N_2928,In_315,In_384);
nor U2929 (N_2929,In_1361,In_1886);
nor U2930 (N_2930,In_477,In_1798);
and U2931 (N_2931,In_1111,In_1159);
xor U2932 (N_2932,In_1285,In_1179);
nor U2933 (N_2933,In_1472,In_2233);
xnor U2934 (N_2934,In_1768,In_2443);
and U2935 (N_2935,In_1618,In_1379);
nor U2936 (N_2936,In_1182,In_750);
or U2937 (N_2937,In_880,In_1805);
and U2938 (N_2938,In_337,In_62);
and U2939 (N_2939,In_831,In_848);
and U2940 (N_2940,In_2381,In_1713);
nand U2941 (N_2941,In_2095,In_453);
nand U2942 (N_2942,In_2204,In_1134);
and U2943 (N_2943,In_1134,In_1142);
and U2944 (N_2944,In_101,In_1019);
or U2945 (N_2945,In_1753,In_1951);
nor U2946 (N_2946,In_2013,In_600);
nand U2947 (N_2947,In_227,In_1501);
nor U2948 (N_2948,In_965,In_1579);
and U2949 (N_2949,In_1516,In_2447);
or U2950 (N_2950,In_1915,In_707);
nand U2951 (N_2951,In_812,In_1880);
or U2952 (N_2952,In_158,In_1925);
nand U2953 (N_2953,In_2278,In_686);
nor U2954 (N_2954,In_2434,In_552);
or U2955 (N_2955,In_217,In_166);
nor U2956 (N_2956,In_443,In_1397);
nor U2957 (N_2957,In_1763,In_1368);
nor U2958 (N_2958,In_2068,In_1712);
nand U2959 (N_2959,In_1031,In_2267);
or U2960 (N_2960,In_2434,In_346);
or U2961 (N_2961,In_661,In_2448);
nor U2962 (N_2962,In_501,In_586);
and U2963 (N_2963,In_529,In_2044);
xor U2964 (N_2964,In_927,In_461);
nor U2965 (N_2965,In_1082,In_932);
nand U2966 (N_2966,In_1899,In_121);
xnor U2967 (N_2967,In_99,In_1901);
or U2968 (N_2968,In_1749,In_799);
or U2969 (N_2969,In_672,In_1215);
and U2970 (N_2970,In_1449,In_1736);
nor U2971 (N_2971,In_2284,In_2381);
and U2972 (N_2972,In_272,In_2315);
and U2973 (N_2973,In_1271,In_1302);
nand U2974 (N_2974,In_1274,In_54);
and U2975 (N_2975,In_2469,In_641);
nand U2976 (N_2976,In_1408,In_1052);
or U2977 (N_2977,In_220,In_774);
and U2978 (N_2978,In_1666,In_2365);
xnor U2979 (N_2979,In_853,In_222);
nor U2980 (N_2980,In_2059,In_632);
nand U2981 (N_2981,In_870,In_89);
or U2982 (N_2982,In_202,In_444);
or U2983 (N_2983,In_1631,In_1467);
nand U2984 (N_2984,In_1146,In_1373);
nand U2985 (N_2985,In_2158,In_2255);
or U2986 (N_2986,In_1685,In_1464);
or U2987 (N_2987,In_1541,In_1969);
nor U2988 (N_2988,In_475,In_330);
or U2989 (N_2989,In_343,In_398);
or U2990 (N_2990,In_1566,In_2082);
nand U2991 (N_2991,In_2343,In_1364);
nor U2992 (N_2992,In_772,In_2013);
and U2993 (N_2993,In_401,In_697);
and U2994 (N_2994,In_1802,In_2326);
and U2995 (N_2995,In_1026,In_1771);
or U2996 (N_2996,In_2056,In_1073);
and U2997 (N_2997,In_1077,In_805);
xnor U2998 (N_2998,In_1662,In_402);
or U2999 (N_2999,In_844,In_1739);
or U3000 (N_3000,In_2340,In_139);
nor U3001 (N_3001,In_2165,In_979);
nand U3002 (N_3002,In_613,In_859);
nand U3003 (N_3003,In_2335,In_942);
xnor U3004 (N_3004,In_2444,In_1189);
nor U3005 (N_3005,In_1441,In_2008);
xor U3006 (N_3006,In_1761,In_2091);
xnor U3007 (N_3007,In_1654,In_1170);
or U3008 (N_3008,In_183,In_2361);
nand U3009 (N_3009,In_735,In_1824);
nand U3010 (N_3010,In_2057,In_1865);
nand U3011 (N_3011,In_384,In_68);
or U3012 (N_3012,In_2365,In_814);
and U3013 (N_3013,In_1285,In_2127);
or U3014 (N_3014,In_1719,In_1036);
nor U3015 (N_3015,In_2109,In_1122);
xor U3016 (N_3016,In_2434,In_2137);
nor U3017 (N_3017,In_325,In_402);
nor U3018 (N_3018,In_1144,In_1733);
nand U3019 (N_3019,In_905,In_837);
nor U3020 (N_3020,In_638,In_863);
nor U3021 (N_3021,In_579,In_1396);
and U3022 (N_3022,In_240,In_703);
nor U3023 (N_3023,In_1223,In_354);
or U3024 (N_3024,In_1105,In_124);
nor U3025 (N_3025,In_2123,In_2275);
nor U3026 (N_3026,In_1713,In_336);
and U3027 (N_3027,In_1065,In_1597);
nor U3028 (N_3028,In_1705,In_2381);
and U3029 (N_3029,In_2044,In_998);
or U3030 (N_3030,In_727,In_1874);
or U3031 (N_3031,In_1577,In_1731);
nor U3032 (N_3032,In_567,In_1267);
and U3033 (N_3033,In_2300,In_332);
xor U3034 (N_3034,In_272,In_601);
or U3035 (N_3035,In_2414,In_2144);
nand U3036 (N_3036,In_361,In_2383);
nor U3037 (N_3037,In_82,In_2029);
or U3038 (N_3038,In_884,In_2258);
and U3039 (N_3039,In_1497,In_393);
nor U3040 (N_3040,In_1465,In_2014);
or U3041 (N_3041,In_1053,In_1236);
or U3042 (N_3042,In_376,In_2049);
and U3043 (N_3043,In_2335,In_269);
xor U3044 (N_3044,In_1752,In_1311);
and U3045 (N_3045,In_1623,In_2440);
nor U3046 (N_3046,In_1623,In_2304);
or U3047 (N_3047,In_660,In_236);
or U3048 (N_3048,In_348,In_1361);
or U3049 (N_3049,In_1718,In_711);
and U3050 (N_3050,In_693,In_935);
nor U3051 (N_3051,In_2168,In_1495);
nor U3052 (N_3052,In_18,In_630);
and U3053 (N_3053,In_48,In_1486);
and U3054 (N_3054,In_681,In_2484);
nor U3055 (N_3055,In_2024,In_1630);
and U3056 (N_3056,In_2424,In_1434);
nor U3057 (N_3057,In_398,In_354);
nor U3058 (N_3058,In_1770,In_1030);
nor U3059 (N_3059,In_98,In_2398);
nand U3060 (N_3060,In_1998,In_666);
nand U3061 (N_3061,In_303,In_1733);
nand U3062 (N_3062,In_1072,In_638);
nor U3063 (N_3063,In_1592,In_220);
nand U3064 (N_3064,In_799,In_1435);
nor U3065 (N_3065,In_1743,In_703);
xnor U3066 (N_3066,In_624,In_1684);
and U3067 (N_3067,In_2004,In_1494);
nand U3068 (N_3068,In_800,In_431);
or U3069 (N_3069,In_1092,In_1147);
and U3070 (N_3070,In_772,In_1790);
or U3071 (N_3071,In_2120,In_531);
and U3072 (N_3072,In_1410,In_1163);
nor U3073 (N_3073,In_1836,In_363);
nand U3074 (N_3074,In_2421,In_2271);
or U3075 (N_3075,In_95,In_2150);
nand U3076 (N_3076,In_706,In_1942);
and U3077 (N_3077,In_539,In_1121);
nor U3078 (N_3078,In_539,In_917);
nand U3079 (N_3079,In_25,In_1372);
or U3080 (N_3080,In_336,In_1346);
and U3081 (N_3081,In_1913,In_1487);
xnor U3082 (N_3082,In_2357,In_175);
nor U3083 (N_3083,In_13,In_770);
nor U3084 (N_3084,In_326,In_1467);
nor U3085 (N_3085,In_950,In_497);
or U3086 (N_3086,In_823,In_159);
nand U3087 (N_3087,In_1376,In_117);
and U3088 (N_3088,In_2481,In_2393);
and U3089 (N_3089,In_2275,In_2476);
nand U3090 (N_3090,In_1857,In_2212);
or U3091 (N_3091,In_2285,In_513);
nor U3092 (N_3092,In_1709,In_544);
or U3093 (N_3093,In_1800,In_279);
nand U3094 (N_3094,In_665,In_573);
nor U3095 (N_3095,In_643,In_644);
and U3096 (N_3096,In_2285,In_598);
nand U3097 (N_3097,In_1387,In_1007);
xnor U3098 (N_3098,In_324,In_652);
or U3099 (N_3099,In_725,In_1700);
nand U3100 (N_3100,In_1391,In_346);
nor U3101 (N_3101,In_2069,In_591);
nor U3102 (N_3102,In_1738,In_2404);
or U3103 (N_3103,In_1742,In_413);
nand U3104 (N_3104,In_2452,In_2187);
xor U3105 (N_3105,In_1579,In_634);
nand U3106 (N_3106,In_1046,In_2338);
nor U3107 (N_3107,In_2320,In_2358);
or U3108 (N_3108,In_1665,In_453);
and U3109 (N_3109,In_383,In_553);
or U3110 (N_3110,In_1719,In_236);
nand U3111 (N_3111,In_2391,In_1086);
nor U3112 (N_3112,In_1365,In_127);
nor U3113 (N_3113,In_1265,In_416);
and U3114 (N_3114,In_357,In_1846);
or U3115 (N_3115,In_2385,In_1629);
or U3116 (N_3116,In_91,In_2250);
or U3117 (N_3117,In_564,In_765);
or U3118 (N_3118,In_1078,In_619);
or U3119 (N_3119,In_330,In_2012);
or U3120 (N_3120,In_1260,In_357);
or U3121 (N_3121,In_1435,In_278);
nand U3122 (N_3122,In_762,In_1263);
nor U3123 (N_3123,In_1912,In_1538);
or U3124 (N_3124,In_1028,In_2452);
nand U3125 (N_3125,In_1618,In_63);
nand U3126 (N_3126,In_441,In_515);
nor U3127 (N_3127,In_2033,In_2314);
and U3128 (N_3128,In_1014,In_1033);
nand U3129 (N_3129,In_1019,In_2084);
xor U3130 (N_3130,In_2379,In_1608);
nor U3131 (N_3131,In_824,In_555);
nand U3132 (N_3132,In_152,In_606);
and U3133 (N_3133,In_1056,In_1454);
or U3134 (N_3134,In_1730,In_296);
nor U3135 (N_3135,In_1699,In_1356);
nand U3136 (N_3136,In_1971,In_992);
xor U3137 (N_3137,In_240,In_724);
and U3138 (N_3138,In_1541,In_929);
or U3139 (N_3139,In_809,In_163);
or U3140 (N_3140,In_706,In_1775);
or U3141 (N_3141,In_2300,In_675);
and U3142 (N_3142,In_1211,In_1975);
nand U3143 (N_3143,In_1973,In_1596);
nor U3144 (N_3144,In_2484,In_175);
and U3145 (N_3145,In_1190,In_2215);
nor U3146 (N_3146,In_1763,In_1418);
xnor U3147 (N_3147,In_1320,In_1415);
and U3148 (N_3148,In_1926,In_153);
and U3149 (N_3149,In_950,In_366);
xor U3150 (N_3150,In_659,In_1063);
nor U3151 (N_3151,In_1198,In_820);
nor U3152 (N_3152,In_1538,In_1587);
nand U3153 (N_3153,In_1226,In_2248);
and U3154 (N_3154,In_1034,In_797);
nand U3155 (N_3155,In_724,In_1050);
and U3156 (N_3156,In_2242,In_1924);
and U3157 (N_3157,In_775,In_324);
and U3158 (N_3158,In_1316,In_624);
or U3159 (N_3159,In_896,In_1993);
or U3160 (N_3160,In_1356,In_1364);
and U3161 (N_3161,In_228,In_1890);
or U3162 (N_3162,In_577,In_2318);
nand U3163 (N_3163,In_573,In_1851);
nor U3164 (N_3164,In_850,In_64);
nand U3165 (N_3165,In_0,In_1563);
xnor U3166 (N_3166,In_1687,In_1433);
or U3167 (N_3167,In_1417,In_842);
nand U3168 (N_3168,In_416,In_1935);
nand U3169 (N_3169,In_302,In_493);
or U3170 (N_3170,In_1326,In_65);
nand U3171 (N_3171,In_422,In_992);
nand U3172 (N_3172,In_1808,In_2161);
nand U3173 (N_3173,In_1718,In_1010);
and U3174 (N_3174,In_855,In_1667);
xnor U3175 (N_3175,In_279,In_47);
and U3176 (N_3176,In_2164,In_396);
and U3177 (N_3177,In_2296,In_2019);
nor U3178 (N_3178,In_608,In_1456);
nor U3179 (N_3179,In_2185,In_1049);
nand U3180 (N_3180,In_1830,In_1265);
xor U3181 (N_3181,In_695,In_1294);
nand U3182 (N_3182,In_1775,In_793);
nand U3183 (N_3183,In_827,In_731);
nand U3184 (N_3184,In_1440,In_1019);
nand U3185 (N_3185,In_1524,In_90);
or U3186 (N_3186,In_312,In_1526);
nand U3187 (N_3187,In_953,In_734);
and U3188 (N_3188,In_665,In_914);
nand U3189 (N_3189,In_1476,In_577);
or U3190 (N_3190,In_2190,In_607);
nor U3191 (N_3191,In_834,In_1451);
nor U3192 (N_3192,In_2068,In_1153);
nand U3193 (N_3193,In_2130,In_2266);
and U3194 (N_3194,In_1771,In_1322);
or U3195 (N_3195,In_1259,In_2114);
or U3196 (N_3196,In_202,In_1355);
nor U3197 (N_3197,In_1714,In_1774);
or U3198 (N_3198,In_1810,In_455);
nand U3199 (N_3199,In_87,In_1139);
nand U3200 (N_3200,In_2171,In_190);
or U3201 (N_3201,In_486,In_1584);
or U3202 (N_3202,In_1024,In_148);
xnor U3203 (N_3203,In_176,In_1794);
or U3204 (N_3204,In_2390,In_2275);
and U3205 (N_3205,In_1749,In_2016);
and U3206 (N_3206,In_1275,In_2030);
and U3207 (N_3207,In_1156,In_918);
nor U3208 (N_3208,In_490,In_291);
nor U3209 (N_3209,In_762,In_394);
nand U3210 (N_3210,In_2067,In_1937);
and U3211 (N_3211,In_1537,In_1718);
or U3212 (N_3212,In_1296,In_817);
and U3213 (N_3213,In_16,In_234);
and U3214 (N_3214,In_452,In_1178);
nor U3215 (N_3215,In_398,In_1562);
and U3216 (N_3216,In_2167,In_2127);
or U3217 (N_3217,In_271,In_998);
and U3218 (N_3218,In_1444,In_1413);
and U3219 (N_3219,In_147,In_462);
or U3220 (N_3220,In_1107,In_756);
nor U3221 (N_3221,In_1462,In_2132);
and U3222 (N_3222,In_1460,In_1956);
and U3223 (N_3223,In_493,In_755);
or U3224 (N_3224,In_277,In_1031);
nor U3225 (N_3225,In_512,In_794);
and U3226 (N_3226,In_1417,In_2092);
and U3227 (N_3227,In_299,In_1905);
nand U3228 (N_3228,In_984,In_1585);
and U3229 (N_3229,In_2455,In_1574);
nand U3230 (N_3230,In_2319,In_598);
and U3231 (N_3231,In_734,In_1104);
nor U3232 (N_3232,In_563,In_1359);
and U3233 (N_3233,In_1330,In_84);
nor U3234 (N_3234,In_1439,In_1275);
and U3235 (N_3235,In_1560,In_166);
xnor U3236 (N_3236,In_423,In_535);
and U3237 (N_3237,In_2072,In_664);
and U3238 (N_3238,In_1406,In_262);
and U3239 (N_3239,In_1975,In_667);
and U3240 (N_3240,In_1506,In_394);
and U3241 (N_3241,In_1177,In_201);
or U3242 (N_3242,In_2271,In_1513);
and U3243 (N_3243,In_2423,In_1294);
xnor U3244 (N_3244,In_2431,In_1679);
nor U3245 (N_3245,In_239,In_308);
nor U3246 (N_3246,In_1710,In_1756);
xnor U3247 (N_3247,In_391,In_965);
xnor U3248 (N_3248,In_708,In_1318);
xor U3249 (N_3249,In_1303,In_1286);
nor U3250 (N_3250,In_876,In_2365);
or U3251 (N_3251,In_1559,In_1774);
nand U3252 (N_3252,In_1607,In_2464);
or U3253 (N_3253,In_2020,In_1802);
nand U3254 (N_3254,In_1886,In_800);
or U3255 (N_3255,In_1688,In_1026);
nand U3256 (N_3256,In_760,In_1894);
and U3257 (N_3257,In_1124,In_1356);
nand U3258 (N_3258,In_446,In_1308);
xor U3259 (N_3259,In_1002,In_128);
nor U3260 (N_3260,In_153,In_1888);
xor U3261 (N_3261,In_2296,In_355);
nand U3262 (N_3262,In_140,In_1516);
nor U3263 (N_3263,In_1717,In_979);
nand U3264 (N_3264,In_1098,In_1345);
nand U3265 (N_3265,In_1611,In_267);
nor U3266 (N_3266,In_1784,In_1522);
nand U3267 (N_3267,In_1931,In_502);
and U3268 (N_3268,In_58,In_1240);
nor U3269 (N_3269,In_1586,In_2372);
or U3270 (N_3270,In_76,In_2040);
xnor U3271 (N_3271,In_592,In_1011);
nand U3272 (N_3272,In_283,In_1095);
xnor U3273 (N_3273,In_323,In_1036);
or U3274 (N_3274,In_1944,In_295);
xor U3275 (N_3275,In_1201,In_823);
and U3276 (N_3276,In_2264,In_1477);
and U3277 (N_3277,In_2056,In_322);
nand U3278 (N_3278,In_2251,In_2265);
and U3279 (N_3279,In_2496,In_537);
xnor U3280 (N_3280,In_443,In_147);
and U3281 (N_3281,In_2164,In_137);
nand U3282 (N_3282,In_1274,In_298);
or U3283 (N_3283,In_1665,In_2036);
nand U3284 (N_3284,In_1963,In_1195);
nand U3285 (N_3285,In_1657,In_552);
or U3286 (N_3286,In_2123,In_539);
or U3287 (N_3287,In_1892,In_1227);
and U3288 (N_3288,In_2496,In_2208);
nor U3289 (N_3289,In_2090,In_514);
or U3290 (N_3290,In_158,In_703);
xnor U3291 (N_3291,In_1686,In_1940);
or U3292 (N_3292,In_1120,In_1470);
nor U3293 (N_3293,In_239,In_2238);
or U3294 (N_3294,In_230,In_972);
or U3295 (N_3295,In_2342,In_479);
xnor U3296 (N_3296,In_369,In_1250);
nor U3297 (N_3297,In_586,In_1311);
xnor U3298 (N_3298,In_535,In_2311);
nand U3299 (N_3299,In_1925,In_1979);
nor U3300 (N_3300,In_413,In_2043);
and U3301 (N_3301,In_852,In_2359);
and U3302 (N_3302,In_999,In_128);
nand U3303 (N_3303,In_1944,In_2357);
and U3304 (N_3304,In_1751,In_2321);
and U3305 (N_3305,In_67,In_920);
nand U3306 (N_3306,In_2384,In_989);
nor U3307 (N_3307,In_375,In_561);
xor U3308 (N_3308,In_1688,In_393);
nor U3309 (N_3309,In_703,In_45);
nand U3310 (N_3310,In_1714,In_2375);
nor U3311 (N_3311,In_566,In_635);
nand U3312 (N_3312,In_1631,In_1664);
nor U3313 (N_3313,In_693,In_1077);
nand U3314 (N_3314,In_611,In_2257);
and U3315 (N_3315,In_1492,In_1821);
nor U3316 (N_3316,In_2303,In_1732);
or U3317 (N_3317,In_2120,In_313);
and U3318 (N_3318,In_2382,In_1717);
nand U3319 (N_3319,In_679,In_53);
xnor U3320 (N_3320,In_529,In_1874);
xor U3321 (N_3321,In_1107,In_1305);
nand U3322 (N_3322,In_1385,In_1920);
nand U3323 (N_3323,In_1658,In_838);
or U3324 (N_3324,In_1993,In_594);
and U3325 (N_3325,In_750,In_1640);
and U3326 (N_3326,In_1140,In_860);
and U3327 (N_3327,In_1841,In_534);
and U3328 (N_3328,In_490,In_2136);
nor U3329 (N_3329,In_1262,In_132);
nor U3330 (N_3330,In_2387,In_1084);
or U3331 (N_3331,In_1123,In_1278);
or U3332 (N_3332,In_168,In_2010);
and U3333 (N_3333,In_1927,In_198);
nand U3334 (N_3334,In_951,In_2008);
and U3335 (N_3335,In_1984,In_2048);
nor U3336 (N_3336,In_1398,In_528);
or U3337 (N_3337,In_2444,In_1841);
or U3338 (N_3338,In_2301,In_438);
and U3339 (N_3339,In_1441,In_1923);
nor U3340 (N_3340,In_1806,In_791);
nand U3341 (N_3341,In_1748,In_753);
or U3342 (N_3342,In_950,In_513);
nand U3343 (N_3343,In_256,In_1267);
or U3344 (N_3344,In_2367,In_1036);
or U3345 (N_3345,In_722,In_1386);
or U3346 (N_3346,In_2340,In_1544);
nor U3347 (N_3347,In_1160,In_351);
or U3348 (N_3348,In_745,In_908);
or U3349 (N_3349,In_470,In_1873);
nand U3350 (N_3350,In_463,In_198);
or U3351 (N_3351,In_1600,In_1788);
or U3352 (N_3352,In_1213,In_659);
xnor U3353 (N_3353,In_1228,In_1262);
and U3354 (N_3354,In_31,In_2216);
nand U3355 (N_3355,In_341,In_2284);
and U3356 (N_3356,In_825,In_1328);
or U3357 (N_3357,In_2404,In_2312);
nor U3358 (N_3358,In_1267,In_625);
or U3359 (N_3359,In_1836,In_773);
or U3360 (N_3360,In_1591,In_726);
xor U3361 (N_3361,In_2151,In_1985);
nor U3362 (N_3362,In_677,In_2128);
nor U3363 (N_3363,In_1786,In_2419);
nand U3364 (N_3364,In_94,In_608);
xnor U3365 (N_3365,In_1533,In_1163);
or U3366 (N_3366,In_1389,In_2425);
or U3367 (N_3367,In_3,In_1415);
and U3368 (N_3368,In_841,In_1642);
nor U3369 (N_3369,In_872,In_1479);
or U3370 (N_3370,In_1800,In_1656);
nor U3371 (N_3371,In_242,In_426);
or U3372 (N_3372,In_935,In_2335);
and U3373 (N_3373,In_1596,In_713);
or U3374 (N_3374,In_1596,In_1370);
nand U3375 (N_3375,In_1444,In_690);
or U3376 (N_3376,In_132,In_1178);
or U3377 (N_3377,In_1533,In_1603);
nor U3378 (N_3378,In_635,In_2177);
nand U3379 (N_3379,In_996,In_2499);
and U3380 (N_3380,In_1886,In_2131);
and U3381 (N_3381,In_548,In_2424);
nor U3382 (N_3382,In_40,In_2255);
or U3383 (N_3383,In_49,In_1431);
nand U3384 (N_3384,In_1035,In_334);
or U3385 (N_3385,In_378,In_611);
nand U3386 (N_3386,In_391,In_815);
nand U3387 (N_3387,In_2396,In_865);
or U3388 (N_3388,In_1807,In_2415);
nand U3389 (N_3389,In_2013,In_1618);
nor U3390 (N_3390,In_131,In_288);
nor U3391 (N_3391,In_804,In_74);
nand U3392 (N_3392,In_342,In_257);
or U3393 (N_3393,In_331,In_885);
and U3394 (N_3394,In_106,In_990);
and U3395 (N_3395,In_698,In_1621);
nand U3396 (N_3396,In_844,In_1653);
or U3397 (N_3397,In_88,In_75);
nand U3398 (N_3398,In_1152,In_281);
nand U3399 (N_3399,In_1012,In_1197);
xnor U3400 (N_3400,In_2290,In_772);
nand U3401 (N_3401,In_968,In_1110);
and U3402 (N_3402,In_2361,In_501);
nor U3403 (N_3403,In_794,In_978);
nand U3404 (N_3404,In_2091,In_286);
or U3405 (N_3405,In_673,In_50);
xor U3406 (N_3406,In_1962,In_764);
or U3407 (N_3407,In_2275,In_777);
or U3408 (N_3408,In_1885,In_1046);
nand U3409 (N_3409,In_873,In_1047);
or U3410 (N_3410,In_2261,In_1310);
nor U3411 (N_3411,In_637,In_2134);
nand U3412 (N_3412,In_34,In_1378);
or U3413 (N_3413,In_2236,In_604);
xnor U3414 (N_3414,In_877,In_1450);
nor U3415 (N_3415,In_1484,In_2063);
or U3416 (N_3416,In_1455,In_1402);
nand U3417 (N_3417,In_1177,In_773);
nor U3418 (N_3418,In_909,In_934);
or U3419 (N_3419,In_1264,In_2360);
nor U3420 (N_3420,In_890,In_1650);
nor U3421 (N_3421,In_1567,In_192);
and U3422 (N_3422,In_810,In_49);
xor U3423 (N_3423,In_2473,In_1950);
and U3424 (N_3424,In_132,In_716);
and U3425 (N_3425,In_1640,In_1371);
xnor U3426 (N_3426,In_2399,In_923);
or U3427 (N_3427,In_2350,In_1218);
or U3428 (N_3428,In_879,In_2461);
nand U3429 (N_3429,In_1316,In_1833);
and U3430 (N_3430,In_481,In_1860);
nor U3431 (N_3431,In_71,In_1233);
or U3432 (N_3432,In_2024,In_2175);
nor U3433 (N_3433,In_1306,In_1656);
nor U3434 (N_3434,In_1916,In_670);
and U3435 (N_3435,In_687,In_1436);
nand U3436 (N_3436,In_1161,In_998);
nor U3437 (N_3437,In_1138,In_287);
nand U3438 (N_3438,In_2138,In_1261);
nand U3439 (N_3439,In_1783,In_420);
and U3440 (N_3440,In_312,In_1344);
and U3441 (N_3441,In_1685,In_1782);
nor U3442 (N_3442,In_1947,In_2365);
nand U3443 (N_3443,In_1644,In_1969);
nand U3444 (N_3444,In_867,In_743);
nor U3445 (N_3445,In_57,In_593);
nor U3446 (N_3446,In_1545,In_662);
and U3447 (N_3447,In_986,In_2001);
and U3448 (N_3448,In_558,In_1256);
nand U3449 (N_3449,In_1496,In_198);
nand U3450 (N_3450,In_2192,In_2461);
nand U3451 (N_3451,In_425,In_1254);
nor U3452 (N_3452,In_1953,In_2380);
and U3453 (N_3453,In_2114,In_1694);
or U3454 (N_3454,In_1451,In_1486);
and U3455 (N_3455,In_1029,In_24);
nor U3456 (N_3456,In_2288,In_23);
nor U3457 (N_3457,In_1404,In_1616);
xnor U3458 (N_3458,In_1561,In_285);
and U3459 (N_3459,In_50,In_448);
nand U3460 (N_3460,In_154,In_1979);
nand U3461 (N_3461,In_698,In_640);
and U3462 (N_3462,In_692,In_177);
nand U3463 (N_3463,In_531,In_2010);
nor U3464 (N_3464,In_932,In_1457);
xor U3465 (N_3465,In_2485,In_1850);
or U3466 (N_3466,In_2137,In_1672);
and U3467 (N_3467,In_1063,In_169);
or U3468 (N_3468,In_2308,In_730);
nor U3469 (N_3469,In_695,In_1195);
and U3470 (N_3470,In_320,In_1922);
xnor U3471 (N_3471,In_139,In_494);
or U3472 (N_3472,In_2018,In_2437);
and U3473 (N_3473,In_243,In_1607);
nand U3474 (N_3474,In_837,In_2078);
and U3475 (N_3475,In_174,In_28);
nand U3476 (N_3476,In_959,In_2173);
nand U3477 (N_3477,In_107,In_2391);
nand U3478 (N_3478,In_1780,In_46);
and U3479 (N_3479,In_613,In_2402);
nand U3480 (N_3480,In_1244,In_450);
nor U3481 (N_3481,In_808,In_2333);
nand U3482 (N_3482,In_2192,In_1524);
and U3483 (N_3483,In_850,In_1164);
nor U3484 (N_3484,In_2002,In_1568);
nand U3485 (N_3485,In_650,In_2233);
or U3486 (N_3486,In_737,In_758);
or U3487 (N_3487,In_166,In_2449);
nor U3488 (N_3488,In_100,In_1554);
and U3489 (N_3489,In_1128,In_2237);
xor U3490 (N_3490,In_802,In_1797);
xnor U3491 (N_3491,In_278,In_1095);
or U3492 (N_3492,In_1160,In_1643);
nor U3493 (N_3493,In_2351,In_1517);
nor U3494 (N_3494,In_1256,In_1032);
nand U3495 (N_3495,In_403,In_1140);
nand U3496 (N_3496,In_1963,In_1421);
and U3497 (N_3497,In_1687,In_1197);
or U3498 (N_3498,In_91,In_555);
nand U3499 (N_3499,In_2058,In_689);
and U3500 (N_3500,In_2192,In_503);
nand U3501 (N_3501,In_2219,In_1867);
or U3502 (N_3502,In_2129,In_1044);
nor U3503 (N_3503,In_924,In_1680);
nand U3504 (N_3504,In_549,In_890);
xnor U3505 (N_3505,In_956,In_2469);
nand U3506 (N_3506,In_1998,In_971);
or U3507 (N_3507,In_300,In_253);
nor U3508 (N_3508,In_780,In_300);
xor U3509 (N_3509,In_2001,In_1221);
nand U3510 (N_3510,In_347,In_2108);
xor U3511 (N_3511,In_1912,In_1603);
nor U3512 (N_3512,In_1841,In_1289);
nor U3513 (N_3513,In_2282,In_1339);
xnor U3514 (N_3514,In_2020,In_913);
or U3515 (N_3515,In_761,In_154);
or U3516 (N_3516,In_863,In_618);
xor U3517 (N_3517,In_219,In_1717);
and U3518 (N_3518,In_1395,In_15);
xor U3519 (N_3519,In_2108,In_1156);
nand U3520 (N_3520,In_1153,In_44);
or U3521 (N_3521,In_2315,In_1022);
and U3522 (N_3522,In_1784,In_1465);
or U3523 (N_3523,In_1684,In_1419);
and U3524 (N_3524,In_2485,In_1919);
and U3525 (N_3525,In_254,In_1366);
nand U3526 (N_3526,In_1298,In_2184);
and U3527 (N_3527,In_1805,In_1167);
or U3528 (N_3528,In_614,In_400);
and U3529 (N_3529,In_1470,In_1688);
nand U3530 (N_3530,In_1583,In_447);
nand U3531 (N_3531,In_1762,In_1048);
and U3532 (N_3532,In_658,In_2458);
or U3533 (N_3533,In_1417,In_100);
or U3534 (N_3534,In_2356,In_255);
nand U3535 (N_3535,In_818,In_129);
nor U3536 (N_3536,In_2262,In_307);
and U3537 (N_3537,In_304,In_651);
nand U3538 (N_3538,In_1765,In_597);
nand U3539 (N_3539,In_1628,In_2071);
nand U3540 (N_3540,In_1324,In_2146);
nand U3541 (N_3541,In_50,In_495);
xor U3542 (N_3542,In_399,In_995);
nand U3543 (N_3543,In_2470,In_2360);
nand U3544 (N_3544,In_300,In_530);
nor U3545 (N_3545,In_1289,In_714);
xor U3546 (N_3546,In_221,In_506);
and U3547 (N_3547,In_2179,In_1155);
xor U3548 (N_3548,In_250,In_1643);
xor U3549 (N_3549,In_2211,In_1866);
nand U3550 (N_3550,In_1580,In_1279);
nor U3551 (N_3551,In_722,In_1876);
nor U3552 (N_3552,In_1979,In_1472);
nor U3553 (N_3553,In_427,In_2177);
nor U3554 (N_3554,In_546,In_607);
and U3555 (N_3555,In_2468,In_927);
or U3556 (N_3556,In_906,In_587);
or U3557 (N_3557,In_83,In_1381);
nand U3558 (N_3558,In_311,In_703);
and U3559 (N_3559,In_955,In_252);
nor U3560 (N_3560,In_340,In_170);
nor U3561 (N_3561,In_1976,In_1272);
or U3562 (N_3562,In_1660,In_1894);
nor U3563 (N_3563,In_2482,In_2471);
nor U3564 (N_3564,In_1462,In_505);
and U3565 (N_3565,In_1067,In_2486);
or U3566 (N_3566,In_1469,In_1911);
or U3567 (N_3567,In_1525,In_1166);
xnor U3568 (N_3568,In_433,In_2055);
nor U3569 (N_3569,In_371,In_2364);
or U3570 (N_3570,In_1334,In_259);
or U3571 (N_3571,In_261,In_1735);
nor U3572 (N_3572,In_373,In_1763);
and U3573 (N_3573,In_2494,In_1255);
xor U3574 (N_3574,In_550,In_535);
xnor U3575 (N_3575,In_1089,In_1213);
xor U3576 (N_3576,In_100,In_1434);
and U3577 (N_3577,In_2406,In_958);
nor U3578 (N_3578,In_1103,In_1106);
xor U3579 (N_3579,In_1912,In_1498);
or U3580 (N_3580,In_80,In_149);
nand U3581 (N_3581,In_1291,In_1698);
and U3582 (N_3582,In_750,In_124);
nor U3583 (N_3583,In_1480,In_2495);
nor U3584 (N_3584,In_1915,In_1408);
and U3585 (N_3585,In_1330,In_824);
nand U3586 (N_3586,In_1614,In_2211);
nand U3587 (N_3587,In_1958,In_1932);
nand U3588 (N_3588,In_469,In_1950);
nor U3589 (N_3589,In_2455,In_1749);
and U3590 (N_3590,In_469,In_1672);
nor U3591 (N_3591,In_2347,In_2488);
nand U3592 (N_3592,In_1044,In_1921);
xor U3593 (N_3593,In_1021,In_148);
nand U3594 (N_3594,In_1192,In_76);
nor U3595 (N_3595,In_1210,In_1246);
or U3596 (N_3596,In_1163,In_6);
nor U3597 (N_3597,In_2350,In_2403);
or U3598 (N_3598,In_314,In_1027);
or U3599 (N_3599,In_866,In_2222);
or U3600 (N_3600,In_809,In_1664);
nor U3601 (N_3601,In_136,In_1432);
xor U3602 (N_3602,In_2006,In_24);
or U3603 (N_3603,In_847,In_596);
nand U3604 (N_3604,In_653,In_2174);
nand U3605 (N_3605,In_1396,In_2026);
and U3606 (N_3606,In_971,In_323);
or U3607 (N_3607,In_1135,In_2117);
nand U3608 (N_3608,In_1419,In_1305);
and U3609 (N_3609,In_996,In_185);
nor U3610 (N_3610,In_450,In_1166);
nand U3611 (N_3611,In_1010,In_72);
nor U3612 (N_3612,In_870,In_735);
or U3613 (N_3613,In_2302,In_1455);
and U3614 (N_3614,In_495,In_2364);
xnor U3615 (N_3615,In_1276,In_1673);
or U3616 (N_3616,In_613,In_721);
nand U3617 (N_3617,In_899,In_262);
nand U3618 (N_3618,In_1793,In_995);
nor U3619 (N_3619,In_299,In_688);
xor U3620 (N_3620,In_1262,In_1149);
xnor U3621 (N_3621,In_1234,In_1385);
nand U3622 (N_3622,In_1535,In_622);
nand U3623 (N_3623,In_383,In_1968);
xnor U3624 (N_3624,In_542,In_1172);
and U3625 (N_3625,In_1938,In_1762);
or U3626 (N_3626,In_289,In_544);
nor U3627 (N_3627,In_217,In_1063);
nor U3628 (N_3628,In_1898,In_1603);
or U3629 (N_3629,In_189,In_1441);
and U3630 (N_3630,In_1996,In_1679);
nor U3631 (N_3631,In_2076,In_1115);
nor U3632 (N_3632,In_574,In_2125);
nand U3633 (N_3633,In_972,In_1217);
or U3634 (N_3634,In_2426,In_1789);
xor U3635 (N_3635,In_96,In_2355);
and U3636 (N_3636,In_438,In_356);
nor U3637 (N_3637,In_1594,In_2349);
or U3638 (N_3638,In_1463,In_1244);
xnor U3639 (N_3639,In_406,In_680);
or U3640 (N_3640,In_1091,In_2116);
and U3641 (N_3641,In_2069,In_95);
or U3642 (N_3642,In_2353,In_992);
and U3643 (N_3643,In_2382,In_1081);
xnor U3644 (N_3644,In_2274,In_1002);
and U3645 (N_3645,In_739,In_744);
nor U3646 (N_3646,In_1733,In_1555);
nor U3647 (N_3647,In_30,In_1136);
xnor U3648 (N_3648,In_2439,In_86);
and U3649 (N_3649,In_1404,In_438);
or U3650 (N_3650,In_2101,In_1964);
and U3651 (N_3651,In_624,In_814);
nand U3652 (N_3652,In_1772,In_1154);
nand U3653 (N_3653,In_452,In_2397);
and U3654 (N_3654,In_605,In_1860);
and U3655 (N_3655,In_1917,In_273);
or U3656 (N_3656,In_399,In_205);
nor U3657 (N_3657,In_385,In_906);
and U3658 (N_3658,In_675,In_1858);
xnor U3659 (N_3659,In_1006,In_1492);
nand U3660 (N_3660,In_313,In_2492);
nor U3661 (N_3661,In_1537,In_2112);
and U3662 (N_3662,In_2465,In_2170);
nand U3663 (N_3663,In_1756,In_2451);
xor U3664 (N_3664,In_1846,In_2172);
nand U3665 (N_3665,In_1660,In_554);
and U3666 (N_3666,In_1621,In_1672);
or U3667 (N_3667,In_545,In_1022);
or U3668 (N_3668,In_1407,In_2415);
and U3669 (N_3669,In_2220,In_2236);
nand U3670 (N_3670,In_1020,In_1070);
nand U3671 (N_3671,In_1541,In_659);
and U3672 (N_3672,In_674,In_1393);
and U3673 (N_3673,In_2266,In_831);
nor U3674 (N_3674,In_1472,In_1905);
nand U3675 (N_3675,In_2087,In_2473);
and U3676 (N_3676,In_1678,In_194);
or U3677 (N_3677,In_2052,In_152);
or U3678 (N_3678,In_2465,In_1480);
xnor U3679 (N_3679,In_685,In_1465);
nor U3680 (N_3680,In_1461,In_356);
or U3681 (N_3681,In_1793,In_1418);
nor U3682 (N_3682,In_296,In_80);
nor U3683 (N_3683,In_2195,In_2121);
or U3684 (N_3684,In_1195,In_1317);
and U3685 (N_3685,In_364,In_1198);
nor U3686 (N_3686,In_1192,In_1617);
xnor U3687 (N_3687,In_1506,In_155);
or U3688 (N_3688,In_1777,In_2419);
or U3689 (N_3689,In_1267,In_2344);
or U3690 (N_3690,In_1227,In_1548);
and U3691 (N_3691,In_2193,In_1048);
and U3692 (N_3692,In_758,In_727);
and U3693 (N_3693,In_1512,In_1104);
xor U3694 (N_3694,In_1730,In_56);
nand U3695 (N_3695,In_784,In_1930);
or U3696 (N_3696,In_1539,In_1780);
and U3697 (N_3697,In_372,In_175);
and U3698 (N_3698,In_1441,In_2074);
nand U3699 (N_3699,In_2215,In_1604);
nand U3700 (N_3700,In_2276,In_206);
nand U3701 (N_3701,In_570,In_1261);
nand U3702 (N_3702,In_1391,In_1418);
and U3703 (N_3703,In_2250,In_2338);
nand U3704 (N_3704,In_1035,In_182);
and U3705 (N_3705,In_1753,In_1136);
nand U3706 (N_3706,In_1719,In_182);
or U3707 (N_3707,In_1087,In_1273);
and U3708 (N_3708,In_2085,In_1220);
nor U3709 (N_3709,In_2283,In_1321);
xor U3710 (N_3710,In_1680,In_317);
xor U3711 (N_3711,In_1708,In_149);
nand U3712 (N_3712,In_33,In_1115);
or U3713 (N_3713,In_419,In_1040);
nand U3714 (N_3714,In_2475,In_1319);
or U3715 (N_3715,In_756,In_1295);
nand U3716 (N_3716,In_483,In_589);
and U3717 (N_3717,In_2060,In_2156);
and U3718 (N_3718,In_2031,In_192);
or U3719 (N_3719,In_1148,In_384);
and U3720 (N_3720,In_1956,In_2227);
nor U3721 (N_3721,In_2325,In_1003);
and U3722 (N_3722,In_95,In_759);
or U3723 (N_3723,In_1592,In_1844);
nand U3724 (N_3724,In_1452,In_1434);
nand U3725 (N_3725,In_1375,In_708);
and U3726 (N_3726,In_856,In_1037);
and U3727 (N_3727,In_1102,In_986);
nor U3728 (N_3728,In_586,In_1121);
xnor U3729 (N_3729,In_2406,In_134);
and U3730 (N_3730,In_75,In_1878);
xnor U3731 (N_3731,In_1126,In_21);
xnor U3732 (N_3732,In_1324,In_974);
and U3733 (N_3733,In_939,In_806);
nor U3734 (N_3734,In_56,In_570);
nor U3735 (N_3735,In_970,In_1657);
or U3736 (N_3736,In_357,In_904);
or U3737 (N_3737,In_1913,In_2421);
or U3738 (N_3738,In_17,In_1670);
nor U3739 (N_3739,In_1886,In_2240);
nand U3740 (N_3740,In_742,In_368);
nand U3741 (N_3741,In_984,In_2459);
or U3742 (N_3742,In_1521,In_927);
and U3743 (N_3743,In_931,In_2323);
nand U3744 (N_3744,In_494,In_1598);
nor U3745 (N_3745,In_66,In_1369);
nor U3746 (N_3746,In_2485,In_967);
or U3747 (N_3747,In_1747,In_849);
or U3748 (N_3748,In_1328,In_832);
nand U3749 (N_3749,In_2479,In_978);
nand U3750 (N_3750,In_2001,In_1098);
nand U3751 (N_3751,In_1580,In_1798);
nor U3752 (N_3752,In_469,In_1555);
nor U3753 (N_3753,In_909,In_599);
or U3754 (N_3754,In_2240,In_793);
and U3755 (N_3755,In_878,In_1676);
nand U3756 (N_3756,In_287,In_1459);
nor U3757 (N_3757,In_1493,In_1109);
and U3758 (N_3758,In_165,In_1987);
nand U3759 (N_3759,In_2224,In_2172);
and U3760 (N_3760,In_1953,In_848);
and U3761 (N_3761,In_103,In_1856);
or U3762 (N_3762,In_2307,In_672);
nor U3763 (N_3763,In_188,In_1542);
xnor U3764 (N_3764,In_1088,In_1933);
nor U3765 (N_3765,In_761,In_1103);
or U3766 (N_3766,In_1032,In_2214);
nor U3767 (N_3767,In_542,In_159);
nor U3768 (N_3768,In_1124,In_1369);
and U3769 (N_3769,In_916,In_1189);
nor U3770 (N_3770,In_44,In_1837);
nor U3771 (N_3771,In_1209,In_434);
nand U3772 (N_3772,In_1428,In_1956);
or U3773 (N_3773,In_1860,In_1066);
or U3774 (N_3774,In_205,In_990);
nor U3775 (N_3775,In_1280,In_975);
and U3776 (N_3776,In_388,In_424);
or U3777 (N_3777,In_1521,In_1924);
and U3778 (N_3778,In_297,In_2228);
nand U3779 (N_3779,In_63,In_2308);
or U3780 (N_3780,In_1042,In_1305);
and U3781 (N_3781,In_1150,In_1228);
nand U3782 (N_3782,In_1310,In_129);
and U3783 (N_3783,In_2115,In_1500);
or U3784 (N_3784,In_684,In_1110);
xor U3785 (N_3785,In_308,In_1049);
and U3786 (N_3786,In_1165,In_861);
nor U3787 (N_3787,In_1310,In_1370);
or U3788 (N_3788,In_487,In_1611);
nor U3789 (N_3789,In_1429,In_266);
or U3790 (N_3790,In_1452,In_1533);
nand U3791 (N_3791,In_1525,In_476);
nor U3792 (N_3792,In_1539,In_1812);
xor U3793 (N_3793,In_999,In_885);
and U3794 (N_3794,In_2400,In_391);
nand U3795 (N_3795,In_1063,In_1087);
or U3796 (N_3796,In_2168,In_1610);
and U3797 (N_3797,In_455,In_173);
nor U3798 (N_3798,In_1180,In_2115);
nand U3799 (N_3799,In_1864,In_2109);
nor U3800 (N_3800,In_1363,In_967);
nand U3801 (N_3801,In_1796,In_1552);
and U3802 (N_3802,In_2202,In_2386);
and U3803 (N_3803,In_1979,In_1606);
nand U3804 (N_3804,In_2087,In_2332);
nand U3805 (N_3805,In_2285,In_123);
nor U3806 (N_3806,In_962,In_1590);
nor U3807 (N_3807,In_470,In_1979);
nor U3808 (N_3808,In_681,In_1080);
nand U3809 (N_3809,In_2167,In_25);
or U3810 (N_3810,In_78,In_1324);
nand U3811 (N_3811,In_2067,In_691);
nor U3812 (N_3812,In_908,In_2264);
or U3813 (N_3813,In_2449,In_1243);
nor U3814 (N_3814,In_50,In_537);
or U3815 (N_3815,In_1427,In_937);
and U3816 (N_3816,In_756,In_1623);
or U3817 (N_3817,In_2147,In_1161);
and U3818 (N_3818,In_857,In_1153);
nand U3819 (N_3819,In_1290,In_1503);
and U3820 (N_3820,In_1506,In_673);
nor U3821 (N_3821,In_2022,In_730);
and U3822 (N_3822,In_206,In_1949);
nand U3823 (N_3823,In_1057,In_2071);
or U3824 (N_3824,In_1683,In_2325);
nand U3825 (N_3825,In_1358,In_1877);
nor U3826 (N_3826,In_2044,In_1327);
nand U3827 (N_3827,In_2389,In_826);
and U3828 (N_3828,In_987,In_191);
nand U3829 (N_3829,In_1427,In_781);
or U3830 (N_3830,In_954,In_1974);
nand U3831 (N_3831,In_1092,In_1074);
nor U3832 (N_3832,In_269,In_1419);
or U3833 (N_3833,In_665,In_618);
and U3834 (N_3834,In_2197,In_1774);
nand U3835 (N_3835,In_1901,In_457);
xnor U3836 (N_3836,In_1593,In_451);
nor U3837 (N_3837,In_207,In_2476);
nand U3838 (N_3838,In_2408,In_1800);
nor U3839 (N_3839,In_1995,In_663);
or U3840 (N_3840,In_2334,In_226);
and U3841 (N_3841,In_420,In_2106);
or U3842 (N_3842,In_233,In_1253);
and U3843 (N_3843,In_2234,In_536);
or U3844 (N_3844,In_463,In_1196);
or U3845 (N_3845,In_2174,In_755);
and U3846 (N_3846,In_58,In_723);
nor U3847 (N_3847,In_148,In_1638);
nor U3848 (N_3848,In_1486,In_465);
xor U3849 (N_3849,In_116,In_135);
and U3850 (N_3850,In_1933,In_1773);
nor U3851 (N_3851,In_1794,In_686);
and U3852 (N_3852,In_2210,In_991);
or U3853 (N_3853,In_2474,In_1260);
nand U3854 (N_3854,In_304,In_2244);
nand U3855 (N_3855,In_1082,In_350);
nor U3856 (N_3856,In_2417,In_631);
nor U3857 (N_3857,In_2125,In_1577);
or U3858 (N_3858,In_1971,In_2052);
nor U3859 (N_3859,In_1192,In_2058);
or U3860 (N_3860,In_828,In_1710);
xnor U3861 (N_3861,In_933,In_1348);
nor U3862 (N_3862,In_1978,In_1896);
nand U3863 (N_3863,In_1867,In_14);
and U3864 (N_3864,In_1148,In_2151);
or U3865 (N_3865,In_780,In_2224);
nand U3866 (N_3866,In_1511,In_1384);
nor U3867 (N_3867,In_424,In_837);
or U3868 (N_3868,In_707,In_1089);
nor U3869 (N_3869,In_327,In_580);
and U3870 (N_3870,In_216,In_1860);
xnor U3871 (N_3871,In_2032,In_2214);
or U3872 (N_3872,In_2155,In_487);
and U3873 (N_3873,In_544,In_1102);
nand U3874 (N_3874,In_2064,In_2024);
and U3875 (N_3875,In_2053,In_1140);
nor U3876 (N_3876,In_334,In_364);
nor U3877 (N_3877,In_262,In_1475);
and U3878 (N_3878,In_2478,In_2056);
and U3879 (N_3879,In_1829,In_2152);
and U3880 (N_3880,In_2363,In_1614);
or U3881 (N_3881,In_2030,In_530);
or U3882 (N_3882,In_1712,In_71);
or U3883 (N_3883,In_324,In_1533);
nor U3884 (N_3884,In_403,In_1595);
nor U3885 (N_3885,In_2230,In_2057);
and U3886 (N_3886,In_1568,In_1452);
or U3887 (N_3887,In_674,In_401);
or U3888 (N_3888,In_1852,In_1561);
nand U3889 (N_3889,In_1327,In_937);
nand U3890 (N_3890,In_824,In_2259);
or U3891 (N_3891,In_1910,In_172);
nand U3892 (N_3892,In_997,In_1410);
or U3893 (N_3893,In_778,In_699);
nand U3894 (N_3894,In_2041,In_870);
and U3895 (N_3895,In_2085,In_2495);
nor U3896 (N_3896,In_1892,In_223);
nand U3897 (N_3897,In_2003,In_545);
and U3898 (N_3898,In_1616,In_1721);
and U3899 (N_3899,In_535,In_1854);
nand U3900 (N_3900,In_1509,In_905);
nor U3901 (N_3901,In_2347,In_723);
xor U3902 (N_3902,In_1834,In_644);
and U3903 (N_3903,In_866,In_1318);
nand U3904 (N_3904,In_2144,In_1191);
and U3905 (N_3905,In_2237,In_1365);
nand U3906 (N_3906,In_2264,In_1049);
and U3907 (N_3907,In_834,In_845);
or U3908 (N_3908,In_2141,In_1392);
nor U3909 (N_3909,In_454,In_1399);
or U3910 (N_3910,In_807,In_2100);
and U3911 (N_3911,In_2065,In_73);
and U3912 (N_3912,In_1772,In_2347);
and U3913 (N_3913,In_118,In_968);
xor U3914 (N_3914,In_1710,In_377);
nand U3915 (N_3915,In_925,In_345);
xor U3916 (N_3916,In_1783,In_1461);
nor U3917 (N_3917,In_2362,In_2123);
nand U3918 (N_3918,In_988,In_1554);
or U3919 (N_3919,In_1812,In_1523);
nand U3920 (N_3920,In_2242,In_529);
nand U3921 (N_3921,In_593,In_772);
nand U3922 (N_3922,In_1370,In_1545);
xor U3923 (N_3923,In_2267,In_44);
nand U3924 (N_3924,In_1926,In_1299);
nor U3925 (N_3925,In_102,In_2428);
or U3926 (N_3926,In_533,In_1914);
xor U3927 (N_3927,In_2273,In_899);
or U3928 (N_3928,In_475,In_2022);
nand U3929 (N_3929,In_217,In_1185);
or U3930 (N_3930,In_2150,In_605);
and U3931 (N_3931,In_976,In_2068);
or U3932 (N_3932,In_86,In_1234);
nor U3933 (N_3933,In_548,In_1028);
or U3934 (N_3934,In_2091,In_2276);
nor U3935 (N_3935,In_177,In_333);
nor U3936 (N_3936,In_1554,In_1494);
and U3937 (N_3937,In_1378,In_1429);
or U3938 (N_3938,In_31,In_1500);
or U3939 (N_3939,In_1501,In_1121);
or U3940 (N_3940,In_1091,In_888);
nor U3941 (N_3941,In_1632,In_78);
nand U3942 (N_3942,In_1679,In_2147);
nor U3943 (N_3943,In_1486,In_313);
and U3944 (N_3944,In_733,In_953);
nor U3945 (N_3945,In_1635,In_2406);
and U3946 (N_3946,In_2,In_2017);
nand U3947 (N_3947,In_1440,In_1990);
and U3948 (N_3948,In_952,In_1663);
or U3949 (N_3949,In_1360,In_639);
xor U3950 (N_3950,In_1891,In_335);
nand U3951 (N_3951,In_1333,In_332);
nand U3952 (N_3952,In_2093,In_949);
and U3953 (N_3953,In_870,In_851);
nand U3954 (N_3954,In_60,In_479);
and U3955 (N_3955,In_945,In_2088);
nand U3956 (N_3956,In_290,In_734);
nor U3957 (N_3957,In_1814,In_171);
or U3958 (N_3958,In_127,In_2020);
and U3959 (N_3959,In_1060,In_451);
nor U3960 (N_3960,In_2330,In_132);
or U3961 (N_3961,In_1284,In_558);
xor U3962 (N_3962,In_197,In_1507);
nand U3963 (N_3963,In_38,In_740);
nand U3964 (N_3964,In_1232,In_865);
nor U3965 (N_3965,In_605,In_954);
nor U3966 (N_3966,In_336,In_428);
xor U3967 (N_3967,In_2024,In_940);
nor U3968 (N_3968,In_2470,In_47);
nor U3969 (N_3969,In_627,In_646);
nand U3970 (N_3970,In_1825,In_1198);
nand U3971 (N_3971,In_782,In_381);
nand U3972 (N_3972,In_1208,In_2099);
xor U3973 (N_3973,In_81,In_1897);
nor U3974 (N_3974,In_84,In_2354);
and U3975 (N_3975,In_995,In_355);
xor U3976 (N_3976,In_1248,In_818);
and U3977 (N_3977,In_456,In_1137);
nor U3978 (N_3978,In_881,In_1199);
and U3979 (N_3979,In_1024,In_711);
nor U3980 (N_3980,In_1515,In_1035);
and U3981 (N_3981,In_124,In_918);
nor U3982 (N_3982,In_2354,In_2479);
nor U3983 (N_3983,In_439,In_2065);
nand U3984 (N_3984,In_2049,In_411);
nand U3985 (N_3985,In_718,In_2418);
nand U3986 (N_3986,In_1035,In_1265);
nor U3987 (N_3987,In_688,In_187);
nand U3988 (N_3988,In_775,In_2227);
or U3989 (N_3989,In_2231,In_1412);
nor U3990 (N_3990,In_1447,In_666);
nand U3991 (N_3991,In_1992,In_1372);
nor U3992 (N_3992,In_2056,In_1303);
and U3993 (N_3993,In_1436,In_1258);
and U3994 (N_3994,In_1370,In_1582);
nor U3995 (N_3995,In_1272,In_772);
nor U3996 (N_3996,In_1453,In_237);
and U3997 (N_3997,In_854,In_802);
and U3998 (N_3998,In_1542,In_466);
and U3999 (N_3999,In_1664,In_823);
nand U4000 (N_4000,In_1195,In_591);
nand U4001 (N_4001,In_799,In_1123);
nand U4002 (N_4002,In_792,In_1327);
xor U4003 (N_4003,In_1,In_1248);
nor U4004 (N_4004,In_1456,In_1007);
or U4005 (N_4005,In_497,In_1433);
nand U4006 (N_4006,In_1191,In_217);
and U4007 (N_4007,In_1681,In_671);
or U4008 (N_4008,In_1347,In_1152);
or U4009 (N_4009,In_1993,In_2202);
nor U4010 (N_4010,In_1607,In_398);
or U4011 (N_4011,In_57,In_40);
or U4012 (N_4012,In_816,In_481);
nor U4013 (N_4013,In_466,In_1574);
or U4014 (N_4014,In_1563,In_2180);
nor U4015 (N_4015,In_1751,In_1742);
or U4016 (N_4016,In_1612,In_1013);
and U4017 (N_4017,In_1278,In_752);
nand U4018 (N_4018,In_1816,In_2372);
and U4019 (N_4019,In_822,In_727);
xor U4020 (N_4020,In_679,In_1605);
xor U4021 (N_4021,In_1013,In_588);
and U4022 (N_4022,In_1321,In_1051);
or U4023 (N_4023,In_1229,In_515);
and U4024 (N_4024,In_2011,In_369);
and U4025 (N_4025,In_2461,In_504);
and U4026 (N_4026,In_447,In_2282);
nand U4027 (N_4027,In_1166,In_660);
and U4028 (N_4028,In_1504,In_1256);
and U4029 (N_4029,In_2284,In_203);
nand U4030 (N_4030,In_1423,In_578);
nand U4031 (N_4031,In_351,In_246);
nor U4032 (N_4032,In_626,In_1971);
and U4033 (N_4033,In_134,In_1824);
and U4034 (N_4034,In_1280,In_2151);
nand U4035 (N_4035,In_536,In_1885);
nand U4036 (N_4036,In_548,In_1289);
nor U4037 (N_4037,In_1623,In_531);
nor U4038 (N_4038,In_1185,In_1133);
or U4039 (N_4039,In_1749,In_618);
xnor U4040 (N_4040,In_822,In_79);
nor U4041 (N_4041,In_2305,In_763);
and U4042 (N_4042,In_1054,In_296);
and U4043 (N_4043,In_1296,In_1705);
nor U4044 (N_4044,In_1227,In_829);
nand U4045 (N_4045,In_1859,In_1297);
nor U4046 (N_4046,In_918,In_1668);
or U4047 (N_4047,In_2289,In_1212);
nand U4048 (N_4048,In_534,In_326);
or U4049 (N_4049,In_2228,In_103);
xnor U4050 (N_4050,In_117,In_2320);
nor U4051 (N_4051,In_118,In_2343);
nor U4052 (N_4052,In_1681,In_501);
nor U4053 (N_4053,In_373,In_1242);
nand U4054 (N_4054,In_17,In_753);
or U4055 (N_4055,In_2057,In_1274);
or U4056 (N_4056,In_2106,In_999);
xor U4057 (N_4057,In_1794,In_340);
and U4058 (N_4058,In_1257,In_253);
or U4059 (N_4059,In_202,In_847);
nor U4060 (N_4060,In_1821,In_300);
and U4061 (N_4061,In_2461,In_182);
or U4062 (N_4062,In_1586,In_1322);
nor U4063 (N_4063,In_1696,In_597);
nor U4064 (N_4064,In_243,In_1765);
nand U4065 (N_4065,In_617,In_23);
or U4066 (N_4066,In_1062,In_2085);
nand U4067 (N_4067,In_2176,In_1620);
or U4068 (N_4068,In_248,In_429);
xor U4069 (N_4069,In_486,In_677);
or U4070 (N_4070,In_498,In_1471);
and U4071 (N_4071,In_1009,In_1098);
nand U4072 (N_4072,In_1667,In_2004);
xnor U4073 (N_4073,In_1197,In_726);
nor U4074 (N_4074,In_1367,In_1698);
or U4075 (N_4075,In_1046,In_2169);
xnor U4076 (N_4076,In_2425,In_191);
or U4077 (N_4077,In_273,In_1874);
xnor U4078 (N_4078,In_1421,In_1348);
or U4079 (N_4079,In_1284,In_203);
nor U4080 (N_4080,In_395,In_1065);
nor U4081 (N_4081,In_1059,In_1574);
or U4082 (N_4082,In_1306,In_130);
and U4083 (N_4083,In_1187,In_1002);
or U4084 (N_4084,In_1673,In_53);
or U4085 (N_4085,In_2303,In_1777);
nand U4086 (N_4086,In_1164,In_1961);
nor U4087 (N_4087,In_1611,In_2222);
nand U4088 (N_4088,In_351,In_859);
or U4089 (N_4089,In_201,In_1140);
and U4090 (N_4090,In_2223,In_2383);
nor U4091 (N_4091,In_1098,In_838);
xnor U4092 (N_4092,In_1338,In_1444);
or U4093 (N_4093,In_580,In_1446);
nand U4094 (N_4094,In_1026,In_702);
nand U4095 (N_4095,In_1104,In_2284);
and U4096 (N_4096,In_925,In_2157);
or U4097 (N_4097,In_688,In_403);
nor U4098 (N_4098,In_601,In_1801);
and U4099 (N_4099,In_2460,In_984);
nor U4100 (N_4100,In_1435,In_981);
and U4101 (N_4101,In_1510,In_625);
nor U4102 (N_4102,In_2282,In_77);
nand U4103 (N_4103,In_494,In_670);
and U4104 (N_4104,In_1319,In_305);
or U4105 (N_4105,In_2473,In_601);
nand U4106 (N_4106,In_527,In_2201);
or U4107 (N_4107,In_2108,In_1972);
or U4108 (N_4108,In_1241,In_2233);
and U4109 (N_4109,In_2089,In_856);
and U4110 (N_4110,In_1510,In_1062);
nand U4111 (N_4111,In_175,In_168);
or U4112 (N_4112,In_1923,In_316);
or U4113 (N_4113,In_2354,In_1246);
and U4114 (N_4114,In_1265,In_2109);
nand U4115 (N_4115,In_127,In_1442);
and U4116 (N_4116,In_1067,In_605);
or U4117 (N_4117,In_1898,In_1097);
xor U4118 (N_4118,In_1962,In_518);
nor U4119 (N_4119,In_284,In_1300);
xnor U4120 (N_4120,In_948,In_1546);
and U4121 (N_4121,In_1853,In_1734);
nand U4122 (N_4122,In_104,In_446);
nand U4123 (N_4123,In_2356,In_1052);
nor U4124 (N_4124,In_1672,In_50);
nor U4125 (N_4125,In_513,In_1769);
nor U4126 (N_4126,In_473,In_505);
or U4127 (N_4127,In_594,In_890);
or U4128 (N_4128,In_1729,In_427);
nor U4129 (N_4129,In_891,In_2336);
and U4130 (N_4130,In_1465,In_1082);
nand U4131 (N_4131,In_1055,In_1676);
xnor U4132 (N_4132,In_336,In_834);
and U4133 (N_4133,In_646,In_31);
or U4134 (N_4134,In_2444,In_1928);
nor U4135 (N_4135,In_1265,In_1588);
nand U4136 (N_4136,In_247,In_1297);
or U4137 (N_4137,In_2138,In_393);
nand U4138 (N_4138,In_48,In_1658);
xor U4139 (N_4139,In_2042,In_1903);
or U4140 (N_4140,In_2462,In_1075);
or U4141 (N_4141,In_1229,In_2357);
or U4142 (N_4142,In_202,In_498);
or U4143 (N_4143,In_891,In_2090);
and U4144 (N_4144,In_2339,In_2246);
nand U4145 (N_4145,In_1269,In_2329);
or U4146 (N_4146,In_1349,In_31);
nand U4147 (N_4147,In_1918,In_325);
nor U4148 (N_4148,In_1593,In_1999);
nor U4149 (N_4149,In_595,In_815);
nand U4150 (N_4150,In_745,In_672);
nand U4151 (N_4151,In_1376,In_1184);
or U4152 (N_4152,In_387,In_574);
and U4153 (N_4153,In_893,In_1429);
xor U4154 (N_4154,In_488,In_47);
or U4155 (N_4155,In_2227,In_545);
nor U4156 (N_4156,In_1145,In_401);
nor U4157 (N_4157,In_1347,In_117);
nor U4158 (N_4158,In_25,In_1419);
or U4159 (N_4159,In_1915,In_1054);
or U4160 (N_4160,In_1457,In_1326);
nor U4161 (N_4161,In_1242,In_2112);
nor U4162 (N_4162,In_2485,In_344);
nand U4163 (N_4163,In_2482,In_2111);
or U4164 (N_4164,In_1153,In_445);
nand U4165 (N_4165,In_475,In_197);
and U4166 (N_4166,In_1918,In_1125);
nand U4167 (N_4167,In_422,In_901);
and U4168 (N_4168,In_2397,In_1614);
nand U4169 (N_4169,In_1789,In_1948);
and U4170 (N_4170,In_970,In_2208);
nor U4171 (N_4171,In_1579,In_820);
nand U4172 (N_4172,In_1862,In_1049);
nor U4173 (N_4173,In_934,In_1804);
or U4174 (N_4174,In_658,In_1572);
or U4175 (N_4175,In_1573,In_1571);
nor U4176 (N_4176,In_559,In_2300);
nor U4177 (N_4177,In_1489,In_936);
nor U4178 (N_4178,In_869,In_601);
or U4179 (N_4179,In_1117,In_1781);
nor U4180 (N_4180,In_57,In_1662);
nand U4181 (N_4181,In_469,In_384);
or U4182 (N_4182,In_1279,In_1445);
nor U4183 (N_4183,In_3,In_2236);
xnor U4184 (N_4184,In_2026,In_2074);
nor U4185 (N_4185,In_484,In_476);
or U4186 (N_4186,In_1218,In_895);
nand U4187 (N_4187,In_54,In_1597);
nor U4188 (N_4188,In_1851,In_1279);
and U4189 (N_4189,In_390,In_344);
or U4190 (N_4190,In_1604,In_1817);
and U4191 (N_4191,In_1171,In_1946);
nor U4192 (N_4192,In_2361,In_508);
nand U4193 (N_4193,In_1083,In_818);
or U4194 (N_4194,In_2332,In_498);
nand U4195 (N_4195,In_1405,In_1640);
and U4196 (N_4196,In_1954,In_645);
and U4197 (N_4197,In_1938,In_2371);
nor U4198 (N_4198,In_2293,In_1911);
nor U4199 (N_4199,In_492,In_664);
xor U4200 (N_4200,In_82,In_2170);
or U4201 (N_4201,In_2425,In_628);
nor U4202 (N_4202,In_856,In_669);
nor U4203 (N_4203,In_1865,In_479);
xor U4204 (N_4204,In_214,In_142);
nand U4205 (N_4205,In_1667,In_1225);
nor U4206 (N_4206,In_1584,In_267);
and U4207 (N_4207,In_991,In_658);
and U4208 (N_4208,In_1675,In_738);
nand U4209 (N_4209,In_1084,In_628);
nor U4210 (N_4210,In_1753,In_2342);
and U4211 (N_4211,In_26,In_684);
nor U4212 (N_4212,In_1345,In_1750);
or U4213 (N_4213,In_1422,In_1998);
and U4214 (N_4214,In_1877,In_381);
nand U4215 (N_4215,In_961,In_829);
and U4216 (N_4216,In_2095,In_889);
xnor U4217 (N_4217,In_1096,In_2216);
and U4218 (N_4218,In_1680,In_1444);
and U4219 (N_4219,In_1147,In_361);
and U4220 (N_4220,In_102,In_1967);
nand U4221 (N_4221,In_755,In_1781);
nor U4222 (N_4222,In_1012,In_1337);
nor U4223 (N_4223,In_1474,In_518);
nor U4224 (N_4224,In_1207,In_2491);
xnor U4225 (N_4225,In_705,In_2213);
nor U4226 (N_4226,In_1863,In_1403);
or U4227 (N_4227,In_2388,In_2172);
nand U4228 (N_4228,In_1414,In_679);
and U4229 (N_4229,In_1804,In_1445);
nor U4230 (N_4230,In_1609,In_1243);
nor U4231 (N_4231,In_607,In_1206);
or U4232 (N_4232,In_2404,In_1671);
nand U4233 (N_4233,In_689,In_581);
nand U4234 (N_4234,In_1343,In_1607);
nand U4235 (N_4235,In_1191,In_1435);
nand U4236 (N_4236,In_226,In_984);
and U4237 (N_4237,In_1816,In_1944);
or U4238 (N_4238,In_194,In_988);
and U4239 (N_4239,In_822,In_2363);
nor U4240 (N_4240,In_1519,In_786);
nor U4241 (N_4241,In_1569,In_493);
or U4242 (N_4242,In_2413,In_1686);
nand U4243 (N_4243,In_497,In_1628);
and U4244 (N_4244,In_1660,In_155);
and U4245 (N_4245,In_1805,In_1976);
nor U4246 (N_4246,In_1451,In_377);
nor U4247 (N_4247,In_1371,In_979);
nand U4248 (N_4248,In_2484,In_408);
or U4249 (N_4249,In_802,In_496);
nor U4250 (N_4250,In_1377,In_1445);
nand U4251 (N_4251,In_646,In_2013);
or U4252 (N_4252,In_131,In_702);
or U4253 (N_4253,In_1520,In_389);
xnor U4254 (N_4254,In_2278,In_1937);
and U4255 (N_4255,In_445,In_2472);
and U4256 (N_4256,In_680,In_2425);
and U4257 (N_4257,In_517,In_419);
and U4258 (N_4258,In_751,In_936);
and U4259 (N_4259,In_1176,In_673);
nand U4260 (N_4260,In_484,In_2285);
nor U4261 (N_4261,In_1890,In_1894);
or U4262 (N_4262,In_2477,In_29);
and U4263 (N_4263,In_245,In_1089);
or U4264 (N_4264,In_241,In_1194);
nand U4265 (N_4265,In_2230,In_907);
nor U4266 (N_4266,In_312,In_551);
nand U4267 (N_4267,In_2279,In_2210);
nand U4268 (N_4268,In_2339,In_1434);
nand U4269 (N_4269,In_391,In_1357);
and U4270 (N_4270,In_1997,In_279);
nor U4271 (N_4271,In_1406,In_1743);
and U4272 (N_4272,In_1676,In_623);
and U4273 (N_4273,In_660,In_774);
nor U4274 (N_4274,In_2254,In_896);
nor U4275 (N_4275,In_1742,In_93);
and U4276 (N_4276,In_2334,In_2075);
or U4277 (N_4277,In_930,In_453);
nor U4278 (N_4278,In_453,In_1390);
or U4279 (N_4279,In_1225,In_2319);
xnor U4280 (N_4280,In_2231,In_1310);
nand U4281 (N_4281,In_1631,In_1434);
nor U4282 (N_4282,In_672,In_209);
and U4283 (N_4283,In_2333,In_1593);
or U4284 (N_4284,In_1481,In_416);
nand U4285 (N_4285,In_719,In_2206);
xor U4286 (N_4286,In_1026,In_733);
or U4287 (N_4287,In_883,In_223);
nor U4288 (N_4288,In_260,In_2254);
xnor U4289 (N_4289,In_1448,In_1377);
and U4290 (N_4290,In_2122,In_649);
or U4291 (N_4291,In_2216,In_1311);
nor U4292 (N_4292,In_2037,In_1814);
xor U4293 (N_4293,In_2375,In_457);
or U4294 (N_4294,In_1228,In_1004);
nor U4295 (N_4295,In_1678,In_2459);
or U4296 (N_4296,In_2398,In_2270);
nor U4297 (N_4297,In_1383,In_706);
or U4298 (N_4298,In_1316,In_1932);
nand U4299 (N_4299,In_2111,In_671);
nor U4300 (N_4300,In_2013,In_91);
nor U4301 (N_4301,In_2178,In_194);
or U4302 (N_4302,In_2237,In_1343);
nand U4303 (N_4303,In_2257,In_100);
and U4304 (N_4304,In_2264,In_425);
and U4305 (N_4305,In_1558,In_1891);
xnor U4306 (N_4306,In_2468,In_926);
and U4307 (N_4307,In_815,In_2136);
or U4308 (N_4308,In_2449,In_802);
nand U4309 (N_4309,In_387,In_1062);
xor U4310 (N_4310,In_120,In_1561);
or U4311 (N_4311,In_2121,In_1787);
and U4312 (N_4312,In_437,In_647);
nand U4313 (N_4313,In_1497,In_558);
nor U4314 (N_4314,In_1234,In_2222);
or U4315 (N_4315,In_647,In_1769);
nor U4316 (N_4316,In_1768,In_2224);
nor U4317 (N_4317,In_1928,In_2079);
or U4318 (N_4318,In_623,In_314);
nor U4319 (N_4319,In_475,In_1648);
nor U4320 (N_4320,In_29,In_830);
nor U4321 (N_4321,In_1370,In_746);
xnor U4322 (N_4322,In_580,In_1928);
nand U4323 (N_4323,In_1046,In_110);
xor U4324 (N_4324,In_743,In_1719);
nand U4325 (N_4325,In_1682,In_2300);
nor U4326 (N_4326,In_2352,In_455);
or U4327 (N_4327,In_494,In_1662);
and U4328 (N_4328,In_241,In_1637);
or U4329 (N_4329,In_981,In_2234);
or U4330 (N_4330,In_198,In_1943);
or U4331 (N_4331,In_897,In_575);
nor U4332 (N_4332,In_66,In_1912);
xor U4333 (N_4333,In_409,In_557);
and U4334 (N_4334,In_537,In_1670);
nor U4335 (N_4335,In_2269,In_2074);
and U4336 (N_4336,In_1361,In_1705);
and U4337 (N_4337,In_2122,In_10);
nand U4338 (N_4338,In_594,In_613);
xnor U4339 (N_4339,In_1692,In_433);
and U4340 (N_4340,In_992,In_1699);
nand U4341 (N_4341,In_1729,In_2107);
nand U4342 (N_4342,In_1224,In_2018);
or U4343 (N_4343,In_1992,In_2331);
xor U4344 (N_4344,In_238,In_1054);
nand U4345 (N_4345,In_467,In_303);
nand U4346 (N_4346,In_762,In_2072);
or U4347 (N_4347,In_2478,In_2166);
nand U4348 (N_4348,In_2472,In_1108);
and U4349 (N_4349,In_1412,In_2299);
or U4350 (N_4350,In_1897,In_1933);
or U4351 (N_4351,In_2301,In_1552);
nor U4352 (N_4352,In_2108,In_2274);
nor U4353 (N_4353,In_118,In_2112);
and U4354 (N_4354,In_2160,In_1613);
and U4355 (N_4355,In_2341,In_382);
nor U4356 (N_4356,In_1886,In_1138);
or U4357 (N_4357,In_1689,In_971);
and U4358 (N_4358,In_2397,In_1382);
nand U4359 (N_4359,In_710,In_1290);
nor U4360 (N_4360,In_577,In_1726);
or U4361 (N_4361,In_1688,In_68);
or U4362 (N_4362,In_1231,In_794);
or U4363 (N_4363,In_327,In_1566);
xnor U4364 (N_4364,In_424,In_2168);
xor U4365 (N_4365,In_959,In_1873);
nand U4366 (N_4366,In_134,In_823);
nand U4367 (N_4367,In_369,In_983);
nand U4368 (N_4368,In_848,In_73);
nand U4369 (N_4369,In_318,In_1564);
or U4370 (N_4370,In_1960,In_1871);
xnor U4371 (N_4371,In_2245,In_1446);
xnor U4372 (N_4372,In_2339,In_1690);
nand U4373 (N_4373,In_2437,In_1287);
or U4374 (N_4374,In_1003,In_441);
xor U4375 (N_4375,In_391,In_813);
and U4376 (N_4376,In_887,In_2418);
or U4377 (N_4377,In_274,In_697);
nor U4378 (N_4378,In_2142,In_1899);
nor U4379 (N_4379,In_2338,In_2473);
xnor U4380 (N_4380,In_2075,In_623);
and U4381 (N_4381,In_2000,In_965);
or U4382 (N_4382,In_266,In_647);
nand U4383 (N_4383,In_882,In_1785);
nor U4384 (N_4384,In_1544,In_787);
or U4385 (N_4385,In_2077,In_1965);
nand U4386 (N_4386,In_715,In_2447);
nor U4387 (N_4387,In_415,In_1108);
nand U4388 (N_4388,In_1709,In_1814);
and U4389 (N_4389,In_77,In_2203);
nor U4390 (N_4390,In_1183,In_1479);
and U4391 (N_4391,In_1304,In_2039);
nand U4392 (N_4392,In_1188,In_2249);
and U4393 (N_4393,In_43,In_2021);
nand U4394 (N_4394,In_2456,In_2110);
nor U4395 (N_4395,In_2116,In_1781);
and U4396 (N_4396,In_682,In_1030);
or U4397 (N_4397,In_1408,In_973);
nand U4398 (N_4398,In_1631,In_583);
nand U4399 (N_4399,In_1761,In_1665);
and U4400 (N_4400,In_2346,In_33);
or U4401 (N_4401,In_1071,In_654);
nor U4402 (N_4402,In_2249,In_2321);
or U4403 (N_4403,In_771,In_2322);
and U4404 (N_4404,In_916,In_2371);
nor U4405 (N_4405,In_627,In_1734);
and U4406 (N_4406,In_1032,In_352);
nor U4407 (N_4407,In_1880,In_1251);
nor U4408 (N_4408,In_1540,In_161);
or U4409 (N_4409,In_1472,In_1020);
nand U4410 (N_4410,In_1741,In_1825);
xnor U4411 (N_4411,In_60,In_97);
and U4412 (N_4412,In_1280,In_2028);
or U4413 (N_4413,In_1614,In_2349);
nor U4414 (N_4414,In_1891,In_2342);
nand U4415 (N_4415,In_98,In_670);
xnor U4416 (N_4416,In_626,In_1406);
or U4417 (N_4417,In_1121,In_79);
or U4418 (N_4418,In_1576,In_886);
and U4419 (N_4419,In_817,In_1543);
nand U4420 (N_4420,In_2105,In_1647);
and U4421 (N_4421,In_1473,In_2343);
or U4422 (N_4422,In_1053,In_2291);
and U4423 (N_4423,In_1365,In_1315);
nor U4424 (N_4424,In_139,In_1726);
and U4425 (N_4425,In_378,In_981);
xnor U4426 (N_4426,In_2111,In_1824);
and U4427 (N_4427,In_2402,In_91);
or U4428 (N_4428,In_1075,In_1429);
nor U4429 (N_4429,In_1788,In_1425);
nand U4430 (N_4430,In_1641,In_860);
and U4431 (N_4431,In_880,In_1347);
and U4432 (N_4432,In_1073,In_30);
or U4433 (N_4433,In_790,In_1335);
and U4434 (N_4434,In_1017,In_1983);
and U4435 (N_4435,In_2169,In_1822);
or U4436 (N_4436,In_1307,In_220);
and U4437 (N_4437,In_786,In_477);
nand U4438 (N_4438,In_1397,In_2191);
nand U4439 (N_4439,In_1099,In_1812);
nor U4440 (N_4440,In_2187,In_1422);
nor U4441 (N_4441,In_1614,In_1900);
or U4442 (N_4442,In_127,In_2324);
and U4443 (N_4443,In_963,In_746);
and U4444 (N_4444,In_1881,In_1329);
nand U4445 (N_4445,In_683,In_830);
and U4446 (N_4446,In_141,In_2004);
and U4447 (N_4447,In_505,In_106);
nor U4448 (N_4448,In_1095,In_2251);
and U4449 (N_4449,In_1721,In_2478);
or U4450 (N_4450,In_976,In_1026);
and U4451 (N_4451,In_2311,In_752);
and U4452 (N_4452,In_180,In_697);
nor U4453 (N_4453,In_1936,In_1615);
nand U4454 (N_4454,In_666,In_1001);
and U4455 (N_4455,In_2416,In_1997);
and U4456 (N_4456,In_247,In_1947);
or U4457 (N_4457,In_2427,In_1711);
or U4458 (N_4458,In_2417,In_128);
or U4459 (N_4459,In_2153,In_1023);
and U4460 (N_4460,In_737,In_1986);
or U4461 (N_4461,In_187,In_482);
and U4462 (N_4462,In_1460,In_207);
nor U4463 (N_4463,In_1435,In_913);
xor U4464 (N_4464,In_1256,In_1803);
nor U4465 (N_4465,In_437,In_840);
nor U4466 (N_4466,In_468,In_582);
nand U4467 (N_4467,In_3,In_1446);
nand U4468 (N_4468,In_1057,In_2186);
or U4469 (N_4469,In_2109,In_2225);
or U4470 (N_4470,In_650,In_555);
xnor U4471 (N_4471,In_1554,In_1251);
nand U4472 (N_4472,In_1280,In_1178);
nor U4473 (N_4473,In_1748,In_2057);
and U4474 (N_4474,In_2072,In_2474);
xor U4475 (N_4475,In_929,In_2461);
or U4476 (N_4476,In_969,In_1373);
and U4477 (N_4477,In_225,In_765);
and U4478 (N_4478,In_420,In_1766);
and U4479 (N_4479,In_67,In_1193);
nand U4480 (N_4480,In_1847,In_702);
and U4481 (N_4481,In_2249,In_85);
and U4482 (N_4482,In_2229,In_870);
nand U4483 (N_4483,In_2039,In_1890);
and U4484 (N_4484,In_1036,In_271);
nand U4485 (N_4485,In_1769,In_1017);
xor U4486 (N_4486,In_1676,In_989);
nor U4487 (N_4487,In_282,In_809);
and U4488 (N_4488,In_1896,In_709);
or U4489 (N_4489,In_656,In_1530);
nor U4490 (N_4490,In_2378,In_756);
nand U4491 (N_4491,In_914,In_1680);
nand U4492 (N_4492,In_1215,In_594);
xor U4493 (N_4493,In_528,In_939);
and U4494 (N_4494,In_1422,In_273);
and U4495 (N_4495,In_1251,In_216);
xor U4496 (N_4496,In_1777,In_0);
nand U4497 (N_4497,In_1806,In_1793);
xor U4498 (N_4498,In_1986,In_1209);
and U4499 (N_4499,In_1624,In_1314);
nor U4500 (N_4500,In_201,In_1082);
xor U4501 (N_4501,In_1782,In_2159);
and U4502 (N_4502,In_1911,In_1113);
xnor U4503 (N_4503,In_1290,In_705);
xor U4504 (N_4504,In_2429,In_1996);
nor U4505 (N_4505,In_422,In_1103);
and U4506 (N_4506,In_2318,In_381);
nor U4507 (N_4507,In_307,In_862);
and U4508 (N_4508,In_134,In_153);
nor U4509 (N_4509,In_1964,In_974);
or U4510 (N_4510,In_768,In_1875);
nand U4511 (N_4511,In_905,In_1649);
nor U4512 (N_4512,In_2031,In_517);
nand U4513 (N_4513,In_1031,In_985);
nor U4514 (N_4514,In_912,In_217);
and U4515 (N_4515,In_766,In_346);
nor U4516 (N_4516,In_1020,In_413);
nor U4517 (N_4517,In_1153,In_751);
xnor U4518 (N_4518,In_2249,In_220);
and U4519 (N_4519,In_79,In_1160);
and U4520 (N_4520,In_2054,In_2430);
or U4521 (N_4521,In_1777,In_289);
nor U4522 (N_4522,In_1434,In_1070);
nor U4523 (N_4523,In_1215,In_1463);
and U4524 (N_4524,In_2374,In_805);
or U4525 (N_4525,In_616,In_490);
or U4526 (N_4526,In_1835,In_2055);
nor U4527 (N_4527,In_1055,In_2061);
or U4528 (N_4528,In_102,In_1995);
nor U4529 (N_4529,In_1819,In_1687);
xor U4530 (N_4530,In_1307,In_1440);
or U4531 (N_4531,In_128,In_1858);
and U4532 (N_4532,In_640,In_2196);
and U4533 (N_4533,In_795,In_780);
nor U4534 (N_4534,In_1621,In_833);
nor U4535 (N_4535,In_400,In_2258);
nor U4536 (N_4536,In_366,In_1233);
or U4537 (N_4537,In_515,In_362);
xnor U4538 (N_4538,In_1294,In_1512);
nor U4539 (N_4539,In_463,In_2069);
and U4540 (N_4540,In_1683,In_1920);
xor U4541 (N_4541,In_1351,In_678);
xnor U4542 (N_4542,In_1257,In_1043);
or U4543 (N_4543,In_1407,In_1546);
or U4544 (N_4544,In_2012,In_77);
nor U4545 (N_4545,In_11,In_1851);
and U4546 (N_4546,In_1162,In_710);
nor U4547 (N_4547,In_2363,In_1593);
or U4548 (N_4548,In_2492,In_810);
or U4549 (N_4549,In_566,In_1375);
nor U4550 (N_4550,In_708,In_668);
nand U4551 (N_4551,In_226,In_1211);
nand U4552 (N_4552,In_1870,In_706);
nor U4553 (N_4553,In_1200,In_816);
nand U4554 (N_4554,In_2097,In_678);
and U4555 (N_4555,In_2098,In_2000);
nand U4556 (N_4556,In_1786,In_1616);
nor U4557 (N_4557,In_1019,In_2488);
nor U4558 (N_4558,In_1206,In_1759);
nor U4559 (N_4559,In_956,In_2093);
or U4560 (N_4560,In_841,In_2372);
nand U4561 (N_4561,In_2203,In_2255);
nor U4562 (N_4562,In_136,In_988);
nand U4563 (N_4563,In_2418,In_2494);
nand U4564 (N_4564,In_152,In_1817);
and U4565 (N_4565,In_1960,In_2431);
nand U4566 (N_4566,In_1535,In_1590);
nor U4567 (N_4567,In_886,In_2123);
nand U4568 (N_4568,In_2098,In_1442);
nor U4569 (N_4569,In_431,In_608);
nor U4570 (N_4570,In_1811,In_413);
or U4571 (N_4571,In_402,In_355);
nor U4572 (N_4572,In_481,In_2227);
and U4573 (N_4573,In_1039,In_755);
nand U4574 (N_4574,In_216,In_2271);
nand U4575 (N_4575,In_2444,In_1490);
and U4576 (N_4576,In_1137,In_1552);
nor U4577 (N_4577,In_986,In_588);
nor U4578 (N_4578,In_2441,In_417);
nor U4579 (N_4579,In_1220,In_630);
nand U4580 (N_4580,In_186,In_2043);
nor U4581 (N_4581,In_1449,In_1640);
xnor U4582 (N_4582,In_380,In_879);
nor U4583 (N_4583,In_1652,In_1822);
or U4584 (N_4584,In_1163,In_1860);
nor U4585 (N_4585,In_338,In_500);
nand U4586 (N_4586,In_1479,In_2277);
or U4587 (N_4587,In_2425,In_992);
nor U4588 (N_4588,In_1515,In_1108);
or U4589 (N_4589,In_699,In_2217);
or U4590 (N_4590,In_1344,In_2173);
and U4591 (N_4591,In_1371,In_742);
or U4592 (N_4592,In_2196,In_83);
xnor U4593 (N_4593,In_2032,In_1768);
nor U4594 (N_4594,In_1673,In_707);
and U4595 (N_4595,In_200,In_859);
nor U4596 (N_4596,In_629,In_1266);
nand U4597 (N_4597,In_1361,In_805);
or U4598 (N_4598,In_1468,In_1828);
xnor U4599 (N_4599,In_861,In_1508);
or U4600 (N_4600,In_1365,In_598);
nor U4601 (N_4601,In_1402,In_1085);
or U4602 (N_4602,In_1493,In_919);
or U4603 (N_4603,In_12,In_1062);
nor U4604 (N_4604,In_664,In_1031);
nor U4605 (N_4605,In_2322,In_1562);
nand U4606 (N_4606,In_2368,In_531);
and U4607 (N_4607,In_1405,In_2201);
nor U4608 (N_4608,In_1905,In_1762);
nand U4609 (N_4609,In_347,In_2329);
nand U4610 (N_4610,In_1632,In_2210);
xor U4611 (N_4611,In_1835,In_90);
or U4612 (N_4612,In_156,In_306);
or U4613 (N_4613,In_969,In_2238);
and U4614 (N_4614,In_816,In_1737);
nand U4615 (N_4615,In_289,In_1060);
xnor U4616 (N_4616,In_356,In_1196);
nand U4617 (N_4617,In_2093,In_1672);
or U4618 (N_4618,In_136,In_1153);
nor U4619 (N_4619,In_1846,In_1148);
or U4620 (N_4620,In_2068,In_594);
nor U4621 (N_4621,In_2377,In_278);
xor U4622 (N_4622,In_2451,In_1778);
and U4623 (N_4623,In_380,In_523);
nand U4624 (N_4624,In_2107,In_1989);
nor U4625 (N_4625,In_2005,In_1699);
and U4626 (N_4626,In_595,In_2061);
nor U4627 (N_4627,In_1677,In_287);
nand U4628 (N_4628,In_2102,In_2422);
and U4629 (N_4629,In_2091,In_1019);
nand U4630 (N_4630,In_933,In_1200);
and U4631 (N_4631,In_1931,In_691);
or U4632 (N_4632,In_1239,In_1987);
nand U4633 (N_4633,In_1495,In_38);
or U4634 (N_4634,In_1802,In_81);
xor U4635 (N_4635,In_58,In_1769);
xnor U4636 (N_4636,In_949,In_1967);
and U4637 (N_4637,In_2231,In_1726);
or U4638 (N_4638,In_1162,In_1748);
or U4639 (N_4639,In_2388,In_1886);
nor U4640 (N_4640,In_50,In_14);
nor U4641 (N_4641,In_212,In_2117);
nand U4642 (N_4642,In_180,In_453);
nand U4643 (N_4643,In_1180,In_137);
or U4644 (N_4644,In_1831,In_1684);
xnor U4645 (N_4645,In_1315,In_1689);
or U4646 (N_4646,In_478,In_2399);
nor U4647 (N_4647,In_2485,In_113);
nor U4648 (N_4648,In_1909,In_1885);
and U4649 (N_4649,In_237,In_160);
and U4650 (N_4650,In_509,In_1414);
or U4651 (N_4651,In_2452,In_1169);
and U4652 (N_4652,In_1069,In_821);
or U4653 (N_4653,In_508,In_1563);
nand U4654 (N_4654,In_2374,In_884);
nor U4655 (N_4655,In_1858,In_1458);
or U4656 (N_4656,In_2252,In_2123);
nand U4657 (N_4657,In_707,In_230);
nand U4658 (N_4658,In_874,In_1052);
nand U4659 (N_4659,In_2039,In_992);
nor U4660 (N_4660,In_1494,In_1171);
nand U4661 (N_4661,In_439,In_1192);
nand U4662 (N_4662,In_451,In_449);
nand U4663 (N_4663,In_856,In_17);
and U4664 (N_4664,In_2312,In_1014);
or U4665 (N_4665,In_1651,In_176);
nand U4666 (N_4666,In_1616,In_1460);
and U4667 (N_4667,In_2136,In_2066);
xnor U4668 (N_4668,In_917,In_1411);
and U4669 (N_4669,In_877,In_1050);
and U4670 (N_4670,In_630,In_611);
nor U4671 (N_4671,In_870,In_356);
nand U4672 (N_4672,In_182,In_1485);
nor U4673 (N_4673,In_1141,In_2265);
nor U4674 (N_4674,In_1794,In_2229);
nand U4675 (N_4675,In_1313,In_912);
nand U4676 (N_4676,In_204,In_1117);
nor U4677 (N_4677,In_1833,In_712);
xnor U4678 (N_4678,In_164,In_2480);
nor U4679 (N_4679,In_61,In_831);
or U4680 (N_4680,In_1916,In_1658);
and U4681 (N_4681,In_2210,In_1959);
or U4682 (N_4682,In_290,In_1017);
and U4683 (N_4683,In_2102,In_601);
nand U4684 (N_4684,In_1275,In_1867);
nor U4685 (N_4685,In_528,In_1254);
nor U4686 (N_4686,In_764,In_201);
nand U4687 (N_4687,In_1211,In_1821);
nand U4688 (N_4688,In_1421,In_1887);
nor U4689 (N_4689,In_1274,In_1729);
and U4690 (N_4690,In_2111,In_2176);
nor U4691 (N_4691,In_1071,In_1856);
xnor U4692 (N_4692,In_237,In_715);
nor U4693 (N_4693,In_1569,In_1972);
nor U4694 (N_4694,In_343,In_2339);
or U4695 (N_4695,In_2216,In_1919);
xor U4696 (N_4696,In_1064,In_1034);
and U4697 (N_4697,In_1418,In_1589);
or U4698 (N_4698,In_433,In_2470);
nand U4699 (N_4699,In_694,In_1073);
nor U4700 (N_4700,In_973,In_1239);
and U4701 (N_4701,In_2101,In_2461);
nand U4702 (N_4702,In_949,In_541);
nand U4703 (N_4703,In_240,In_312);
and U4704 (N_4704,In_1081,In_209);
nand U4705 (N_4705,In_2026,In_728);
and U4706 (N_4706,In_741,In_114);
or U4707 (N_4707,In_2370,In_1207);
or U4708 (N_4708,In_20,In_2169);
or U4709 (N_4709,In_2215,In_2012);
or U4710 (N_4710,In_2085,In_405);
nand U4711 (N_4711,In_1284,In_1598);
and U4712 (N_4712,In_671,In_2022);
or U4713 (N_4713,In_14,In_1274);
or U4714 (N_4714,In_1724,In_1642);
or U4715 (N_4715,In_938,In_2238);
and U4716 (N_4716,In_2455,In_2039);
nor U4717 (N_4717,In_52,In_1100);
nand U4718 (N_4718,In_1307,In_1223);
nor U4719 (N_4719,In_878,In_1545);
and U4720 (N_4720,In_695,In_2495);
or U4721 (N_4721,In_623,In_223);
or U4722 (N_4722,In_1451,In_1390);
or U4723 (N_4723,In_1685,In_2008);
nor U4724 (N_4724,In_1534,In_1928);
or U4725 (N_4725,In_864,In_199);
or U4726 (N_4726,In_1803,In_470);
or U4727 (N_4727,In_489,In_160);
or U4728 (N_4728,In_1082,In_336);
nor U4729 (N_4729,In_1538,In_2451);
xnor U4730 (N_4730,In_319,In_2220);
or U4731 (N_4731,In_1031,In_2332);
nand U4732 (N_4732,In_496,In_1332);
nand U4733 (N_4733,In_943,In_1255);
and U4734 (N_4734,In_2417,In_191);
xnor U4735 (N_4735,In_1617,In_186);
or U4736 (N_4736,In_38,In_1064);
nand U4737 (N_4737,In_285,In_154);
nand U4738 (N_4738,In_574,In_1496);
nor U4739 (N_4739,In_528,In_517);
or U4740 (N_4740,In_482,In_1989);
or U4741 (N_4741,In_288,In_1002);
nand U4742 (N_4742,In_1517,In_2373);
and U4743 (N_4743,In_443,In_1096);
and U4744 (N_4744,In_2225,In_336);
nor U4745 (N_4745,In_1030,In_1519);
nand U4746 (N_4746,In_1434,In_1982);
nor U4747 (N_4747,In_374,In_127);
nand U4748 (N_4748,In_1903,In_226);
nor U4749 (N_4749,In_2148,In_144);
and U4750 (N_4750,In_445,In_1513);
or U4751 (N_4751,In_752,In_1924);
nand U4752 (N_4752,In_751,In_914);
or U4753 (N_4753,In_779,In_503);
nand U4754 (N_4754,In_125,In_2062);
or U4755 (N_4755,In_1511,In_791);
nand U4756 (N_4756,In_2135,In_1326);
or U4757 (N_4757,In_48,In_744);
nand U4758 (N_4758,In_382,In_138);
nor U4759 (N_4759,In_1652,In_579);
or U4760 (N_4760,In_998,In_1332);
or U4761 (N_4761,In_2217,In_1933);
nor U4762 (N_4762,In_2110,In_829);
or U4763 (N_4763,In_966,In_54);
nor U4764 (N_4764,In_849,In_2144);
nor U4765 (N_4765,In_109,In_2330);
and U4766 (N_4766,In_1183,In_2024);
and U4767 (N_4767,In_595,In_419);
nor U4768 (N_4768,In_2096,In_1998);
or U4769 (N_4769,In_1022,In_697);
nor U4770 (N_4770,In_1116,In_1756);
xor U4771 (N_4771,In_1437,In_209);
nand U4772 (N_4772,In_513,In_475);
or U4773 (N_4773,In_686,In_1314);
nor U4774 (N_4774,In_1665,In_1141);
or U4775 (N_4775,In_688,In_695);
and U4776 (N_4776,In_1558,In_807);
or U4777 (N_4777,In_1115,In_393);
nor U4778 (N_4778,In_730,In_218);
or U4779 (N_4779,In_1795,In_479);
and U4780 (N_4780,In_2328,In_485);
nand U4781 (N_4781,In_1323,In_2302);
nor U4782 (N_4782,In_1019,In_872);
xor U4783 (N_4783,In_645,In_107);
and U4784 (N_4784,In_673,In_2498);
nand U4785 (N_4785,In_795,In_1455);
or U4786 (N_4786,In_1038,In_1821);
or U4787 (N_4787,In_177,In_1428);
or U4788 (N_4788,In_1617,In_1101);
nor U4789 (N_4789,In_2309,In_1260);
nand U4790 (N_4790,In_455,In_1041);
and U4791 (N_4791,In_1900,In_2311);
and U4792 (N_4792,In_682,In_349);
or U4793 (N_4793,In_2212,In_2002);
nand U4794 (N_4794,In_840,In_195);
nor U4795 (N_4795,In_503,In_606);
or U4796 (N_4796,In_253,In_555);
or U4797 (N_4797,In_1701,In_1959);
or U4798 (N_4798,In_1799,In_1198);
or U4799 (N_4799,In_1714,In_2012);
nand U4800 (N_4800,In_39,In_1318);
nor U4801 (N_4801,In_207,In_684);
or U4802 (N_4802,In_1592,In_1112);
nand U4803 (N_4803,In_1608,In_1776);
and U4804 (N_4804,In_1989,In_2293);
nor U4805 (N_4805,In_235,In_1892);
and U4806 (N_4806,In_2415,In_1594);
or U4807 (N_4807,In_1796,In_1648);
nor U4808 (N_4808,In_1021,In_356);
and U4809 (N_4809,In_2044,In_770);
xnor U4810 (N_4810,In_1156,In_1618);
nand U4811 (N_4811,In_1447,In_692);
nand U4812 (N_4812,In_770,In_1531);
and U4813 (N_4813,In_1522,In_1487);
or U4814 (N_4814,In_131,In_1942);
and U4815 (N_4815,In_1803,In_790);
nor U4816 (N_4816,In_168,In_2134);
and U4817 (N_4817,In_2283,In_1532);
nand U4818 (N_4818,In_670,In_2307);
nor U4819 (N_4819,In_412,In_1072);
or U4820 (N_4820,In_1771,In_2411);
and U4821 (N_4821,In_682,In_1080);
nor U4822 (N_4822,In_2312,In_858);
xor U4823 (N_4823,In_1860,In_845);
nor U4824 (N_4824,In_1125,In_1355);
and U4825 (N_4825,In_679,In_215);
nand U4826 (N_4826,In_2028,In_735);
xor U4827 (N_4827,In_1544,In_1357);
nor U4828 (N_4828,In_2403,In_247);
nor U4829 (N_4829,In_2474,In_1928);
nor U4830 (N_4830,In_804,In_1902);
xnor U4831 (N_4831,In_2305,In_1102);
xnor U4832 (N_4832,In_188,In_182);
nand U4833 (N_4833,In_1512,In_1713);
xor U4834 (N_4834,In_2081,In_232);
or U4835 (N_4835,In_867,In_1936);
nand U4836 (N_4836,In_1641,In_975);
nand U4837 (N_4837,In_51,In_1492);
xor U4838 (N_4838,In_1964,In_2406);
nor U4839 (N_4839,In_1426,In_2038);
and U4840 (N_4840,In_2349,In_141);
nand U4841 (N_4841,In_2336,In_404);
nor U4842 (N_4842,In_646,In_1817);
xnor U4843 (N_4843,In_921,In_476);
and U4844 (N_4844,In_761,In_683);
and U4845 (N_4845,In_2473,In_1435);
nor U4846 (N_4846,In_1944,In_1365);
or U4847 (N_4847,In_998,In_2012);
nand U4848 (N_4848,In_595,In_2347);
xor U4849 (N_4849,In_2377,In_2434);
or U4850 (N_4850,In_1189,In_2484);
or U4851 (N_4851,In_120,In_53);
or U4852 (N_4852,In_2010,In_744);
nor U4853 (N_4853,In_1838,In_1576);
and U4854 (N_4854,In_1920,In_591);
and U4855 (N_4855,In_1732,In_1698);
xnor U4856 (N_4856,In_739,In_534);
nand U4857 (N_4857,In_1836,In_545);
or U4858 (N_4858,In_1056,In_190);
or U4859 (N_4859,In_2100,In_1579);
nand U4860 (N_4860,In_2200,In_855);
or U4861 (N_4861,In_2001,In_1717);
nor U4862 (N_4862,In_61,In_1026);
or U4863 (N_4863,In_2431,In_176);
or U4864 (N_4864,In_2270,In_1040);
and U4865 (N_4865,In_650,In_126);
nand U4866 (N_4866,In_1545,In_2103);
nor U4867 (N_4867,In_128,In_825);
nor U4868 (N_4868,In_1531,In_1968);
and U4869 (N_4869,In_1124,In_2329);
nand U4870 (N_4870,In_2460,In_1794);
nand U4871 (N_4871,In_1287,In_267);
and U4872 (N_4872,In_766,In_849);
nor U4873 (N_4873,In_1815,In_326);
and U4874 (N_4874,In_2272,In_892);
nor U4875 (N_4875,In_733,In_1150);
and U4876 (N_4876,In_1998,In_865);
nand U4877 (N_4877,In_1733,In_2401);
xor U4878 (N_4878,In_874,In_2007);
and U4879 (N_4879,In_2267,In_642);
or U4880 (N_4880,In_969,In_2333);
or U4881 (N_4881,In_1043,In_2498);
xnor U4882 (N_4882,In_2467,In_1749);
and U4883 (N_4883,In_224,In_147);
or U4884 (N_4884,In_2204,In_1848);
xnor U4885 (N_4885,In_2257,In_1904);
and U4886 (N_4886,In_2188,In_74);
nand U4887 (N_4887,In_330,In_1996);
and U4888 (N_4888,In_1723,In_138);
nand U4889 (N_4889,In_214,In_1402);
or U4890 (N_4890,In_1734,In_219);
nand U4891 (N_4891,In_388,In_492);
nand U4892 (N_4892,In_993,In_998);
or U4893 (N_4893,In_832,In_1614);
nand U4894 (N_4894,In_670,In_1338);
or U4895 (N_4895,In_217,In_192);
xnor U4896 (N_4896,In_1203,In_936);
and U4897 (N_4897,In_2102,In_787);
nand U4898 (N_4898,In_675,In_1043);
nand U4899 (N_4899,In_1181,In_804);
or U4900 (N_4900,In_1208,In_1231);
nor U4901 (N_4901,In_100,In_2002);
and U4902 (N_4902,In_2382,In_1308);
or U4903 (N_4903,In_599,In_1680);
or U4904 (N_4904,In_1584,In_1508);
nor U4905 (N_4905,In_1998,In_550);
nand U4906 (N_4906,In_2282,In_691);
nor U4907 (N_4907,In_1718,In_559);
nand U4908 (N_4908,In_224,In_2202);
and U4909 (N_4909,In_1140,In_1760);
or U4910 (N_4910,In_801,In_51);
nor U4911 (N_4911,In_1498,In_1196);
or U4912 (N_4912,In_2346,In_1177);
or U4913 (N_4913,In_663,In_1107);
nand U4914 (N_4914,In_2312,In_449);
nand U4915 (N_4915,In_1744,In_2475);
nor U4916 (N_4916,In_1128,In_211);
and U4917 (N_4917,In_661,In_1734);
nand U4918 (N_4918,In_1773,In_19);
nor U4919 (N_4919,In_1260,In_1852);
or U4920 (N_4920,In_2291,In_580);
and U4921 (N_4921,In_608,In_1190);
nor U4922 (N_4922,In_1275,In_991);
nor U4923 (N_4923,In_643,In_2135);
xnor U4924 (N_4924,In_1990,In_2476);
nor U4925 (N_4925,In_117,In_2221);
or U4926 (N_4926,In_1749,In_1312);
nor U4927 (N_4927,In_896,In_1069);
nor U4928 (N_4928,In_910,In_1015);
xnor U4929 (N_4929,In_317,In_529);
or U4930 (N_4930,In_820,In_839);
xor U4931 (N_4931,In_1033,In_1681);
or U4932 (N_4932,In_308,In_1453);
nor U4933 (N_4933,In_1639,In_2269);
nand U4934 (N_4934,In_1277,In_627);
or U4935 (N_4935,In_1452,In_357);
nor U4936 (N_4936,In_753,In_2149);
nor U4937 (N_4937,In_988,In_110);
or U4938 (N_4938,In_573,In_1314);
nand U4939 (N_4939,In_1736,In_1336);
nor U4940 (N_4940,In_1599,In_2256);
nand U4941 (N_4941,In_767,In_10);
xnor U4942 (N_4942,In_1298,In_2395);
nor U4943 (N_4943,In_1341,In_563);
nand U4944 (N_4944,In_1948,In_372);
or U4945 (N_4945,In_1939,In_2046);
nor U4946 (N_4946,In_1614,In_2025);
nand U4947 (N_4947,In_16,In_502);
nand U4948 (N_4948,In_2388,In_315);
and U4949 (N_4949,In_1761,In_1222);
nand U4950 (N_4950,In_1089,In_2289);
nand U4951 (N_4951,In_769,In_988);
nand U4952 (N_4952,In_681,In_1972);
nor U4953 (N_4953,In_1556,In_807);
nor U4954 (N_4954,In_1259,In_1871);
and U4955 (N_4955,In_1093,In_1329);
xor U4956 (N_4956,In_1971,In_1813);
nand U4957 (N_4957,In_2233,In_394);
nand U4958 (N_4958,In_1716,In_1565);
or U4959 (N_4959,In_1959,In_1286);
and U4960 (N_4960,In_2467,In_557);
xor U4961 (N_4961,In_141,In_2392);
nand U4962 (N_4962,In_2137,In_1583);
xnor U4963 (N_4963,In_2344,In_1822);
or U4964 (N_4964,In_1778,In_670);
or U4965 (N_4965,In_2339,In_249);
and U4966 (N_4966,In_345,In_2065);
or U4967 (N_4967,In_1087,In_1283);
and U4968 (N_4968,In_1196,In_820);
nor U4969 (N_4969,In_647,In_1266);
or U4970 (N_4970,In_328,In_537);
or U4971 (N_4971,In_1859,In_2408);
nand U4972 (N_4972,In_1121,In_1158);
and U4973 (N_4973,In_2175,In_348);
nor U4974 (N_4974,In_2389,In_2023);
nor U4975 (N_4975,In_244,In_2395);
nand U4976 (N_4976,In_1225,In_1562);
and U4977 (N_4977,In_10,In_2333);
and U4978 (N_4978,In_950,In_541);
nor U4979 (N_4979,In_887,In_1493);
nand U4980 (N_4980,In_522,In_444);
nor U4981 (N_4981,In_1584,In_2018);
xor U4982 (N_4982,In_2072,In_1317);
nand U4983 (N_4983,In_851,In_1211);
nand U4984 (N_4984,In_1307,In_653);
nor U4985 (N_4985,In_503,In_2310);
xnor U4986 (N_4986,In_2234,In_105);
xor U4987 (N_4987,In_2397,In_704);
and U4988 (N_4988,In_2138,In_826);
nand U4989 (N_4989,In_1852,In_269);
and U4990 (N_4990,In_97,In_382);
xnor U4991 (N_4991,In_928,In_2370);
nand U4992 (N_4992,In_2062,In_731);
nor U4993 (N_4993,In_1731,In_994);
nand U4994 (N_4994,In_2197,In_2215);
or U4995 (N_4995,In_373,In_252);
xnor U4996 (N_4996,In_1987,In_1594);
nor U4997 (N_4997,In_50,In_724);
nor U4998 (N_4998,In_413,In_1342);
or U4999 (N_4999,In_1921,In_238);
nand U5000 (N_5000,In_131,In_1592);
and U5001 (N_5001,In_1989,In_2213);
nor U5002 (N_5002,In_993,In_2086);
nor U5003 (N_5003,In_1668,In_342);
nand U5004 (N_5004,In_1187,In_1756);
and U5005 (N_5005,In_2330,In_406);
nand U5006 (N_5006,In_1370,In_2205);
or U5007 (N_5007,In_1697,In_113);
nand U5008 (N_5008,In_1201,In_680);
nor U5009 (N_5009,In_2093,In_1424);
or U5010 (N_5010,In_583,In_2282);
or U5011 (N_5011,In_1225,In_1362);
or U5012 (N_5012,In_1580,In_727);
nor U5013 (N_5013,In_564,In_470);
or U5014 (N_5014,In_1667,In_2239);
or U5015 (N_5015,In_251,In_2460);
nor U5016 (N_5016,In_38,In_2018);
nor U5017 (N_5017,In_2405,In_274);
xnor U5018 (N_5018,In_837,In_815);
and U5019 (N_5019,In_1933,In_1461);
and U5020 (N_5020,In_72,In_1237);
xor U5021 (N_5021,In_196,In_1456);
and U5022 (N_5022,In_2345,In_1737);
nand U5023 (N_5023,In_19,In_1495);
or U5024 (N_5024,In_2062,In_60);
and U5025 (N_5025,In_879,In_2283);
nor U5026 (N_5026,In_492,In_2176);
nor U5027 (N_5027,In_117,In_1718);
nor U5028 (N_5028,In_784,In_1312);
or U5029 (N_5029,In_267,In_1500);
nor U5030 (N_5030,In_1935,In_2116);
and U5031 (N_5031,In_1268,In_264);
or U5032 (N_5032,In_744,In_1749);
and U5033 (N_5033,In_108,In_1303);
and U5034 (N_5034,In_947,In_429);
or U5035 (N_5035,In_247,In_380);
xor U5036 (N_5036,In_2102,In_401);
and U5037 (N_5037,In_634,In_51);
or U5038 (N_5038,In_1095,In_1398);
nand U5039 (N_5039,In_1585,In_388);
or U5040 (N_5040,In_388,In_1002);
nor U5041 (N_5041,In_305,In_1937);
nor U5042 (N_5042,In_2488,In_55);
and U5043 (N_5043,In_181,In_1950);
xor U5044 (N_5044,In_2212,In_450);
or U5045 (N_5045,In_2177,In_44);
nor U5046 (N_5046,In_1508,In_1123);
nand U5047 (N_5047,In_1567,In_2332);
nand U5048 (N_5048,In_1475,In_646);
nand U5049 (N_5049,In_1082,In_1548);
xnor U5050 (N_5050,In_2483,In_873);
nor U5051 (N_5051,In_2159,In_129);
and U5052 (N_5052,In_403,In_453);
nor U5053 (N_5053,In_1783,In_2135);
nand U5054 (N_5054,In_2359,In_627);
nand U5055 (N_5055,In_1067,In_1226);
xnor U5056 (N_5056,In_1137,In_453);
and U5057 (N_5057,In_1806,In_468);
nand U5058 (N_5058,In_671,In_227);
nor U5059 (N_5059,In_1371,In_1787);
nor U5060 (N_5060,In_308,In_1286);
nor U5061 (N_5061,In_66,In_1506);
and U5062 (N_5062,In_642,In_2195);
or U5063 (N_5063,In_1365,In_1897);
nor U5064 (N_5064,In_2279,In_1557);
or U5065 (N_5065,In_848,In_679);
nand U5066 (N_5066,In_1914,In_148);
nand U5067 (N_5067,In_1843,In_366);
nand U5068 (N_5068,In_1119,In_2390);
and U5069 (N_5069,In_455,In_1280);
nand U5070 (N_5070,In_1774,In_2126);
nor U5071 (N_5071,In_1407,In_78);
nand U5072 (N_5072,In_1800,In_2215);
or U5073 (N_5073,In_696,In_2453);
or U5074 (N_5074,In_1641,In_2118);
and U5075 (N_5075,In_142,In_38);
or U5076 (N_5076,In_2281,In_1064);
nor U5077 (N_5077,In_1679,In_1920);
and U5078 (N_5078,In_1207,In_373);
xor U5079 (N_5079,In_13,In_1918);
nand U5080 (N_5080,In_2203,In_1300);
nand U5081 (N_5081,In_68,In_676);
and U5082 (N_5082,In_1693,In_173);
or U5083 (N_5083,In_1341,In_1014);
and U5084 (N_5084,In_120,In_127);
and U5085 (N_5085,In_2264,In_1750);
nand U5086 (N_5086,In_1230,In_1570);
or U5087 (N_5087,In_1428,In_1918);
nand U5088 (N_5088,In_1480,In_2420);
or U5089 (N_5089,In_989,In_341);
and U5090 (N_5090,In_2093,In_979);
xnor U5091 (N_5091,In_1535,In_2484);
or U5092 (N_5092,In_155,In_1779);
nor U5093 (N_5093,In_442,In_241);
nor U5094 (N_5094,In_1608,In_1541);
nor U5095 (N_5095,In_2147,In_264);
nand U5096 (N_5096,In_1578,In_1030);
or U5097 (N_5097,In_2372,In_1022);
or U5098 (N_5098,In_2085,In_10);
nand U5099 (N_5099,In_1156,In_2039);
xor U5100 (N_5100,In_1163,In_1980);
nor U5101 (N_5101,In_1719,In_191);
nor U5102 (N_5102,In_565,In_1816);
nor U5103 (N_5103,In_1880,In_55);
nand U5104 (N_5104,In_864,In_2271);
nor U5105 (N_5105,In_2175,In_1835);
xor U5106 (N_5106,In_1150,In_1607);
nand U5107 (N_5107,In_191,In_1863);
nand U5108 (N_5108,In_1991,In_1743);
or U5109 (N_5109,In_1098,In_2423);
nand U5110 (N_5110,In_1292,In_1963);
nor U5111 (N_5111,In_1427,In_2101);
and U5112 (N_5112,In_1913,In_746);
nand U5113 (N_5113,In_1612,In_1243);
or U5114 (N_5114,In_1302,In_199);
or U5115 (N_5115,In_483,In_566);
or U5116 (N_5116,In_2393,In_1463);
nand U5117 (N_5117,In_2338,In_756);
nor U5118 (N_5118,In_1071,In_953);
nor U5119 (N_5119,In_1798,In_1313);
xnor U5120 (N_5120,In_1720,In_1859);
and U5121 (N_5121,In_1613,In_1602);
nor U5122 (N_5122,In_585,In_1986);
nand U5123 (N_5123,In_1355,In_1411);
nand U5124 (N_5124,In_498,In_194);
nor U5125 (N_5125,In_48,In_1142);
xor U5126 (N_5126,In_416,In_220);
nand U5127 (N_5127,In_206,In_1649);
and U5128 (N_5128,In_1871,In_2406);
nand U5129 (N_5129,In_1791,In_1340);
or U5130 (N_5130,In_1723,In_783);
nor U5131 (N_5131,In_198,In_635);
xnor U5132 (N_5132,In_1091,In_8);
nor U5133 (N_5133,In_1274,In_1089);
nand U5134 (N_5134,In_165,In_2167);
xor U5135 (N_5135,In_1402,In_600);
nand U5136 (N_5136,In_1994,In_1872);
xnor U5137 (N_5137,In_2409,In_849);
nand U5138 (N_5138,In_404,In_2250);
and U5139 (N_5139,In_1212,In_1324);
nor U5140 (N_5140,In_1849,In_200);
and U5141 (N_5141,In_1095,In_1071);
nor U5142 (N_5142,In_1545,In_744);
xor U5143 (N_5143,In_1338,In_1915);
and U5144 (N_5144,In_1604,In_1056);
xnor U5145 (N_5145,In_1356,In_2222);
nand U5146 (N_5146,In_1353,In_1743);
xnor U5147 (N_5147,In_2428,In_69);
nor U5148 (N_5148,In_1067,In_418);
nand U5149 (N_5149,In_704,In_894);
nor U5150 (N_5150,In_1527,In_535);
nor U5151 (N_5151,In_4,In_1376);
nor U5152 (N_5152,In_1484,In_606);
xnor U5153 (N_5153,In_132,In_498);
xnor U5154 (N_5154,In_160,In_998);
nand U5155 (N_5155,In_2495,In_2178);
nor U5156 (N_5156,In_536,In_1992);
and U5157 (N_5157,In_763,In_2373);
or U5158 (N_5158,In_1665,In_1790);
nand U5159 (N_5159,In_958,In_1209);
or U5160 (N_5160,In_882,In_303);
or U5161 (N_5161,In_2412,In_1535);
nand U5162 (N_5162,In_1003,In_404);
nor U5163 (N_5163,In_2445,In_1166);
and U5164 (N_5164,In_403,In_1862);
nor U5165 (N_5165,In_1768,In_1121);
or U5166 (N_5166,In_195,In_2027);
nand U5167 (N_5167,In_468,In_1657);
nand U5168 (N_5168,In_2360,In_1465);
or U5169 (N_5169,In_719,In_1357);
nand U5170 (N_5170,In_746,In_1156);
nor U5171 (N_5171,In_950,In_30);
or U5172 (N_5172,In_2022,In_1051);
nor U5173 (N_5173,In_167,In_171);
nand U5174 (N_5174,In_1639,In_206);
xor U5175 (N_5175,In_1471,In_1728);
nor U5176 (N_5176,In_283,In_2176);
nand U5177 (N_5177,In_713,In_1723);
nand U5178 (N_5178,In_2072,In_2382);
and U5179 (N_5179,In_326,In_473);
nand U5180 (N_5180,In_2446,In_1104);
nor U5181 (N_5181,In_527,In_1523);
and U5182 (N_5182,In_1780,In_2078);
or U5183 (N_5183,In_497,In_1904);
or U5184 (N_5184,In_989,In_666);
nor U5185 (N_5185,In_403,In_96);
nand U5186 (N_5186,In_1830,In_1178);
and U5187 (N_5187,In_575,In_604);
nand U5188 (N_5188,In_2229,In_1307);
xor U5189 (N_5189,In_1171,In_63);
nand U5190 (N_5190,In_1513,In_1204);
and U5191 (N_5191,In_2016,In_902);
nand U5192 (N_5192,In_117,In_29);
nor U5193 (N_5193,In_425,In_113);
nand U5194 (N_5194,In_644,In_729);
nand U5195 (N_5195,In_681,In_1445);
and U5196 (N_5196,In_224,In_1575);
nor U5197 (N_5197,In_1496,In_1101);
nor U5198 (N_5198,In_1532,In_283);
and U5199 (N_5199,In_1324,In_905);
nor U5200 (N_5200,In_732,In_1199);
nand U5201 (N_5201,In_215,In_1786);
nor U5202 (N_5202,In_807,In_763);
and U5203 (N_5203,In_1724,In_2404);
nand U5204 (N_5204,In_898,In_1454);
and U5205 (N_5205,In_2345,In_1623);
nand U5206 (N_5206,In_2167,In_889);
nor U5207 (N_5207,In_916,In_2016);
and U5208 (N_5208,In_967,In_91);
nand U5209 (N_5209,In_499,In_2209);
and U5210 (N_5210,In_1697,In_114);
and U5211 (N_5211,In_312,In_2064);
nor U5212 (N_5212,In_2452,In_87);
nor U5213 (N_5213,In_339,In_1970);
or U5214 (N_5214,In_1413,In_1765);
xor U5215 (N_5215,In_1322,In_2003);
nor U5216 (N_5216,In_1224,In_471);
and U5217 (N_5217,In_1224,In_98);
and U5218 (N_5218,In_1235,In_2144);
nor U5219 (N_5219,In_2481,In_30);
nand U5220 (N_5220,In_1773,In_1598);
or U5221 (N_5221,In_1402,In_623);
or U5222 (N_5222,In_839,In_2008);
nand U5223 (N_5223,In_2236,In_504);
or U5224 (N_5224,In_922,In_2049);
nand U5225 (N_5225,In_1587,In_894);
nor U5226 (N_5226,In_578,In_958);
and U5227 (N_5227,In_1286,In_1672);
xor U5228 (N_5228,In_406,In_943);
and U5229 (N_5229,In_743,In_1635);
nor U5230 (N_5230,In_1824,In_1233);
and U5231 (N_5231,In_122,In_1792);
nor U5232 (N_5232,In_981,In_2160);
xnor U5233 (N_5233,In_829,In_1156);
xor U5234 (N_5234,In_501,In_2016);
or U5235 (N_5235,In_819,In_984);
nand U5236 (N_5236,In_167,In_1954);
and U5237 (N_5237,In_1822,In_213);
nand U5238 (N_5238,In_2343,In_956);
nor U5239 (N_5239,In_1906,In_1827);
nor U5240 (N_5240,In_1998,In_710);
nand U5241 (N_5241,In_339,In_1947);
and U5242 (N_5242,In_1684,In_706);
or U5243 (N_5243,In_1064,In_1212);
and U5244 (N_5244,In_107,In_572);
nor U5245 (N_5245,In_1325,In_1247);
nor U5246 (N_5246,In_1346,In_1104);
nor U5247 (N_5247,In_582,In_1057);
nor U5248 (N_5248,In_1569,In_2371);
and U5249 (N_5249,In_389,In_2463);
or U5250 (N_5250,In_2472,In_2141);
or U5251 (N_5251,In_2041,In_207);
or U5252 (N_5252,In_2034,In_2132);
nand U5253 (N_5253,In_742,In_56);
or U5254 (N_5254,In_325,In_1490);
nand U5255 (N_5255,In_204,In_1930);
and U5256 (N_5256,In_188,In_618);
nand U5257 (N_5257,In_1860,In_740);
nand U5258 (N_5258,In_1717,In_108);
or U5259 (N_5259,In_1807,In_1633);
nand U5260 (N_5260,In_1830,In_1821);
nand U5261 (N_5261,In_1502,In_410);
nor U5262 (N_5262,In_2367,In_1612);
xnor U5263 (N_5263,In_1311,In_767);
or U5264 (N_5264,In_2006,In_29);
xor U5265 (N_5265,In_1575,In_2250);
or U5266 (N_5266,In_2491,In_2323);
nand U5267 (N_5267,In_590,In_774);
xnor U5268 (N_5268,In_657,In_434);
nor U5269 (N_5269,In_86,In_366);
xnor U5270 (N_5270,In_1275,In_922);
nand U5271 (N_5271,In_1410,In_2259);
nand U5272 (N_5272,In_1511,In_706);
nand U5273 (N_5273,In_68,In_2289);
or U5274 (N_5274,In_2270,In_190);
nand U5275 (N_5275,In_25,In_1479);
or U5276 (N_5276,In_1587,In_675);
and U5277 (N_5277,In_577,In_1413);
or U5278 (N_5278,In_235,In_2117);
or U5279 (N_5279,In_915,In_2196);
and U5280 (N_5280,In_986,In_47);
nand U5281 (N_5281,In_1394,In_575);
nor U5282 (N_5282,In_918,In_1458);
nand U5283 (N_5283,In_2422,In_352);
and U5284 (N_5284,In_541,In_2137);
nand U5285 (N_5285,In_56,In_165);
xnor U5286 (N_5286,In_1257,In_1859);
nor U5287 (N_5287,In_357,In_1379);
xor U5288 (N_5288,In_907,In_461);
nor U5289 (N_5289,In_409,In_827);
and U5290 (N_5290,In_639,In_1296);
or U5291 (N_5291,In_1213,In_736);
nand U5292 (N_5292,In_1953,In_1888);
and U5293 (N_5293,In_105,In_632);
nor U5294 (N_5294,In_948,In_1078);
or U5295 (N_5295,In_414,In_2411);
nand U5296 (N_5296,In_16,In_1998);
and U5297 (N_5297,In_1151,In_585);
nor U5298 (N_5298,In_682,In_1957);
and U5299 (N_5299,In_52,In_2325);
nor U5300 (N_5300,In_553,In_816);
or U5301 (N_5301,In_50,In_435);
or U5302 (N_5302,In_998,In_2021);
and U5303 (N_5303,In_2255,In_1548);
or U5304 (N_5304,In_419,In_327);
or U5305 (N_5305,In_1347,In_2419);
or U5306 (N_5306,In_395,In_53);
and U5307 (N_5307,In_1462,In_2374);
nand U5308 (N_5308,In_356,In_984);
and U5309 (N_5309,In_1791,In_2034);
nor U5310 (N_5310,In_106,In_637);
nand U5311 (N_5311,In_557,In_1485);
nor U5312 (N_5312,In_338,In_1884);
xor U5313 (N_5313,In_2185,In_2018);
nand U5314 (N_5314,In_402,In_1938);
nand U5315 (N_5315,In_1638,In_2011);
and U5316 (N_5316,In_1773,In_1497);
nand U5317 (N_5317,In_1872,In_597);
or U5318 (N_5318,In_1632,In_700);
nor U5319 (N_5319,In_114,In_2339);
or U5320 (N_5320,In_991,In_338);
or U5321 (N_5321,In_801,In_2323);
and U5322 (N_5322,In_2039,In_1495);
nor U5323 (N_5323,In_543,In_312);
nand U5324 (N_5324,In_2232,In_1910);
or U5325 (N_5325,In_1306,In_1441);
and U5326 (N_5326,In_952,In_2222);
xor U5327 (N_5327,In_1109,In_443);
nand U5328 (N_5328,In_2311,In_2118);
or U5329 (N_5329,In_1140,In_103);
xor U5330 (N_5330,In_2051,In_1335);
nand U5331 (N_5331,In_462,In_890);
nor U5332 (N_5332,In_1680,In_1301);
or U5333 (N_5333,In_1280,In_2269);
nor U5334 (N_5334,In_265,In_2425);
nand U5335 (N_5335,In_897,In_2281);
nand U5336 (N_5336,In_195,In_1987);
nor U5337 (N_5337,In_1153,In_256);
or U5338 (N_5338,In_124,In_1917);
nand U5339 (N_5339,In_1480,In_485);
or U5340 (N_5340,In_1635,In_1843);
and U5341 (N_5341,In_2016,In_300);
or U5342 (N_5342,In_230,In_115);
and U5343 (N_5343,In_23,In_1831);
nor U5344 (N_5344,In_736,In_2491);
and U5345 (N_5345,In_1131,In_39);
xor U5346 (N_5346,In_21,In_1257);
nor U5347 (N_5347,In_1785,In_263);
nand U5348 (N_5348,In_508,In_1094);
xnor U5349 (N_5349,In_1529,In_734);
and U5350 (N_5350,In_1727,In_1082);
or U5351 (N_5351,In_662,In_1021);
or U5352 (N_5352,In_2340,In_456);
and U5353 (N_5353,In_1661,In_89);
and U5354 (N_5354,In_372,In_2332);
or U5355 (N_5355,In_2408,In_774);
xnor U5356 (N_5356,In_1282,In_1911);
or U5357 (N_5357,In_1154,In_460);
nor U5358 (N_5358,In_2032,In_1296);
or U5359 (N_5359,In_2297,In_2413);
nand U5360 (N_5360,In_1144,In_922);
xor U5361 (N_5361,In_1545,In_1007);
nand U5362 (N_5362,In_1515,In_625);
and U5363 (N_5363,In_2036,In_1200);
nand U5364 (N_5364,In_868,In_217);
and U5365 (N_5365,In_1897,In_205);
nor U5366 (N_5366,In_210,In_1313);
nand U5367 (N_5367,In_151,In_1193);
nor U5368 (N_5368,In_952,In_1166);
xnor U5369 (N_5369,In_2385,In_1253);
or U5370 (N_5370,In_1724,In_228);
nor U5371 (N_5371,In_1539,In_1427);
or U5372 (N_5372,In_760,In_383);
and U5373 (N_5373,In_1026,In_18);
nand U5374 (N_5374,In_1999,In_1950);
or U5375 (N_5375,In_2363,In_1156);
and U5376 (N_5376,In_2260,In_2251);
or U5377 (N_5377,In_2338,In_853);
nand U5378 (N_5378,In_2218,In_1125);
nor U5379 (N_5379,In_1364,In_1083);
and U5380 (N_5380,In_884,In_2180);
nor U5381 (N_5381,In_1627,In_29);
nand U5382 (N_5382,In_2243,In_1803);
and U5383 (N_5383,In_1339,In_1385);
nand U5384 (N_5384,In_2376,In_2295);
nand U5385 (N_5385,In_897,In_989);
or U5386 (N_5386,In_735,In_1346);
or U5387 (N_5387,In_2463,In_2395);
nor U5388 (N_5388,In_1926,In_1850);
or U5389 (N_5389,In_205,In_1366);
xor U5390 (N_5390,In_782,In_1810);
and U5391 (N_5391,In_2194,In_669);
nand U5392 (N_5392,In_24,In_410);
or U5393 (N_5393,In_282,In_867);
nand U5394 (N_5394,In_456,In_1191);
and U5395 (N_5395,In_1479,In_2297);
or U5396 (N_5396,In_2228,In_812);
nand U5397 (N_5397,In_850,In_2361);
or U5398 (N_5398,In_545,In_209);
nor U5399 (N_5399,In_1023,In_1889);
or U5400 (N_5400,In_1420,In_1945);
and U5401 (N_5401,In_860,In_722);
or U5402 (N_5402,In_101,In_1677);
or U5403 (N_5403,In_41,In_2440);
nor U5404 (N_5404,In_1632,In_1808);
xor U5405 (N_5405,In_539,In_1965);
nor U5406 (N_5406,In_2194,In_3);
and U5407 (N_5407,In_1017,In_621);
or U5408 (N_5408,In_919,In_99);
or U5409 (N_5409,In_769,In_1303);
nor U5410 (N_5410,In_296,In_94);
and U5411 (N_5411,In_557,In_2264);
or U5412 (N_5412,In_1178,In_768);
or U5413 (N_5413,In_2359,In_1397);
xnor U5414 (N_5414,In_837,In_1734);
nor U5415 (N_5415,In_1265,In_1673);
nand U5416 (N_5416,In_851,In_1695);
nor U5417 (N_5417,In_1068,In_2053);
nand U5418 (N_5418,In_1742,In_1514);
xor U5419 (N_5419,In_1472,In_379);
nor U5420 (N_5420,In_2074,In_2219);
and U5421 (N_5421,In_1776,In_199);
nand U5422 (N_5422,In_2030,In_1296);
nor U5423 (N_5423,In_2028,In_1023);
nor U5424 (N_5424,In_2284,In_995);
or U5425 (N_5425,In_529,In_834);
or U5426 (N_5426,In_1728,In_2400);
nand U5427 (N_5427,In_1161,In_2416);
nor U5428 (N_5428,In_2123,In_1315);
nor U5429 (N_5429,In_1989,In_2065);
nand U5430 (N_5430,In_2392,In_2305);
or U5431 (N_5431,In_2439,In_92);
and U5432 (N_5432,In_1051,In_1056);
nand U5433 (N_5433,In_277,In_2370);
xor U5434 (N_5434,In_1412,In_831);
nand U5435 (N_5435,In_16,In_400);
and U5436 (N_5436,In_964,In_68);
nand U5437 (N_5437,In_1889,In_1814);
or U5438 (N_5438,In_753,In_996);
nor U5439 (N_5439,In_1539,In_1883);
xnor U5440 (N_5440,In_1019,In_106);
nor U5441 (N_5441,In_526,In_1732);
or U5442 (N_5442,In_2464,In_798);
nand U5443 (N_5443,In_459,In_1824);
and U5444 (N_5444,In_602,In_1047);
or U5445 (N_5445,In_543,In_1338);
nand U5446 (N_5446,In_269,In_731);
and U5447 (N_5447,In_1433,In_126);
and U5448 (N_5448,In_1573,In_186);
and U5449 (N_5449,In_1192,In_253);
and U5450 (N_5450,In_2130,In_1020);
nand U5451 (N_5451,In_65,In_883);
nand U5452 (N_5452,In_2287,In_1856);
or U5453 (N_5453,In_249,In_1645);
nand U5454 (N_5454,In_1383,In_1277);
and U5455 (N_5455,In_703,In_876);
nand U5456 (N_5456,In_690,In_2364);
and U5457 (N_5457,In_1622,In_1308);
or U5458 (N_5458,In_1920,In_847);
nor U5459 (N_5459,In_243,In_822);
and U5460 (N_5460,In_1503,In_2268);
and U5461 (N_5461,In_414,In_264);
xnor U5462 (N_5462,In_1743,In_273);
or U5463 (N_5463,In_1132,In_1388);
nand U5464 (N_5464,In_1273,In_1652);
and U5465 (N_5465,In_1235,In_997);
nor U5466 (N_5466,In_2156,In_1352);
or U5467 (N_5467,In_1649,In_2076);
nor U5468 (N_5468,In_680,In_1963);
and U5469 (N_5469,In_908,In_919);
nor U5470 (N_5470,In_1223,In_1333);
nor U5471 (N_5471,In_2230,In_918);
or U5472 (N_5472,In_48,In_334);
and U5473 (N_5473,In_808,In_2469);
nor U5474 (N_5474,In_310,In_120);
nor U5475 (N_5475,In_432,In_857);
nand U5476 (N_5476,In_457,In_1455);
and U5477 (N_5477,In_833,In_2364);
and U5478 (N_5478,In_2142,In_673);
and U5479 (N_5479,In_1172,In_474);
and U5480 (N_5480,In_1479,In_2415);
or U5481 (N_5481,In_980,In_765);
xor U5482 (N_5482,In_166,In_1547);
nand U5483 (N_5483,In_1248,In_2363);
nor U5484 (N_5484,In_483,In_1888);
nor U5485 (N_5485,In_521,In_1263);
and U5486 (N_5486,In_790,In_2286);
nand U5487 (N_5487,In_1876,In_1965);
xnor U5488 (N_5488,In_289,In_2075);
nor U5489 (N_5489,In_2229,In_1073);
or U5490 (N_5490,In_916,In_1085);
nor U5491 (N_5491,In_1682,In_78);
and U5492 (N_5492,In_182,In_1915);
nand U5493 (N_5493,In_1145,In_107);
xor U5494 (N_5494,In_1358,In_1977);
xnor U5495 (N_5495,In_2426,In_1578);
nor U5496 (N_5496,In_1533,In_362);
xor U5497 (N_5497,In_1603,In_803);
xor U5498 (N_5498,In_1534,In_544);
nand U5499 (N_5499,In_1871,In_1885);
and U5500 (N_5500,In_1982,In_674);
nor U5501 (N_5501,In_2072,In_110);
xor U5502 (N_5502,In_425,In_1761);
nor U5503 (N_5503,In_2386,In_1759);
nor U5504 (N_5504,In_1740,In_1212);
or U5505 (N_5505,In_1245,In_1116);
xnor U5506 (N_5506,In_1556,In_579);
nand U5507 (N_5507,In_511,In_484);
xnor U5508 (N_5508,In_1339,In_868);
or U5509 (N_5509,In_1035,In_205);
and U5510 (N_5510,In_1400,In_615);
nand U5511 (N_5511,In_780,In_484);
or U5512 (N_5512,In_650,In_757);
and U5513 (N_5513,In_1029,In_1952);
nand U5514 (N_5514,In_967,In_894);
nor U5515 (N_5515,In_1683,In_1349);
or U5516 (N_5516,In_1282,In_1511);
or U5517 (N_5517,In_1421,In_2408);
or U5518 (N_5518,In_348,In_50);
nand U5519 (N_5519,In_2211,In_2424);
and U5520 (N_5520,In_615,In_1110);
or U5521 (N_5521,In_673,In_216);
or U5522 (N_5522,In_2295,In_442);
nor U5523 (N_5523,In_1658,In_419);
and U5524 (N_5524,In_1857,In_2026);
or U5525 (N_5525,In_558,In_1690);
nor U5526 (N_5526,In_1522,In_570);
nor U5527 (N_5527,In_600,In_291);
nor U5528 (N_5528,In_1863,In_2431);
nor U5529 (N_5529,In_1450,In_2401);
nor U5530 (N_5530,In_11,In_1256);
xnor U5531 (N_5531,In_82,In_267);
nor U5532 (N_5532,In_793,In_1063);
nor U5533 (N_5533,In_1417,In_1847);
and U5534 (N_5534,In_853,In_1281);
and U5535 (N_5535,In_1069,In_1430);
nor U5536 (N_5536,In_2149,In_405);
nor U5537 (N_5537,In_899,In_508);
and U5538 (N_5538,In_1860,In_2180);
and U5539 (N_5539,In_2243,In_1359);
nand U5540 (N_5540,In_2397,In_1937);
nand U5541 (N_5541,In_331,In_976);
or U5542 (N_5542,In_702,In_1833);
nor U5543 (N_5543,In_1595,In_2342);
nor U5544 (N_5544,In_2215,In_1597);
xnor U5545 (N_5545,In_2197,In_195);
or U5546 (N_5546,In_328,In_739);
or U5547 (N_5547,In_1736,In_1337);
or U5548 (N_5548,In_2448,In_1115);
nand U5549 (N_5549,In_1865,In_550);
nor U5550 (N_5550,In_2409,In_751);
or U5551 (N_5551,In_124,In_1749);
or U5552 (N_5552,In_890,In_668);
or U5553 (N_5553,In_972,In_2018);
or U5554 (N_5554,In_905,In_1506);
nand U5555 (N_5555,In_1880,In_764);
xor U5556 (N_5556,In_448,In_293);
nand U5557 (N_5557,In_2094,In_2235);
nand U5558 (N_5558,In_1014,In_1358);
or U5559 (N_5559,In_1212,In_1930);
nor U5560 (N_5560,In_123,In_1431);
nand U5561 (N_5561,In_2158,In_1881);
and U5562 (N_5562,In_33,In_2192);
or U5563 (N_5563,In_1691,In_2194);
or U5564 (N_5564,In_581,In_628);
or U5565 (N_5565,In_1171,In_1210);
or U5566 (N_5566,In_904,In_1125);
and U5567 (N_5567,In_39,In_2416);
nor U5568 (N_5568,In_15,In_1553);
and U5569 (N_5569,In_382,In_708);
and U5570 (N_5570,In_1214,In_535);
or U5571 (N_5571,In_1095,In_2324);
nor U5572 (N_5572,In_1509,In_1666);
nand U5573 (N_5573,In_437,In_742);
and U5574 (N_5574,In_2230,In_65);
xnor U5575 (N_5575,In_805,In_1940);
or U5576 (N_5576,In_1023,In_2208);
and U5577 (N_5577,In_1230,In_2386);
and U5578 (N_5578,In_1694,In_1168);
and U5579 (N_5579,In_1661,In_126);
nor U5580 (N_5580,In_1563,In_1973);
and U5581 (N_5581,In_1218,In_1983);
and U5582 (N_5582,In_1065,In_2381);
or U5583 (N_5583,In_1826,In_2050);
nor U5584 (N_5584,In_1802,In_2251);
nand U5585 (N_5585,In_2326,In_1483);
xnor U5586 (N_5586,In_2455,In_2487);
and U5587 (N_5587,In_2075,In_1831);
nand U5588 (N_5588,In_1858,In_2365);
nor U5589 (N_5589,In_1076,In_2292);
nand U5590 (N_5590,In_1481,In_2035);
and U5591 (N_5591,In_1585,In_2173);
and U5592 (N_5592,In_1561,In_840);
nand U5593 (N_5593,In_393,In_2395);
xnor U5594 (N_5594,In_1695,In_915);
xor U5595 (N_5595,In_1047,In_2065);
or U5596 (N_5596,In_1063,In_868);
nand U5597 (N_5597,In_1982,In_1994);
and U5598 (N_5598,In_358,In_2387);
or U5599 (N_5599,In_1993,In_984);
nor U5600 (N_5600,In_2032,In_1346);
nand U5601 (N_5601,In_1449,In_1283);
nor U5602 (N_5602,In_1890,In_28);
nand U5603 (N_5603,In_246,In_2393);
and U5604 (N_5604,In_932,In_2042);
and U5605 (N_5605,In_112,In_1915);
and U5606 (N_5606,In_333,In_2039);
nand U5607 (N_5607,In_692,In_1056);
or U5608 (N_5608,In_611,In_2168);
nor U5609 (N_5609,In_663,In_1460);
or U5610 (N_5610,In_794,In_1992);
and U5611 (N_5611,In_127,In_1091);
and U5612 (N_5612,In_2218,In_2292);
or U5613 (N_5613,In_175,In_1692);
or U5614 (N_5614,In_828,In_1461);
or U5615 (N_5615,In_516,In_1097);
nor U5616 (N_5616,In_406,In_2054);
xor U5617 (N_5617,In_80,In_217);
xor U5618 (N_5618,In_154,In_1815);
or U5619 (N_5619,In_645,In_574);
nand U5620 (N_5620,In_2352,In_637);
xnor U5621 (N_5621,In_2185,In_1240);
and U5622 (N_5622,In_908,In_1875);
xor U5623 (N_5623,In_772,In_1466);
xnor U5624 (N_5624,In_70,In_2043);
and U5625 (N_5625,In_2432,In_644);
xor U5626 (N_5626,In_2369,In_2305);
nor U5627 (N_5627,In_2112,In_1971);
nor U5628 (N_5628,In_213,In_2070);
and U5629 (N_5629,In_1546,In_1688);
or U5630 (N_5630,In_367,In_396);
or U5631 (N_5631,In_1297,In_1882);
nand U5632 (N_5632,In_1861,In_1555);
and U5633 (N_5633,In_342,In_981);
nand U5634 (N_5634,In_1657,In_109);
or U5635 (N_5635,In_1745,In_144);
or U5636 (N_5636,In_1525,In_236);
nand U5637 (N_5637,In_365,In_991);
nor U5638 (N_5638,In_1508,In_656);
nand U5639 (N_5639,In_1026,In_1773);
or U5640 (N_5640,In_1763,In_291);
xor U5641 (N_5641,In_1072,In_1826);
nor U5642 (N_5642,In_1384,In_1926);
nor U5643 (N_5643,In_853,In_2191);
and U5644 (N_5644,In_362,In_2184);
or U5645 (N_5645,In_1926,In_701);
xor U5646 (N_5646,In_857,In_345);
or U5647 (N_5647,In_2236,In_1974);
or U5648 (N_5648,In_897,In_588);
and U5649 (N_5649,In_1315,In_1313);
nor U5650 (N_5650,In_331,In_1435);
or U5651 (N_5651,In_2024,In_638);
or U5652 (N_5652,In_225,In_1513);
nor U5653 (N_5653,In_182,In_1370);
nand U5654 (N_5654,In_874,In_523);
nor U5655 (N_5655,In_300,In_1184);
nor U5656 (N_5656,In_633,In_973);
nor U5657 (N_5657,In_2084,In_1005);
xor U5658 (N_5658,In_409,In_1577);
nand U5659 (N_5659,In_1479,In_1894);
nand U5660 (N_5660,In_481,In_2492);
nand U5661 (N_5661,In_196,In_1145);
or U5662 (N_5662,In_1015,In_1943);
nand U5663 (N_5663,In_209,In_981);
nor U5664 (N_5664,In_1384,In_1976);
nand U5665 (N_5665,In_2170,In_735);
and U5666 (N_5666,In_2311,In_209);
or U5667 (N_5667,In_436,In_764);
nand U5668 (N_5668,In_62,In_1180);
xor U5669 (N_5669,In_1422,In_186);
xnor U5670 (N_5670,In_1096,In_2332);
and U5671 (N_5671,In_1449,In_1124);
or U5672 (N_5672,In_993,In_2147);
or U5673 (N_5673,In_2294,In_553);
and U5674 (N_5674,In_1375,In_1057);
nor U5675 (N_5675,In_350,In_305);
nand U5676 (N_5676,In_1398,In_80);
nor U5677 (N_5677,In_1625,In_637);
nor U5678 (N_5678,In_1067,In_406);
or U5679 (N_5679,In_2098,In_1660);
or U5680 (N_5680,In_699,In_1701);
nor U5681 (N_5681,In_2312,In_116);
nor U5682 (N_5682,In_105,In_1550);
and U5683 (N_5683,In_1043,In_2228);
nor U5684 (N_5684,In_1345,In_814);
xor U5685 (N_5685,In_2169,In_647);
nand U5686 (N_5686,In_1524,In_412);
nand U5687 (N_5687,In_2136,In_580);
and U5688 (N_5688,In_1037,In_982);
and U5689 (N_5689,In_713,In_869);
or U5690 (N_5690,In_1723,In_1405);
or U5691 (N_5691,In_1441,In_1267);
nand U5692 (N_5692,In_1076,In_2146);
nor U5693 (N_5693,In_1977,In_244);
nand U5694 (N_5694,In_715,In_360);
or U5695 (N_5695,In_349,In_1834);
nand U5696 (N_5696,In_699,In_335);
or U5697 (N_5697,In_2048,In_2185);
nor U5698 (N_5698,In_1410,In_792);
and U5699 (N_5699,In_797,In_1759);
and U5700 (N_5700,In_1044,In_2017);
or U5701 (N_5701,In_1307,In_257);
or U5702 (N_5702,In_925,In_1584);
and U5703 (N_5703,In_163,In_83);
nor U5704 (N_5704,In_1770,In_860);
and U5705 (N_5705,In_237,In_1621);
nor U5706 (N_5706,In_229,In_686);
or U5707 (N_5707,In_1069,In_585);
xnor U5708 (N_5708,In_897,In_2166);
nor U5709 (N_5709,In_506,In_1012);
nand U5710 (N_5710,In_421,In_1613);
xnor U5711 (N_5711,In_1047,In_1234);
or U5712 (N_5712,In_2251,In_1226);
and U5713 (N_5713,In_188,In_1381);
nor U5714 (N_5714,In_2035,In_830);
nor U5715 (N_5715,In_1175,In_756);
nand U5716 (N_5716,In_1919,In_2282);
and U5717 (N_5717,In_1134,In_1090);
or U5718 (N_5718,In_1986,In_525);
nor U5719 (N_5719,In_980,In_368);
nand U5720 (N_5720,In_165,In_2375);
nand U5721 (N_5721,In_907,In_1129);
nand U5722 (N_5722,In_1465,In_1458);
or U5723 (N_5723,In_1606,In_2101);
nor U5724 (N_5724,In_1181,In_2262);
nand U5725 (N_5725,In_504,In_2287);
or U5726 (N_5726,In_319,In_114);
and U5727 (N_5727,In_2016,In_1799);
nand U5728 (N_5728,In_634,In_710);
or U5729 (N_5729,In_1681,In_1649);
nor U5730 (N_5730,In_707,In_2025);
nor U5731 (N_5731,In_1202,In_849);
and U5732 (N_5732,In_1342,In_2310);
or U5733 (N_5733,In_2167,In_929);
and U5734 (N_5734,In_481,In_1136);
and U5735 (N_5735,In_296,In_476);
nor U5736 (N_5736,In_2054,In_1103);
and U5737 (N_5737,In_862,In_2383);
nand U5738 (N_5738,In_2210,In_1907);
nand U5739 (N_5739,In_1763,In_1732);
or U5740 (N_5740,In_1842,In_1300);
and U5741 (N_5741,In_732,In_2135);
nand U5742 (N_5742,In_1153,In_1545);
nor U5743 (N_5743,In_1919,In_761);
and U5744 (N_5744,In_2141,In_256);
or U5745 (N_5745,In_1289,In_1589);
and U5746 (N_5746,In_329,In_1495);
xnor U5747 (N_5747,In_1177,In_2041);
nor U5748 (N_5748,In_2247,In_1616);
and U5749 (N_5749,In_52,In_460);
and U5750 (N_5750,In_1961,In_1813);
nor U5751 (N_5751,In_94,In_1506);
xor U5752 (N_5752,In_2184,In_1779);
nand U5753 (N_5753,In_1987,In_249);
and U5754 (N_5754,In_1871,In_1644);
or U5755 (N_5755,In_238,In_1425);
and U5756 (N_5756,In_1185,In_1590);
nor U5757 (N_5757,In_36,In_2245);
nor U5758 (N_5758,In_317,In_2147);
nand U5759 (N_5759,In_1085,In_510);
or U5760 (N_5760,In_2296,In_2064);
or U5761 (N_5761,In_209,In_1112);
nand U5762 (N_5762,In_1373,In_1598);
nor U5763 (N_5763,In_2420,In_2431);
or U5764 (N_5764,In_252,In_269);
nand U5765 (N_5765,In_192,In_713);
or U5766 (N_5766,In_1034,In_1272);
or U5767 (N_5767,In_2470,In_985);
nand U5768 (N_5768,In_1806,In_1227);
or U5769 (N_5769,In_2321,In_325);
nand U5770 (N_5770,In_1871,In_1442);
and U5771 (N_5771,In_632,In_1330);
nor U5772 (N_5772,In_2362,In_875);
and U5773 (N_5773,In_1329,In_1040);
and U5774 (N_5774,In_2368,In_1322);
and U5775 (N_5775,In_1412,In_1306);
or U5776 (N_5776,In_301,In_2184);
xor U5777 (N_5777,In_1038,In_638);
nor U5778 (N_5778,In_1138,In_1384);
or U5779 (N_5779,In_909,In_1785);
nor U5780 (N_5780,In_998,In_806);
nor U5781 (N_5781,In_2117,In_1812);
nand U5782 (N_5782,In_2112,In_128);
xor U5783 (N_5783,In_162,In_598);
and U5784 (N_5784,In_315,In_1619);
nand U5785 (N_5785,In_835,In_992);
xnor U5786 (N_5786,In_1106,In_1743);
nor U5787 (N_5787,In_2429,In_880);
nand U5788 (N_5788,In_449,In_1218);
or U5789 (N_5789,In_1177,In_2111);
and U5790 (N_5790,In_1798,In_1278);
and U5791 (N_5791,In_1255,In_881);
nand U5792 (N_5792,In_437,In_878);
or U5793 (N_5793,In_827,In_1237);
nor U5794 (N_5794,In_962,In_1911);
or U5795 (N_5795,In_395,In_1147);
or U5796 (N_5796,In_780,In_2144);
and U5797 (N_5797,In_450,In_1101);
and U5798 (N_5798,In_2063,In_2354);
and U5799 (N_5799,In_1084,In_32);
or U5800 (N_5800,In_2000,In_749);
xnor U5801 (N_5801,In_966,In_727);
or U5802 (N_5802,In_964,In_92);
xnor U5803 (N_5803,In_1422,In_960);
xnor U5804 (N_5804,In_2376,In_903);
or U5805 (N_5805,In_992,In_1534);
xor U5806 (N_5806,In_254,In_558);
and U5807 (N_5807,In_652,In_1622);
nand U5808 (N_5808,In_1475,In_1151);
and U5809 (N_5809,In_574,In_1669);
or U5810 (N_5810,In_1389,In_2216);
and U5811 (N_5811,In_467,In_1756);
nand U5812 (N_5812,In_1308,In_2128);
and U5813 (N_5813,In_2113,In_2428);
nand U5814 (N_5814,In_2109,In_1747);
nor U5815 (N_5815,In_761,In_923);
nand U5816 (N_5816,In_1205,In_1170);
nor U5817 (N_5817,In_544,In_1725);
nor U5818 (N_5818,In_862,In_1120);
and U5819 (N_5819,In_2395,In_173);
nand U5820 (N_5820,In_2482,In_460);
or U5821 (N_5821,In_893,In_1829);
nand U5822 (N_5822,In_2146,In_1517);
nand U5823 (N_5823,In_396,In_1128);
nand U5824 (N_5824,In_1382,In_308);
nand U5825 (N_5825,In_1858,In_157);
nand U5826 (N_5826,In_1313,In_2407);
or U5827 (N_5827,In_2155,In_2393);
or U5828 (N_5828,In_605,In_471);
nand U5829 (N_5829,In_1332,In_2011);
nor U5830 (N_5830,In_2027,In_825);
and U5831 (N_5831,In_1585,In_2028);
and U5832 (N_5832,In_949,In_527);
nor U5833 (N_5833,In_1554,In_947);
or U5834 (N_5834,In_527,In_1638);
and U5835 (N_5835,In_1489,In_722);
xor U5836 (N_5836,In_2412,In_2201);
and U5837 (N_5837,In_49,In_1489);
nor U5838 (N_5838,In_1473,In_2443);
nor U5839 (N_5839,In_551,In_2150);
nor U5840 (N_5840,In_2209,In_917);
xor U5841 (N_5841,In_754,In_1758);
nor U5842 (N_5842,In_1346,In_1351);
nand U5843 (N_5843,In_1842,In_1376);
xnor U5844 (N_5844,In_22,In_1940);
nor U5845 (N_5845,In_1097,In_2252);
or U5846 (N_5846,In_751,In_1373);
nor U5847 (N_5847,In_2091,In_777);
nor U5848 (N_5848,In_682,In_2032);
nand U5849 (N_5849,In_826,In_728);
nand U5850 (N_5850,In_494,In_2292);
nand U5851 (N_5851,In_1742,In_1044);
nand U5852 (N_5852,In_830,In_1256);
or U5853 (N_5853,In_947,In_400);
nor U5854 (N_5854,In_771,In_733);
or U5855 (N_5855,In_1326,In_2065);
nand U5856 (N_5856,In_4,In_1477);
or U5857 (N_5857,In_432,In_1761);
xnor U5858 (N_5858,In_834,In_311);
nor U5859 (N_5859,In_766,In_63);
nor U5860 (N_5860,In_884,In_1847);
nor U5861 (N_5861,In_331,In_228);
nor U5862 (N_5862,In_1224,In_567);
and U5863 (N_5863,In_916,In_1807);
nand U5864 (N_5864,In_1459,In_2232);
nor U5865 (N_5865,In_2287,In_2494);
nor U5866 (N_5866,In_823,In_1477);
or U5867 (N_5867,In_1543,In_540);
and U5868 (N_5868,In_1908,In_2217);
xor U5869 (N_5869,In_243,In_2309);
nor U5870 (N_5870,In_2484,In_304);
and U5871 (N_5871,In_1575,In_2341);
nor U5872 (N_5872,In_1896,In_124);
nor U5873 (N_5873,In_410,In_76);
and U5874 (N_5874,In_656,In_394);
and U5875 (N_5875,In_2169,In_279);
or U5876 (N_5876,In_1790,In_1332);
or U5877 (N_5877,In_1651,In_198);
and U5878 (N_5878,In_1547,In_368);
and U5879 (N_5879,In_2386,In_772);
nor U5880 (N_5880,In_1055,In_107);
and U5881 (N_5881,In_427,In_111);
nor U5882 (N_5882,In_886,In_1448);
nor U5883 (N_5883,In_973,In_2306);
xor U5884 (N_5884,In_961,In_1009);
or U5885 (N_5885,In_1053,In_2024);
or U5886 (N_5886,In_1045,In_317);
or U5887 (N_5887,In_211,In_2067);
and U5888 (N_5888,In_1373,In_2257);
nand U5889 (N_5889,In_656,In_74);
or U5890 (N_5890,In_1884,In_810);
xor U5891 (N_5891,In_2079,In_1803);
and U5892 (N_5892,In_2269,In_538);
and U5893 (N_5893,In_1979,In_1196);
nand U5894 (N_5894,In_631,In_2124);
or U5895 (N_5895,In_1778,In_957);
and U5896 (N_5896,In_1162,In_825);
nand U5897 (N_5897,In_2334,In_1907);
or U5898 (N_5898,In_2421,In_1858);
nor U5899 (N_5899,In_360,In_684);
or U5900 (N_5900,In_2069,In_956);
nand U5901 (N_5901,In_1926,In_1330);
xnor U5902 (N_5902,In_1625,In_1570);
or U5903 (N_5903,In_1672,In_120);
nor U5904 (N_5904,In_1505,In_2305);
and U5905 (N_5905,In_906,In_470);
and U5906 (N_5906,In_1794,In_2245);
and U5907 (N_5907,In_1879,In_1560);
nand U5908 (N_5908,In_1987,In_1536);
nand U5909 (N_5909,In_1959,In_1424);
nand U5910 (N_5910,In_686,In_2);
nor U5911 (N_5911,In_1250,In_1659);
or U5912 (N_5912,In_2209,In_923);
or U5913 (N_5913,In_252,In_1791);
or U5914 (N_5914,In_2470,In_1176);
nor U5915 (N_5915,In_884,In_469);
xor U5916 (N_5916,In_1963,In_1135);
and U5917 (N_5917,In_433,In_2169);
nor U5918 (N_5918,In_1587,In_2125);
nor U5919 (N_5919,In_746,In_179);
nor U5920 (N_5920,In_1013,In_1267);
nor U5921 (N_5921,In_609,In_1024);
nand U5922 (N_5922,In_1808,In_117);
nor U5923 (N_5923,In_156,In_25);
and U5924 (N_5924,In_1176,In_1500);
nor U5925 (N_5925,In_39,In_1226);
nand U5926 (N_5926,In_1787,In_1215);
or U5927 (N_5927,In_1248,In_268);
nand U5928 (N_5928,In_1167,In_878);
or U5929 (N_5929,In_1275,In_753);
and U5930 (N_5930,In_2335,In_936);
and U5931 (N_5931,In_179,In_86);
nor U5932 (N_5932,In_4,In_1968);
nor U5933 (N_5933,In_458,In_2094);
xnor U5934 (N_5934,In_2065,In_794);
and U5935 (N_5935,In_472,In_869);
or U5936 (N_5936,In_1116,In_1908);
and U5937 (N_5937,In_1713,In_1843);
xor U5938 (N_5938,In_1838,In_1369);
xor U5939 (N_5939,In_141,In_675);
nor U5940 (N_5940,In_1561,In_2084);
xor U5941 (N_5941,In_2284,In_1379);
or U5942 (N_5942,In_775,In_1182);
and U5943 (N_5943,In_935,In_461);
or U5944 (N_5944,In_207,In_1847);
nor U5945 (N_5945,In_930,In_1092);
and U5946 (N_5946,In_886,In_2177);
nor U5947 (N_5947,In_1310,In_15);
nand U5948 (N_5948,In_1937,In_1663);
and U5949 (N_5949,In_1990,In_284);
nor U5950 (N_5950,In_299,In_2045);
or U5951 (N_5951,In_1485,In_1779);
or U5952 (N_5952,In_1772,In_1072);
xnor U5953 (N_5953,In_374,In_907);
nand U5954 (N_5954,In_2101,In_698);
nand U5955 (N_5955,In_2218,In_2350);
and U5956 (N_5956,In_599,In_587);
nand U5957 (N_5957,In_123,In_722);
nand U5958 (N_5958,In_1028,In_1363);
nor U5959 (N_5959,In_1832,In_1947);
nand U5960 (N_5960,In_1099,In_333);
or U5961 (N_5961,In_642,In_1765);
nand U5962 (N_5962,In_1412,In_713);
and U5963 (N_5963,In_2123,In_1162);
xnor U5964 (N_5964,In_2198,In_1106);
or U5965 (N_5965,In_2118,In_642);
and U5966 (N_5966,In_39,In_719);
or U5967 (N_5967,In_2256,In_1732);
and U5968 (N_5968,In_2099,In_708);
or U5969 (N_5969,In_696,In_1037);
or U5970 (N_5970,In_727,In_1561);
nor U5971 (N_5971,In_1871,In_813);
or U5972 (N_5972,In_800,In_54);
or U5973 (N_5973,In_2080,In_1559);
nand U5974 (N_5974,In_1569,In_1718);
xnor U5975 (N_5975,In_1380,In_1057);
and U5976 (N_5976,In_1236,In_2215);
nor U5977 (N_5977,In_404,In_1713);
nor U5978 (N_5978,In_313,In_1066);
and U5979 (N_5979,In_1455,In_527);
or U5980 (N_5980,In_658,In_612);
and U5981 (N_5981,In_1327,In_710);
and U5982 (N_5982,In_1306,In_201);
and U5983 (N_5983,In_1595,In_195);
or U5984 (N_5984,In_653,In_1369);
nand U5985 (N_5985,In_953,In_716);
or U5986 (N_5986,In_2060,In_123);
and U5987 (N_5987,In_708,In_2198);
or U5988 (N_5988,In_1835,In_1821);
and U5989 (N_5989,In_1073,In_2181);
xnor U5990 (N_5990,In_1040,In_2103);
nor U5991 (N_5991,In_1144,In_555);
or U5992 (N_5992,In_1052,In_1140);
and U5993 (N_5993,In_630,In_1236);
xnor U5994 (N_5994,In_17,In_1879);
or U5995 (N_5995,In_1198,In_2389);
or U5996 (N_5996,In_1590,In_153);
nand U5997 (N_5997,In_1711,In_2495);
nand U5998 (N_5998,In_1344,In_287);
or U5999 (N_5999,In_1802,In_2259);
nand U6000 (N_6000,In_1455,In_71);
nor U6001 (N_6001,In_2308,In_2356);
or U6002 (N_6002,In_1603,In_1729);
and U6003 (N_6003,In_632,In_603);
nand U6004 (N_6004,In_2121,In_374);
and U6005 (N_6005,In_763,In_1372);
nand U6006 (N_6006,In_902,In_1066);
or U6007 (N_6007,In_1271,In_285);
nor U6008 (N_6008,In_931,In_2037);
nor U6009 (N_6009,In_346,In_1244);
and U6010 (N_6010,In_742,In_1978);
nor U6011 (N_6011,In_672,In_1941);
nor U6012 (N_6012,In_187,In_1278);
nand U6013 (N_6013,In_1142,In_2079);
xor U6014 (N_6014,In_2107,In_1945);
and U6015 (N_6015,In_1716,In_1547);
or U6016 (N_6016,In_1853,In_259);
nor U6017 (N_6017,In_1644,In_1182);
or U6018 (N_6018,In_1786,In_1293);
nor U6019 (N_6019,In_1820,In_2105);
nand U6020 (N_6020,In_1047,In_158);
or U6021 (N_6021,In_1271,In_1442);
nand U6022 (N_6022,In_2030,In_2063);
or U6023 (N_6023,In_1385,In_198);
nand U6024 (N_6024,In_2497,In_1905);
or U6025 (N_6025,In_133,In_1401);
or U6026 (N_6026,In_275,In_1100);
or U6027 (N_6027,In_38,In_935);
or U6028 (N_6028,In_1529,In_1883);
and U6029 (N_6029,In_378,In_105);
nand U6030 (N_6030,In_2060,In_922);
nor U6031 (N_6031,In_2332,In_1375);
or U6032 (N_6032,In_196,In_1688);
and U6033 (N_6033,In_1059,In_710);
or U6034 (N_6034,In_2323,In_647);
and U6035 (N_6035,In_1475,In_2480);
nor U6036 (N_6036,In_555,In_29);
xor U6037 (N_6037,In_397,In_528);
or U6038 (N_6038,In_417,In_542);
nor U6039 (N_6039,In_1238,In_1163);
and U6040 (N_6040,In_288,In_1133);
nor U6041 (N_6041,In_2461,In_1320);
nor U6042 (N_6042,In_426,In_2001);
and U6043 (N_6043,In_515,In_1408);
nand U6044 (N_6044,In_1798,In_497);
nand U6045 (N_6045,In_1220,In_653);
nor U6046 (N_6046,In_1657,In_915);
or U6047 (N_6047,In_1274,In_512);
xnor U6048 (N_6048,In_1968,In_1221);
and U6049 (N_6049,In_2204,In_2054);
nor U6050 (N_6050,In_1732,In_2285);
or U6051 (N_6051,In_1908,In_408);
nand U6052 (N_6052,In_853,In_95);
and U6053 (N_6053,In_2376,In_1384);
nor U6054 (N_6054,In_2205,In_1037);
or U6055 (N_6055,In_45,In_1537);
and U6056 (N_6056,In_1093,In_2479);
or U6057 (N_6057,In_919,In_1247);
nor U6058 (N_6058,In_1646,In_877);
nand U6059 (N_6059,In_2163,In_1780);
nor U6060 (N_6060,In_137,In_305);
xnor U6061 (N_6061,In_242,In_309);
or U6062 (N_6062,In_1382,In_1366);
nand U6063 (N_6063,In_583,In_1673);
and U6064 (N_6064,In_2324,In_1713);
nand U6065 (N_6065,In_1583,In_629);
nand U6066 (N_6066,In_747,In_1537);
or U6067 (N_6067,In_1296,In_1970);
nor U6068 (N_6068,In_1283,In_1978);
nor U6069 (N_6069,In_278,In_2233);
nand U6070 (N_6070,In_2287,In_1289);
nor U6071 (N_6071,In_84,In_378);
xor U6072 (N_6072,In_1587,In_2490);
nor U6073 (N_6073,In_1242,In_1453);
xor U6074 (N_6074,In_1319,In_1677);
nor U6075 (N_6075,In_962,In_1983);
nor U6076 (N_6076,In_661,In_711);
or U6077 (N_6077,In_2357,In_1298);
or U6078 (N_6078,In_2095,In_2397);
nor U6079 (N_6079,In_1394,In_1422);
and U6080 (N_6080,In_1680,In_389);
and U6081 (N_6081,In_575,In_347);
or U6082 (N_6082,In_1240,In_1216);
nor U6083 (N_6083,In_1113,In_1881);
and U6084 (N_6084,In_1877,In_895);
nor U6085 (N_6085,In_2317,In_1765);
nor U6086 (N_6086,In_2096,In_1138);
and U6087 (N_6087,In_1572,In_502);
or U6088 (N_6088,In_683,In_1270);
nand U6089 (N_6089,In_646,In_1890);
and U6090 (N_6090,In_2374,In_980);
and U6091 (N_6091,In_732,In_225);
nor U6092 (N_6092,In_1318,In_789);
or U6093 (N_6093,In_2017,In_1657);
nand U6094 (N_6094,In_2455,In_239);
nand U6095 (N_6095,In_2000,In_2437);
or U6096 (N_6096,In_1516,In_1963);
nand U6097 (N_6097,In_802,In_1414);
and U6098 (N_6098,In_1015,In_2418);
or U6099 (N_6099,In_1173,In_1287);
nand U6100 (N_6100,In_2286,In_361);
and U6101 (N_6101,In_1877,In_713);
xor U6102 (N_6102,In_1441,In_420);
and U6103 (N_6103,In_1866,In_378);
nand U6104 (N_6104,In_1625,In_1934);
and U6105 (N_6105,In_2106,In_70);
nor U6106 (N_6106,In_1046,In_1551);
and U6107 (N_6107,In_1954,In_368);
nand U6108 (N_6108,In_1152,In_2057);
nor U6109 (N_6109,In_1888,In_579);
and U6110 (N_6110,In_1151,In_396);
nor U6111 (N_6111,In_790,In_1708);
nor U6112 (N_6112,In_1149,In_1693);
nand U6113 (N_6113,In_267,In_2381);
and U6114 (N_6114,In_1847,In_279);
or U6115 (N_6115,In_2059,In_1254);
and U6116 (N_6116,In_273,In_992);
nand U6117 (N_6117,In_2159,In_2251);
nand U6118 (N_6118,In_1881,In_2338);
nand U6119 (N_6119,In_545,In_698);
or U6120 (N_6120,In_796,In_1764);
nor U6121 (N_6121,In_1231,In_1663);
or U6122 (N_6122,In_1394,In_2079);
nor U6123 (N_6123,In_1956,In_1585);
nor U6124 (N_6124,In_1665,In_832);
nand U6125 (N_6125,In_1168,In_1623);
nand U6126 (N_6126,In_662,In_51);
nand U6127 (N_6127,In_1122,In_188);
or U6128 (N_6128,In_1664,In_1426);
or U6129 (N_6129,In_2363,In_11);
nor U6130 (N_6130,In_1284,In_2026);
and U6131 (N_6131,In_1346,In_1382);
nor U6132 (N_6132,In_447,In_2162);
and U6133 (N_6133,In_193,In_2188);
or U6134 (N_6134,In_2169,In_1557);
and U6135 (N_6135,In_294,In_920);
and U6136 (N_6136,In_761,In_227);
nor U6137 (N_6137,In_2346,In_1068);
and U6138 (N_6138,In_1385,In_1689);
nor U6139 (N_6139,In_1108,In_753);
and U6140 (N_6140,In_1210,In_928);
xor U6141 (N_6141,In_870,In_2182);
and U6142 (N_6142,In_408,In_1913);
nor U6143 (N_6143,In_2176,In_1818);
or U6144 (N_6144,In_1069,In_1413);
and U6145 (N_6145,In_504,In_700);
nor U6146 (N_6146,In_2311,In_804);
and U6147 (N_6147,In_108,In_1431);
nor U6148 (N_6148,In_1855,In_1431);
and U6149 (N_6149,In_1875,In_194);
and U6150 (N_6150,In_1019,In_2308);
nand U6151 (N_6151,In_1254,In_2439);
or U6152 (N_6152,In_2283,In_443);
or U6153 (N_6153,In_1596,In_1730);
xnor U6154 (N_6154,In_2336,In_751);
and U6155 (N_6155,In_1899,In_1444);
nor U6156 (N_6156,In_1721,In_846);
nor U6157 (N_6157,In_879,In_954);
nand U6158 (N_6158,In_449,In_1790);
and U6159 (N_6159,In_1997,In_1297);
xor U6160 (N_6160,In_2215,In_2093);
nand U6161 (N_6161,In_1428,In_82);
nor U6162 (N_6162,In_1170,In_1520);
and U6163 (N_6163,In_2414,In_2232);
or U6164 (N_6164,In_285,In_1147);
or U6165 (N_6165,In_2009,In_794);
xor U6166 (N_6166,In_538,In_1853);
nor U6167 (N_6167,In_1371,In_1265);
xnor U6168 (N_6168,In_542,In_1923);
or U6169 (N_6169,In_1330,In_2147);
nor U6170 (N_6170,In_1001,In_1365);
or U6171 (N_6171,In_1348,In_1167);
or U6172 (N_6172,In_1575,In_450);
nand U6173 (N_6173,In_166,In_906);
or U6174 (N_6174,In_1060,In_2315);
or U6175 (N_6175,In_1313,In_1548);
or U6176 (N_6176,In_1182,In_778);
or U6177 (N_6177,In_79,In_1427);
or U6178 (N_6178,In_669,In_1893);
or U6179 (N_6179,In_2003,In_505);
and U6180 (N_6180,In_857,In_6);
nand U6181 (N_6181,In_2093,In_2056);
xor U6182 (N_6182,In_7,In_1698);
nor U6183 (N_6183,In_285,In_2135);
xor U6184 (N_6184,In_826,In_2222);
or U6185 (N_6185,In_1917,In_1844);
and U6186 (N_6186,In_2118,In_2148);
nand U6187 (N_6187,In_2332,In_1685);
nor U6188 (N_6188,In_1834,In_548);
nand U6189 (N_6189,In_487,In_342);
and U6190 (N_6190,In_1925,In_2488);
nor U6191 (N_6191,In_752,In_883);
and U6192 (N_6192,In_861,In_1761);
nor U6193 (N_6193,In_1103,In_1785);
nor U6194 (N_6194,In_1604,In_2446);
or U6195 (N_6195,In_10,In_2386);
and U6196 (N_6196,In_1121,In_1775);
or U6197 (N_6197,In_1153,In_1704);
nand U6198 (N_6198,In_969,In_925);
nor U6199 (N_6199,In_1278,In_709);
nand U6200 (N_6200,In_620,In_278);
nor U6201 (N_6201,In_2117,In_1329);
or U6202 (N_6202,In_1517,In_1333);
nor U6203 (N_6203,In_2035,In_2290);
nand U6204 (N_6204,In_1407,In_1109);
nor U6205 (N_6205,In_2260,In_1608);
or U6206 (N_6206,In_2059,In_883);
or U6207 (N_6207,In_1964,In_178);
nor U6208 (N_6208,In_717,In_711);
or U6209 (N_6209,In_2211,In_258);
nand U6210 (N_6210,In_500,In_1819);
or U6211 (N_6211,In_1136,In_1621);
nor U6212 (N_6212,In_1825,In_81);
and U6213 (N_6213,In_963,In_1517);
nand U6214 (N_6214,In_449,In_150);
xnor U6215 (N_6215,In_2333,In_668);
and U6216 (N_6216,In_2468,In_1933);
and U6217 (N_6217,In_34,In_1919);
and U6218 (N_6218,In_1969,In_151);
nor U6219 (N_6219,In_528,In_1853);
nand U6220 (N_6220,In_2221,In_1646);
and U6221 (N_6221,In_1793,In_986);
nor U6222 (N_6222,In_462,In_2155);
nor U6223 (N_6223,In_330,In_2201);
nand U6224 (N_6224,In_683,In_1155);
and U6225 (N_6225,In_2410,In_1155);
nand U6226 (N_6226,In_2193,In_423);
and U6227 (N_6227,In_689,In_397);
xor U6228 (N_6228,In_521,In_842);
nand U6229 (N_6229,In_700,In_1508);
nand U6230 (N_6230,In_2465,In_582);
nand U6231 (N_6231,In_1488,In_1425);
nor U6232 (N_6232,In_2088,In_774);
or U6233 (N_6233,In_1128,In_1925);
nor U6234 (N_6234,In_1656,In_941);
or U6235 (N_6235,In_2385,In_2330);
nand U6236 (N_6236,In_1084,In_587);
nand U6237 (N_6237,In_850,In_1394);
nand U6238 (N_6238,In_1204,In_1325);
nor U6239 (N_6239,In_1992,In_448);
or U6240 (N_6240,In_2158,In_1888);
and U6241 (N_6241,In_1698,In_354);
nand U6242 (N_6242,In_132,In_1535);
or U6243 (N_6243,In_1662,In_1418);
nand U6244 (N_6244,In_2172,In_2465);
or U6245 (N_6245,In_2273,In_1661);
nor U6246 (N_6246,In_1421,In_941);
nor U6247 (N_6247,In_1243,In_2248);
nor U6248 (N_6248,In_478,In_1384);
nand U6249 (N_6249,In_622,In_943);
xnor U6250 (N_6250,N_2775,N_3885);
and U6251 (N_6251,N_2509,N_3051);
and U6252 (N_6252,N_3679,N_4618);
nand U6253 (N_6253,N_5123,N_4504);
and U6254 (N_6254,N_5373,N_1920);
or U6255 (N_6255,N_4837,N_5712);
and U6256 (N_6256,N_3862,N_4942);
xor U6257 (N_6257,N_2979,N_1072);
nand U6258 (N_6258,N_4763,N_388);
xnor U6259 (N_6259,N_1437,N_2967);
or U6260 (N_6260,N_830,N_1832);
nand U6261 (N_6261,N_1674,N_4620);
and U6262 (N_6262,N_3800,N_4143);
nor U6263 (N_6263,N_5028,N_733);
or U6264 (N_6264,N_4779,N_5549);
or U6265 (N_6265,N_597,N_309);
nor U6266 (N_6266,N_2095,N_5249);
nor U6267 (N_6267,N_3280,N_1107);
or U6268 (N_6268,N_2001,N_4909);
or U6269 (N_6269,N_104,N_5739);
nor U6270 (N_6270,N_4768,N_886);
or U6271 (N_6271,N_5466,N_2200);
nor U6272 (N_6272,N_3557,N_478);
nand U6273 (N_6273,N_4315,N_5576);
and U6274 (N_6274,N_2487,N_2286);
or U6275 (N_6275,N_5047,N_1543);
and U6276 (N_6276,N_4794,N_2124);
or U6277 (N_6277,N_6197,N_1830);
nor U6278 (N_6278,N_3855,N_4156);
and U6279 (N_6279,N_4722,N_383);
nand U6280 (N_6280,N_4624,N_1536);
and U6281 (N_6281,N_617,N_1957);
nor U6282 (N_6282,N_2619,N_2941);
and U6283 (N_6283,N_422,N_3389);
nor U6284 (N_6284,N_3619,N_804);
nand U6285 (N_6285,N_5207,N_4895);
nor U6286 (N_6286,N_344,N_5338);
nor U6287 (N_6287,N_1296,N_3154);
nor U6288 (N_6288,N_2350,N_4542);
or U6289 (N_6289,N_696,N_223);
or U6290 (N_6290,N_3661,N_3024);
and U6291 (N_6291,N_955,N_3041);
nand U6292 (N_6292,N_1394,N_5565);
or U6293 (N_6293,N_3572,N_2503);
nand U6294 (N_6294,N_4865,N_45);
xor U6295 (N_6295,N_6096,N_576);
nand U6296 (N_6296,N_3350,N_1804);
nand U6297 (N_6297,N_559,N_1639);
and U6298 (N_6298,N_2860,N_2249);
xnor U6299 (N_6299,N_1343,N_2910);
and U6300 (N_6300,N_6043,N_2114);
nor U6301 (N_6301,N_789,N_2376);
or U6302 (N_6302,N_937,N_4258);
xor U6303 (N_6303,N_2752,N_5305);
nor U6304 (N_6304,N_4426,N_1602);
or U6305 (N_6305,N_4372,N_4662);
and U6306 (N_6306,N_3006,N_4547);
nor U6307 (N_6307,N_3502,N_5837);
or U6308 (N_6308,N_869,N_2318);
nand U6309 (N_6309,N_3105,N_3636);
nor U6310 (N_6310,N_4767,N_5720);
or U6311 (N_6311,N_6149,N_5064);
nor U6312 (N_6312,N_2292,N_2966);
nand U6313 (N_6313,N_5529,N_2531);
nor U6314 (N_6314,N_5211,N_1635);
and U6315 (N_6315,N_3137,N_2595);
nor U6316 (N_6316,N_2079,N_379);
xnor U6317 (N_6317,N_834,N_3090);
nor U6318 (N_6318,N_1211,N_5450);
and U6319 (N_6319,N_2485,N_4911);
or U6320 (N_6320,N_5954,N_2477);
nor U6321 (N_6321,N_4700,N_5875);
nand U6322 (N_6322,N_82,N_3171);
or U6323 (N_6323,N_2794,N_289);
xor U6324 (N_6324,N_1295,N_2605);
nand U6325 (N_6325,N_5031,N_5844);
xor U6326 (N_6326,N_2285,N_4864);
and U6327 (N_6327,N_1553,N_4020);
or U6328 (N_6328,N_5803,N_5397);
nor U6329 (N_6329,N_115,N_2068);
or U6330 (N_6330,N_5796,N_4607);
xnor U6331 (N_6331,N_3963,N_103);
nor U6332 (N_6332,N_5806,N_5676);
nand U6333 (N_6333,N_3829,N_1098);
or U6334 (N_6334,N_6203,N_4306);
or U6335 (N_6335,N_4399,N_1392);
nand U6336 (N_6336,N_978,N_1722);
nand U6337 (N_6337,N_5560,N_4245);
and U6338 (N_6338,N_5000,N_1627);
nor U6339 (N_6339,N_34,N_6116);
nor U6340 (N_6340,N_1452,N_4450);
nand U6341 (N_6341,N_4925,N_831);
nor U6342 (N_6342,N_6156,N_753);
nor U6343 (N_6343,N_1003,N_3040);
xnor U6344 (N_6344,N_1236,N_1310);
nor U6345 (N_6345,N_2626,N_3003);
and U6346 (N_6346,N_3723,N_5876);
or U6347 (N_6347,N_3846,N_4995);
or U6348 (N_6348,N_4378,N_4192);
nor U6349 (N_6349,N_3352,N_1616);
or U6350 (N_6350,N_5361,N_4477);
or U6351 (N_6351,N_1378,N_4047);
and U6352 (N_6352,N_612,N_1008);
nand U6353 (N_6353,N_349,N_432);
nor U6354 (N_6354,N_4848,N_2521);
and U6355 (N_6355,N_1477,N_469);
or U6356 (N_6356,N_4751,N_6076);
or U6357 (N_6357,N_137,N_4968);
nand U6358 (N_6358,N_2107,N_5180);
nand U6359 (N_6359,N_3929,N_4106);
nand U6360 (N_6360,N_5777,N_2528);
nor U6361 (N_6361,N_1807,N_2909);
xnor U6362 (N_6362,N_2141,N_3703);
nor U6363 (N_6363,N_248,N_4736);
nand U6364 (N_6364,N_4010,N_1658);
nor U6365 (N_6365,N_3711,N_2137);
nand U6366 (N_6366,N_3663,N_4976);
nand U6367 (N_6367,N_3984,N_6169);
or U6368 (N_6368,N_5723,N_5307);
and U6369 (N_6369,N_1117,N_3252);
nand U6370 (N_6370,N_748,N_2188);
nor U6371 (N_6371,N_2706,N_4654);
or U6372 (N_6372,N_2639,N_4184);
nand U6373 (N_6373,N_3841,N_3744);
and U6374 (N_6374,N_993,N_3313);
nand U6375 (N_6375,N_3191,N_3119);
nor U6376 (N_6376,N_35,N_3382);
and U6377 (N_6377,N_5581,N_6142);
or U6378 (N_6378,N_5497,N_3604);
and U6379 (N_6379,N_2519,N_5944);
nor U6380 (N_6380,N_2482,N_3466);
nand U6381 (N_6381,N_1710,N_2307);
nor U6382 (N_6382,N_215,N_4612);
nand U6383 (N_6383,N_4369,N_1732);
and U6384 (N_6384,N_4539,N_6123);
nor U6385 (N_6385,N_393,N_4127);
or U6386 (N_6386,N_4469,N_4592);
nor U6387 (N_6387,N_287,N_3290);
nor U6388 (N_6388,N_5543,N_970);
nor U6389 (N_6389,N_6029,N_2510);
or U6390 (N_6390,N_1007,N_722);
nor U6391 (N_6391,N_4064,N_5569);
nor U6392 (N_6392,N_909,N_5515);
nand U6393 (N_6393,N_1390,N_6082);
and U6394 (N_6394,N_2683,N_5807);
and U6395 (N_6395,N_2102,N_2214);
nand U6396 (N_6396,N_3315,N_2208);
nor U6397 (N_6397,N_1141,N_4559);
nor U6398 (N_6398,N_2974,N_2806);
or U6399 (N_6399,N_589,N_2555);
or U6400 (N_6400,N_2624,N_3305);
or U6401 (N_6401,N_4596,N_4648);
or U6402 (N_6402,N_6120,N_2237);
nand U6403 (N_6403,N_3426,N_5978);
nor U6404 (N_6404,N_163,N_945);
and U6405 (N_6405,N_2197,N_15);
nor U6406 (N_6406,N_854,N_2828);
nand U6407 (N_6407,N_3153,N_3416);
xor U6408 (N_6408,N_4550,N_210);
xnor U6409 (N_6409,N_3458,N_3949);
nor U6410 (N_6410,N_4820,N_2646);
or U6411 (N_6411,N_2972,N_2106);
nor U6412 (N_6412,N_4874,N_1179);
xnor U6413 (N_6413,N_1982,N_3671);
xor U6414 (N_6414,N_4214,N_1865);
nor U6415 (N_6415,N_3830,N_4876);
or U6416 (N_6416,N_5622,N_3825);
nand U6417 (N_6417,N_3785,N_1103);
nand U6418 (N_6418,N_3344,N_2354);
or U6419 (N_6419,N_3774,N_4919);
and U6420 (N_6420,N_4021,N_4923);
nand U6421 (N_6421,N_683,N_601);
nor U6422 (N_6422,N_4415,N_592);
and U6423 (N_6423,N_5069,N_6212);
and U6424 (N_6424,N_4471,N_21);
xnor U6425 (N_6425,N_2699,N_3658);
or U6426 (N_6426,N_5275,N_4553);
nand U6427 (N_6427,N_1403,N_2193);
or U6428 (N_6428,N_4797,N_5282);
nor U6429 (N_6429,N_2695,N_906);
and U6430 (N_6430,N_38,N_418);
nand U6431 (N_6431,N_4501,N_1245);
xnor U6432 (N_6432,N_3307,N_3987);
nand U6433 (N_6433,N_2504,N_4734);
and U6434 (N_6434,N_1829,N_1596);
and U6435 (N_6435,N_2623,N_4357);
nand U6436 (N_6436,N_3113,N_2257);
or U6437 (N_6437,N_1540,N_3092);
or U6438 (N_6438,N_5388,N_4176);
and U6439 (N_6439,N_2118,N_2568);
or U6440 (N_6440,N_5360,N_1928);
and U6441 (N_6441,N_5879,N_439);
or U6442 (N_6442,N_2344,N_1479);
xnor U6443 (N_6443,N_5034,N_3775);
nor U6444 (N_6444,N_5626,N_4151);
or U6445 (N_6445,N_936,N_5118);
xor U6446 (N_6446,N_4237,N_3245);
and U6447 (N_6447,N_4094,N_2147);
and U6448 (N_6448,N_1538,N_1905);
nor U6449 (N_6449,N_2630,N_278);
or U6450 (N_6450,N_843,N_4628);
nand U6451 (N_6451,N_4500,N_3194);
nand U6452 (N_6452,N_2332,N_3170);
or U6453 (N_6453,N_914,N_868);
and U6454 (N_6454,N_6119,N_5753);
nor U6455 (N_6455,N_5598,N_2043);
nand U6456 (N_6456,N_4702,N_1853);
xor U6457 (N_6457,N_5802,N_2406);
or U6458 (N_6458,N_5415,N_2685);
nor U6459 (N_6459,N_810,N_5218);
nand U6460 (N_6460,N_1426,N_520);
xnor U6461 (N_6461,N_308,N_579);
and U6462 (N_6462,N_5062,N_4470);
or U6463 (N_6463,N_5080,N_4247);
or U6464 (N_6464,N_5903,N_3962);
and U6465 (N_6465,N_4377,N_4164);
and U6466 (N_6466,N_515,N_341);
nand U6467 (N_6467,N_1660,N_2557);
nor U6468 (N_6468,N_1498,N_1637);
nand U6469 (N_6469,N_3385,N_2917);
nor U6470 (N_6470,N_5268,N_0);
nand U6471 (N_6471,N_2898,N_4045);
and U6472 (N_6472,N_259,N_1719);
and U6473 (N_6473,N_3147,N_706);
nand U6474 (N_6474,N_5151,N_5328);
and U6475 (N_6475,N_4342,N_4479);
and U6476 (N_6476,N_4849,N_6041);
nor U6477 (N_6477,N_4997,N_4059);
xor U6478 (N_6478,N_3882,N_3014);
xor U6479 (N_6479,N_5910,N_5181);
nand U6480 (N_6480,N_3367,N_3716);
and U6481 (N_6481,N_5776,N_1899);
nor U6482 (N_6482,N_4095,N_5446);
or U6483 (N_6483,N_1551,N_1988);
and U6484 (N_6484,N_76,N_5434);
nand U6485 (N_6485,N_5725,N_3048);
or U6486 (N_6486,N_5502,N_3169);
or U6487 (N_6487,N_3083,N_5773);
nand U6488 (N_6488,N_1778,N_3594);
nand U6489 (N_6489,N_5744,N_5857);
and U6490 (N_6490,N_1466,N_2842);
and U6491 (N_6491,N_5110,N_3116);
or U6492 (N_6492,N_3750,N_5436);
and U6493 (N_6493,N_2621,N_5286);
and U6494 (N_6494,N_1385,N_508);
or U6495 (N_6495,N_2629,N_5669);
or U6496 (N_6496,N_5741,N_1872);
xor U6497 (N_6497,N_5510,N_3482);
and U6498 (N_6498,N_3700,N_5940);
nor U6499 (N_6499,N_1401,N_1659);
nor U6500 (N_6500,N_2361,N_386);
nand U6501 (N_6501,N_2936,N_6221);
and U6502 (N_6502,N_4616,N_2186);
or U6503 (N_6503,N_1070,N_3507);
or U6504 (N_6504,N_2539,N_197);
nand U6505 (N_6505,N_3889,N_2299);
nand U6506 (N_6506,N_2881,N_1562);
and U6507 (N_6507,N_4979,N_4460);
or U6508 (N_6508,N_3141,N_3600);
and U6509 (N_6509,N_5912,N_5748);
nand U6510 (N_6510,N_3834,N_5824);
xnor U6511 (N_6511,N_5981,N_5775);
and U6512 (N_6512,N_2378,N_2349);
and U6513 (N_6513,N_981,N_2236);
or U6514 (N_6514,N_790,N_3017);
nand U6515 (N_6515,N_74,N_2494);
and U6516 (N_6516,N_2261,N_3251);
and U6517 (N_6517,N_3945,N_4326);
nand U6518 (N_6518,N_2665,N_4368);
xnor U6519 (N_6519,N_4379,N_5813);
nand U6520 (N_6520,N_3523,N_802);
nor U6521 (N_6521,N_4103,N_2949);
xor U6522 (N_6522,N_853,N_258);
nand U6523 (N_6523,N_4906,N_2224);
nor U6524 (N_6524,N_1874,N_5325);
nor U6525 (N_6525,N_2761,N_3522);
and U6526 (N_6526,N_561,N_4945);
and U6527 (N_6527,N_2222,N_986);
xnor U6528 (N_6528,N_95,N_2758);
nand U6529 (N_6529,N_879,N_3802);
xnor U6530 (N_6530,N_1011,N_6248);
or U6531 (N_6531,N_3735,N_5461);
nor U6532 (N_6532,N_3903,N_3418);
nor U6533 (N_6533,N_6154,N_898);
or U6534 (N_6534,N_252,N_3563);
nand U6535 (N_6535,N_3743,N_6222);
and U6536 (N_6536,N_5804,N_2462);
nand U6537 (N_6537,N_5304,N_54);
or U6538 (N_6538,N_5900,N_972);
nor U6539 (N_6539,N_5977,N_2074);
and U6540 (N_6540,N_2204,N_1279);
nand U6541 (N_6541,N_4370,N_1699);
nor U6542 (N_6542,N_3104,N_4586);
nand U6543 (N_6543,N_3964,N_6239);
nor U6544 (N_6544,N_6025,N_4916);
nand U6545 (N_6545,N_364,N_5052);
or U6546 (N_6546,N_5347,N_5293);
and U6547 (N_6547,N_1074,N_5234);
or U6548 (N_6548,N_2862,N_5699);
or U6549 (N_6549,N_3731,N_4673);
nand U6550 (N_6550,N_4299,N_5623);
nor U6551 (N_6551,N_2723,N_484);
and U6552 (N_6552,N_4135,N_4287);
nand U6553 (N_6553,N_3863,N_25);
nand U6554 (N_6554,N_3215,N_4692);
nor U6555 (N_6555,N_784,N_660);
and U6556 (N_6556,N_2496,N_1788);
and U6557 (N_6557,N_97,N_1673);
and U6558 (N_6558,N_2316,N_4381);
nand U6559 (N_6559,N_4220,N_5367);
nor U6560 (N_6560,N_4271,N_6118);
nor U6561 (N_6561,N_2081,N_1075);
and U6562 (N_6562,N_3796,N_4527);
nor U6563 (N_6563,N_3675,N_3577);
nor U6564 (N_6564,N_4867,N_3438);
nor U6565 (N_6565,N_2438,N_581);
and U6566 (N_6566,N_6134,N_166);
xor U6567 (N_6567,N_300,N_5170);
or U6568 (N_6568,N_4255,N_5897);
nor U6569 (N_6569,N_984,N_4729);
or U6570 (N_6570,N_3339,N_4826);
or U6571 (N_6571,N_1305,N_608);
nor U6572 (N_6572,N_497,N_5649);
or U6573 (N_6573,N_1294,N_4549);
nand U6574 (N_6574,N_3455,N_1340);
and U6575 (N_6575,N_1453,N_1791);
or U6576 (N_6576,N_5274,N_1055);
nand U6577 (N_6577,N_4157,N_1285);
nand U6578 (N_6578,N_3901,N_119);
xor U6579 (N_6579,N_889,N_1106);
nand U6580 (N_6580,N_1777,N_4562);
nor U6581 (N_6581,N_5348,N_3471);
nand U6582 (N_6582,N_912,N_5345);
nor U6583 (N_6583,N_4614,N_5054);
nand U6584 (N_6584,N_6168,N_2045);
nor U6585 (N_6585,N_2433,N_5276);
or U6586 (N_6586,N_4108,N_4811);
xor U6587 (N_6587,N_141,N_3612);
xor U6588 (N_6588,N_3032,N_4728);
nand U6589 (N_6589,N_5866,N_57);
or U6590 (N_6590,N_151,N_5511);
nor U6591 (N_6591,N_1984,N_2122);
and U6592 (N_6592,N_4711,N_3505);
or U6593 (N_6593,N_1787,N_2090);
nor U6594 (N_6594,N_1123,N_2947);
or U6595 (N_6595,N_3564,N_5480);
xor U6596 (N_6596,N_5376,N_4420);
nand U6597 (N_6597,N_4955,N_3826);
or U6598 (N_6598,N_1578,N_2817);
or U6599 (N_6599,N_4615,N_1092);
nor U6600 (N_6600,N_1181,N_5183);
or U6601 (N_6601,N_4611,N_5267);
or U6602 (N_6602,N_2712,N_443);
or U6603 (N_6603,N_686,N_250);
xnor U6604 (N_6604,N_4881,N_4641);
and U6605 (N_6605,N_5172,N_1393);
nand U6606 (N_6606,N_1516,N_1603);
or U6607 (N_6607,N_963,N_5101);
and U6608 (N_6608,N_845,N_631);
nand U6609 (N_6609,N_5186,N_5240);
nor U6610 (N_6610,N_5722,N_2182);
nand U6611 (N_6611,N_5377,N_1135);
nand U6612 (N_6612,N_348,N_3887);
nor U6613 (N_6613,N_4522,N_4209);
or U6614 (N_6614,N_5290,N_2034);
and U6615 (N_6615,N_1046,N_950);
nand U6616 (N_6616,N_1360,N_5849);
xor U6617 (N_6617,N_883,N_3866);
or U6618 (N_6618,N_2044,N_1449);
or U6619 (N_6619,N_5996,N_5874);
or U6620 (N_6620,N_5136,N_806);
xor U6621 (N_6621,N_2388,N_3073);
or U6622 (N_6622,N_72,N_3506);
and U6623 (N_6623,N_5209,N_3983);
xor U6624 (N_6624,N_3956,N_172);
nand U6625 (N_6625,N_5507,N_5258);
xor U6626 (N_6626,N_5877,N_958);
or U6627 (N_6627,N_3157,N_267);
nor U6628 (N_6628,N_771,N_650);
and U6629 (N_6629,N_1170,N_4969);
xnor U6630 (N_6630,N_3645,N_5167);
nor U6631 (N_6631,N_1156,N_4782);
and U6632 (N_6632,N_616,N_5087);
and U6633 (N_6633,N_2781,N_3388);
or U6634 (N_6634,N_5627,N_850);
xor U6635 (N_6635,N_4425,N_5068);
nor U6636 (N_6636,N_136,N_375);
or U6637 (N_6637,N_1595,N_4502);
nor U6638 (N_6638,N_1078,N_4203);
or U6639 (N_6639,N_4484,N_2322);
and U6640 (N_6640,N_5506,N_5533);
or U6641 (N_6641,N_5930,N_6100);
and U6642 (N_6642,N_5455,N_2310);
or U6643 (N_6643,N_3749,N_1570);
nand U6644 (N_6644,N_2542,N_2488);
and U6645 (N_6645,N_1,N_2337);
nor U6646 (N_6646,N_5327,N_3688);
or U6647 (N_6647,N_2324,N_3100);
or U6648 (N_6648,N_5432,N_2096);
and U6649 (N_6649,N_1324,N_1272);
and U6650 (N_6650,N_1025,N_664);
and U6651 (N_6651,N_1921,N_1020);
nor U6652 (N_6652,N_198,N_40);
and U6653 (N_6653,N_4065,N_3115);
or U6654 (N_6654,N_1473,N_3241);
nor U6655 (N_6655,N_395,N_1851);
or U6656 (N_6656,N_5764,N_2108);
or U6657 (N_6657,N_1806,N_4558);
and U6658 (N_6658,N_1204,N_4427);
nand U6659 (N_6659,N_5901,N_5179);
nor U6660 (N_6660,N_377,N_4311);
and U6661 (N_6661,N_1188,N_6034);
or U6662 (N_6662,N_931,N_4960);
and U6663 (N_6663,N_2530,N_833);
and U6664 (N_6664,N_3609,N_6018);
nand U6665 (N_6665,N_3286,N_2328);
nor U6666 (N_6666,N_1102,N_1776);
xnor U6667 (N_6667,N_3682,N_4771);
nand U6668 (N_6668,N_4257,N_3268);
or U6669 (N_6669,N_4686,N_3478);
or U6670 (N_6670,N_3935,N_1246);
or U6671 (N_6671,N_2335,N_4971);
nand U6672 (N_6672,N_994,N_2801);
nor U6673 (N_6673,N_3182,N_4079);
nand U6674 (N_6674,N_3538,N_4605);
and U6675 (N_6675,N_5521,N_3786);
nor U6676 (N_6676,N_3222,N_4190);
nor U6677 (N_6677,N_3881,N_3155);
or U6678 (N_6678,N_3871,N_1446);
or U6679 (N_6679,N_5379,N_4468);
and U6680 (N_6680,N_1047,N_2341);
nor U6681 (N_6681,N_2975,N_2668);
nor U6682 (N_6682,N_935,N_5848);
and U6683 (N_6683,N_4147,N_6081);
or U6684 (N_6684,N_4320,N_874);
and U6685 (N_6685,N_3427,N_3257);
nand U6686 (N_6686,N_408,N_2678);
nor U6687 (N_6687,N_5614,N_3644);
and U6688 (N_6688,N_3597,N_4749);
and U6689 (N_6689,N_1044,N_1149);
nand U6690 (N_6690,N_799,N_4392);
or U6691 (N_6691,N_3321,N_3234);
nor U6692 (N_6692,N_5675,N_5225);
nand U6693 (N_6693,N_3780,N_3621);
or U6694 (N_6694,N_1654,N_638);
nor U6695 (N_6695,N_4684,N_2374);
nand U6696 (N_6696,N_233,N_3988);
nand U6697 (N_6697,N_1024,N_5872);
and U6698 (N_6698,N_3472,N_4590);
nor U6699 (N_6699,N_47,N_3);
nor U6700 (N_6700,N_5261,N_1462);
or U6701 (N_6701,N_5688,N_6104);
or U6702 (N_6702,N_4571,N_4694);
nor U6703 (N_6703,N_5702,N_5652);
and U6704 (N_6704,N_4123,N_5093);
or U6705 (N_6705,N_2814,N_2436);
nor U6706 (N_6706,N_3263,N_3611);
or U6707 (N_6707,N_1618,N_1409);
nor U6708 (N_6708,N_4980,N_1610);
and U6709 (N_6709,N_3072,N_1789);
nor U6710 (N_6710,N_3031,N_4310);
nand U6711 (N_6711,N_4827,N_4319);
and U6712 (N_6712,N_1889,N_4987);
or U6713 (N_6713,N_1239,N_871);
nand U6714 (N_6714,N_1233,N_4169);
nor U6715 (N_6715,N_3308,N_3550);
or U6716 (N_6716,N_5449,N_3993);
and U6717 (N_6717,N_1738,N_5009);
xnor U6718 (N_6718,N_3560,N_5193);
xor U6719 (N_6719,N_4754,N_78);
nand U6720 (N_6720,N_2737,N_3149);
and U6721 (N_6721,N_5458,N_5260);
xnor U6722 (N_6722,N_5931,N_2772);
or U6723 (N_6723,N_1849,N_5043);
or U6724 (N_6724,N_893,N_3250);
or U6725 (N_6725,N_2732,N_4914);
and U6726 (N_6726,N_2120,N_5154);
nor U6727 (N_6727,N_1898,N_6042);
nand U6728 (N_6728,N_5830,N_4132);
nand U6729 (N_6729,N_5314,N_3088);
nand U6730 (N_6730,N_552,N_2779);
and U6731 (N_6731,N_4073,N_5650);
nor U6732 (N_6732,N_4179,N_2207);
nand U6733 (N_6733,N_1749,N_2168);
and U6734 (N_6734,N_5474,N_5019);
nor U6735 (N_6735,N_2968,N_3973);
nor U6736 (N_6736,N_2988,N_345);
nor U6737 (N_6737,N_4516,N_2038);
nor U6738 (N_6738,N_90,N_723);
xor U6739 (N_6739,N_3705,N_3405);
or U6740 (N_6740,N_2133,N_490);
nor U6741 (N_6741,N_2019,N_4557);
nor U6742 (N_6742,N_4882,N_1461);
nor U6743 (N_6743,N_1545,N_148);
nand U6744 (N_6744,N_2183,N_1765);
or U6745 (N_6745,N_5916,N_4602);
or U6746 (N_6746,N_335,N_3199);
xnor U6747 (N_6747,N_306,N_5359);
xnor U6748 (N_6748,N_4276,N_3904);
xor U6749 (N_6749,N_6107,N_6143);
nand U6750 (N_6750,N_785,N_756);
nor U6751 (N_6751,N_1704,N_2245);
nor U6752 (N_6752,N_3186,N_4232);
nor U6753 (N_6753,N_1095,N_3428);
or U6754 (N_6754,N_691,N_5421);
nand U6755 (N_6755,N_1359,N_2437);
nand U6756 (N_6756,N_3091,N_3913);
xnor U6757 (N_6757,N_4185,N_3314);
nand U6758 (N_6758,N_3664,N_4078);
or U6759 (N_6759,N_3680,N_769);
or U6760 (N_6760,N_3287,N_4060);
xnor U6761 (N_6761,N_2961,N_4048);
or U6762 (N_6762,N_2953,N_1669);
nor U6763 (N_6763,N_6181,N_596);
nand U6764 (N_6764,N_5503,N_4125);
and U6765 (N_6765,N_2417,N_5337);
nand U6766 (N_6766,N_6158,N_6140);
nand U6767 (N_6767,N_568,N_2875);
and U6768 (N_6768,N_2375,N_5891);
and U6769 (N_6769,N_3409,N_4639);
nor U6770 (N_6770,N_5715,N_5681);
nor U6771 (N_6771,N_3236,N_3531);
or U6772 (N_6772,N_292,N_1508);
nand U6773 (N_6773,N_1624,N_2535);
and U6774 (N_6774,N_1825,N_1128);
nor U6775 (N_6775,N_2870,N_352);
nand U6776 (N_6776,N_3821,N_63);
and U6777 (N_6777,N_1754,N_3566);
or U6778 (N_6778,N_3328,N_4234);
nor U6779 (N_6779,N_2002,N_2109);
or U6780 (N_6780,N_2041,N_2423);
nor U6781 (N_6781,N_2701,N_3126);
or U6782 (N_6782,N_4894,N_3148);
and U6783 (N_6783,N_2746,N_270);
nor U6784 (N_6784,N_1283,N_1623);
nand U6785 (N_6785,N_2896,N_3767);
nand U6786 (N_6786,N_1506,N_1897);
nand U6787 (N_6787,N_713,N_1541);
nand U6788 (N_6788,N_274,N_211);
nand U6789 (N_6789,N_2424,N_1376);
xor U6790 (N_6790,N_3442,N_1199);
nor U6791 (N_6791,N_5657,N_891);
and U6792 (N_6792,N_1867,N_4747);
nor U6793 (N_6793,N_385,N_1460);
or U6794 (N_6794,N_5355,N_3473);
nand U6795 (N_6795,N_3867,N_389);
xor U6796 (N_6796,N_2872,N_4606);
and U6797 (N_6797,N_164,N_4941);
nor U6798 (N_6798,N_2522,N_5417);
nor U6799 (N_6799,N_659,N_654);
or U6800 (N_6800,N_525,N_5735);
or U6801 (N_6801,N_3080,N_7);
nor U6802 (N_6802,N_3637,N_1922);
or U6803 (N_6803,N_3578,N_594);
xor U6804 (N_6804,N_3030,N_1143);
or U6805 (N_6805,N_1282,N_933);
xnor U6806 (N_6806,N_5726,N_3527);
and U6807 (N_6807,N_3860,N_2944);
xor U6808 (N_6808,N_828,N_712);
and U6809 (N_6809,N_2931,N_2067);
or U6810 (N_6810,N_1432,N_5058);
nor U6811 (N_6811,N_89,N_5997);
nand U6812 (N_6812,N_1794,N_526);
and U6813 (N_6813,N_3582,N_4657);
or U6814 (N_6814,N_4939,N_1118);
nor U6815 (N_6815,N_4149,N_4746);
nor U6816 (N_6816,N_52,N_4859);
and U6817 (N_6817,N_1041,N_888);
nand U6818 (N_6818,N_2529,N_3589);
or U6819 (N_6819,N_5835,N_2072);
or U6820 (N_6820,N_523,N_1967);
nand U6821 (N_6821,N_382,N_2240);
nor U6822 (N_6822,N_1912,N_1517);
and U6823 (N_6823,N_825,N_661);
or U6824 (N_6824,N_3195,N_5917);
or U6825 (N_6825,N_1902,N_5370);
or U6826 (N_6826,N_5315,N_5678);
and U6827 (N_6827,N_3736,N_6215);
nor U6828 (N_6828,N_2527,N_139);
and U6829 (N_6829,N_5298,N_1225);
nand U6830 (N_6830,N_5887,N_531);
nand U6831 (N_6831,N_5423,N_5541);
nand U6832 (N_6832,N_3768,N_585);
nor U6833 (N_6833,N_2161,N_4431);
and U6834 (N_6834,N_4003,N_218);
xor U6835 (N_6835,N_1743,N_1194);
nor U6836 (N_6836,N_3961,N_6190);
or U6837 (N_6837,N_3260,N_882);
nor U6838 (N_6838,N_239,N_4845);
xor U6839 (N_6839,N_2525,N_5400);
nand U6840 (N_6840,N_3050,N_4927);
and U6841 (N_6841,N_3310,N_4810);
and U6842 (N_6842,N_3642,N_2869);
and U6843 (N_6843,N_5587,N_2368);
or U6844 (N_6844,N_1230,N_1599);
or U6845 (N_6845,N_448,N_6233);
xor U6846 (N_6846,N_4990,N_3812);
nand U6847 (N_6847,N_4396,N_4889);
and U6848 (N_6848,N_6068,N_623);
or U6849 (N_6849,N_3135,N_100);
nor U6850 (N_6850,N_2989,N_1081);
or U6851 (N_6851,N_1125,N_532);
nand U6852 (N_6852,N_1489,N_629);
nor U6853 (N_6853,N_1625,N_548);
and U6854 (N_6854,N_4296,N_4608);
nand U6855 (N_6855,N_818,N_2134);
nand U6856 (N_6856,N_2831,N_506);
nand U6857 (N_6857,N_6136,N_2533);
nor U6858 (N_6858,N_1580,N_1910);
or U6859 (N_6859,N_2065,N_3179);
or U6860 (N_6860,N_3976,N_798);
nor U6861 (N_6861,N_6179,N_2130);
and U6862 (N_6862,N_4595,N_3647);
nand U6863 (N_6863,N_5442,N_6094);
nand U6864 (N_6864,N_5077,N_5422);
nor U6865 (N_6865,N_6022,N_5021);
and U6866 (N_6866,N_2370,N_4111);
xnor U6867 (N_6867,N_4540,N_2243);
or U6868 (N_6868,N_5152,N_1567);
xor U6869 (N_6869,N_3299,N_66);
xnor U6870 (N_6870,N_5178,N_3704);
nand U6871 (N_6871,N_2929,N_1227);
nand U6872 (N_6872,N_2942,N_2778);
xor U6873 (N_6873,N_3108,N_2991);
or U6874 (N_6874,N_2631,N_1981);
nand U6875 (N_6875,N_4327,N_4703);
or U6876 (N_6876,N_1956,N_3127);
or U6877 (N_6877,N_555,N_4343);
and U6878 (N_6878,N_5869,N_2302);
nor U6879 (N_6879,N_2359,N_1307);
nor U6880 (N_6880,N_1725,N_3226);
or U6881 (N_6881,N_4948,N_5907);
and U6882 (N_6882,N_3086,N_4601);
or U6883 (N_6883,N_5612,N_181);
nand U6884 (N_6884,N_1601,N_2054);
nor U6885 (N_6885,N_39,N_2728);
or U6886 (N_6886,N_2003,N_4635);
and U6887 (N_6887,N_1191,N_2666);
xnor U6888 (N_6888,N_5718,N_2708);
and U6889 (N_6889,N_5245,N_4198);
nor U6890 (N_6890,N_3386,N_2252);
nand U6891 (N_6891,N_6183,N_2835);
nor U6892 (N_6892,N_206,N_567);
nor U6893 (N_6893,N_5295,N_3575);
and U6894 (N_6894,N_5611,N_837);
or U6895 (N_6895,N_2803,N_5424);
or U6896 (N_6896,N_2807,N_1677);
nand U6897 (N_6897,N_6157,N_1613);
and U6898 (N_6898,N_4796,N_3320);
xor U6899 (N_6899,N_5752,N_991);
nor U6900 (N_6900,N_68,N_5620);
or U6901 (N_6901,N_2866,N_1679);
nand U6902 (N_6902,N_4053,N_2753);
nand U6903 (N_6903,N_3914,N_1050);
nand U6904 (N_6904,N_3519,N_5984);
nand U6905 (N_6905,N_1254,N_116);
or U6906 (N_6906,N_1268,N_3803);
nor U6907 (N_6907,N_5696,N_1848);
nand U6908 (N_6908,N_865,N_2087);
and U6909 (N_6909,N_5670,N_3192);
nor U6910 (N_6910,N_431,N_5624);
or U6911 (N_6911,N_6247,N_3132);
nor U6912 (N_6912,N_4638,N_1638);
xnor U6913 (N_6913,N_873,N_5842);
nor U6914 (N_6914,N_5285,N_1309);
nor U6915 (N_6915,N_684,N_4617);
nand U6916 (N_6916,N_3469,N_2042);
or U6917 (N_6917,N_5629,N_3021);
nand U6918 (N_6918,N_2308,N_5750);
and U6919 (N_6919,N_5112,N_938);
nor U6920 (N_6920,N_5871,N_407);
nand U6921 (N_6921,N_5772,N_979);
or U6922 (N_6922,N_135,N_1693);
and U6923 (N_6923,N_3383,N_757);
nor U6924 (N_6924,N_1259,N_2452);
and U6925 (N_6925,N_29,N_900);
nor U6926 (N_6926,N_3552,N_3403);
nor U6927 (N_6927,N_876,N_4254);
nand U6928 (N_6928,N_2458,N_1033);
or U6929 (N_6929,N_1816,N_1260);
and U6930 (N_6930,N_5829,N_3225);
nor U6931 (N_6931,N_4546,N_1263);
and U6932 (N_6932,N_602,N_2590);
nand U6933 (N_6933,N_2442,N_173);
xor U6934 (N_6934,N_4301,N_4281);
nor U6935 (N_6935,N_1702,N_1249);
or U6936 (N_6936,N_3259,N_6173);
or U6937 (N_6937,N_5411,N_2809);
nor U6938 (N_6938,N_1844,N_2060);
nor U6939 (N_6939,N_3946,N_4362);
or U6940 (N_6940,N_1594,N_2562);
and U6941 (N_6941,N_1941,N_5852);
and U6942 (N_6942,N_6206,N_3358);
nor U6943 (N_6943,N_4455,N_3122);
and U6944 (N_6944,N_102,N_194);
nand U6945 (N_6945,N_2730,N_1326);
or U6946 (N_6946,N_2997,N_3447);
and U6947 (N_6947,N_4698,N_2690);
and U6948 (N_6948,N_3978,N_5554);
and U6949 (N_6949,N_1427,N_5029);
nor U6950 (N_6950,N_2650,N_464);
or U6951 (N_6951,N_4024,N_3659);
nand U6952 (N_6952,N_2719,N_4757);
or U6953 (N_6953,N_3591,N_146);
or U6954 (N_6954,N_4759,N_1582);
nand U6955 (N_6955,N_144,N_254);
xnor U6956 (N_6956,N_4821,N_3533);
nor U6957 (N_6957,N_2653,N_2849);
or U6958 (N_6958,N_3133,N_406);
nand U6959 (N_6959,N_3301,N_2675);
or U6960 (N_6960,N_3989,N_992);
nor U6961 (N_6961,N_3540,N_416);
nor U6962 (N_6962,N_1375,N_6069);
nor U6963 (N_6963,N_4878,N_5216);
or U6964 (N_6964,N_4262,N_6147);
nor U6965 (N_6965,N_907,N_3770);
and U6966 (N_6966,N_1809,N_1132);
nor U6967 (N_6967,N_4414,N_2689);
and U6968 (N_6968,N_1958,N_5710);
and U6969 (N_6969,N_5386,N_4272);
nand U6970 (N_6970,N_2838,N_2396);
and U6971 (N_6971,N_2269,N_5477);
nand U6972 (N_6972,N_4062,N_280);
nor U6973 (N_6973,N_613,N_3276);
nand U6974 (N_6974,N_2587,N_112);
or U6975 (N_6975,N_5289,N_5237);
xor U6976 (N_6976,N_1017,N_1676);
nor U6977 (N_6977,N_5892,N_5143);
nand U6978 (N_6978,N_3844,N_4708);
nand U6979 (N_6979,N_1766,N_249);
and U6980 (N_6980,N_4809,N_3754);
nor U6981 (N_6981,N_2589,N_2925);
nor U6982 (N_6982,N_3781,N_1989);
nand U6983 (N_6983,N_4256,N_228);
nor U6984 (N_6984,N_1171,N_2230);
xor U6985 (N_6985,N_3475,N_4439);
nor U6986 (N_6986,N_70,N_4795);
or U6987 (N_6987,N_2805,N_2478);
or U6988 (N_6988,N_1864,N_92);
and U6989 (N_6989,N_332,N_2418);
xor U6990 (N_6990,N_2507,N_120);
xnor U6991 (N_6991,N_343,N_2339);
and U6992 (N_6992,N_6037,N_483);
and U6993 (N_6993,N_5044,N_5583);
and U6994 (N_6994,N_5672,N_896);
nand U6995 (N_6995,N_4267,N_527);
or U6996 (N_6996,N_3559,N_6007);
nand U6997 (N_6997,N_5572,N_2755);
nor U6998 (N_6998,N_1406,N_692);
nor U6999 (N_6999,N_5202,N_3425);
and U7000 (N_7000,N_2747,N_4693);
nand U7001 (N_7001,N_149,N_545);
nand U7002 (N_7002,N_1110,N_2037);
xor U7003 (N_7003,N_496,N_2393);
and U7004 (N_7004,N_5165,N_3343);
or U7005 (N_7005,N_5632,N_5001);
and U7006 (N_7006,N_4261,N_3691);
and U7007 (N_7007,N_6242,N_3623);
nor U7008 (N_7008,N_4629,N_5595);
or U7009 (N_7009,N_4748,N_5965);
nor U7010 (N_7010,N_6121,N_626);
or U7011 (N_7011,N_5113,N_5816);
or U7012 (N_7012,N_4609,N_1850);
nor U7013 (N_7013,N_1189,N_2085);
nor U7014 (N_7014,N_1416,N_5730);
and U7015 (N_7015,N_4483,N_5055);
nor U7016 (N_7016,N_1895,N_2795);
nand U7017 (N_7017,N_5318,N_2721);
or U7018 (N_7018,N_2456,N_3831);
nor U7019 (N_7019,N_380,N_26);
xor U7020 (N_7020,N_5945,N_5647);
and U7021 (N_7021,N_3870,N_4581);
nand U7022 (N_7022,N_5224,N_4446);
and U7023 (N_7023,N_2847,N_4588);
nand U7024 (N_7024,N_5535,N_316);
nor U7025 (N_7025,N_3955,N_2804);
nand U7026 (N_7026,N_1563,N_4853);
nor U7027 (N_7027,N_2647,N_3532);
nor U7028 (N_7028,N_1907,N_1998);
nor U7029 (N_7029,N_1711,N_3034);
nand U7030 (N_7030,N_2360,N_1924);
or U7031 (N_7031,N_4699,N_5066);
and U7032 (N_7032,N_5390,N_5173);
nor U7033 (N_7033,N_536,N_4380);
and U7034 (N_7034,N_1652,N_1433);
nor U7035 (N_7035,N_3638,N_2352);
and U7036 (N_7036,N_240,N_5861);
and U7037 (N_7037,N_2572,N_3783);
nor U7038 (N_7038,N_5201,N_560);
nand U7039 (N_7039,N_1287,N_4631);
or U7040 (N_7040,N_3586,N_5433);
and U7041 (N_7041,N_3244,N_2963);
nand U7042 (N_7042,N_4983,N_4875);
or U7043 (N_7043,N_1820,N_2569);
nand U7044 (N_7044,N_2154,N_1940);
nor U7045 (N_7045,N_2179,N_2315);
nand U7046 (N_7046,N_3200,N_928);
or U7047 (N_7047,N_1965,N_5399);
xor U7048 (N_7048,N_620,N_5993);
or U7049 (N_7049,N_5357,N_2499);
or U7050 (N_7050,N_4801,N_651);
nor U7051 (N_7051,N_4489,N_499);
and U7052 (N_7052,N_3927,N_4839);
nand U7053 (N_7053,N_5287,N_456);
xor U7054 (N_7054,N_1184,N_5156);
nand U7055 (N_7055,N_5004,N_2213);
or U7056 (N_7056,N_5006,N_1009);
nand U7057 (N_7057,N_142,N_5233);
xor U7058 (N_7058,N_391,N_6108);
or U7059 (N_7059,N_5841,N_482);
and U7060 (N_7060,N_1105,N_961);
nor U7061 (N_7061,N_1647,N_5762);
nor U7062 (N_7062,N_14,N_1815);
xnor U7063 (N_7063,N_4511,N_3681);
and U7064 (N_7064,N_2448,N_51);
nand U7065 (N_7065,N_2945,N_2715);
or U7066 (N_7066,N_75,N_5578);
xor U7067 (N_7067,N_703,N_1785);
xor U7068 (N_7068,N_4915,N_5740);
nand U7069 (N_7069,N_2140,N_5677);
nor U7070 (N_7070,N_1687,N_1917);
nand U7071 (N_7071,N_2965,N_1499);
nor U7072 (N_7072,N_367,N_1483);
or U7073 (N_7073,N_605,N_2928);
nand U7074 (N_7074,N_977,N_366);
and U7075 (N_7075,N_360,N_2220);
or U7076 (N_7076,N_3207,N_3778);
nor U7077 (N_7077,N_178,N_1004);
nand U7078 (N_7078,N_1334,N_5760);
and U7079 (N_7079,N_1023,N_1773);
nor U7080 (N_7080,N_5589,N_4856);
or U7081 (N_7081,N_4107,N_71);
or U7082 (N_7082,N_5071,N_3701);
and U7083 (N_7083,N_3371,N_3511);
and U7084 (N_7084,N_6060,N_2904);
nand U7085 (N_7085,N_3602,N_1311);
or U7086 (N_7086,N_486,N_5880);
nand U7087 (N_7087,N_3390,N_774);
nand U7088 (N_7088,N_6148,N_3347);
xnor U7089 (N_7089,N_1976,N_5317);
nand U7090 (N_7090,N_4998,N_5405);
nand U7091 (N_7091,N_3546,N_5020);
and U7092 (N_7092,N_1834,N_3453);
xor U7093 (N_7093,N_3916,N_5539);
and U7094 (N_7094,N_4030,N_6209);
and U7095 (N_7095,N_1420,N_5065);
nand U7096 (N_7096,N_1482,N_4871);
nor U7097 (N_7097,N_4740,N_1503);
nor U7098 (N_7098,N_705,N_4400);
or U7099 (N_7099,N_5107,N_276);
or U7100 (N_7100,N_5478,N_1366);
or U7101 (N_7101,N_4696,N_5420);
xnor U7102 (N_7102,N_4634,N_3018);
nor U7103 (N_7103,N_2545,N_645);
and U7104 (N_7104,N_98,N_4695);
nand U7105 (N_7105,N_4764,N_1534);
and U7106 (N_7106,N_1474,N_5256);
and U7107 (N_7107,N_5365,N_5545);
nand U7108 (N_7108,N_1250,N_5695);
nor U7109 (N_7109,N_212,N_6224);
and U7110 (N_7110,N_5103,N_5662);
xnor U7111 (N_7111,N_1495,N_489);
xnor U7112 (N_7112,N_1488,N_668);
nor U7113 (N_7113,N_1137,N_3334);
or U7114 (N_7114,N_3922,N_6161);
and U7115 (N_7115,N_5099,N_1728);
xor U7116 (N_7116,N_1884,N_4374);
and U7117 (N_7117,N_3218,N_3931);
nor U7118 (N_7118,N_3158,N_3592);
and U7119 (N_7119,N_4096,N_3777);
and U7120 (N_7120,N_5383,N_444);
or U7121 (N_7121,N_1944,N_6178);
nand U7122 (N_7122,N_5392,N_3166);
or U7123 (N_7123,N_1026,N_2206);
nor U7124 (N_7124,N_3441,N_2276);
xnor U7125 (N_7125,N_134,N_2272);
nor U7126 (N_7126,N_3534,N_378);
nand U7127 (N_7127,N_5607,N_2672);
nand U7128 (N_7128,N_2634,N_2082);
nor U7129 (N_7129,N_803,N_3485);
and U7130 (N_7130,N_2117,N_1695);
xor U7131 (N_7131,N_3608,N_1380);
nor U7132 (N_7132,N_384,N_2460);
nor U7133 (N_7133,N_2145,N_140);
nand U7134 (N_7134,N_2296,N_376);
nor U7135 (N_7135,N_3980,N_1750);
and U7136 (N_7136,N_768,N_419);
xor U7137 (N_7137,N_1196,N_5683);
or U7138 (N_7138,N_2850,N_36);
nand U7139 (N_7139,N_2607,N_4852);
or U7140 (N_7140,N_3029,N_3355);
or U7141 (N_7141,N_3724,N_5961);
and U7142 (N_7142,N_1678,N_2383);
nor U7143 (N_7143,N_4075,N_3198);
nand U7144 (N_7144,N_4816,N_3864);
or U7145 (N_7145,N_1388,N_5326);
or U7146 (N_7146,N_2408,N_1680);
xor U7147 (N_7147,N_6056,N_2582);
nand U7148 (N_7148,N_1299,N_3574);
or U7149 (N_7149,N_2776,N_1980);
xnor U7150 (N_7150,N_1140,N_3196);
and U7151 (N_7151,N_5527,N_1344);
and U7152 (N_7152,N_1528,N_244);
and U7153 (N_7153,N_2673,N_3397);
nor U7154 (N_7154,N_633,N_5255);
or U7155 (N_7155,N_4999,N_2912);
nor U7156 (N_7156,N_582,N_985);
or U7157 (N_7157,N_4403,N_5610);
nor U7158 (N_7158,N_4838,N_2115);
and U7159 (N_7159,N_3391,N_2167);
and U7160 (N_7160,N_4704,N_6214);
or U7161 (N_7161,N_583,N_4528);
and U7162 (N_7162,N_2023,N_4181);
nand U7163 (N_7163,N_2384,N_1253);
or U7164 (N_7164,N_2932,N_5994);
or U7165 (N_7165,N_5518,N_2825);
nor U7166 (N_7166,N_1932,N_1772);
nor U7167 (N_7167,N_5500,N_1621);
nor U7168 (N_7168,N_2741,N_2667);
or U7169 (N_7169,N_5943,N_2610);
or U7170 (N_7170,N_4585,N_4544);
or U7171 (N_7171,N_1860,N_6207);
and U7172 (N_7172,N_2314,N_3246);
or U7173 (N_7173,N_3561,N_4497);
nor U7174 (N_7174,N_2094,N_4456);
or U7175 (N_7175,N_1177,N_411);
nor U7176 (N_7176,N_2158,N_4126);
nor U7177 (N_7177,N_916,N_3618);
or U7178 (N_7178,N_3937,N_3833);
or U7179 (N_7179,N_4011,N_3242);
or U7180 (N_7180,N_1331,N_521);
xor U7181 (N_7181,N_1212,N_3275);
nor U7182 (N_7182,N_3378,N_4309);
nand U7183 (N_7183,N_4317,N_4872);
and U7184 (N_7184,N_3460,N_3784);
and U7185 (N_7185,N_2579,N_5306);
and U7186 (N_7186,N_3555,N_5732);
or U7187 (N_7187,N_5540,N_1491);
or U7188 (N_7188,N_5653,N_923);
nor U7189 (N_7189,N_5825,N_3430);
nor U7190 (N_7190,N_5457,N_3950);
and U7191 (N_7191,N_5479,N_4910);
and U7192 (N_7192,N_5697,N_5135);
nand U7193 (N_7193,N_4862,N_1111);
or U7194 (N_7194,N_2994,N_1573);
nor U7195 (N_7195,N_2465,N_1206);
xnor U7196 (N_7196,N_3180,N_124);
and U7197 (N_7197,N_5435,N_4623);
and U7198 (N_7198,N_2628,N_674);
nand U7199 (N_7199,N_5641,N_18);
or U7200 (N_7200,N_811,N_1001);
and U7201 (N_7201,N_3000,N_1139);
nand U7202 (N_7202,N_1597,N_2680);
nor U7203 (N_7203,N_441,N_1060);
nand U7204 (N_7204,N_5139,N_5228);
nor U7205 (N_7205,N_2857,N_3010);
nor U7206 (N_7206,N_2718,N_510);
nand U7207 (N_7207,N_2015,N_2822);
and U7208 (N_7208,N_247,N_3793);
or U7209 (N_7209,N_724,N_3598);
nand U7210 (N_7210,N_2427,N_4228);
or U7211 (N_7211,N_209,N_5344);
or U7212 (N_7212,N_4937,N_5429);
and U7213 (N_7213,N_934,N_6102);
xor U7214 (N_7214,N_6166,N_663);
or U7215 (N_7215,N_4284,N_6128);
or U7216 (N_7216,N_1672,N_4721);
xor U7217 (N_7217,N_4089,N_4672);
nand U7218 (N_7218,N_4346,N_848);
and U7219 (N_7219,N_5097,N_4683);
nand U7220 (N_7220,N_410,N_2575);
or U7221 (N_7221,N_6196,N_4367);
nor U7222 (N_7222,N_4467,N_989);
nand U7223 (N_7223,N_4025,N_1266);
and U7224 (N_7224,N_1389,N_2709);
xnor U7225 (N_7225,N_2165,N_5684);
or U7226 (N_7226,N_982,N_1911);
nand U7227 (N_7227,N_3078,N_2209);
nor U7228 (N_7228,N_3570,N_161);
and U7229 (N_7229,N_2258,N_3738);
and U7230 (N_7230,N_3272,N_5666);
nor U7231 (N_7231,N_1575,N_1893);
and U7232 (N_7232,N_4052,N_4449);
xor U7233 (N_7233,N_473,N_4042);
nand U7234 (N_7234,N_5594,N_4627);
or U7235 (N_7235,N_1683,N_1598);
nor U7236 (N_7236,N_1763,N_4017);
and U7237 (N_7237,N_5133,N_3982);
nor U7238 (N_7238,N_4642,N_4285);
or U7239 (N_7239,N_734,N_5980);
xnor U7240 (N_7240,N_5472,N_1837);
nand U7241 (N_7241,N_566,N_4512);
and U7242 (N_7242,N_2430,N_3813);
and U7243 (N_7243,N_5036,N_5593);
nor U7244 (N_7244,N_3859,N_2098);
and U7245 (N_7245,N_1057,N_3693);
nand U7246 (N_7246,N_5942,N_1643);
and U7247 (N_7247,N_114,N_6205);
xor U7248 (N_7248,N_5196,N_3631);
or U7249 (N_7249,N_2774,N_3038);
or U7250 (N_7250,N_5878,N_3284);
nor U7251 (N_7251,N_6111,N_1737);
or U7252 (N_7252,N_4807,N_2025);
or U7253 (N_7253,N_6078,N_4888);
xor U7254 (N_7254,N_3884,N_3992);
nor U7255 (N_7255,N_2513,N_4167);
nor U7256 (N_7256,N_1226,N_763);
and U7257 (N_7257,N_586,N_3852);
and U7258 (N_7258,N_5079,N_3486);
and U7259 (N_7259,N_2643,N_4036);
nand U7260 (N_7260,N_5208,N_3452);
and U7261 (N_7261,N_2655,N_949);
and U7262 (N_7262,N_3037,N_1288);
nand U7263 (N_7263,N_2852,N_41);
xor U7264 (N_7264,N_1162,N_4411);
xor U7265 (N_7265,N_4249,N_4944);
xnor U7266 (N_7266,N_5229,N_2093);
and U7267 (N_7267,N_4398,N_3312);
nand U7268 (N_7268,N_123,N_2566);
and U7269 (N_7269,N_4982,N_4651);
or U7270 (N_7270,N_5462,N_2111);
and U7271 (N_7271,N_4177,N_2006);
xor U7272 (N_7272,N_1537,N_2964);
xor U7273 (N_7273,N_6199,N_826);
nand U7274 (N_7274,N_3408,N_1866);
nand U7275 (N_7275,N_6159,N_5160);
and U7276 (N_7276,N_6138,N_2777);
and U7277 (N_7277,N_5812,N_4793);
nor U7278 (N_7278,N_4776,N_3954);
and U7279 (N_7279,N_2560,N_5979);
nor U7280 (N_7280,N_5767,N_4733);
and U7281 (N_7281,N_59,N_4129);
or U7282 (N_7282,N_3213,N_2483);
and U7283 (N_7283,N_911,N_5687);
nand U7284 (N_7284,N_3820,N_4067);
nor U7285 (N_7285,N_4967,N_746);
nor U7286 (N_7286,N_1634,N_1337);
and U7287 (N_7287,N_85,N_3082);
nor U7288 (N_7288,N_1030,N_6085);
nand U7289 (N_7289,N_1325,N_318);
nor U7290 (N_7290,N_191,N_1747);
or U7291 (N_7291,N_2927,N_1962);
and U7292 (N_7292,N_2446,N_1803);
or U7293 (N_7293,N_310,N_2810);
xor U7294 (N_7294,N_1109,N_953);
or U7295 (N_7295,N_2585,N_4823);
and U7296 (N_7296,N_3203,N_5297);
and U7297 (N_7297,N_4402,N_5372);
xor U7298 (N_7298,N_5731,N_1938);
or U7299 (N_7299,N_964,N_5665);
or U7300 (N_7300,N_4752,N_3836);
or U7301 (N_7301,N_5,N_3727);
or U7302 (N_7302,N_6139,N_4899);
xor U7303 (N_7303,N_5637,N_603);
or U7304 (N_7304,N_2544,N_2993);
nand U7305 (N_7305,N_5470,N_2882);
or U7306 (N_7306,N_6164,N_4972);
xor U7307 (N_7307,N_1209,N_3095);
and U7308 (N_7308,N_1756,N_2009);
nand U7309 (N_7309,N_1301,N_4259);
and U7310 (N_7310,N_4421,N_3888);
nor U7311 (N_7311,N_1906,N_2916);
and U7312 (N_7312,N_5033,N_2297);
and U7313 (N_7313,N_326,N_4071);
or U7314 (N_7314,N_3480,N_3123);
nor U7315 (N_7315,N_3026,N_3818);
nand U7316 (N_7316,N_4221,N_4200);
nor U7317 (N_7317,N_3739,N_2669);
nor U7318 (N_7318,N_1373,N_138);
or U7319 (N_7319,N_781,N_2434);
nor U7320 (N_7320,N_1396,N_4753);
and U7321 (N_7321,N_5788,N_1972);
nor U7322 (N_7322,N_1130,N_4928);
or U7323 (N_7323,N_2893,N_6210);
nor U7324 (N_7324,N_1255,N_5310);
nor U7325 (N_7325,N_1913,N_5106);
and U7326 (N_7326,N_5691,N_1441);
and U7327 (N_7327,N_2724,N_48);
or U7328 (N_7328,N_5924,N_2026);
and U7329 (N_7329,N_4289,N_159);
nand U7330 (N_7330,N_5443,N_902);
nor U7331 (N_7331,N_1458,N_1951);
xor U7332 (N_7332,N_5492,N_3853);
nand U7333 (N_7333,N_169,N_6131);
nor U7334 (N_7334,N_2159,N_5040);
nor U7335 (N_7335,N_2398,N_2760);
xnor U7336 (N_7336,N_402,N_3265);
and U7337 (N_7337,N_4850,N_3401);
nand U7338 (N_7338,N_2820,N_2196);
nand U7339 (N_7339,N_5438,N_2738);
or U7340 (N_7340,N_4706,N_5704);
nor U7341 (N_7341,N_1694,N_4294);
nor U7342 (N_7342,N_4719,N_5418);
nor U7343 (N_7343,N_2788,N_918);
nor U7344 (N_7344,N_5519,N_2780);
xnor U7345 (N_7345,N_5416,N_6208);
or U7346 (N_7346,N_5212,N_5013);
and U7347 (N_7347,N_3049,N_5319);
or U7348 (N_7348,N_976,N_2811);
or U7349 (N_7349,N_512,N_5805);
nand U7350 (N_7350,N_2930,N_959);
nand U7351 (N_7351,N_1208,N_3878);
or U7352 (N_7352,N_3990,N_787);
or U7353 (N_7353,N_1190,N_1615);
nor U7354 (N_7354,N_3827,N_4758);
xnor U7355 (N_7355,N_3677,N_2355);
nand U7356 (N_7356,N_236,N_4116);
nand U7357 (N_7357,N_4155,N_4389);
and U7358 (N_7358,N_6088,N_28);
xnor U7359 (N_7359,N_3938,N_2698);
or U7360 (N_7360,N_2497,N_3799);
nand U7361 (N_7361,N_1028,N_4007);
xor U7362 (N_7362,N_5551,N_1338);
and U7363 (N_7363,N_5476,N_3641);
nor U7364 (N_7364,N_3733,N_5007);
nand U7365 (N_7365,N_69,N_657);
or U7366 (N_7366,N_1016,N_3064);
and U7367 (N_7367,N_5407,N_4689);
xnor U7368 (N_7368,N_1306,N_4714);
nor U7369 (N_7369,N_2686,N_1723);
or U7370 (N_7370,N_2382,N_1995);
nor U7371 (N_7371,N_5264,N_1670);
nor U7372 (N_7372,N_4207,N_1317);
and U7373 (N_7373,N_5491,N_1280);
xor U7374 (N_7374,N_6027,N_956);
and U7375 (N_7375,N_3766,N_6033);
nor U7376 (N_7376,N_4243,N_2565);
and U7377 (N_7377,N_4033,N_1795);
nor U7378 (N_7378,N_3634,N_2472);
or U7379 (N_7379,N_2336,N_3883);
nor U7380 (N_7380,N_2696,N_4388);
xor U7381 (N_7381,N_4461,N_1515);
or U7382 (N_7382,N_5395,N_1646);
or U7383 (N_7383,N_3905,N_1439);
or U7384 (N_7384,N_263,N_2664);
nand U7385 (N_7385,N_3610,N_2014);
or U7386 (N_7386,N_1415,N_5269);
or U7387 (N_7387,N_5920,N_2867);
nand U7388 (N_7388,N_3854,N_4172);
nor U7389 (N_7389,N_425,N_238);
nand U7390 (N_7390,N_1169,N_1410);
and U7391 (N_7391,N_987,N_5198);
and U7392 (N_7392,N_5995,N_4238);
xnor U7393 (N_7393,N_1792,N_5656);
nand U7394 (N_7394,N_615,N_960);
xor U7395 (N_7395,N_3580,N_5588);
or U7396 (N_7396,N_5811,N_3293);
or U7397 (N_7397,N_220,N_5182);
and U7398 (N_7398,N_3062,N_3872);
and U7399 (N_7399,N_4105,N_1147);
nand U7400 (N_7400,N_479,N_2116);
and U7401 (N_7401,N_513,N_4330);
or U7402 (N_7402,N_1769,N_1690);
nand U7403 (N_7403,N_4938,N_1550);
nand U7404 (N_7404,N_477,N_2687);
or U7405 (N_7405,N_1119,N_4705);
and U7406 (N_7406,N_5408,N_2883);
or U7407 (N_7407,N_5389,N_6052);
nand U7408 (N_7408,N_2040,N_4216);
nand U7409 (N_7409,N_1080,N_4194);
or U7410 (N_7410,N_4924,N_3759);
and U7411 (N_7411,N_2306,N_1216);
nand U7412 (N_7412,N_5296,N_606);
nand U7413 (N_7413,N_1355,N_5197);
and U7414 (N_7414,N_5532,N_2129);
or U7415 (N_7415,N_3969,N_1240);
nand U7416 (N_7416,N_3067,N_1422);
xor U7417 (N_7417,N_2886,N_2616);
nand U7418 (N_7418,N_4292,N_4956);
or U7419 (N_7419,N_2808,N_3518);
xnor U7420 (N_7420,N_3948,N_3285);
and U7421 (N_7421,N_6125,N_3742);
nor U7422 (N_7422,N_3354,N_314);
nor U7423 (N_7423,N_1656,N_3649);
and U7424 (N_7424,N_5642,N_731);
nand U7425 (N_7425,N_3857,N_1244);
or U7426 (N_7426,N_1955,N_2091);
and U7427 (N_7427,N_488,N_5692);
or U7428 (N_7428,N_1811,N_1247);
or U7429 (N_7429,N_5597,N_295);
and U7430 (N_7430,N_3968,N_5736);
and U7431 (N_7431,N_285,N_3847);
nand U7432 (N_7432,N_3576,N_648);
and U7433 (N_7433,N_5863,N_800);
and U7434 (N_7434,N_5884,N_4433);
and U7435 (N_7435,N_1478,N_2295);
or U7436 (N_7436,N_4325,N_1312);
nand U7437 (N_7437,N_3396,N_1475);
nand U7438 (N_7438,N_4121,N_3331);
nand U7439 (N_7439,N_5313,N_4744);
or U7440 (N_7440,N_4404,N_3861);
and U7441 (N_7441,N_1757,N_1636);
nand U7442 (N_7442,N_1713,N_453);
or U7443 (N_7443,N_2745,N_5671);
nor U7444 (N_7444,N_4037,N_4857);
nand U7445 (N_7445,N_2956,N_2089);
nor U7446 (N_7446,N_4579,N_3046);
nand U7447 (N_7447,N_6184,N_4307);
nand U7448 (N_7448,N_2216,N_1440);
xnor U7449 (N_7449,N_2317,N_131);
nand U7450 (N_7450,N_4263,N_4709);
and U7451 (N_7451,N_1855,N_1559);
xor U7452 (N_7452,N_6011,N_242);
and U7453 (N_7453,N_6091,N_3628);
or U7454 (N_7454,N_863,N_442);
nor U7455 (N_7455,N_3606,N_1833);
and U7456 (N_7456,N_3548,N_334);
xor U7457 (N_7457,N_3721,N_5445);
and U7458 (N_7458,N_5108,N_951);
nand U7459 (N_7459,N_899,N_4034);
xor U7460 (N_7460,N_5991,N_1930);
or U7461 (N_7461,N_2278,N_3209);
nor U7462 (N_7462,N_4049,N_2681);
nor U7463 (N_7463,N_3646,N_5941);
and U7464 (N_7464,N_5563,N_5430);
nand U7465 (N_7465,N_5145,N_294);
nor U7466 (N_7466,N_3940,N_4732);
xnor U7467 (N_7467,N_4074,N_2717);
nand U7468 (N_7468,N_6237,N_1509);
or U7469 (N_7469,N_689,N_5440);
or U7470 (N_7470,N_4266,N_1952);
nand U7471 (N_7471,N_3456,N_4290);
or U7472 (N_7472,N_4395,N_919);
or U7473 (N_7473,N_1168,N_2873);
and U7474 (N_7474,N_5222,N_656);
nand U7475 (N_7475,N_2946,N_1182);
or U7476 (N_7476,N_1963,N_5014);
or U7477 (N_7477,N_541,N_1160);
nand U7478 (N_7478,N_5316,N_2789);
or U7479 (N_7479,N_866,N_1298);
or U7480 (N_7480,N_2432,N_587);
nor U7481 (N_7481,N_1178,N_3921);
nor U7482 (N_7482,N_196,N_4959);
nand U7483 (N_7483,N_1042,N_4561);
or U7484 (N_7484,N_2540,N_5714);
or U7485 (N_7485,N_4622,N_4000);
nand U7486 (N_7486,N_3161,N_1076);
nor U7487 (N_7487,N_730,N_2289);
and U7488 (N_7488,N_3084,N_2851);
or U7489 (N_7489,N_1734,N_925);
or U7490 (N_7490,N_655,N_4725);
and U7491 (N_7491,N_1090,N_2181);
nor U7492 (N_7492,N_4117,N_177);
or U7493 (N_7493,N_2618,N_2978);
nor U7494 (N_7494,N_1115,N_1036);
nor U7495 (N_7495,N_5795,N_2048);
or U7496 (N_7496,N_4419,N_1985);
and U7497 (N_7497,N_2532,N_3694);
nor U7498 (N_7498,N_857,N_572);
or U7499 (N_7499,N_2505,N_2453);
nor U7500 (N_7500,N_3128,N_303);
nor U7501 (N_7501,N_625,N_3685);
or U7502 (N_7502,N_5465,N_5035);
nand U7503 (N_7503,N_5894,N_5129);
and U7504 (N_7504,N_3269,N_4966);
nand U7505 (N_7505,N_1935,N_2399);
nor U7506 (N_7506,N_1752,N_2273);
nor U7507 (N_7507,N_1186,N_4081);
and U7508 (N_7508,N_3635,N_2640);
and U7509 (N_7509,N_5867,N_4454);
nor U7510 (N_7510,N_2232,N_4068);
nor U7511 (N_7511,N_1198,N_6145);
xor U7512 (N_7512,N_3655,N_4687);
and U7513 (N_7513,N_5493,N_5771);
and U7514 (N_7514,N_32,N_4970);
and U7515 (N_7515,N_1293,N_2506);
and U7516 (N_7516,N_2301,N_4908);
and U7517 (N_7517,N_226,N_3690);
xor U7518 (N_7518,N_1726,N_4929);
nor U7519 (N_7519,N_5577,N_3816);
xor U7520 (N_7520,N_1120,N_4278);
nand U7521 (N_7521,N_4685,N_2251);
or U7522 (N_7522,N_922,N_634);
and U7523 (N_7523,N_1187,N_4336);
nor U7524 (N_7524,N_2550,N_480);
nor U7525 (N_7525,N_1675,N_5571);
or U7526 (N_7526,N_5738,N_365);
nor U7527 (N_7527,N_1869,N_2325);
and U7528 (N_7528,N_1767,N_1261);
or U7529 (N_7529,N_3267,N_1448);
or U7530 (N_7530,N_1566,N_742);
nand U7531 (N_7531,N_4741,N_1796);
and U7532 (N_7532,N_5553,N_4250);
and U7533 (N_7533,N_653,N_179);
xnor U7534 (N_7534,N_4224,N_5768);
and U7535 (N_7535,N_5766,N_3228);
xor U7536 (N_7536,N_699,N_130);
xnor U7537 (N_7537,N_4935,N_6182);
nand U7538 (N_7538,N_2899,N_1327);
and U7539 (N_7539,N_1316,N_1049);
and U7540 (N_7540,N_5487,N_5719);
nand U7541 (N_7541,N_1413,N_4900);
xnor U7542 (N_7542,N_9,N_574);
nor U7543 (N_7543,N_5673,N_1842);
nand U7544 (N_7544,N_1289,N_4361);
and U7545 (N_7545,N_4165,N_5617);
nand U7546 (N_7546,N_1157,N_715);
nor U7547 (N_7547,N_966,N_208);
or U7548 (N_7548,N_856,N_3376);
and U7549 (N_7549,N_5708,N_4229);
or U7550 (N_7550,N_3707,N_1435);
nor U7551 (N_7551,N_6101,N_3789);
nand U7552 (N_7552,N_5339,N_5356);
nor U7553 (N_7553,N_3230,N_2123);
nand U7554 (N_7554,N_2797,N_4727);
nand U7555 (N_7555,N_1826,N_4984);
nand U7556 (N_7556,N_5219,N_3717);
xnor U7557 (N_7557,N_6047,N_312);
or U7558 (N_7558,N_338,N_1745);
nand U7559 (N_7559,N_3233,N_1961);
nand U7560 (N_7560,N_192,N_540);
and U7561 (N_7561,N_2416,N_4498);
and U7562 (N_7562,N_2962,N_2773);
or U7563 (N_7563,N_3782,N_1167);
xor U7564 (N_7564,N_5003,N_2304);
nor U7565 (N_7565,N_4087,N_4556);
and U7566 (N_7566,N_1841,N_1217);
nand U7567 (N_7567,N_2262,N_2404);
and U7568 (N_7568,N_5147,N_1349);
and U7569 (N_7569,N_5266,N_3459);
nor U7570 (N_7570,N_5241,N_5050);
and U7571 (N_7571,N_1192,N_4174);
nor U7572 (N_7572,N_1501,N_2620);
nand U7573 (N_7573,N_2369,N_5177);
or U7574 (N_7574,N_3463,N_4445);
nor U7575 (N_7575,N_4577,N_1183);
xnor U7576 (N_7576,N_6057,N_1619);
nand U7577 (N_7577,N_2139,N_627);
xnor U7578 (N_7578,N_2148,N_6175);
xor U7579 (N_7579,N_3542,N_2793);
nor U7580 (N_7580,N_3737,N_5494);
nand U7581 (N_7581,N_1999,N_5926);
nand U7582 (N_7582,N_5265,N_4582);
and U7583 (N_7583,N_152,N_4697);
nor U7584 (N_7584,N_665,N_30);
or U7585 (N_7585,N_1925,N_2722);
nor U7586 (N_7586,N_3227,N_4656);
nand U7587 (N_7587,N_1456,N_3136);
nor U7588 (N_7588,N_357,N_1423);
nand U7589 (N_7589,N_3928,N_449);
and U7590 (N_7590,N_3056,N_4555);
nand U7591 (N_7591,N_875,N_4348);
nor U7592 (N_7592,N_4070,N_4);
nor U7593 (N_7593,N_1062,N_5709);
nor U7594 (N_7594,N_2635,N_2469);
or U7595 (N_7595,N_5127,N_782);
or U7596 (N_7596,N_1133,N_2415);
or U7597 (N_7597,N_2663,N_4360);
or U7598 (N_7598,N_5088,N_5070);
or U7599 (N_7599,N_3772,N_4166);
or U7600 (N_7600,N_4091,N_3009);
and U7601 (N_7601,N_4828,N_2981);
nand U7602 (N_7602,N_3342,N_5950);
or U7603 (N_7603,N_2670,N_4097);
nor U7604 (N_7604,N_1121,N_544);
nor U7605 (N_7605,N_1808,N_4275);
and U7606 (N_7606,N_4619,N_4975);
nor U7607 (N_7607,N_1352,N_975);
xor U7608 (N_7608,N_1395,N_4225);
nand U7609 (N_7609,N_3567,N_6141);
and U7610 (N_7610,N_4632,N_5204);
nor U7611 (N_7611,N_2227,N_3380);
and U7612 (N_7612,N_4755,N_524);
nand U7613 (N_7613,N_2787,N_2783);
or U7614 (N_7614,N_6087,N_1224);
nand U7615 (N_7615,N_5826,N_2588);
nor U7616 (N_7616,N_6023,N_5056);
nor U7617 (N_7617,N_1444,N_3341);
nand U7618 (N_7618,N_1136,N_1530);
nor U7619 (N_7619,N_3134,N_927);
and U7620 (N_7620,N_2281,N_232);
nor U7621 (N_7621,N_1265,N_3316);
or U7622 (N_7622,N_229,N_1994);
nand U7623 (N_7623,N_1620,N_1753);
or U7624 (N_7624,N_3353,N_1116);
nand U7625 (N_7625,N_1918,N_4015);
nor U7626 (N_7626,N_3924,N_4526);
xor U7627 (N_7627,N_1323,N_4236);
or U7628 (N_7628,N_5929,N_5815);
and U7629 (N_7629,N_1604,N_5616);
and U7630 (N_7630,N_1455,N_4405);
xnor U7631 (N_7631,N_2467,N_1069);
or U7632 (N_7632,N_5555,N_643);
nor U7633 (N_7633,N_5437,N_4679);
and U7634 (N_7634,N_754,N_6045);
nor U7635 (N_7635,N_2935,N_636);
xnor U7636 (N_7636,N_4297,N_4248);
nor U7637 (N_7637,N_3933,N_4001);
or U7638 (N_7638,N_738,N_3792);
or U7639 (N_7639,N_4390,N_3238);
xor U7640 (N_7640,N_646,N_1937);
or U7641 (N_7641,N_1043,N_2798);
nand U7642 (N_7642,N_3167,N_5174);
xnor U7643 (N_7643,N_1810,N_3692);
or U7644 (N_7644,N_4653,N_932);
and U7645 (N_7645,N_5575,N_761);
or U7646 (N_7646,N_1471,N_3985);
and U7647 (N_7647,N_4814,N_1447);
nor U7648 (N_7648,N_4476,N_188);
and U7649 (N_7649,N_1346,N_3510);
and U7650 (N_7650,N_1412,N_4494);
or U7651 (N_7651,N_4675,N_2799);
or U7652 (N_7652,N_1302,N_4023);
and U7653 (N_7653,N_3605,N_3981);
or U7654 (N_7654,N_5404,N_6019);
nor U7655 (N_7655,N_4148,N_4530);
nor U7656 (N_7656,N_3377,N_2604);
xnor U7657 (N_7657,N_27,N_4843);
nand U7658 (N_7658,N_2648,N_679);
nand U7659 (N_7659,N_4204,N_3790);
xnor U7660 (N_7660,N_3488,N_5398);
nor U7661 (N_7661,N_1600,N_1035);
and U7662 (N_7662,N_5959,N_2474);
nand U7663 (N_7663,N_46,N_2707);
or U7664 (N_7664,N_2493,N_6040);
and U7665 (N_7665,N_1707,N_2064);
and U7666 (N_7666,N_87,N_5638);
or U7667 (N_7667,N_5886,N_4082);
nor U7668 (N_7668,N_5301,N_1048);
nand U7669 (N_7669,N_3524,N_5814);
nand U7670 (N_7670,N_6016,N_4773);
xor U7671 (N_7671,N_718,N_1701);
and U7672 (N_7672,N_405,N_1950);
and U7673 (N_7673,N_1494,N_1661);
and U7674 (N_7674,N_4946,N_1203);
and U7675 (N_7675,N_3558,N_3824);
nand U7676 (N_7676,N_2740,N_6193);
nand U7677 (N_7677,N_1056,N_84);
nand U7678 (N_7678,N_5621,N_2594);
nor U7679 (N_7679,N_5082,N_5223);
nand U7680 (N_7680,N_182,N_3457);
nor U7681 (N_7681,N_6163,N_415);
and U7682 (N_7682,N_4707,N_2018);
nor U7683 (N_7683,N_1088,N_2032);
nand U7684 (N_7684,N_4440,N_354);
xnor U7685 (N_7685,N_4787,N_2466);
or U7686 (N_7686,N_2939,N_221);
or U7687 (N_7687,N_607,N_1445);
xor U7688 (N_7688,N_6077,N_5935);
nand U7689 (N_7689,N_4713,N_4780);
nor U7690 (N_7690,N_1313,N_4358);
nand U7691 (N_7691,N_1012,N_3725);
nand U7692 (N_7692,N_1739,N_822);
nor U7693 (N_7693,N_4226,N_2385);
nor U7694 (N_7694,N_511,N_1153);
and U7695 (N_7695,N_6226,N_4661);
or U7696 (N_7696,N_4069,N_3709);
or U7697 (N_7697,N_1681,N_5171);
and U7698 (N_7698,N_4613,N_1793);
or U7699 (N_7699,N_5199,N_5985);
nand U7700 (N_7700,N_4359,N_3330);
or U7701 (N_7701,N_3052,N_635);
or U7702 (N_7702,N_4934,N_5431);
and U7703 (N_7703,N_5528,N_1665);
nor U7704 (N_7704,N_745,N_3468);
or U7705 (N_7705,N_1367,N_519);
or U7706 (N_7706,N_5045,N_6004);
nand U7707 (N_7707,N_2425,N_780);
or U7708 (N_7708,N_1696,N_714);
and U7709 (N_7709,N_6188,N_5862);
or U7710 (N_7710,N_4219,N_1657);
or U7711 (N_7711,N_5393,N_5955);
nor U7712 (N_7712,N_6218,N_2950);
nand U7713 (N_7713,N_1871,N_4974);
or U7714 (N_7714,N_5221,N_426);
and U7715 (N_7715,N_577,N_1361);
and U7716 (N_7716,N_5419,N_6109);
nand U7717 (N_7717,N_272,N_1824);
and U7718 (N_7718,N_1840,N_3384);
nor U7719 (N_7719,N_4525,N_2517);
nor U7720 (N_7720,N_1510,N_2101);
xnor U7721 (N_7721,N_1549,N_2329);
or U7722 (N_7722,N_1322,N_2767);
nor U7723 (N_7723,N_2671,N_42);
nand U7724 (N_7724,N_2104,N_3039);
nor U7725 (N_7725,N_5217,N_492);
nor U7726 (N_7726,N_565,N_4193);
nand U7727 (N_7727,N_323,N_5590);
and U7728 (N_7728,N_5084,N_5596);
or U7729 (N_7729,N_1096,N_5988);
nand U7730 (N_7730,N_3311,N_1520);
and U7731 (N_7731,N_3173,N_1052);
nand U7732 (N_7732,N_2574,N_5368);
and U7733 (N_7733,N_1469,N_4416);
and U7734 (N_7734,N_4589,N_2030);
nand U7735 (N_7735,N_4851,N_767);
nor U7736 (N_7736,N_5958,N_766);
and U7737 (N_7737,N_6249,N_4329);
nand U7738 (N_7738,N_4603,N_2400);
nand U7739 (N_7739,N_3719,N_1879);
nor U7740 (N_7740,N_1402,N_5375);
and U7741 (N_7741,N_1708,N_3893);
and U7742 (N_7742,N_305,N_744);
and U7743 (N_7743,N_6064,N_2070);
and U7744 (N_7744,N_2682,N_704);
or U7745 (N_7745,N_5089,N_4520);
and U7746 (N_7746,N_4806,N_5584);
xor U7747 (N_7747,N_3217,N_3918);
xnor U7748 (N_7748,N_3868,N_3848);
nor U7749 (N_7749,N_1341,N_2312);
or U7750 (N_7750,N_1997,N_5974);
nand U7751 (N_7751,N_4621,N_903);
and U7752 (N_7752,N_2326,N_6032);
or U7753 (N_7753,N_4808,N_6113);
nand U7754 (N_7754,N_5114,N_5075);
nor U7755 (N_7755,N_3007,N_4335);
or U7756 (N_7756,N_1214,N_3753);
or U7757 (N_7757,N_1101,N_427);
nor U7758 (N_7758,N_2246,N_1000);
or U7759 (N_7759,N_737,N_4175);
or U7760 (N_7760,N_5495,N_2570);
and U7761 (N_7761,N_5206,N_6176);
nor U7762 (N_7762,N_5786,N_1277);
and U7763 (N_7763,N_4212,N_1942);
nand U7764 (N_7764,N_2922,N_5743);
or U7765 (N_7765,N_5161,N_399);
nor U7766 (N_7766,N_320,N_6126);
nor U7767 (N_7767,N_268,N_5190);
nor U7768 (N_7768,N_2693,N_1274);
nand U7769 (N_7769,N_1304,N_1609);
nand U7770 (N_7770,N_2162,N_1751);
or U7771 (N_7771,N_2063,N_5526);
or U7772 (N_7772,N_64,N_3930);
nor U7773 (N_7773,N_5483,N_5403);
or U7774 (N_7774,N_4575,N_1085);
or U7775 (N_7775,N_3670,N_2877);
and U7776 (N_7776,N_5333,N_4834);
nand U7777 (N_7777,N_4804,N_2066);
xor U7778 (N_7778,N_5349,N_2419);
nand U7779 (N_7779,N_3615,N_537);
nor U7780 (N_7780,N_507,N_4710);
or U7781 (N_7781,N_3417,N_920);
nor U7782 (N_7782,N_1173,N_4847);
nand U7783 (N_7783,N_4424,N_1276);
nor U7784 (N_7784,N_5189,N_4481);
nand U7785 (N_7785,N_5116,N_2536);
and U7786 (N_7786,N_2625,N_3099);
nor U7787 (N_7787,N_328,N_1010);
and U7788 (N_7788,N_1258,N_3065);
nand U7789 (N_7789,N_1436,N_2290);
xor U7790 (N_7790,N_2450,N_4737);
and U7791 (N_7791,N_4678,N_4897);
nor U7792 (N_7792,N_1805,N_1991);
nand U7793 (N_7793,N_2919,N_3496);
and U7794 (N_7794,N_4926,N_4836);
and U7795 (N_7795,N_167,N_4533);
nand U7796 (N_7796,N_3529,N_2484);
nand U7797 (N_7797,N_4139,N_5332);
nand U7798 (N_7798,N_6186,N_3189);
and U7799 (N_7799,N_1398,N_4459);
nand U7800 (N_7800,N_5059,N_1195);
xor U7801 (N_7801,N_5387,N_3470);
nand U7802 (N_7802,N_2642,N_2157);
nor U7803 (N_7803,N_4269,N_1926);
or U7804 (N_7804,N_6189,N_4833);
or U7805 (N_7805,N_424,N_1242);
xnor U7806 (N_7806,N_4018,N_5864);
or U7807 (N_7807,N_3481,N_2241);
nand U7808 (N_7808,N_3562,N_3448);
nor U7809 (N_7809,N_2283,N_4447);
or U7810 (N_7810,N_1154,N_4905);
xor U7811 (N_7811,N_5363,N_2225);
xor U7812 (N_7812,N_4978,N_4818);
xnor U7813 (N_7813,N_322,N_4805);
or U7814 (N_7814,N_4058,N_710);
and U7815 (N_7815,N_2121,N_5284);
nor U7816 (N_7816,N_2138,N_398);
nor U7817 (N_7817,N_2564,N_1588);
nand U7818 (N_7818,N_2358,N_3966);
nor U7819 (N_7819,N_758,N_4765);
nor U7820 (N_7820,N_5851,N_2785);
and U7821 (N_7821,N_49,N_6129);
nand U7822 (N_7822,N_4401,N_458);
and U7823 (N_7823,N_2476,N_5409);
and U7824 (N_7824,N_622,N_4182);
or U7825 (N_7825,N_4141,N_143);
and U7826 (N_7826,N_260,N_475);
nand U7827 (N_7827,N_4774,N_1365);
and U7828 (N_7828,N_5700,N_5489);
nand U7829 (N_7829,N_4962,N_3755);
and U7830 (N_7830,N_2511,N_3392);
or U7831 (N_7831,N_3512,N_5919);
or U7832 (N_7832,N_4432,N_1112);
nand U7833 (N_7833,N_1873,N_1064);
or U7834 (N_7834,N_4163,N_3678);
nand U7835 (N_7835,N_5257,N_3974);
nand U7836 (N_7836,N_4084,N_476);
xnor U7837 (N_7837,N_842,N_3261);
and U7838 (N_7838,N_4154,N_3120);
and U7839 (N_7839,N_6067,N_1533);
nand U7840 (N_7840,N_4723,N_5591);
nand U7841 (N_7841,N_468,N_2311);
and U7842 (N_7842,N_1574,N_1243);
nand U7843 (N_7843,N_778,N_5556);
or U7844 (N_7844,N_397,N_290);
xor U7845 (N_7845,N_2340,N_4667);
nand U7846 (N_7846,N_1948,N_5090);
and U7847 (N_7847,N_3372,N_2395);
or U7848 (N_7848,N_447,N_6243);
or U7849 (N_7849,N_2342,N_3220);
nor U7850 (N_7850,N_193,N_4196);
and U7851 (N_7851,N_2127,N_470);
or U7852 (N_7852,N_1418,N_2859);
and U7853 (N_7853,N_5947,N_619);
nand U7854 (N_7854,N_551,N_231);
nand U7855 (N_7855,N_995,N_5606);
xnor U7856 (N_7856,N_207,N_3728);
nand U7857 (N_7857,N_662,N_3573);
nand U7858 (N_7858,N_6122,N_1146);
nand U7859 (N_7859,N_265,N_158);
nand U7860 (N_7860,N_4537,N_19);
nand U7861 (N_7861,N_5302,N_4570);
and U7862 (N_7862,N_5475,N_5288);
xor U7863 (N_7863,N_5948,N_1519);
nand U7864 (N_7864,N_264,N_3216);
and U7865 (N_7865,N_4300,N_4393);
or U7866 (N_7866,N_5724,N_3164);
nand U7867 (N_7867,N_3156,N_4005);
xor U7868 (N_7868,N_3146,N_2174);
nand U7869 (N_7869,N_4055,N_213);
or U7870 (N_7870,N_5490,N_5235);
nor U7871 (N_7871,N_4451,N_4418);
and U7872 (N_7872,N_1885,N_2428);
xnor U7873 (N_7873,N_94,N_1063);
nor U7874 (N_7874,N_3568,N_5248);
and U7875 (N_7875,N_190,N_6219);
and U7876 (N_7876,N_3520,N_3054);
nor U7877 (N_7877,N_5414,N_829);
nor U7878 (N_7878,N_4186,N_1193);
nor U7879 (N_7879,N_1612,N_3131);
and U7880 (N_7880,N_2959,N_5406);
and U7881 (N_7881,N_1251,N_1321);
nand U7882 (N_7882,N_2843,N_3748);
nand U7883 (N_7883,N_4735,N_3345);
and U7884 (N_7884,N_2323,N_16);
and U7885 (N_7885,N_3625,N_6054);
nand U7886 (N_7886,N_2253,N_1821);
and U7887 (N_7887,N_2858,N_1232);
or U7888 (N_7888,N_1770,N_815);
or U7889 (N_7889,N_1165,N_2756);
nor U7890 (N_7890,N_4016,N_4988);
nor U7891 (N_7891,N_3449,N_5982);
nand U7892 (N_7892,N_13,N_6174);
nand U7893 (N_7893,N_1529,N_1134);
and U7894 (N_7894,N_2000,N_156);
xnor U7895 (N_7895,N_3150,N_942);
nand U7896 (N_7896,N_5818,N_5496);
xor U7897 (N_7897,N_1585,N_5157);
nand U7898 (N_7898,N_3231,N_3282);
nand U7899 (N_7899,N_2046,N_3214);
nand U7900 (N_7900,N_2923,N_543);
nand U7901 (N_7901,N_3876,N_4322);
or U7902 (N_7902,N_5015,N_4239);
xnor U7903 (N_7903,N_3909,N_1568);
nor U7904 (N_7904,N_4986,N_420);
and U7905 (N_7905,N_1724,N_3650);
and U7906 (N_7906,N_5323,N_3665);
nor U7907 (N_7907,N_2163,N_5279);
or U7908 (N_7908,N_1218,N_3111);
nand U7909 (N_7909,N_81,N_4499);
nand U7910 (N_7910,N_4407,N_2461);
nor U7911 (N_7911,N_2890,N_503);
or U7912 (N_7912,N_3279,N_3603);
and U7913 (N_7913,N_1058,N_974);
or U7914 (N_7914,N_2234,N_4356);
and U7915 (N_7915,N_5717,N_5117);
and U7916 (N_7916,N_3745,N_1626);
or U7917 (N_7917,N_3751,N_832);
or U7918 (N_7918,N_3798,N_5504);
nand U7919 (N_7919,N_3773,N_5635);
and U7920 (N_7920,N_1554,N_5278);
and U7921 (N_7921,N_3839,N_2691);
xor U7922 (N_7922,N_2543,N_4223);
or U7923 (N_7923,N_374,N_5674);
or U7924 (N_7924,N_1966,N_2279);
and U7925 (N_7925,N_2309,N_4345);
nor U7926 (N_7926,N_6127,N_3627);
nor U7927 (N_7927,N_4548,N_145);
and U7928 (N_7928,N_4485,N_1086);
or U7929 (N_7929,N_154,N_1235);
nand U7930 (N_7930,N_2733,N_2219);
nand U7931 (N_7931,N_1915,N_3483);
and U7932 (N_7932,N_4855,N_5072);
nand U7933 (N_7933,N_776,N_3565);
nor U7934 (N_7934,N_5130,N_6230);
and U7935 (N_7935,N_1505,N_2854);
and U7936 (N_7936,N_6098,N_3817);
and U7937 (N_7937,N_4312,N_5544);
or U7938 (N_7938,N_1159,N_3337);
or U7939 (N_7939,N_1027,N_4363);
nand U7940 (N_7940,N_5049,N_1490);
nor U7941 (N_7941,N_5953,N_2739);
xor U7942 (N_7942,N_5745,N_2198);
xnor U7943 (N_7943,N_4870,N_6137);
xor U7944 (N_7944,N_735,N_6039);
or U7945 (N_7945,N_6017,N_2602);
or U7946 (N_7946,N_3446,N_5968);
nor U7947 (N_7947,N_4514,N_1114);
nor U7948 (N_7948,N_227,N_330);
and U7949 (N_7949,N_2152,N_275);
nand U7950 (N_7950,N_5073,N_5412);
and U7951 (N_7951,N_202,N_2447);
xnor U7952 (N_7952,N_2146,N_2887);
or U7953 (N_7953,N_3915,N_199);
or U7954 (N_7954,N_6021,N_2175);
and U7955 (N_7955,N_4231,N_3071);
or U7956 (N_7956,N_4012,N_3891);
or U7957 (N_7957,N_6051,N_5794);
or U7958 (N_7958,N_3823,N_5336);
xnor U7959 (N_7959,N_1231,N_4644);
or U7960 (N_7960,N_4466,N_2888);
nand U7961 (N_7961,N_852,N_1689);
or U7962 (N_7962,N_5076,N_1464);
nand U7963 (N_7963,N_2713,N_3077);
xnor U7964 (N_7964,N_2255,N_3406);
and U7965 (N_7965,N_6079,N_3795);
nor U7966 (N_7966,N_2934,N_2823);
nand U7967 (N_7967,N_4943,N_2229);
nand U7968 (N_7968,N_3184,N_5115);
xor U7969 (N_7969,N_4188,N_6097);
nand U7970 (N_7970,N_6211,N_369);
or U7971 (N_7971,N_4191,N_1700);
xor U7972 (N_7972,N_5351,N_593);
nand U7973 (N_7973,N_739,N_4576);
nor U7974 (N_7974,N_4486,N_4785);
and U7975 (N_7975,N_924,N_2573);
and U7976 (N_7976,N_6213,N_5558);
nor U7977 (N_7977,N_2649,N_5646);
xnor U7978 (N_7978,N_4473,N_2031);
xor U7979 (N_7979,N_1784,N_2514);
nand U7980 (N_7980,N_3900,N_1587);
and U7981 (N_7981,N_4032,N_4217);
nand U7982 (N_7982,N_5951,N_3439);
or U7983 (N_7983,N_262,N_1786);
or U7984 (N_7984,N_5239,N_2143);
nor U7985 (N_7985,N_3660,N_2184);
xnor U7986 (N_7986,N_3633,N_5883);
nor U7987 (N_7987,N_2422,N_4283);
or U7988 (N_7988,N_4211,N_462);
nand U7989 (N_7989,N_2459,N_1197);
xnor U7990 (N_7990,N_3840,N_3497);
and U7991 (N_7991,N_3819,N_2131);
nand U7992 (N_7992,N_3210,N_939);
and U7993 (N_7993,N_4215,N_2612);
nor U7994 (N_7994,N_1584,N_2853);
nor U7995 (N_7995,N_4538,N_4417);
nand U7996 (N_7996,N_546,N_2900);
or U7997 (N_7997,N_6170,N_658);
nor U7998 (N_7998,N_400,N_4880);
and U7999 (N_7999,N_516,N_2861);
nor U8000 (N_8000,N_1631,N_4681);
nor U8001 (N_8001,N_1548,N_4022);
or U8002 (N_8002,N_3101,N_1087);
nor U8003 (N_8003,N_2215,N_4208);
or U8004 (N_8004,N_1649,N_728);
and U8005 (N_8005,N_4658,N_5155);
or U8006 (N_8006,N_1839,N_1630);
nand U8007 (N_8007,N_2552,N_1904);
and U8008 (N_8008,N_4671,N_3526);
nand U8009 (N_8009,N_2411,N_2839);
or U8010 (N_8010,N_2563,N_5454);
nor U8011 (N_8011,N_3047,N_5784);
nand U8012 (N_8012,N_2099,N_4738);
nor U8013 (N_8013,N_1022,N_4444);
nand U8014 (N_8014,N_2547,N_3539);
nor U8015 (N_8015,N_3614,N_3593);
or U8016 (N_8016,N_2386,N_1845);
or U8017 (N_8017,N_4961,N_3490);
xnor U8018 (N_8018,N_465,N_2710);
nand U8019 (N_8019,N_553,N_500);
and U8020 (N_8020,N_5469,N_107);
or U8021 (N_8021,N_1213,N_5060);
nor U8022 (N_8022,N_3023,N_1560);
nor U8023 (N_8023,N_549,N_5548);
xnor U8024 (N_8024,N_4316,N_4604);
or U8025 (N_8025,N_111,N_6010);
nor U8026 (N_8026,N_2534,N_741);
nor U8027 (N_8027,N_6024,N_5573);
nor U8028 (N_8028,N_2254,N_2380);
or U8029 (N_8029,N_3240,N_3324);
or U8030 (N_8030,N_2856,N_3765);
and U8031 (N_8031,N_2676,N_5999);
nand U8032 (N_8032,N_5168,N_5983);
and U8033 (N_8033,N_1256,N_3657);
xnor U8034 (N_8034,N_1397,N_1903);
or U8035 (N_8035,N_5973,N_946);
nor U8036 (N_8036,N_5246,N_2880);
nand U8037 (N_8037,N_4178,N_6229);
nor U8038 (N_8038,N_435,N_749);
or U8039 (N_8039,N_864,N_3925);
or U8040 (N_8040,N_1496,N_6059);
nand U8041 (N_8041,N_5914,N_3489);
nand U8042 (N_8042,N_2320,N_609);
xnor U8043 (N_8043,N_2264,N_1066);
or U8044 (N_8044,N_1535,N_86);
and U8045 (N_8045,N_2802,N_3939);
nor U8046 (N_8046,N_786,N_277);
or U8047 (N_8047,N_5909,N_3298);
nor U8048 (N_8048,N_3121,N_4046);
or U8049 (N_8049,N_5989,N_3493);
nand U8050 (N_8050,N_3303,N_2136);
or U8051 (N_8051,N_6228,N_2008);
nand U8052 (N_8052,N_2840,N_5016);
nor U8053 (N_8053,N_2387,N_1400);
xor U8054 (N_8054,N_4887,N_529);
nand U8055 (N_8055,N_6133,N_2057);
nand U8056 (N_8056,N_53,N_5085);
nand U8057 (N_8057,N_253,N_1782);
nand U8058 (N_8058,N_2986,N_562);
and U8059 (N_8059,N_1131,N_4260);
and U8060 (N_8060,N_4013,N_6);
nor U8061 (N_8061,N_5105,N_313);
and U8062 (N_8062,N_1220,N_6005);
and U8063 (N_8063,N_2097,N_5330);
and U8064 (N_8064,N_4305,N_1648);
and U8065 (N_8065,N_1151,N_813);
and U8066 (N_8066,N_3201,N_452);
nor U8067 (N_8067,N_1822,N_4088);
nor U8068 (N_8068,N_3002,N_3070);
nand U8069 (N_8069,N_2489,N_910);
nor U8070 (N_8070,N_4936,N_4531);
nand U8071 (N_8071,N_1653,N_3431);
and U8072 (N_8072,N_2371,N_5881);
nor U8073 (N_8073,N_2834,N_6238);
nand U8074 (N_8074,N_2645,N_1174);
and U8075 (N_8075,N_5585,N_1544);
and U8076 (N_8076,N_600,N_3494);
nand U8077 (N_8077,N_4790,N_1252);
nor U8078 (N_8078,N_1172,N_1561);
nor U8079 (N_8079,N_5651,N_846);
or U8080 (N_8080,N_417,N_5176);
nand U8081 (N_8081,N_3322,N_1571);
or U8082 (N_8082,N_255,N_4441);
nor U8083 (N_8083,N_5095,N_2757);
nor U8084 (N_8084,N_3920,N_5238);
and U8085 (N_8085,N_5801,N_1978);
nor U8086 (N_8086,N_3718,N_752);
xor U8087 (N_8087,N_2313,N_127);
nand U8088 (N_8088,N_2202,N_2440);
nor U8089 (N_8089,N_588,N_2454);
and U8090 (N_8090,N_2990,N_2221);
and U8091 (N_8091,N_4435,N_4731);
nor U8092 (N_8092,N_3333,N_5600);
or U8093 (N_8093,N_412,N_5550);
or U8094 (N_8094,N_4778,N_4750);
nand U8095 (N_8095,N_4896,N_245);
nand U8096 (N_8096,N_3243,N_4201);
or U8097 (N_8097,N_4474,N_4085);
nand U8098 (N_8098,N_6165,N_1591);
or U8099 (N_8099,N_1442,N_5986);
nand U8100 (N_8100,N_5536,N_1799);
nor U8101 (N_8101,N_2475,N_2305);
nand U8102 (N_8102,N_1697,N_3035);
and U8103 (N_8103,N_4406,N_2660);
nor U8104 (N_8104,N_282,N_4324);
or U8105 (N_8105,N_1686,N_317);
nand U8106 (N_8106,N_5855,N_3892);
and U8107 (N_8107,N_1717,N_1959);
nand U8108 (N_8108,N_392,N_847);
or U8109 (N_8109,N_2277,N_5661);
nand U8110 (N_8110,N_3151,N_4491);
xor U8111 (N_8111,N_4098,N_2766);
or U8112 (N_8112,N_3926,N_4490);
nand U8113 (N_8113,N_2084,N_3528);
nor U8114 (N_8114,N_3902,N_1381);
nand U8115 (N_8115,N_2591,N_872);
xnor U8116 (N_8116,N_880,N_4567);
nor U8117 (N_8117,N_3629,N_171);
nor U8118 (N_8118,N_2363,N_3710);
and U8119 (N_8119,N_1709,N_599);
nor U8120 (N_8120,N_6144,N_2836);
nor U8121 (N_8121,N_2558,N_4505);
or U8122 (N_8122,N_4985,N_4830);
nor U8123 (N_8123,N_4138,N_4868);
nand U8124 (N_8124,N_6061,N_1655);
nand U8125 (N_8125,N_4572,N_430);
or U8126 (N_8126,N_2409,N_5200);
nor U8127 (N_8127,N_917,N_1472);
nor U8128 (N_8128,N_721,N_5761);
nor U8129 (N_8129,N_693,N_1859);
or U8130 (N_8130,N_1556,N_6074);
nand U8131 (N_8131,N_3801,N_5512);
nor U8132 (N_8132,N_3175,N_5309);
nor U8133 (N_8133,N_5780,N_2327);
or U8134 (N_8134,N_4545,N_3110);
xor U8135 (N_8135,N_1565,N_3856);
and U8136 (N_8136,N_2703,N_795);
and U8137 (N_8137,N_2180,N_6180);
nand U8138 (N_8138,N_3525,N_6135);
xnor U8139 (N_8139,N_5230,N_673);
and U8140 (N_8140,N_1163,N_1099);
or U8141 (N_8141,N_5520,N_5754);
or U8142 (N_8142,N_3467,N_495);
and U8143 (N_8143,N_4340,N_2592);
and U8144 (N_8144,N_5324,N_5727);
or U8145 (N_8145,N_1434,N_1371);
nor U8146 (N_8146,N_436,N_4660);
and U8147 (N_8147,N_4218,N_1223);
nand U8148 (N_8148,N_701,N_671);
nor U8149 (N_8149,N_611,N_855);
nor U8150 (N_8150,N_4674,N_2926);
xnor U8151 (N_8151,N_1527,N_3996);
nand U8152 (N_8152,N_4387,N_3036);
nand U8153 (N_8153,N_5783,N_884);
nand U8154 (N_8154,N_4383,N_2603);
or U8155 (N_8155,N_2971,N_915);
nor U8156 (N_8156,N_5012,N_2786);
nor U8157 (N_8157,N_2039,N_878);
and U8158 (N_8158,N_840,N_3934);
nor U8159 (N_8159,N_1290,N_3185);
nor U8160 (N_8160,N_4035,N_3398);
nand U8161 (N_8161,N_3306,N_666);
or U8162 (N_8162,N_3814,N_4130);
nand U8163 (N_8163,N_1607,N_3221);
and U8164 (N_8164,N_3256,N_4730);
and U8165 (N_8165,N_630,N_1947);
xnor U8166 (N_8166,N_4131,N_2903);
or U8167 (N_8167,N_1431,N_4565);
nor U8168 (N_8168,N_321,N_3336);
or U8169 (N_8169,N_3266,N_584);
nor U8170 (N_8170,N_1180,N_4770);
and U8171 (N_8171,N_358,N_639);
and U8172 (N_8172,N_3329,N_3159);
and U8173 (N_8173,N_2356,N_237);
nand U8174 (N_8174,N_2516,N_6162);
or U8175 (N_8175,N_3756,N_1760);
nand U8176 (N_8176,N_5291,N_1108);
nor U8177 (N_8177,N_3420,N_3294);
nand U8178 (N_8178,N_2561,N_6124);
and U8179 (N_8179,N_1547,N_1854);
nand U8180 (N_8180,N_3951,N_6146);
and U8181 (N_8181,N_2600,N_3434);
nand U8182 (N_8182,N_394,N_3504);
nand U8183 (N_8183,N_3106,N_5792);
or U8184 (N_8184,N_203,N_4724);
and U8185 (N_8185,N_2353,N_3359);
nand U8186 (N_8186,N_1546,N_4195);
nor U8187 (N_8187,N_2011,N_5032);
nor U8188 (N_8188,N_3254,N_2199);
nor U8189 (N_8189,N_5644,N_6114);
nor U8190 (N_8190,N_952,N_4173);
nor U8191 (N_8191,N_1097,N_176);
nand U8192 (N_8192,N_5428,N_362);
nor U8193 (N_8193,N_3432,N_5498);
nand U8194 (N_8194,N_2751,N_5378);
nand U8195 (N_8195,N_4521,N_5362);
or U8196 (N_8196,N_3919,N_4092);
or U8197 (N_8197,N_6026,N_2661);
nor U8198 (N_8198,N_4354,N_580);
or U8199 (N_8199,N_1731,N_759);
nand U8200 (N_8200,N_1318,N_1524);
nand U8201 (N_8201,N_1262,N_5394);
and U8202 (N_8202,N_1934,N_3264);
nand U8203 (N_8203,N_4600,N_2464);
and U8204 (N_8204,N_2871,N_4028);
nor U8205 (N_8205,N_5898,N_5381);
or U8206 (N_8206,N_4413,N_6071);
xnor U8207 (N_8207,N_3491,N_750);
and U8208 (N_8208,N_1531,N_2829);
and U8209 (N_8209,N_4496,N_4409);
nand U8210 (N_8210,N_2725,N_1200);
nand U8211 (N_8211,N_862,N_1735);
or U8212 (N_8212,N_860,N_1838);
or U8213 (N_8213,N_3212,N_4280);
nand U8214 (N_8214,N_5402,N_2846);
and U8215 (N_8215,N_2812,N_1569);
or U8216 (N_8216,N_827,N_4464);
nor U8217 (N_8217,N_2915,N_4841);
xnor U8218 (N_8218,N_2731,N_5053);
nand U8219 (N_8219,N_5499,N_501);
nand U8220 (N_8220,N_2298,N_2902);
and U8221 (N_8221,N_3058,N_688);
nor U8222 (N_8222,N_2878,N_5122);
or U8223 (N_8223,N_3484,N_1387);
xnor U8224 (N_8224,N_3632,N_5932);
nand U8225 (N_8225,N_4328,N_5413);
nor U8226 (N_8226,N_3277,N_905);
nand U8227 (N_8227,N_2201,N_3364);
nor U8228 (N_8228,N_816,N_302);
nor U8229 (N_8229,N_2677,N_2250);
nor U8230 (N_8230,N_5808,N_4423);
and U8231 (N_8231,N_5353,N_3579);
xnor U8232 (N_8232,N_5523,N_1946);
nor U8233 (N_8233,N_5840,N_687);
or U8234 (N_8234,N_1617,N_1663);
nor U8235 (N_8235,N_3535,N_4488);
or U8236 (N_8236,N_792,N_1405);
xor U8237 (N_8237,N_1968,N_4578);
nor U8238 (N_8238,N_1742,N_1819);
nand U8239 (N_8239,N_5538,N_1315);
or U8240 (N_8240,N_1668,N_4128);
nor U8241 (N_8241,N_4099,N_2364);
nor U8242 (N_8242,N_1977,N_2259);
and U8243 (N_8243,N_1964,N_5138);
and U8244 (N_8244,N_62,N_4762);
nand U8245 (N_8245,N_556,N_155);
nand U8246 (N_8246,N_2176,N_5949);
and U8247 (N_8247,N_3706,N_2113);
nor U8248 (N_8248,N_2062,N_5486);
nor U8249 (N_8249,N_764,N_3869);
nor U8250 (N_8250,N_812,N_775);
and U8251 (N_8251,N_4274,N_2012);
or U8252 (N_8252,N_5925,N_5698);
nor U8253 (N_8253,N_3124,N_4783);
and U8254 (N_8254,N_3433,N_4002);
nor U8255 (N_8255,N_5976,N_5481);
and U8256 (N_8256,N_1067,N_361);
or U8257 (N_8257,N_4883,N_5271);
or U8258 (N_8258,N_467,N_5828);
nand U8259 (N_8259,N_3947,N_3089);
or U8260 (N_8260,N_1715,N_2749);
nor U8261 (N_8261,N_3828,N_3295);
or U8262 (N_8262,N_1774,N_2194);
nand U8263 (N_8263,N_3672,N_5827);
and U8264 (N_8264,N_2744,N_299);
and U8265 (N_8265,N_624,N_3761);
nand U8266 (N_8266,N_5957,N_2242);
nand U8267 (N_8267,N_5937,N_337);
or U8268 (N_8268,N_6038,N_554);
and U8269 (N_8269,N_2056,N_5658);
and U8270 (N_8270,N_1892,N_1622);
or U8271 (N_8271,N_5721,N_4086);
nand U8272 (N_8272,N_3596,N_5092);
nor U8273 (N_8273,N_5838,N_1943);
nand U8274 (N_8274,N_3255,N_5158);
xor U8275 (N_8275,N_4523,N_1379);
nand U8276 (N_8276,N_563,N_3910);
xor U8277 (N_8277,N_128,N_4534);
or U8278 (N_8278,N_6216,N_2347);
or U8279 (N_8279,N_2333,N_2059);
nor U8280 (N_8280,N_3292,N_2284);
nor U8281 (N_8281,N_4150,N_3270);
or U8282 (N_8282,N_4480,N_5913);
nor U8283 (N_8283,N_5643,N_6028);
or U8284 (N_8284,N_3936,N_4076);
nand U8285 (N_8285,N_1425,N_4524);
nand U8286 (N_8286,N_1013,N_4951);
or U8287 (N_8287,N_4640,N_445);
xnor U8288 (N_8288,N_2763,N_3229);
and U8289 (N_8289,N_4109,N_2256);
or U8290 (N_8290,N_4408,N_5615);
and U8291 (N_8291,N_5008,N_4382);
xnor U8292 (N_8292,N_5220,N_3726);
and U8293 (N_8293,N_1358,N_3451);
and U8294 (N_8294,N_4508,N_5253);
or U8295 (N_8295,N_2546,N_5444);
nor U8296 (N_8296,N_2855,N_2576);
nor U8297 (N_8297,N_4994,N_1939);
and U8298 (N_8298,N_3521,N_5559);
nand U8299 (N_8299,N_2523,N_1931);
nor U8300 (N_8300,N_359,N_5568);
and U8301 (N_8301,N_3368,N_5659);
xnor U8302 (N_8302,N_4077,N_4886);
or U8303 (N_8303,N_2049,N_429);
or U8304 (N_8304,N_340,N_2233);
and U8305 (N_8305,N_2228,N_4554);
or U8306 (N_8306,N_2924,N_4688);
nand U8307 (N_8307,N_1579,N_1082);
and U8308 (N_8308,N_2231,N_1862);
and U8309 (N_8309,N_3569,N_2244);
and U8310 (N_8310,N_1145,N_3360);
xor U8311 (N_8311,N_2524,N_329);
or U8312 (N_8312,N_4462,N_6167);
and U8313 (N_8313,N_4349,N_5121);
and U8314 (N_8314,N_2889,N_2362);
nand U8315 (N_8315,N_1264,N_533);
nor U8316 (N_8316,N_5163,N_1369);
xnor U8317 (N_8317,N_2940,N_5525);
nor U8318 (N_8318,N_3219,N_2128);
nor U8319 (N_8319,N_3076,N_4429);
xor U8320 (N_8320,N_5299,N_1933);
nor U8321 (N_8321,N_4858,N_1858);
nand U8322 (N_8322,N_5508,N_2486);
or U8323 (N_8323,N_4206,N_5514);
or U8324 (N_8324,N_3053,N_1476);
nor U8325 (N_8325,N_1590,N_4277);
and U8326 (N_8326,N_669,N_5552);
nor U8327 (N_8327,N_3995,N_708);
and U8328 (N_8328,N_2150,N_4597);
nor U8329 (N_8329,N_5836,N_2559);
nand U8330 (N_8330,N_3325,N_2754);
nor U8331 (N_8331,N_988,N_4366);
nor U8332 (N_8332,N_3517,N_2125);
nand U8333 (N_8333,N_3022,N_2022);
or U8334 (N_8334,N_4230,N_3740);
or U8335 (N_8335,N_3232,N_5119);
nor U8336 (N_8336,N_2366,N_2596);
and U8337 (N_8337,N_3043,N_3890);
nand U8338 (N_8338,N_3722,N_4503);
and U8339 (N_8339,N_2463,N_3943);
nand U8340 (N_8340,N_2837,N_5439);
and U8341 (N_8341,N_1522,N_2958);
xor U8342 (N_8342,N_1019,N_6160);
or U8343 (N_8343,N_3666,N_5737);
or U8344 (N_8344,N_5273,N_5566);
or U8345 (N_8345,N_1364,N_117);
nor U8346 (N_8346,N_1916,N_4799);
or U8347 (N_8347,N_1150,N_1271);
or U8348 (N_8348,N_2998,N_4669);
nand U8349 (N_8349,N_5153,N_5870);
or U8350 (N_8350,N_2495,N_881);
nand U8351 (N_8351,N_4279,N_3013);
xnor U8352 (N_8352,N_2470,N_3394);
nand U8353 (N_8353,N_4981,N_6044);
or U8354 (N_8354,N_1888,N_5148);
or U8355 (N_8355,N_796,N_3262);
and U8356 (N_8356,N_4659,N_4008);
nand U8357 (N_8357,N_4246,N_24);
or U8358 (N_8358,N_4812,N_4788);
nand U8359 (N_8359,N_2952,N_6225);
and U8360 (N_8360,N_1857,N_5799);
or U8361 (N_8361,N_297,N_1990);
nand U8362 (N_8362,N_4690,N_4993);
and U8363 (N_8363,N_3163,N_3544);
nand U8364 (N_8364,N_2556,N_3140);
nand U8365 (N_8365,N_5501,N_5061);
or U8366 (N_8366,N_3399,N_2365);
or U8367 (N_8367,N_5817,N_5969);
nor U8368 (N_8368,N_4063,N_5205);
nand U8369 (N_8369,N_3332,N_6046);
and U8370 (N_8370,N_3172,N_409);
nor U8371 (N_8371,N_2391,N_50);
and U8372 (N_8372,N_2656,N_509);
nand U8373 (N_8373,N_4813,N_353);
nor U8374 (N_8374,N_222,N_189);
nor U8375 (N_8375,N_4314,N_4760);
nand U8376 (N_8376,N_6063,N_4375);
xnor U8377 (N_8377,N_2832,N_5244);
nand U8378 (N_8378,N_1176,N_4122);
nor U8379 (N_8379,N_2445,N_2156);
nand U8380 (N_8380,N_904,N_4680);
or U8381 (N_8381,N_6009,N_421);
nor U8382 (N_8382,N_5905,N_6105);
nor U8383 (N_8383,N_5194,N_1628);
or U8384 (N_8384,N_4302,N_1504);
and U8385 (N_8385,N_1241,N_1093);
and U8386 (N_8386,N_632,N_2617);
or U8387 (N_8387,N_861,N_1927);
nor U8388 (N_8388,N_284,N_4846);
and U8389 (N_8389,N_859,N_1748);
and U8390 (N_8390,N_4949,N_1581);
xor U8391 (N_8391,N_2441,N_5104);
and U8392 (N_8392,N_5227,N_5705);
nor U8393 (N_8393,N_1006,N_3501);
nor U8394 (N_8394,N_5485,N_2300);
nand U8395 (N_8395,N_3912,N_2571);
and U8396 (N_8396,N_3811,N_3415);
nand U8397 (N_8397,N_5800,N_2638);
and U8398 (N_8398,N_5972,N_4066);
and U8399 (N_8399,N_4422,N_3975);
nand U8400 (N_8400,N_777,N_1417);
or U8401 (N_8401,N_2033,N_3291);
nor U8402 (N_8402,N_2271,N_1138);
and U8403 (N_8403,N_2238,N_4529);
or U8404 (N_8404,N_1513,N_5187);
nand U8405 (N_8405,N_4136,N_342);
or U8406 (N_8406,N_821,N_3296);
and U8407 (N_8407,N_2658,N_5734);
and U8408 (N_8408,N_3357,N_3402);
nor U8409 (N_8409,N_2471,N_6093);
nor U8410 (N_8410,N_4594,N_793);
or U8411 (N_8411,N_1847,N_5856);
or U8412 (N_8412,N_983,N_184);
nand U8413 (N_8413,N_2821,N_1500);
or U8414 (N_8414,N_2268,N_3874);
and U8415 (N_8415,N_6112,N_685);
nand U8416 (N_8416,N_3178,N_370);
nor U8417 (N_8417,N_2173,N_5706);
and U8418 (N_8418,N_33,N_1764);
xnor U8419 (N_8419,N_3129,N_3374);
nand U8420 (N_8420,N_5809,N_5831);
or U8421 (N_8421,N_6130,N_6013);
or U8422 (N_8422,N_3541,N_1831);
nor U8423 (N_8423,N_5460,N_1234);
nand U8424 (N_8424,N_1363,N_2970);
nor U8425 (N_8425,N_967,N_4472);
or U8426 (N_8426,N_887,N_217);
nand U8427 (N_8427,N_4436,N_3822);
nor U8428 (N_8428,N_3094,N_1877);
nand U8429 (N_8429,N_4802,N_4006);
nor U8430 (N_8430,N_3055,N_4482);
nor U8431 (N_8431,N_3708,N_2479);
nand U8432 (N_8432,N_5839,N_2538);
nor U8433 (N_8433,N_5048,N_2636);
nand U8434 (N_8434,N_5210,N_498);
nor U8435 (N_8435,N_5964,N_4893);
nor U8436 (N_8436,N_2013,N_4142);
and U8437 (N_8437,N_153,N_4933);
and U8438 (N_8438,N_817,N_2551);
nor U8439 (N_8439,N_3879,N_4869);
and U8440 (N_8440,N_542,N_528);
nor U8441 (N_8441,N_4691,N_716);
xor U8442 (N_8442,N_2957,N_5505);
and U8443 (N_8443,N_2613,N_3323);
or U8444 (N_8444,N_2110,N_5654);
and U8445 (N_8445,N_2007,N_4766);
nor U8446 (N_8446,N_4112,N_5693);
or U8447 (N_8447,N_1059,N_4940);
or U8448 (N_8448,N_5579,N_1727);
nor U8449 (N_8449,N_1682,N_1039);
nor U8450 (N_8450,N_1514,N_5547);
xor U8451 (N_8451,N_1487,N_4726);
nor U8452 (N_8452,N_4161,N_755);
nand U8453 (N_8453,N_4437,N_61);
and U8454 (N_8454,N_929,N_2218);
nand U8455 (N_8455,N_2205,N_4119);
and U8456 (N_8456,N_20,N_5701);
and U8457 (N_8457,N_2674,N_5630);
and U8458 (N_8458,N_434,N_3273);
and U8459 (N_8459,N_4664,N_1034);
nor U8460 (N_8460,N_3247,N_5655);
nand U8461 (N_8461,N_4120,N_1328);
or U8462 (N_8462,N_80,N_3098);
or U8463 (N_8463,N_3365,N_4831);
nor U8464 (N_8464,N_6227,N_637);
nand U8465 (N_8465,N_3300,N_3139);
or U8466 (N_8466,N_3838,N_487);
or U8467 (N_8467,N_717,N_4114);
nor U8468 (N_8468,N_4391,N_6150);
nand U8469 (N_8469,N_6195,N_2734);
and U8470 (N_8470,N_779,N_5679);
and U8471 (N_8471,N_1611,N_11);
or U8472 (N_8472,N_4197,N_5557);
nand U8473 (N_8473,N_2153,N_205);
nand U8474 (N_8474,N_1465,N_3514);
nand U8475 (N_8475,N_4918,N_3005);
and U8476 (N_8476,N_2407,N_2498);
or U8477 (N_8477,N_4769,N_2818);
or U8478 (N_8478,N_2457,N_4341);
xor U8479 (N_8479,N_2879,N_2999);
nand U8480 (N_8480,N_3145,N_2921);
xnor U8481 (N_8481,N_1880,N_3601);
nand U8482 (N_8482,N_301,N_4668);
and U8483 (N_8483,N_4323,N_10);
nand U8484 (N_8484,N_6073,N_37);
xnor U8485 (N_8485,N_539,N_5277);
nor U8486 (N_8486,N_3205,N_5128);
or U8487 (N_8487,N_3165,N_5694);
nand U8488 (N_8488,N_3712,N_3536);
and U8489 (N_8489,N_4610,N_5396);
nand U8490 (N_8490,N_2303,N_4371);
nand U8491 (N_8491,N_5051,N_4140);
nor U8492 (N_8492,N_96,N_2586);
or U8493 (N_8493,N_5960,N_5975);
xor U8494 (N_8494,N_5757,N_1852);
nand U8495 (N_8495,N_4947,N_573);
xor U8496 (N_8496,N_319,N_1901);
or U8497 (N_8497,N_6234,N_3118);
nand U8498 (N_8498,N_4376,N_4134);
and U8499 (N_8499,N_3809,N_5648);
nor U8500 (N_8500,N_1974,N_644);
xor U8501 (N_8501,N_3085,N_440);
nor U8502 (N_8502,N_91,N_2100);
and U8503 (N_8503,N_2577,N_2481);
nand U8504 (N_8504,N_5441,N_1936);
or U8505 (N_8505,N_1493,N_1688);
nand U8506 (N_8506,N_4438,N_4050);
nand U8507 (N_8507,N_2247,N_4854);
nand U8508 (N_8508,N_390,N_2581);
or U8509 (N_8509,N_3093,N_3197);
and U8510 (N_8510,N_5231,N_3697);
nor U8511 (N_8511,N_3807,N_5109);
and U8512 (N_8512,N_1248,N_1051);
or U8513 (N_8513,N_6058,N_4532);
nor U8514 (N_8514,N_1891,N_4829);
and U8515 (N_8515,N_2548,N_3837);
and U8516 (N_8516,N_4781,N_5707);
nor U8517 (N_8517,N_2637,N_808);
and U8518 (N_8518,N_5184,N_1644);
and U8519 (N_8519,N_336,N_1664);
nand U8520 (N_8520,N_1979,N_2973);
and U8521 (N_8521,N_5236,N_1771);
and U8522 (N_8522,N_6151,N_79);
or U8523 (N_8523,N_2914,N_2784);
nor U8524 (N_8524,N_3590,N_3476);
xnor U8525 (N_8525,N_5922,N_1155);
or U8526 (N_8526,N_438,N_4241);
or U8527 (N_8527,N_3462,N_4384);
nand U8528 (N_8528,N_2977,N_2553);
nor U8529 (N_8529,N_6030,N_877);
and U8530 (N_8530,N_4004,N_4321);
and U8531 (N_8531,N_2700,N_1945);
and U8532 (N_8532,N_1065,N_3059);
nand U8533 (N_8533,N_3732,N_3763);
or U8534 (N_8534,N_2813,N_999);
and U8535 (N_8535,N_3288,N_4351);
nand U8536 (N_8536,N_4866,N_678);
nor U8537 (N_8537,N_3653,N_2092);
nand U8538 (N_8538,N_3503,N_3674);
xor U8539 (N_8539,N_4715,N_4568);
and U8540 (N_8540,N_4043,N_2845);
nand U8541 (N_8541,N_457,N_5283);
nor U8542 (N_8542,N_3581,N_4303);
or U8543 (N_8543,N_1291,N_2735);
nor U8544 (N_8544,N_3249,N_1781);
nor U8545 (N_8545,N_1377,N_5303);
and U8546 (N_8546,N_1876,N_1856);
xor U8547 (N_8547,N_1175,N_2692);
or U8548 (N_8548,N_2748,N_5522);
nand U8549 (N_8549,N_5250,N_4288);
or U8550 (N_8550,N_450,N_5854);
xnor U8551 (N_8551,N_2863,N_1468);
and U8552 (N_8552,N_201,N_1029);
nor U8553 (N_8553,N_1404,N_3849);
or U8554 (N_8554,N_930,N_5618);
nand U8555 (N_8555,N_4210,N_3381);
and U8556 (N_8556,N_3075,N_3613);
nand U8557 (N_8557,N_4973,N_3114);
or U8558 (N_8558,N_575,N_680);
and U8559 (N_8559,N_1229,N_1949);
or U8560 (N_8560,N_2050,N_3001);
and U8561 (N_8561,N_5663,N_5473);
nor U8562 (N_8562,N_2736,N_4051);
nand U8563 (N_8563,N_2260,N_836);
nand U8564 (N_8564,N_4244,N_4739);
nor U8565 (N_8565,N_610,N_2274);
or U8566 (N_8566,N_3125,N_125);
xor U8567 (N_8567,N_3373,N_2622);
nor U8568 (N_8568,N_1015,N_2321);
nor U8569 (N_8569,N_3842,N_4040);
nor U8570 (N_8570,N_5294,N_4863);
and U8571 (N_8571,N_5562,N_485);
xnor U8572 (N_8572,N_4093,N_5858);
and U8573 (N_8573,N_3585,N_2501);
nand U8574 (N_8574,N_3498,N_4410);
or U8575 (N_8575,N_4931,N_5765);
or U8576 (N_8576,N_2053,N_446);
nor U8577 (N_8577,N_493,N_2187);
nor U8578 (N_8578,N_3696,N_4222);
nand U8579 (N_8579,N_2028,N_4213);
nand U8580 (N_8580,N_4083,N_6031);
nor U8581 (N_8581,N_22,N_1215);
nand U8582 (N_8582,N_350,N_2688);
or U8583 (N_8583,N_5272,N_941);
nand U8584 (N_8584,N_5542,N_1332);
or U8585 (N_8585,N_5126,N_700);
or U8586 (N_8586,N_3806,N_2742);
xor U8587 (N_8587,N_4510,N_437);
and U8588 (N_8588,N_1512,N_4825);
or U8589 (N_8589,N_1645,N_3835);
nand U8590 (N_8590,N_518,N_105);
and U8591 (N_8591,N_2435,N_3068);
nor U8592 (N_8592,N_3317,N_5091);
nand U8593 (N_8593,N_214,N_3443);
nand U8594 (N_8594,N_1286,N_2189);
nand U8595 (N_8595,N_4877,N_2549);
nand U8596 (N_8596,N_363,N_1555);
and U8597 (N_8597,N_1651,N_5232);
nand U8598 (N_8598,N_2016,N_5341);
and U8599 (N_8599,N_373,N_5259);
or U8600 (N_8600,N_2841,N_3714);
nand U8601 (N_8601,N_4574,N_4101);
or U8602 (N_8602,N_2266,N_1736);
and U8603 (N_8603,N_4599,N_2069);
nor U8604 (N_8604,N_550,N_368);
nor U8605 (N_8605,N_5369,N_849);
xnor U8606 (N_8606,N_3683,N_5782);
xnor U8607 (N_8607,N_3069,N_1577);
nor U8608 (N_8608,N_1339,N_604);
and U8609 (N_8609,N_3994,N_4913);
or U8610 (N_8610,N_5364,N_325);
or U8611 (N_8611,N_3999,N_3412);
or U8612 (N_8612,N_3624,N_3607);
xor U8613 (N_8613,N_4162,N_6132);
nor U8614 (N_8614,N_4775,N_2679);
or U8615 (N_8615,N_2443,N_4054);
or U8616 (N_8616,N_2455,N_3970);
nand U8617 (N_8617,N_3622,N_2897);
nand U8618 (N_8618,N_2876,N_2901);
or U8619 (N_8619,N_195,N_901);
and U8620 (N_8620,N_3654,N_1558);
nor U8621 (N_8621,N_2770,N_5608);
xnor U8622 (N_8622,N_1987,N_3015);
nand U8623 (N_8623,N_6083,N_4452);
and U8624 (N_8624,N_3896,N_1428);
and U8625 (N_8625,N_4720,N_3224);
nor U8626 (N_8626,N_6200,N_2657);
and U8627 (N_8627,N_1894,N_3138);
nand U8628 (N_8628,N_1861,N_2554);
nor U8629 (N_8629,N_3202,N_2235);
nor U8630 (N_8630,N_3107,N_2537);
or U8631 (N_8631,N_1005,N_5195);
nor U8632 (N_8632,N_3959,N_3117);
nor U8633 (N_8633,N_3850,N_3366);
nor U8634 (N_8634,N_454,N_5134);
nor U8635 (N_8635,N_2759,N_3858);
and U8636 (N_8636,N_4026,N_4791);
or U8637 (N_8637,N_4264,N_522);
and U8638 (N_8638,N_2895,N_481);
or U8639 (N_8639,N_5484,N_1091);
nor U8640 (N_8640,N_618,N_2819);
or U8641 (N_8641,N_4443,N_3851);
and U8642 (N_8642,N_1384,N_5938);
xor U8643 (N_8643,N_954,N_3020);
and U8644 (N_8644,N_1351,N_1411);
nand U8645 (N_8645,N_3340,N_1650);
nand U8646 (N_8646,N_3477,N_187);
or U8647 (N_8647,N_4756,N_4989);
nor U8648 (N_8648,N_3626,N_2906);
xor U8649 (N_8649,N_4583,N_3686);
or U8650 (N_8650,N_2982,N_5384);
xor U8651 (N_8651,N_147,N_279);
and U8652 (N_8652,N_3941,N_3016);
or U8653 (N_8653,N_2058,N_246);
nand U8654 (N_8654,N_5164,N_5667);
nand U8655 (N_8655,N_3066,N_1526);
or U8656 (N_8656,N_2593,N_2195);
nor U8657 (N_8657,N_3584,N_4965);
nand U8658 (N_8658,N_2694,N_3465);
nand U8659 (N_8659,N_5682,N_2086);
or U8660 (N_8660,N_2149,N_5464);
and U8661 (N_8661,N_3019,N_3444);
or U8662 (N_8662,N_3667,N_2911);
nor U8663 (N_8663,N_4282,N_1846);
and U8664 (N_8664,N_2343,N_251);
nor U8665 (N_8665,N_908,N_641);
nand U8666 (N_8666,N_1741,N_1100);
or U8667 (N_8667,N_1319,N_505);
nor U8668 (N_8668,N_697,N_5425);
and U8669 (N_8669,N_5895,N_4920);
nand U8670 (N_8670,N_6117,N_1161);
and U8671 (N_8671,N_4517,N_1761);
nor U8672 (N_8672,N_4100,N_2294);
nand U8673 (N_8673,N_99,N_5038);
and U8674 (N_8674,N_5041,N_126);
nor U8675 (N_8675,N_2792,N_4932);
and U8676 (N_8676,N_3720,N_1835);
nand U8677 (N_8677,N_6065,N_1762);
nand U8678 (N_8678,N_5226,N_3953);
nor U8679 (N_8679,N_2397,N_4199);
or U8680 (N_8680,N_3595,N_4591);
nand U8681 (N_8681,N_4891,N_4412);
or U8682 (N_8682,N_12,N_2492);
and U8683 (N_8683,N_1814,N_2954);
or U8684 (N_8684,N_3979,N_3081);
or U8685 (N_8685,N_2697,N_5252);
nand U8686 (N_8686,N_4844,N_4242);
or U8687 (N_8687,N_4475,N_5755);
nor U8688 (N_8688,N_5026,N_2119);
nand U8689 (N_8689,N_5203,N_1463);
or U8690 (N_8690,N_3087,N_5371);
or U8691 (N_8691,N_5790,N_3474);
xor U8692 (N_8692,N_3762,N_3549);
or U8693 (N_8693,N_3461,N_1698);
xnor U8694 (N_8694,N_5380,N_2609);
and U8695 (N_8695,N_4313,N_694);
nor U8696 (N_8696,N_5703,N_5785);
and U8697 (N_8697,N_1800,N_5120);
and U8698 (N_8698,N_3897,N_670);
xor U8699 (N_8699,N_4160,N_283);
nand U8700 (N_8700,N_1113,N_709);
or U8701 (N_8701,N_1758,N_3177);
nand U8702 (N_8702,N_2892,N_1185);
nand U8703 (N_8703,N_2984,N_3429);
xnor U8704 (N_8704,N_2969,N_5509);
nand U8705 (N_8705,N_4884,N_346);
nor U8706 (N_8706,N_428,N_1836);
nor U8707 (N_8707,N_4044,N_1348);
nand U8708 (N_8708,N_5280,N_5564);
nand U8709 (N_8709,N_5102,N_6020);
nor U8710 (N_8710,N_3923,N_2047);
nand U8711 (N_8711,N_1586,N_6075);
nor U8712 (N_8712,N_1408,N_1257);
nand U8713 (N_8713,N_3500,N_6172);
and U8714 (N_8714,N_2061,N_1443);
or U8715 (N_8715,N_971,N_1783);
xor U8716 (N_8716,N_396,N_897);
nand U8717 (N_8717,N_3283,N_5447);
xnor U8718 (N_8718,N_2144,N_760);
nand U8719 (N_8719,N_3097,N_5850);
nand U8720 (N_8720,N_3057,N_2980);
nand U8721 (N_8721,N_762,N_997);
and U8722 (N_8722,N_113,N_2288);
nand U8723 (N_8723,N_3907,N_5759);
xnor U8724 (N_8724,N_4347,N_1608);
or U8725 (N_8725,N_6204,N_3351);
nor U8726 (N_8726,N_5531,N_1202);
or U8727 (N_8727,N_1744,N_83);
or U8728 (N_8728,N_3684,N_4991);
nor U8729 (N_8729,N_4041,N_5952);
and U8730 (N_8730,N_5751,N_5459);
or U8731 (N_8731,N_2599,N_1881);
or U8732 (N_8732,N_5599,N_6220);
or U8733 (N_8733,N_6072,N_6153);
nor U8734 (N_8734,N_3318,N_858);
or U8735 (N_8735,N_4543,N_1040);
nor U8736 (N_8736,N_4718,N_4080);
and U8737 (N_8737,N_2051,N_3363);
and U8738 (N_8738,N_4110,N_4515);
or U8739 (N_8739,N_55,N_4434);
or U8740 (N_8740,N_4977,N_998);
xnor U8741 (N_8741,N_5605,N_3997);
xor U8742 (N_8742,N_2995,N_2217);
nor U8743 (N_8743,N_5592,N_474);
nor U8744 (N_8744,N_3045,N_6053);
and U8745 (N_8745,N_3414,N_814);
and U8746 (N_8746,N_980,N_5005);
nor U8747 (N_8747,N_5074,N_1127);
and U8748 (N_8748,N_5166,N_2105);
or U8749 (N_8749,N_667,N_4952);
or U8750 (N_8750,N_1883,N_824);
nand U8751 (N_8751,N_3102,N_1228);
or U8752 (N_8752,N_3656,N_5146);
nand U8753 (N_8753,N_4842,N_965);
nor U8754 (N_8754,N_2608,N_2078);
xnor U8755 (N_8755,N_947,N_5343);
nand U8756 (N_8756,N_943,N_2597);
and U8757 (N_8757,N_2160,N_200);
or U8758 (N_8758,N_2868,N_5131);
or U8759 (N_8759,N_1671,N_273);
nor U8760 (N_8760,N_3174,N_1878);
and U8761 (N_8761,N_5570,N_4745);
nor U8762 (N_8762,N_2379,N_6000);
nor U8763 (N_8763,N_491,N_3734);
and U8764 (N_8764,N_809,N_5604);
and U8765 (N_8765,N_2865,N_2908);
xnor U8766 (N_8766,N_3142,N_423);
nand U8767 (N_8767,N_2348,N_530);
nand U8768 (N_8768,N_2429,N_682);
nor U8769 (N_8769,N_5335,N_4251);
or U8770 (N_8770,N_4716,N_3771);
or U8771 (N_8771,N_4901,N_5868);
nand U8772 (N_8772,N_621,N_1863);
xnor U8773 (N_8773,N_614,N_4536);
xnor U8774 (N_8774,N_2976,N_4252);
or U8775 (N_8775,N_2791,N_43);
xor U8776 (N_8776,N_4633,N_1430);
or U8777 (N_8777,N_2905,N_5561);
nand U8778 (N_8778,N_3932,N_459);
and U8779 (N_8779,N_4442,N_5834);
nand U8780 (N_8780,N_3698,N_5427);
or U8781 (N_8781,N_1362,N_3271);
xor U8782 (N_8782,N_5322,N_4677);
and U8783 (N_8783,N_5689,N_2293);
nor U8784 (N_8784,N_2265,N_3335);
and U8785 (N_8785,N_5311,N_5482);
and U8786 (N_8786,N_6106,N_204);
or U8787 (N_8787,N_2405,N_5934);
and U8788 (N_8788,N_5191,N_3587);
and U8789 (N_8789,N_647,N_4922);
and U8790 (N_8790,N_4665,N_4124);
or U8791 (N_8791,N_77,N_2394);
nand U8792 (N_8792,N_5791,N_5609);
nor U8793 (N_8793,N_3309,N_2702);
xnor U8794 (N_8794,N_3730,N_472);
or U8795 (N_8795,N_1718,N_1054);
nand U8796 (N_8796,N_3880,N_4513);
xor U8797 (N_8797,N_4786,N_1164);
or U8798 (N_8798,N_1662,N_5729);
and U8799 (N_8799,N_1077,N_65);
nor U8800 (N_8800,N_1729,N_2580);
or U8801 (N_8801,N_5096,N_5882);
nand U8802 (N_8802,N_3421,N_2684);
or U8803 (N_8803,N_4903,N_3958);
and U8804 (N_8804,N_1798,N_2010);
and U8805 (N_8805,N_3758,N_4463);
nor U8806 (N_8806,N_1914,N_2800);
nor U8807 (N_8807,N_3411,N_743);
or U8808 (N_8808,N_3875,N_3545);
xor U8809 (N_8809,N_2796,N_4171);
nor U8810 (N_8810,N_5018,N_2178);
nor U8811 (N_8811,N_3699,N_5448);
nor U8812 (N_8812,N_3752,N_4453);
and U8813 (N_8813,N_839,N_2088);
nand U8814 (N_8814,N_5142,N_1954);
nor U8815 (N_8815,N_3509,N_3588);
or U8816 (N_8816,N_2824,N_150);
and U8817 (N_8817,N_6191,N_698);
and U8818 (N_8818,N_3304,N_4233);
or U8819 (N_8819,N_1502,N_6055);
nand U8820 (N_8820,N_347,N_895);
nand U8821 (N_8821,N_1592,N_1706);
and U8822 (N_8822,N_2508,N_1221);
nand U8823 (N_8823,N_2291,N_1158);
or U8824 (N_8824,N_5385,N_1539);
or U8825 (N_8825,N_5011,N_1641);
xnor U8826 (N_8826,N_5254,N_3669);
and U8827 (N_8827,N_5057,N_4029);
and U8828 (N_8828,N_4742,N_5601);
or U8829 (N_8829,N_162,N_3369);
and U8830 (N_8830,N_1451,N_844);
xor U8831 (N_8831,N_1919,N_5810);
or U8832 (N_8832,N_711,N_1986);
nand U8833 (N_8833,N_5037,N_3944);
nor U8834 (N_8834,N_2420,N_4902);
or U8835 (N_8835,N_990,N_175);
and U8836 (N_8836,N_1333,N_3911);
or U8837 (N_8837,N_1484,N_1045);
or U8838 (N_8838,N_3639,N_570);
or U8839 (N_8839,N_23,N_6236);
or U8840 (N_8840,N_1061,N_4950);
nand U8841 (N_8841,N_5690,N_1605);
nor U8842 (N_8842,N_3042,N_4832);
nand U8843 (N_8843,N_4636,N_1497);
nor U8844 (N_8844,N_3689,N_2480);
nor U8845 (N_8845,N_4145,N_3440);
nor U8846 (N_8846,N_940,N_5192);
nand U8847 (N_8847,N_5214,N_4996);
and U8848 (N_8848,N_969,N_2764);
nand U8849 (N_8849,N_6084,N_6201);
or U8850 (N_8850,N_640,N_3895);
nand U8851 (N_8851,N_4385,N_2920);
or U8852 (N_8852,N_890,N_1275);
nand U8853 (N_8853,N_4227,N_433);
or U8854 (N_8854,N_3356,N_4815);
or U8855 (N_8855,N_2816,N_4333);
and U8856 (N_8856,N_2239,N_4646);
nand U8857 (N_8857,N_331,N_4587);
nand U8858 (N_8858,N_5463,N_1354);
nand U8859 (N_8859,N_3630,N_3788);
nand U8860 (N_8860,N_1802,N_3404);
or U8861 (N_8861,N_3208,N_6152);
and U8862 (N_8862,N_2052,N_5358);
and U8863 (N_8863,N_5453,N_4183);
nor U8864 (N_8864,N_1053,N_3547);
or U8865 (N_8865,N_1421,N_5971);
nand U8866 (N_8866,N_5962,N_1896);
nor U8867 (N_8867,N_1399,N_3651);
and U8868 (N_8868,N_2578,N_6240);
xor U8869 (N_8869,N_3437,N_3516);
nor U8870 (N_8870,N_1481,N_590);
or U8871 (N_8871,N_2848,N_957);
xor U8872 (N_8872,N_132,N_1797);
nor U8873 (N_8873,N_5843,N_4273);
and U8874 (N_8874,N_2704,N_5488);
and U8875 (N_8875,N_3986,N_5787);
nand U8876 (N_8876,N_2662,N_6245);
nor U8877 (N_8877,N_121,N_4761);
xor U8878 (N_8878,N_4772,N_4268);
xor U8879 (N_8879,N_5915,N_1572);
nor U8880 (N_8880,N_6115,N_4907);
or U8881 (N_8881,N_996,N_3464);
nand U8882 (N_8882,N_5685,N_2937);
nand U8883 (N_8883,N_67,N_1237);
or U8884 (N_8884,N_5789,N_2330);
nor U8885 (N_8885,N_1273,N_772);
or U8886 (N_8886,N_535,N_5634);
nand U8887 (N_8887,N_2830,N_3702);
or U8888 (N_8888,N_867,N_5410);
and U8889 (N_8889,N_3387,N_4180);
or U8890 (N_8890,N_2771,N_2345);
and U8891 (N_8891,N_3513,N_4353);
or U8892 (N_8892,N_4598,N_5888);
and U8893 (N_8893,N_2077,N_293);
and U8894 (N_8894,N_1303,N_1281);
and U8895 (N_8895,N_3715,N_5763);
xor U8896 (N_8896,N_2073,N_3991);
or U8897 (N_8897,N_5467,N_4146);
nor U8898 (N_8898,N_5859,N_652);
xor U8899 (N_8899,N_1828,N_5921);
and U8900 (N_8900,N_1450,N_2346);
nor U8901 (N_8901,N_1969,N_1692);
or U8902 (N_8902,N_1270,N_5819);
or U8903 (N_8903,N_740,N_2171);
nand U8904 (N_8904,N_4331,N_3515);
nand U8905 (N_8905,N_17,N_6049);
nand U8906 (N_8906,N_870,N_4240);
nand U8907 (N_8907,N_5574,N_5456);
nand U8908 (N_8908,N_3258,N_1759);
or U8909 (N_8909,N_3349,N_973);
nand U8910 (N_8910,N_5017,N_311);
and U8911 (N_8911,N_160,N_5631);
or U8912 (N_8912,N_307,N_339);
nand U8913 (N_8913,N_4584,N_6223);
nand U8914 (N_8914,N_2996,N_1459);
and U8915 (N_8915,N_256,N_3027);
xor U8916 (N_8916,N_2864,N_4202);
nand U8917 (N_8917,N_5797,N_6185);
xor U8918 (N_8918,N_3410,N_3957);
and U8919 (N_8919,N_2414,N_921);
or U8920 (N_8920,N_6002,N_2389);
and U8921 (N_8921,N_1126,N_3779);
nor U8922 (N_8922,N_823,N_6092);
xor U8923 (N_8923,N_269,N_6241);
nor U8924 (N_8924,N_2750,N_4552);
nand U8925 (N_8925,N_2372,N_186);
nor U8926 (N_8926,N_5619,N_6103);
nor U8927 (N_8927,N_5320,N_3908);
and U8928 (N_8928,N_3445,N_3436);
or U8929 (N_8929,N_3253,N_3942);
and U8930 (N_8930,N_3998,N_5946);
nor U8931 (N_8931,N_5778,N_1037);
nor U8932 (N_8932,N_2421,N_2743);
and U8933 (N_8933,N_3297,N_298);
nor U8934 (N_8934,N_6036,N_2601);
xnor U8935 (N_8935,N_296,N_315);
nor U8936 (N_8936,N_3193,N_5159);
or U8937 (N_8937,N_4090,N_2983);
or U8938 (N_8938,N_4792,N_1953);
and U8939 (N_8939,N_1970,N_5331);
or U8940 (N_8940,N_4964,N_4917);
nor U8941 (N_8941,N_3583,N_5987);
or U8942 (N_8942,N_5270,N_60);
nor U8943 (N_8943,N_5063,N_1813);
nor U8944 (N_8944,N_1201,N_118);
or U8945 (N_8945,N_3395,N_3289);
nor U8946 (N_8946,N_1887,N_5111);
nand U8947 (N_8947,N_4953,N_819);
and U8948 (N_8948,N_403,N_3326);
nor U8949 (N_8949,N_1457,N_5350);
nand U8950 (N_8950,N_1386,N_4295);
nand U8951 (N_8951,N_5896,N_3965);
and U8952 (N_8952,N_288,N_5998);
nand U8953 (N_8953,N_4541,N_1314);
nor U8954 (N_8954,N_3899,N_3144);
nand U8955 (N_8955,N_2518,N_2726);
nor U8956 (N_8956,N_3152,N_5781);
nor U8957 (N_8957,N_5039,N_1768);
and U8958 (N_8958,N_5918,N_2203);
xnor U8959 (N_8959,N_6006,N_3729);
or U8960 (N_8960,N_401,N_4626);
or U8961 (N_8961,N_5046,N_3204);
and U8962 (N_8962,N_5906,N_5094);
xnor U8963 (N_8963,N_1335,N_2491);
xor U8964 (N_8964,N_1031,N_4332);
or U8965 (N_8965,N_414,N_2267);
nor U8966 (N_8966,N_2891,N_4009);
xnor U8967 (N_8967,N_3886,N_5141);
or U8968 (N_8968,N_1720,N_224);
and U8969 (N_8969,N_5213,N_1614);
nor U8970 (N_8970,N_3972,N_835);
nor U8971 (N_8971,N_1973,N_4803);
nor U8972 (N_8972,N_3898,N_1868);
nor U8973 (N_8973,N_1079,N_2541);
nand U8974 (N_8974,N_2606,N_2377);
and U8975 (N_8975,N_1089,N_3843);
or U8976 (N_8976,N_4518,N_1470);
or U8977 (N_8977,N_4159,N_1552);
and U8978 (N_8978,N_5822,N_5300);
or U8979 (N_8979,N_6003,N_3393);
xnor U8980 (N_8980,N_2782,N_3648);
nor U8981 (N_8981,N_1152,N_1356);
xor U8982 (N_8982,N_6099,N_2826);
and U8983 (N_8983,N_5242,N_4819);
or U8984 (N_8984,N_3074,N_3422);
and U8985 (N_8985,N_6244,N_2705);
or U8986 (N_8986,N_4652,N_751);
and U8987 (N_8987,N_5716,N_8);
nand U8988 (N_8988,N_4428,N_885);
and U8989 (N_8989,N_5169,N_2142);
nor U8990 (N_8990,N_2151,N_5023);
nor U8991 (N_8991,N_4682,N_281);
xnor U8992 (N_8992,N_4465,N_1038);
and U8993 (N_8993,N_732,N_1576);
nand U8994 (N_8994,N_3537,N_4027);
nor U8995 (N_8995,N_1507,N_534);
nand U8996 (N_8996,N_93,N_110);
and U8997 (N_8997,N_2027,N_948);
nor U8998 (N_8998,N_2126,N_4798);
or U8999 (N_8999,N_5893,N_2473);
and U9000 (N_9000,N_4153,N_690);
or U9001 (N_9001,N_598,N_5963);
or U9002 (N_9002,N_3361,N_2762);
nand U9003 (N_9003,N_3302,N_6050);
nand U9004 (N_9004,N_1642,N_6155);
and U9005 (N_9005,N_5513,N_5468);
nand U9006 (N_9006,N_6095,N_4133);
and U9007 (N_9007,N_4743,N_5042);
and U9008 (N_9008,N_2402,N_4365);
nand U9009 (N_9009,N_5188,N_2381);
nand U9010 (N_9010,N_4487,N_5902);
and U9011 (N_9011,N_4800,N_356);
and U9012 (N_9012,N_3791,N_4835);
nand U9013 (N_9013,N_820,N_1667);
nand U9014 (N_9014,N_3130,N_4457);
xor U9015 (N_9015,N_2641,N_1971);
nor U9016 (N_9016,N_2987,N_2907);
nor U9017 (N_9017,N_1297,N_4563);
or U9018 (N_9018,N_5749,N_2338);
nand U9019 (N_9019,N_1124,N_1219);
or U9020 (N_9020,N_4509,N_3877);
nor U9021 (N_9021,N_3370,N_1267);
nand U9022 (N_9022,N_5911,N_5967);
or U9023 (N_9023,N_5366,N_2190);
and U9024 (N_9024,N_1336,N_3797);
nand U9025 (N_9025,N_2210,N_797);
nand U9026 (N_9026,N_4430,N_557);
nor U9027 (N_9027,N_5516,N_5992);
or U9028 (N_9028,N_372,N_944);
xnor U9029 (N_9029,N_3079,N_807);
and U9030 (N_9030,N_1703,N_3551);
nand U9031 (N_9031,N_1454,N_2029);
nand U9032 (N_9032,N_1511,N_261);
nand U9033 (N_9033,N_558,N_1370);
nand U9034 (N_9034,N_3400,N_1740);
xor U9035 (N_9035,N_5124,N_4298);
or U9036 (N_9036,N_4507,N_5939);
and U9037 (N_9037,N_3435,N_2512);
nor U9038 (N_9038,N_4253,N_1368);
xor U9039 (N_9039,N_4394,N_2992);
nand U9040 (N_9040,N_504,N_5660);
nor U9041 (N_9041,N_4187,N_1353);
and U9042 (N_9042,N_266,N_5081);
nor U9043 (N_9043,N_791,N_5582);
nor U9044 (N_9044,N_4308,N_1142);
and U9045 (N_9045,N_5426,N_4506);
or U9046 (N_9046,N_3808,N_5382);
xor U9047 (N_9047,N_702,N_2526);
nor U9048 (N_9048,N_3741,N_4373);
and U9049 (N_9049,N_3492,N_2567);
nor U9050 (N_9050,N_1094,N_4717);
nand U9051 (N_9051,N_2223,N_2439);
or U9052 (N_9052,N_1419,N_4573);
nor U9053 (N_9053,N_6090,N_3011);
and U9054 (N_9054,N_3640,N_1975);
and U9055 (N_9055,N_5308,N_461);
or U9056 (N_9056,N_3620,N_719);
nor U9057 (N_9057,N_5889,N_4676);
nand U9058 (N_9058,N_3804,N_6086);
and U9059 (N_9059,N_1525,N_2172);
and U9060 (N_9060,N_4364,N_56);
xor U9061 (N_9061,N_5680,N_2769);
nand U9062 (N_9062,N_5885,N_1812);
or U9063 (N_9063,N_5793,N_3643);
and U9064 (N_9064,N_5567,N_5640);
nor U9065 (N_9065,N_2884,N_4784);
nor U9066 (N_9066,N_5928,N_4824);
and U9067 (N_9067,N_1210,N_2212);
xnor U9068 (N_9068,N_4137,N_108);
and U9069 (N_9069,N_695,N_404);
nand U9070 (N_9070,N_1929,N_1632);
xnor U9071 (N_9071,N_4670,N_3424);
nor U9072 (N_9072,N_234,N_6192);
nor U9073 (N_9073,N_1775,N_2155);
or U9074 (N_9074,N_463,N_5823);
and U9075 (N_9075,N_327,N_3143);
and U9076 (N_9076,N_4645,N_3327);
or U9077 (N_9077,N_5534,N_5125);
nor U9078 (N_9078,N_460,N_73);
nand U9079 (N_9079,N_1593,N_2410);
xnor U9080 (N_9080,N_4386,N_3673);
xor U9081 (N_9081,N_381,N_3617);
xor U9082 (N_9082,N_2431,N_1716);
nor U9083 (N_9083,N_4593,N_3237);
nor U9084 (N_9084,N_4650,N_517);
nor U9085 (N_9085,N_4102,N_1144);
or U9086 (N_9086,N_1684,N_133);
nor U9087 (N_9087,N_2071,N_2894);
or U9088 (N_9088,N_3413,N_2720);
nor U9089 (N_9089,N_3499,N_2401);
nor U9090 (N_9090,N_1557,N_2632);
nand U9091 (N_9091,N_3794,N_3348);
nor U9092 (N_9092,N_1308,N_241);
and U9093 (N_9093,N_5340,N_1480);
or U9094 (N_9094,N_5098,N_4637);
and U9095 (N_9095,N_1083,N_5645);
nor U9096 (N_9096,N_3379,N_1438);
and U9097 (N_9097,N_5546,N_88);
nand U9098 (N_9098,N_5770,N_1996);
or U9099 (N_9099,N_235,N_1801);
nor U9100 (N_9100,N_6110,N_2280);
nand U9101 (N_9101,N_4397,N_1523);
nor U9102 (N_9102,N_165,N_3235);
nand U9103 (N_9103,N_6012,N_2827);
nor U9104 (N_9104,N_1746,N_3181);
or U9105 (N_9105,N_5010,N_5027);
nor U9106 (N_9106,N_1992,N_1345);
nor U9107 (N_9107,N_109,N_5346);
nand U9108 (N_9108,N_788,N_413);
nor U9109 (N_9109,N_578,N_4890);
nand U9110 (N_9110,N_5185,N_4663);
nand U9111 (N_9111,N_2390,N_514);
and U9112 (N_9112,N_2017,N_4168);
nor U9113 (N_9113,N_1122,N_5452);
nor U9114 (N_9114,N_6035,N_3278);
nor U9115 (N_9115,N_2844,N_371);
or U9116 (N_9116,N_4031,N_6217);
or U9117 (N_9117,N_5636,N_2164);
nor U9118 (N_9118,N_5342,N_5956);
nand U9119 (N_9119,N_2615,N_2651);
or U9120 (N_9120,N_6171,N_569);
or U9121 (N_9121,N_3652,N_747);
xnor U9122 (N_9122,N_1207,N_3873);
xor U9123 (N_9123,N_3168,N_2270);
xor U9124 (N_9124,N_725,N_2021);
and U9125 (N_9125,N_2334,N_5821);
xor U9126 (N_9126,N_4235,N_3599);
or U9127 (N_9127,N_451,N_1486);
or U9128 (N_9128,N_4912,N_4291);
or U9129 (N_9129,N_6001,N_773);
nand U9130 (N_9130,N_3556,N_5774);
or U9131 (N_9131,N_3338,N_4666);
or U9132 (N_9132,N_5334,N_4056);
or U9133 (N_9133,N_2611,N_1407);
or U9134 (N_9134,N_5150,N_1372);
xor U9135 (N_9135,N_5923,N_4495);
xnor U9136 (N_9136,N_225,N_4647);
and U9137 (N_9137,N_736,N_1330);
nor U9138 (N_9138,N_257,N_1492);
or U9139 (N_9139,N_1779,N_5281);
nor U9140 (N_9140,N_4904,N_1278);
and U9141 (N_9141,N_5927,N_1993);
or U9142 (N_9142,N_1900,N_1564);
or U9143 (N_9143,N_3616,N_5686);
and U9144 (N_9144,N_3787,N_3554);
nor U9145 (N_9145,N_1817,N_1542);
or U9146 (N_9146,N_5756,N_2035);
or U9147 (N_9147,N_1983,N_2468);
xnor U9148 (N_9148,N_2444,N_6062);
or U9149 (N_9149,N_2075,N_2135);
xor U9150 (N_9150,N_1148,N_892);
and U9151 (N_9151,N_2500,N_4873);
and U9152 (N_9152,N_2502,N_6246);
or U9153 (N_9153,N_5471,N_1357);
nand U9154 (N_9154,N_4930,N_3776);
or U9155 (N_9155,N_3450,N_3687);
xnor U9156 (N_9156,N_4189,N_2103);
and U9157 (N_9157,N_6089,N_106);
or U9158 (N_9158,N_5742,N_5078);
nand U9159 (N_9159,N_3183,N_5908);
nor U9160 (N_9160,N_2132,N_5613);
nor U9161 (N_9161,N_2226,N_4954);
or U9162 (N_9162,N_4630,N_2);
or U9163 (N_9163,N_2815,N_1002);
nand U9164 (N_9164,N_174,N_351);
xnor U9165 (N_9165,N_4118,N_1424);
nand U9166 (N_9166,N_2833,N_122);
nor U9167 (N_9167,N_2112,N_3061);
or U9168 (N_9168,N_5022,N_2644);
xnor U9169 (N_9169,N_5517,N_1032);
and U9170 (N_9170,N_3454,N_2036);
or U9171 (N_9171,N_649,N_4344);
nand U9172 (N_9172,N_1666,N_5354);
nand U9173 (N_9173,N_2357,N_2170);
nand U9174 (N_9174,N_5586,N_1429);
nor U9175 (N_9175,N_538,N_5251);
nand U9176 (N_9176,N_2933,N_4649);
or U9177 (N_9177,N_1084,N_726);
nand U9178 (N_9178,N_2913,N_324);
or U9179 (N_9179,N_3695,N_2287);
or U9180 (N_9180,N_3917,N_2449);
nand U9181 (N_9181,N_591,N_3060);
nor U9182 (N_9182,N_2938,N_3764);
and U9183 (N_9183,N_3008,N_5990);
nand U9184 (N_9184,N_5391,N_4963);
nand U9185 (N_9185,N_4205,N_5243);
xor U9186 (N_9186,N_5137,N_5329);
nand U9187 (N_9187,N_4580,N_6187);
or U9188 (N_9188,N_4019,N_2659);
and U9189 (N_9189,N_5149,N_3239);
nand U9190 (N_9190,N_2955,N_4840);
xnor U9191 (N_9191,N_1691,N_1014);
and U9192 (N_9192,N_4478,N_1347);
or U9193 (N_9193,N_4655,N_3160);
xnor U9194 (N_9194,N_4879,N_3508);
nand U9195 (N_9195,N_4569,N_4519);
xor U9196 (N_9196,N_3407,N_3894);
and U9197 (N_9197,N_2192,N_5728);
xor U9198 (N_9198,N_5664,N_5853);
or U9199 (N_9199,N_5144,N_2652);
and U9200 (N_9200,N_5537,N_3033);
xnor U9201 (N_9201,N_1730,N_5263);
or U9202 (N_9202,N_1467,N_1909);
or U9203 (N_9203,N_1640,N_2263);
nand U9204 (N_9204,N_6048,N_4158);
or U9205 (N_9205,N_3495,N_2654);
nand U9206 (N_9206,N_4265,N_183);
nor U9207 (N_9207,N_3815,N_219);
or U9208 (N_9208,N_5132,N_4061);
and U9209 (N_9209,N_727,N_672);
and U9210 (N_9210,N_2020,N_58);
and U9211 (N_9211,N_6070,N_4337);
xnor U9212 (N_9212,N_5746,N_1583);
and U9213 (N_9213,N_3362,N_5899);
and U9214 (N_9214,N_3190,N_2005);
nand U9215 (N_9215,N_4057,N_2614);
nand U9216 (N_9216,N_2584,N_3713);
nand U9217 (N_9217,N_3028,N_3805);
and U9218 (N_9218,N_6198,N_129);
xnor U9219 (N_9219,N_841,N_5030);
and U9220 (N_9220,N_4286,N_913);
and U9221 (N_9221,N_3103,N_5769);
nand U9222 (N_9222,N_3162,N_1374);
and U9223 (N_9223,N_170,N_3865);
nand U9224 (N_9224,N_4072,N_2211);
nor U9225 (N_9225,N_5966,N_333);
or U9226 (N_9226,N_1205,N_851);
nor U9227 (N_9227,N_2960,N_5292);
or U9228 (N_9228,N_1890,N_1521);
and U9229 (N_9229,N_6232,N_2765);
xnor U9230 (N_9230,N_6015,N_4152);
or U9231 (N_9231,N_2055,N_5603);
xnor U9232 (N_9232,N_3977,N_894);
and U9233 (N_9233,N_2426,N_243);
and U9234 (N_9234,N_4560,N_4170);
or U9235 (N_9235,N_471,N_4352);
xnor U9236 (N_9236,N_681,N_5779);
or U9237 (N_9237,N_5733,N_1383);
xor U9238 (N_9238,N_2373,N_729);
and U9239 (N_9239,N_4339,N_3676);
nor U9240 (N_9240,N_1350,N_4535);
nand U9241 (N_9241,N_168,N_3746);
and U9242 (N_9242,N_2412,N_5025);
xor U9243 (N_9243,N_2451,N_4350);
or U9244 (N_9244,N_5747,N_2403);
nand U9245 (N_9245,N_5633,N_1269);
and U9246 (N_9246,N_1908,N_2583);
nand U9247 (N_9247,N_720,N_101);
nor U9248 (N_9248,N_2351,N_3967);
and U9249 (N_9249,N_5865,N_1923);
or U9250 (N_9250,N_6014,N_5639);
nand U9251 (N_9251,N_3063,N_5580);
or U9252 (N_9252,N_5845,N_1629);
or U9253 (N_9253,N_3096,N_5247);
xnor U9254 (N_9254,N_4860,N_4270);
and U9255 (N_9255,N_1073,N_5970);
nand U9256 (N_9256,N_1342,N_4104);
and U9257 (N_9257,N_1382,N_5162);
or U9258 (N_9258,N_4566,N_3530);
and U9259 (N_9259,N_2490,N_2711);
or U9260 (N_9260,N_1485,N_4921);
nor U9261 (N_9261,N_3662,N_3004);
nor U9262 (N_9262,N_1166,N_4898);
or U9263 (N_9263,N_4334,N_286);
nand U9264 (N_9264,N_4293,N_5711);
nand U9265 (N_9265,N_5002,N_2729);
and U9266 (N_9266,N_5625,N_31);
and U9267 (N_9267,N_6066,N_5933);
or U9268 (N_9268,N_5352,N_304);
or U9269 (N_9269,N_3319,N_3044);
and U9270 (N_9270,N_5904,N_1960);
and U9271 (N_9271,N_1414,N_6008);
nor U9272 (N_9272,N_1129,N_3960);
and U9273 (N_9273,N_5321,N_2004);
or U9274 (N_9274,N_5820,N_2185);
nand U9275 (N_9275,N_1284,N_4318);
or U9276 (N_9276,N_5524,N_4777);
nand U9277 (N_9277,N_1712,N_838);
or U9278 (N_9278,N_3025,N_2413);
nor U9279 (N_9279,N_2727,N_968);
nand U9280 (N_9280,N_2392,N_1292);
nor U9281 (N_9281,N_783,N_1875);
nor U9282 (N_9282,N_770,N_2790);
and U9283 (N_9283,N_4712,N_2331);
and U9284 (N_9284,N_1755,N_2169);
and U9285 (N_9285,N_494,N_1300);
nand U9286 (N_9286,N_1705,N_547);
or U9287 (N_9287,N_3543,N_4551);
nand U9288 (N_9288,N_3012,N_3971);
nor U9289 (N_9289,N_3211,N_2083);
nand U9290 (N_9290,N_387,N_3757);
or U9291 (N_9291,N_1886,N_4492);
xnor U9292 (N_9292,N_4817,N_2885);
nand U9293 (N_9293,N_1685,N_2248);
nand U9294 (N_9294,N_3375,N_6202);
nor U9295 (N_9295,N_2275,N_2076);
nand U9296 (N_9296,N_185,N_44);
nand U9297 (N_9297,N_5936,N_1714);
nand U9298 (N_9298,N_794,N_2598);
xor U9299 (N_9299,N_6231,N_3419);
nand U9300 (N_9300,N_707,N_4338);
nor U9301 (N_9301,N_3188,N_642);
or U9302 (N_9302,N_676,N_2918);
or U9303 (N_9303,N_5668,N_355);
and U9304 (N_9304,N_3248,N_3223);
or U9305 (N_9305,N_3346,N_3487);
nor U9306 (N_9306,N_1391,N_6080);
nor U9307 (N_9307,N_5832,N_5401);
xor U9308 (N_9308,N_4458,N_2520);
and U9309 (N_9309,N_6235,N_5100);
nand U9310 (N_9310,N_1222,N_1606);
and U9311 (N_9311,N_291,N_1870);
or U9312 (N_9312,N_5215,N_4113);
and U9313 (N_9313,N_1238,N_5067);
nand U9314 (N_9314,N_3810,N_5628);
or U9315 (N_9315,N_2627,N_230);
nand U9316 (N_9316,N_962,N_3760);
and U9317 (N_9317,N_5846,N_2319);
nand U9318 (N_9318,N_5374,N_3845);
and U9319 (N_9319,N_4885,N_5451);
or U9320 (N_9320,N_157,N_5024);
nand U9321 (N_9321,N_6177,N_4957);
nand U9322 (N_9322,N_5530,N_4355);
and U9323 (N_9323,N_466,N_4564);
nand U9324 (N_9324,N_271,N_2024);
or U9325 (N_9325,N_5262,N_4039);
nand U9326 (N_9326,N_4822,N_5602);
nor U9327 (N_9327,N_2282,N_3281);
or U9328 (N_9328,N_3571,N_4144);
and U9329 (N_9329,N_564,N_4861);
nand U9330 (N_9330,N_3274,N_1320);
or U9331 (N_9331,N_2951,N_4014);
xor U9332 (N_9332,N_3553,N_1823);
nand U9333 (N_9333,N_1518,N_765);
or U9334 (N_9334,N_1882,N_6194);
nand U9335 (N_9335,N_4789,N_2768);
nand U9336 (N_9336,N_5860,N_3952);
or U9337 (N_9337,N_4643,N_5175);
or U9338 (N_9338,N_3187,N_3769);
or U9339 (N_9339,N_1018,N_1633);
and U9340 (N_9340,N_5798,N_3747);
and U9341 (N_9341,N_3906,N_1843);
nor U9342 (N_9342,N_5847,N_677);
nand U9343 (N_9343,N_3423,N_1329);
and U9344 (N_9344,N_2080,N_2191);
nand U9345 (N_9345,N_1818,N_4493);
and U9346 (N_9346,N_502,N_5086);
nand U9347 (N_9347,N_1068,N_2166);
nor U9348 (N_9348,N_1721,N_2367);
nand U9349 (N_9349,N_2943,N_1733);
or U9350 (N_9350,N_1021,N_801);
nor U9351 (N_9351,N_3668,N_1790);
nand U9352 (N_9352,N_1827,N_5713);
or U9353 (N_9353,N_3112,N_1780);
nand U9354 (N_9354,N_2633,N_2985);
nand U9355 (N_9355,N_2177,N_4992);
or U9356 (N_9356,N_3832,N_4892);
nand U9357 (N_9357,N_2714,N_4448);
xnor U9358 (N_9358,N_4625,N_1589);
xnor U9359 (N_9359,N_628,N_180);
nand U9360 (N_9360,N_595,N_1532);
nor U9361 (N_9361,N_2515,N_926);
or U9362 (N_9362,N_3109,N_4958);
or U9363 (N_9363,N_5833,N_4304);
nor U9364 (N_9364,N_216,N_4701);
or U9365 (N_9365,N_805,N_5890);
nand U9366 (N_9366,N_571,N_2716);
nand U9367 (N_9367,N_3176,N_5083);
xor U9368 (N_9368,N_1071,N_1104);
nor U9369 (N_9369,N_5758,N_5140);
or U9370 (N_9370,N_2948,N_675);
or U9371 (N_9371,N_3206,N_455);
and U9372 (N_9372,N_4115,N_4038);
or U9373 (N_9373,N_3479,N_5312);
or U9374 (N_9374,N_5873,N_2874);
or U9375 (N_9375,N_4709,N_6221);
nand U9376 (N_9376,N_1974,N_4250);
nand U9377 (N_9377,N_1896,N_2067);
nor U9378 (N_9378,N_1002,N_4868);
and U9379 (N_9379,N_3267,N_3261);
xor U9380 (N_9380,N_4798,N_6054);
or U9381 (N_9381,N_2082,N_2885);
and U9382 (N_9382,N_2610,N_5906);
nand U9383 (N_9383,N_34,N_5668);
and U9384 (N_9384,N_3037,N_2070);
or U9385 (N_9385,N_3441,N_4990);
or U9386 (N_9386,N_5624,N_5653);
nand U9387 (N_9387,N_3579,N_4032);
and U9388 (N_9388,N_346,N_3810);
or U9389 (N_9389,N_4888,N_6224);
nor U9390 (N_9390,N_4214,N_3439);
or U9391 (N_9391,N_4092,N_716);
or U9392 (N_9392,N_4880,N_5194);
nor U9393 (N_9393,N_2169,N_2409);
nor U9394 (N_9394,N_374,N_4135);
nand U9395 (N_9395,N_5282,N_5116);
or U9396 (N_9396,N_4529,N_6094);
and U9397 (N_9397,N_3936,N_1250);
nand U9398 (N_9398,N_2202,N_2212);
or U9399 (N_9399,N_4533,N_4068);
or U9400 (N_9400,N_3187,N_2044);
or U9401 (N_9401,N_1419,N_2043);
or U9402 (N_9402,N_5817,N_4552);
or U9403 (N_9403,N_5983,N_2892);
or U9404 (N_9404,N_1186,N_2793);
nor U9405 (N_9405,N_2665,N_1128);
and U9406 (N_9406,N_5156,N_1075);
or U9407 (N_9407,N_5048,N_5152);
xnor U9408 (N_9408,N_780,N_6145);
nand U9409 (N_9409,N_2264,N_465);
or U9410 (N_9410,N_6199,N_5577);
nand U9411 (N_9411,N_1791,N_1644);
nand U9412 (N_9412,N_2845,N_4166);
nor U9413 (N_9413,N_1205,N_2656);
nor U9414 (N_9414,N_3031,N_614);
nor U9415 (N_9415,N_4441,N_5487);
nand U9416 (N_9416,N_2338,N_5361);
xnor U9417 (N_9417,N_4048,N_3456);
or U9418 (N_9418,N_5946,N_1211);
and U9419 (N_9419,N_3417,N_3519);
nand U9420 (N_9420,N_6142,N_4385);
and U9421 (N_9421,N_1518,N_4848);
nor U9422 (N_9422,N_4243,N_4481);
nand U9423 (N_9423,N_5235,N_2255);
xnor U9424 (N_9424,N_1980,N_2055);
xnor U9425 (N_9425,N_4831,N_158);
xor U9426 (N_9426,N_1266,N_341);
nor U9427 (N_9427,N_61,N_3038);
xor U9428 (N_9428,N_5014,N_3652);
or U9429 (N_9429,N_682,N_3515);
nand U9430 (N_9430,N_3497,N_1454);
and U9431 (N_9431,N_1925,N_5239);
nor U9432 (N_9432,N_496,N_1016);
nand U9433 (N_9433,N_2150,N_6221);
nor U9434 (N_9434,N_3983,N_3066);
nor U9435 (N_9435,N_5606,N_756);
xnor U9436 (N_9436,N_4490,N_1953);
and U9437 (N_9437,N_2954,N_3291);
nand U9438 (N_9438,N_1560,N_2124);
or U9439 (N_9439,N_2027,N_4127);
nand U9440 (N_9440,N_4912,N_5585);
and U9441 (N_9441,N_1992,N_4356);
nand U9442 (N_9442,N_1608,N_5300);
nor U9443 (N_9443,N_1457,N_5579);
nor U9444 (N_9444,N_2997,N_2711);
xor U9445 (N_9445,N_2625,N_5897);
and U9446 (N_9446,N_1827,N_808);
and U9447 (N_9447,N_2633,N_1974);
nor U9448 (N_9448,N_5036,N_6154);
nand U9449 (N_9449,N_6110,N_4638);
nand U9450 (N_9450,N_2179,N_5816);
nand U9451 (N_9451,N_5894,N_1070);
nor U9452 (N_9452,N_2305,N_4539);
and U9453 (N_9453,N_961,N_1351);
or U9454 (N_9454,N_4873,N_5523);
and U9455 (N_9455,N_542,N_1210);
and U9456 (N_9456,N_3197,N_6082);
or U9457 (N_9457,N_4017,N_4208);
nor U9458 (N_9458,N_3986,N_3232);
or U9459 (N_9459,N_2429,N_385);
nor U9460 (N_9460,N_1265,N_425);
nand U9461 (N_9461,N_1130,N_6056);
xor U9462 (N_9462,N_5805,N_862);
and U9463 (N_9463,N_6246,N_440);
and U9464 (N_9464,N_715,N_3270);
and U9465 (N_9465,N_187,N_1811);
nor U9466 (N_9466,N_5774,N_5683);
and U9467 (N_9467,N_2530,N_300);
nor U9468 (N_9468,N_2174,N_5481);
nor U9469 (N_9469,N_219,N_2620);
xor U9470 (N_9470,N_6243,N_2544);
or U9471 (N_9471,N_1808,N_2787);
and U9472 (N_9472,N_3759,N_1013);
nand U9473 (N_9473,N_5225,N_4684);
nor U9474 (N_9474,N_4224,N_3889);
or U9475 (N_9475,N_4821,N_5728);
nand U9476 (N_9476,N_2877,N_3478);
and U9477 (N_9477,N_4365,N_4058);
nor U9478 (N_9478,N_3885,N_5715);
or U9479 (N_9479,N_5640,N_254);
nand U9480 (N_9480,N_76,N_1809);
and U9481 (N_9481,N_1738,N_6214);
nand U9482 (N_9482,N_1910,N_958);
nand U9483 (N_9483,N_4466,N_3287);
and U9484 (N_9484,N_2379,N_270);
nand U9485 (N_9485,N_5297,N_3337);
nand U9486 (N_9486,N_1893,N_5008);
or U9487 (N_9487,N_2796,N_2372);
or U9488 (N_9488,N_2267,N_1475);
nand U9489 (N_9489,N_2241,N_2528);
or U9490 (N_9490,N_5505,N_2134);
nand U9491 (N_9491,N_2886,N_4693);
nand U9492 (N_9492,N_5138,N_3322);
xor U9493 (N_9493,N_630,N_6029);
nor U9494 (N_9494,N_1677,N_4944);
and U9495 (N_9495,N_3814,N_3205);
nor U9496 (N_9496,N_1208,N_4026);
and U9497 (N_9497,N_1985,N_2992);
or U9498 (N_9498,N_4484,N_4153);
and U9499 (N_9499,N_5253,N_3649);
nor U9500 (N_9500,N_3710,N_5301);
nor U9501 (N_9501,N_3857,N_4982);
xnor U9502 (N_9502,N_5435,N_4721);
and U9503 (N_9503,N_2768,N_2009);
xor U9504 (N_9504,N_4440,N_1821);
and U9505 (N_9505,N_6075,N_3060);
xnor U9506 (N_9506,N_4165,N_5146);
xor U9507 (N_9507,N_2848,N_4174);
or U9508 (N_9508,N_5955,N_2625);
and U9509 (N_9509,N_2916,N_1067);
or U9510 (N_9510,N_5214,N_2349);
or U9511 (N_9511,N_575,N_4814);
xor U9512 (N_9512,N_1146,N_3097);
or U9513 (N_9513,N_398,N_1344);
or U9514 (N_9514,N_4902,N_4303);
nor U9515 (N_9515,N_3163,N_2017);
and U9516 (N_9516,N_956,N_5063);
and U9517 (N_9517,N_5889,N_4153);
nand U9518 (N_9518,N_639,N_1251);
or U9519 (N_9519,N_243,N_4894);
nor U9520 (N_9520,N_5258,N_326);
or U9521 (N_9521,N_2480,N_1286);
and U9522 (N_9522,N_5674,N_3526);
nand U9523 (N_9523,N_1755,N_515);
nor U9524 (N_9524,N_3786,N_4609);
xnor U9525 (N_9525,N_5087,N_4298);
or U9526 (N_9526,N_2311,N_4437);
xnor U9527 (N_9527,N_796,N_4190);
or U9528 (N_9528,N_5479,N_5778);
or U9529 (N_9529,N_3262,N_4845);
xor U9530 (N_9530,N_4630,N_961);
or U9531 (N_9531,N_3051,N_5525);
xnor U9532 (N_9532,N_411,N_5850);
or U9533 (N_9533,N_3791,N_222);
and U9534 (N_9534,N_1207,N_2078);
xor U9535 (N_9535,N_3965,N_2290);
or U9536 (N_9536,N_4478,N_5891);
nor U9537 (N_9537,N_2020,N_2619);
or U9538 (N_9538,N_1085,N_829);
nand U9539 (N_9539,N_5914,N_166);
or U9540 (N_9540,N_4474,N_522);
nor U9541 (N_9541,N_4506,N_21);
nor U9542 (N_9542,N_1986,N_1717);
nand U9543 (N_9543,N_4484,N_111);
or U9544 (N_9544,N_477,N_5225);
nand U9545 (N_9545,N_4994,N_6184);
xor U9546 (N_9546,N_3839,N_5097);
nor U9547 (N_9547,N_3827,N_1157);
nor U9548 (N_9548,N_3601,N_5775);
or U9549 (N_9549,N_2565,N_5123);
xor U9550 (N_9550,N_3085,N_1060);
nor U9551 (N_9551,N_212,N_4960);
and U9552 (N_9552,N_1284,N_4899);
xnor U9553 (N_9553,N_1020,N_5648);
nor U9554 (N_9554,N_3982,N_3909);
xor U9555 (N_9555,N_2516,N_3030);
xor U9556 (N_9556,N_1176,N_3226);
or U9557 (N_9557,N_1425,N_4511);
or U9558 (N_9558,N_1096,N_6183);
and U9559 (N_9559,N_294,N_3617);
nor U9560 (N_9560,N_3873,N_2627);
nand U9561 (N_9561,N_5469,N_3559);
and U9562 (N_9562,N_5979,N_5074);
nor U9563 (N_9563,N_2215,N_2564);
xor U9564 (N_9564,N_3093,N_5983);
nor U9565 (N_9565,N_5741,N_6114);
xnor U9566 (N_9566,N_2582,N_3544);
or U9567 (N_9567,N_376,N_4898);
nand U9568 (N_9568,N_2949,N_5735);
and U9569 (N_9569,N_2134,N_567);
nor U9570 (N_9570,N_4573,N_4924);
or U9571 (N_9571,N_2315,N_2673);
nand U9572 (N_9572,N_288,N_4774);
nand U9573 (N_9573,N_2057,N_2765);
nor U9574 (N_9574,N_2504,N_1074);
or U9575 (N_9575,N_2719,N_3907);
nand U9576 (N_9576,N_4462,N_1477);
and U9577 (N_9577,N_1944,N_3892);
nand U9578 (N_9578,N_1535,N_1268);
nor U9579 (N_9579,N_4243,N_4496);
and U9580 (N_9580,N_2856,N_5197);
and U9581 (N_9581,N_4093,N_3529);
nor U9582 (N_9582,N_4886,N_5832);
nor U9583 (N_9583,N_3881,N_2403);
nor U9584 (N_9584,N_1437,N_2365);
or U9585 (N_9585,N_6105,N_4141);
and U9586 (N_9586,N_5114,N_3416);
nor U9587 (N_9587,N_1200,N_1377);
and U9588 (N_9588,N_4161,N_4461);
nand U9589 (N_9589,N_5871,N_4193);
nor U9590 (N_9590,N_3255,N_3458);
and U9591 (N_9591,N_2549,N_5802);
nor U9592 (N_9592,N_607,N_4709);
nor U9593 (N_9593,N_194,N_733);
or U9594 (N_9594,N_3529,N_2907);
nand U9595 (N_9595,N_4294,N_4389);
nor U9596 (N_9596,N_4871,N_2825);
and U9597 (N_9597,N_4240,N_5329);
nand U9598 (N_9598,N_1815,N_328);
xor U9599 (N_9599,N_5059,N_4008);
and U9600 (N_9600,N_4098,N_5861);
and U9601 (N_9601,N_3377,N_2161);
nand U9602 (N_9602,N_2394,N_1189);
xor U9603 (N_9603,N_1449,N_2229);
xnor U9604 (N_9604,N_993,N_3393);
and U9605 (N_9605,N_5929,N_4477);
or U9606 (N_9606,N_1274,N_4655);
nand U9607 (N_9607,N_3918,N_4937);
or U9608 (N_9608,N_5073,N_3079);
and U9609 (N_9609,N_4633,N_149);
nor U9610 (N_9610,N_1254,N_1286);
nand U9611 (N_9611,N_5146,N_3244);
or U9612 (N_9612,N_1081,N_554);
nor U9613 (N_9613,N_4008,N_3899);
or U9614 (N_9614,N_4161,N_2982);
or U9615 (N_9615,N_4768,N_3699);
or U9616 (N_9616,N_3712,N_2046);
nand U9617 (N_9617,N_177,N_6138);
and U9618 (N_9618,N_3876,N_1043);
nand U9619 (N_9619,N_2895,N_442);
nand U9620 (N_9620,N_1962,N_49);
or U9621 (N_9621,N_1086,N_6099);
nor U9622 (N_9622,N_4470,N_3774);
nand U9623 (N_9623,N_5984,N_1166);
and U9624 (N_9624,N_4552,N_5152);
nand U9625 (N_9625,N_2111,N_6106);
or U9626 (N_9626,N_6158,N_4642);
xnor U9627 (N_9627,N_4859,N_3018);
or U9628 (N_9628,N_797,N_3657);
or U9629 (N_9629,N_5627,N_165);
nand U9630 (N_9630,N_2436,N_2494);
nand U9631 (N_9631,N_4834,N_2604);
and U9632 (N_9632,N_4554,N_1849);
nand U9633 (N_9633,N_1682,N_1903);
nand U9634 (N_9634,N_6165,N_4751);
nor U9635 (N_9635,N_4720,N_5070);
nand U9636 (N_9636,N_5100,N_5946);
xor U9637 (N_9637,N_50,N_1466);
or U9638 (N_9638,N_3248,N_5300);
or U9639 (N_9639,N_3517,N_3820);
nor U9640 (N_9640,N_3457,N_1880);
or U9641 (N_9641,N_4106,N_2602);
xnor U9642 (N_9642,N_6130,N_1635);
or U9643 (N_9643,N_6234,N_4151);
xor U9644 (N_9644,N_2410,N_1713);
xnor U9645 (N_9645,N_4799,N_570);
or U9646 (N_9646,N_5450,N_777);
nor U9647 (N_9647,N_673,N_1499);
nand U9648 (N_9648,N_78,N_2120);
and U9649 (N_9649,N_3752,N_827);
nor U9650 (N_9650,N_592,N_91);
nor U9651 (N_9651,N_663,N_1145);
xnor U9652 (N_9652,N_2017,N_3930);
or U9653 (N_9653,N_3054,N_5194);
and U9654 (N_9654,N_2659,N_2308);
nand U9655 (N_9655,N_5779,N_2765);
nor U9656 (N_9656,N_882,N_372);
nand U9657 (N_9657,N_4982,N_5258);
xor U9658 (N_9658,N_90,N_2500);
nand U9659 (N_9659,N_2912,N_3668);
nand U9660 (N_9660,N_6157,N_2826);
xnor U9661 (N_9661,N_26,N_484);
nor U9662 (N_9662,N_5666,N_667);
nor U9663 (N_9663,N_244,N_6221);
or U9664 (N_9664,N_179,N_611);
nand U9665 (N_9665,N_3604,N_6008);
and U9666 (N_9666,N_852,N_98);
or U9667 (N_9667,N_3898,N_15);
nor U9668 (N_9668,N_3516,N_4936);
and U9669 (N_9669,N_897,N_5595);
nand U9670 (N_9670,N_4679,N_1843);
nand U9671 (N_9671,N_3767,N_673);
nand U9672 (N_9672,N_5824,N_167);
nand U9673 (N_9673,N_1938,N_5140);
nor U9674 (N_9674,N_5835,N_4779);
xor U9675 (N_9675,N_2461,N_2465);
or U9676 (N_9676,N_4341,N_1740);
and U9677 (N_9677,N_5858,N_3472);
nor U9678 (N_9678,N_4084,N_1104);
nand U9679 (N_9679,N_2766,N_255);
and U9680 (N_9680,N_2888,N_4566);
nand U9681 (N_9681,N_5481,N_5800);
or U9682 (N_9682,N_495,N_4061);
and U9683 (N_9683,N_3919,N_5847);
or U9684 (N_9684,N_2073,N_1764);
xnor U9685 (N_9685,N_5049,N_3289);
and U9686 (N_9686,N_5302,N_2445);
nand U9687 (N_9687,N_641,N_3563);
and U9688 (N_9688,N_4851,N_1063);
or U9689 (N_9689,N_1632,N_5528);
or U9690 (N_9690,N_5532,N_134);
nor U9691 (N_9691,N_4114,N_5084);
nor U9692 (N_9692,N_877,N_4325);
nor U9693 (N_9693,N_1878,N_2198);
and U9694 (N_9694,N_5498,N_5622);
nor U9695 (N_9695,N_5993,N_1024);
or U9696 (N_9696,N_536,N_988);
or U9697 (N_9697,N_296,N_3488);
nand U9698 (N_9698,N_5101,N_5342);
and U9699 (N_9699,N_1143,N_2471);
nand U9700 (N_9700,N_5424,N_873);
nor U9701 (N_9701,N_5700,N_2720);
and U9702 (N_9702,N_6026,N_5608);
nor U9703 (N_9703,N_2329,N_5313);
nor U9704 (N_9704,N_1728,N_3904);
nand U9705 (N_9705,N_1891,N_4375);
or U9706 (N_9706,N_4317,N_277);
or U9707 (N_9707,N_1108,N_3632);
nand U9708 (N_9708,N_4831,N_3010);
and U9709 (N_9709,N_2600,N_2772);
nand U9710 (N_9710,N_3551,N_1573);
nor U9711 (N_9711,N_2020,N_4759);
or U9712 (N_9712,N_1424,N_6014);
nor U9713 (N_9713,N_3837,N_3342);
xor U9714 (N_9714,N_720,N_3088);
or U9715 (N_9715,N_2693,N_2460);
nand U9716 (N_9716,N_4792,N_227);
or U9717 (N_9717,N_3083,N_4060);
or U9718 (N_9718,N_4249,N_2446);
nor U9719 (N_9719,N_2105,N_2821);
and U9720 (N_9720,N_451,N_3453);
and U9721 (N_9721,N_3155,N_3901);
nor U9722 (N_9722,N_4783,N_3812);
xnor U9723 (N_9723,N_4998,N_4180);
nand U9724 (N_9724,N_1154,N_161);
or U9725 (N_9725,N_5485,N_964);
nor U9726 (N_9726,N_5772,N_2146);
nor U9727 (N_9727,N_4276,N_515);
and U9728 (N_9728,N_2129,N_3495);
xnor U9729 (N_9729,N_5932,N_3260);
nor U9730 (N_9730,N_2090,N_1324);
nor U9731 (N_9731,N_1202,N_3257);
nand U9732 (N_9732,N_4793,N_3768);
and U9733 (N_9733,N_1049,N_3381);
or U9734 (N_9734,N_6092,N_1086);
or U9735 (N_9735,N_570,N_1432);
and U9736 (N_9736,N_3877,N_3378);
nor U9737 (N_9737,N_5423,N_5644);
nand U9738 (N_9738,N_2343,N_5250);
nand U9739 (N_9739,N_3299,N_2203);
nor U9740 (N_9740,N_5903,N_4460);
or U9741 (N_9741,N_6231,N_4145);
nand U9742 (N_9742,N_2845,N_3455);
nand U9743 (N_9743,N_898,N_4235);
nand U9744 (N_9744,N_5211,N_1181);
or U9745 (N_9745,N_3761,N_5659);
nor U9746 (N_9746,N_2770,N_1438);
nor U9747 (N_9747,N_5249,N_3129);
nor U9748 (N_9748,N_2530,N_4631);
nand U9749 (N_9749,N_4066,N_361);
xor U9750 (N_9750,N_197,N_5261);
or U9751 (N_9751,N_3396,N_1240);
and U9752 (N_9752,N_2204,N_4451);
xor U9753 (N_9753,N_2904,N_3115);
nor U9754 (N_9754,N_4058,N_5759);
and U9755 (N_9755,N_497,N_2680);
nand U9756 (N_9756,N_3452,N_56);
and U9757 (N_9757,N_709,N_1271);
or U9758 (N_9758,N_6229,N_171);
nand U9759 (N_9759,N_358,N_723);
nand U9760 (N_9760,N_411,N_1);
and U9761 (N_9761,N_973,N_5374);
and U9762 (N_9762,N_3300,N_5559);
nor U9763 (N_9763,N_4248,N_5920);
or U9764 (N_9764,N_3271,N_52);
and U9765 (N_9765,N_43,N_3144);
nor U9766 (N_9766,N_5389,N_1805);
nor U9767 (N_9767,N_432,N_5978);
xor U9768 (N_9768,N_3019,N_2198);
nand U9769 (N_9769,N_2082,N_4147);
nor U9770 (N_9770,N_5381,N_250);
or U9771 (N_9771,N_5274,N_471);
nor U9772 (N_9772,N_2933,N_1301);
nand U9773 (N_9773,N_6196,N_2846);
or U9774 (N_9774,N_5928,N_292);
nor U9775 (N_9775,N_5020,N_4298);
or U9776 (N_9776,N_5070,N_3637);
or U9777 (N_9777,N_1501,N_3887);
and U9778 (N_9778,N_631,N_5189);
and U9779 (N_9779,N_5322,N_5970);
or U9780 (N_9780,N_366,N_2099);
and U9781 (N_9781,N_4556,N_5765);
and U9782 (N_9782,N_1290,N_1555);
nand U9783 (N_9783,N_177,N_2052);
or U9784 (N_9784,N_2620,N_2347);
and U9785 (N_9785,N_5491,N_2361);
nor U9786 (N_9786,N_6159,N_5707);
and U9787 (N_9787,N_1474,N_3450);
nand U9788 (N_9788,N_2202,N_5342);
and U9789 (N_9789,N_3521,N_4550);
nor U9790 (N_9790,N_4405,N_4669);
nor U9791 (N_9791,N_2622,N_4561);
xnor U9792 (N_9792,N_1525,N_3225);
and U9793 (N_9793,N_2117,N_903);
nor U9794 (N_9794,N_5342,N_3294);
and U9795 (N_9795,N_5963,N_2818);
nor U9796 (N_9796,N_2804,N_6184);
nand U9797 (N_9797,N_2044,N_3998);
or U9798 (N_9798,N_2975,N_4086);
nor U9799 (N_9799,N_2089,N_1085);
and U9800 (N_9800,N_451,N_4584);
xnor U9801 (N_9801,N_3702,N_5038);
or U9802 (N_9802,N_2371,N_555);
nor U9803 (N_9803,N_3770,N_4682);
nand U9804 (N_9804,N_872,N_3547);
or U9805 (N_9805,N_3456,N_3515);
or U9806 (N_9806,N_1227,N_3462);
nor U9807 (N_9807,N_3339,N_6184);
nor U9808 (N_9808,N_4741,N_5938);
nand U9809 (N_9809,N_3758,N_5351);
or U9810 (N_9810,N_4599,N_3572);
or U9811 (N_9811,N_2020,N_715);
xnor U9812 (N_9812,N_4247,N_5967);
or U9813 (N_9813,N_3701,N_5792);
nor U9814 (N_9814,N_5582,N_2673);
nand U9815 (N_9815,N_2555,N_3617);
or U9816 (N_9816,N_5667,N_1248);
nor U9817 (N_9817,N_1070,N_2717);
or U9818 (N_9818,N_2280,N_5505);
nand U9819 (N_9819,N_6006,N_1837);
nand U9820 (N_9820,N_4736,N_5652);
nand U9821 (N_9821,N_2985,N_6040);
nor U9822 (N_9822,N_505,N_2628);
or U9823 (N_9823,N_1275,N_3257);
and U9824 (N_9824,N_58,N_2684);
and U9825 (N_9825,N_2430,N_282);
or U9826 (N_9826,N_1104,N_5423);
nor U9827 (N_9827,N_4660,N_1729);
nand U9828 (N_9828,N_5698,N_4269);
nand U9829 (N_9829,N_1641,N_5749);
or U9830 (N_9830,N_1315,N_820);
or U9831 (N_9831,N_3638,N_6216);
nor U9832 (N_9832,N_3560,N_4178);
nand U9833 (N_9833,N_3543,N_5249);
nor U9834 (N_9834,N_5255,N_2530);
nand U9835 (N_9835,N_3283,N_3261);
or U9836 (N_9836,N_2727,N_5801);
or U9837 (N_9837,N_5919,N_5129);
nor U9838 (N_9838,N_1414,N_2835);
nand U9839 (N_9839,N_1180,N_1722);
or U9840 (N_9840,N_990,N_1783);
nor U9841 (N_9841,N_2497,N_1418);
and U9842 (N_9842,N_1596,N_2976);
and U9843 (N_9843,N_545,N_1658);
nor U9844 (N_9844,N_6244,N_4372);
nor U9845 (N_9845,N_2630,N_3662);
xnor U9846 (N_9846,N_858,N_3162);
or U9847 (N_9847,N_5286,N_4667);
nor U9848 (N_9848,N_408,N_104);
or U9849 (N_9849,N_3771,N_1452);
or U9850 (N_9850,N_2302,N_3054);
and U9851 (N_9851,N_3927,N_3028);
and U9852 (N_9852,N_4406,N_3633);
or U9853 (N_9853,N_6127,N_5399);
and U9854 (N_9854,N_2657,N_3379);
nor U9855 (N_9855,N_4594,N_2127);
or U9856 (N_9856,N_3240,N_3454);
nor U9857 (N_9857,N_5450,N_539);
and U9858 (N_9858,N_2530,N_5614);
and U9859 (N_9859,N_5426,N_309);
or U9860 (N_9860,N_3201,N_4088);
nand U9861 (N_9861,N_4800,N_3855);
nor U9862 (N_9862,N_1284,N_3611);
and U9863 (N_9863,N_1250,N_5814);
xor U9864 (N_9864,N_4473,N_2167);
and U9865 (N_9865,N_939,N_4922);
nor U9866 (N_9866,N_780,N_5746);
nand U9867 (N_9867,N_1275,N_722);
xnor U9868 (N_9868,N_1895,N_162);
nor U9869 (N_9869,N_40,N_5966);
or U9870 (N_9870,N_4274,N_314);
nand U9871 (N_9871,N_1586,N_4291);
or U9872 (N_9872,N_4411,N_3728);
nor U9873 (N_9873,N_393,N_3120);
nand U9874 (N_9874,N_5961,N_1652);
xor U9875 (N_9875,N_1812,N_5517);
nor U9876 (N_9876,N_3454,N_1333);
and U9877 (N_9877,N_4262,N_1534);
nand U9878 (N_9878,N_3039,N_5567);
nand U9879 (N_9879,N_1230,N_2231);
nand U9880 (N_9880,N_4586,N_3349);
and U9881 (N_9881,N_4559,N_2475);
nand U9882 (N_9882,N_3826,N_3028);
or U9883 (N_9883,N_486,N_3240);
or U9884 (N_9884,N_2256,N_3811);
and U9885 (N_9885,N_1896,N_4991);
nand U9886 (N_9886,N_768,N_4004);
xnor U9887 (N_9887,N_2426,N_4207);
or U9888 (N_9888,N_572,N_6223);
or U9889 (N_9889,N_2445,N_2892);
and U9890 (N_9890,N_803,N_3739);
and U9891 (N_9891,N_1177,N_5520);
or U9892 (N_9892,N_3013,N_3875);
or U9893 (N_9893,N_1000,N_1768);
nor U9894 (N_9894,N_1340,N_1200);
nor U9895 (N_9895,N_2645,N_337);
nor U9896 (N_9896,N_2370,N_190);
or U9897 (N_9897,N_1380,N_3529);
and U9898 (N_9898,N_4856,N_6018);
xor U9899 (N_9899,N_5721,N_3965);
nor U9900 (N_9900,N_809,N_3986);
or U9901 (N_9901,N_1360,N_5403);
and U9902 (N_9902,N_4777,N_308);
nor U9903 (N_9903,N_5472,N_592);
or U9904 (N_9904,N_23,N_1726);
nand U9905 (N_9905,N_2281,N_125);
xnor U9906 (N_9906,N_5270,N_2694);
or U9907 (N_9907,N_5917,N_5797);
nor U9908 (N_9908,N_246,N_5717);
nor U9909 (N_9909,N_2456,N_469);
xor U9910 (N_9910,N_1473,N_5280);
or U9911 (N_9911,N_3145,N_4733);
nor U9912 (N_9912,N_3207,N_5898);
nand U9913 (N_9913,N_784,N_5576);
or U9914 (N_9914,N_1960,N_194);
and U9915 (N_9915,N_608,N_483);
nor U9916 (N_9916,N_4877,N_4686);
nand U9917 (N_9917,N_4534,N_2969);
and U9918 (N_9918,N_5154,N_1647);
nand U9919 (N_9919,N_5355,N_2481);
xnor U9920 (N_9920,N_624,N_5453);
nor U9921 (N_9921,N_2051,N_5677);
nand U9922 (N_9922,N_2980,N_5833);
and U9923 (N_9923,N_2856,N_5676);
nand U9924 (N_9924,N_3926,N_2749);
or U9925 (N_9925,N_4835,N_834);
nor U9926 (N_9926,N_1169,N_3885);
nor U9927 (N_9927,N_5951,N_921);
xor U9928 (N_9928,N_3938,N_908);
or U9929 (N_9929,N_2074,N_3336);
nand U9930 (N_9930,N_3304,N_2364);
nand U9931 (N_9931,N_2088,N_6170);
or U9932 (N_9932,N_635,N_2812);
or U9933 (N_9933,N_265,N_4473);
and U9934 (N_9934,N_2327,N_409);
nand U9935 (N_9935,N_5289,N_1226);
nand U9936 (N_9936,N_6053,N_2572);
nor U9937 (N_9937,N_4206,N_2099);
and U9938 (N_9938,N_4365,N_4255);
or U9939 (N_9939,N_2394,N_5498);
or U9940 (N_9940,N_3249,N_4758);
or U9941 (N_9941,N_4227,N_1651);
nor U9942 (N_9942,N_1759,N_5839);
and U9943 (N_9943,N_3594,N_3954);
nor U9944 (N_9944,N_2164,N_5219);
nand U9945 (N_9945,N_411,N_3076);
and U9946 (N_9946,N_178,N_3077);
or U9947 (N_9947,N_1164,N_3474);
or U9948 (N_9948,N_4215,N_950);
nor U9949 (N_9949,N_3798,N_4655);
nand U9950 (N_9950,N_5519,N_1597);
nor U9951 (N_9951,N_3809,N_495);
and U9952 (N_9952,N_5572,N_3457);
and U9953 (N_9953,N_3040,N_3105);
nor U9954 (N_9954,N_5707,N_1871);
nor U9955 (N_9955,N_2284,N_2170);
or U9956 (N_9956,N_4639,N_817);
and U9957 (N_9957,N_6074,N_2492);
and U9958 (N_9958,N_5823,N_1203);
and U9959 (N_9959,N_6138,N_627);
nand U9960 (N_9960,N_4289,N_1262);
nor U9961 (N_9961,N_2410,N_4037);
nand U9962 (N_9962,N_573,N_5624);
and U9963 (N_9963,N_2430,N_5767);
or U9964 (N_9964,N_2346,N_773);
nor U9965 (N_9965,N_890,N_1903);
or U9966 (N_9966,N_1317,N_2434);
or U9967 (N_9967,N_1654,N_1508);
nand U9968 (N_9968,N_5433,N_1851);
or U9969 (N_9969,N_6227,N_1538);
nand U9970 (N_9970,N_2587,N_6237);
and U9971 (N_9971,N_4368,N_2723);
nand U9972 (N_9972,N_540,N_823);
nand U9973 (N_9973,N_1102,N_208);
nand U9974 (N_9974,N_1026,N_555);
nand U9975 (N_9975,N_1375,N_3588);
nand U9976 (N_9976,N_239,N_3879);
and U9977 (N_9977,N_5751,N_2756);
and U9978 (N_9978,N_2339,N_778);
nor U9979 (N_9979,N_5088,N_5591);
nor U9980 (N_9980,N_1054,N_6173);
or U9981 (N_9981,N_2717,N_4906);
or U9982 (N_9982,N_5224,N_126);
or U9983 (N_9983,N_3890,N_414);
and U9984 (N_9984,N_4938,N_4252);
nor U9985 (N_9985,N_2592,N_901);
and U9986 (N_9986,N_2421,N_3565);
or U9987 (N_9987,N_3769,N_3753);
or U9988 (N_9988,N_5649,N_6055);
and U9989 (N_9989,N_4929,N_5507);
nor U9990 (N_9990,N_1908,N_647);
nor U9991 (N_9991,N_5589,N_2459);
or U9992 (N_9992,N_4642,N_633);
nor U9993 (N_9993,N_1881,N_4536);
nor U9994 (N_9994,N_473,N_1455);
or U9995 (N_9995,N_3692,N_3874);
xnor U9996 (N_9996,N_1150,N_2032);
nor U9997 (N_9997,N_4009,N_124);
xor U9998 (N_9998,N_4480,N_4648);
or U9999 (N_9999,N_6185,N_2327);
xnor U10000 (N_10000,N_2732,N_3190);
and U10001 (N_10001,N_441,N_1011);
nor U10002 (N_10002,N_6101,N_3615);
and U10003 (N_10003,N_2197,N_1711);
or U10004 (N_10004,N_5917,N_736);
and U10005 (N_10005,N_1690,N_1901);
xor U10006 (N_10006,N_1695,N_3418);
xnor U10007 (N_10007,N_3730,N_3124);
and U10008 (N_10008,N_4782,N_833);
nor U10009 (N_10009,N_2661,N_2129);
or U10010 (N_10010,N_3182,N_1338);
nand U10011 (N_10011,N_581,N_1291);
nor U10012 (N_10012,N_3618,N_1554);
nor U10013 (N_10013,N_1985,N_4818);
and U10014 (N_10014,N_1402,N_4484);
and U10015 (N_10015,N_3021,N_5742);
nand U10016 (N_10016,N_2694,N_1330);
and U10017 (N_10017,N_3011,N_274);
nand U10018 (N_10018,N_708,N_2480);
nand U10019 (N_10019,N_5370,N_1046);
xor U10020 (N_10020,N_2437,N_4279);
xnor U10021 (N_10021,N_5962,N_4168);
nor U10022 (N_10022,N_5614,N_3067);
nand U10023 (N_10023,N_4812,N_3863);
nor U10024 (N_10024,N_3906,N_2825);
nor U10025 (N_10025,N_3740,N_5401);
or U10026 (N_10026,N_1743,N_399);
or U10027 (N_10027,N_4236,N_5114);
or U10028 (N_10028,N_979,N_5076);
or U10029 (N_10029,N_4938,N_1101);
or U10030 (N_10030,N_4571,N_2863);
and U10031 (N_10031,N_1148,N_2896);
or U10032 (N_10032,N_1958,N_83);
nand U10033 (N_10033,N_1454,N_1562);
nor U10034 (N_10034,N_2171,N_555);
xor U10035 (N_10035,N_889,N_3462);
and U10036 (N_10036,N_4999,N_4493);
nand U10037 (N_10037,N_3903,N_4406);
nand U10038 (N_10038,N_2287,N_3521);
nand U10039 (N_10039,N_4347,N_552);
xor U10040 (N_10040,N_287,N_694);
nand U10041 (N_10041,N_4211,N_1622);
or U10042 (N_10042,N_1227,N_1031);
xnor U10043 (N_10043,N_2725,N_579);
and U10044 (N_10044,N_1207,N_845);
nand U10045 (N_10045,N_1105,N_6046);
nor U10046 (N_10046,N_6233,N_636);
nand U10047 (N_10047,N_958,N_5694);
and U10048 (N_10048,N_2454,N_2483);
xor U10049 (N_10049,N_1611,N_2217);
or U10050 (N_10050,N_3189,N_1001);
and U10051 (N_10051,N_1090,N_5317);
and U10052 (N_10052,N_791,N_1840);
or U10053 (N_10053,N_3980,N_3105);
and U10054 (N_10054,N_4250,N_854);
and U10055 (N_10055,N_2922,N_39);
nand U10056 (N_10056,N_1258,N_3855);
nand U10057 (N_10057,N_239,N_153);
and U10058 (N_10058,N_5221,N_5104);
and U10059 (N_10059,N_189,N_3663);
or U10060 (N_10060,N_2375,N_5621);
and U10061 (N_10061,N_5669,N_5283);
nand U10062 (N_10062,N_284,N_4096);
and U10063 (N_10063,N_3376,N_3080);
nand U10064 (N_10064,N_5455,N_6245);
and U10065 (N_10065,N_4248,N_5138);
and U10066 (N_10066,N_1560,N_1873);
nand U10067 (N_10067,N_5480,N_4084);
xnor U10068 (N_10068,N_4963,N_4750);
nor U10069 (N_10069,N_3302,N_2968);
or U10070 (N_10070,N_2585,N_6230);
and U10071 (N_10071,N_4714,N_3049);
nand U10072 (N_10072,N_4025,N_3702);
or U10073 (N_10073,N_4355,N_5731);
nor U10074 (N_10074,N_1181,N_2372);
and U10075 (N_10075,N_4826,N_5885);
and U10076 (N_10076,N_3280,N_174);
or U10077 (N_10077,N_4922,N_1638);
and U10078 (N_10078,N_3299,N_3593);
nor U10079 (N_10079,N_136,N_1942);
nand U10080 (N_10080,N_2979,N_4884);
nor U10081 (N_10081,N_2727,N_5765);
xnor U10082 (N_10082,N_4643,N_5594);
or U10083 (N_10083,N_1884,N_3822);
and U10084 (N_10084,N_2922,N_4405);
nor U10085 (N_10085,N_1531,N_1934);
nor U10086 (N_10086,N_1339,N_3255);
and U10087 (N_10087,N_1612,N_5808);
or U10088 (N_10088,N_4254,N_6244);
xnor U10089 (N_10089,N_4135,N_5418);
and U10090 (N_10090,N_2428,N_4297);
nand U10091 (N_10091,N_4990,N_3385);
nand U10092 (N_10092,N_4111,N_4572);
nor U10093 (N_10093,N_5575,N_1803);
nand U10094 (N_10094,N_2928,N_3539);
or U10095 (N_10095,N_5773,N_3459);
nand U10096 (N_10096,N_1544,N_3542);
nor U10097 (N_10097,N_144,N_2630);
nor U10098 (N_10098,N_452,N_2817);
or U10099 (N_10099,N_2741,N_3401);
xnor U10100 (N_10100,N_2518,N_5001);
and U10101 (N_10101,N_6008,N_4097);
and U10102 (N_10102,N_672,N_1245);
nor U10103 (N_10103,N_2787,N_2617);
or U10104 (N_10104,N_720,N_4392);
and U10105 (N_10105,N_1040,N_4772);
nand U10106 (N_10106,N_3234,N_3164);
and U10107 (N_10107,N_1572,N_5227);
nand U10108 (N_10108,N_393,N_3924);
xor U10109 (N_10109,N_2000,N_537);
and U10110 (N_10110,N_5738,N_4369);
nor U10111 (N_10111,N_5622,N_2090);
nand U10112 (N_10112,N_2258,N_3350);
and U10113 (N_10113,N_526,N_5561);
or U10114 (N_10114,N_609,N_1438);
and U10115 (N_10115,N_1490,N_3118);
and U10116 (N_10116,N_6038,N_5344);
or U10117 (N_10117,N_4793,N_4627);
xor U10118 (N_10118,N_2400,N_6057);
xnor U10119 (N_10119,N_2573,N_5474);
and U10120 (N_10120,N_1942,N_2091);
xnor U10121 (N_10121,N_427,N_1371);
or U10122 (N_10122,N_4733,N_5439);
and U10123 (N_10123,N_3625,N_3825);
nand U10124 (N_10124,N_11,N_5051);
and U10125 (N_10125,N_2352,N_4115);
and U10126 (N_10126,N_3656,N_5291);
nand U10127 (N_10127,N_3800,N_5576);
or U10128 (N_10128,N_4002,N_2828);
nor U10129 (N_10129,N_3827,N_4570);
nor U10130 (N_10130,N_1529,N_2176);
and U10131 (N_10131,N_3820,N_1004);
and U10132 (N_10132,N_5552,N_3686);
xor U10133 (N_10133,N_2570,N_354);
nand U10134 (N_10134,N_3651,N_3869);
nor U10135 (N_10135,N_2318,N_3855);
nand U10136 (N_10136,N_3678,N_3617);
or U10137 (N_10137,N_1323,N_4545);
nor U10138 (N_10138,N_11,N_4160);
or U10139 (N_10139,N_1205,N_442);
nor U10140 (N_10140,N_144,N_3717);
and U10141 (N_10141,N_444,N_5364);
nand U10142 (N_10142,N_5358,N_4016);
or U10143 (N_10143,N_5456,N_6223);
nor U10144 (N_10144,N_3025,N_4655);
nor U10145 (N_10145,N_4680,N_841);
or U10146 (N_10146,N_2760,N_1445);
nor U10147 (N_10147,N_3256,N_972);
or U10148 (N_10148,N_3474,N_4064);
nor U10149 (N_10149,N_4661,N_489);
or U10150 (N_10150,N_3135,N_5219);
nand U10151 (N_10151,N_664,N_4812);
nor U10152 (N_10152,N_5594,N_4008);
and U10153 (N_10153,N_5691,N_5971);
or U10154 (N_10154,N_943,N_3883);
nand U10155 (N_10155,N_3827,N_1748);
or U10156 (N_10156,N_2155,N_2950);
or U10157 (N_10157,N_4597,N_3165);
nand U10158 (N_10158,N_2446,N_4033);
or U10159 (N_10159,N_702,N_2202);
nand U10160 (N_10160,N_4269,N_3681);
and U10161 (N_10161,N_2108,N_1388);
nor U10162 (N_10162,N_2547,N_5494);
nor U10163 (N_10163,N_1308,N_2158);
or U10164 (N_10164,N_2059,N_5488);
xnor U10165 (N_10165,N_2835,N_5219);
nand U10166 (N_10166,N_5437,N_1649);
or U10167 (N_10167,N_677,N_4004);
and U10168 (N_10168,N_2494,N_5014);
and U10169 (N_10169,N_2137,N_3303);
or U10170 (N_10170,N_5736,N_291);
nand U10171 (N_10171,N_2430,N_2268);
or U10172 (N_10172,N_2905,N_1161);
and U10173 (N_10173,N_2248,N_300);
and U10174 (N_10174,N_441,N_1884);
or U10175 (N_10175,N_4071,N_1270);
xnor U10176 (N_10176,N_3393,N_597);
nor U10177 (N_10177,N_4345,N_2556);
nor U10178 (N_10178,N_3058,N_864);
nor U10179 (N_10179,N_863,N_4565);
nand U10180 (N_10180,N_4023,N_5369);
and U10181 (N_10181,N_794,N_4894);
nand U10182 (N_10182,N_5946,N_1270);
nand U10183 (N_10183,N_2355,N_2263);
xor U10184 (N_10184,N_916,N_846);
nor U10185 (N_10185,N_3872,N_1567);
and U10186 (N_10186,N_1045,N_4637);
nor U10187 (N_10187,N_3852,N_4616);
xor U10188 (N_10188,N_1902,N_2785);
nand U10189 (N_10189,N_3298,N_1049);
nand U10190 (N_10190,N_698,N_5561);
nor U10191 (N_10191,N_2188,N_2346);
xor U10192 (N_10192,N_3179,N_6084);
and U10193 (N_10193,N_3520,N_4018);
nor U10194 (N_10194,N_5175,N_261);
or U10195 (N_10195,N_4646,N_353);
nor U10196 (N_10196,N_2186,N_2539);
nand U10197 (N_10197,N_2848,N_3871);
xnor U10198 (N_10198,N_1877,N_1776);
nor U10199 (N_10199,N_2097,N_4257);
nor U10200 (N_10200,N_1045,N_5337);
nand U10201 (N_10201,N_200,N_5421);
nand U10202 (N_10202,N_969,N_852);
nand U10203 (N_10203,N_2370,N_1731);
nor U10204 (N_10204,N_5087,N_3562);
or U10205 (N_10205,N_5889,N_2983);
or U10206 (N_10206,N_4622,N_584);
nand U10207 (N_10207,N_1618,N_5114);
nor U10208 (N_10208,N_5571,N_4423);
or U10209 (N_10209,N_2898,N_3474);
nor U10210 (N_10210,N_5613,N_3975);
xnor U10211 (N_10211,N_4193,N_5874);
xnor U10212 (N_10212,N_4485,N_5920);
or U10213 (N_10213,N_5385,N_1083);
xnor U10214 (N_10214,N_524,N_5461);
nor U10215 (N_10215,N_2858,N_4954);
and U10216 (N_10216,N_5167,N_5530);
nor U10217 (N_10217,N_3490,N_320);
nand U10218 (N_10218,N_801,N_2664);
nor U10219 (N_10219,N_3288,N_4542);
xnor U10220 (N_10220,N_6068,N_1834);
nand U10221 (N_10221,N_4239,N_1977);
and U10222 (N_10222,N_4097,N_5468);
nor U10223 (N_10223,N_3998,N_1495);
nor U10224 (N_10224,N_6206,N_511);
nor U10225 (N_10225,N_2922,N_1006);
and U10226 (N_10226,N_4865,N_286);
and U10227 (N_10227,N_366,N_2878);
nand U10228 (N_10228,N_2441,N_3438);
and U10229 (N_10229,N_5292,N_717);
and U10230 (N_10230,N_459,N_2548);
or U10231 (N_10231,N_3056,N_5466);
and U10232 (N_10232,N_3041,N_1474);
nor U10233 (N_10233,N_1276,N_6116);
and U10234 (N_10234,N_1256,N_5688);
xor U10235 (N_10235,N_4613,N_1944);
or U10236 (N_10236,N_51,N_545);
and U10237 (N_10237,N_2634,N_5715);
xor U10238 (N_10238,N_4485,N_4521);
and U10239 (N_10239,N_3470,N_429);
and U10240 (N_10240,N_3055,N_3735);
nand U10241 (N_10241,N_1009,N_3265);
nor U10242 (N_10242,N_5131,N_3930);
and U10243 (N_10243,N_5120,N_411);
nor U10244 (N_10244,N_4924,N_2672);
nor U10245 (N_10245,N_6068,N_5555);
nor U10246 (N_10246,N_2813,N_3825);
or U10247 (N_10247,N_1609,N_5799);
and U10248 (N_10248,N_2540,N_527);
or U10249 (N_10249,N_5480,N_578);
nand U10250 (N_10250,N_834,N_2278);
and U10251 (N_10251,N_1342,N_5817);
and U10252 (N_10252,N_5277,N_1096);
or U10253 (N_10253,N_2219,N_2447);
nor U10254 (N_10254,N_4118,N_2849);
xnor U10255 (N_10255,N_2837,N_5218);
xor U10256 (N_10256,N_2691,N_852);
and U10257 (N_10257,N_4798,N_2234);
nor U10258 (N_10258,N_2389,N_311);
xor U10259 (N_10259,N_5457,N_437);
nor U10260 (N_10260,N_1671,N_1372);
or U10261 (N_10261,N_1131,N_3860);
nor U10262 (N_10262,N_2424,N_2665);
or U10263 (N_10263,N_2251,N_1020);
xor U10264 (N_10264,N_5856,N_4273);
nor U10265 (N_10265,N_4543,N_2235);
xor U10266 (N_10266,N_797,N_5055);
or U10267 (N_10267,N_2351,N_5740);
xor U10268 (N_10268,N_4762,N_633);
and U10269 (N_10269,N_5881,N_1255);
nor U10270 (N_10270,N_5793,N_5806);
nor U10271 (N_10271,N_603,N_227);
xnor U10272 (N_10272,N_3017,N_3574);
and U10273 (N_10273,N_5045,N_1886);
or U10274 (N_10274,N_2528,N_3631);
nand U10275 (N_10275,N_4460,N_1831);
nand U10276 (N_10276,N_5358,N_434);
or U10277 (N_10277,N_1653,N_5130);
or U10278 (N_10278,N_2326,N_3353);
nor U10279 (N_10279,N_5466,N_4468);
or U10280 (N_10280,N_3319,N_1758);
nand U10281 (N_10281,N_1616,N_33);
and U10282 (N_10282,N_3128,N_2825);
nand U10283 (N_10283,N_4906,N_5503);
nand U10284 (N_10284,N_5116,N_917);
and U10285 (N_10285,N_3000,N_4122);
nand U10286 (N_10286,N_1116,N_3588);
nor U10287 (N_10287,N_3328,N_814);
xor U10288 (N_10288,N_1323,N_4886);
nand U10289 (N_10289,N_2105,N_3650);
or U10290 (N_10290,N_6127,N_2840);
xnor U10291 (N_10291,N_1577,N_3344);
and U10292 (N_10292,N_2089,N_4455);
nor U10293 (N_10293,N_648,N_4138);
nor U10294 (N_10294,N_1530,N_2214);
xnor U10295 (N_10295,N_3483,N_155);
nor U10296 (N_10296,N_2597,N_2811);
and U10297 (N_10297,N_611,N_3736);
nor U10298 (N_10298,N_4580,N_5461);
and U10299 (N_10299,N_441,N_598);
or U10300 (N_10300,N_814,N_2770);
nor U10301 (N_10301,N_330,N_3825);
nand U10302 (N_10302,N_4197,N_5459);
and U10303 (N_10303,N_931,N_6057);
and U10304 (N_10304,N_4193,N_4272);
nor U10305 (N_10305,N_1167,N_1180);
nand U10306 (N_10306,N_1696,N_5848);
nand U10307 (N_10307,N_330,N_380);
and U10308 (N_10308,N_443,N_3549);
and U10309 (N_10309,N_1061,N_4369);
or U10310 (N_10310,N_1019,N_266);
and U10311 (N_10311,N_1935,N_1168);
or U10312 (N_10312,N_3954,N_4253);
or U10313 (N_10313,N_5022,N_3615);
nor U10314 (N_10314,N_4098,N_5073);
or U10315 (N_10315,N_1365,N_5822);
or U10316 (N_10316,N_5076,N_2674);
nor U10317 (N_10317,N_2881,N_3063);
or U10318 (N_10318,N_5287,N_5917);
nand U10319 (N_10319,N_327,N_5413);
and U10320 (N_10320,N_5710,N_508);
or U10321 (N_10321,N_2909,N_2697);
or U10322 (N_10322,N_204,N_3351);
xor U10323 (N_10323,N_6084,N_741);
or U10324 (N_10324,N_4167,N_5610);
nand U10325 (N_10325,N_2237,N_1802);
or U10326 (N_10326,N_5500,N_4666);
and U10327 (N_10327,N_5504,N_2694);
and U10328 (N_10328,N_5069,N_610);
nor U10329 (N_10329,N_3881,N_3326);
nor U10330 (N_10330,N_4783,N_1669);
nor U10331 (N_10331,N_5582,N_5361);
nand U10332 (N_10332,N_2375,N_3421);
xor U10333 (N_10333,N_5361,N_293);
or U10334 (N_10334,N_3967,N_569);
nand U10335 (N_10335,N_3401,N_4540);
xnor U10336 (N_10336,N_932,N_4228);
and U10337 (N_10337,N_4412,N_3601);
and U10338 (N_10338,N_1169,N_2562);
nand U10339 (N_10339,N_1304,N_4762);
nor U10340 (N_10340,N_203,N_1158);
nor U10341 (N_10341,N_5562,N_5520);
xor U10342 (N_10342,N_4211,N_38);
and U10343 (N_10343,N_4125,N_5128);
xnor U10344 (N_10344,N_5902,N_3524);
nand U10345 (N_10345,N_5846,N_3082);
nor U10346 (N_10346,N_3345,N_3191);
nand U10347 (N_10347,N_5799,N_1619);
and U10348 (N_10348,N_4371,N_2500);
nor U10349 (N_10349,N_197,N_581);
nand U10350 (N_10350,N_595,N_3386);
or U10351 (N_10351,N_1033,N_3603);
or U10352 (N_10352,N_3144,N_5293);
or U10353 (N_10353,N_1551,N_2106);
nand U10354 (N_10354,N_104,N_981);
nor U10355 (N_10355,N_2905,N_4024);
nand U10356 (N_10356,N_5951,N_1724);
or U10357 (N_10357,N_395,N_702);
nand U10358 (N_10358,N_1076,N_3410);
nor U10359 (N_10359,N_551,N_1936);
or U10360 (N_10360,N_5572,N_5868);
and U10361 (N_10361,N_5140,N_491);
nor U10362 (N_10362,N_3910,N_3544);
xnor U10363 (N_10363,N_695,N_3571);
and U10364 (N_10364,N_2986,N_584);
and U10365 (N_10365,N_5294,N_4524);
or U10366 (N_10366,N_2938,N_5330);
nor U10367 (N_10367,N_1073,N_2659);
nand U10368 (N_10368,N_2818,N_1013);
nor U10369 (N_10369,N_1749,N_2982);
nor U10370 (N_10370,N_2793,N_4668);
or U10371 (N_10371,N_6076,N_157);
and U10372 (N_10372,N_2121,N_2850);
and U10373 (N_10373,N_2971,N_300);
and U10374 (N_10374,N_2240,N_5749);
and U10375 (N_10375,N_893,N_2908);
xor U10376 (N_10376,N_265,N_3092);
nor U10377 (N_10377,N_4731,N_5633);
or U10378 (N_10378,N_5110,N_5780);
or U10379 (N_10379,N_4671,N_1429);
or U10380 (N_10380,N_2169,N_4660);
or U10381 (N_10381,N_3325,N_3468);
nand U10382 (N_10382,N_3945,N_864);
and U10383 (N_10383,N_1459,N_2479);
or U10384 (N_10384,N_4700,N_5447);
nand U10385 (N_10385,N_5380,N_5341);
nor U10386 (N_10386,N_251,N_1550);
and U10387 (N_10387,N_5751,N_4711);
nor U10388 (N_10388,N_5475,N_447);
xnor U10389 (N_10389,N_3816,N_5087);
or U10390 (N_10390,N_193,N_1262);
nor U10391 (N_10391,N_4315,N_4377);
nand U10392 (N_10392,N_5572,N_4301);
nand U10393 (N_10393,N_3518,N_5094);
nand U10394 (N_10394,N_2112,N_2616);
nor U10395 (N_10395,N_2665,N_1502);
nor U10396 (N_10396,N_3780,N_1965);
and U10397 (N_10397,N_4235,N_283);
xnor U10398 (N_10398,N_1320,N_4138);
nand U10399 (N_10399,N_5167,N_1950);
xnor U10400 (N_10400,N_1003,N_5989);
or U10401 (N_10401,N_2904,N_2580);
nand U10402 (N_10402,N_4222,N_4876);
nand U10403 (N_10403,N_3093,N_2053);
and U10404 (N_10404,N_5391,N_464);
nor U10405 (N_10405,N_4289,N_5391);
nor U10406 (N_10406,N_1888,N_3962);
nand U10407 (N_10407,N_1345,N_362);
nor U10408 (N_10408,N_4749,N_3450);
and U10409 (N_10409,N_2488,N_1890);
nand U10410 (N_10410,N_6033,N_3490);
or U10411 (N_10411,N_5238,N_3681);
or U10412 (N_10412,N_541,N_2527);
and U10413 (N_10413,N_4681,N_1925);
nor U10414 (N_10414,N_4304,N_1918);
nand U10415 (N_10415,N_1784,N_1564);
nand U10416 (N_10416,N_4144,N_5199);
nand U10417 (N_10417,N_3631,N_2292);
or U10418 (N_10418,N_342,N_2015);
nand U10419 (N_10419,N_6045,N_3203);
nor U10420 (N_10420,N_4065,N_4267);
nor U10421 (N_10421,N_1188,N_555);
and U10422 (N_10422,N_2498,N_3814);
and U10423 (N_10423,N_1874,N_415);
nor U10424 (N_10424,N_5302,N_3112);
or U10425 (N_10425,N_1520,N_4572);
and U10426 (N_10426,N_5390,N_5735);
or U10427 (N_10427,N_759,N_4992);
nor U10428 (N_10428,N_4740,N_3827);
or U10429 (N_10429,N_6225,N_1326);
nor U10430 (N_10430,N_2285,N_3107);
or U10431 (N_10431,N_825,N_4099);
and U10432 (N_10432,N_5086,N_2283);
nor U10433 (N_10433,N_1874,N_142);
and U10434 (N_10434,N_500,N_3289);
and U10435 (N_10435,N_764,N_1155);
and U10436 (N_10436,N_2080,N_2132);
and U10437 (N_10437,N_4215,N_6072);
xnor U10438 (N_10438,N_1419,N_2746);
nand U10439 (N_10439,N_2766,N_5067);
or U10440 (N_10440,N_2042,N_4288);
or U10441 (N_10441,N_6128,N_3666);
and U10442 (N_10442,N_4918,N_5612);
or U10443 (N_10443,N_4550,N_489);
nand U10444 (N_10444,N_155,N_1366);
nand U10445 (N_10445,N_3968,N_2038);
and U10446 (N_10446,N_3415,N_3657);
nor U10447 (N_10447,N_4039,N_2233);
or U10448 (N_10448,N_1284,N_4593);
or U10449 (N_10449,N_6039,N_4476);
nor U10450 (N_10450,N_1031,N_3725);
nand U10451 (N_10451,N_4659,N_874);
and U10452 (N_10452,N_5675,N_3906);
and U10453 (N_10453,N_2764,N_2530);
or U10454 (N_10454,N_601,N_6079);
xnor U10455 (N_10455,N_1551,N_1939);
xnor U10456 (N_10456,N_3249,N_4913);
nand U10457 (N_10457,N_3509,N_3913);
nor U10458 (N_10458,N_4038,N_4567);
nand U10459 (N_10459,N_1679,N_2185);
xnor U10460 (N_10460,N_1091,N_4095);
nand U10461 (N_10461,N_3729,N_5064);
and U10462 (N_10462,N_5678,N_4616);
nand U10463 (N_10463,N_1286,N_3338);
or U10464 (N_10464,N_924,N_1798);
and U10465 (N_10465,N_1451,N_4000);
or U10466 (N_10466,N_4146,N_2849);
nand U10467 (N_10467,N_466,N_4364);
and U10468 (N_10468,N_1394,N_3145);
and U10469 (N_10469,N_3015,N_1280);
and U10470 (N_10470,N_3794,N_1048);
nand U10471 (N_10471,N_1541,N_5642);
nor U10472 (N_10472,N_954,N_4517);
or U10473 (N_10473,N_2723,N_4630);
or U10474 (N_10474,N_5805,N_4388);
xnor U10475 (N_10475,N_1732,N_5834);
nand U10476 (N_10476,N_3313,N_4662);
xnor U10477 (N_10477,N_264,N_688);
nand U10478 (N_10478,N_5543,N_4622);
nor U10479 (N_10479,N_1875,N_5193);
or U10480 (N_10480,N_2888,N_119);
or U10481 (N_10481,N_3349,N_4194);
or U10482 (N_10482,N_1668,N_6057);
or U10483 (N_10483,N_1868,N_253);
nor U10484 (N_10484,N_3957,N_5752);
and U10485 (N_10485,N_327,N_3650);
and U10486 (N_10486,N_40,N_4563);
and U10487 (N_10487,N_3555,N_4636);
nor U10488 (N_10488,N_1860,N_1134);
or U10489 (N_10489,N_2549,N_902);
xor U10490 (N_10490,N_4434,N_5112);
xor U10491 (N_10491,N_2145,N_6109);
or U10492 (N_10492,N_2966,N_905);
or U10493 (N_10493,N_153,N_5986);
nand U10494 (N_10494,N_920,N_1604);
and U10495 (N_10495,N_3090,N_4786);
and U10496 (N_10496,N_3735,N_795);
and U10497 (N_10497,N_5367,N_6141);
nor U10498 (N_10498,N_2810,N_1401);
or U10499 (N_10499,N_2559,N_3608);
and U10500 (N_10500,N_1203,N_3971);
nor U10501 (N_10501,N_1703,N_6063);
nand U10502 (N_10502,N_780,N_2385);
or U10503 (N_10503,N_1090,N_2575);
nor U10504 (N_10504,N_5155,N_3823);
and U10505 (N_10505,N_1985,N_1121);
nand U10506 (N_10506,N_1915,N_5502);
xnor U10507 (N_10507,N_3838,N_5872);
or U10508 (N_10508,N_406,N_1055);
xor U10509 (N_10509,N_5692,N_2833);
and U10510 (N_10510,N_611,N_389);
or U10511 (N_10511,N_5480,N_2482);
and U10512 (N_10512,N_66,N_1512);
or U10513 (N_10513,N_2659,N_6220);
or U10514 (N_10514,N_6216,N_2130);
and U10515 (N_10515,N_943,N_286);
nand U10516 (N_10516,N_5483,N_883);
nor U10517 (N_10517,N_1672,N_5334);
and U10518 (N_10518,N_5404,N_5849);
nand U10519 (N_10519,N_979,N_363);
and U10520 (N_10520,N_2418,N_5453);
xor U10521 (N_10521,N_4380,N_4206);
nor U10522 (N_10522,N_3642,N_444);
nand U10523 (N_10523,N_5339,N_6218);
nor U10524 (N_10524,N_3954,N_5804);
or U10525 (N_10525,N_5280,N_4734);
nor U10526 (N_10526,N_1391,N_872);
or U10527 (N_10527,N_1281,N_4186);
and U10528 (N_10528,N_1551,N_3511);
nand U10529 (N_10529,N_3470,N_3456);
xor U10530 (N_10530,N_1833,N_3469);
and U10531 (N_10531,N_1276,N_2559);
xor U10532 (N_10532,N_3140,N_1861);
and U10533 (N_10533,N_3770,N_5154);
nand U10534 (N_10534,N_139,N_795);
nand U10535 (N_10535,N_37,N_2060);
and U10536 (N_10536,N_2825,N_2911);
nand U10537 (N_10537,N_4602,N_678);
or U10538 (N_10538,N_1324,N_4708);
or U10539 (N_10539,N_5296,N_4447);
or U10540 (N_10540,N_5365,N_3114);
or U10541 (N_10541,N_882,N_389);
and U10542 (N_10542,N_5387,N_1443);
nor U10543 (N_10543,N_6110,N_352);
nor U10544 (N_10544,N_119,N_1565);
nand U10545 (N_10545,N_986,N_3974);
xnor U10546 (N_10546,N_202,N_1155);
and U10547 (N_10547,N_4615,N_135);
and U10548 (N_10548,N_4631,N_1048);
nor U10549 (N_10549,N_2812,N_6033);
or U10550 (N_10550,N_4874,N_2385);
nand U10551 (N_10551,N_2604,N_3472);
and U10552 (N_10552,N_5090,N_671);
nor U10553 (N_10553,N_3025,N_6040);
and U10554 (N_10554,N_4989,N_1610);
and U10555 (N_10555,N_2958,N_867);
nand U10556 (N_10556,N_4652,N_3132);
nor U10557 (N_10557,N_490,N_5066);
nand U10558 (N_10558,N_1141,N_4783);
and U10559 (N_10559,N_3146,N_5053);
or U10560 (N_10560,N_4386,N_5631);
xor U10561 (N_10561,N_790,N_4380);
or U10562 (N_10562,N_5611,N_3516);
nand U10563 (N_10563,N_618,N_447);
or U10564 (N_10564,N_3741,N_513);
or U10565 (N_10565,N_5955,N_5780);
nand U10566 (N_10566,N_1156,N_1836);
and U10567 (N_10567,N_4503,N_4680);
nand U10568 (N_10568,N_4280,N_6236);
and U10569 (N_10569,N_3159,N_2575);
nor U10570 (N_10570,N_3265,N_2639);
nor U10571 (N_10571,N_4182,N_1196);
and U10572 (N_10572,N_2551,N_690);
nand U10573 (N_10573,N_2739,N_5617);
nand U10574 (N_10574,N_6189,N_13);
xnor U10575 (N_10575,N_1910,N_4048);
and U10576 (N_10576,N_5683,N_3042);
nand U10577 (N_10577,N_822,N_1081);
and U10578 (N_10578,N_581,N_1419);
nor U10579 (N_10579,N_2753,N_2030);
nand U10580 (N_10580,N_4362,N_3139);
or U10581 (N_10581,N_1441,N_585);
or U10582 (N_10582,N_3872,N_2997);
and U10583 (N_10583,N_5962,N_1061);
nor U10584 (N_10584,N_3189,N_3104);
or U10585 (N_10585,N_4830,N_1894);
nor U10586 (N_10586,N_2276,N_4065);
nor U10587 (N_10587,N_469,N_2798);
nand U10588 (N_10588,N_4284,N_2502);
or U10589 (N_10589,N_768,N_194);
or U10590 (N_10590,N_3411,N_1158);
and U10591 (N_10591,N_5134,N_5895);
and U10592 (N_10592,N_3389,N_3319);
or U10593 (N_10593,N_2994,N_3556);
nor U10594 (N_10594,N_432,N_3119);
xor U10595 (N_10595,N_2864,N_5411);
nor U10596 (N_10596,N_310,N_519);
and U10597 (N_10597,N_5724,N_1974);
and U10598 (N_10598,N_3960,N_5740);
nand U10599 (N_10599,N_1856,N_2818);
nor U10600 (N_10600,N_645,N_3595);
or U10601 (N_10601,N_545,N_5051);
and U10602 (N_10602,N_2177,N_4298);
and U10603 (N_10603,N_90,N_5436);
and U10604 (N_10604,N_966,N_5406);
nor U10605 (N_10605,N_3273,N_1215);
xor U10606 (N_10606,N_1674,N_1912);
or U10607 (N_10607,N_2871,N_4442);
or U10608 (N_10608,N_2118,N_5261);
and U10609 (N_10609,N_5518,N_4284);
xnor U10610 (N_10610,N_989,N_5437);
and U10611 (N_10611,N_2997,N_5483);
nor U10612 (N_10612,N_353,N_746);
nand U10613 (N_10613,N_3685,N_3321);
nand U10614 (N_10614,N_2931,N_2430);
and U10615 (N_10615,N_5285,N_6017);
nand U10616 (N_10616,N_5287,N_2793);
or U10617 (N_10617,N_1846,N_1319);
nand U10618 (N_10618,N_3185,N_5304);
nand U10619 (N_10619,N_5154,N_5173);
and U10620 (N_10620,N_3401,N_2609);
nor U10621 (N_10621,N_4067,N_3754);
nand U10622 (N_10622,N_4256,N_1379);
nand U10623 (N_10623,N_2218,N_3577);
nand U10624 (N_10624,N_4789,N_5156);
and U10625 (N_10625,N_3965,N_1119);
nand U10626 (N_10626,N_4718,N_1361);
nor U10627 (N_10627,N_289,N_1842);
nor U10628 (N_10628,N_2595,N_3831);
nor U10629 (N_10629,N_4301,N_2290);
or U10630 (N_10630,N_1496,N_4678);
and U10631 (N_10631,N_6095,N_3920);
nand U10632 (N_10632,N_2178,N_2225);
xnor U10633 (N_10633,N_4216,N_5491);
nand U10634 (N_10634,N_5804,N_4094);
nand U10635 (N_10635,N_5474,N_5195);
nor U10636 (N_10636,N_5385,N_5407);
or U10637 (N_10637,N_4792,N_4093);
nand U10638 (N_10638,N_2423,N_4484);
and U10639 (N_10639,N_1126,N_2759);
and U10640 (N_10640,N_3784,N_1643);
or U10641 (N_10641,N_561,N_2604);
and U10642 (N_10642,N_4411,N_2662);
nor U10643 (N_10643,N_412,N_3300);
nand U10644 (N_10644,N_2199,N_165);
and U10645 (N_10645,N_1361,N_3524);
or U10646 (N_10646,N_1513,N_5586);
nor U10647 (N_10647,N_5179,N_3229);
and U10648 (N_10648,N_6016,N_5316);
nand U10649 (N_10649,N_996,N_1802);
and U10650 (N_10650,N_5747,N_2593);
nand U10651 (N_10651,N_5154,N_2507);
nand U10652 (N_10652,N_5450,N_3802);
nor U10653 (N_10653,N_3975,N_5246);
nand U10654 (N_10654,N_2715,N_379);
nand U10655 (N_10655,N_1953,N_1542);
nor U10656 (N_10656,N_5634,N_4309);
or U10657 (N_10657,N_3115,N_1521);
nor U10658 (N_10658,N_827,N_2741);
nor U10659 (N_10659,N_5834,N_2101);
nand U10660 (N_10660,N_1904,N_3851);
or U10661 (N_10661,N_2882,N_5404);
or U10662 (N_10662,N_2473,N_5597);
nand U10663 (N_10663,N_5067,N_1303);
and U10664 (N_10664,N_5774,N_610);
nor U10665 (N_10665,N_1855,N_5165);
nor U10666 (N_10666,N_1516,N_4562);
xor U10667 (N_10667,N_3588,N_3714);
xnor U10668 (N_10668,N_1501,N_3668);
or U10669 (N_10669,N_1531,N_5025);
nand U10670 (N_10670,N_1997,N_77);
nand U10671 (N_10671,N_4730,N_5358);
or U10672 (N_10672,N_4421,N_6050);
nor U10673 (N_10673,N_5806,N_3892);
and U10674 (N_10674,N_4206,N_5878);
and U10675 (N_10675,N_5821,N_2544);
nor U10676 (N_10676,N_2238,N_4826);
or U10677 (N_10677,N_4074,N_2635);
xnor U10678 (N_10678,N_978,N_4369);
or U10679 (N_10679,N_5305,N_3881);
xnor U10680 (N_10680,N_2800,N_6037);
and U10681 (N_10681,N_287,N_1508);
nand U10682 (N_10682,N_2680,N_4375);
xor U10683 (N_10683,N_919,N_2958);
and U10684 (N_10684,N_5790,N_4495);
nor U10685 (N_10685,N_3828,N_32);
nor U10686 (N_10686,N_3146,N_70);
nor U10687 (N_10687,N_2809,N_2243);
nor U10688 (N_10688,N_3568,N_5659);
or U10689 (N_10689,N_1445,N_1465);
or U10690 (N_10690,N_823,N_3274);
or U10691 (N_10691,N_6073,N_986);
xnor U10692 (N_10692,N_1924,N_5093);
or U10693 (N_10693,N_1937,N_3305);
nand U10694 (N_10694,N_3011,N_5545);
nor U10695 (N_10695,N_5094,N_422);
nand U10696 (N_10696,N_6056,N_2986);
nor U10697 (N_10697,N_4522,N_5096);
and U10698 (N_10698,N_3438,N_5108);
or U10699 (N_10699,N_5591,N_3211);
nand U10700 (N_10700,N_4770,N_3969);
xor U10701 (N_10701,N_3261,N_2496);
or U10702 (N_10702,N_3189,N_4320);
nand U10703 (N_10703,N_5201,N_4088);
or U10704 (N_10704,N_227,N_5334);
or U10705 (N_10705,N_5829,N_4555);
xnor U10706 (N_10706,N_3047,N_2829);
xor U10707 (N_10707,N_5286,N_3757);
or U10708 (N_10708,N_748,N_1636);
xnor U10709 (N_10709,N_2170,N_3314);
and U10710 (N_10710,N_1574,N_2755);
nor U10711 (N_10711,N_3965,N_102);
and U10712 (N_10712,N_4776,N_2890);
nor U10713 (N_10713,N_4152,N_1966);
and U10714 (N_10714,N_774,N_5851);
nor U10715 (N_10715,N_5317,N_4559);
and U10716 (N_10716,N_1368,N_3629);
or U10717 (N_10717,N_446,N_4006);
or U10718 (N_10718,N_235,N_3681);
nand U10719 (N_10719,N_5090,N_4338);
xor U10720 (N_10720,N_3247,N_5259);
and U10721 (N_10721,N_4486,N_191);
nand U10722 (N_10722,N_5508,N_5035);
and U10723 (N_10723,N_3634,N_2852);
and U10724 (N_10724,N_3806,N_1832);
nor U10725 (N_10725,N_6051,N_5024);
and U10726 (N_10726,N_3053,N_3593);
and U10727 (N_10727,N_5598,N_2355);
nor U10728 (N_10728,N_5850,N_5719);
and U10729 (N_10729,N_3307,N_579);
or U10730 (N_10730,N_664,N_2017);
nand U10731 (N_10731,N_5648,N_2174);
or U10732 (N_10732,N_3410,N_5360);
or U10733 (N_10733,N_1515,N_3671);
nand U10734 (N_10734,N_761,N_2352);
and U10735 (N_10735,N_4066,N_6209);
nor U10736 (N_10736,N_2647,N_5343);
nor U10737 (N_10737,N_2155,N_2449);
nand U10738 (N_10738,N_377,N_2079);
nand U10739 (N_10739,N_1715,N_3768);
and U10740 (N_10740,N_4327,N_3276);
nand U10741 (N_10741,N_6198,N_2849);
or U10742 (N_10742,N_1073,N_587);
nand U10743 (N_10743,N_5412,N_5441);
nand U10744 (N_10744,N_5209,N_3673);
and U10745 (N_10745,N_2018,N_6093);
nor U10746 (N_10746,N_4965,N_2106);
nor U10747 (N_10747,N_143,N_5493);
or U10748 (N_10748,N_3071,N_6130);
nand U10749 (N_10749,N_4485,N_3422);
or U10750 (N_10750,N_6132,N_1986);
nand U10751 (N_10751,N_4995,N_3631);
or U10752 (N_10752,N_6107,N_4607);
or U10753 (N_10753,N_5897,N_4217);
xnor U10754 (N_10754,N_5677,N_1548);
or U10755 (N_10755,N_4771,N_1611);
or U10756 (N_10756,N_4369,N_678);
or U10757 (N_10757,N_2391,N_1624);
nand U10758 (N_10758,N_2610,N_4538);
and U10759 (N_10759,N_2511,N_5485);
nand U10760 (N_10760,N_6160,N_5805);
nand U10761 (N_10761,N_2794,N_542);
or U10762 (N_10762,N_235,N_5242);
nand U10763 (N_10763,N_4790,N_4655);
nand U10764 (N_10764,N_5886,N_925);
or U10765 (N_10765,N_4031,N_1073);
nand U10766 (N_10766,N_953,N_4419);
nor U10767 (N_10767,N_4092,N_2334);
nor U10768 (N_10768,N_4157,N_646);
nor U10769 (N_10769,N_2505,N_816);
nor U10770 (N_10770,N_1577,N_5041);
nor U10771 (N_10771,N_1664,N_6103);
nor U10772 (N_10772,N_136,N_1116);
nand U10773 (N_10773,N_4519,N_5788);
nand U10774 (N_10774,N_4912,N_2806);
and U10775 (N_10775,N_2024,N_2601);
nand U10776 (N_10776,N_479,N_3415);
nand U10777 (N_10777,N_3143,N_2714);
or U10778 (N_10778,N_5003,N_3069);
or U10779 (N_10779,N_2515,N_5696);
xor U10780 (N_10780,N_4671,N_1697);
xnor U10781 (N_10781,N_4431,N_4221);
or U10782 (N_10782,N_4802,N_763);
or U10783 (N_10783,N_754,N_3751);
nor U10784 (N_10784,N_3193,N_4056);
nand U10785 (N_10785,N_2059,N_5428);
nor U10786 (N_10786,N_4970,N_153);
nor U10787 (N_10787,N_3968,N_1473);
and U10788 (N_10788,N_5860,N_737);
nand U10789 (N_10789,N_1818,N_4330);
and U10790 (N_10790,N_2455,N_4149);
nor U10791 (N_10791,N_1181,N_36);
nor U10792 (N_10792,N_1686,N_2287);
and U10793 (N_10793,N_2732,N_3295);
or U10794 (N_10794,N_4067,N_758);
and U10795 (N_10795,N_5205,N_2439);
xnor U10796 (N_10796,N_5213,N_1448);
nor U10797 (N_10797,N_944,N_3785);
nand U10798 (N_10798,N_6117,N_1202);
nand U10799 (N_10799,N_5240,N_4325);
and U10800 (N_10800,N_1729,N_5005);
or U10801 (N_10801,N_6012,N_1932);
or U10802 (N_10802,N_5144,N_3965);
and U10803 (N_10803,N_5146,N_1860);
nand U10804 (N_10804,N_5655,N_3397);
nor U10805 (N_10805,N_3210,N_2055);
or U10806 (N_10806,N_2995,N_5978);
or U10807 (N_10807,N_5705,N_4504);
or U10808 (N_10808,N_542,N_1303);
and U10809 (N_10809,N_195,N_5511);
nand U10810 (N_10810,N_2496,N_2105);
nor U10811 (N_10811,N_3097,N_2404);
nand U10812 (N_10812,N_2738,N_5170);
nand U10813 (N_10813,N_5459,N_5994);
xnor U10814 (N_10814,N_1781,N_4192);
or U10815 (N_10815,N_5310,N_3129);
nor U10816 (N_10816,N_5931,N_2348);
nand U10817 (N_10817,N_2760,N_3195);
xnor U10818 (N_10818,N_2299,N_5002);
nand U10819 (N_10819,N_2955,N_5658);
nand U10820 (N_10820,N_1332,N_4050);
nand U10821 (N_10821,N_5994,N_4614);
nor U10822 (N_10822,N_3057,N_1012);
xnor U10823 (N_10823,N_2497,N_1617);
or U10824 (N_10824,N_666,N_4505);
nand U10825 (N_10825,N_3745,N_3766);
nor U10826 (N_10826,N_5646,N_2252);
or U10827 (N_10827,N_1811,N_5626);
or U10828 (N_10828,N_2468,N_4836);
nor U10829 (N_10829,N_5453,N_438);
and U10830 (N_10830,N_4992,N_1290);
or U10831 (N_10831,N_4508,N_5758);
or U10832 (N_10832,N_4518,N_4360);
or U10833 (N_10833,N_2463,N_2536);
nand U10834 (N_10834,N_2257,N_4663);
and U10835 (N_10835,N_137,N_4215);
and U10836 (N_10836,N_4382,N_1443);
nor U10837 (N_10837,N_4218,N_2749);
nand U10838 (N_10838,N_3195,N_5468);
nor U10839 (N_10839,N_5996,N_4094);
or U10840 (N_10840,N_4777,N_312);
xor U10841 (N_10841,N_5820,N_5970);
or U10842 (N_10842,N_2815,N_713);
and U10843 (N_10843,N_4097,N_71);
and U10844 (N_10844,N_5297,N_2215);
nand U10845 (N_10845,N_368,N_5055);
xnor U10846 (N_10846,N_4973,N_1775);
or U10847 (N_10847,N_399,N_166);
xnor U10848 (N_10848,N_3302,N_79);
nand U10849 (N_10849,N_5754,N_4424);
nand U10850 (N_10850,N_5652,N_5531);
nor U10851 (N_10851,N_4423,N_6112);
nor U10852 (N_10852,N_1044,N_890);
nor U10853 (N_10853,N_514,N_4152);
nor U10854 (N_10854,N_1709,N_2632);
or U10855 (N_10855,N_3415,N_5612);
or U10856 (N_10856,N_2174,N_5784);
nor U10857 (N_10857,N_3637,N_3032);
and U10858 (N_10858,N_6006,N_5927);
or U10859 (N_10859,N_3874,N_2476);
nor U10860 (N_10860,N_5717,N_5937);
and U10861 (N_10861,N_195,N_3167);
xnor U10862 (N_10862,N_3879,N_2813);
nor U10863 (N_10863,N_29,N_468);
xnor U10864 (N_10864,N_2785,N_4929);
nand U10865 (N_10865,N_6207,N_5868);
or U10866 (N_10866,N_3666,N_4411);
nand U10867 (N_10867,N_2699,N_1168);
xor U10868 (N_10868,N_4455,N_272);
nand U10869 (N_10869,N_978,N_455);
xor U10870 (N_10870,N_1557,N_60);
nand U10871 (N_10871,N_4143,N_4412);
nand U10872 (N_10872,N_491,N_1953);
nand U10873 (N_10873,N_2414,N_5029);
and U10874 (N_10874,N_472,N_4532);
nand U10875 (N_10875,N_5456,N_4753);
xor U10876 (N_10876,N_157,N_4336);
xor U10877 (N_10877,N_4762,N_183);
nand U10878 (N_10878,N_3112,N_1090);
or U10879 (N_10879,N_3039,N_2210);
nand U10880 (N_10880,N_3373,N_4119);
and U10881 (N_10881,N_779,N_1389);
and U10882 (N_10882,N_5448,N_2091);
nor U10883 (N_10883,N_4705,N_3487);
xor U10884 (N_10884,N_5314,N_5041);
xnor U10885 (N_10885,N_387,N_2869);
nor U10886 (N_10886,N_3329,N_578);
nor U10887 (N_10887,N_5401,N_3526);
nor U10888 (N_10888,N_3656,N_2174);
and U10889 (N_10889,N_2442,N_5718);
nand U10890 (N_10890,N_4995,N_2909);
or U10891 (N_10891,N_1885,N_1864);
and U10892 (N_10892,N_5467,N_3342);
xnor U10893 (N_10893,N_6000,N_1733);
nand U10894 (N_10894,N_2910,N_2852);
nor U10895 (N_10895,N_3677,N_1029);
and U10896 (N_10896,N_3727,N_4523);
xnor U10897 (N_10897,N_121,N_3886);
and U10898 (N_10898,N_2108,N_3843);
nor U10899 (N_10899,N_5861,N_5220);
nor U10900 (N_10900,N_17,N_3186);
nor U10901 (N_10901,N_5490,N_3698);
nand U10902 (N_10902,N_179,N_6224);
nand U10903 (N_10903,N_1042,N_2546);
nand U10904 (N_10904,N_5253,N_6231);
xor U10905 (N_10905,N_293,N_4435);
or U10906 (N_10906,N_3904,N_5309);
and U10907 (N_10907,N_2149,N_2695);
nor U10908 (N_10908,N_1521,N_3910);
nor U10909 (N_10909,N_1534,N_935);
nor U10910 (N_10910,N_599,N_5689);
nor U10911 (N_10911,N_4632,N_2159);
nand U10912 (N_10912,N_5643,N_3414);
nand U10913 (N_10913,N_879,N_576);
nor U10914 (N_10914,N_2762,N_4868);
nor U10915 (N_10915,N_4789,N_3503);
and U10916 (N_10916,N_931,N_2232);
or U10917 (N_10917,N_691,N_1915);
and U10918 (N_10918,N_1351,N_3851);
or U10919 (N_10919,N_4936,N_5548);
nand U10920 (N_10920,N_5084,N_1182);
xor U10921 (N_10921,N_139,N_2762);
nand U10922 (N_10922,N_3365,N_3290);
nand U10923 (N_10923,N_2218,N_4625);
and U10924 (N_10924,N_2119,N_5758);
xnor U10925 (N_10925,N_441,N_1473);
nor U10926 (N_10926,N_2492,N_4663);
or U10927 (N_10927,N_5586,N_4601);
nor U10928 (N_10928,N_385,N_2277);
or U10929 (N_10929,N_977,N_70);
xnor U10930 (N_10930,N_4235,N_5401);
or U10931 (N_10931,N_5719,N_2685);
nor U10932 (N_10932,N_5888,N_5579);
xor U10933 (N_10933,N_935,N_4907);
and U10934 (N_10934,N_570,N_602);
xor U10935 (N_10935,N_205,N_117);
or U10936 (N_10936,N_6187,N_3933);
nand U10937 (N_10937,N_2721,N_1308);
nand U10938 (N_10938,N_2309,N_3326);
and U10939 (N_10939,N_789,N_4018);
xnor U10940 (N_10940,N_696,N_5226);
and U10941 (N_10941,N_3815,N_5315);
and U10942 (N_10942,N_4948,N_3648);
and U10943 (N_10943,N_1688,N_4147);
or U10944 (N_10944,N_5977,N_2772);
or U10945 (N_10945,N_832,N_3748);
xor U10946 (N_10946,N_4364,N_3173);
or U10947 (N_10947,N_3709,N_310);
or U10948 (N_10948,N_4864,N_4568);
nor U10949 (N_10949,N_5675,N_5458);
or U10950 (N_10950,N_4812,N_3535);
and U10951 (N_10951,N_5249,N_4221);
and U10952 (N_10952,N_1740,N_5000);
nand U10953 (N_10953,N_2380,N_3096);
nand U10954 (N_10954,N_3672,N_5883);
nand U10955 (N_10955,N_613,N_2345);
nor U10956 (N_10956,N_61,N_2533);
nor U10957 (N_10957,N_4794,N_349);
nor U10958 (N_10958,N_4433,N_1254);
xnor U10959 (N_10959,N_3168,N_1655);
and U10960 (N_10960,N_294,N_2343);
nand U10961 (N_10961,N_1875,N_5686);
or U10962 (N_10962,N_5913,N_570);
nand U10963 (N_10963,N_2908,N_3118);
or U10964 (N_10964,N_5526,N_109);
nor U10965 (N_10965,N_1749,N_2769);
xnor U10966 (N_10966,N_1016,N_2118);
nand U10967 (N_10967,N_2849,N_3818);
and U10968 (N_10968,N_405,N_3613);
nor U10969 (N_10969,N_3280,N_1130);
xor U10970 (N_10970,N_5505,N_4277);
nor U10971 (N_10971,N_964,N_328);
and U10972 (N_10972,N_6163,N_5429);
nor U10973 (N_10973,N_3050,N_2300);
nand U10974 (N_10974,N_5328,N_1263);
and U10975 (N_10975,N_282,N_1942);
nand U10976 (N_10976,N_1285,N_5783);
xnor U10977 (N_10977,N_3461,N_237);
nand U10978 (N_10978,N_2931,N_3283);
nand U10979 (N_10979,N_2583,N_4545);
nand U10980 (N_10980,N_773,N_690);
nor U10981 (N_10981,N_3767,N_1326);
and U10982 (N_10982,N_1698,N_3785);
xnor U10983 (N_10983,N_1594,N_4022);
or U10984 (N_10984,N_2215,N_832);
nor U10985 (N_10985,N_1111,N_4133);
nor U10986 (N_10986,N_831,N_4938);
nand U10987 (N_10987,N_1449,N_4299);
nor U10988 (N_10988,N_3942,N_6109);
xnor U10989 (N_10989,N_5708,N_1921);
nor U10990 (N_10990,N_5218,N_3317);
or U10991 (N_10991,N_3983,N_1157);
or U10992 (N_10992,N_3207,N_4860);
nor U10993 (N_10993,N_1981,N_4804);
xor U10994 (N_10994,N_4470,N_3614);
nand U10995 (N_10995,N_3788,N_3489);
and U10996 (N_10996,N_4846,N_5687);
xnor U10997 (N_10997,N_6164,N_4388);
and U10998 (N_10998,N_2483,N_157);
nand U10999 (N_10999,N_4467,N_6003);
and U11000 (N_11000,N_5803,N_2884);
xnor U11001 (N_11001,N_1434,N_1911);
nand U11002 (N_11002,N_2345,N_293);
nand U11003 (N_11003,N_2746,N_3562);
nor U11004 (N_11004,N_5930,N_1209);
nand U11005 (N_11005,N_5101,N_2307);
nor U11006 (N_11006,N_4201,N_5890);
nand U11007 (N_11007,N_264,N_80);
or U11008 (N_11008,N_4964,N_1947);
or U11009 (N_11009,N_2572,N_1143);
nor U11010 (N_11010,N_6177,N_5342);
xnor U11011 (N_11011,N_5915,N_3111);
xor U11012 (N_11012,N_2851,N_2329);
nand U11013 (N_11013,N_2893,N_1707);
nor U11014 (N_11014,N_5813,N_719);
and U11015 (N_11015,N_1438,N_2701);
nand U11016 (N_11016,N_5736,N_1324);
or U11017 (N_11017,N_2270,N_4430);
nand U11018 (N_11018,N_4075,N_1998);
or U11019 (N_11019,N_631,N_1689);
and U11020 (N_11020,N_289,N_641);
nor U11021 (N_11021,N_3622,N_2203);
and U11022 (N_11022,N_5451,N_1847);
and U11023 (N_11023,N_401,N_3424);
or U11024 (N_11024,N_1328,N_3094);
nand U11025 (N_11025,N_5548,N_468);
nor U11026 (N_11026,N_5462,N_3413);
or U11027 (N_11027,N_4119,N_5156);
and U11028 (N_11028,N_335,N_4491);
nor U11029 (N_11029,N_5199,N_3660);
and U11030 (N_11030,N_5285,N_4579);
nor U11031 (N_11031,N_1565,N_416);
and U11032 (N_11032,N_160,N_5755);
and U11033 (N_11033,N_1763,N_1900);
xor U11034 (N_11034,N_2649,N_238);
and U11035 (N_11035,N_4224,N_2082);
nor U11036 (N_11036,N_839,N_5863);
nand U11037 (N_11037,N_5936,N_2424);
nand U11038 (N_11038,N_858,N_4643);
or U11039 (N_11039,N_1895,N_3905);
and U11040 (N_11040,N_5049,N_4493);
or U11041 (N_11041,N_4752,N_405);
nor U11042 (N_11042,N_2440,N_4412);
and U11043 (N_11043,N_1556,N_5542);
or U11044 (N_11044,N_4576,N_2533);
or U11045 (N_11045,N_74,N_5656);
nor U11046 (N_11046,N_5491,N_1252);
nor U11047 (N_11047,N_2167,N_3841);
or U11048 (N_11048,N_1064,N_2942);
nand U11049 (N_11049,N_5060,N_4791);
nor U11050 (N_11050,N_5248,N_3628);
nor U11051 (N_11051,N_3757,N_3297);
nor U11052 (N_11052,N_5876,N_1402);
or U11053 (N_11053,N_482,N_1119);
nor U11054 (N_11054,N_3470,N_1911);
and U11055 (N_11055,N_2245,N_5784);
or U11056 (N_11056,N_5100,N_1939);
or U11057 (N_11057,N_2415,N_4536);
or U11058 (N_11058,N_3705,N_2447);
nand U11059 (N_11059,N_2746,N_5186);
nand U11060 (N_11060,N_2350,N_1416);
xnor U11061 (N_11061,N_5955,N_3135);
and U11062 (N_11062,N_1211,N_719);
and U11063 (N_11063,N_3404,N_5470);
xnor U11064 (N_11064,N_6205,N_2239);
and U11065 (N_11065,N_5855,N_45);
nor U11066 (N_11066,N_3479,N_2248);
xnor U11067 (N_11067,N_3331,N_3518);
or U11068 (N_11068,N_825,N_5337);
and U11069 (N_11069,N_1078,N_348);
nand U11070 (N_11070,N_5790,N_2304);
nand U11071 (N_11071,N_5040,N_480);
nand U11072 (N_11072,N_3517,N_4679);
nand U11073 (N_11073,N_3510,N_3646);
and U11074 (N_11074,N_1942,N_331);
nor U11075 (N_11075,N_3841,N_190);
and U11076 (N_11076,N_2624,N_5546);
nor U11077 (N_11077,N_1105,N_5632);
nand U11078 (N_11078,N_86,N_1114);
or U11079 (N_11079,N_189,N_5594);
xnor U11080 (N_11080,N_5607,N_4237);
and U11081 (N_11081,N_6049,N_512);
or U11082 (N_11082,N_737,N_1308);
or U11083 (N_11083,N_4868,N_3753);
or U11084 (N_11084,N_4061,N_3433);
and U11085 (N_11085,N_6195,N_5746);
nand U11086 (N_11086,N_3826,N_3227);
xnor U11087 (N_11087,N_2046,N_3808);
or U11088 (N_11088,N_1486,N_2684);
or U11089 (N_11089,N_1041,N_3054);
and U11090 (N_11090,N_876,N_1950);
nor U11091 (N_11091,N_2585,N_5593);
nor U11092 (N_11092,N_1625,N_4113);
nand U11093 (N_11093,N_1933,N_2416);
nor U11094 (N_11094,N_4854,N_2726);
or U11095 (N_11095,N_6032,N_5339);
or U11096 (N_11096,N_5349,N_4250);
or U11097 (N_11097,N_4622,N_2836);
nand U11098 (N_11098,N_4336,N_4739);
and U11099 (N_11099,N_5431,N_5622);
and U11100 (N_11100,N_5129,N_3988);
or U11101 (N_11101,N_4322,N_1746);
xor U11102 (N_11102,N_4205,N_1708);
xnor U11103 (N_11103,N_1161,N_3161);
nand U11104 (N_11104,N_592,N_889);
nand U11105 (N_11105,N_5369,N_1416);
or U11106 (N_11106,N_4919,N_5235);
nand U11107 (N_11107,N_157,N_2954);
and U11108 (N_11108,N_3218,N_39);
and U11109 (N_11109,N_1473,N_326);
or U11110 (N_11110,N_1560,N_4906);
xor U11111 (N_11111,N_2769,N_656);
xnor U11112 (N_11112,N_5526,N_4814);
and U11113 (N_11113,N_2067,N_2700);
and U11114 (N_11114,N_5535,N_1261);
xor U11115 (N_11115,N_4701,N_3032);
or U11116 (N_11116,N_1025,N_2123);
nand U11117 (N_11117,N_271,N_4148);
nor U11118 (N_11118,N_3999,N_2278);
or U11119 (N_11119,N_3367,N_2133);
nor U11120 (N_11120,N_675,N_849);
nand U11121 (N_11121,N_775,N_472);
xor U11122 (N_11122,N_4926,N_915);
nand U11123 (N_11123,N_4627,N_2536);
nor U11124 (N_11124,N_4631,N_323);
nand U11125 (N_11125,N_5061,N_2153);
nor U11126 (N_11126,N_4728,N_4319);
or U11127 (N_11127,N_5292,N_162);
and U11128 (N_11128,N_953,N_6038);
nor U11129 (N_11129,N_703,N_1755);
nor U11130 (N_11130,N_4794,N_4514);
nor U11131 (N_11131,N_2366,N_985);
and U11132 (N_11132,N_3103,N_2049);
nor U11133 (N_11133,N_5592,N_2448);
or U11134 (N_11134,N_204,N_3654);
nand U11135 (N_11135,N_3364,N_826);
and U11136 (N_11136,N_5677,N_1244);
or U11137 (N_11137,N_951,N_5813);
and U11138 (N_11138,N_2892,N_5624);
nor U11139 (N_11139,N_4931,N_4791);
or U11140 (N_11140,N_3234,N_2718);
nand U11141 (N_11141,N_1608,N_831);
and U11142 (N_11142,N_3024,N_5479);
or U11143 (N_11143,N_1245,N_4377);
nand U11144 (N_11144,N_1820,N_5920);
xor U11145 (N_11145,N_3816,N_3581);
nor U11146 (N_11146,N_917,N_2309);
nand U11147 (N_11147,N_1079,N_6094);
nor U11148 (N_11148,N_4446,N_4767);
nor U11149 (N_11149,N_5869,N_2698);
nand U11150 (N_11150,N_1741,N_4110);
nand U11151 (N_11151,N_1765,N_5643);
nor U11152 (N_11152,N_3661,N_214);
or U11153 (N_11153,N_4678,N_1287);
nor U11154 (N_11154,N_5492,N_1020);
or U11155 (N_11155,N_4767,N_1521);
or U11156 (N_11156,N_870,N_5902);
and U11157 (N_11157,N_2581,N_2184);
nand U11158 (N_11158,N_6118,N_1502);
nor U11159 (N_11159,N_799,N_5896);
or U11160 (N_11160,N_1571,N_2706);
xor U11161 (N_11161,N_317,N_5471);
nand U11162 (N_11162,N_3646,N_58);
nand U11163 (N_11163,N_346,N_2561);
or U11164 (N_11164,N_2433,N_4054);
or U11165 (N_11165,N_4033,N_4924);
and U11166 (N_11166,N_3594,N_2299);
nor U11167 (N_11167,N_1608,N_6084);
nor U11168 (N_11168,N_3324,N_2889);
and U11169 (N_11169,N_1686,N_3537);
and U11170 (N_11170,N_5878,N_2785);
xnor U11171 (N_11171,N_5419,N_1805);
nor U11172 (N_11172,N_5255,N_3152);
nand U11173 (N_11173,N_5496,N_4707);
or U11174 (N_11174,N_5262,N_4258);
nand U11175 (N_11175,N_3111,N_4775);
nor U11176 (N_11176,N_1538,N_5419);
or U11177 (N_11177,N_5851,N_2705);
or U11178 (N_11178,N_2754,N_2045);
and U11179 (N_11179,N_4659,N_5080);
and U11180 (N_11180,N_3627,N_513);
or U11181 (N_11181,N_1278,N_2346);
or U11182 (N_11182,N_664,N_1348);
nor U11183 (N_11183,N_1354,N_1547);
and U11184 (N_11184,N_663,N_340);
and U11185 (N_11185,N_2906,N_4615);
or U11186 (N_11186,N_5306,N_5194);
nand U11187 (N_11187,N_5821,N_4873);
xor U11188 (N_11188,N_990,N_1455);
nand U11189 (N_11189,N_4278,N_2081);
or U11190 (N_11190,N_6086,N_25);
or U11191 (N_11191,N_2266,N_4243);
or U11192 (N_11192,N_3933,N_5603);
nand U11193 (N_11193,N_3435,N_2876);
nor U11194 (N_11194,N_672,N_5349);
or U11195 (N_11195,N_6244,N_821);
nor U11196 (N_11196,N_6004,N_5227);
xor U11197 (N_11197,N_4948,N_3467);
nor U11198 (N_11198,N_5920,N_4300);
or U11199 (N_11199,N_4792,N_2481);
and U11200 (N_11200,N_1774,N_3443);
xor U11201 (N_11201,N_3908,N_1163);
and U11202 (N_11202,N_1309,N_1971);
nor U11203 (N_11203,N_2992,N_1352);
nand U11204 (N_11204,N_4736,N_2847);
nand U11205 (N_11205,N_2868,N_2541);
or U11206 (N_11206,N_1146,N_3192);
nor U11207 (N_11207,N_5939,N_5861);
nor U11208 (N_11208,N_4147,N_5710);
nor U11209 (N_11209,N_707,N_5400);
nor U11210 (N_11210,N_5074,N_6223);
xnor U11211 (N_11211,N_4933,N_2158);
and U11212 (N_11212,N_4377,N_2606);
nor U11213 (N_11213,N_5580,N_2120);
xor U11214 (N_11214,N_5138,N_5741);
or U11215 (N_11215,N_5969,N_4266);
nor U11216 (N_11216,N_4005,N_5411);
nand U11217 (N_11217,N_5398,N_2013);
nand U11218 (N_11218,N_3789,N_2747);
nor U11219 (N_11219,N_3384,N_546);
nand U11220 (N_11220,N_2681,N_659);
nor U11221 (N_11221,N_3186,N_191);
or U11222 (N_11222,N_4642,N_2014);
nor U11223 (N_11223,N_5558,N_77);
nor U11224 (N_11224,N_4126,N_1569);
nand U11225 (N_11225,N_2549,N_4822);
and U11226 (N_11226,N_1587,N_612);
and U11227 (N_11227,N_1289,N_5956);
or U11228 (N_11228,N_2793,N_588);
nor U11229 (N_11229,N_6092,N_1101);
xor U11230 (N_11230,N_2562,N_5063);
or U11231 (N_11231,N_5992,N_4066);
nor U11232 (N_11232,N_1681,N_5898);
and U11233 (N_11233,N_2727,N_2807);
or U11234 (N_11234,N_2140,N_2339);
nor U11235 (N_11235,N_4299,N_3869);
and U11236 (N_11236,N_4215,N_2529);
nand U11237 (N_11237,N_6061,N_4298);
or U11238 (N_11238,N_4969,N_2654);
or U11239 (N_11239,N_1088,N_2581);
nand U11240 (N_11240,N_2909,N_6193);
and U11241 (N_11241,N_326,N_4524);
nand U11242 (N_11242,N_2158,N_4280);
and U11243 (N_11243,N_2681,N_3385);
and U11244 (N_11244,N_2320,N_3577);
xnor U11245 (N_11245,N_4455,N_3103);
nand U11246 (N_11246,N_2895,N_1519);
or U11247 (N_11247,N_2212,N_5914);
or U11248 (N_11248,N_4568,N_1500);
and U11249 (N_11249,N_856,N_3798);
nor U11250 (N_11250,N_5658,N_566);
nand U11251 (N_11251,N_2961,N_1035);
nand U11252 (N_11252,N_3094,N_5167);
nor U11253 (N_11253,N_3626,N_3342);
xor U11254 (N_11254,N_4941,N_1133);
and U11255 (N_11255,N_5396,N_1221);
and U11256 (N_11256,N_2707,N_5371);
or U11257 (N_11257,N_2786,N_631);
and U11258 (N_11258,N_2037,N_3980);
and U11259 (N_11259,N_2655,N_1637);
nand U11260 (N_11260,N_600,N_2408);
nand U11261 (N_11261,N_3976,N_3861);
nand U11262 (N_11262,N_1828,N_965);
and U11263 (N_11263,N_2876,N_1648);
nand U11264 (N_11264,N_2425,N_1497);
and U11265 (N_11265,N_2144,N_2722);
and U11266 (N_11266,N_806,N_3503);
xor U11267 (N_11267,N_401,N_4990);
or U11268 (N_11268,N_4142,N_841);
and U11269 (N_11269,N_4840,N_4343);
nor U11270 (N_11270,N_3952,N_267);
and U11271 (N_11271,N_5518,N_4337);
or U11272 (N_11272,N_5610,N_3697);
nor U11273 (N_11273,N_126,N_2966);
nor U11274 (N_11274,N_2981,N_4451);
nor U11275 (N_11275,N_2350,N_2761);
nand U11276 (N_11276,N_4079,N_3537);
or U11277 (N_11277,N_632,N_2496);
and U11278 (N_11278,N_5756,N_4341);
or U11279 (N_11279,N_4629,N_2513);
nand U11280 (N_11280,N_4223,N_4467);
nor U11281 (N_11281,N_1913,N_5675);
or U11282 (N_11282,N_1659,N_4623);
and U11283 (N_11283,N_5309,N_1120);
nor U11284 (N_11284,N_5326,N_5291);
nand U11285 (N_11285,N_6008,N_5417);
and U11286 (N_11286,N_5475,N_2486);
nand U11287 (N_11287,N_831,N_4322);
nand U11288 (N_11288,N_3288,N_3964);
xor U11289 (N_11289,N_3594,N_5373);
and U11290 (N_11290,N_1777,N_5975);
or U11291 (N_11291,N_2332,N_5079);
nor U11292 (N_11292,N_502,N_4921);
and U11293 (N_11293,N_1437,N_100);
or U11294 (N_11294,N_4929,N_4367);
or U11295 (N_11295,N_1031,N_980);
nand U11296 (N_11296,N_3750,N_4703);
or U11297 (N_11297,N_839,N_3339);
nand U11298 (N_11298,N_362,N_4679);
nor U11299 (N_11299,N_3854,N_5538);
nand U11300 (N_11300,N_6000,N_3200);
nand U11301 (N_11301,N_1875,N_5432);
xnor U11302 (N_11302,N_2554,N_365);
nor U11303 (N_11303,N_1165,N_2467);
xnor U11304 (N_11304,N_3741,N_5420);
nor U11305 (N_11305,N_4656,N_3021);
nand U11306 (N_11306,N_2624,N_1116);
nand U11307 (N_11307,N_138,N_4782);
nor U11308 (N_11308,N_4657,N_870);
nand U11309 (N_11309,N_6208,N_4988);
or U11310 (N_11310,N_6193,N_3902);
and U11311 (N_11311,N_4389,N_6070);
nor U11312 (N_11312,N_1534,N_3247);
or U11313 (N_11313,N_5627,N_5887);
and U11314 (N_11314,N_4375,N_5139);
and U11315 (N_11315,N_3328,N_4755);
nor U11316 (N_11316,N_2036,N_2386);
nor U11317 (N_11317,N_5041,N_3006);
nor U11318 (N_11318,N_2093,N_5526);
and U11319 (N_11319,N_2762,N_2268);
xor U11320 (N_11320,N_3297,N_3652);
and U11321 (N_11321,N_5272,N_5222);
nand U11322 (N_11322,N_3822,N_2311);
or U11323 (N_11323,N_2492,N_3003);
and U11324 (N_11324,N_439,N_6238);
or U11325 (N_11325,N_6134,N_1321);
nand U11326 (N_11326,N_849,N_338);
nand U11327 (N_11327,N_2820,N_5323);
and U11328 (N_11328,N_1364,N_3133);
and U11329 (N_11329,N_3973,N_4168);
and U11330 (N_11330,N_1662,N_1401);
nor U11331 (N_11331,N_4288,N_2102);
nor U11332 (N_11332,N_5718,N_3854);
xnor U11333 (N_11333,N_2445,N_2321);
nand U11334 (N_11334,N_3697,N_248);
nor U11335 (N_11335,N_2821,N_2738);
xnor U11336 (N_11336,N_3841,N_2894);
xor U11337 (N_11337,N_4034,N_646);
nand U11338 (N_11338,N_6021,N_1423);
xnor U11339 (N_11339,N_1287,N_1058);
nor U11340 (N_11340,N_2482,N_5585);
nand U11341 (N_11341,N_2060,N_365);
nor U11342 (N_11342,N_5404,N_6121);
nor U11343 (N_11343,N_1133,N_3138);
and U11344 (N_11344,N_4551,N_959);
nor U11345 (N_11345,N_4960,N_4382);
xor U11346 (N_11346,N_5877,N_4187);
nor U11347 (N_11347,N_3601,N_5383);
xor U11348 (N_11348,N_1008,N_5407);
nor U11349 (N_11349,N_3260,N_678);
nor U11350 (N_11350,N_2836,N_1729);
nand U11351 (N_11351,N_3448,N_3855);
or U11352 (N_11352,N_4089,N_2719);
nor U11353 (N_11353,N_420,N_2079);
or U11354 (N_11354,N_176,N_3338);
nor U11355 (N_11355,N_3268,N_1382);
nor U11356 (N_11356,N_3672,N_3212);
nand U11357 (N_11357,N_4549,N_5273);
nor U11358 (N_11358,N_4968,N_4571);
nor U11359 (N_11359,N_1020,N_3104);
nor U11360 (N_11360,N_2077,N_3760);
nand U11361 (N_11361,N_5670,N_483);
and U11362 (N_11362,N_4428,N_2112);
nand U11363 (N_11363,N_570,N_1688);
nand U11364 (N_11364,N_5856,N_6152);
nand U11365 (N_11365,N_4322,N_3638);
and U11366 (N_11366,N_2424,N_2519);
nor U11367 (N_11367,N_4698,N_4165);
xnor U11368 (N_11368,N_4026,N_432);
nand U11369 (N_11369,N_6032,N_3692);
nand U11370 (N_11370,N_130,N_4842);
or U11371 (N_11371,N_4142,N_698);
xnor U11372 (N_11372,N_3851,N_277);
nor U11373 (N_11373,N_4281,N_825);
nor U11374 (N_11374,N_3612,N_1071);
and U11375 (N_11375,N_5319,N_4888);
nand U11376 (N_11376,N_3623,N_1825);
nand U11377 (N_11377,N_2927,N_5129);
nand U11378 (N_11378,N_3857,N_5078);
and U11379 (N_11379,N_2643,N_5674);
nand U11380 (N_11380,N_1967,N_5114);
nand U11381 (N_11381,N_3784,N_5959);
nor U11382 (N_11382,N_3003,N_5893);
and U11383 (N_11383,N_4890,N_2478);
nor U11384 (N_11384,N_5764,N_3616);
or U11385 (N_11385,N_2706,N_5487);
nand U11386 (N_11386,N_1534,N_3152);
nor U11387 (N_11387,N_5080,N_405);
nand U11388 (N_11388,N_1199,N_3269);
nand U11389 (N_11389,N_3893,N_4374);
nand U11390 (N_11390,N_3182,N_5828);
xor U11391 (N_11391,N_3535,N_3322);
nand U11392 (N_11392,N_5983,N_1839);
nand U11393 (N_11393,N_3983,N_1673);
or U11394 (N_11394,N_3388,N_6046);
or U11395 (N_11395,N_5815,N_44);
nand U11396 (N_11396,N_8,N_3641);
xnor U11397 (N_11397,N_5817,N_30);
nor U11398 (N_11398,N_4441,N_4724);
or U11399 (N_11399,N_2432,N_2525);
or U11400 (N_11400,N_4850,N_5821);
nor U11401 (N_11401,N_6195,N_6030);
nor U11402 (N_11402,N_2189,N_4630);
nor U11403 (N_11403,N_5226,N_1540);
and U11404 (N_11404,N_1943,N_5080);
and U11405 (N_11405,N_4054,N_4696);
nand U11406 (N_11406,N_4963,N_3449);
nand U11407 (N_11407,N_5879,N_4401);
nor U11408 (N_11408,N_4203,N_3093);
and U11409 (N_11409,N_5317,N_1057);
xor U11410 (N_11410,N_5735,N_4757);
nand U11411 (N_11411,N_314,N_5295);
or U11412 (N_11412,N_5708,N_1874);
and U11413 (N_11413,N_5663,N_5214);
xnor U11414 (N_11414,N_329,N_5133);
or U11415 (N_11415,N_5067,N_3764);
nor U11416 (N_11416,N_681,N_495);
nand U11417 (N_11417,N_4825,N_2260);
nand U11418 (N_11418,N_2462,N_3318);
nor U11419 (N_11419,N_2532,N_1914);
nand U11420 (N_11420,N_3668,N_1055);
nand U11421 (N_11421,N_5389,N_1936);
nand U11422 (N_11422,N_1978,N_3123);
or U11423 (N_11423,N_5227,N_2127);
nor U11424 (N_11424,N_1368,N_4833);
nor U11425 (N_11425,N_4330,N_5116);
xnor U11426 (N_11426,N_5106,N_2470);
nand U11427 (N_11427,N_4300,N_1492);
nand U11428 (N_11428,N_4061,N_5011);
and U11429 (N_11429,N_1762,N_4852);
and U11430 (N_11430,N_601,N_133);
and U11431 (N_11431,N_2451,N_1187);
xnor U11432 (N_11432,N_6161,N_1704);
xnor U11433 (N_11433,N_4512,N_5598);
and U11434 (N_11434,N_3183,N_3420);
nand U11435 (N_11435,N_3478,N_5948);
nor U11436 (N_11436,N_336,N_6149);
and U11437 (N_11437,N_2781,N_2382);
nand U11438 (N_11438,N_2098,N_5939);
nor U11439 (N_11439,N_4386,N_4503);
nor U11440 (N_11440,N_3877,N_4057);
and U11441 (N_11441,N_56,N_4104);
and U11442 (N_11442,N_4480,N_599);
xnor U11443 (N_11443,N_6055,N_755);
nor U11444 (N_11444,N_4091,N_258);
or U11445 (N_11445,N_2898,N_1230);
xor U11446 (N_11446,N_517,N_3637);
nor U11447 (N_11447,N_6107,N_2488);
nand U11448 (N_11448,N_5911,N_1090);
and U11449 (N_11449,N_4907,N_2616);
and U11450 (N_11450,N_4532,N_2556);
and U11451 (N_11451,N_2693,N_2703);
or U11452 (N_11452,N_62,N_839);
and U11453 (N_11453,N_614,N_4498);
or U11454 (N_11454,N_5789,N_2695);
nand U11455 (N_11455,N_3973,N_5049);
nand U11456 (N_11456,N_4217,N_2001);
nor U11457 (N_11457,N_6246,N_1691);
and U11458 (N_11458,N_319,N_5738);
or U11459 (N_11459,N_2406,N_4570);
xor U11460 (N_11460,N_2720,N_2200);
and U11461 (N_11461,N_2290,N_2708);
nand U11462 (N_11462,N_2320,N_4391);
nor U11463 (N_11463,N_4700,N_1967);
nand U11464 (N_11464,N_3428,N_5838);
and U11465 (N_11465,N_2663,N_182);
and U11466 (N_11466,N_1873,N_1828);
or U11467 (N_11467,N_3087,N_5446);
nand U11468 (N_11468,N_2158,N_855);
or U11469 (N_11469,N_1023,N_6112);
nand U11470 (N_11470,N_2078,N_727);
or U11471 (N_11471,N_5290,N_5157);
nor U11472 (N_11472,N_2764,N_309);
nor U11473 (N_11473,N_3493,N_5202);
nor U11474 (N_11474,N_5331,N_3161);
or U11475 (N_11475,N_229,N_5144);
nor U11476 (N_11476,N_5596,N_4927);
or U11477 (N_11477,N_5627,N_982);
nor U11478 (N_11478,N_3387,N_6063);
nor U11479 (N_11479,N_5726,N_2652);
xor U11480 (N_11480,N_5639,N_5541);
or U11481 (N_11481,N_5049,N_5293);
and U11482 (N_11482,N_1497,N_1973);
and U11483 (N_11483,N_2888,N_2523);
nor U11484 (N_11484,N_3784,N_4219);
nor U11485 (N_11485,N_3217,N_231);
or U11486 (N_11486,N_5966,N_1389);
or U11487 (N_11487,N_2362,N_5902);
nor U11488 (N_11488,N_3295,N_183);
or U11489 (N_11489,N_1017,N_466);
and U11490 (N_11490,N_1283,N_4589);
or U11491 (N_11491,N_59,N_128);
nand U11492 (N_11492,N_6194,N_119);
or U11493 (N_11493,N_283,N_2376);
xnor U11494 (N_11494,N_1959,N_725);
nor U11495 (N_11495,N_2284,N_106);
nor U11496 (N_11496,N_516,N_5860);
xor U11497 (N_11497,N_493,N_3083);
nand U11498 (N_11498,N_4158,N_164);
or U11499 (N_11499,N_3478,N_960);
and U11500 (N_11500,N_2099,N_1381);
and U11501 (N_11501,N_3575,N_1967);
nand U11502 (N_11502,N_1500,N_3417);
or U11503 (N_11503,N_4525,N_2744);
or U11504 (N_11504,N_3877,N_307);
or U11505 (N_11505,N_748,N_6044);
nand U11506 (N_11506,N_3634,N_1320);
nand U11507 (N_11507,N_850,N_3229);
and U11508 (N_11508,N_1300,N_3690);
and U11509 (N_11509,N_1946,N_3205);
or U11510 (N_11510,N_5659,N_3978);
nand U11511 (N_11511,N_1140,N_791);
and U11512 (N_11512,N_2433,N_3164);
and U11513 (N_11513,N_1716,N_6008);
and U11514 (N_11514,N_2384,N_63);
xnor U11515 (N_11515,N_5891,N_2457);
xor U11516 (N_11516,N_1940,N_3798);
and U11517 (N_11517,N_4457,N_789);
or U11518 (N_11518,N_3572,N_5824);
and U11519 (N_11519,N_592,N_2483);
or U11520 (N_11520,N_5536,N_5939);
nor U11521 (N_11521,N_350,N_665);
xor U11522 (N_11522,N_1370,N_5683);
nand U11523 (N_11523,N_558,N_2998);
and U11524 (N_11524,N_5391,N_6077);
and U11525 (N_11525,N_5180,N_1053);
or U11526 (N_11526,N_1618,N_1467);
nand U11527 (N_11527,N_897,N_4986);
or U11528 (N_11528,N_3277,N_2872);
nand U11529 (N_11529,N_370,N_2594);
and U11530 (N_11530,N_5916,N_2587);
and U11531 (N_11531,N_3016,N_5764);
nor U11532 (N_11532,N_1052,N_4061);
and U11533 (N_11533,N_345,N_6047);
and U11534 (N_11534,N_2744,N_260);
nand U11535 (N_11535,N_4731,N_4196);
nor U11536 (N_11536,N_3273,N_3735);
or U11537 (N_11537,N_2829,N_38);
and U11538 (N_11538,N_1263,N_2504);
xnor U11539 (N_11539,N_3779,N_11);
and U11540 (N_11540,N_1330,N_5186);
or U11541 (N_11541,N_4104,N_1969);
nand U11542 (N_11542,N_5242,N_6237);
nor U11543 (N_11543,N_2400,N_179);
and U11544 (N_11544,N_1291,N_6008);
and U11545 (N_11545,N_4896,N_2298);
nor U11546 (N_11546,N_5484,N_3285);
nand U11547 (N_11547,N_3145,N_2822);
nand U11548 (N_11548,N_2964,N_4829);
or U11549 (N_11549,N_1102,N_6150);
and U11550 (N_11550,N_4616,N_499);
or U11551 (N_11551,N_1980,N_565);
and U11552 (N_11552,N_2683,N_215);
xor U11553 (N_11553,N_4606,N_5515);
nor U11554 (N_11554,N_1322,N_4041);
or U11555 (N_11555,N_4864,N_4140);
or U11556 (N_11556,N_1877,N_5812);
xnor U11557 (N_11557,N_6113,N_6170);
or U11558 (N_11558,N_2461,N_2483);
or U11559 (N_11559,N_5301,N_3475);
nor U11560 (N_11560,N_4851,N_2660);
and U11561 (N_11561,N_4391,N_5552);
and U11562 (N_11562,N_5589,N_2786);
and U11563 (N_11563,N_4174,N_3999);
and U11564 (N_11564,N_5152,N_3556);
xor U11565 (N_11565,N_5523,N_5434);
nor U11566 (N_11566,N_3786,N_8);
or U11567 (N_11567,N_4313,N_3534);
and U11568 (N_11568,N_4167,N_5697);
nor U11569 (N_11569,N_2033,N_4960);
or U11570 (N_11570,N_3257,N_1041);
nor U11571 (N_11571,N_5406,N_5231);
and U11572 (N_11572,N_3774,N_3306);
nor U11573 (N_11573,N_4758,N_4348);
nand U11574 (N_11574,N_940,N_3149);
xor U11575 (N_11575,N_2959,N_2104);
nand U11576 (N_11576,N_468,N_1835);
and U11577 (N_11577,N_4494,N_3565);
or U11578 (N_11578,N_775,N_92);
nor U11579 (N_11579,N_6137,N_1871);
and U11580 (N_11580,N_2351,N_3565);
nor U11581 (N_11581,N_3256,N_2815);
or U11582 (N_11582,N_4709,N_1703);
nor U11583 (N_11583,N_148,N_2658);
nor U11584 (N_11584,N_4163,N_4365);
and U11585 (N_11585,N_2570,N_2489);
and U11586 (N_11586,N_5649,N_3345);
xor U11587 (N_11587,N_1666,N_6109);
xor U11588 (N_11588,N_5262,N_5986);
or U11589 (N_11589,N_5467,N_6042);
nand U11590 (N_11590,N_2557,N_3936);
nor U11591 (N_11591,N_4302,N_5817);
nor U11592 (N_11592,N_3937,N_1714);
nand U11593 (N_11593,N_134,N_3122);
or U11594 (N_11594,N_4419,N_4188);
or U11595 (N_11595,N_3337,N_5500);
nand U11596 (N_11596,N_899,N_2661);
nand U11597 (N_11597,N_2114,N_4837);
and U11598 (N_11598,N_1308,N_1598);
or U11599 (N_11599,N_4611,N_2163);
nand U11600 (N_11600,N_1115,N_3783);
or U11601 (N_11601,N_3995,N_1913);
nor U11602 (N_11602,N_764,N_5525);
and U11603 (N_11603,N_3488,N_4814);
and U11604 (N_11604,N_376,N_3922);
or U11605 (N_11605,N_2205,N_2799);
or U11606 (N_11606,N_2157,N_5867);
nand U11607 (N_11607,N_4131,N_4289);
xnor U11608 (N_11608,N_5100,N_1238);
and U11609 (N_11609,N_1950,N_2781);
or U11610 (N_11610,N_2443,N_3388);
nand U11611 (N_11611,N_6170,N_3074);
nand U11612 (N_11612,N_2773,N_306);
xnor U11613 (N_11613,N_5798,N_5426);
or U11614 (N_11614,N_4795,N_5659);
nand U11615 (N_11615,N_5911,N_5195);
nor U11616 (N_11616,N_1575,N_1423);
nand U11617 (N_11617,N_5853,N_2587);
nand U11618 (N_11618,N_573,N_3582);
nand U11619 (N_11619,N_3304,N_1389);
or U11620 (N_11620,N_2481,N_2675);
or U11621 (N_11621,N_4309,N_5441);
and U11622 (N_11622,N_5434,N_2250);
nor U11623 (N_11623,N_1388,N_537);
xnor U11624 (N_11624,N_5910,N_1332);
and U11625 (N_11625,N_205,N_4442);
nor U11626 (N_11626,N_921,N_3747);
and U11627 (N_11627,N_4787,N_5573);
nor U11628 (N_11628,N_2766,N_5553);
or U11629 (N_11629,N_330,N_2818);
nand U11630 (N_11630,N_272,N_516);
or U11631 (N_11631,N_2427,N_5679);
or U11632 (N_11632,N_750,N_4492);
nand U11633 (N_11633,N_1247,N_4287);
and U11634 (N_11634,N_3368,N_1041);
or U11635 (N_11635,N_86,N_1964);
xor U11636 (N_11636,N_525,N_967);
or U11637 (N_11637,N_1840,N_1301);
or U11638 (N_11638,N_4430,N_928);
and U11639 (N_11639,N_48,N_2929);
nand U11640 (N_11640,N_6115,N_582);
nand U11641 (N_11641,N_1604,N_4677);
nand U11642 (N_11642,N_2674,N_6148);
and U11643 (N_11643,N_1029,N_5299);
or U11644 (N_11644,N_5440,N_2092);
nor U11645 (N_11645,N_1881,N_5708);
nor U11646 (N_11646,N_4473,N_6015);
and U11647 (N_11647,N_4284,N_2793);
nand U11648 (N_11648,N_3149,N_3179);
nand U11649 (N_11649,N_2664,N_3992);
nor U11650 (N_11650,N_4422,N_247);
and U11651 (N_11651,N_5004,N_5634);
xor U11652 (N_11652,N_2409,N_2761);
and U11653 (N_11653,N_217,N_723);
nor U11654 (N_11654,N_4774,N_5990);
nor U11655 (N_11655,N_3050,N_3128);
and U11656 (N_11656,N_59,N_2561);
nor U11657 (N_11657,N_2168,N_4344);
nor U11658 (N_11658,N_3632,N_2155);
and U11659 (N_11659,N_1920,N_693);
xnor U11660 (N_11660,N_2522,N_5344);
nand U11661 (N_11661,N_5177,N_1538);
nand U11662 (N_11662,N_23,N_4711);
nand U11663 (N_11663,N_5181,N_170);
and U11664 (N_11664,N_1288,N_1055);
or U11665 (N_11665,N_2850,N_2364);
or U11666 (N_11666,N_4271,N_3585);
or U11667 (N_11667,N_3769,N_6048);
nor U11668 (N_11668,N_1628,N_318);
or U11669 (N_11669,N_2236,N_2114);
nor U11670 (N_11670,N_2375,N_4512);
nor U11671 (N_11671,N_4405,N_1317);
or U11672 (N_11672,N_3578,N_3300);
xnor U11673 (N_11673,N_1827,N_5887);
and U11674 (N_11674,N_3090,N_1430);
xor U11675 (N_11675,N_5489,N_246);
and U11676 (N_11676,N_2788,N_5873);
and U11677 (N_11677,N_622,N_4378);
xnor U11678 (N_11678,N_587,N_5508);
nor U11679 (N_11679,N_3997,N_3086);
nand U11680 (N_11680,N_199,N_2992);
or U11681 (N_11681,N_3401,N_6072);
or U11682 (N_11682,N_4394,N_5320);
or U11683 (N_11683,N_5920,N_3538);
nor U11684 (N_11684,N_4187,N_5116);
xnor U11685 (N_11685,N_1480,N_3423);
nand U11686 (N_11686,N_5368,N_1854);
and U11687 (N_11687,N_3369,N_4844);
xor U11688 (N_11688,N_4530,N_2416);
nor U11689 (N_11689,N_2932,N_4808);
nor U11690 (N_11690,N_2223,N_1142);
nor U11691 (N_11691,N_2341,N_6210);
or U11692 (N_11692,N_2937,N_1954);
and U11693 (N_11693,N_4634,N_2861);
nor U11694 (N_11694,N_5476,N_4436);
nand U11695 (N_11695,N_5517,N_4759);
and U11696 (N_11696,N_1849,N_6170);
nand U11697 (N_11697,N_5444,N_3431);
nor U11698 (N_11698,N_428,N_5139);
and U11699 (N_11699,N_1548,N_1071);
xor U11700 (N_11700,N_5039,N_3744);
nand U11701 (N_11701,N_1389,N_3105);
or U11702 (N_11702,N_2962,N_5628);
and U11703 (N_11703,N_5822,N_359);
nand U11704 (N_11704,N_4693,N_1782);
nand U11705 (N_11705,N_5495,N_3453);
nor U11706 (N_11706,N_4782,N_1177);
or U11707 (N_11707,N_3098,N_5672);
xnor U11708 (N_11708,N_4393,N_5340);
nand U11709 (N_11709,N_2353,N_2675);
or U11710 (N_11710,N_877,N_5064);
nor U11711 (N_11711,N_5568,N_5053);
and U11712 (N_11712,N_4754,N_2260);
and U11713 (N_11713,N_2850,N_4501);
nor U11714 (N_11714,N_4931,N_722);
nor U11715 (N_11715,N_1658,N_4276);
or U11716 (N_11716,N_2212,N_424);
nand U11717 (N_11717,N_856,N_1271);
nand U11718 (N_11718,N_4649,N_3146);
nor U11719 (N_11719,N_2123,N_1572);
or U11720 (N_11720,N_3466,N_1802);
and U11721 (N_11721,N_436,N_4160);
and U11722 (N_11722,N_1493,N_570);
and U11723 (N_11723,N_996,N_4340);
or U11724 (N_11724,N_677,N_904);
nor U11725 (N_11725,N_4673,N_462);
nor U11726 (N_11726,N_5600,N_4276);
nand U11727 (N_11727,N_5624,N_5028);
xnor U11728 (N_11728,N_1781,N_2927);
nor U11729 (N_11729,N_761,N_2904);
nor U11730 (N_11730,N_969,N_6075);
nor U11731 (N_11731,N_4322,N_5310);
nor U11732 (N_11732,N_910,N_5796);
nand U11733 (N_11733,N_3215,N_3786);
and U11734 (N_11734,N_779,N_955);
nand U11735 (N_11735,N_4263,N_663);
xnor U11736 (N_11736,N_4802,N_3647);
and U11737 (N_11737,N_2857,N_4597);
or U11738 (N_11738,N_4844,N_1479);
nor U11739 (N_11739,N_1406,N_1691);
nor U11740 (N_11740,N_2139,N_1377);
nand U11741 (N_11741,N_568,N_3784);
nor U11742 (N_11742,N_3670,N_2402);
nor U11743 (N_11743,N_3338,N_2823);
nor U11744 (N_11744,N_5569,N_6083);
and U11745 (N_11745,N_6248,N_4632);
nor U11746 (N_11746,N_1992,N_1048);
nand U11747 (N_11747,N_723,N_6227);
or U11748 (N_11748,N_5339,N_5901);
nor U11749 (N_11749,N_5536,N_5358);
and U11750 (N_11750,N_1070,N_5079);
or U11751 (N_11751,N_1162,N_3504);
and U11752 (N_11752,N_4630,N_657);
nand U11753 (N_11753,N_1536,N_554);
and U11754 (N_11754,N_2919,N_1818);
and U11755 (N_11755,N_3617,N_2755);
nor U11756 (N_11756,N_5001,N_2881);
xnor U11757 (N_11757,N_4817,N_310);
nand U11758 (N_11758,N_2326,N_3598);
and U11759 (N_11759,N_4276,N_875);
and U11760 (N_11760,N_2210,N_2762);
nor U11761 (N_11761,N_3787,N_4560);
nand U11762 (N_11762,N_5059,N_2654);
xor U11763 (N_11763,N_2376,N_1257);
nand U11764 (N_11764,N_2014,N_1033);
and U11765 (N_11765,N_5350,N_5845);
nand U11766 (N_11766,N_5982,N_1794);
and U11767 (N_11767,N_2141,N_4741);
nor U11768 (N_11768,N_3723,N_2964);
nand U11769 (N_11769,N_618,N_3984);
and U11770 (N_11770,N_1766,N_5611);
xnor U11771 (N_11771,N_355,N_1814);
and U11772 (N_11772,N_2684,N_589);
nand U11773 (N_11773,N_119,N_4577);
nor U11774 (N_11774,N_6102,N_4635);
or U11775 (N_11775,N_5923,N_1342);
or U11776 (N_11776,N_5059,N_491);
nand U11777 (N_11777,N_2394,N_5081);
nand U11778 (N_11778,N_4268,N_4713);
nor U11779 (N_11779,N_4267,N_5509);
nand U11780 (N_11780,N_2999,N_571);
nand U11781 (N_11781,N_5097,N_3725);
and U11782 (N_11782,N_4590,N_4237);
nor U11783 (N_11783,N_337,N_350);
nor U11784 (N_11784,N_6059,N_3234);
nand U11785 (N_11785,N_118,N_4830);
nand U11786 (N_11786,N_1927,N_5909);
nand U11787 (N_11787,N_2510,N_2372);
and U11788 (N_11788,N_4053,N_937);
nor U11789 (N_11789,N_3354,N_1440);
or U11790 (N_11790,N_694,N_3581);
nor U11791 (N_11791,N_1430,N_5416);
and U11792 (N_11792,N_5544,N_5898);
or U11793 (N_11793,N_2443,N_1904);
and U11794 (N_11794,N_2370,N_2158);
xor U11795 (N_11795,N_6225,N_65);
nor U11796 (N_11796,N_2606,N_3220);
nand U11797 (N_11797,N_4865,N_2318);
nor U11798 (N_11798,N_3044,N_5761);
nand U11799 (N_11799,N_5160,N_1446);
nand U11800 (N_11800,N_5871,N_4683);
nor U11801 (N_11801,N_2063,N_1000);
nand U11802 (N_11802,N_2703,N_5016);
nor U11803 (N_11803,N_2538,N_3360);
or U11804 (N_11804,N_1718,N_3735);
or U11805 (N_11805,N_2027,N_676);
nand U11806 (N_11806,N_1126,N_3625);
and U11807 (N_11807,N_4560,N_3138);
or U11808 (N_11808,N_4337,N_6164);
and U11809 (N_11809,N_6043,N_3710);
nor U11810 (N_11810,N_1802,N_3223);
xnor U11811 (N_11811,N_2279,N_1530);
nand U11812 (N_11812,N_4047,N_4178);
and U11813 (N_11813,N_117,N_390);
and U11814 (N_11814,N_271,N_467);
and U11815 (N_11815,N_2253,N_2702);
nand U11816 (N_11816,N_1660,N_2470);
nor U11817 (N_11817,N_2967,N_3434);
or U11818 (N_11818,N_4760,N_3234);
or U11819 (N_11819,N_4955,N_2610);
or U11820 (N_11820,N_53,N_1023);
nand U11821 (N_11821,N_2814,N_582);
or U11822 (N_11822,N_1984,N_3585);
nand U11823 (N_11823,N_5401,N_4019);
xor U11824 (N_11824,N_3690,N_5647);
nand U11825 (N_11825,N_2478,N_499);
nand U11826 (N_11826,N_4352,N_5874);
nor U11827 (N_11827,N_3391,N_5202);
nand U11828 (N_11828,N_6085,N_6183);
and U11829 (N_11829,N_258,N_4132);
or U11830 (N_11830,N_2788,N_2007);
or U11831 (N_11831,N_6209,N_1345);
and U11832 (N_11832,N_4589,N_2692);
and U11833 (N_11833,N_800,N_533);
or U11834 (N_11834,N_2158,N_5150);
nor U11835 (N_11835,N_21,N_998);
nand U11836 (N_11836,N_4555,N_3617);
nand U11837 (N_11837,N_3457,N_2637);
and U11838 (N_11838,N_4182,N_4318);
and U11839 (N_11839,N_3329,N_5751);
and U11840 (N_11840,N_6021,N_3283);
nor U11841 (N_11841,N_929,N_72);
nand U11842 (N_11842,N_4163,N_3776);
and U11843 (N_11843,N_2140,N_409);
or U11844 (N_11844,N_3624,N_3874);
and U11845 (N_11845,N_58,N_5664);
or U11846 (N_11846,N_330,N_3630);
xor U11847 (N_11847,N_4224,N_5944);
or U11848 (N_11848,N_5004,N_2796);
and U11849 (N_11849,N_741,N_4656);
nand U11850 (N_11850,N_2722,N_1049);
and U11851 (N_11851,N_2951,N_471);
or U11852 (N_11852,N_1872,N_1363);
nor U11853 (N_11853,N_3367,N_4967);
and U11854 (N_11854,N_6148,N_169);
and U11855 (N_11855,N_2359,N_659);
nor U11856 (N_11856,N_5753,N_3070);
and U11857 (N_11857,N_4746,N_457);
or U11858 (N_11858,N_89,N_6062);
nand U11859 (N_11859,N_1145,N_3228);
nor U11860 (N_11860,N_6207,N_1504);
nand U11861 (N_11861,N_2551,N_1862);
xor U11862 (N_11862,N_5882,N_3881);
and U11863 (N_11863,N_4402,N_4882);
and U11864 (N_11864,N_4152,N_5368);
nand U11865 (N_11865,N_1048,N_5585);
nor U11866 (N_11866,N_3060,N_1328);
xor U11867 (N_11867,N_3192,N_1871);
nand U11868 (N_11868,N_4602,N_5044);
and U11869 (N_11869,N_5765,N_5098);
nand U11870 (N_11870,N_1262,N_3920);
and U11871 (N_11871,N_5049,N_441);
nand U11872 (N_11872,N_5135,N_907);
nand U11873 (N_11873,N_4905,N_5131);
nand U11874 (N_11874,N_647,N_6145);
xor U11875 (N_11875,N_5327,N_2131);
nor U11876 (N_11876,N_1168,N_2151);
nand U11877 (N_11877,N_1915,N_3844);
or U11878 (N_11878,N_6233,N_6124);
nor U11879 (N_11879,N_860,N_1363);
and U11880 (N_11880,N_1747,N_1677);
nor U11881 (N_11881,N_4727,N_4475);
nor U11882 (N_11882,N_1966,N_4958);
or U11883 (N_11883,N_4843,N_1255);
nor U11884 (N_11884,N_2262,N_49);
and U11885 (N_11885,N_670,N_2236);
or U11886 (N_11886,N_5498,N_1523);
nor U11887 (N_11887,N_5928,N_5560);
nand U11888 (N_11888,N_408,N_3612);
and U11889 (N_11889,N_4287,N_2978);
nor U11890 (N_11890,N_5503,N_4700);
and U11891 (N_11891,N_5330,N_5577);
nand U11892 (N_11892,N_2016,N_3439);
nor U11893 (N_11893,N_5986,N_606);
nor U11894 (N_11894,N_1643,N_2760);
or U11895 (N_11895,N_4869,N_2924);
or U11896 (N_11896,N_3760,N_2159);
and U11897 (N_11897,N_1068,N_4267);
and U11898 (N_11898,N_6171,N_1886);
nand U11899 (N_11899,N_988,N_5554);
and U11900 (N_11900,N_2135,N_3629);
and U11901 (N_11901,N_6212,N_5838);
or U11902 (N_11902,N_4278,N_5511);
nor U11903 (N_11903,N_4804,N_5636);
and U11904 (N_11904,N_175,N_4758);
nor U11905 (N_11905,N_2317,N_965);
or U11906 (N_11906,N_371,N_1695);
or U11907 (N_11907,N_896,N_1264);
nand U11908 (N_11908,N_2134,N_4734);
and U11909 (N_11909,N_2258,N_5612);
or U11910 (N_11910,N_120,N_869);
or U11911 (N_11911,N_2499,N_352);
nand U11912 (N_11912,N_242,N_231);
nand U11913 (N_11913,N_474,N_2506);
nand U11914 (N_11914,N_311,N_4040);
xor U11915 (N_11915,N_3359,N_674);
or U11916 (N_11916,N_5042,N_5553);
or U11917 (N_11917,N_3020,N_4199);
and U11918 (N_11918,N_80,N_2410);
nand U11919 (N_11919,N_5026,N_900);
or U11920 (N_11920,N_1487,N_4132);
nor U11921 (N_11921,N_1643,N_3415);
nor U11922 (N_11922,N_5802,N_4538);
and U11923 (N_11923,N_4113,N_1484);
nor U11924 (N_11924,N_5152,N_2676);
or U11925 (N_11925,N_6196,N_2541);
or U11926 (N_11926,N_2119,N_634);
nor U11927 (N_11927,N_2668,N_1987);
and U11928 (N_11928,N_4342,N_4989);
nor U11929 (N_11929,N_3146,N_3708);
nor U11930 (N_11930,N_5896,N_5823);
or U11931 (N_11931,N_1881,N_4278);
xnor U11932 (N_11932,N_413,N_515);
or U11933 (N_11933,N_2252,N_1238);
nor U11934 (N_11934,N_4363,N_60);
or U11935 (N_11935,N_2477,N_191);
nor U11936 (N_11936,N_331,N_6113);
or U11937 (N_11937,N_712,N_3479);
nand U11938 (N_11938,N_3732,N_86);
xnor U11939 (N_11939,N_2048,N_63);
nand U11940 (N_11940,N_4428,N_558);
nor U11941 (N_11941,N_5449,N_753);
xor U11942 (N_11942,N_3864,N_718);
nor U11943 (N_11943,N_4864,N_490);
or U11944 (N_11944,N_1172,N_2173);
and U11945 (N_11945,N_4035,N_365);
and U11946 (N_11946,N_5588,N_4934);
xnor U11947 (N_11947,N_5233,N_4908);
and U11948 (N_11948,N_922,N_2586);
and U11949 (N_11949,N_5693,N_2638);
and U11950 (N_11950,N_345,N_5965);
nand U11951 (N_11951,N_6096,N_2727);
nand U11952 (N_11952,N_513,N_3189);
and U11953 (N_11953,N_2973,N_6235);
or U11954 (N_11954,N_31,N_3023);
nor U11955 (N_11955,N_5780,N_2674);
nand U11956 (N_11956,N_983,N_1472);
nand U11957 (N_11957,N_3720,N_934);
or U11958 (N_11958,N_2241,N_3997);
or U11959 (N_11959,N_3093,N_1908);
nand U11960 (N_11960,N_2831,N_1830);
nand U11961 (N_11961,N_1206,N_5853);
or U11962 (N_11962,N_773,N_1080);
or U11963 (N_11963,N_3954,N_2890);
and U11964 (N_11964,N_1899,N_2874);
xor U11965 (N_11965,N_3615,N_334);
and U11966 (N_11966,N_5253,N_605);
nor U11967 (N_11967,N_2383,N_824);
xor U11968 (N_11968,N_4307,N_4450);
nand U11969 (N_11969,N_6106,N_5599);
or U11970 (N_11970,N_5578,N_1593);
or U11971 (N_11971,N_579,N_5299);
and U11972 (N_11972,N_3953,N_1514);
nor U11973 (N_11973,N_741,N_5913);
or U11974 (N_11974,N_2115,N_5424);
xnor U11975 (N_11975,N_3726,N_946);
xor U11976 (N_11976,N_247,N_6220);
and U11977 (N_11977,N_5937,N_5510);
nand U11978 (N_11978,N_2470,N_4103);
nor U11979 (N_11979,N_4633,N_1882);
nor U11980 (N_11980,N_1809,N_5112);
nor U11981 (N_11981,N_1313,N_3799);
nand U11982 (N_11982,N_5481,N_2587);
and U11983 (N_11983,N_1037,N_4181);
nor U11984 (N_11984,N_4768,N_1106);
and U11985 (N_11985,N_5418,N_1596);
nand U11986 (N_11986,N_6217,N_36);
nor U11987 (N_11987,N_837,N_5303);
or U11988 (N_11988,N_590,N_108);
or U11989 (N_11989,N_4075,N_677);
nor U11990 (N_11990,N_1286,N_2874);
or U11991 (N_11991,N_4260,N_2156);
nand U11992 (N_11992,N_187,N_4876);
nand U11993 (N_11993,N_2653,N_1823);
and U11994 (N_11994,N_4286,N_4841);
or U11995 (N_11995,N_2736,N_4460);
or U11996 (N_11996,N_3063,N_2988);
or U11997 (N_11997,N_3100,N_5987);
nand U11998 (N_11998,N_3644,N_2841);
nand U11999 (N_11999,N_3973,N_1088);
xnor U12000 (N_12000,N_630,N_2851);
nor U12001 (N_12001,N_1879,N_1841);
xor U12002 (N_12002,N_5669,N_1635);
or U12003 (N_12003,N_3933,N_263);
nand U12004 (N_12004,N_2239,N_5749);
nor U12005 (N_12005,N_4552,N_1086);
nand U12006 (N_12006,N_2230,N_1339);
nor U12007 (N_12007,N_2445,N_1152);
nor U12008 (N_12008,N_1214,N_6114);
nor U12009 (N_12009,N_52,N_5221);
and U12010 (N_12010,N_4770,N_3716);
or U12011 (N_12011,N_1436,N_6245);
or U12012 (N_12012,N_251,N_6001);
and U12013 (N_12013,N_6114,N_4597);
or U12014 (N_12014,N_5273,N_2285);
or U12015 (N_12015,N_4599,N_6007);
or U12016 (N_12016,N_522,N_1031);
or U12017 (N_12017,N_3769,N_4866);
nand U12018 (N_12018,N_1911,N_65);
or U12019 (N_12019,N_4151,N_2086);
nand U12020 (N_12020,N_1022,N_4020);
nand U12021 (N_12021,N_5269,N_5069);
or U12022 (N_12022,N_3853,N_5375);
nand U12023 (N_12023,N_1853,N_3562);
nand U12024 (N_12024,N_5627,N_3854);
xor U12025 (N_12025,N_2254,N_3540);
and U12026 (N_12026,N_4652,N_1522);
nand U12027 (N_12027,N_6103,N_499);
and U12028 (N_12028,N_4483,N_4811);
nand U12029 (N_12029,N_5923,N_3187);
and U12030 (N_12030,N_6192,N_3010);
nor U12031 (N_12031,N_647,N_6056);
or U12032 (N_12032,N_2459,N_1838);
nand U12033 (N_12033,N_65,N_213);
nor U12034 (N_12034,N_2736,N_5279);
nand U12035 (N_12035,N_4758,N_4039);
and U12036 (N_12036,N_1796,N_3187);
or U12037 (N_12037,N_5215,N_1189);
or U12038 (N_12038,N_6038,N_2037);
xnor U12039 (N_12039,N_1685,N_603);
nor U12040 (N_12040,N_4817,N_4561);
and U12041 (N_12041,N_370,N_1814);
xnor U12042 (N_12042,N_460,N_756);
or U12043 (N_12043,N_62,N_3767);
and U12044 (N_12044,N_6176,N_5905);
xnor U12045 (N_12045,N_61,N_835);
or U12046 (N_12046,N_3967,N_3737);
nand U12047 (N_12047,N_4101,N_1526);
or U12048 (N_12048,N_798,N_3983);
nand U12049 (N_12049,N_845,N_1018);
nor U12050 (N_12050,N_3431,N_603);
or U12051 (N_12051,N_1607,N_6045);
or U12052 (N_12052,N_3136,N_4035);
nor U12053 (N_12053,N_5141,N_4137);
nor U12054 (N_12054,N_2752,N_1590);
or U12055 (N_12055,N_1947,N_421);
nor U12056 (N_12056,N_1870,N_2637);
or U12057 (N_12057,N_5084,N_1227);
nand U12058 (N_12058,N_479,N_267);
nor U12059 (N_12059,N_2570,N_1688);
nand U12060 (N_12060,N_3788,N_2377);
nand U12061 (N_12061,N_3655,N_5311);
and U12062 (N_12062,N_3387,N_1538);
or U12063 (N_12063,N_598,N_2639);
xor U12064 (N_12064,N_1646,N_2061);
nor U12065 (N_12065,N_3447,N_3143);
or U12066 (N_12066,N_4886,N_660);
nand U12067 (N_12067,N_277,N_2439);
xor U12068 (N_12068,N_4239,N_2897);
nand U12069 (N_12069,N_5934,N_1756);
xnor U12070 (N_12070,N_4483,N_710);
nor U12071 (N_12071,N_6047,N_1316);
xor U12072 (N_12072,N_4350,N_4407);
and U12073 (N_12073,N_4658,N_5311);
nor U12074 (N_12074,N_1017,N_4615);
nand U12075 (N_12075,N_1165,N_2796);
and U12076 (N_12076,N_6130,N_3676);
or U12077 (N_12077,N_3923,N_1669);
or U12078 (N_12078,N_4236,N_3148);
nand U12079 (N_12079,N_6203,N_4985);
nor U12080 (N_12080,N_2125,N_7);
or U12081 (N_12081,N_5729,N_4275);
and U12082 (N_12082,N_124,N_2958);
nor U12083 (N_12083,N_2752,N_237);
nor U12084 (N_12084,N_3625,N_5537);
nor U12085 (N_12085,N_5982,N_4063);
xnor U12086 (N_12086,N_2133,N_3395);
and U12087 (N_12087,N_150,N_307);
xor U12088 (N_12088,N_2631,N_673);
nand U12089 (N_12089,N_4241,N_5394);
nor U12090 (N_12090,N_3107,N_2043);
nor U12091 (N_12091,N_3826,N_6215);
or U12092 (N_12092,N_2121,N_2988);
or U12093 (N_12093,N_4880,N_3677);
nand U12094 (N_12094,N_2535,N_5020);
nand U12095 (N_12095,N_2429,N_1877);
xnor U12096 (N_12096,N_3087,N_4255);
or U12097 (N_12097,N_5907,N_3773);
or U12098 (N_12098,N_2099,N_6004);
and U12099 (N_12099,N_5894,N_4628);
nor U12100 (N_12100,N_4362,N_4441);
or U12101 (N_12101,N_6029,N_4351);
nand U12102 (N_12102,N_5112,N_2798);
nand U12103 (N_12103,N_3362,N_4814);
and U12104 (N_12104,N_294,N_3229);
or U12105 (N_12105,N_2876,N_4446);
and U12106 (N_12106,N_3683,N_26);
or U12107 (N_12107,N_5342,N_4331);
nor U12108 (N_12108,N_2420,N_3651);
nand U12109 (N_12109,N_4956,N_3517);
or U12110 (N_12110,N_2306,N_3463);
or U12111 (N_12111,N_2187,N_5529);
nor U12112 (N_12112,N_4699,N_1419);
nand U12113 (N_12113,N_6117,N_4184);
and U12114 (N_12114,N_3087,N_540);
nor U12115 (N_12115,N_2028,N_5902);
or U12116 (N_12116,N_823,N_636);
xor U12117 (N_12117,N_5426,N_1417);
nor U12118 (N_12118,N_4470,N_1767);
or U12119 (N_12119,N_5803,N_3083);
nor U12120 (N_12120,N_1166,N_2778);
nand U12121 (N_12121,N_3906,N_1290);
and U12122 (N_12122,N_1806,N_1372);
or U12123 (N_12123,N_5084,N_4630);
nor U12124 (N_12124,N_4963,N_4334);
nand U12125 (N_12125,N_5544,N_2464);
and U12126 (N_12126,N_1592,N_3055);
xor U12127 (N_12127,N_2598,N_2622);
xnor U12128 (N_12128,N_1912,N_947);
and U12129 (N_12129,N_1843,N_415);
and U12130 (N_12130,N_551,N_6048);
and U12131 (N_12131,N_996,N_1180);
or U12132 (N_12132,N_808,N_2433);
or U12133 (N_12133,N_2676,N_1317);
or U12134 (N_12134,N_2096,N_4179);
nand U12135 (N_12135,N_4512,N_3604);
nand U12136 (N_12136,N_2436,N_3778);
and U12137 (N_12137,N_4625,N_4472);
or U12138 (N_12138,N_1152,N_3129);
or U12139 (N_12139,N_3114,N_1287);
nor U12140 (N_12140,N_2817,N_4431);
nor U12141 (N_12141,N_3529,N_3397);
and U12142 (N_12142,N_4799,N_5287);
and U12143 (N_12143,N_3750,N_3492);
nor U12144 (N_12144,N_4184,N_3325);
nand U12145 (N_12145,N_2759,N_847);
and U12146 (N_12146,N_2138,N_5231);
and U12147 (N_12147,N_6021,N_4694);
and U12148 (N_12148,N_4046,N_5394);
and U12149 (N_12149,N_2224,N_2649);
or U12150 (N_12150,N_4631,N_5835);
or U12151 (N_12151,N_5012,N_4897);
nand U12152 (N_12152,N_3772,N_5867);
or U12153 (N_12153,N_2186,N_383);
or U12154 (N_12154,N_3312,N_3793);
and U12155 (N_12155,N_2197,N_3333);
nor U12156 (N_12156,N_5915,N_5212);
nand U12157 (N_12157,N_5666,N_2894);
or U12158 (N_12158,N_1614,N_460);
or U12159 (N_12159,N_2196,N_3577);
nand U12160 (N_12160,N_4586,N_3264);
and U12161 (N_12161,N_335,N_5061);
and U12162 (N_12162,N_3911,N_5796);
and U12163 (N_12163,N_6039,N_2030);
and U12164 (N_12164,N_5519,N_3839);
or U12165 (N_12165,N_5805,N_374);
nor U12166 (N_12166,N_5582,N_3586);
nand U12167 (N_12167,N_3162,N_4565);
nor U12168 (N_12168,N_4294,N_5850);
or U12169 (N_12169,N_3128,N_125);
nor U12170 (N_12170,N_2792,N_1889);
or U12171 (N_12171,N_1537,N_4473);
and U12172 (N_12172,N_2588,N_5155);
and U12173 (N_12173,N_3359,N_6077);
nand U12174 (N_12174,N_664,N_858);
or U12175 (N_12175,N_772,N_963);
and U12176 (N_12176,N_3252,N_5297);
or U12177 (N_12177,N_5002,N_2558);
nand U12178 (N_12178,N_5849,N_4023);
or U12179 (N_12179,N_4701,N_1426);
nor U12180 (N_12180,N_3055,N_318);
and U12181 (N_12181,N_1164,N_4235);
and U12182 (N_12182,N_4313,N_4588);
nand U12183 (N_12183,N_4365,N_2223);
nand U12184 (N_12184,N_1729,N_1444);
and U12185 (N_12185,N_3622,N_526);
or U12186 (N_12186,N_1253,N_3795);
nand U12187 (N_12187,N_5448,N_5769);
nand U12188 (N_12188,N_4975,N_2494);
nand U12189 (N_12189,N_4946,N_4372);
nor U12190 (N_12190,N_4196,N_5056);
nand U12191 (N_12191,N_4199,N_5835);
or U12192 (N_12192,N_3449,N_3693);
or U12193 (N_12193,N_1526,N_2481);
xnor U12194 (N_12194,N_5228,N_3303);
or U12195 (N_12195,N_650,N_854);
and U12196 (N_12196,N_1902,N_5929);
nand U12197 (N_12197,N_4903,N_1120);
xor U12198 (N_12198,N_4453,N_5257);
and U12199 (N_12199,N_2821,N_5106);
nand U12200 (N_12200,N_5244,N_3133);
nand U12201 (N_12201,N_1299,N_3109);
or U12202 (N_12202,N_4087,N_759);
and U12203 (N_12203,N_4611,N_1720);
and U12204 (N_12204,N_372,N_327);
nor U12205 (N_12205,N_4954,N_2075);
nor U12206 (N_12206,N_1833,N_3144);
nor U12207 (N_12207,N_5176,N_2355);
nand U12208 (N_12208,N_360,N_1305);
nor U12209 (N_12209,N_3565,N_2179);
xnor U12210 (N_12210,N_4653,N_2863);
and U12211 (N_12211,N_5471,N_2489);
nor U12212 (N_12212,N_5968,N_2227);
and U12213 (N_12213,N_4759,N_3193);
xor U12214 (N_12214,N_1351,N_5341);
nor U12215 (N_12215,N_3483,N_537);
xnor U12216 (N_12216,N_5775,N_4800);
xor U12217 (N_12217,N_5451,N_5955);
or U12218 (N_12218,N_5903,N_1075);
or U12219 (N_12219,N_2212,N_3533);
nand U12220 (N_12220,N_4866,N_4364);
xnor U12221 (N_12221,N_926,N_4847);
or U12222 (N_12222,N_2706,N_4373);
nor U12223 (N_12223,N_5916,N_4137);
nand U12224 (N_12224,N_516,N_3483);
and U12225 (N_12225,N_1464,N_2376);
nor U12226 (N_12226,N_2258,N_3836);
or U12227 (N_12227,N_4275,N_559);
nand U12228 (N_12228,N_1101,N_2844);
nand U12229 (N_12229,N_5181,N_2616);
or U12230 (N_12230,N_1218,N_5236);
nor U12231 (N_12231,N_4834,N_5481);
nor U12232 (N_12232,N_6069,N_3016);
nand U12233 (N_12233,N_4270,N_3863);
nand U12234 (N_12234,N_3792,N_2011);
and U12235 (N_12235,N_3623,N_5348);
and U12236 (N_12236,N_4592,N_2474);
and U12237 (N_12237,N_1101,N_2523);
nor U12238 (N_12238,N_5422,N_2661);
or U12239 (N_12239,N_1829,N_658);
nand U12240 (N_12240,N_2686,N_2325);
and U12241 (N_12241,N_2222,N_4545);
nor U12242 (N_12242,N_4478,N_5024);
or U12243 (N_12243,N_4972,N_2591);
or U12244 (N_12244,N_3321,N_4044);
nand U12245 (N_12245,N_4331,N_5678);
nand U12246 (N_12246,N_2766,N_858);
xor U12247 (N_12247,N_3800,N_4075);
nor U12248 (N_12248,N_709,N_5222);
and U12249 (N_12249,N_2730,N_4081);
nand U12250 (N_12250,N_3386,N_4093);
nand U12251 (N_12251,N_4991,N_5390);
or U12252 (N_12252,N_1937,N_3632);
nand U12253 (N_12253,N_5856,N_5610);
nand U12254 (N_12254,N_5540,N_5897);
xnor U12255 (N_12255,N_5590,N_1771);
nand U12256 (N_12256,N_526,N_5287);
nand U12257 (N_12257,N_2660,N_4819);
nand U12258 (N_12258,N_870,N_443);
or U12259 (N_12259,N_4981,N_529);
nor U12260 (N_12260,N_4448,N_955);
or U12261 (N_12261,N_5270,N_2925);
nand U12262 (N_12262,N_5171,N_3424);
or U12263 (N_12263,N_5496,N_3746);
xnor U12264 (N_12264,N_578,N_4502);
nor U12265 (N_12265,N_2840,N_1914);
nand U12266 (N_12266,N_710,N_2782);
nand U12267 (N_12267,N_3157,N_5126);
nand U12268 (N_12268,N_3247,N_3226);
and U12269 (N_12269,N_3999,N_2146);
nand U12270 (N_12270,N_1499,N_1087);
nor U12271 (N_12271,N_4667,N_2185);
nand U12272 (N_12272,N_5163,N_3082);
nor U12273 (N_12273,N_3852,N_2125);
nor U12274 (N_12274,N_1479,N_3209);
and U12275 (N_12275,N_3808,N_5868);
and U12276 (N_12276,N_2079,N_3540);
or U12277 (N_12277,N_2762,N_3879);
nand U12278 (N_12278,N_1556,N_98);
and U12279 (N_12279,N_633,N_735);
and U12280 (N_12280,N_1050,N_1005);
or U12281 (N_12281,N_3076,N_4877);
nor U12282 (N_12282,N_2277,N_3447);
nor U12283 (N_12283,N_184,N_2467);
nor U12284 (N_12284,N_2963,N_3749);
and U12285 (N_12285,N_65,N_1901);
nand U12286 (N_12286,N_3777,N_1487);
nand U12287 (N_12287,N_4614,N_5723);
and U12288 (N_12288,N_4510,N_1178);
xor U12289 (N_12289,N_5231,N_5609);
nor U12290 (N_12290,N_44,N_3613);
nor U12291 (N_12291,N_3789,N_5658);
or U12292 (N_12292,N_307,N_2927);
or U12293 (N_12293,N_5009,N_2099);
and U12294 (N_12294,N_494,N_3985);
nor U12295 (N_12295,N_5108,N_2194);
nand U12296 (N_12296,N_402,N_2358);
and U12297 (N_12297,N_2709,N_144);
xnor U12298 (N_12298,N_5180,N_3430);
or U12299 (N_12299,N_5409,N_515);
xor U12300 (N_12300,N_4601,N_1252);
and U12301 (N_12301,N_1292,N_3420);
nor U12302 (N_12302,N_741,N_1035);
or U12303 (N_12303,N_4261,N_2783);
nor U12304 (N_12304,N_1731,N_4077);
nand U12305 (N_12305,N_545,N_3257);
or U12306 (N_12306,N_4552,N_1300);
nor U12307 (N_12307,N_2728,N_3064);
nor U12308 (N_12308,N_956,N_6231);
nand U12309 (N_12309,N_2199,N_5935);
nor U12310 (N_12310,N_2774,N_5236);
nor U12311 (N_12311,N_3201,N_4943);
or U12312 (N_12312,N_5222,N_2795);
nand U12313 (N_12313,N_2727,N_5482);
or U12314 (N_12314,N_2178,N_4265);
nand U12315 (N_12315,N_3063,N_391);
nor U12316 (N_12316,N_3000,N_94);
nand U12317 (N_12317,N_4868,N_3752);
nor U12318 (N_12318,N_4428,N_1635);
or U12319 (N_12319,N_2606,N_3342);
or U12320 (N_12320,N_1295,N_3565);
nand U12321 (N_12321,N_3280,N_4101);
nand U12322 (N_12322,N_5411,N_4808);
and U12323 (N_12323,N_3774,N_605);
nand U12324 (N_12324,N_4009,N_3095);
nand U12325 (N_12325,N_525,N_1145);
nor U12326 (N_12326,N_2626,N_2817);
nor U12327 (N_12327,N_5026,N_3842);
or U12328 (N_12328,N_4453,N_5685);
nor U12329 (N_12329,N_4712,N_495);
or U12330 (N_12330,N_344,N_2544);
nand U12331 (N_12331,N_1679,N_1023);
and U12332 (N_12332,N_2199,N_601);
nor U12333 (N_12333,N_1034,N_1989);
and U12334 (N_12334,N_818,N_4929);
and U12335 (N_12335,N_3374,N_979);
or U12336 (N_12336,N_3088,N_2502);
and U12337 (N_12337,N_768,N_4867);
nor U12338 (N_12338,N_3726,N_769);
and U12339 (N_12339,N_5229,N_5345);
or U12340 (N_12340,N_3107,N_2900);
and U12341 (N_12341,N_1412,N_1720);
xnor U12342 (N_12342,N_3107,N_5665);
xnor U12343 (N_12343,N_4268,N_589);
or U12344 (N_12344,N_5183,N_2738);
or U12345 (N_12345,N_3398,N_5477);
or U12346 (N_12346,N_4958,N_5492);
nand U12347 (N_12347,N_3695,N_4841);
xor U12348 (N_12348,N_4673,N_5715);
and U12349 (N_12349,N_3761,N_2343);
or U12350 (N_12350,N_5214,N_1805);
and U12351 (N_12351,N_4039,N_1630);
and U12352 (N_12352,N_3313,N_2240);
and U12353 (N_12353,N_5028,N_4124);
nand U12354 (N_12354,N_4313,N_1201);
or U12355 (N_12355,N_3333,N_1909);
or U12356 (N_12356,N_2934,N_2967);
nand U12357 (N_12357,N_2360,N_5981);
nor U12358 (N_12358,N_3952,N_4414);
nor U12359 (N_12359,N_4055,N_5);
nand U12360 (N_12360,N_924,N_2251);
and U12361 (N_12361,N_2613,N_1263);
and U12362 (N_12362,N_3635,N_3993);
nand U12363 (N_12363,N_5089,N_982);
or U12364 (N_12364,N_1875,N_1797);
and U12365 (N_12365,N_615,N_1846);
nor U12366 (N_12366,N_4047,N_687);
and U12367 (N_12367,N_1209,N_160);
nor U12368 (N_12368,N_336,N_3222);
nor U12369 (N_12369,N_2789,N_3072);
nor U12370 (N_12370,N_5846,N_4393);
and U12371 (N_12371,N_295,N_4494);
or U12372 (N_12372,N_3013,N_3894);
nand U12373 (N_12373,N_4872,N_2612);
or U12374 (N_12374,N_941,N_5374);
or U12375 (N_12375,N_4325,N_6195);
and U12376 (N_12376,N_259,N_1817);
nand U12377 (N_12377,N_4065,N_1883);
nor U12378 (N_12378,N_5747,N_5501);
xor U12379 (N_12379,N_4515,N_3442);
nand U12380 (N_12380,N_4431,N_3835);
nand U12381 (N_12381,N_2978,N_1302);
nor U12382 (N_12382,N_2343,N_2632);
and U12383 (N_12383,N_1014,N_489);
or U12384 (N_12384,N_1694,N_6044);
or U12385 (N_12385,N_3676,N_3674);
or U12386 (N_12386,N_1049,N_3530);
or U12387 (N_12387,N_2621,N_1735);
nand U12388 (N_12388,N_2474,N_3602);
nor U12389 (N_12389,N_2267,N_1029);
nand U12390 (N_12390,N_2857,N_5568);
and U12391 (N_12391,N_5683,N_2380);
or U12392 (N_12392,N_4174,N_304);
nor U12393 (N_12393,N_5918,N_4577);
and U12394 (N_12394,N_3613,N_3030);
or U12395 (N_12395,N_5332,N_4726);
nor U12396 (N_12396,N_5913,N_5214);
and U12397 (N_12397,N_5896,N_2596);
nor U12398 (N_12398,N_2826,N_440);
nand U12399 (N_12399,N_81,N_4678);
and U12400 (N_12400,N_1506,N_5970);
or U12401 (N_12401,N_5433,N_2872);
nor U12402 (N_12402,N_2506,N_3616);
or U12403 (N_12403,N_1926,N_4835);
nand U12404 (N_12404,N_4333,N_5546);
and U12405 (N_12405,N_4207,N_5110);
nand U12406 (N_12406,N_5162,N_1026);
or U12407 (N_12407,N_180,N_5953);
or U12408 (N_12408,N_1971,N_6027);
and U12409 (N_12409,N_4262,N_1978);
or U12410 (N_12410,N_1273,N_6247);
nand U12411 (N_12411,N_4153,N_3852);
nand U12412 (N_12412,N_1389,N_229);
nor U12413 (N_12413,N_5297,N_1800);
xor U12414 (N_12414,N_3858,N_97);
nand U12415 (N_12415,N_4519,N_2250);
or U12416 (N_12416,N_5944,N_2399);
xnor U12417 (N_12417,N_4590,N_806);
nor U12418 (N_12418,N_5361,N_4162);
xor U12419 (N_12419,N_2892,N_1011);
nand U12420 (N_12420,N_2627,N_1090);
xnor U12421 (N_12421,N_2010,N_5234);
and U12422 (N_12422,N_3653,N_3611);
or U12423 (N_12423,N_3705,N_2696);
and U12424 (N_12424,N_3138,N_4502);
nor U12425 (N_12425,N_3283,N_5641);
nand U12426 (N_12426,N_1172,N_1206);
nor U12427 (N_12427,N_2723,N_2911);
nor U12428 (N_12428,N_3702,N_5630);
nor U12429 (N_12429,N_2812,N_4330);
nand U12430 (N_12430,N_5806,N_3721);
and U12431 (N_12431,N_5499,N_1120);
nor U12432 (N_12432,N_1211,N_5072);
nand U12433 (N_12433,N_5573,N_1852);
nand U12434 (N_12434,N_3688,N_3698);
nor U12435 (N_12435,N_518,N_1979);
nor U12436 (N_12436,N_4531,N_2674);
nor U12437 (N_12437,N_2726,N_3370);
and U12438 (N_12438,N_3238,N_6201);
nand U12439 (N_12439,N_5739,N_5176);
or U12440 (N_12440,N_2348,N_6237);
xnor U12441 (N_12441,N_3205,N_3312);
nand U12442 (N_12442,N_3025,N_1339);
xnor U12443 (N_12443,N_599,N_3252);
nor U12444 (N_12444,N_4360,N_3888);
nand U12445 (N_12445,N_143,N_5721);
nor U12446 (N_12446,N_3785,N_679);
nor U12447 (N_12447,N_488,N_3560);
nand U12448 (N_12448,N_3894,N_3655);
or U12449 (N_12449,N_5552,N_763);
or U12450 (N_12450,N_3711,N_6115);
nand U12451 (N_12451,N_4794,N_5425);
xnor U12452 (N_12452,N_3639,N_2053);
nor U12453 (N_12453,N_3996,N_5780);
or U12454 (N_12454,N_4165,N_1322);
nor U12455 (N_12455,N_515,N_4053);
and U12456 (N_12456,N_2313,N_4276);
xor U12457 (N_12457,N_3620,N_3274);
xnor U12458 (N_12458,N_6025,N_1183);
nor U12459 (N_12459,N_3270,N_41);
xnor U12460 (N_12460,N_602,N_2897);
or U12461 (N_12461,N_1354,N_1965);
or U12462 (N_12462,N_3830,N_491);
or U12463 (N_12463,N_1522,N_2067);
nand U12464 (N_12464,N_2673,N_1907);
or U12465 (N_12465,N_3457,N_1933);
and U12466 (N_12466,N_699,N_3277);
and U12467 (N_12467,N_808,N_6139);
nor U12468 (N_12468,N_4000,N_5225);
or U12469 (N_12469,N_44,N_1175);
nor U12470 (N_12470,N_1542,N_482);
and U12471 (N_12471,N_4912,N_1527);
and U12472 (N_12472,N_4308,N_2280);
nand U12473 (N_12473,N_1757,N_981);
nor U12474 (N_12474,N_5555,N_4176);
or U12475 (N_12475,N_5824,N_4492);
nand U12476 (N_12476,N_2198,N_848);
nand U12477 (N_12477,N_6025,N_788);
nor U12478 (N_12478,N_768,N_4112);
and U12479 (N_12479,N_5259,N_256);
and U12480 (N_12480,N_306,N_4924);
nor U12481 (N_12481,N_3258,N_1379);
xor U12482 (N_12482,N_545,N_1403);
or U12483 (N_12483,N_5832,N_5615);
or U12484 (N_12484,N_1647,N_944);
or U12485 (N_12485,N_6132,N_2373);
nand U12486 (N_12486,N_5404,N_4071);
and U12487 (N_12487,N_3041,N_5775);
or U12488 (N_12488,N_4166,N_4179);
nor U12489 (N_12489,N_634,N_1566);
nand U12490 (N_12490,N_511,N_3275);
or U12491 (N_12491,N_5358,N_6181);
xor U12492 (N_12492,N_5756,N_3507);
nand U12493 (N_12493,N_4791,N_5099);
nand U12494 (N_12494,N_4695,N_2737);
nand U12495 (N_12495,N_2474,N_3533);
nor U12496 (N_12496,N_1385,N_5968);
nand U12497 (N_12497,N_2029,N_2949);
or U12498 (N_12498,N_3627,N_4202);
or U12499 (N_12499,N_4878,N_1200);
nand U12500 (N_12500,N_11712,N_11399);
nor U12501 (N_12501,N_7587,N_11202);
nor U12502 (N_12502,N_8174,N_9834);
nand U12503 (N_12503,N_11014,N_7744);
xnor U12504 (N_12504,N_9345,N_8418);
and U12505 (N_12505,N_11992,N_9688);
nand U12506 (N_12506,N_7457,N_11122);
nand U12507 (N_12507,N_6699,N_7957);
nor U12508 (N_12508,N_9281,N_10780);
xnor U12509 (N_12509,N_7043,N_12364);
and U12510 (N_12510,N_8498,N_10013);
or U12511 (N_12511,N_7946,N_11969);
nand U12512 (N_12512,N_11934,N_6692);
nor U12513 (N_12513,N_11935,N_10650);
nor U12514 (N_12514,N_12149,N_11586);
and U12515 (N_12515,N_12082,N_10579);
and U12516 (N_12516,N_10114,N_12092);
and U12517 (N_12517,N_9122,N_9203);
and U12518 (N_12518,N_7080,N_7368);
nor U12519 (N_12519,N_6460,N_8647);
xor U12520 (N_12520,N_10876,N_10739);
nor U12521 (N_12521,N_8526,N_10944);
and U12522 (N_12522,N_9803,N_10524);
nand U12523 (N_12523,N_11405,N_7428);
and U12524 (N_12524,N_12337,N_11303);
nor U12525 (N_12525,N_11048,N_10246);
nor U12526 (N_12526,N_10460,N_12150);
and U12527 (N_12527,N_11849,N_8827);
nor U12528 (N_12528,N_10840,N_9426);
nor U12529 (N_12529,N_8266,N_8606);
or U12530 (N_12530,N_12379,N_11352);
or U12531 (N_12531,N_7842,N_7093);
nand U12532 (N_12532,N_7046,N_7445);
and U12533 (N_12533,N_11836,N_7944);
and U12534 (N_12534,N_12418,N_11464);
nor U12535 (N_12535,N_11862,N_6402);
and U12536 (N_12536,N_12493,N_6573);
xor U12537 (N_12537,N_9313,N_7877);
nor U12538 (N_12538,N_9805,N_11580);
nor U12539 (N_12539,N_10490,N_6802);
nand U12540 (N_12540,N_10554,N_11851);
or U12541 (N_12541,N_9985,N_9319);
and U12542 (N_12542,N_9033,N_10311);
nand U12543 (N_12543,N_10005,N_12461);
and U12544 (N_12544,N_6723,N_6394);
nand U12545 (N_12545,N_6697,N_9637);
nand U12546 (N_12546,N_7699,N_9726);
nand U12547 (N_12547,N_6343,N_10585);
and U12548 (N_12548,N_11337,N_10727);
and U12549 (N_12549,N_12141,N_12319);
nor U12550 (N_12550,N_10115,N_10865);
nand U12551 (N_12551,N_9740,N_12458);
or U12552 (N_12552,N_10428,N_8662);
and U12553 (N_12553,N_9562,N_8106);
and U12554 (N_12554,N_12153,N_6786);
and U12555 (N_12555,N_11133,N_10623);
and U12556 (N_12556,N_11788,N_10238);
and U12557 (N_12557,N_7548,N_8254);
or U12558 (N_12558,N_9933,N_8987);
and U12559 (N_12559,N_9755,N_9452);
nand U12560 (N_12560,N_8719,N_7212);
or U12561 (N_12561,N_11302,N_7666);
nand U12562 (N_12562,N_6761,N_11694);
and U12563 (N_12563,N_12283,N_11530);
nor U12564 (N_12564,N_8824,N_11560);
nor U12565 (N_12565,N_12087,N_6937);
or U12566 (N_12566,N_9139,N_7621);
nor U12567 (N_12567,N_10297,N_9018);
nand U12568 (N_12568,N_10410,N_6878);
nand U12569 (N_12569,N_9996,N_10257);
nand U12570 (N_12570,N_8380,N_7175);
nor U12571 (N_12571,N_10863,N_10300);
nand U12572 (N_12572,N_12413,N_7658);
and U12573 (N_12573,N_12290,N_8041);
xor U12574 (N_12574,N_9647,N_11706);
nand U12575 (N_12575,N_10157,N_9550);
nor U12576 (N_12576,N_9915,N_6589);
nand U12577 (N_12577,N_8387,N_10872);
and U12578 (N_12578,N_6680,N_7302);
nand U12579 (N_12579,N_6832,N_10450);
or U12580 (N_12580,N_9476,N_7198);
xor U12581 (N_12581,N_10139,N_9750);
and U12582 (N_12582,N_6622,N_9106);
nor U12583 (N_12583,N_11168,N_9083);
and U12584 (N_12584,N_8287,N_9062);
xnor U12585 (N_12585,N_12330,N_12088);
and U12586 (N_12586,N_9797,N_6946);
xnor U12587 (N_12587,N_8938,N_11430);
xnor U12588 (N_12588,N_10642,N_8724);
nand U12589 (N_12589,N_8807,N_8375);
or U12590 (N_12590,N_8805,N_8502);
nor U12591 (N_12591,N_11717,N_9751);
or U12592 (N_12592,N_6899,N_8016);
nand U12593 (N_12593,N_9055,N_8810);
and U12594 (N_12594,N_8323,N_8439);
and U12595 (N_12595,N_7624,N_7760);
and U12596 (N_12596,N_10716,N_10708);
and U12597 (N_12597,N_8709,N_7793);
or U12598 (N_12598,N_11483,N_10845);
and U12599 (N_12599,N_11402,N_6731);
and U12600 (N_12600,N_12253,N_11299);
nand U12601 (N_12601,N_11901,N_7274);
and U12602 (N_12602,N_10160,N_11845);
nand U12603 (N_12603,N_10662,N_9618);
or U12604 (N_12604,N_6848,N_10955);
xnor U12605 (N_12605,N_11091,N_11132);
nand U12606 (N_12606,N_9419,N_10888);
or U12607 (N_12607,N_8753,N_7722);
or U12608 (N_12608,N_7253,N_10413);
or U12609 (N_12609,N_8042,N_10105);
and U12610 (N_12610,N_6547,N_7843);
and U12611 (N_12611,N_11237,N_7854);
or U12612 (N_12612,N_6433,N_9651);
nor U12613 (N_12613,N_7257,N_9232);
nor U12614 (N_12614,N_10893,N_6423);
nand U12615 (N_12615,N_6552,N_7614);
and U12616 (N_12616,N_9259,N_11798);
nor U12617 (N_12617,N_8152,N_6850);
or U12618 (N_12618,N_7585,N_11711);
nand U12619 (N_12619,N_9277,N_8221);
nand U12620 (N_12620,N_12297,N_8204);
and U12621 (N_12621,N_10804,N_7285);
nor U12622 (N_12622,N_11595,N_10758);
nor U12623 (N_12623,N_9839,N_7465);
nand U12624 (N_12624,N_9328,N_7040);
xor U12625 (N_12625,N_6774,N_8994);
xnor U12626 (N_12626,N_7815,N_8012);
or U12627 (N_12627,N_11608,N_8472);
and U12628 (N_12628,N_6755,N_6951);
nand U12629 (N_12629,N_6930,N_11701);
or U12630 (N_12630,N_8906,N_9470);
xor U12631 (N_12631,N_7995,N_7458);
and U12632 (N_12632,N_11439,N_9764);
or U12633 (N_12633,N_6868,N_7791);
or U12634 (N_12634,N_10763,N_10933);
nand U12635 (N_12635,N_11092,N_8172);
nor U12636 (N_12636,N_9733,N_6756);
nand U12637 (N_12637,N_7307,N_6505);
nor U12638 (N_12638,N_8487,N_10578);
xor U12639 (N_12639,N_10236,N_9813);
nand U12640 (N_12640,N_7738,N_6655);
and U12641 (N_12641,N_12397,N_9086);
or U12642 (N_12642,N_8252,N_12248);
nor U12643 (N_12643,N_7436,N_8836);
or U12644 (N_12644,N_8713,N_11419);
nand U12645 (N_12645,N_7128,N_9218);
nand U12646 (N_12646,N_8651,N_10978);
nor U12647 (N_12647,N_6792,N_6492);
nor U12648 (N_12648,N_10277,N_7499);
nor U12649 (N_12649,N_6443,N_11428);
or U12650 (N_12650,N_10332,N_9308);
or U12651 (N_12651,N_7862,N_8817);
xor U12652 (N_12652,N_11172,N_8674);
nand U12653 (N_12653,N_8077,N_8269);
nor U12654 (N_12654,N_11317,N_7534);
nor U12655 (N_12655,N_11774,N_8435);
and U12656 (N_12656,N_11520,N_11787);
nand U12657 (N_12657,N_11697,N_10477);
nor U12658 (N_12658,N_11425,N_9511);
nand U12659 (N_12659,N_9780,N_7091);
and U12660 (N_12660,N_12184,N_8990);
or U12661 (N_12661,N_8296,N_7129);
nand U12662 (N_12662,N_10607,N_9807);
and U12663 (N_12663,N_8108,N_7454);
or U12664 (N_12664,N_9997,N_10880);
and U12665 (N_12665,N_9979,N_11401);
nor U12666 (N_12666,N_8073,N_6744);
or U12667 (N_12667,N_11020,N_8761);
nand U12668 (N_12668,N_8071,N_9167);
or U12669 (N_12669,N_9207,N_7771);
or U12670 (N_12670,N_7663,N_11816);
and U12671 (N_12671,N_12207,N_12155);
nand U12672 (N_12672,N_6777,N_9204);
or U12673 (N_12673,N_10839,N_8253);
nor U12674 (N_12674,N_10778,N_8302);
or U12675 (N_12675,N_9987,N_12177);
nor U12676 (N_12676,N_10797,N_8934);
or U12677 (N_12677,N_6252,N_11897);
and U12678 (N_12678,N_9513,N_8960);
nand U12679 (N_12679,N_7340,N_7498);
nor U12680 (N_12680,N_8667,N_8594);
and U12681 (N_12681,N_10186,N_8864);
nor U12682 (N_12682,N_6334,N_9198);
nand U12683 (N_12683,N_6500,N_9903);
or U12684 (N_12684,N_8796,N_11331);
or U12685 (N_12685,N_9349,N_7078);
or U12686 (N_12686,N_7341,N_8013);
nor U12687 (N_12687,N_11461,N_6788);
nor U12688 (N_12688,N_9876,N_8843);
nor U12689 (N_12689,N_7715,N_11702);
nand U12690 (N_12690,N_7896,N_9197);
and U12691 (N_12691,N_6508,N_7549);
and U12692 (N_12692,N_8219,N_7144);
or U12693 (N_12693,N_9000,N_12056);
or U12694 (N_12694,N_12308,N_8227);
and U12695 (N_12695,N_7582,N_6475);
nand U12696 (N_12696,N_11366,N_9599);
and U12697 (N_12697,N_9245,N_11081);
nor U12698 (N_12698,N_12091,N_9311);
nand U12699 (N_12699,N_12108,N_6940);
and U12700 (N_12700,N_10270,N_9827);
and U12701 (N_12701,N_11398,N_11271);
nor U12702 (N_12702,N_10020,N_10902);
nor U12703 (N_12703,N_8479,N_9925);
nand U12704 (N_12704,N_9555,N_9624);
xor U12705 (N_12705,N_8362,N_10420);
nand U12706 (N_12706,N_9019,N_8121);
nor U12707 (N_12707,N_9283,N_12080);
nor U12708 (N_12708,N_7476,N_7471);
and U12709 (N_12709,N_11307,N_6368);
or U12710 (N_12710,N_9710,N_11118);
xnor U12711 (N_12711,N_8804,N_8169);
or U12712 (N_12712,N_12479,N_9474);
nor U12713 (N_12713,N_8188,N_7934);
nand U12714 (N_12714,N_10854,N_12366);
nand U12715 (N_12715,N_6550,N_12264);
and U12716 (N_12716,N_11869,N_6586);
nor U12717 (N_12717,N_11657,N_9022);
and U12718 (N_12718,N_8292,N_10453);
or U12719 (N_12719,N_9446,N_6570);
nor U12720 (N_12720,N_7105,N_6734);
nor U12721 (N_12721,N_10027,N_10909);
nand U12722 (N_12722,N_11388,N_10634);
and U12723 (N_12723,N_9079,N_12162);
and U12724 (N_12724,N_7677,N_8705);
nand U12725 (N_12725,N_6440,N_7455);
or U12726 (N_12726,N_7994,N_8235);
or U12727 (N_12727,N_7770,N_7878);
xor U12728 (N_12728,N_10941,N_7038);
or U12729 (N_12729,N_10781,N_6863);
and U12730 (N_12730,N_9802,N_10390);
and U12731 (N_12731,N_8966,N_10345);
xor U12732 (N_12732,N_8712,N_8337);
nor U12733 (N_12733,N_10523,N_12231);
nand U12734 (N_12734,N_12383,N_9307);
nand U12735 (N_12735,N_6927,N_11727);
and U12736 (N_12736,N_10671,N_10196);
nand U12737 (N_12737,N_10260,N_9141);
and U12738 (N_12738,N_8033,N_9380);
nor U12739 (N_12739,N_10684,N_9905);
or U12740 (N_12740,N_11039,N_12224);
nor U12741 (N_12741,N_12057,N_6254);
or U12742 (N_12742,N_12440,N_11714);
or U12743 (N_12743,N_10809,N_6280);
nand U12744 (N_12744,N_6604,N_12168);
and U12745 (N_12745,N_6370,N_7185);
and U12746 (N_12746,N_11753,N_9456);
and U12747 (N_12747,N_10220,N_9427);
and U12748 (N_12748,N_9842,N_11370);
nand U12749 (N_12749,N_9159,N_8461);
nand U12750 (N_12750,N_12093,N_10400);
nand U12751 (N_12751,N_7623,N_11834);
and U12752 (N_12752,N_7673,N_9926);
and U12753 (N_12753,N_8240,N_8257);
nor U12754 (N_12754,N_10088,N_10614);
nor U12755 (N_12755,N_8282,N_9093);
or U12756 (N_12756,N_11134,N_8223);
or U12757 (N_12757,N_8999,N_9772);
nand U12758 (N_12758,N_10030,N_8626);
nor U12759 (N_12759,N_11561,N_7618);
nor U12760 (N_12760,N_8772,N_6873);
nand U12761 (N_12761,N_9350,N_7537);
or U12762 (N_12762,N_7230,N_10859);
nand U12763 (N_12763,N_11531,N_8773);
nor U12764 (N_12764,N_7087,N_7339);
and U12765 (N_12765,N_9039,N_9065);
or U12766 (N_12766,N_8480,N_7086);
or U12767 (N_12767,N_9629,N_12174);
and U12768 (N_12768,N_11462,N_8940);
and U12769 (N_12769,N_9316,N_10406);
and U12770 (N_12770,N_12215,N_9450);
or U12771 (N_12771,N_12315,N_10016);
and U12772 (N_12772,N_7342,N_12267);
and U12773 (N_12773,N_7565,N_6795);
nand U12774 (N_12774,N_9270,N_10603);
xnor U12775 (N_12775,N_9447,N_7903);
nand U12776 (N_12776,N_9028,N_7372);
nor U12777 (N_12777,N_7167,N_9187);
and U12778 (N_12778,N_11999,N_8231);
and U12779 (N_12779,N_8403,N_11945);
nor U12780 (N_12780,N_9354,N_8086);
nand U12781 (N_12781,N_6569,N_9542);
nor U12782 (N_12782,N_9692,N_7330);
and U12783 (N_12783,N_11339,N_8320);
nand U12784 (N_12784,N_8920,N_10365);
nand U12785 (N_12785,N_7158,N_11394);
nand U12786 (N_12786,N_10461,N_9011);
or U12787 (N_12787,N_10571,N_9586);
or U12788 (N_12788,N_8588,N_11078);
nor U12789 (N_12789,N_7765,N_10372);
xor U12790 (N_12790,N_9889,N_6561);
nand U12791 (N_12791,N_6427,N_8612);
nand U12792 (N_12792,N_9382,N_7984);
nand U12793 (N_12793,N_8853,N_12166);
or U12794 (N_12794,N_6938,N_10041);
nand U12795 (N_12795,N_9801,N_10548);
nand U12796 (N_12796,N_7874,N_9649);
xor U12797 (N_12797,N_10281,N_11255);
or U12798 (N_12798,N_10950,N_9519);
nor U12799 (N_12799,N_9571,N_6853);
nor U12800 (N_12800,N_7197,N_11547);
nor U12801 (N_12801,N_12367,N_10207);
nand U12802 (N_12802,N_8275,N_7234);
nand U12803 (N_12803,N_9041,N_10808);
nand U12804 (N_12804,N_10163,N_7392);
nand U12805 (N_12805,N_10562,N_6536);
and U12806 (N_12806,N_11976,N_6292);
nand U12807 (N_12807,N_11682,N_11319);
nand U12808 (N_12808,N_9874,N_11350);
xnor U12809 (N_12809,N_9305,N_9901);
or U12810 (N_12810,N_7047,N_9583);
nand U12811 (N_12811,N_8683,N_7865);
nand U12812 (N_12812,N_7683,N_8813);
nor U12813 (N_12813,N_12157,N_11076);
or U12814 (N_12814,N_12400,N_10681);
nor U12815 (N_12815,N_10071,N_8104);
and U12816 (N_12816,N_10544,N_12134);
nor U12817 (N_12817,N_12328,N_6556);
and U12818 (N_12818,N_8707,N_7360);
or U12819 (N_12819,N_7605,N_8448);
nand U12820 (N_12820,N_11323,N_9239);
or U12821 (N_12821,N_12273,N_9385);
nand U12822 (N_12822,N_8161,N_7682);
nor U12823 (N_12823,N_10028,N_12299);
nand U12824 (N_12824,N_11433,N_8618);
and U12825 (N_12825,N_7220,N_7408);
nor U12826 (N_12826,N_12284,N_8420);
nand U12827 (N_12827,N_7398,N_8144);
and U12828 (N_12828,N_12279,N_11848);
or U12829 (N_12829,N_9054,N_11918);
xor U12830 (N_12830,N_7556,N_12278);
nand U12831 (N_12831,N_11120,N_7976);
nor U12832 (N_12832,N_10683,N_10226);
nor U12833 (N_12833,N_10098,N_8038);
xnor U12834 (N_12834,N_7469,N_10458);
and U12835 (N_12835,N_7259,N_9091);
nor U12836 (N_12836,N_12104,N_10328);
nand U12837 (N_12837,N_7998,N_12132);
and U12838 (N_12838,N_9982,N_11431);
and U12839 (N_12839,N_8535,N_9670);
and U12840 (N_12840,N_9192,N_7089);
nand U12841 (N_12841,N_9002,N_11742);
nor U12842 (N_12842,N_11658,N_9396);
nor U12843 (N_12843,N_10120,N_12498);
or U12844 (N_12844,N_7875,N_8488);
nor U12845 (N_12845,N_8779,N_11932);
nor U12846 (N_12846,N_12237,N_8694);
nor U12847 (N_12847,N_9128,N_8276);
nor U12848 (N_12848,N_9561,N_7162);
nand U12849 (N_12849,N_6714,N_11173);
and U12850 (N_12850,N_11625,N_12409);
nor U12851 (N_12851,N_10796,N_8316);
nand U12852 (N_12852,N_10802,N_11971);
nor U12853 (N_12853,N_9379,N_6882);
or U12854 (N_12854,N_7665,N_8000);
nor U12855 (N_12855,N_12357,N_9704);
or U12856 (N_12856,N_11664,N_8870);
nand U12857 (N_12857,N_10875,N_6912);
nor U12858 (N_12858,N_10405,N_9588);
nor U12859 (N_12859,N_7418,N_11813);
and U12860 (N_12860,N_9071,N_11963);
xor U12861 (N_12861,N_8128,N_9407);
nor U12862 (N_12862,N_8841,N_8019);
or U12863 (N_12863,N_10656,N_9698);
nor U12864 (N_12864,N_8645,N_6408);
or U12865 (N_12865,N_10636,N_11357);
nand U12866 (N_12866,N_8604,N_12426);
nor U12867 (N_12867,N_7391,N_11991);
nand U12868 (N_12868,N_11231,N_6485);
nand U12869 (N_12869,N_11384,N_11227);
nand U12870 (N_12870,N_12223,N_10990);
and U12871 (N_12871,N_10732,N_8236);
nand U12872 (N_12872,N_9040,N_10706);
or U12873 (N_12873,N_11387,N_9709);
nand U12874 (N_12874,N_6746,N_10689);
nor U12875 (N_12875,N_10900,N_9340);
or U12876 (N_12876,N_7786,N_7907);
nor U12877 (N_12877,N_11894,N_9824);
nor U12878 (N_12878,N_11659,N_8742);
or U12879 (N_12879,N_11735,N_11652);
and U12880 (N_12880,N_11011,N_11094);
and U12881 (N_12881,N_6305,N_7241);
nor U12882 (N_12882,N_7366,N_7505);
nand U12883 (N_12883,N_6354,N_11484);
nor U12884 (N_12884,N_8392,N_9165);
nor U12885 (N_12885,N_7400,N_11044);
and U12886 (N_12886,N_10767,N_9492);
and U12887 (N_12887,N_10530,N_10630);
nor U12888 (N_12888,N_8595,N_7237);
or U12889 (N_12889,N_9421,N_7045);
or U12890 (N_12890,N_8196,N_9875);
nand U12891 (N_12891,N_9715,N_12476);
nand U12892 (N_12892,N_12487,N_11599);
and U12893 (N_12893,N_6648,N_11511);
nand U12894 (N_12894,N_11465,N_11435);
or U12895 (N_12895,N_12301,N_6640);
and U12896 (N_12896,N_10230,N_8965);
and U12897 (N_12897,N_7076,N_6548);
nor U12898 (N_12898,N_10653,N_6486);
nand U12899 (N_12899,N_8159,N_11089);
xnor U12900 (N_12900,N_7531,N_9904);
or U12901 (N_12901,N_7920,N_11084);
nor U12902 (N_12902,N_9540,N_10657);
nand U12903 (N_12903,N_9417,N_8786);
or U12904 (N_12904,N_8358,N_9983);
nand U12905 (N_12905,N_10890,N_6607);
or U12906 (N_12906,N_11494,N_9989);
and U12907 (N_12907,N_9856,N_6635);
nand U12908 (N_12908,N_9254,N_9746);
or U12909 (N_12909,N_11614,N_7561);
nand U12910 (N_12910,N_6403,N_11905);
or U12911 (N_12911,N_11310,N_6865);
nand U12912 (N_12912,N_6487,N_6884);
or U12913 (N_12913,N_8556,N_6818);
nand U12914 (N_12914,N_6299,N_12130);
nor U12915 (N_12915,N_7664,N_10306);
xor U12916 (N_12916,N_8497,N_12466);
and U12917 (N_12917,N_7603,N_11931);
and U12918 (N_12918,N_8330,N_7138);
nor U12919 (N_12919,N_6941,N_7141);
and U12920 (N_12920,N_12407,N_6609);
and U12921 (N_12921,N_8902,N_8765);
and U12922 (N_12922,N_6285,N_10976);
nor U12923 (N_12923,N_7914,N_10963);
and U12924 (N_12924,N_7810,N_7935);
xor U12925 (N_12925,N_6702,N_9587);
or U12926 (N_12926,N_7217,N_8539);
nor U12927 (N_12927,N_10275,N_11995);
nand U12928 (N_12928,N_12478,N_7169);
nand U12929 (N_12929,N_8312,N_9836);
nand U12930 (N_12930,N_9858,N_10515);
nor U12931 (N_12931,N_9635,N_6456);
or U12932 (N_12932,N_9654,N_8289);
nand U12933 (N_12933,N_10487,N_7503);
nand U12934 (N_12934,N_7337,N_9366);
xnor U12935 (N_12935,N_7371,N_8964);
or U12936 (N_12936,N_7216,N_6530);
nand U12937 (N_12937,N_6498,N_9318);
or U12938 (N_12938,N_8037,N_11422);
or U12939 (N_12939,N_7578,N_8143);
nor U12940 (N_12940,N_8284,N_8268);
nor U12941 (N_12941,N_7140,N_11156);
or U12942 (N_12942,N_8344,N_11391);
or U12943 (N_12943,N_8541,N_10033);
nand U12944 (N_12944,N_8098,N_11167);
nand U12945 (N_12945,N_10652,N_10244);
nand U12946 (N_12946,N_8768,N_10521);
nand U12947 (N_12947,N_7739,N_10058);
nand U12948 (N_12948,N_6274,N_11300);
or U12949 (N_12949,N_8536,N_9809);
xnor U12950 (N_12950,N_10253,N_11928);
and U12951 (N_12951,N_7879,N_11259);
nor U12952 (N_12952,N_7598,N_11042);
nor U12953 (N_12953,N_10946,N_7426);
or U12954 (N_12954,N_7160,N_8346);
nor U12955 (N_12955,N_7807,N_12051);
nand U12956 (N_12956,N_9943,N_8162);
nor U12957 (N_12957,N_8054,N_12396);
nor U12958 (N_12958,N_7316,N_9310);
or U12959 (N_12959,N_11597,N_10510);
nor U12960 (N_12960,N_10188,N_10715);
and U12961 (N_12961,N_6693,N_9515);
nand U12962 (N_12962,N_10171,N_6494);
xor U12963 (N_12963,N_9430,N_9449);
and U12964 (N_12964,N_8814,N_11601);
nor U12965 (N_12965,N_11284,N_9063);
nand U12966 (N_12966,N_10137,N_10309);
nor U12967 (N_12967,N_6303,N_7423);
nand U12968 (N_12968,N_6711,N_8122);
and U12969 (N_12969,N_10367,N_10308);
nand U12970 (N_12970,N_11047,N_6908);
or U12971 (N_12971,N_8295,N_11279);
and U12972 (N_12972,N_10125,N_10668);
nand U12973 (N_12973,N_8905,N_9974);
nor U12974 (N_12974,N_7075,N_11872);
and U12975 (N_12975,N_7861,N_8774);
nor U12976 (N_12976,N_8518,N_10516);
nand U12977 (N_12977,N_7497,N_7858);
nand U12978 (N_12978,N_11616,N_8191);
nor U12979 (N_12979,N_9778,N_8373);
xnor U12980 (N_12980,N_12246,N_7749);
nand U12981 (N_12981,N_8288,N_9848);
or U12982 (N_12982,N_6690,N_7152);
xor U12983 (N_12983,N_6890,N_9415);
and U12984 (N_12984,N_7460,N_8551);
nand U12985 (N_12985,N_12336,N_6339);
and U12986 (N_12986,N_8001,N_9945);
or U12987 (N_12987,N_11192,N_8918);
nor U12988 (N_12988,N_8656,N_7612);
nor U12989 (N_12989,N_12238,N_6328);
and U12990 (N_12990,N_10432,N_8688);
or U12991 (N_12991,N_10853,N_11062);
xnor U12992 (N_12992,N_10378,N_10182);
and U12993 (N_12993,N_6533,N_7209);
and U12994 (N_12994,N_11961,N_9570);
or U12995 (N_12995,N_7628,N_9553);
or U12996 (N_12996,N_11233,N_6834);
nand U12997 (N_12997,N_9672,N_8405);
and U12998 (N_12998,N_12280,N_12033);
xnor U12999 (N_12999,N_10380,N_9200);
nor U13000 (N_13000,N_8771,N_10788);
nor U13001 (N_13001,N_8102,N_8428);
and U13002 (N_13002,N_7074,N_11032);
and U13003 (N_13003,N_8904,N_7122);
and U13004 (N_13004,N_6910,N_8570);
nand U13005 (N_13005,N_8022,N_11543);
and U13006 (N_13006,N_7344,N_10324);
nand U13007 (N_13007,N_10654,N_8600);
nor U13008 (N_13008,N_9359,N_11794);
nor U13009 (N_13009,N_11215,N_8675);
nand U13010 (N_13010,N_12100,N_8599);
or U13011 (N_13011,N_7975,N_11882);
nand U13012 (N_13012,N_9600,N_9590);
or U13013 (N_13013,N_7702,N_7928);
nor U13014 (N_13014,N_6265,N_9510);
nor U13015 (N_13015,N_6256,N_12454);
and U13016 (N_13016,N_7778,N_9249);
nand U13017 (N_13017,N_10228,N_10001);
and U13018 (N_13018,N_6519,N_8897);
xor U13019 (N_13019,N_7432,N_11559);
or U13020 (N_13020,N_6849,N_11059);
or U13021 (N_13021,N_6646,N_8725);
nor U13022 (N_13022,N_8752,N_8631);
or U13023 (N_13023,N_6988,N_10736);
and U13024 (N_13024,N_11236,N_8024);
nor U13025 (N_13025,N_6759,N_8875);
nor U13026 (N_13026,N_9279,N_11311);
nor U13027 (N_13027,N_8134,N_8715);
and U13028 (N_13028,N_11238,N_9678);
xnor U13029 (N_13029,N_9367,N_7627);
or U13030 (N_13030,N_8261,N_7062);
xor U13031 (N_13031,N_12042,N_9508);
or U13032 (N_13032,N_11157,N_6923);
nand U13033 (N_13033,N_12311,N_8802);
nor U13034 (N_13034,N_7610,N_11630);
and U13035 (N_13035,N_8800,N_11407);
nand U13036 (N_13036,N_6700,N_11103);
or U13037 (N_13037,N_11557,N_10723);
nor U13038 (N_13038,N_7676,N_7056);
nor U13039 (N_13039,N_7215,N_9639);
and U13040 (N_13040,N_10731,N_12183);
and U13041 (N_13041,N_8424,N_10874);
or U13042 (N_13042,N_8690,N_8265);
and U13043 (N_13043,N_9917,N_10801);
xor U13044 (N_13044,N_7938,N_6659);
nor U13045 (N_13045,N_8972,N_6316);
nor U13046 (N_13046,N_7159,N_8821);
nand U13047 (N_13047,N_6482,N_6342);
or U13048 (N_13048,N_8294,N_12252);
and U13049 (N_13049,N_12142,N_9835);
xor U13050 (N_13050,N_6879,N_11591);
or U13051 (N_13051,N_11954,N_11676);
nor U13052 (N_13052,N_9924,N_9468);
nand U13053 (N_13053,N_10936,N_10419);
nand U13054 (N_13054,N_10957,N_9595);
nand U13055 (N_13055,N_12034,N_10059);
nor U13056 (N_13056,N_7801,N_10785);
or U13057 (N_13057,N_8971,N_7500);
nand U13058 (N_13058,N_8281,N_6804);
and U13059 (N_13059,N_10701,N_12074);
and U13060 (N_13060,N_8861,N_8482);
or U13061 (N_13061,N_7592,N_11396);
or U13062 (N_13062,N_8568,N_9263);
and U13063 (N_13063,N_7918,N_9477);
and U13064 (N_13064,N_12327,N_9505);
xor U13065 (N_13065,N_8140,N_6517);
nor U13066 (N_13066,N_8082,N_10979);
or U13067 (N_13067,N_8005,N_12325);
or U13068 (N_13068,N_11330,N_6445);
nand U13069 (N_13069,N_11606,N_12355);
or U13070 (N_13070,N_8200,N_11245);
nor U13071 (N_13071,N_9406,N_10503);
or U13072 (N_13072,N_6404,N_10482);
xnor U13073 (N_13073,N_12119,N_6600);
nor U13074 (N_13074,N_9643,N_7059);
or U13075 (N_13075,N_8232,N_7524);
nor U13076 (N_13076,N_6939,N_7973);
nand U13077 (N_13077,N_12024,N_12123);
or U13078 (N_13078,N_11124,N_11959);
nor U13079 (N_13079,N_12111,N_7965);
nand U13080 (N_13080,N_9258,N_7743);
or U13081 (N_13081,N_10827,N_6840);
xnor U13082 (N_13082,N_6450,N_12342);
and U13083 (N_13083,N_6534,N_9716);
or U13084 (N_13084,N_7964,N_10189);
and U13085 (N_13085,N_11612,N_9742);
and U13086 (N_13086,N_6341,N_11924);
or U13087 (N_13087,N_7369,N_9615);
nand U13088 (N_13088,N_11035,N_6833);
nand U13089 (N_13089,N_11734,N_11796);
or U13090 (N_13090,N_11509,N_7950);
and U13091 (N_13091,N_10143,N_6758);
and U13092 (N_13092,N_9864,N_8021);
or U13093 (N_13093,N_8212,N_9936);
nor U13094 (N_13094,N_10597,N_7651);
nor U13095 (N_13095,N_11501,N_9206);
nand U13096 (N_13096,N_10745,N_9865);
nor U13097 (N_13097,N_10089,N_11950);
and U13098 (N_13098,N_8913,N_10465);
and U13099 (N_13099,N_7235,N_11194);
nand U13100 (N_13100,N_7252,N_7039);
and U13101 (N_13101,N_11418,N_9286);
nor U13102 (N_13102,N_11269,N_9284);
xnor U13103 (N_13103,N_6599,N_9910);
or U13104 (N_13104,N_6728,N_11978);
or U13105 (N_13105,N_8815,N_12485);
nor U13106 (N_13106,N_9923,N_8978);
and U13107 (N_13107,N_12185,N_9358);
or U13108 (N_13108,N_6918,N_6617);
xor U13109 (N_13109,N_6660,N_8311);
xor U13110 (N_13110,N_8233,N_6822);
nand U13111 (N_13111,N_10357,N_7293);
nand U13112 (N_13112,N_8566,N_10794);
or U13113 (N_13113,N_11251,N_7750);
nand U13114 (N_13114,N_11282,N_7297);
nor U13115 (N_13115,N_6806,N_10444);
xnor U13116 (N_13116,N_10968,N_9500);
xnor U13117 (N_13117,N_11438,N_9955);
nand U13118 (N_13118,N_6410,N_9816);
nor U13119 (N_13119,N_8049,N_6459);
nor U13120 (N_13120,N_9804,N_6351);
and U13121 (N_13121,N_9662,N_7014);
nor U13122 (N_13122,N_9375,N_6881);
xor U13123 (N_13123,N_7978,N_7573);
or U13124 (N_13124,N_9666,N_10212);
or U13125 (N_13125,N_8579,N_11180);
xnor U13126 (N_13126,N_9617,N_8854);
and U13127 (N_13127,N_8522,N_10205);
and U13128 (N_13128,N_7792,N_7178);
nand U13129 (N_13129,N_12241,N_8446);
and U13130 (N_13130,N_11525,N_10006);
xor U13131 (N_13131,N_7856,N_11353);
or U13132 (N_13132,N_8438,N_8856);
nor U13133 (N_13133,N_10855,N_8666);
and U13134 (N_13134,N_7814,N_10296);
or U13135 (N_13135,N_8400,N_8164);
or U13136 (N_13136,N_7839,N_12265);
nand U13137 (N_13137,N_8943,N_7917);
or U13138 (N_13138,N_10312,N_6675);
and U13139 (N_13139,N_10851,N_8510);
and U13140 (N_13140,N_8034,N_8090);
or U13141 (N_13141,N_8863,N_6545);
and U13142 (N_13142,N_7101,N_10920);
and U13143 (N_13143,N_10416,N_7602);
or U13144 (N_13144,N_11771,N_10046);
xor U13145 (N_13145,N_6616,N_7669);
and U13146 (N_13146,N_11739,N_7272);
nand U13147 (N_13147,N_11449,N_12002);
and U13148 (N_13148,N_6914,N_11104);
nor U13149 (N_13149,N_12167,N_12110);
xor U13150 (N_13150,N_10532,N_12020);
nand U13151 (N_13151,N_6364,N_12014);
and U13152 (N_13152,N_9321,N_10966);
or U13153 (N_13153,N_8349,N_10231);
nand U13154 (N_13154,N_9527,N_11964);
and U13155 (N_13155,N_7442,N_6346);
nor U13156 (N_13156,N_9361,N_9413);
nor U13157 (N_13157,N_8153,N_8989);
nand U13158 (N_13158,N_11321,N_12410);
nand U13159 (N_13159,N_8529,N_9660);
nand U13160 (N_13160,N_7103,N_11554);
or U13161 (N_13161,N_7630,N_10539);
nor U13162 (N_13162,N_7633,N_12258);
and U13163 (N_13163,N_9798,N_12482);
nor U13164 (N_13164,N_11055,N_6778);
and U13165 (N_13165,N_9828,N_9191);
nor U13166 (N_13166,N_9657,N_8189);
xor U13167 (N_13167,N_9580,N_10560);
xnor U13168 (N_13168,N_6499,N_12199);
or U13169 (N_13169,N_7294,N_8309);
and U13170 (N_13170,N_9053,N_11286);
or U13171 (N_13171,N_8669,N_11814);
and U13172 (N_13172,N_11646,N_9362);
xnor U13173 (N_13173,N_10629,N_7980);
and U13174 (N_13174,N_11772,N_6898);
xor U13175 (N_13175,N_7326,N_6708);
nand U13176 (N_13176,N_11653,N_6580);
xnor U13177 (N_13177,N_12424,N_7006);
nor U13178 (N_13178,N_11143,N_11548);
nand U13179 (N_13179,N_9212,N_11631);
nor U13180 (N_13180,N_10339,N_10691);
or U13181 (N_13181,N_12154,N_11113);
or U13182 (N_13182,N_12124,N_11718);
or U13183 (N_13183,N_10138,N_10782);
nor U13184 (N_13184,N_7113,N_6284);
or U13185 (N_13185,N_7414,N_8347);
nor U13186 (N_13186,N_9490,N_6987);
nand U13187 (N_13187,N_10729,N_6541);
nand U13188 (N_13188,N_6824,N_9922);
and U13189 (N_13189,N_10133,N_8561);
nor U13190 (N_13190,N_11807,N_8895);
xnor U13191 (N_13191,N_10100,N_7381);
nand U13192 (N_13192,N_11539,N_7639);
nor U13193 (N_13193,N_7021,N_9029);
and U13194 (N_13194,N_12209,N_6794);
nand U13195 (N_13195,N_7845,N_10437);
and U13196 (N_13196,N_10329,N_9566);
nor U13197 (N_13197,N_8372,N_7620);
and U13198 (N_13198,N_7824,N_8736);
or U13199 (N_13199,N_8374,N_7795);
xnor U13200 (N_13200,N_9965,N_12144);
or U13201 (N_13201,N_9155,N_7788);
or U13202 (N_13202,N_11679,N_10402);
nand U13203 (N_13203,N_6842,N_12362);
and U13204 (N_13204,N_10847,N_8426);
and U13205 (N_13205,N_11201,N_7846);
nor U13206 (N_13206,N_10619,N_9403);
nor U13207 (N_13207,N_12102,N_9188);
or U13208 (N_13208,N_8589,N_6762);
nand U13209 (N_13209,N_7567,N_11674);
nand U13210 (N_13210,N_9723,N_9058);
or U13211 (N_13211,N_7745,N_6729);
nand U13212 (N_13212,N_8925,N_10087);
xor U13213 (N_13213,N_10083,N_8723);
and U13214 (N_13214,N_8496,N_8941);
nand U13215 (N_13215,N_8171,N_7443);
xnor U13216 (N_13216,N_10857,N_11638);
and U13217 (N_13217,N_9495,N_6817);
nand U13218 (N_13218,N_11996,N_11629);
nand U13219 (N_13219,N_9517,N_6955);
and U13220 (N_13220,N_8201,N_10427);
nor U13221 (N_13221,N_6811,N_8544);
nand U13222 (N_13222,N_8910,N_8676);
nand U13223 (N_13223,N_8381,N_12276);
or U13224 (N_13224,N_7026,N_7389);
nand U13225 (N_13225,N_11648,N_11949);
xnor U13226 (N_13226,N_10074,N_12012);
and U13227 (N_13227,N_7174,N_10463);
and U13228 (N_13228,N_10867,N_10775);
and U13229 (N_13229,N_12349,N_6666);
and U13230 (N_13230,N_8930,N_6730);
nand U13231 (N_13231,N_10099,N_9815);
and U13232 (N_13232,N_9006,N_7656);
xnor U13233 (N_13233,N_7301,N_11555);
nand U13234 (N_13234,N_7143,N_6812);
nand U13235 (N_13235,N_10881,N_8871);
or U13236 (N_13236,N_12353,N_8124);
nor U13237 (N_13237,N_12081,N_9080);
nor U13238 (N_13238,N_11220,N_9478);
nor U13239 (N_13239,N_7177,N_8525);
nand U13240 (N_13240,N_12391,N_6613);
or U13241 (N_13241,N_9329,N_9652);
and U13242 (N_13242,N_8702,N_9946);
nor U13243 (N_13243,N_9202,N_12442);
and U13244 (N_13244,N_10386,N_8413);
and U13245 (N_13245,N_11598,N_7805);
or U13246 (N_13246,N_12483,N_8078);
nand U13247 (N_13247,N_6420,N_11294);
nor U13248 (N_13248,N_12392,N_7002);
or U13249 (N_13249,N_6261,N_9213);
nand U13250 (N_13250,N_6654,N_9701);
nand U13251 (N_13251,N_12416,N_9256);
and U13252 (N_13252,N_10269,N_9738);
nor U13253 (N_13253,N_7401,N_10919);
nor U13254 (N_13254,N_10170,N_9509);
or U13255 (N_13255,N_7033,N_6979);
or U13256 (N_13256,N_10756,N_7179);
or U13257 (N_13257,N_11239,N_11188);
and U13258 (N_13258,N_7733,N_9576);
and U13259 (N_13259,N_7009,N_9309);
xor U13260 (N_13260,N_7886,N_7092);
and U13261 (N_13261,N_7876,N_10553);
and U13262 (N_13262,N_6395,N_10960);
or U13263 (N_13263,N_8247,N_6747);
nand U13264 (N_13264,N_11095,N_8301);
nor U13265 (N_13265,N_8641,N_11948);
and U13266 (N_13266,N_8043,N_6283);
nor U13267 (N_13267,N_7960,N_10566);
or U13268 (N_13268,N_7619,N_10905);
nand U13269 (N_13269,N_9633,N_9219);
or U13270 (N_13270,N_6703,N_11823);
or U13271 (N_13271,N_7483,N_9104);
nand U13272 (N_13272,N_8523,N_6752);
and U13273 (N_13273,N_8307,N_7527);
or U13274 (N_13274,N_11636,N_7962);
nor U13275 (N_13275,N_8578,N_7310);
nor U13276 (N_13276,N_10047,N_9404);
and U13277 (N_13277,N_9304,N_7591);
or U13278 (N_13278,N_10518,N_8067);
and U13279 (N_13279,N_6393,N_12028);
nand U13280 (N_13280,N_11274,N_11691);
and U13281 (N_13281,N_9111,N_12007);
or U13282 (N_13282,N_8035,N_8336);
nand U13283 (N_13283,N_11109,N_9373);
and U13284 (N_13284,N_11650,N_9050);
and U13285 (N_13285,N_11781,N_10724);
nor U13286 (N_13286,N_8516,N_9882);
xor U13287 (N_13287,N_12245,N_9169);
or U13288 (N_13288,N_9124,N_11510);
nand U13289 (N_13289,N_11016,N_9073);
or U13290 (N_13290,N_11859,N_8462);
nand U13291 (N_13291,N_12216,N_10878);
nand U13292 (N_13292,N_8701,N_7490);
nand U13293 (N_13293,N_9433,N_9869);
or U13294 (N_13294,N_6511,N_11364);
and U13295 (N_13295,N_11527,N_12382);
nor U13296 (N_13296,N_7632,N_7100);
or U13297 (N_13297,N_9240,N_7767);
xnor U13298 (N_13298,N_12445,N_9800);
and U13299 (N_13299,N_7256,N_8613);
and U13300 (N_13300,N_10287,N_10543);
nor U13301 (N_13301,N_7568,N_8787);
nand U13302 (N_13302,N_7127,N_9383);
or U13303 (N_13303,N_8687,N_9211);
nand U13304 (N_13304,N_8313,N_9290);
or U13305 (N_13305,N_7599,N_8650);
nor U13306 (N_13306,N_11850,N_7611);
nand U13307 (N_13307,N_9153,N_8452);
xor U13308 (N_13308,N_10301,N_7732);
nand U13309 (N_13309,N_11356,N_8534);
nor U13310 (N_13310,N_9573,N_6350);
and U13311 (N_13311,N_9374,N_11618);
xnor U13312 (N_13312,N_9810,N_7168);
nand U13313 (N_13313,N_8872,N_11345);
nand U13314 (N_13314,N_11835,N_7149);
nand U13315 (N_13315,N_9988,N_11252);
and U13316 (N_13316,N_6453,N_11556);
or U13317 (N_13317,N_7108,N_11135);
xor U13318 (N_13318,N_10039,N_10791);
and U13319 (N_13319,N_11822,N_8089);
or U13320 (N_13320,N_8512,N_12305);
xnor U13321 (N_13321,N_8503,N_7513);
and U13322 (N_13322,N_8339,N_6546);
or U13323 (N_13323,N_9247,N_6887);
nor U13324 (N_13324,N_9530,N_12289);
nor U13325 (N_13325,N_12052,N_9126);
or U13326 (N_13326,N_8209,N_6269);
nor U13327 (N_13327,N_6584,N_11746);
nand U13328 (N_13328,N_7948,N_7759);
nor U13329 (N_13329,N_10737,N_12447);
and U13330 (N_13330,N_8590,N_8803);
nor U13331 (N_13331,N_7584,N_8602);
nor U13332 (N_13332,N_8192,N_7533);
nand U13333 (N_13333,N_9538,N_11611);
and U13334 (N_13334,N_6643,N_8286);
and U13335 (N_13335,N_12272,N_9957);
and U13336 (N_13336,N_8831,N_9606);
or U13337 (N_13337,N_9663,N_7834);
nand U13338 (N_13338,N_12345,N_8799);
nor U13339 (N_13339,N_8758,N_12107);
and U13340 (N_13340,N_11375,N_6514);
xnor U13341 (N_13341,N_11729,N_7358);
nand U13342 (N_13342,N_11196,N_11840);
and U13343 (N_13343,N_9012,N_10967);
and U13344 (N_13344,N_11204,N_9017);
and U13345 (N_13345,N_8660,N_8975);
nor U13346 (N_13346,N_6323,N_10744);
nand U13347 (N_13347,N_7945,N_8992);
and U13348 (N_13348,N_9103,N_7117);
and U13349 (N_13349,N_8649,N_11666);
or U13350 (N_13350,N_12182,N_10823);
nand U13351 (N_13351,N_11593,N_9101);
or U13352 (N_13352,N_9085,N_8315);
and U13353 (N_13353,N_11979,N_9113);
or U13354 (N_13354,N_9143,N_10848);
nand U13355 (N_13355,N_7336,N_6973);
or U13356 (N_13356,N_6984,N_10505);
nand U13357 (N_13357,N_11363,N_10015);
nand U13358 (N_13358,N_7208,N_6845);
xnor U13359 (N_13359,N_7899,N_8291);
or U13360 (N_13360,N_10568,N_8747);
and U13361 (N_13361,N_10352,N_9830);
nand U13362 (N_13362,N_8834,N_9773);
xnor U13363 (N_13363,N_11589,N_10174);
nor U13364 (N_13364,N_8317,N_11187);
nor U13365 (N_13365,N_7203,N_11455);
xor U13366 (N_13366,N_7910,N_10971);
nor U13367 (N_13367,N_10672,N_9930);
xnor U13368 (N_13368,N_6789,N_8530);
and U13369 (N_13369,N_6773,N_7468);
and U13370 (N_13370,N_8132,N_9424);
and U13371 (N_13371,N_11804,N_8110);
nor U13372 (N_13372,N_9868,N_8889);
and U13373 (N_13373,N_9897,N_7184);
nand U13374 (N_13374,N_10822,N_12312);
or U13375 (N_13375,N_9276,N_10925);
nor U13376 (N_13376,N_7011,N_6807);
nor U13377 (N_13377,N_11692,N_9675);
nor U13378 (N_13378,N_8207,N_9440);
and U13379 (N_13379,N_11833,N_10079);
nand U13380 (N_13380,N_10564,N_10319);
nor U13381 (N_13381,N_10741,N_10825);
and U13382 (N_13382,N_10838,N_9001);
or U13383 (N_13383,N_11726,N_8837);
nand U13384 (N_13384,N_10768,N_9401);
nor U13385 (N_13385,N_11668,N_8783);
or U13386 (N_13386,N_7827,N_11451);
and U13387 (N_13387,N_6713,N_11985);
nor U13388 (N_13388,N_9646,N_7125);
xnor U13389 (N_13389,N_12180,N_12048);
or U13390 (N_13390,N_10779,N_6779);
and U13391 (N_13391,N_6872,N_7949);
xor U13392 (N_13392,N_11819,N_10563);
and U13393 (N_13393,N_8449,N_10155);
and U13394 (N_13394,N_8250,N_9049);
and U13395 (N_13395,N_7338,N_11662);
or U13396 (N_13396,N_10526,N_7485);
nand U13397 (N_13397,N_10141,N_8592);
and U13398 (N_13398,N_10930,N_11671);
xnor U13399 (N_13399,N_10468,N_9234);
nor U13400 (N_13400,N_12191,N_8117);
nor U13401 (N_13401,N_10486,N_12156);
nand U13402 (N_13402,N_11359,N_11492);
nand U13403 (N_13403,N_6799,N_12044);
nor U13404 (N_13404,N_7161,N_11161);
nor U13405 (N_13405,N_11003,N_9994);
nand U13406 (N_13406,N_6380,N_7595);
and U13407 (N_13407,N_6645,N_9448);
and U13408 (N_13408,N_9330,N_11355);
nor U13409 (N_13409,N_10673,N_11318);
nor U13410 (N_13410,N_11904,N_10820);
and U13411 (N_13411,N_8668,N_9089);
nand U13412 (N_13412,N_10556,N_10166);
or U13413 (N_13413,N_8477,N_7295);
and U13414 (N_13414,N_10592,N_11828);
nor U13415 (N_13415,N_6302,N_9556);
nand U13416 (N_13416,N_6419,N_9781);
nand U13417 (N_13417,N_10861,N_8412);
and U13418 (N_13418,N_9250,N_12170);
nand U13419 (N_13419,N_11477,N_8341);
nand U13420 (N_13420,N_8460,N_10666);
nor U13421 (N_13421,N_11056,N_10907);
and U13422 (N_13422,N_6471,N_8072);
and U13423 (N_13423,N_8002,N_11728);
and U13424 (N_13424,N_11825,N_8272);
xor U13425 (N_13425,N_12322,N_11123);
and U13426 (N_13426,N_12398,N_12036);
nand U13427 (N_13427,N_9272,N_9368);
and U13428 (N_13428,N_7034,N_9422);
nor U13429 (N_13429,N_6431,N_9112);
nor U13430 (N_13430,N_12288,N_10134);
nand U13431 (N_13431,N_7273,N_6748);
or U13432 (N_13432,N_10024,N_7357);
nand U13433 (N_13433,N_7799,N_8156);
nor U13434 (N_13434,N_11686,N_10121);
or U13435 (N_13435,N_12423,N_9339);
xnor U13436 (N_13436,N_7313,N_9156);
nand U13437 (N_13437,N_7835,N_10826);
nor U13438 (N_13438,N_9078,N_9575);
xor U13439 (N_13439,N_9533,N_10877);
or U13440 (N_13440,N_7941,N_8246);
or U13441 (N_13441,N_9466,N_10646);
xor U13442 (N_13442,N_9630,N_12371);
and U13443 (N_13443,N_9845,N_11857);
nor U13444 (N_13444,N_10215,N_8163);
or U13445 (N_13445,N_6531,N_8698);
nand U13446 (N_13446,N_9978,N_8494);
nor U13447 (N_13447,N_9770,N_9854);
and U13448 (N_13448,N_10102,N_12148);
nand U13449 (N_13449,N_7653,N_8700);
nand U13450 (N_13450,N_6425,N_9981);
or U13451 (N_13451,N_11065,N_7229);
or U13452 (N_13452,N_7521,N_6591);
nor U13453 (N_13453,N_10485,N_7951);
and U13454 (N_13454,N_11175,N_12137);
or U13455 (N_13455,N_10803,N_6264);
or U13456 (N_13456,N_11602,N_10730);
and U13457 (N_13457,N_10254,N_11913);
and U13458 (N_13458,N_10784,N_8050);
xnor U13459 (N_13459,N_11607,N_12160);
xnor U13460 (N_13460,N_8944,N_10858);
nand U13461 (N_13461,N_8909,N_11116);
or U13462 (N_13462,N_6847,N_8443);
and U13463 (N_13463,N_12084,N_11800);
nor U13464 (N_13464,N_8573,N_7031);
nand U13465 (N_13465,N_7115,N_7992);
or U13466 (N_13466,N_11622,N_11360);
nor U13467 (N_13467,N_8355,N_11875);
and U13468 (N_13468,N_9162,N_9669);
and U13469 (N_13469,N_7440,N_10922);
and U13470 (N_13470,N_9880,N_9293);
nand U13471 (N_13471,N_10752,N_9627);
and U13472 (N_13472,N_10494,N_10123);
and U13473 (N_13473,N_11420,N_6830);
nand U13474 (N_13474,N_8968,N_10509);
nand U13475 (N_13475,N_10986,N_8572);
nand U13476 (N_13476,N_6583,N_9271);
xnor U13477 (N_13477,N_11853,N_9451);
nor U13478 (N_13478,N_6357,N_12172);
nor U13479 (N_13479,N_7982,N_10399);
and U13480 (N_13480,N_9991,N_11214);
and U13481 (N_13481,N_8213,N_9133);
and U13482 (N_13482,N_6532,N_7254);
or U13483 (N_13483,N_8696,N_7095);
or U13484 (N_13484,N_9105,N_8995);
nand U13485 (N_13485,N_11393,N_6495);
nor U13486 (N_13486,N_8961,N_9969);
nand U13487 (N_13487,N_11460,N_7729);
nor U13488 (N_13488,N_9567,N_9488);
and U13489 (N_13489,N_7322,N_10814);
and U13490 (N_13490,N_8878,N_11756);
nor U13491 (N_13491,N_11329,N_10124);
nor U13492 (N_13492,N_6490,N_8119);
nor U13493 (N_13493,N_8951,N_6684);
nor U13494 (N_13494,N_8574,N_9944);
or U13495 (N_13495,N_10349,N_12009);
nor U13496 (N_13496,N_7487,N_8376);
or U13497 (N_13497,N_10981,N_11975);
nand U13498 (N_13498,N_6594,N_9786);
nand U13499 (N_13499,N_9759,N_9941);
and U13500 (N_13500,N_8520,N_9873);
xnor U13501 (N_13501,N_10200,N_6696);
and U13502 (N_13502,N_7311,N_7354);
nand U13503 (N_13503,N_7124,N_10488);
and U13504 (N_13504,N_11160,N_12256);
or U13505 (N_13505,N_11414,N_7700);
nor U13506 (N_13506,N_7233,N_8193);
and U13507 (N_13507,N_9962,N_9097);
nand U13508 (N_13508,N_10392,N_12126);
xor U13509 (N_13509,N_6437,N_12444);
and U13510 (N_13510,N_8453,N_9887);
and U13511 (N_13511,N_9458,N_11562);
nand U13512 (N_13512,N_8777,N_7564);
or U13513 (N_13513,N_8963,N_9363);
xor U13514 (N_13514,N_11342,N_9337);
or U13515 (N_13515,N_10846,N_7754);
nand U13516 (N_13516,N_10637,N_7331);
or U13517 (N_13517,N_10007,N_8532);
or U13518 (N_13518,N_8504,N_12329);
nor U13519 (N_13519,N_6481,N_7720);
nor U13520 (N_13520,N_6373,N_6528);
nand U13521 (N_13521,N_10204,N_7748);
nor U13522 (N_13522,N_9867,N_12159);
nor U13523 (N_13523,N_10280,N_10962);
or U13524 (N_13524,N_7554,N_7889);
or U13525 (N_13525,N_7866,N_6719);
xnor U13526 (N_13526,N_11665,N_11731);
and U13527 (N_13527,N_11797,N_9844);
and U13528 (N_13528,N_9948,N_10355);
nor U13529 (N_13529,N_10029,N_11149);
and U13530 (N_13530,N_9730,N_11754);
or U13531 (N_13531,N_10443,N_6526);
nor U13532 (N_13532,N_8798,N_9190);
or U13533 (N_13533,N_11349,N_8830);
or U13534 (N_13534,N_9544,N_12486);
nand U13535 (N_13535,N_10927,N_11021);
or U13536 (N_13536,N_8825,N_11027);
and U13537 (N_13537,N_7210,N_12099);
nand U13538 (N_13538,N_8531,N_10103);
nand U13539 (N_13539,N_8959,N_9431);
xnor U13540 (N_13540,N_8637,N_8478);
nor U13541 (N_13541,N_10710,N_8793);
and U13542 (N_13542,N_9631,N_9879);
or U13543 (N_13543,N_7692,N_9853);
or U13544 (N_13544,N_6816,N_7983);
and U13545 (N_13545,N_12380,N_9268);
nand U13546 (N_13546,N_7981,N_10926);
nor U13547 (N_13547,N_7853,N_7844);
and U13548 (N_13548,N_10886,N_11644);
nand U13549 (N_13549,N_6455,N_10262);
or U13550 (N_13550,N_9958,N_12058);
nand U13551 (N_13551,N_9523,N_11899);
nand U13552 (N_13552,N_12112,N_7512);
nand U13553 (N_13553,N_12286,N_7061);
nor U13554 (N_13554,N_8671,N_11240);
or U13555 (N_13555,N_8950,N_10842);
and U13556 (N_13556,N_7085,N_6383);
or U13557 (N_13557,N_9360,N_8063);
and U13558 (N_13558,N_6577,N_8404);
xor U13559 (N_13559,N_8585,N_9531);
and U13560 (N_13560,N_6467,N_9885);
nand U13561 (N_13561,N_10132,N_8826);
nor U13562 (N_13562,N_11478,N_12049);
nor U13563 (N_13563,N_9300,N_6651);
or U13564 (N_13564,N_11956,N_8896);
nor U13565 (N_13565,N_8241,N_10620);
nor U13566 (N_13566,N_9966,N_10197);
nand U13567 (N_13567,N_11289,N_8167);
and U13568 (N_13568,N_9487,N_7897);
xnor U13569 (N_13569,N_8202,N_10651);
or U13570 (N_13570,N_10602,N_11139);
nor U13571 (N_13571,N_7306,N_7131);
nor U13572 (N_13572,N_9658,N_7435);
or U13573 (N_13573,N_8464,N_11581);
nor U13574 (N_13574,N_11941,N_12307);
nor U13575 (N_13575,N_10830,N_12321);
xnor U13576 (N_13576,N_11847,N_11685);
xor U13577 (N_13577,N_10496,N_7409);
nand U13578 (N_13578,N_9411,N_11265);
xor U13579 (N_13579,N_9731,N_6916);
and U13580 (N_13580,N_11368,N_12255);
and U13581 (N_13581,N_7608,N_8775);
nor U13582 (N_13582,N_6396,N_7735);
xnor U13583 (N_13583,N_6275,N_7588);
nand U13584 (N_13584,N_6791,N_6787);
xnor U13585 (N_13585,N_8194,N_12213);
xnor U13586 (N_13586,N_7546,N_7437);
nor U13587 (N_13587,N_11246,N_6614);
and U13588 (N_13588,N_12062,N_10381);
and U13589 (N_13589,N_12384,N_9753);
xnor U13590 (N_13590,N_10423,N_11534);
and U13591 (N_13591,N_12105,N_7199);
nand U13592 (N_13592,N_9975,N_12316);
xnor U13593 (N_13593,N_12067,N_9236);
or U13594 (N_13594,N_11110,N_11040);
nor U13595 (N_13595,N_9481,N_11184);
or U13596 (N_13596,N_8629,N_11010);
or U13597 (N_13597,N_11324,N_11390);
nor U13598 (N_13598,N_9964,N_11812);
xnor U13599 (N_13599,N_8757,N_7626);
or U13600 (N_13600,N_8238,N_6889);
nand U13601 (N_13601,N_7183,N_12352);
and U13602 (N_13602,N_10806,N_7888);
or U13603 (N_13603,N_10003,N_12054);
nand U13604 (N_13604,N_6751,N_8596);
or U13605 (N_13605,N_9014,N_11695);
nor U13606 (N_13606,N_8789,N_8155);
nand U13607 (N_13607,N_8980,N_9840);
or U13608 (N_13608,N_10935,N_12401);
and U13609 (N_13609,N_8237,N_6780);
and U13610 (N_13610,N_10167,N_7987);
nor U13611 (N_13611,N_8273,N_8222);
and U13612 (N_13612,N_7016,N_7239);
nand U13613 (N_13613,N_6253,N_10605);
and U13614 (N_13614,N_7139,N_6619);
nand U13615 (N_13615,N_9118,N_8886);
or U13616 (N_13616,N_11837,N_8957);
xor U13617 (N_13617,N_6694,N_7363);
or U13618 (N_13618,N_8109,N_11827);
or U13619 (N_13619,N_7332,N_10394);
nor U13620 (N_13620,N_8801,N_7044);
nor U13621 (N_13621,N_6953,N_8094);
and U13622 (N_13622,N_7236,N_10733);
and U13623 (N_13623,N_6994,N_11481);
nand U13624 (N_13624,N_9116,N_6353);
and U13625 (N_13625,N_11502,N_6764);
nand U13626 (N_13626,N_12326,N_8224);
nand U13627 (N_13627,N_10685,N_11403);
nand U13628 (N_13628,N_12193,N_7974);
or U13629 (N_13629,N_8370,N_6388);
xnor U13630 (N_13630,N_11429,N_7728);
and U13631 (N_13631,N_8081,N_6438);
or U13632 (N_13632,N_10241,N_11408);
and U13633 (N_13633,N_8458,N_9823);
nor U13634 (N_13634,N_12227,N_8970);
and U13635 (N_13635,N_6484,N_9784);
nand U13636 (N_13636,N_9090,N_7659);
nand U13637 (N_13637,N_8481,N_9727);
or U13638 (N_13638,N_11106,N_9612);
or U13639 (N_13639,N_9779,N_10162);
nand U13640 (N_13640,N_8180,N_9724);
or U13641 (N_13641,N_6964,N_9389);
xnor U13642 (N_13642,N_6785,N_9076);
nor U13643 (N_13643,N_9163,N_9687);
nand U13644 (N_13644,N_6861,N_12068);
and U13645 (N_13645,N_10067,N_11009);
nor U13646 (N_13646,N_8216,N_8621);
and U13647 (N_13647,N_8378,N_9348);
and U13648 (N_13648,N_6413,N_6917);
and U13649 (N_13649,N_6281,N_8652);
or U13650 (N_13650,N_10892,N_12165);
nand U13651 (N_13651,N_8084,N_7395);
or U13652 (N_13652,N_9928,N_10446);
nor U13653 (N_13653,N_6776,N_11015);
nand U13654 (N_13654,N_6333,N_10433);
and U13655 (N_13655,N_6603,N_10415);
nand U13656 (N_13656,N_7121,N_12350);
nand U13657 (N_13657,N_11573,N_9094);
or U13658 (N_13658,N_8264,N_10628);
and U13659 (N_13659,N_7329,N_9394);
xnor U13660 (N_13660,N_10235,N_9603);
and U13661 (N_13661,N_11489,N_6473);
and U13662 (N_13662,N_11558,N_11655);
nor U13663 (N_13663,N_7406,N_10343);
and U13664 (N_13664,N_11203,N_6856);
nand U13665 (N_13665,N_9620,N_11376);
and U13666 (N_13666,N_10080,N_8447);
nand U13667 (N_13667,N_11953,N_12497);
xor U13668 (N_13668,N_6338,N_11333);
or U13669 (N_13669,N_7689,N_7507);
nor U13670 (N_13670,N_6470,N_8457);
nor U13671 (N_13671,N_12437,N_7721);
nand U13672 (N_13672,N_7650,N_12143);
nor U13673 (N_13673,N_7480,N_8350);
or U13674 (N_13674,N_8738,N_11624);
nand U13675 (N_13675,N_7961,N_7249);
and U13676 (N_13676,N_6966,N_9507);
or U13677 (N_13677,N_11463,N_12274);
nor U13678 (N_13678,N_12344,N_11456);
nand U13679 (N_13679,N_10816,N_10600);
nand U13680 (N_13680,N_8135,N_10032);
or U13681 (N_13681,N_6544,N_7849);
nor U13682 (N_13682,N_8695,N_10849);
and U13683 (N_13683,N_9420,N_6854);
nor U13684 (N_13684,N_7390,N_8025);
xnor U13685 (N_13685,N_6539,N_7712);
xnor U13686 (N_13686,N_7334,N_12356);
nor U13687 (N_13687,N_10835,N_9241);
nor U13688 (N_13688,N_7794,N_7266);
nor U13689 (N_13689,N_10678,N_10757);
or U13690 (N_13690,N_10403,N_8492);
nor U13691 (N_13691,N_8490,N_7997);
nand U13692 (N_13692,N_11574,N_8114);
or U13693 (N_13693,N_6836,N_10263);
or U13694 (N_13694,N_7018,N_7264);
xnor U13695 (N_13695,N_9961,N_7416);
and U13696 (N_13696,N_9036,N_8314);
or U13697 (N_13697,N_10680,N_10540);
xor U13698 (N_13698,N_9501,N_10665);
or U13699 (N_13699,N_9176,N_11871);
and U13700 (N_13700,N_7566,N_6883);
nand U13701 (N_13701,N_8879,N_6362);
xnor U13702 (N_13702,N_9909,N_8061);
and U13703 (N_13703,N_7394,N_6463);
nor U13704 (N_13704,N_8023,N_11908);
and U13705 (N_13705,N_11254,N_11280);
nor U13706 (N_13706,N_9502,N_7508);
or U13707 (N_13707,N_11079,N_7022);
nor U13708 (N_13708,N_11105,N_7300);
nand U13709 (N_13709,N_8862,N_8845);
xnor U13710 (N_13710,N_11958,N_6562);
xor U13711 (N_13711,N_10422,N_8141);
nor U13712 (N_13712,N_11965,N_6324);
nor U13713 (N_13713,N_7774,N_6503);
and U13714 (N_13714,N_12259,N_10868);
nand U13715 (N_13715,N_6523,N_8440);
nand U13716 (N_13716,N_6796,N_9525);
nand U13717 (N_13717,N_12197,N_11334);
or U13718 (N_13718,N_11900,N_11870);
nand U13719 (N_13719,N_10686,N_10031);
nor U13720 (N_13720,N_6258,N_6943);
nor U13721 (N_13721,N_7477,N_6657);
nand U13722 (N_13722,N_8682,N_6430);
xor U13723 (N_13723,N_11541,N_7283);
or U13724 (N_13724,N_10417,N_8858);
or U13725 (N_13725,N_9386,N_7456);
or U13726 (N_13726,N_7378,N_7991);
nand U13727 (N_13727,N_11936,N_11937);
nand U13728 (N_13728,N_9397,N_8657);
nor U13729 (N_13729,N_8327,N_6678);
and U13730 (N_13730,N_11434,N_12187);
nand U13731 (N_13731,N_8470,N_12277);
nor U13732 (N_13732,N_11778,N_12136);
and U13733 (N_13733,N_10844,N_6981);
or U13734 (N_13734,N_11766,N_7966);
nor U13735 (N_13735,N_12306,N_11565);
and U13736 (N_13736,N_7425,N_10298);
nand U13737 (N_13737,N_10789,N_7580);
nand U13738 (N_13738,N_10363,N_7224);
nand U13739 (N_13739,N_8105,N_12460);
or U13740 (N_13740,N_7270,N_7756);
and U13741 (N_13741,N_11545,N_10202);
nand U13742 (N_13742,N_10702,N_12334);
and U13743 (N_13743,N_8360,N_6911);
nand U13744 (N_13744,N_10489,N_8946);
or U13745 (N_13745,N_8507,N_8728);
and U13746 (N_13746,N_12491,N_6461);
and U13747 (N_13747,N_6452,N_12065);
or U13748 (N_13748,N_8397,N_10873);
nand U13749 (N_13749,N_11441,N_7859);
xnor U13750 (N_13750,N_9653,N_7488);
or U13751 (N_13751,N_11305,N_6626);
nand U13752 (N_13752,N_11775,N_10916);
nand U13753 (N_13753,N_9127,N_9266);
and U13754 (N_13754,N_8407,N_10704);
xor U13755 (N_13755,N_6720,N_9082);
nand U13756 (N_13756,N_11445,N_7867);
or U13757 (N_13757,N_11838,N_9109);
nand U13758 (N_13758,N_12338,N_8369);
nor U13759 (N_13759,N_7060,N_6417);
and U13760 (N_13760,N_12378,N_8678);
nand U13761 (N_13761,N_8636,N_7764);
or U13762 (N_13762,N_9622,N_7746);
or U13763 (N_13763,N_6772,N_9125);
and U13764 (N_13764,N_11503,N_7969);
nor U13765 (N_13765,N_8969,N_12363);
and U13766 (N_13766,N_6716,N_12310);
nor U13767 (N_13767,N_8809,N_8874);
or U13768 (N_13768,N_11725,N_6293);
nand U13769 (N_13769,N_11432,N_11290);
or U13770 (N_13770,N_11656,N_8655);
nor U13771 (N_13771,N_12425,N_6564);
or U13772 (N_13772,N_6477,N_7586);
or U13773 (N_13773,N_6507,N_7054);
and U13774 (N_13774,N_7134,N_10621);
and U13775 (N_13775,N_9775,N_8003);
and U13776 (N_13776,N_9463,N_9043);
xnor U13777 (N_13777,N_9584,N_9973);
or U13778 (N_13778,N_6466,N_6745);
and U13779 (N_13779,N_9061,N_11675);
xnor U13780 (N_13780,N_12218,N_8411);
nor U13781 (N_13781,N_11450,N_11906);
nand U13782 (N_13782,N_6372,N_8907);
or U13783 (N_13783,N_11448,N_6952);
nor U13784 (N_13784,N_7373,N_10177);
xor U13785 (N_13785,N_8151,N_10513);
or U13786 (N_13786,N_10615,N_10787);
or U13787 (N_13787,N_9837,N_8484);
xnor U13788 (N_13788,N_8026,N_11444);
or U13789 (N_13789,N_11779,N_9132);
nand U13790 (N_13790,N_6989,N_6725);
nor U13791 (N_13791,N_8953,N_10720);
and U13792 (N_13792,N_10376,N_8759);
and U13793 (N_13793,N_10889,N_9483);
and U13794 (N_13794,N_9857,N_11423);
nand U13795 (N_13795,N_12451,N_10747);
and U13796 (N_13796,N_10836,N_11803);
nor U13797 (N_13797,N_9843,N_9384);
nand U13798 (N_13798,N_6465,N_8342);
xor U13799 (N_13799,N_11997,N_12208);
nand U13800 (N_13800,N_7120,N_12075);
nor U13801 (N_13801,N_6961,N_7309);
or U13802 (N_13802,N_9034,N_10774);
nand U13803 (N_13803,N_10346,N_11865);
and U13804 (N_13804,N_8177,N_9025);
nand U13805 (N_13805,N_8560,N_11672);
and U13806 (N_13806,N_12304,N_11190);
nand U13807 (N_13807,N_6742,N_10070);
nand U13808 (N_13808,N_6913,N_9769);
and U13809 (N_13809,N_10914,N_8146);
or U13810 (N_13810,N_6891,N_6768);
nor U13811 (N_13811,N_10576,N_8818);
nand U13812 (N_13812,N_7238,N_10832);
or U13813 (N_13813,N_6462,N_7491);
xor U13814 (N_13814,N_8409,N_12415);
nand U13815 (N_13815,N_6661,N_9037);
and U13816 (N_13816,N_6441,N_9287);
nand U13817 (N_13817,N_10441,N_10705);
and U13818 (N_13818,N_8593,N_11670);
nor U13819 (N_13819,N_10096,N_8251);
and U13820 (N_13820,N_7761,N_9808);
nor U13821 (N_13821,N_6880,N_9110);
xor U13822 (N_13822,N_9794,N_11752);
nand U13823 (N_13823,N_7540,N_8868);
nand U13824 (N_13824,N_9668,N_10687);
nand U13825 (N_13825,N_11546,N_9585);
nor U13826 (N_13826,N_10947,N_10866);
nand U13827 (N_13827,N_8947,N_7698);
xor U13828 (N_13828,N_10140,N_10958);
nor U13829 (N_13829,N_10764,N_7622);
and U13830 (N_13830,N_8611,N_12389);
or U13831 (N_13831,N_7459,N_10447);
nor U13832 (N_13832,N_9068,N_10193);
nor U13833 (N_13833,N_9331,N_11902);
nand U13834 (N_13834,N_11066,N_8684);
and U13835 (N_13835,N_10094,N_7562);
or U13836 (N_13836,N_9766,N_10284);
or U13837 (N_13837,N_9543,N_9214);
nor U13838 (N_13838,N_10066,N_9021);
nor U13839 (N_13839,N_6317,N_7967);
and U13840 (N_13840,N_7971,N_9173);
xnor U13841 (N_13841,N_9393,N_8278);
nor U13842 (N_13842,N_10869,N_11385);
and U13843 (N_13843,N_11594,N_7711);
nor U13844 (N_13844,N_11517,N_11377);
nor U13845 (N_13845,N_9825,N_11243);
nand U13846 (N_13846,N_10897,N_11911);
nor U13847 (N_13847,N_9027,N_10793);
xor U13848 (N_13848,N_12135,N_11165);
and U13849 (N_13849,N_9486,N_9898);
nor U13850 (N_13850,N_8422,N_7526);
nand U13851 (N_13851,N_9280,N_9664);
nand U13852 (N_13852,N_7678,N_8808);
nor U13853 (N_13853,N_11642,N_9160);
and U13854 (N_13854,N_10698,N_11689);
nand U13855 (N_13855,N_10495,N_10703);
and U13856 (N_13856,N_9790,N_10753);
nor U13857 (N_13857,N_8080,N_10517);
or U13858 (N_13858,N_8755,N_7410);
or U13859 (N_13859,N_8693,N_11267);
nor U13860 (N_13860,N_11479,N_7636);
xor U13861 (N_13861,N_7708,N_10776);
and U13862 (N_13862,N_8811,N_9044);
or U13863 (N_13863,N_8004,N_7447);
nor U13864 (N_13864,N_7204,N_11987);
and U13865 (N_13865,N_8039,N_11004);
or U13866 (N_13866,N_12496,N_12147);
nand U13867 (N_13867,N_6361,N_10442);
xor U13868 (N_13868,N_10800,N_10159);
nand U13869 (N_13869,N_11519,N_8473);
nand U13870 (N_13870,N_6313,N_11085);
and U13871 (N_13871,N_11473,N_7977);
or U13872 (N_13872,N_6416,N_8985);
xnor U13873 (N_13873,N_8181,N_7218);
nor U13874 (N_13874,N_10921,N_12282);
nor U13875 (N_13875,N_7462,N_6876);
nor U13876 (N_13876,N_8822,N_11343);
or U13877 (N_13877,N_7701,N_8425);
nor U13878 (N_13878,N_7696,N_9614);
nand U13879 (N_13879,N_7084,N_7223);
or U13880 (N_13880,N_8499,N_10484);
xor U13881 (N_13881,N_8131,N_8483);
nor U13882 (N_13882,N_11696,N_8466);
and U13883 (N_13883,N_10466,N_8737);
nand U13884 (N_13884,N_11874,N_11272);
or U13885 (N_13885,N_8672,N_9785);
or U13886 (N_13886,N_7279,N_9292);
or U13887 (N_13887,N_8706,N_11909);
or U13888 (N_13888,N_6945,N_11802);
or U13889 (N_13889,N_10599,N_8983);
nor U13890 (N_13890,N_9952,N_8170);
and U13891 (N_13891,N_11107,N_11715);
nand U13892 (N_13892,N_9931,N_12235);
nand U13893 (N_13893,N_10214,N_6348);
nand U13894 (N_13894,N_10915,N_6598);
and U13895 (N_13895,N_7262,N_8976);
and U13896 (N_13896,N_12053,N_8633);
and U13897 (N_13897,N_10130,N_11292);
nor U13898 (N_13898,N_12120,N_7841);
nor U13899 (N_13899,N_7291,N_8542);
and U13900 (N_13900,N_7088,N_10475);
nand U13901 (N_13901,N_6770,N_7434);
nor U13902 (N_13902,N_11892,N_10772);
or U13903 (N_13903,N_7130,N_11563);
or U13904 (N_13904,N_6982,N_10213);
nor U13905 (N_13905,N_8399,N_6344);
or U13906 (N_13906,N_9179,N_8894);
and U13907 (N_13907,N_7486,N_9536);
xnor U13908 (N_13908,N_11758,N_7905);
nor U13909 (N_13909,N_12263,N_9526);
nor U13910 (N_13910,N_7857,N_10670);
or U13911 (N_13911,N_9518,N_7193);
or U13912 (N_13912,N_11513,N_12006);
and U13913 (N_13913,N_6814,N_10856);
nand U13914 (N_13914,N_10633,N_12113);
and U13915 (N_13915,N_7051,N_10388);
or U13916 (N_13916,N_10908,N_9681);
nand U13917 (N_13917,N_11683,N_10250);
or U13918 (N_13918,N_6950,N_10973);
nor U13919 (N_13919,N_9217,N_10021);
or U13920 (N_13920,N_11174,N_9225);
nor U13921 (N_13921,N_11293,N_10341);
or U13922 (N_13922,N_9423,N_9574);
or U13923 (N_13923,N_7731,N_10326);
and U13924 (N_13924,N_9516,N_12096);
nand U13925 (N_13925,N_10954,N_6321);
xnor U13926 (N_13926,N_10850,N_9009);
or U13927 (N_13927,N_10340,N_7923);
xnor U13928 (N_13928,N_11732,N_10101);
and U13929 (N_13929,N_10887,N_11801);
xnor U13930 (N_13930,N_10078,N_7221);
nor U13931 (N_13931,N_9623,N_6506);
or U13932 (N_13932,N_8145,N_9564);
and U13933 (N_13933,N_6501,N_7855);
nor U13934 (N_13934,N_7350,N_6521);
xnor U13935 (N_13935,N_6954,N_6790);
and U13936 (N_13936,N_12175,N_10917);
nand U13937 (N_13937,N_8298,N_6999);
and U13938 (N_13938,N_6414,N_11306);
nor U13939 (N_13939,N_6540,N_12029);
xnor U13940 (N_13940,N_8933,N_8324);
and U13941 (N_13941,N_9673,N_7913);
and U13942 (N_13942,N_9180,N_6740);
nand U13943 (N_13943,N_10473,N_6905);
and U13944 (N_13944,N_7826,N_9095);
nor U13945 (N_13945,N_12196,N_6798);
or U13946 (N_13946,N_10136,N_7637);
and U13947 (N_13947,N_8113,N_8476);
xnor U13948 (N_13948,N_11383,N_6732);
or U13949 (N_13949,N_10828,N_8059);
nand U13950 (N_13950,N_12186,N_9317);
or U13951 (N_13951,N_9342,N_9534);
nand U13952 (N_13952,N_12027,N_6272);
nor U13953 (N_13953,N_10310,N_12139);
or U13954 (N_13954,N_12375,N_8377);
nor U13955 (N_13955,N_9528,N_6307);
nor U13956 (N_13956,N_6763,N_6502);
nand U13957 (N_13957,N_11549,N_7804);
nand U13958 (N_13958,N_9465,N_10192);
nor U13959 (N_13959,N_7003,N_8996);
and U13960 (N_13960,N_10478,N_10761);
xnor U13961 (N_13961,N_10810,N_10722);
and U13962 (N_13962,N_6559,N_11074);
nor U13963 (N_13963,N_10351,N_12464);
and U13964 (N_13964,N_10728,N_11162);
or U13965 (N_13965,N_7687,N_10766);
and U13966 (N_13966,N_9684,N_10282);
nor U13967 (N_13967,N_8942,N_12484);
nor U13968 (N_13968,N_7343,N_12341);
nand U13969 (N_13969,N_6996,N_10165);
and U13970 (N_13970,N_6921,N_8047);
xor U13971 (N_13971,N_9819,N_9157);
nand U13972 (N_13972,N_12066,N_8263);
nand U13973 (N_13973,N_10939,N_9168);
nor U13974 (N_13974,N_7164,N_11071);
xnor U13975 (N_13975,N_9229,N_7570);
and U13976 (N_13976,N_9625,N_10536);
or U13977 (N_13977,N_6743,N_9506);
and U13978 (N_13978,N_9439,N_6681);
or U13979 (N_13979,N_7379,N_11998);
or U13980 (N_13980,N_10949,N_8459);
nor U13981 (N_13981,N_6642,N_12047);
and U13982 (N_13982,N_10293,N_8984);
or U13983 (N_13983,N_8351,N_7154);
nor U13984 (N_13984,N_7137,N_9795);
nor U13985 (N_13985,N_11424,N_11893);
and U13986 (N_13986,N_6271,N_12402);
xnor U13987 (N_13987,N_10091,N_6529);
or U13988 (N_13988,N_9154,N_8220);
nor U13989 (N_13989,N_6658,N_7001);
nor U13990 (N_13990,N_7106,N_10535);
xnor U13991 (N_13991,N_8419,N_9485);
xor U13992 (N_13992,N_9429,N_7123);
and U13993 (N_13993,N_8361,N_10038);
nor U13994 (N_13994,N_6563,N_11216);
or U13995 (N_13995,N_11183,N_10060);
nor U13996 (N_13996,N_9806,N_12189);
and U13997 (N_13997,N_6476,N_8717);
or U13998 (N_13998,N_9064,N_10233);
and U13999 (N_13999,N_10097,N_11053);
nand U14000 (N_14000,N_12495,N_8008);
nor U14001 (N_14001,N_6415,N_11535);
nor U14002 (N_14002,N_8748,N_11583);
xor U14003 (N_14003,N_11362,N_9960);
nor U14004 (N_14004,N_10210,N_7151);
nand U14005 (N_14005,N_8259,N_9472);
nand U14006 (N_14006,N_11304,N_11068);
nand U14007 (N_14007,N_6892,N_11129);
or U14008 (N_14008,N_8186,N_12412);
nor U14009 (N_14009,N_12249,N_12490);
xor U14010 (N_14010,N_7333,N_11386);
nand U14011 (N_14011,N_9209,N_7452);
nand U14012 (N_14012,N_7383,N_11413);
nor U14013 (N_14013,N_10895,N_8463);
nand U14014 (N_14014,N_7008,N_11505);
and U14015 (N_14015,N_8860,N_7642);
and U14016 (N_14016,N_9707,N_12204);
xor U14017 (N_14017,N_11680,N_10815);
nor U14018 (N_14018,N_6813,N_10675);
nor U14019 (N_14019,N_6448,N_8303);
xor U14020 (N_14020,N_10179,N_8892);
and U14021 (N_14021,N_8076,N_12473);
nand U14022 (N_14022,N_7315,N_9752);
and U14023 (N_14023,N_8563,N_11793);
nor U14024 (N_14024,N_8070,N_11883);
or U14025 (N_14025,N_11576,N_7032);
xnor U14026 (N_14026,N_11811,N_7572);
and U14027 (N_14027,N_7496,N_9832);
and U14028 (N_14028,N_10044,N_9336);
and U14029 (N_14029,N_9851,N_9720);
xnor U14030 (N_14030,N_11736,N_10268);
and U14031 (N_14031,N_11528,N_10837);
nor U14032 (N_14032,N_11205,N_9355);
nor U14033 (N_14033,N_8670,N_7353);
xor U14034 (N_14034,N_10559,N_6378);
and U14035 (N_14035,N_12302,N_9438);
and U14036 (N_14036,N_10110,N_9565);
or U14037 (N_14037,N_11846,N_6457);
nand U14038 (N_14038,N_7644,N_11960);
or U14039 (N_14039,N_9323,N_8203);
nand U14040 (N_14040,N_8107,N_10561);
nor U14041 (N_14041,N_8781,N_10649);
and U14042 (N_14042,N_8795,N_10508);
nor U14043 (N_14043,N_12331,N_11713);
or U14044 (N_14044,N_6574,N_7908);
nand U14045 (N_14045,N_8628,N_8883);
nor U14046 (N_14046,N_11647,N_10385);
nor U14047 (N_14047,N_8686,N_12046);
nand U14048 (N_14048,N_7544,N_11588);
and U14049 (N_14049,N_9855,N_12431);
or U14050 (N_14050,N_7019,N_9371);
and U14051 (N_14051,N_8888,N_10575);
and U14052 (N_14052,N_8338,N_11256);
or U14053 (N_14053,N_11392,N_11885);
nand U14054 (N_14054,N_12295,N_10790);
nor U14055 (N_14055,N_8103,N_8348);
and U14056 (N_14056,N_9782,N_10551);
nor U14057 (N_14057,N_11747,N_7399);
nand U14058 (N_14058,N_10471,N_9434);
or U14059 (N_14059,N_9273,N_11693);
nor U14060 (N_14060,N_8756,N_7066);
and U14061 (N_14061,N_8720,N_9498);
nand U14062 (N_14062,N_8926,N_8445);
nand U14063 (N_14063,N_7707,N_7364);
nor U14064 (N_14064,N_12019,N_10734);
nand U14065 (N_14065,N_9471,N_6782);
nand U14066 (N_14066,N_10217,N_10053);
and U14067 (N_14067,N_9812,N_7887);
or U14068 (N_14068,N_11127,N_8993);
or U14069 (N_14069,N_11030,N_8558);
nor U14070 (N_14070,N_9178,N_11012);
or U14071 (N_14071,N_7940,N_8639);
xnor U14072 (N_14072,N_9005,N_10606);
or U14073 (N_14073,N_11115,N_8395);
nand U14074 (N_14074,N_8215,N_12181);
nor U14075 (N_14075,N_6827,N_7347);
and U14076 (N_14076,N_7670,N_9696);
and U14077 (N_14077,N_6449,N_10391);
and U14078 (N_14078,N_7142,N_6468);
nand U14079 (N_14079,N_10932,N_11632);
nand U14080 (N_14080,N_8559,N_8924);
or U14081 (N_14081,N_11189,N_12164);
and U14082 (N_14082,N_12405,N_10350);
nor U14083 (N_14083,N_6653,N_12050);
and U14084 (N_14084,N_8096,N_7883);
or U14085 (N_14085,N_10208,N_8634);
and U14086 (N_14086,N_10256,N_11268);
or U14087 (N_14087,N_7470,N_9123);
or U14088 (N_14088,N_12488,N_10045);
nand U14089 (N_14089,N_10726,N_7036);
and U14090 (N_14090,N_7681,N_12179);
or U14091 (N_14091,N_11022,N_7396);
or U14092 (N_14092,N_11200,N_6509);
or U14093 (N_14093,N_12031,N_8900);
nor U14094 (N_14094,N_8028,N_10942);
nand U14095 (N_14095,N_11453,N_6689);
or U14096 (N_14096,N_10106,N_10502);
xor U14097 (N_14097,N_7317,N_9338);
or U14098 (N_14098,N_9285,N_6901);
and U14099 (N_14099,N_8160,N_6291);
and U14100 (N_14100,N_6775,N_9577);
or U14101 (N_14101,N_9369,N_11613);
or U14102 (N_14102,N_12387,N_6565);
or U14103 (N_14103,N_11990,N_8383);
nor U14104 (N_14104,N_11724,N_6558);
nor U14105 (N_14105,N_9294,N_7335);
nand U14106 (N_14106,N_7245,N_7355);
nor U14107 (N_14107,N_11166,N_7709);
nor U14108 (N_14108,N_10387,N_9894);
or U14109 (N_14109,N_11111,N_10824);
or U14110 (N_14110,N_6895,N_6513);
nor U14111 (N_14111,N_10085,N_7559);
or U14112 (N_14112,N_10449,N_8125);
or U14113 (N_14113,N_9697,N_9569);
nor U14114 (N_14114,N_10469,N_6588);
or U14115 (N_14115,N_10118,N_8876);
nor U14116 (N_14116,N_6733,N_11101);
or U14117 (N_14117,N_12463,N_10320);
nor U14118 (N_14118,N_11575,N_11197);
nor U14119 (N_14119,N_6933,N_7150);
and U14120 (N_14120,N_11745,N_10799);
nand U14121 (N_14121,N_6520,N_11206);
nor U14122 (N_14122,N_7489,N_11536);
or U14123 (N_14123,N_6972,N_6340);
and U14124 (N_14124,N_12004,N_7365);
xnor U14125 (N_14125,N_10327,N_7348);
nand U14126 (N_14126,N_7680,N_7155);
nor U14127 (N_14127,N_7830,N_7438);
or U14128 (N_14128,N_7135,N_8867);
and U14129 (N_14129,N_10617,N_11472);
nand U14130 (N_14130,N_10147,N_10004);
or U14131 (N_14131,N_9016,N_10276);
nor U14132 (N_14132,N_10126,N_11361);
nand U14133 (N_14133,N_10913,N_8763);
xor U14134 (N_14134,N_11347,N_6637);
nand U14135 (N_14135,N_9264,N_11699);
xor U14136 (N_14136,N_7649,N_11263);
nor U14137 (N_14137,N_10267,N_6371);
nor U14138 (N_14138,N_12043,N_8899);
nor U14139 (N_14139,N_12270,N_9060);
nor U14140 (N_14140,N_10537,N_9072);
nor U14141 (N_14141,N_7020,N_7502);
or U14142 (N_14142,N_10223,N_10258);
and U14143 (N_14143,N_7823,N_8335);
nand U14144 (N_14144,N_12268,N_6590);
nand U14145 (N_14145,N_9013,N_11346);
nand U14146 (N_14146,N_11641,N_6924);
or U14147 (N_14147,N_9023,N_11486);
nand U14148 (N_14148,N_9826,N_9661);
and U14149 (N_14149,N_7202,N_12059);
xnor U14150 (N_14150,N_10538,N_9140);
or U14151 (N_14151,N_7375,N_11914);
or U14152 (N_14152,N_9052,N_9084);
or U14153 (N_14153,N_7860,N_8956);
xnor U14154 (N_14154,N_10522,N_7989);
nand U14155 (N_14155,N_11213,N_8432);
xnor U14156 (N_14156,N_7523,N_7146);
and U14157 (N_14157,N_10292,N_8075);
or U14158 (N_14158,N_7284,N_7387);
and U14159 (N_14159,N_8962,N_7251);
or U14160 (N_14160,N_8545,N_9892);
and U14161 (N_14161,N_11296,N_9454);
nor U14162 (N_14162,N_11596,N_11844);
nor U14163 (N_14163,N_12097,N_11516);
nor U14164 (N_14164,N_8587,N_10911);
nand U14165 (N_14165,N_8306,N_12374);
or U14166 (N_14166,N_7574,N_6722);
or U14167 (N_14167,N_6871,N_6389);
or U14168 (N_14168,N_8485,N_10330);
or U14169 (N_14169,N_10054,N_8099);
or U14170 (N_14170,N_7504,N_8111);
or U14171 (N_14171,N_6377,N_8321);
or U14172 (N_14172,N_10588,N_7494);
or U14173 (N_14173,N_7004,N_10552);
nor U14174 (N_14174,N_10612,N_9469);
and U14175 (N_14175,N_12118,N_7930);
or U14176 (N_14176,N_7871,N_11326);
and U14177 (N_14177,N_10694,N_10395);
nor U14178 (N_14178,N_7495,N_10751);
and U14179 (N_14179,N_6356,N_6846);
nand U14180 (N_14180,N_10176,N_7370);
nor U14181 (N_14181,N_9096,N_9260);
and U14182 (N_14182,N_9344,N_9714);
xor U14183 (N_14183,N_6638,N_9333);
or U14184 (N_14184,N_7538,N_10008);
or U14185 (N_14185,N_7482,N_10811);
or U14186 (N_14186,N_8027,N_7718);
nor U14187 (N_14187,N_12025,N_9895);
xor U14188 (N_14188,N_12450,N_8785);
nand U14189 (N_14189,N_10022,N_7190);
nand U14190 (N_14190,N_9522,N_7118);
and U14191 (N_14191,N_10408,N_9376);
and U14192 (N_14192,N_9818,N_7444);
or U14193 (N_14193,N_12469,N_9634);
nor U14194 (N_14194,N_7027,N_6797);
xnor U14195 (N_14195,N_11843,N_6935);
and U14196 (N_14196,N_11585,N_11177);
and U14197 (N_14197,N_7710,N_7784);
and U14198 (N_14198,N_12381,N_6835);
nor U14199 (N_14199,N_12347,N_10528);
nand U14200 (N_14200,N_10459,N_8205);
and U14201 (N_14201,N_11061,N_9282);
and U14202 (N_14202,N_10931,N_10721);
or U14203 (N_14203,N_10242,N_11169);
or U14204 (N_14204,N_7615,N_8467);
nand U14205 (N_14205,N_12261,N_9900);
nand U14206 (N_14206,N_7402,N_10500);
nor U14207 (N_14207,N_7747,N_10593);
or U14208 (N_14208,N_10545,N_6629);
and U14209 (N_14209,N_8486,N_9799);
nor U14210 (N_14210,N_11114,N_12403);
nand U14211 (N_14211,N_11763,N_7136);
nand U14212 (N_14212,N_11687,N_7882);
and U14213 (N_14213,N_6575,N_11817);
nand U14214 (N_14214,N_8245,N_9789);
or U14215 (N_14215,N_10695,N_7532);
and U14216 (N_14216,N_8493,N_8776);
nand U14217 (N_14217,N_7970,N_9954);
nand U14218 (N_14218,N_8353,N_9693);
nand U14219 (N_14219,N_8591,N_11582);
or U14220 (N_14220,N_6976,N_11993);
nand U14221 (N_14221,N_10073,N_6557);
nand U14222 (N_14222,N_6706,N_7613);
nand U14223 (N_14223,N_12257,N_10331);
and U14224 (N_14224,N_11765,N_10243);
nand U14225 (N_14225,N_10937,N_11476);
nand U14226 (N_14226,N_11038,N_11939);
and U14227 (N_14227,N_7430,N_10759);
or U14228 (N_14228,N_6906,N_6611);
and U14229 (N_14229,N_6360,N_12254);
nor U14230 (N_14230,N_7796,N_7589);
nor U14231 (N_14231,N_9521,N_6874);
and U14232 (N_14232,N_6820,N_10591);
nor U14233 (N_14233,N_8100,N_9201);
nor U14234 (N_14234,N_7450,N_10584);
xnor U14235 (N_14235,N_9174,N_12089);
or U14236 (N_14236,N_6809,N_12194);
or U14237 (N_14237,N_11072,N_8521);
or U14238 (N_14238,N_9237,N_7467);
nor U14239 (N_14239,N_6823,N_6392);
nand U14240 (N_14240,N_8991,N_10128);
xnor U14241 (N_14241,N_8127,N_10108);
and U14242 (N_14242,N_9004,N_9706);
nor U14243 (N_14243,N_10470,N_10573);
or U14244 (N_14244,N_6886,N_9998);
nor U14245 (N_14245,N_6667,N_8007);
xnor U14246 (N_14246,N_11700,N_8912);
and U14247 (N_14247,N_9007,N_7030);
or U14248 (N_14248,N_7116,N_10965);
nand U14249 (N_14249,N_8365,N_7631);
and U14250 (N_14250,N_7852,N_9114);
or U14251 (N_14251,N_9741,N_9177);
and U14252 (N_14252,N_11678,N_9605);
or U14253 (N_14253,N_9196,N_10520);
and U14254 (N_14254,N_9607,N_10116);
xor U14255 (N_14255,N_10992,N_10371);
nor U14256 (N_14256,N_9582,N_10251);
or U14257 (N_14257,N_12467,N_7647);
and U14258 (N_14258,N_10982,N_10714);
and U14259 (N_14259,N_9145,N_8052);
and U14260 (N_14260,N_11437,N_8624);
xnor U14261 (N_14261,N_10299,N_8414);
and U14262 (N_14262,N_9591,N_8388);
and U14263 (N_14263,N_9761,N_12260);
or U14264 (N_14264,N_10501,N_7777);
xnor U14265 (N_14265,N_8708,N_7509);
nand U14266 (N_14266,N_10366,N_11442);
nand U14267 (N_14267,N_9891,N_8066);
and U14268 (N_14268,N_7010,N_11784);
xnor U14269 (N_14269,N_10993,N_10316);
nand U14270 (N_14270,N_7110,N_6401);
nor U14271 (N_14271,N_9721,N_12101);
nand U14272 (N_14272,N_11262,N_6929);
and U14273 (N_14273,N_9841,N_12429);
nor U14274 (N_14274,N_8884,N_12211);
nor U14275 (N_14275,N_9092,N_11195);
or U14276 (N_14276,N_7481,N_12203);
or U14277 (N_14277,N_7017,N_10393);
nand U14278 (N_14278,N_7029,N_7634);
nand U14279 (N_14279,N_11064,N_10818);
nor U14280 (N_14280,N_7265,N_10896);
nand U14281 (N_14281,N_8986,N_8010);
or U14282 (N_14282,N_9267,N_7660);
nor U14283 (N_14283,N_12109,N_11917);
nor U14284 (N_14284,N_6542,N_11572);
xnor U14285 (N_14285,N_7833,N_11193);
nor U14286 (N_14286,N_6864,N_10912);
nand U14287 (N_14287,N_9667,N_9717);
nor U14288 (N_14288,N_7956,N_7163);
or U14289 (N_14289,N_10198,N_11273);
xnor U14290 (N_14290,N_6426,N_10272);
nor U14291 (N_14291,N_11261,N_8857);
and U14292 (N_14292,N_6390,N_6384);
nor U14293 (N_14293,N_10081,N_11567);
nor U14294 (N_14294,N_6429,N_9152);
nor U14295 (N_14295,N_7023,N_12222);
xnor U14296 (N_14296,N_12070,N_10813);
nand U14297 (N_14297,N_7828,N_8509);
or U14298 (N_14298,N_12361,N_8394);
and U14299 (N_14299,N_11830,N_7832);
nand U14300 (N_14300,N_7171,N_11221);
or U14301 (N_14301,N_6893,N_9067);
xor U14302 (N_14302,N_6903,N_10610);
and U14303 (N_14303,N_11443,N_9414);
or U14304 (N_14304,N_6636,N_11962);
nor U14305 (N_14305,N_9597,N_9735);
nand U14306 (N_14306,N_10129,N_11507);
and U14307 (N_14307,N_8258,N_7714);
nor U14308 (N_14308,N_7067,N_11568);
or U14309 (N_14309,N_8654,N_11351);
and U14310 (N_14310,N_9436,N_11229);
and U14311 (N_14311,N_11667,N_11491);
and U14312 (N_14312,N_7384,N_12393);
nand U14313 (N_14313,N_11873,N_9222);
xor U14314 (N_14314,N_8471,N_10295);
or U14315 (N_14315,N_11131,N_7648);
and U14316 (N_14316,N_9269,N_12376);
xnor U14317 (N_14317,N_8450,N_11723);
or U14318 (N_14318,N_10590,N_8508);
xor U14319 (N_14319,N_10401,N_8416);
or U14320 (N_14320,N_8197,N_10674);
and U14321 (N_14321,N_9402,N_10655);
xnor U14322 (N_14322,N_12372,N_10519);
nor U14323 (N_14323,N_11454,N_9739);
or U14324 (N_14324,N_9228,N_10952);
or U14325 (N_14325,N_12026,N_6688);
or U14326 (N_14326,N_6327,N_11224);
nand U14327 (N_14327,N_8093,N_9563);
nand U14328 (N_14328,N_8326,N_7986);
or U14329 (N_14329,N_11235,N_8550);
nand U14330 (N_14330,N_9473,N_9392);
nor U14331 (N_14331,N_11219,N_8423);
and U14332 (N_14332,N_9343,N_6398);
and U14333 (N_14333,N_10245,N_7816);
or U14334 (N_14334,N_11799,N_6326);
and U14335 (N_14335,N_10719,N_9993);
and U14336 (N_14336,N_11749,N_12406);
and U14337 (N_14337,N_12438,N_11762);
nand U14338 (N_14338,N_11379,N_8967);
nand U14339 (N_14339,N_11707,N_11406);
nor U14340 (N_14340,N_7323,N_11086);
or U14341 (N_14341,N_10304,N_10334);
or U14342 (N_14342,N_8408,N_7693);
nor U14343 (N_14343,N_10452,N_7943);
or U14344 (N_14344,N_11532,N_6620);
and U14345 (N_14345,N_10583,N_6644);
or U14346 (N_14346,N_8718,N_12038);
or U14347 (N_14347,N_10504,N_11923);
or U14348 (N_14348,N_10834,N_9768);
nor U14349 (N_14349,N_7096,N_11780);
and U14350 (N_14350,N_7881,N_7356);
or U14351 (N_14351,N_7643,N_9183);
nor U14352 (N_14352,N_6566,N_11584);
and U14353 (N_14353,N_6320,N_8364);
nor U14354 (N_14354,N_6387,N_8929);
or U14355 (N_14355,N_6512,N_10023);
and U14356 (N_14356,N_12226,N_10172);
nor U14357 (N_14357,N_12386,N_7898);
nor U14358 (N_14358,N_9677,N_8505);
or U14359 (N_14359,N_11806,N_6516);
or U14360 (N_14360,N_7590,N_9443);
or U14361 (N_14361,N_9918,N_11211);
nor U14362 (N_14362,N_11153,N_9935);
nor U14363 (N_14363,N_10567,N_12127);
nor U14364 (N_14364,N_10248,N_11228);
and U14365 (N_14365,N_8974,N_11126);
or U14366 (N_14366,N_11058,N_9871);
and U14367 (N_14367,N_11708,N_6947);
nand U14368 (N_14368,N_10337,N_8184);
nand U14369 (N_14369,N_10901,N_6535);
or U14370 (N_14370,N_9722,N_8681);
and U14371 (N_14371,N_11087,N_8101);
and U14372 (N_14372,N_8017,N_11829);
or U14373 (N_14373,N_8527,N_11427);
nand U14374 (N_14374,N_7411,N_11957);
nor U14375 (N_14375,N_9026,N_7514);
nand U14376 (N_14376,N_9497,N_6363);
xor U14377 (N_14377,N_11920,N_7727);
nand U14378 (N_14378,N_6631,N_10829);
nand U14379 (N_14379,N_9291,N_8540);
nand U14380 (N_14380,N_7937,N_11645);
nor U14381 (N_14381,N_11117,N_7575);
and U14382 (N_14382,N_10525,N_7466);
nand U14383 (N_14383,N_9902,N_6858);
nor U14384 (N_14384,N_11426,N_12022);
nand U14385 (N_14385,N_9347,N_11002);
nor U14386 (N_14386,N_11164,N_12188);
and U14387 (N_14387,N_9863,N_8921);
nand U14388 (N_14388,N_8256,N_11234);
or U14389 (N_14389,N_8112,N_9326);
nor U14390 (N_14390,N_7112,N_8782);
and U14391 (N_14391,N_10451,N_8147);
nor U14392 (N_14392,N_6993,N_11551);
nor U14393 (N_14393,N_9621,N_8625);
and U14394 (N_14394,N_7424,N_11447);
nor U14395 (N_14395,N_12085,N_12428);
xnor U14396 (N_14396,N_7694,N_12358);
xnor U14397 (N_14397,N_9144,N_8332);
nor U14398 (N_14398,N_11028,N_11592);
nor U14399 (N_14399,N_9238,N_8555);
or U14400 (N_14400,N_7818,N_10373);
xnor U14401 (N_14401,N_8060,N_11705);
and U14402 (N_14402,N_10397,N_11852);
xnor U14403 (N_14403,N_6765,N_9298);
nor U14404 (N_14404,N_6995,N_7755);
xnor U14405 (N_14405,N_7278,N_7187);
and U14406 (N_14406,N_8382,N_8087);
nand U14407 (N_14407,N_8733,N_12176);
nand U14408 (N_14408,N_10589,N_8095);
nor U14409 (N_14409,N_11867,N_7181);
or U14410 (N_14410,N_6801,N_10409);
nor U14411 (N_14411,N_6624,N_8511);
nand U14412 (N_14412,N_9608,N_11372);
nand U14413 (N_14413,N_11170,N_11266);
and U14414 (N_14414,N_10596,N_7263);
or U14415 (N_14415,N_10279,N_11929);
nand U14416 (N_14416,N_9610,N_11041);
or U14417 (N_14417,N_11332,N_10454);
nor U14418 (N_14418,N_7811,N_10457);
xnor U14419 (N_14419,N_6560,N_10640);
and U14420 (N_14420,N_11538,N_6958);
nor U14421 (N_14421,N_9748,N_11005);
or U14422 (N_14422,N_6968,N_8547);
nand U14423 (N_14423,N_7684,N_7188);
nor U14424 (N_14424,N_11025,N_10369);
nand U14425 (N_14425,N_7780,N_8270);
nand U14426 (N_14426,N_11881,N_10870);
or U14427 (N_14427,N_8739,N_7013);
and U14428 (N_14428,N_10414,N_9546);
nand U14429 (N_14429,N_11716,N_8434);
nor U14430 (N_14430,N_9579,N_10358);
nor U14431 (N_14431,N_7473,N_9520);
nand U14432 (N_14432,N_7180,N_8363);
nor U14433 (N_14433,N_12008,N_11288);
nor U14434 (N_14434,N_9725,N_11121);
nor U14435 (N_14435,N_10676,N_10511);
and U14436 (N_14436,N_10970,N_12296);
nand U14437 (N_14437,N_10699,N_7939);
or U14438 (N_14438,N_7242,N_10613);
or U14439 (N_14439,N_8234,N_10113);
or U14440 (N_14440,N_12433,N_7276);
nor U14441 (N_14441,N_6287,N_10425);
nor U14442 (N_14442,N_12435,N_7851);
nor U14443 (N_14443,N_11308,N_9767);
or U14444 (N_14444,N_12420,N_7247);
or U14445 (N_14445,N_11052,N_11951);
and U14446 (N_14446,N_8704,N_10273);
and U14447 (N_14447,N_12449,N_10404);
nor U14448 (N_14448,N_6625,N_10547);
nor U14449 (N_14449,N_7479,N_6337);
and U14450 (N_14450,N_6896,N_9295);
or U14451 (N_14451,N_11017,N_6349);
and U14452 (N_14452,N_6405,N_6963);
xnor U14453 (N_14453,N_11182,N_9896);
nor U14454 (N_14454,N_11367,N_11008);
xnor U14455 (N_14455,N_7346,N_9408);
nand U14456 (N_14456,N_6985,N_11809);
xor U14457 (N_14457,N_11145,N_6650);
or U14458 (N_14458,N_7560,N_8729);
or U14459 (N_14459,N_10209,N_6634);
or U14460 (N_14460,N_7890,N_11698);
nor U14461 (N_14461,N_7248,N_12045);
or U14462 (N_14462,N_7114,N_9619);
nor U14463 (N_14463,N_12243,N_12419);
xnor U14464 (N_14464,N_9215,N_7543);
xnor U14465 (N_14465,N_9893,N_7200);
nand U14466 (N_14466,N_11230,N_8891);
nand U14467 (N_14467,N_7277,N_8046);
or U14468 (N_14468,N_11673,N_10194);
nor U14469 (N_14469,N_8123,N_7990);
and U14470 (N_14470,N_6922,N_10777);
nor U14471 (N_14471,N_9908,N_11590);
nand U14472 (N_14472,N_8762,N_9425);
nor U14473 (N_14473,N_8949,N_7094);
nand U14474 (N_14474,N_11831,N_8784);
nand U14475 (N_14475,N_6990,N_7282);
or U14476 (N_14476,N_9322,N_6266);
and U14477 (N_14477,N_12385,N_8794);
and U14478 (N_14478,N_8869,N_7968);
or U14479 (N_14479,N_7377,N_11181);
nand U14480 (N_14480,N_7064,N_10156);
or U14481 (N_14481,N_9749,N_11191);
and U14482 (N_14482,N_6959,N_7519);
nor U14483 (N_14483,N_10356,N_11327);
and U14484 (N_14484,N_9971,N_7713);
xor U14485 (N_14485,N_8538,N_9437);
or U14486 (N_14486,N_7156,N_12169);
and U14487 (N_14487,N_10587,N_8945);
nand U14488 (N_14488,N_7769,N_11257);
nor U14489 (N_14489,N_12474,N_7916);
xnor U14490 (N_14490,N_6268,N_7176);
nand U14491 (N_14491,N_9391,N_10631);
nor U14492 (N_14492,N_7601,N_12303);
nor U14493 (N_14493,N_9604,N_8138);
nor U14494 (N_14494,N_7232,N_7147);
nor U14495 (N_14495,N_6828,N_8064);
xor U14496 (N_14496,N_6931,N_8285);
or U14497 (N_14497,N_7596,N_12055);
and U14498 (N_14498,N_11148,N_6969);
nand U14499 (N_14499,N_11029,N_7314);
nor U14500 (N_14500,N_11297,N_9199);
or U14501 (N_14501,N_7803,N_6608);
nand U14502 (N_14502,N_9680,N_9650);
or U14503 (N_14503,N_8819,N_9758);
or U14504 (N_14504,N_9846,N_8429);
xor U14505 (N_14505,N_9947,N_10232);
xnor U14506 (N_14506,N_9906,N_7895);
or U14507 (N_14507,N_7717,N_10347);
nand U14508 (N_14508,N_7652,N_8609);
nor U14509 (N_14509,N_6260,N_7269);
nand U14510 (N_14510,N_8619,N_10448);
or U14511 (N_14511,N_11496,N_12205);
xnor U14512 (N_14512,N_8136,N_9460);
nor U14513 (N_14513,N_10375,N_11322);
and U14514 (N_14514,N_10894,N_10462);
nor U14515 (N_14515,N_11088,N_10711);
xnor U14516 (N_14516,N_10491,N_8833);
nand U14517 (N_14517,N_6718,N_6948);
nand U14518 (N_14518,N_12318,N_7719);
nand U14519 (N_14519,N_7255,N_8973);
nand U14520 (N_14520,N_12010,N_10667);
and U14521 (N_14521,N_7478,N_6421);
nor U14522 (N_14522,N_8293,N_6259);
or U14523 (N_14523,N_11270,N_11898);
nor U14524 (N_14524,N_12079,N_6297);
or U14525 (N_14525,N_6568,N_9231);
nor U14526 (N_14526,N_8557,N_12131);
or U14527 (N_14527,N_7616,N_8354);
xnor U14528 (N_14528,N_9024,N_11096);
or U14529 (N_14529,N_6641,N_9679);
nand U14530 (N_14530,N_9655,N_11773);
or U14531 (N_14531,N_10164,N_7813);
or U14532 (N_14532,N_11617,N_6579);
nor U14533 (N_14533,N_9557,N_9545);
nor U14534 (N_14534,N_8691,N_11751);
or U14535 (N_14535,N_8928,N_8371);
nor U14536 (N_14536,N_6860,N_6843);
xnor U14537 (N_14537,N_9046,N_10626);
and U14538 (N_14538,N_6949,N_9296);
or U14539 (N_14539,N_7625,N_6925);
nand U14540 (N_14540,N_7148,N_12041);
xnor U14541 (N_14541,N_10956,N_11338);
and U14542 (N_14542,N_8415,N_12494);
nor U14543 (N_14543,N_7775,N_8179);
xor U14544 (N_14544,N_8714,N_12472);
xor U14545 (N_14545,N_10111,N_10643);
or U14546 (N_14546,N_10773,N_9554);
or U14547 (N_14547,N_8917,N_8638);
nor U14548 (N_14548,N_12171,N_11077);
nand U14549 (N_14549,N_7312,N_8519);
xor U14550 (N_14550,N_11344,N_6412);
xor U14551 (N_14551,N_9151,N_7600);
or U14552 (N_14552,N_7397,N_9792);
nand U14553 (N_14553,N_10180,N_9911);
nor U14554 (N_14554,N_8749,N_9560);
or U14555 (N_14555,N_7880,N_7952);
and U14556 (N_14556,N_10988,N_7107);
and U14557 (N_14557,N_10906,N_9927);
or U14558 (N_14558,N_11488,N_6904);
nand U14559 (N_14559,N_9378,N_12465);
and U14560 (N_14560,N_7063,N_12129);
nor U14561 (N_14561,N_11054,N_10755);
nor U14562 (N_14562,N_10899,N_8431);
nor U14563 (N_14563,N_7558,N_12430);
and U14564 (N_14564,N_9791,N_10361);
nor U14565 (N_14565,N_10742,N_9186);
nor U14566 (N_14566,N_11023,N_6737);
or U14567 (N_14567,N_8495,N_11661);
nor U14568 (N_14568,N_11382,N_12201);
or U14569 (N_14569,N_10184,N_11395);
or U14570 (N_14570,N_8620,N_12446);
nor U14571 (N_14571,N_10224,N_9645);
or U14572 (N_14572,N_8919,N_9866);
and U14573 (N_14573,N_8850,N_11930);
nor U14574 (N_14574,N_6632,N_8368);
and U14575 (N_14575,N_11858,N_9194);
nor U14576 (N_14576,N_7005,N_12408);
nor U14577 (N_14577,N_11336,N_7734);
nand U14578 (N_14578,N_7194,N_8778);
or U14579 (N_14579,N_9705,N_7779);
and U14580 (N_14580,N_12339,N_10412);
nand U14581 (N_14581,N_7475,N_9760);
nor U14582 (N_14582,N_9255,N_7679);
nand U14583 (N_14583,N_6738,N_10291);
and U14584 (N_14584,N_7553,N_8770);
or U14585 (N_14585,N_9861,N_6649);
nand U14586 (N_14586,N_10439,N_11839);
or U14587 (N_14587,N_11417,N_9445);
or U14588 (N_14588,N_8398,N_9814);
or U14589 (N_14589,N_10498,N_10529);
nor U14590 (N_14590,N_12001,N_6705);
nand U14591 (N_14591,N_8977,N_9117);
xnor U14592 (N_14592,N_6587,N_10661);
nor U14593 (N_14593,N_10481,N_7847);
and U14594 (N_14594,N_6623,N_11643);
nor U14595 (N_14595,N_12121,N_11738);
and U14596 (N_14596,N_8277,N_12195);
and U14597 (N_14597,N_11070,N_9467);
nor U14598 (N_14598,N_11577,N_8780);
nor U14599 (N_14599,N_7919,N_12161);
and U14600 (N_14600,N_8036,N_12035);
xor U14601 (N_14601,N_9777,N_6704);
and U14602 (N_14602,N_10871,N_8903);
nor U14603 (N_14603,N_10145,N_11217);
nand U14604 (N_14604,N_11452,N_11777);
and U14605 (N_14605,N_9762,N_9626);
nor U14606 (N_14606,N_12395,N_10679);
and U14607 (N_14607,N_10862,N_7933);
or U14608 (N_14608,N_8703,N_11018);
xor U14609 (N_14609,N_12090,N_10249);
xnor U14610 (N_14610,N_10512,N_8267);
nor U14611 (N_14611,N_11412,N_9246);
or U14612 (N_14612,N_6288,N_7691);
nor U14613 (N_14613,N_12298,N_6942);
nand U14614 (N_14614,N_9970,N_7261);
nor U14615 (N_14615,N_7518,N_7099);
nor U14616 (N_14616,N_12477,N_9686);
and U14617 (N_14617,N_10010,N_10805);
nor U14618 (N_14618,N_11944,N_6318);
xnor U14619 (N_14619,N_10983,N_11495);
or U14620 (N_14620,N_7736,N_8129);
and U14621 (N_14621,N_6592,N_8548);
nor U14622 (N_14622,N_8954,N_9899);
and U14623 (N_14623,N_10178,N_7361);
nand U14624 (N_14624,N_11927,N_11946);
or U14625 (N_14625,N_7607,N_6406);
nand U14626 (N_14626,N_7820,N_7892);
xnor U14627 (N_14627,N_11060,N_7963);
nand U14628 (N_14628,N_11365,N_8401);
and U14629 (N_14629,N_9038,N_9479);
and U14630 (N_14630,N_11791,N_10090);
and U14631 (N_14631,N_10075,N_12221);
and U14632 (N_14632,N_8847,N_9388);
nor U14633 (N_14633,N_8988,N_8433);
or U14634 (N_14634,N_9275,N_6844);
or U14635 (N_14635,N_11471,N_12077);
nor U14636 (N_14636,N_10725,N_6400);
nand U14637 (N_14637,N_6257,N_8659);
nor U14638 (N_14638,N_10812,N_9995);
nor U14639 (N_14639,N_7806,N_6478);
nor U14640 (N_14640,N_7510,N_7529);
nor U14641 (N_14641,N_8406,N_11832);
nor U14642 (N_14642,N_7662,N_9959);
and U14643 (N_14643,N_6837,N_11635);
xor U14644 (N_14644,N_12163,N_7109);
nor U14645 (N_14645,N_12233,N_6630);
or U14646 (N_14646,N_7145,N_11090);
and U14647 (N_14647,N_7904,N_7420);
and U14648 (N_14648,N_10154,N_6329);
nand U14649 (N_14649,N_8217,N_10266);
nor U14650 (N_14650,N_8840,N_11212);
xor U14651 (N_14651,N_8157,N_8142);
nand U14652 (N_14652,N_7072,N_10082);
nor U14653 (N_14653,N_9493,N_6712);
and U14654 (N_14654,N_7787,N_9703);
and U14655 (N_14655,N_8711,N_12404);
or U14656 (N_14656,N_11940,N_9166);
nor U14657 (N_14657,N_8083,N_11242);
or U14658 (N_14658,N_9548,N_10664);
or U14659 (N_14659,N_10975,N_8297);
and U14660 (N_14660,N_7571,N_7173);
and U14661 (N_14661,N_7104,N_10492);
nand U14662 (N_14662,N_10084,N_7797);
nand U14663 (N_14663,N_8058,N_6894);
nor U14664 (N_14664,N_12285,N_11475);
xnor U14665 (N_14665,N_9811,N_6446);
and U14666 (N_14666,N_7581,N_7550);
nand U14667 (N_14667,N_12251,N_7798);
and U14668 (N_14668,N_11415,N_9640);
or U14669 (N_14669,N_9035,N_11730);
and U14670 (N_14670,N_10996,N_12343);
nor U14671 (N_14671,N_9859,N_11264);
and U14672 (N_14672,N_8500,N_8182);
nand U14673 (N_14673,N_10807,N_10531);
and U14674 (N_14674,N_8554,N_10229);
nor U14675 (N_14675,N_10183,N_7213);
nor U14676 (N_14676,N_11571,N_9594);
nand U14677 (N_14677,N_10037,N_7393);
nand U14678 (N_14678,N_7742,N_8760);
or U14679 (N_14679,N_10318,N_11163);
and U14680 (N_14680,N_7925,N_10142);
nand U14681 (N_14681,N_6867,N_8304);
and U14682 (N_14682,N_8385,N_12448);
and U14683 (N_14683,N_7320,N_11760);
nand U14684 (N_14684,N_12456,N_8630);
and U14685 (N_14685,N_11826,N_9262);
and U14686 (N_14686,N_10690,N_8389);
nand U14687 (N_14687,N_8658,N_11033);
and U14688 (N_14688,N_6877,N_7448);
nor U14689 (N_14689,N_11980,N_8766);
or U14690 (N_14690,N_7706,N_6250);
xor U14691 (N_14691,N_11922,N_10852);
nor U14692 (N_14692,N_9921,N_9914);
and U14693 (N_14693,N_7730,N_11521);
and U14694 (N_14694,N_10076,N_11876);
or U14695 (N_14695,N_12063,N_9020);
and U14696 (N_14696,N_10411,N_11320);
xor U14697 (N_14697,N_6691,N_9457);
nor U14698 (N_14698,N_9578,N_6596);
and U14699 (N_14699,N_11972,N_7380);
nand U14700 (N_14700,N_9205,N_7359);
and U14701 (N_14701,N_11138,N_11067);
nand U14702 (N_14702,N_11276,N_6407);
nor U14703 (N_14703,N_7304,N_12271);
or U14704 (N_14704,N_12432,N_11287);
and U14705 (N_14705,N_12365,N_7958);
nand U14706 (N_14706,N_7525,N_9683);
or U14707 (N_14707,N_10221,N_6578);
nand U14708 (N_14708,N_11410,N_11112);
nand U14709 (N_14709,N_10325,N_12351);
or U14710 (N_14710,N_8183,N_11210);
or U14711 (N_14711,N_6497,N_9793);
nor U14712 (N_14712,N_6312,N_10333);
and U14713 (N_14713,N_9107,N_12394);
nor U14714 (N_14714,N_8552,N_11285);
nor U14715 (N_14715,N_11063,N_9077);
nor U14716 (N_14716,N_11150,N_8665);
xor U14717 (N_14717,N_6627,N_10009);
nand U14718 (N_14718,N_11036,N_12320);
or U14719 (N_14719,N_12439,N_6304);
and U14720 (N_14720,N_9694,N_12000);
nor U14721 (N_14721,N_9820,N_6428);
xor U14722 (N_14722,N_9031,N_11049);
nand U14723 (N_14723,N_9771,N_11907);
nand U14724 (N_14724,N_10910,N_10307);
and U14725 (N_14725,N_7751,N_9728);
and U14726 (N_14726,N_10904,N_10370);
or U14727 (N_14727,N_7783,N_9747);
and U14728 (N_14728,N_9098,N_7836);
and U14729 (N_14729,N_6902,N_9164);
nor U14730 (N_14730,N_6282,N_10977);
nand U14731 (N_14731,N_7429,N_6278);
nor U14732 (N_14732,N_9150,N_9324);
and U14733 (N_14733,N_7819,N_10222);
and U14734 (N_14734,N_10426,N_9491);
nor U14735 (N_14735,N_9335,N_7226);
nor U14736 (N_14736,N_8014,N_11854);
and U14737 (N_14737,N_8190,N_8710);
or U14738 (N_14738,N_9175,N_10572);
nand U14739 (N_14739,N_8020,N_11553);
and U14740 (N_14740,N_8031,N_8730);
xnor U14741 (N_14741,N_9676,N_6496);
or U14742 (N_14742,N_7522,N_7165);
nor U14743 (N_14743,N_10750,N_6277);
nand U14744 (N_14744,N_10018,N_9535);
or U14745 (N_14745,N_6409,N_11073);
or U14746 (N_14746,N_10359,N_10286);
or U14747 (N_14747,N_7593,N_6670);
nor U14748 (N_14748,N_7240,N_9636);
nand U14749 (N_14749,N_8939,N_9700);
or U14750 (N_14750,N_8208,N_12060);
or U14751 (N_14751,N_10289,N_10945);
or U14752 (N_14752,N_6510,N_9977);
xnor U14753 (N_14753,N_6610,N_10682);
and U14754 (N_14754,N_10700,N_6582);
nor U14755 (N_14755,N_12212,N_11522);
and U14756 (N_14756,N_11880,N_6749);
nor U14757 (N_14757,N_8150,N_10040);
or U14758 (N_14758,N_8743,N_7922);
nand U14759 (N_14759,N_8791,N_6359);
nand U14760 (N_14760,N_8249,N_7640);
and U14761 (N_14761,N_10338,N_8130);
or U14762 (N_14762,N_7049,N_7345);
nand U14763 (N_14763,N_11623,N_7413);
nor U14764 (N_14764,N_11878,N_12240);
nor U14765 (N_14765,N_12335,N_8640);
nor U14766 (N_14766,N_11487,N_11782);
nor U14767 (N_14767,N_11690,N_9734);
or U14768 (N_14768,N_11141,N_9920);
xnor U14769 (N_14769,N_8754,N_7012);
nand U14770 (N_14770,N_9514,N_12236);
and U14771 (N_14771,N_12146,N_10991);
and U14772 (N_14772,N_6621,N_11034);
or U14773 (N_14773,N_10052,N_6633);
xnor U14774 (N_14774,N_11890,N_8334);
nand U14775 (N_14775,N_7214,N_11710);
nor U14776 (N_14776,N_10924,N_7070);
nor U14777 (N_14777,N_6432,N_6685);
nand U14778 (N_14778,N_10792,N_10064);
nor U14779 (N_14779,N_11783,N_9121);
or U14780 (N_14780,N_9251,N_7376);
or U14781 (N_14781,N_7723,N_12234);
or U14782 (N_14782,N_7321,N_12225);
and U14783 (N_14783,N_7222,N_9659);
nor U14784 (N_14784,N_10989,N_8206);
or U14785 (N_14785,N_9257,N_9390);
nand U14786 (N_14786,N_9418,N_10061);
and U14787 (N_14787,N_9539,N_10831);
nand U14788 (N_14788,N_12116,N_9999);
nand U14789 (N_14789,N_10313,N_6656);
xor U14790 (N_14790,N_8308,N_6998);
and U14791 (N_14791,N_11024,N_7290);
or U14792 (N_14792,N_6385,N_10929);
nor U14793 (N_14793,N_11312,N_9048);
nand U14794 (N_14794,N_11457,N_8882);
nor U14795 (N_14795,N_6808,N_10632);
nor U14796 (N_14796,N_11381,N_8053);
or U14797 (N_14797,N_9193,N_8322);
or U14798 (N_14798,N_8139,N_11916);
nand U14799 (N_14799,N_11721,N_11142);
or U14800 (N_14800,N_7885,N_9030);
and U14801 (N_14801,N_7541,N_11250);
or U14802 (N_14802,N_11468,N_6736);
and U14803 (N_14803,N_6369,N_7225);
nand U14804 (N_14804,N_12468,N_6335);
nand U14805 (N_14805,N_7604,N_7419);
or U14806 (N_14806,N_7891,N_9299);
nand U14807 (N_14807,N_9289,N_10999);
or U14808 (N_14808,N_9210,N_8623);
and U14809 (N_14809,N_12421,N_9712);
nor U14810 (N_14810,N_8421,N_7954);
nand U14811 (N_14811,N_7097,N_6639);
and U14812 (N_14812,N_7228,N_10265);
and U14813 (N_14813,N_11440,N_6757);
nand U14814 (N_14814,N_7516,N_12346);
nand U14815 (N_14815,N_9216,N_6549);
and U14816 (N_14816,N_12061,N_9489);
and U14817 (N_14817,N_10938,N_8396);
or U14818 (N_14818,N_7848,N_9788);
or U14819 (N_14819,N_6279,N_12269);
and U14820 (N_14820,N_10598,N_9644);
or U14821 (N_14821,N_7057,N_11298);
or U14822 (N_14822,N_11868,N_10383);
or U14823 (N_14823,N_10051,N_12443);
nor U14824 (N_14824,N_8873,N_10036);
xor U14825 (N_14825,N_7996,N_9265);
or U14826 (N_14826,N_8393,N_11108);
and U14827 (N_14827,N_8305,N_8154);
nor U14828 (N_14828,N_9671,N_10608);
nand U14829 (N_14829,N_7753,N_11649);
or U14830 (N_14830,N_6479,N_7367);
or U14831 (N_14831,N_12294,N_8225);
or U14832 (N_14832,N_9512,N_9149);
and U14833 (N_14833,N_9208,N_7884);
nand U14834 (N_14834,N_9737,N_8958);
or U14835 (N_14835,N_9907,N_10771);
or U14836 (N_14836,N_8823,N_8262);
or U14837 (N_14837,N_10765,N_11400);
nor U14838 (N_14838,N_11232,N_7909);
nor U14839 (N_14839,N_9032,N_6286);
and U14840 (N_14840,N_9558,N_9817);
nand U14841 (N_14841,N_8011,N_8069);
nor U14842 (N_14842,N_9088,N_10203);
nor U14843 (N_14843,N_8732,N_12309);
nand U14844 (N_14844,N_11514,N_6472);
or U14845 (N_14845,N_8583,N_7403);
nor U14846 (N_14846,N_8468,N_7298);
nand U14847 (N_14847,N_9939,N_11421);
or U14848 (N_14848,N_9136,N_8040);
nor U14849 (N_14849,N_9185,N_9475);
and U14850 (N_14850,N_9852,N_9736);
and U14851 (N_14851,N_9968,N_11681);
nand U14852 (N_14852,N_11761,N_8610);
and U14853 (N_14853,N_7606,N_8226);
nor U14854 (N_14854,N_11140,N_10025);
and U14855 (N_14855,N_10884,N_8632);
nand U14856 (N_14856,N_7703,N_10864);
nor U14857 (N_14857,N_11281,N_9529);
or U14858 (N_14858,N_10014,N_9346);
xnor U14859 (N_14859,N_6314,N_7539);
or U14860 (N_14860,N_8565,N_11605);
nor U14861 (N_14861,N_10271,N_9435);
nand U14862 (N_14862,N_10168,N_9913);
nor U14863 (N_14863,N_11031,N_7153);
nand U14864 (N_14864,N_8564,N_11247);
nand U14865 (N_14865,N_8274,N_8055);
and U14866 (N_14866,N_10746,N_8513);
and U14867 (N_14867,N_6518,N_6821);
and U14868 (N_14868,N_10641,N_9377);
and U14869 (N_14869,N_10998,N_9937);
or U14870 (N_14870,N_10527,N_11609);
nor U14871 (N_14871,N_7271,N_6815);
nor U14872 (N_14872,N_7170,N_10709);
and U14873 (N_14873,N_10972,N_12217);
nor U14874 (N_14874,N_7501,N_11790);
and U14875 (N_14875,N_10002,N_7528);
or U14876 (N_14876,N_8441,N_9932);
nand U14877 (N_14877,N_11970,N_9691);
nand U14878 (N_14878,N_12173,N_8280);
or U14879 (N_14879,N_10445,N_10994);
or U14880 (N_14880,N_7451,N_7947);
nor U14881 (N_14881,N_11512,N_6543);
nor U14882 (N_14882,N_11639,N_12422);
or U14883 (N_14883,N_9189,N_12489);
xor U14884 (N_14884,N_8384,N_6602);
nand U14885 (N_14885,N_11043,N_11619);
or U14886 (N_14886,N_12228,N_11504);
and U14887 (N_14887,N_11380,N_11977);
and U14888 (N_14888,N_10012,N_12011);
nor U14889 (N_14889,N_8158,N_10056);
xnor U14890 (N_14890,N_10019,N_6986);
or U14891 (N_14891,N_8663,N_7058);
and U14892 (N_14892,N_9850,N_7025);
xnor U14893 (N_14893,N_7102,N_7762);
xnor U14894 (N_14894,N_8491,N_9003);
nor U14895 (N_14895,N_9134,N_7863);
and U14896 (N_14896,N_8726,N_7132);
and U14897 (N_14897,N_8936,N_8601);
nand U14898 (N_14898,N_9066,N_6934);
nand U14899 (N_14899,N_11733,N_9524);
nor U14900 (N_14900,N_8855,N_8797);
xnor U14901 (N_14901,N_11099,N_6647);
or U14902 (N_14902,N_11805,N_11497);
and U14903 (N_14903,N_10961,N_6825);
xnor U14904 (N_14904,N_6671,N_9685);
and U14905 (N_14905,N_8880,N_9364);
nand U14906 (N_14906,N_12455,N_8469);
and U14907 (N_14907,N_8165,N_6308);
and U14908 (N_14908,N_8244,N_10940);
xor U14909 (N_14909,N_7829,N_10616);
xnor U14910 (N_14910,N_7201,N_7050);
or U14911 (N_14911,N_9315,N_10997);
xor U14912 (N_14912,N_8952,N_8319);
xor U14913 (N_14913,N_7894,N_8790);
xor U14914 (N_14914,N_6663,N_7065);
xor U14915 (N_14915,N_8979,N_8097);
and U14916 (N_14916,N_6926,N_11295);
or U14917 (N_14917,N_10483,N_6411);
and U14918 (N_14918,N_8923,N_7287);
nand U14919 (N_14919,N_11684,N_8386);
and U14920 (N_14920,N_11178,N_11895);
and U14921 (N_14921,N_9699,N_8581);
nand U14922 (N_14922,N_10322,N_10497);
nand U14923 (N_14923,N_7433,N_7260);
nor U14924 (N_14924,N_7069,N_11309);
nand U14925 (N_14925,N_7250,N_6524);
xor U14926 (N_14926,N_9877,N_10294);
or U14927 (N_14927,N_9656,N_10903);
nand U14928 (N_14928,N_10542,N_9226);
nand U14929 (N_14929,N_10429,N_9847);
xnor U14930 (N_14930,N_10577,N_8584);
or U14931 (N_14931,N_10923,N_9306);
nor U14932 (N_14932,N_7646,N_10146);
and U14933 (N_14933,N_12452,N_9056);
and U14934 (N_14934,N_7206,N_6315);
nand U14935 (N_14935,N_7351,N_10506);
and U14936 (N_14936,N_11051,N_8764);
and U14937 (N_14937,N_10259,N_10580);
nor U14938 (N_14938,N_10817,N_11808);
nor U14939 (N_14939,N_9115,N_11566);
nand U14940 (N_14940,N_12190,N_10743);
or U14941 (N_14941,N_10274,N_12005);
nand U14942 (N_14942,N_9765,N_6932);
nor U14943 (N_14943,N_11842,N_11552);
nand U14944 (N_14944,N_8622,N_11378);
nor U14945 (N_14945,N_11389,N_9334);
nand U14946 (N_14946,N_8528,N_10493);
or U14947 (N_14947,N_10095,N_8390);
nand U14948 (N_14948,N_8175,N_9822);
nand U14949 (N_14949,N_6345,N_6907);
nor U14950 (N_14950,N_7195,N_7716);
nor U14951 (N_14951,N_8537,N_7052);
nand U14952 (N_14952,N_11523,N_8417);
or U14953 (N_14953,N_7126,N_8006);
xor U14954 (N_14954,N_7493,N_6980);
or U14955 (N_14955,N_12239,N_9729);
nand U14956 (N_14956,N_9956,N_6296);
nor U14957 (N_14957,N_7671,N_7790);
and U14958 (N_14958,N_12317,N_10190);
and U14959 (N_14959,N_8852,N_7772);
or U14960 (N_14960,N_7474,N_9074);
or U14961 (N_14961,N_10104,N_11526);
or U14962 (N_14962,N_9552,N_8018);
nor U14963 (N_14963,N_7404,N_10748);
and U14964 (N_14964,N_10314,N_10601);
nor U14965 (N_14965,N_11877,N_10718);
xor U14966 (N_14966,N_10149,N_10918);
and U14967 (N_14967,N_9992,N_11994);
nor U14968 (N_14968,N_7921,N_11277);
nand U14969 (N_14969,N_9244,N_6739);
nor U14970 (N_14970,N_8057,N_10305);
xnor U14971 (N_14971,N_10362,N_10288);
xor U14972 (N_14972,N_9142,N_8436);
nor U14973 (N_14973,N_9878,N_8402);
or U14974 (N_14974,N_11125,N_6301);
or U14975 (N_14975,N_9301,N_11942);
nor U14976 (N_14976,N_7583,N_9754);
nor U14977 (N_14977,N_8699,N_8849);
nor U14978 (N_14978,N_10264,N_11542);
nor U14979 (N_14979,N_6451,N_10435);
nor U14980 (N_14980,N_9227,N_7082);
and U14981 (N_14981,N_9547,N_8916);
xor U14982 (N_14982,N_11057,N_9195);
or U14983 (N_14983,N_8553,N_6628);
and U14984 (N_14984,N_11841,N_12200);
nand U14985 (N_14985,N_9059,N_10216);
and U14986 (N_14986,N_11855,N_8032);
nand U14987 (N_14987,N_8079,N_10713);
nor U14988 (N_14988,N_9504,N_7555);
xor U14989 (N_14989,N_10985,N_11436);
nor U14990 (N_14990,N_11093,N_8318);
nand U14991 (N_14991,N_7024,N_6839);
nand U14992 (N_14992,N_6581,N_7192);
xor U14993 (N_14993,N_9833,N_7825);
and U14994 (N_14994,N_11137,N_6434);
or U14995 (N_14995,N_11128,N_9559);
xnor U14996 (N_14996,N_11146,N_8242);
nor U14997 (N_14997,N_8750,N_12470);
or U14998 (N_14998,N_9883,N_11884);
and U14999 (N_14999,N_6493,N_10173);
nor U15000 (N_15000,N_11075,N_11818);
or U15001 (N_15001,N_11896,N_8543);
nand U15002 (N_15002,N_7999,N_9010);
and U15003 (N_15003,N_8243,N_10712);
or U15004 (N_15004,N_6365,N_8091);
nor U15005 (N_15005,N_9398,N_11776);
nand U15006 (N_15006,N_11152,N_6983);
and U15007 (N_15007,N_6263,N_11082);
xnor U15008 (N_15008,N_7231,N_11968);
nand U15009 (N_15009,N_8692,N_7275);
or U15010 (N_15010,N_9332,N_10175);
and U15011 (N_15011,N_10377,N_9702);
nand U15012 (N_15012,N_10283,N_11249);
nor U15013 (N_15013,N_7906,N_6862);
nand U15014 (N_15014,N_6803,N_11888);
xnor U15015 (N_15015,N_7542,N_12262);
and U15016 (N_15016,N_10211,N_9632);
or U15017 (N_15017,N_11703,N_9158);
or U15018 (N_15018,N_8198,N_10191);
or U15019 (N_15019,N_8605,N_8352);
nand U15020 (N_15020,N_7545,N_7205);
or U15021 (N_15021,N_7415,N_10396);
nand U15022 (N_15022,N_11861,N_7758);
nand U15023 (N_15023,N_8575,N_9787);
and U15024 (N_15024,N_10467,N_8948);
nand U15025 (N_15025,N_9395,N_8214);
xor U15026 (N_15026,N_11397,N_6956);
and U15027 (N_15027,N_8325,N_11943);
nor U15028 (N_15028,N_7901,N_10586);
nand U15029 (N_15029,N_8751,N_6606);
or U15030 (N_15030,N_9459,N_7872);
nor U15031 (N_15031,N_7028,N_7453);
or U15032 (N_15032,N_11910,N_8030);
or U15033 (N_15033,N_10049,N_9351);
nor U15034 (N_15034,N_12333,N_9353);
or U15035 (N_15035,N_6397,N_11603);
or U15036 (N_15036,N_9008,N_6537);
nor U15037 (N_15037,N_8646,N_7597);
nor U15038 (N_15038,N_8661,N_8410);
xnor U15039 (N_15039,N_10057,N_11767);
and U15040 (N_15040,N_10622,N_6491);
nand U15041 (N_15041,N_10017,N_10063);
nor U15042 (N_15042,N_7349,N_12125);
or U15043 (N_15043,N_9261,N_9416);
nor U15044 (N_15044,N_8279,N_12039);
nand U15045 (N_15045,N_9129,N_7972);
nand U15046 (N_15046,N_11770,N_8741);
nand U15047 (N_15047,N_11314,N_9976);
and U15048 (N_15048,N_11226,N_9370);
or U15049 (N_15049,N_7405,N_10234);
and U15050 (N_15050,N_9235,N_7243);
and U15051 (N_15051,N_7258,N_8029);
and U15052 (N_15052,N_6841,N_7800);
or U15053 (N_15053,N_6554,N_9719);
nor U15054 (N_15054,N_6885,N_8166);
nand U15055 (N_15055,N_12360,N_10624);
or U15056 (N_15056,N_9352,N_6727);
xnor U15057 (N_15057,N_6612,N_9120);
or U15058 (N_15058,N_12291,N_10969);
xnor U15059 (N_15059,N_10974,N_7119);
nor U15060 (N_15060,N_11926,N_9242);
and U15061 (N_15061,N_12072,N_11147);
nand U15062 (N_15062,N_10795,N_7015);
and U15063 (N_15063,N_7822,N_11786);
nor U15064 (N_15064,N_8239,N_9015);
or U15065 (N_15065,N_6852,N_11083);
nand U15066 (N_15066,N_10951,N_12244);
or U15067 (N_15067,N_11856,N_9929);
xor U15068 (N_15068,N_10161,N_6674);
or U15069 (N_15069,N_10201,N_7635);
and U15070 (N_15070,N_9302,N_11119);
or U15071 (N_15071,N_12017,N_6919);
nand U15072 (N_15072,N_12115,N_12013);
or U15073 (N_15073,N_9482,N_8427);
or U15074 (N_15074,N_6375,N_7511);
nor U15075 (N_15075,N_10117,N_9860);
nor U15076 (N_15076,N_8391,N_12219);
nand U15077 (N_15077,N_7431,N_9356);
and U15078 (N_15078,N_8228,N_10644);
nand U15079 (N_15079,N_6754,N_8379);
and U15080 (N_15080,N_7055,N_10464);
or U15081 (N_15081,N_11677,N_10421);
xor U15082 (N_15082,N_12281,N_11260);
nor U15083 (N_15083,N_11171,N_7182);
nand U15084 (N_15084,N_9763,N_11222);
and U15085 (N_15085,N_6977,N_12313);
or U15086 (N_15086,N_7515,N_6273);
nor U15087 (N_15087,N_7388,N_6687);
nand U15088 (N_15088,N_10227,N_10987);
and U15089 (N_15089,N_9409,N_10158);
and U15090 (N_15090,N_12198,N_6447);
nand U15091 (N_15091,N_7667,N_7083);
or U15092 (N_15092,N_11755,N_10119);
nor U15093 (N_15093,N_9224,N_6458);
nor U15094 (N_15094,N_7757,N_10474);
nor U15095 (N_15095,N_6538,N_10638);
and U15096 (N_15096,N_8927,N_7042);
nand U15097 (N_15097,N_11741,N_8603);
or U15098 (N_15098,N_11544,N_7172);
nand U15099 (N_15099,N_8982,N_9148);
nor U15100 (N_15100,N_12323,N_9665);
or U15101 (N_15101,N_7547,N_11938);
nand U15102 (N_15102,N_11984,N_8562);
or U15103 (N_15103,N_7207,N_8932);
nor U15104 (N_15104,N_10948,N_11498);
nor U15105 (N_15105,N_11815,N_11241);
or U15106 (N_15106,N_7873,N_10430);
xor U15107 (N_15107,N_9963,N_10760);
nor U15108 (N_15108,N_9796,N_10821);
or U15109 (N_15109,N_9312,N_8788);
or U15110 (N_15110,N_12117,N_8881);
and U15111 (N_15111,N_8740,N_11933);
and U15112 (N_15112,N_8580,N_10456);
nand U15113 (N_15113,N_10499,N_10980);
or U15114 (N_15114,N_6267,N_11768);
nand U15115 (N_15115,N_6831,N_7915);
or U15116 (N_15116,N_9320,N_11097);
xor U15117 (N_15117,N_7821,N_9303);
and U15118 (N_15118,N_10384,N_9453);
nand U15119 (N_15119,N_11374,N_7328);
and U15120 (N_15120,N_10122,N_8721);
or U15121 (N_15121,N_8126,N_6585);
nor U15122 (N_15122,N_7812,N_9732);
xnor U15123 (N_15123,N_8567,N_9100);
nand U15124 (N_15124,N_7688,N_10112);
and U15125 (N_15125,N_6251,N_6781);
nor U15126 (N_15126,N_6859,N_7286);
or U15127 (N_15127,N_10151,N_6668);
nand U15128 (N_15128,N_10625,N_9441);
or U15129 (N_15129,N_12128,N_11626);
or U15130 (N_15130,N_10660,N_11973);
or U15131 (N_15131,N_9942,N_6442);
nand U15132 (N_15132,N_9243,N_12145);
and U15133 (N_15133,N_6682,N_6686);
and U15134 (N_15134,N_10026,N_8173);
or U15135 (N_15135,N_11863,N_10169);
nor U15136 (N_15136,N_10480,N_11474);
nand U15137 (N_15137,N_6970,N_11886);
xor U15138 (N_15138,N_11660,N_6347);
nand U15139 (N_15139,N_9252,N_11301);
nand U15140 (N_15140,N_12106,N_12247);
nor U15141 (N_15141,N_8437,N_11743);
nor U15142 (N_15142,N_10717,N_11080);
nor U15143 (N_15143,N_9949,N_9641);
nor U15144 (N_15144,N_11506,N_11789);
nand U15145 (N_15145,N_7219,N_6717);
and U15146 (N_15146,N_7166,N_10011);
nand U15147 (N_15147,N_12368,N_7303);
and U15148 (N_15148,N_6978,N_8328);
and U15149 (N_15149,N_10533,N_8248);
and U15150 (N_15150,N_8697,N_8642);
nor U15151 (N_15151,N_9757,N_11704);
and U15152 (N_15152,N_9137,N_12417);
nor U15153 (N_15153,N_11719,N_10335);
and U15154 (N_15154,N_7657,N_6735);
and U15155 (N_15155,N_8582,N_12037);
nor U15156 (N_15156,N_8820,N_9274);
and U15157 (N_15157,N_10152,N_6769);
nor U15158 (N_15158,N_8607,N_7850);
nand U15159 (N_15159,N_7985,N_6992);
nor U15160 (N_15160,N_10042,N_10696);
nor U15161 (N_15161,N_7577,N_10199);
and U15162 (N_15162,N_9047,N_9593);
nand U15163 (N_15163,N_11982,N_10000);
and U15164 (N_15164,N_6553,N_11912);
or U15165 (N_15165,N_6352,N_9598);
nor U15166 (N_15166,N_8015,N_6571);
nor U15167 (N_15167,N_7308,N_6897);
and U15168 (N_15168,N_8456,N_12152);
xnor U15169 (N_15169,N_11722,N_6358);
nand U15170 (N_15170,N_7705,N_10879);
nand U15171 (N_15171,N_11579,N_7563);
nor U15172 (N_15172,N_7695,N_10436);
or U15173 (N_15173,N_12324,N_9233);
and U15174 (N_15174,N_9744,N_10255);
or U15175 (N_15175,N_7053,N_11001);
or U15176 (N_15176,N_6857,N_12480);
nor U15177 (N_15177,N_11578,N_8615);
nand U15178 (N_15178,N_8056,N_11810);
or U15179 (N_15179,N_6605,N_7840);
nor U15180 (N_15180,N_9984,N_10738);
nor U15181 (N_15181,N_9119,N_8068);
or U15182 (N_15182,N_7289,N_6572);
and U15183 (N_15183,N_11316,N_11821);
or U15184 (N_15184,N_11785,N_11275);
and U15185 (N_15185,N_9327,N_12206);
or U15186 (N_15186,N_6771,N_7924);
nor U15187 (N_15187,N_10697,N_7189);
xnor U15188 (N_15188,N_11348,N_11209);
nor U15189 (N_15189,N_7041,N_10581);
and U15190 (N_15190,N_11130,N_9138);
xnor U15191 (N_15191,N_10707,N_7817);
and U15192 (N_15192,N_8356,N_11709);
or U15193 (N_15193,N_8767,N_9184);
nand U15194 (N_15194,N_6920,N_9181);
and U15195 (N_15195,N_12003,N_12314);
xor U15196 (N_15196,N_9432,N_9297);
nor U15197 (N_15197,N_8846,N_12040);
and U15198 (N_15198,N_7506,N_7421);
or U15199 (N_15199,N_10055,N_11411);
or U15200 (N_15200,N_7661,N_10135);
nand U15201 (N_15201,N_10303,N_11879);
and U15202 (N_15202,N_6869,N_7077);
or U15203 (N_15203,N_9613,N_10093);
nor U15204 (N_15204,N_6488,N_10594);
nand U15205 (N_15205,N_6665,N_7461);
nand U15206 (N_15206,N_8885,N_7936);
nor U15207 (N_15207,N_6391,N_8685);
and U15208 (N_15208,N_9821,N_10749);
nand U15209 (N_15209,N_6707,N_8569);
nor U15210 (N_15210,N_10570,N_7668);
xnor U15211 (N_15211,N_6669,N_6767);
and U15212 (N_15212,N_11919,N_11325);
nor U15213 (N_15213,N_8260,N_10181);
or U15214 (N_15214,N_10239,N_7697);
nor U15215 (N_15215,N_11750,N_11570);
or U15216 (N_15216,N_12192,N_8088);
nor U15217 (N_15217,N_11278,N_8442);
nor U15218 (N_15218,N_12076,N_7472);
or U15219 (N_15219,N_6753,N_12232);
nor U15220 (N_15220,N_12388,N_11046);
xor U15221 (N_15221,N_9146,N_9934);
and U15222 (N_15222,N_11633,N_12453);
nor U15223 (N_15223,N_6309,N_8085);
nand U15224 (N_15224,N_9549,N_9986);
and U15225 (N_15225,N_7808,N_6331);
nand U15226 (N_15226,N_8549,N_9938);
and U15227 (N_15227,N_9990,N_9950);
nand U15228 (N_15228,N_11493,N_10225);
and U15229 (N_15229,N_8290,N_11966);
and U15230 (N_15230,N_10786,N_10569);
or U15231 (N_15231,N_8627,N_10754);
or U15232 (N_15232,N_9951,N_7090);
nand U15233 (N_15233,N_8673,N_10557);
and U15234 (N_15234,N_8048,N_8185);
nor U15235 (N_15235,N_8816,N_10153);
nand U15236 (N_15236,N_10479,N_7594);
nor U15237 (N_15237,N_6483,N_7299);
nor U15238 (N_15238,N_11915,N_11610);
or U15239 (N_15239,N_12390,N_12499);
and U15240 (N_15240,N_6424,N_6336);
or U15241 (N_15241,N_10582,N_11889);
nor U15242 (N_15242,N_8210,N_7932);
nor U15243 (N_15243,N_11824,N_11769);
and U15244 (N_15244,N_8137,N_6838);
or U15245 (N_15245,N_11654,N_7802);
nor U15246 (N_15246,N_6310,N_11155);
nor U15247 (N_15247,N_9171,N_7530);
nand U15248 (N_15248,N_10315,N_11983);
nor U15249 (N_15249,N_8501,N_7704);
nand U15250 (N_15250,N_11185,N_7638);
and U15251 (N_15251,N_8062,N_9387);
nor U15252 (N_15252,N_9572,N_7785);
nand U15253 (N_15253,N_6418,N_10639);
and U15254 (N_15254,N_11569,N_10507);
nor U15255 (N_15255,N_8168,N_10514);
nand U15256 (N_15256,N_6760,N_12023);
and U15257 (N_15257,N_8997,N_8329);
nor U15258 (N_15258,N_10206,N_8465);
or U15259 (N_15259,N_8877,N_11663);
nand U15260 (N_15260,N_10431,N_7288);
nor U15261 (N_15261,N_11891,N_7551);
nand U15262 (N_15262,N_7726,N_6724);
xor U15263 (N_15263,N_11208,N_7305);
nand U15264 (N_15264,N_9400,N_10077);
and U15265 (N_15265,N_8635,N_7781);
nor U15266 (N_15266,N_10247,N_8981);
or U15267 (N_15267,N_8908,N_10407);
and U15268 (N_15268,N_11620,N_11019);
and U15269 (N_15269,N_11026,N_11482);
xor U15270 (N_15270,N_6805,N_7686);
and U15271 (N_15271,N_7098,N_6928);
nor U15272 (N_15272,N_12369,N_7629);
and U15273 (N_15273,N_11634,N_12073);
and U15274 (N_15274,N_10693,N_9972);
nor U15275 (N_15275,N_10150,N_9081);
and U15276 (N_15276,N_6875,N_8333);
or U15277 (N_15277,N_12475,N_7492);
or U15278 (N_15278,N_10072,N_7868);
or U15279 (N_15279,N_10555,N_8300);
or U15280 (N_15280,N_7837,N_10062);
or U15281 (N_15281,N_9365,N_12230);
xor U15282 (N_15282,N_10943,N_9708);
nand U15283 (N_15283,N_6480,N_8474);
or U15284 (N_15284,N_7035,N_10237);
and U15285 (N_15285,N_11223,N_7763);
and U15286 (N_15286,N_11283,N_7362);
or U15287 (N_15287,N_7244,N_9568);
nand U15288 (N_15288,N_7675,N_6695);
or U15289 (N_15289,N_11989,N_11154);
nand U15290 (N_15290,N_6962,N_10131);
and U15291 (N_15291,N_9045,N_8310);
nor U15292 (N_15292,N_12114,N_6672);
and U15293 (N_15293,N_7325,N_9886);
nand U15294 (N_15294,N_6298,N_11485);
or U15295 (N_15295,N_9638,N_7073);
xnor U15296 (N_15296,N_10353,N_6294);
nand U15297 (N_15297,N_9745,N_12287);
nor U15298 (N_15298,N_9480,N_10953);
and U15299 (N_15299,N_8931,N_9689);
nand U15300 (N_15300,N_8935,N_11533);
nand U15301 (N_15301,N_6522,N_10278);
nand U15302 (N_15302,N_9461,N_11748);
or U15303 (N_15303,N_10092,N_8255);
and U15304 (N_15304,N_9220,N_6974);
or U15305 (N_15305,N_11144,N_8722);
nor U15306 (N_15306,N_8218,N_8828);
nor U15307 (N_15307,N_7191,N_8998);
nor U15308 (N_15308,N_11974,N_11354);
or U15309 (N_15309,N_10546,N_6710);
nand U15310 (N_15310,N_6991,N_12083);
nor U15311 (N_15311,N_10885,N_7267);
nand U15312 (N_15312,N_11315,N_6915);
nand U15313 (N_15313,N_10048,N_8359);
or U15314 (N_15314,N_10558,N_12210);
nand U15315 (N_15315,N_12348,N_9783);
and U15316 (N_15316,N_10762,N_12457);
nor U15317 (N_15317,N_9131,N_9674);
or U15318 (N_15318,N_12359,N_10344);
xnor U15319 (N_15319,N_7385,N_12459);
or U15320 (N_15320,N_11136,N_11369);
nand U15321 (N_15321,N_9601,N_6399);
and U15322 (N_15322,N_9980,N_9890);
and U15323 (N_15323,N_7912,N_8848);
xnor U15324 (N_15324,N_10618,N_10891);
nor U15325 (N_15325,N_7654,N_10645);
nor U15326 (N_15326,N_11615,N_7809);
nand U15327 (N_15327,N_7609,N_7412);
nor U15328 (N_15328,N_10148,N_10261);
nand U15329 (N_15329,N_8937,N_10035);
xnor U15330 (N_15330,N_10833,N_11744);
or U15331 (N_15331,N_9916,N_8648);
nor U15332 (N_15332,N_12071,N_10379);
or U15333 (N_15333,N_6595,N_9428);
xor U15334 (N_15334,N_12266,N_10455);
nand U15335 (N_15335,N_6306,N_9912);
or U15336 (N_15336,N_10364,N_6701);
and U15337 (N_15337,N_7296,N_7740);
and U15338 (N_15338,N_10883,N_10185);
nand U15339 (N_15339,N_7979,N_6255);
nand U15340 (N_15340,N_11651,N_12242);
and U15341 (N_15341,N_11007,N_8806);
nand U15342 (N_15342,N_9410,N_9057);
and U15343 (N_15343,N_11515,N_9592);
and U15344 (N_15344,N_7741,N_8835);
nand U15345 (N_15345,N_7617,N_11470);
or U15346 (N_15346,N_10984,N_12078);
or U15347 (N_15347,N_6909,N_8734);
nand U15348 (N_15348,N_7535,N_11986);
and U15349 (N_15349,N_8653,N_7831);
nand U15350 (N_15350,N_8345,N_8367);
and U15351 (N_15351,N_12220,N_8366);
xor U15352 (N_15352,N_9223,N_8283);
nor U15353 (N_15353,N_9161,N_10658);
and U15354 (N_15354,N_8727,N_10050);
nor U15355 (N_15355,N_9532,N_7157);
nor U15356 (N_15356,N_8211,N_11921);
nor U15357 (N_15357,N_11955,N_10611);
or U15358 (N_15358,N_6601,N_6381);
nand U15359 (N_15359,N_6319,N_9596);
nor U15360 (N_15360,N_10574,N_6290);
xor U15361 (N_15361,N_6527,N_10550);
and U15362 (N_15362,N_8489,N_9718);
and U15363 (N_15363,N_7227,N_6851);
xor U15364 (N_15364,N_6975,N_7517);
xor U15365 (N_15365,N_11446,N_9953);
nor U15366 (N_15366,N_9455,N_10783);
nand U15367 (N_15367,N_7552,N_7068);
and U15368 (N_15368,N_11550,N_6597);
nand U15369 (N_15369,N_11159,N_9616);
and U15370 (N_15370,N_6355,N_10144);
and U15371 (N_15371,N_7324,N_11313);
nand U15372 (N_15372,N_11518,N_6330);
or U15373 (N_15373,N_10541,N_8195);
nor U15374 (N_15374,N_9496,N_12133);
nand U15375 (N_15375,N_9870,N_6454);
or U15376 (N_15376,N_10240,N_9831);
nor U15377 (N_15377,N_11947,N_9499);
nor U15378 (N_15378,N_11176,N_9484);
nor U15379 (N_15379,N_7893,N_8898);
xor U15380 (N_15380,N_8608,N_9182);
and U15381 (N_15381,N_10336,N_10898);
nor U15382 (N_15382,N_12481,N_6855);
xor U15383 (N_15383,N_6900,N_12354);
and U15384 (N_15384,N_12462,N_7902);
xnor U15385 (N_15385,N_12151,N_10476);
or U15386 (N_15386,N_10290,N_10438);
nand U15387 (N_15387,N_7766,N_8430);
nand U15388 (N_15388,N_7926,N_8115);
nand U15389 (N_15389,N_7789,N_9464);
or U15390 (N_15390,N_10218,N_9743);
nor U15391 (N_15391,N_12140,N_12434);
nand U15392 (N_15392,N_9589,N_10663);
nor U15393 (N_15393,N_10109,N_8643);
nand U15394 (N_15394,N_9756,N_11416);
xnor U15395 (N_15395,N_8571,N_11604);
nand U15396 (N_15396,N_8340,N_6741);
and U15397 (N_15397,N_10317,N_10841);
nand U15398 (N_15398,N_12138,N_11458);
xor U15399 (N_15399,N_9642,N_7374);
nor U15400 (N_15400,N_12399,N_9278);
xnor U15401 (N_15401,N_7672,N_12250);
and U15402 (N_15402,N_9713,N_9230);
and U15403 (N_15403,N_10595,N_8680);
nor U15404 (N_15404,N_9609,N_10360);
and U15405 (N_15405,N_10819,N_6422);
nor U15406 (N_15406,N_9253,N_6766);
or U15407 (N_15407,N_6936,N_12202);
nor U15408 (N_15408,N_7319,N_11600);
nand U15409 (N_15409,N_10069,N_7111);
nand U15410 (N_15410,N_10843,N_6750);
or U15411 (N_15411,N_10434,N_12122);
nor U15412 (N_15412,N_7911,N_8455);
nand U15413 (N_15413,N_7211,N_9102);
or U15414 (N_15414,N_11341,N_11737);
nor U15415 (N_15415,N_10354,N_6464);
and U15416 (N_15416,N_9881,N_8769);
and U15417 (N_15417,N_9551,N_11540);
nand U15418 (N_15418,N_11480,N_11248);
xnor U15419 (N_15419,N_7674,N_10609);
and U15420 (N_15420,N_12015,N_9069);
nand U15421 (N_15421,N_12370,N_10740);
and U15422 (N_15422,N_11459,N_7645);
xor U15423 (N_15423,N_11795,N_7869);
nor U15424 (N_15424,N_8922,N_7579);
nand U15425 (N_15425,N_7768,N_6332);
nand U15426 (N_15426,N_7427,N_8120);
and U15427 (N_15427,N_8044,N_11467);
xnor U15428 (N_15428,N_8844,N_11490);
and U15429 (N_15429,N_8118,N_9967);
nor U15430 (N_15430,N_10302,N_6676);
and U15431 (N_15431,N_10769,N_8343);
nand U15432 (N_15432,N_9170,N_6593);
xnor U15433 (N_15433,N_10252,N_9442);
or U15434 (N_15434,N_9172,N_7449);
and U15435 (N_15435,N_7352,N_11759);
or U15436 (N_15436,N_10321,N_9399);
and U15437 (N_15437,N_8901,N_10127);
or U15438 (N_15438,N_8065,N_8199);
nor U15439 (N_15439,N_7782,N_9288);
or U15440 (N_15440,N_6376,N_6673);
and U15441 (N_15441,N_8859,N_7000);
nand U15442 (N_15442,N_7724,N_11045);
xor U15443 (N_15443,N_11524,N_11564);
and U15444 (N_15444,N_7464,N_11179);
or U15445 (N_15445,N_8229,N_11587);
and U15446 (N_15446,N_11500,N_6295);
nand U15447 (N_15447,N_8838,N_11151);
or U15448 (N_15448,N_8148,N_9341);
nor U15449 (N_15449,N_6965,N_7737);
or U15450 (N_15450,N_8731,N_6652);
xor U15451 (N_15451,N_8074,N_11792);
nor U15452 (N_15452,N_10323,N_7725);
nor U15453 (N_15453,N_9648,N_7318);
xor U15454 (N_15454,N_11967,N_8133);
or U15455 (N_15455,N_11757,N_10565);
nand U15456 (N_15456,N_7569,N_9872);
xnor U15457 (N_15457,N_7133,N_8616);
xnor U15458 (N_15458,N_10688,N_10995);
and U15459 (N_15459,N_7655,N_10342);
nand U15460 (N_15460,N_11198,N_10389);
and U15461 (N_15461,N_12094,N_9444);
nor U15462 (N_15462,N_9940,N_11186);
and U15463 (N_15463,N_6276,N_10659);
or U15464 (N_15464,N_8689,N_9628);
or U15465 (N_15465,N_11328,N_6709);
nor U15466 (N_15466,N_9051,N_8577);
nor U15467 (N_15467,N_7838,N_9494);
nand U15468 (N_15468,N_9372,N_10285);
nand U15469 (N_15469,N_9581,N_9602);
nor U15470 (N_15470,N_11903,N_6504);
nand U15471 (N_15471,N_9042,N_9221);
and U15472 (N_15472,N_10604,N_9862);
and U15473 (N_15473,N_9838,N_6469);
nor U15474 (N_15474,N_6960,N_6662);
xor U15475 (N_15475,N_10549,N_11050);
nor U15476 (N_15476,N_10068,N_7407);
or U15477 (N_15477,N_7484,N_11688);
xnor U15478 (N_15478,N_11864,N_8745);
xor U15479 (N_15479,N_10677,N_12229);
or U15480 (N_15480,N_6444,N_7281);
nand U15481 (N_15481,N_9611,N_10959);
or U15482 (N_15482,N_6677,N_11529);
nor U15483 (N_15483,N_10418,N_11158);
nor U15484 (N_15484,N_11981,N_6567);
or U15485 (N_15485,N_9248,N_10195);
nor U15486 (N_15486,N_12016,N_8617);
xnor U15487 (N_15487,N_11013,N_10692);
or U15488 (N_15488,N_11102,N_11669);
and U15489 (N_15489,N_10348,N_8792);
nand U15490 (N_15490,N_6721,N_7576);
or U15491 (N_15491,N_6944,N_8677);
nor U15492 (N_15492,N_11720,N_12178);
nor U15493 (N_15493,N_12436,N_8506);
and U15494 (N_15494,N_8893,N_8051);
and U15495 (N_15495,N_7446,N_8454);
nor U15496 (N_15496,N_6679,N_6664);
nand U15497 (N_15497,N_10107,N_7280);
or U15498 (N_15498,N_10534,N_10472);
nor U15499 (N_15499,N_11628,N_7037);
or U15500 (N_15500,N_8679,N_10440);
or U15501 (N_15501,N_7942,N_8475);
xor U15502 (N_15502,N_9314,N_12018);
nand U15503 (N_15503,N_6366,N_11621);
nand U15504 (N_15504,N_12293,N_12064);
nand U15505 (N_15505,N_6289,N_7955);
and U15506 (N_15506,N_8911,N_7292);
and U15507 (N_15507,N_7382,N_8116);
nor U15508 (N_15508,N_6322,N_8865);
nand U15509 (N_15509,N_10043,N_8299);
nand U15510 (N_15510,N_6382,N_6683);
or U15511 (N_15511,N_11358,N_12086);
and U15512 (N_15512,N_10735,N_8597);
and U15513 (N_15513,N_9774,N_10647);
nor U15514 (N_15514,N_8832,N_11335);
nand U15515 (N_15515,N_6800,N_8598);
xnor U15516 (N_15516,N_9537,N_9888);
nor U15517 (N_15517,N_8357,N_11207);
nand U15518 (N_15518,N_11627,N_11258);
and U15519 (N_15519,N_12300,N_7864);
or U15520 (N_15520,N_6379,N_10648);
and U15521 (N_15521,N_9135,N_11037);
or U15522 (N_15522,N_7931,N_10934);
nor U15523 (N_15523,N_9130,N_10219);
nor U15524 (N_15524,N_11340,N_11887);
and U15525 (N_15525,N_7929,N_8955);
and U15526 (N_15526,N_10635,N_11640);
nor U15527 (N_15527,N_9412,N_11199);
and U15528 (N_15528,N_10860,N_6957);
or U15529 (N_15529,N_9711,N_6793);
or U15530 (N_15530,N_7959,N_8271);
or U15531 (N_15531,N_8839,N_9405);
nand U15532 (N_15532,N_10086,N_7463);
or U15533 (N_15533,N_11925,N_8517);
and U15534 (N_15534,N_7993,N_6726);
or U15535 (N_15535,N_10382,N_9849);
nor U15536 (N_15536,N_11069,N_6525);
nor U15537 (N_15537,N_9829,N_8586);
xor U15538 (N_15538,N_9357,N_6819);
nand U15539 (N_15539,N_7439,N_6436);
nor U15540 (N_15540,N_8614,N_9462);
nand U15541 (N_15541,N_9503,N_10424);
and U15542 (N_15542,N_8451,N_9695);
nand U15543 (N_15543,N_7417,N_6698);
nand U15544 (N_15544,N_7641,N_12032);
or U15545 (N_15545,N_11006,N_12214);
nand U15546 (N_15546,N_6300,N_7246);
or U15547 (N_15547,N_6784,N_8915);
and U15548 (N_15548,N_6311,N_12069);
nor U15549 (N_15549,N_7441,N_6615);
nor U15550 (N_15550,N_8045,N_8735);
nand U15551 (N_15551,N_8746,N_8851);
or U15552 (N_15552,N_7386,N_11404);
nand U15553 (N_15553,N_6435,N_8829);
nor U15554 (N_15554,N_6386,N_6270);
nand U15555 (N_15555,N_6810,N_11866);
nand U15556 (N_15556,N_6367,N_12095);
nor U15557 (N_15557,N_11988,N_11537);
or U15558 (N_15558,N_8887,N_8546);
or U15559 (N_15559,N_12292,N_10669);
and U15560 (N_15560,N_8515,N_11469);
or U15561 (N_15561,N_12414,N_9070);
and U15562 (N_15562,N_7690,N_8533);
and U15563 (N_15563,N_6555,N_10187);
nor U15564 (N_15564,N_7557,N_7685);
and U15565 (N_15565,N_12340,N_6967);
or U15566 (N_15566,N_8092,N_10964);
and U15567 (N_15567,N_11100,N_7776);
nor U15568 (N_15568,N_9108,N_10627);
and U15569 (N_15569,N_12377,N_11225);
or U15570 (N_15570,N_7048,N_10928);
nand U15571 (N_15571,N_11499,N_7953);
xnor U15572 (N_15572,N_12103,N_11860);
and U15573 (N_15573,N_8914,N_10034);
nand U15574 (N_15574,N_6870,N_8178);
or U15575 (N_15575,N_6866,N_9682);
nor U15576 (N_15576,N_8524,N_11508);
nor U15577 (N_15577,N_11000,N_6551);
nor U15578 (N_15578,N_11244,N_7900);
and U15579 (N_15579,N_10882,N_12427);
nor U15580 (N_15580,N_6515,N_10798);
or U15581 (N_15581,N_9325,N_7327);
or U15582 (N_15582,N_8744,N_11371);
or U15583 (N_15583,N_11291,N_11373);
nor U15584 (N_15584,N_10368,N_7536);
and U15585 (N_15585,N_6374,N_8230);
nor U15586 (N_15586,N_11409,N_6829);
nor U15587 (N_15587,N_7079,N_10374);
nand U15588 (N_15588,N_8176,N_7773);
and U15589 (N_15589,N_7196,N_8444);
and U15590 (N_15590,N_7870,N_6618);
or U15591 (N_15591,N_9381,N_11952);
or U15592 (N_15592,N_7988,N_9776);
or U15593 (N_15593,N_9147,N_8812);
nand U15594 (N_15594,N_12471,N_12021);
nor U15595 (N_15595,N_6997,N_9690);
or U15596 (N_15596,N_10065,N_8866);
and U15597 (N_15597,N_6576,N_12373);
nand U15598 (N_15598,N_10770,N_7071);
nor U15599 (N_15599,N_6489,N_8664);
or U15600 (N_15600,N_9099,N_8187);
or U15601 (N_15601,N_9884,N_7520);
and U15602 (N_15602,N_11764,N_7186);
nand U15603 (N_15603,N_12158,N_6826);
and U15604 (N_15604,N_12492,N_8576);
nor U15605 (N_15605,N_6715,N_12332);
and U15606 (N_15606,N_8514,N_12030);
nor U15607 (N_15607,N_8716,N_9075);
and U15608 (N_15608,N_8890,N_11740);
nor U15609 (N_15609,N_6783,N_6325);
and U15610 (N_15610,N_7268,N_8842);
or U15611 (N_15611,N_7752,N_11218);
nor U15612 (N_15612,N_12098,N_7927);
and U15613 (N_15613,N_6474,N_11820);
nand U15614 (N_15614,N_7422,N_12411);
and U15615 (N_15615,N_9919,N_6888);
and U15616 (N_15616,N_9087,N_6971);
or U15617 (N_15617,N_8009,N_10398);
xnor U15618 (N_15618,N_11253,N_8644);
nor U15619 (N_15619,N_12275,N_6262);
and U15620 (N_15620,N_7081,N_11637);
and U15621 (N_15621,N_6439,N_11466);
nand U15622 (N_15622,N_12441,N_9541);
nand U15623 (N_15623,N_7007,N_8149);
or U15624 (N_15624,N_11098,N_8331);
or U15625 (N_15625,N_10194,N_7148);
nand U15626 (N_15626,N_6602,N_6371);
nand U15627 (N_15627,N_7337,N_11780);
and U15628 (N_15628,N_8312,N_6575);
or U15629 (N_15629,N_9884,N_8745);
or U15630 (N_15630,N_8899,N_6633);
or U15631 (N_15631,N_10199,N_11732);
nand U15632 (N_15632,N_10973,N_12308);
nand U15633 (N_15633,N_7897,N_11052);
or U15634 (N_15634,N_9626,N_10497);
and U15635 (N_15635,N_8080,N_6443);
nor U15636 (N_15636,N_9774,N_7054);
nand U15637 (N_15637,N_10153,N_10402);
nor U15638 (N_15638,N_6697,N_8650);
nand U15639 (N_15639,N_12294,N_11074);
and U15640 (N_15640,N_10272,N_8383);
and U15641 (N_15641,N_6304,N_7913);
nand U15642 (N_15642,N_10852,N_9504);
or U15643 (N_15643,N_8218,N_11990);
nor U15644 (N_15644,N_7077,N_12181);
nor U15645 (N_15645,N_10215,N_9167);
nor U15646 (N_15646,N_6972,N_8417);
nand U15647 (N_15647,N_6944,N_12002);
nand U15648 (N_15648,N_7532,N_11775);
nand U15649 (N_15649,N_7035,N_10742);
and U15650 (N_15650,N_9674,N_6301);
or U15651 (N_15651,N_9214,N_7889);
nor U15652 (N_15652,N_7286,N_11789);
or U15653 (N_15653,N_11599,N_7161);
nor U15654 (N_15654,N_11224,N_12386);
or U15655 (N_15655,N_10222,N_9976);
nand U15656 (N_15656,N_10323,N_11866);
nor U15657 (N_15657,N_11346,N_9147);
nor U15658 (N_15658,N_10315,N_11226);
and U15659 (N_15659,N_9594,N_9210);
nor U15660 (N_15660,N_9517,N_6322);
nand U15661 (N_15661,N_7363,N_6605);
and U15662 (N_15662,N_9042,N_8446);
or U15663 (N_15663,N_10697,N_9509);
nor U15664 (N_15664,N_9026,N_9952);
nor U15665 (N_15665,N_12179,N_8863);
and U15666 (N_15666,N_9100,N_6977);
xnor U15667 (N_15667,N_10961,N_8231);
and U15668 (N_15668,N_8151,N_6654);
nand U15669 (N_15669,N_12289,N_7228);
and U15670 (N_15670,N_9083,N_11740);
and U15671 (N_15671,N_8938,N_8133);
nor U15672 (N_15672,N_8488,N_7736);
and U15673 (N_15673,N_7718,N_7953);
and U15674 (N_15674,N_9033,N_8997);
xnor U15675 (N_15675,N_7390,N_8174);
nand U15676 (N_15676,N_9187,N_7180);
nand U15677 (N_15677,N_7682,N_8376);
or U15678 (N_15678,N_6449,N_10455);
nand U15679 (N_15679,N_11357,N_9144);
nand U15680 (N_15680,N_6944,N_6395);
or U15681 (N_15681,N_10825,N_10169);
nand U15682 (N_15682,N_10257,N_10505);
xnor U15683 (N_15683,N_11496,N_8538);
and U15684 (N_15684,N_7154,N_8992);
and U15685 (N_15685,N_6550,N_12483);
and U15686 (N_15686,N_8586,N_6384);
nor U15687 (N_15687,N_11070,N_11304);
nor U15688 (N_15688,N_10599,N_7133);
or U15689 (N_15689,N_9275,N_11433);
nand U15690 (N_15690,N_7545,N_7453);
and U15691 (N_15691,N_6258,N_7112);
nor U15692 (N_15692,N_11858,N_12114);
or U15693 (N_15693,N_9121,N_10675);
or U15694 (N_15694,N_11780,N_6828);
xor U15695 (N_15695,N_6947,N_12332);
and U15696 (N_15696,N_10341,N_9419);
nand U15697 (N_15697,N_10165,N_6947);
or U15698 (N_15698,N_8519,N_9765);
xnor U15699 (N_15699,N_8565,N_10148);
nor U15700 (N_15700,N_11248,N_7200);
and U15701 (N_15701,N_8305,N_9728);
nand U15702 (N_15702,N_7385,N_8693);
xor U15703 (N_15703,N_10872,N_12278);
nor U15704 (N_15704,N_10530,N_11686);
or U15705 (N_15705,N_7425,N_10274);
nor U15706 (N_15706,N_10333,N_6658);
and U15707 (N_15707,N_10912,N_6394);
xor U15708 (N_15708,N_6984,N_9668);
or U15709 (N_15709,N_7520,N_8928);
nand U15710 (N_15710,N_8932,N_11660);
and U15711 (N_15711,N_6299,N_9022);
or U15712 (N_15712,N_9736,N_11697);
nor U15713 (N_15713,N_11800,N_9111);
nor U15714 (N_15714,N_6449,N_6882);
or U15715 (N_15715,N_7289,N_8374);
or U15716 (N_15716,N_10507,N_6302);
nand U15717 (N_15717,N_9362,N_11066);
and U15718 (N_15718,N_6303,N_10331);
nor U15719 (N_15719,N_9559,N_11974);
xor U15720 (N_15720,N_12226,N_12254);
nor U15721 (N_15721,N_7293,N_11027);
xnor U15722 (N_15722,N_7955,N_9644);
and U15723 (N_15723,N_6543,N_12053);
or U15724 (N_15724,N_7603,N_7580);
and U15725 (N_15725,N_10157,N_7576);
nand U15726 (N_15726,N_11386,N_9294);
and U15727 (N_15727,N_8058,N_9334);
and U15728 (N_15728,N_8255,N_11795);
or U15729 (N_15729,N_9972,N_6375);
nand U15730 (N_15730,N_10239,N_10353);
nor U15731 (N_15731,N_10632,N_10934);
nor U15732 (N_15732,N_9582,N_9452);
and U15733 (N_15733,N_9855,N_8720);
or U15734 (N_15734,N_6318,N_10984);
nand U15735 (N_15735,N_8520,N_8241);
and U15736 (N_15736,N_11456,N_7213);
nor U15737 (N_15737,N_10637,N_7136);
nor U15738 (N_15738,N_8741,N_11251);
or U15739 (N_15739,N_8545,N_10023);
and U15740 (N_15740,N_6288,N_8968);
and U15741 (N_15741,N_11099,N_8026);
or U15742 (N_15742,N_6853,N_9640);
or U15743 (N_15743,N_8164,N_9480);
nor U15744 (N_15744,N_11841,N_7089);
and U15745 (N_15745,N_8942,N_6775);
nand U15746 (N_15746,N_8775,N_7014);
nor U15747 (N_15747,N_10409,N_11190);
nor U15748 (N_15748,N_10099,N_9704);
or U15749 (N_15749,N_6408,N_12370);
or U15750 (N_15750,N_11942,N_12055);
nand U15751 (N_15751,N_12021,N_11782);
nand U15752 (N_15752,N_7190,N_7737);
nor U15753 (N_15753,N_9093,N_9545);
and U15754 (N_15754,N_11542,N_9982);
or U15755 (N_15755,N_10219,N_12114);
nand U15756 (N_15756,N_8784,N_7683);
nor U15757 (N_15757,N_8610,N_10177);
nand U15758 (N_15758,N_8736,N_11840);
nand U15759 (N_15759,N_8343,N_6333);
nor U15760 (N_15760,N_8660,N_7843);
nand U15761 (N_15761,N_9545,N_11834);
or U15762 (N_15762,N_8236,N_9366);
xnor U15763 (N_15763,N_7145,N_7306);
and U15764 (N_15764,N_7322,N_11079);
nor U15765 (N_15765,N_7632,N_12041);
nand U15766 (N_15766,N_11696,N_6289);
and U15767 (N_15767,N_11133,N_8061);
or U15768 (N_15768,N_9656,N_9867);
and U15769 (N_15769,N_11757,N_9081);
nand U15770 (N_15770,N_10721,N_10199);
nor U15771 (N_15771,N_12303,N_6575);
nand U15772 (N_15772,N_6744,N_6785);
or U15773 (N_15773,N_12248,N_8191);
or U15774 (N_15774,N_10692,N_10147);
nor U15775 (N_15775,N_7458,N_11344);
nor U15776 (N_15776,N_10162,N_9538);
or U15777 (N_15777,N_11494,N_9528);
xor U15778 (N_15778,N_8652,N_10742);
or U15779 (N_15779,N_10244,N_11509);
nor U15780 (N_15780,N_12037,N_10348);
nand U15781 (N_15781,N_7836,N_9004);
or U15782 (N_15782,N_11765,N_12394);
nand U15783 (N_15783,N_11496,N_10939);
nand U15784 (N_15784,N_12408,N_9175);
xor U15785 (N_15785,N_9888,N_10080);
and U15786 (N_15786,N_11203,N_11924);
and U15787 (N_15787,N_11279,N_11332);
and U15788 (N_15788,N_7598,N_8906);
and U15789 (N_15789,N_10620,N_7411);
and U15790 (N_15790,N_6657,N_8126);
nand U15791 (N_15791,N_6678,N_11110);
or U15792 (N_15792,N_11804,N_6919);
and U15793 (N_15793,N_11783,N_11823);
xnor U15794 (N_15794,N_10377,N_9071);
nor U15795 (N_15795,N_9267,N_9613);
and U15796 (N_15796,N_11701,N_10122);
nand U15797 (N_15797,N_7038,N_11431);
nor U15798 (N_15798,N_8892,N_10725);
and U15799 (N_15799,N_10182,N_6866);
nand U15800 (N_15800,N_6795,N_7502);
nor U15801 (N_15801,N_12256,N_10693);
or U15802 (N_15802,N_8985,N_8920);
or U15803 (N_15803,N_11817,N_7836);
or U15804 (N_15804,N_7006,N_7399);
nor U15805 (N_15805,N_11334,N_10719);
nand U15806 (N_15806,N_12369,N_10723);
xnor U15807 (N_15807,N_12347,N_10601);
nor U15808 (N_15808,N_6768,N_7029);
or U15809 (N_15809,N_12192,N_11559);
or U15810 (N_15810,N_9896,N_11974);
nand U15811 (N_15811,N_9769,N_8606);
nand U15812 (N_15812,N_8478,N_12281);
nor U15813 (N_15813,N_7049,N_12439);
and U15814 (N_15814,N_8748,N_7787);
nor U15815 (N_15815,N_7068,N_9495);
or U15816 (N_15816,N_11257,N_7233);
and U15817 (N_15817,N_9173,N_6412);
or U15818 (N_15818,N_12168,N_11145);
nor U15819 (N_15819,N_10958,N_7116);
or U15820 (N_15820,N_6986,N_8967);
and U15821 (N_15821,N_9202,N_10812);
or U15822 (N_15822,N_9211,N_7827);
nand U15823 (N_15823,N_8955,N_7720);
nor U15824 (N_15824,N_8411,N_11711);
xnor U15825 (N_15825,N_7381,N_11505);
and U15826 (N_15826,N_7476,N_10105);
or U15827 (N_15827,N_9231,N_8566);
and U15828 (N_15828,N_7155,N_8409);
and U15829 (N_15829,N_6931,N_8342);
or U15830 (N_15830,N_12105,N_11469);
xnor U15831 (N_15831,N_8796,N_7577);
or U15832 (N_15832,N_9016,N_9970);
nand U15833 (N_15833,N_6461,N_8190);
xor U15834 (N_15834,N_7892,N_8244);
nor U15835 (N_15835,N_10114,N_10936);
xnor U15836 (N_15836,N_11523,N_8609);
nand U15837 (N_15837,N_8155,N_12465);
nor U15838 (N_15838,N_11781,N_6664);
and U15839 (N_15839,N_8660,N_9355);
xor U15840 (N_15840,N_6308,N_6816);
nand U15841 (N_15841,N_8105,N_6896);
nor U15842 (N_15842,N_11056,N_12483);
nor U15843 (N_15843,N_10727,N_8915);
or U15844 (N_15844,N_7509,N_9919);
and U15845 (N_15845,N_10412,N_6808);
or U15846 (N_15846,N_9219,N_8565);
nor U15847 (N_15847,N_11526,N_7822);
nand U15848 (N_15848,N_8053,N_11695);
or U15849 (N_15849,N_10601,N_9114);
xnor U15850 (N_15850,N_10602,N_9077);
and U15851 (N_15851,N_11901,N_10788);
nand U15852 (N_15852,N_6970,N_10581);
xor U15853 (N_15853,N_9391,N_10550);
and U15854 (N_15854,N_11656,N_10848);
and U15855 (N_15855,N_8613,N_7529);
or U15856 (N_15856,N_6436,N_12469);
and U15857 (N_15857,N_8751,N_12199);
nand U15858 (N_15858,N_9393,N_9074);
nor U15859 (N_15859,N_7773,N_9466);
nor U15860 (N_15860,N_8598,N_11345);
or U15861 (N_15861,N_6760,N_6693);
and U15862 (N_15862,N_7348,N_6780);
and U15863 (N_15863,N_10417,N_9387);
and U15864 (N_15864,N_11868,N_10930);
nor U15865 (N_15865,N_9365,N_6633);
nand U15866 (N_15866,N_6987,N_7864);
nor U15867 (N_15867,N_11680,N_7836);
or U15868 (N_15868,N_10605,N_10174);
nand U15869 (N_15869,N_8261,N_7486);
nor U15870 (N_15870,N_8828,N_9104);
or U15871 (N_15871,N_10322,N_9302);
or U15872 (N_15872,N_12282,N_8443);
and U15873 (N_15873,N_10688,N_10983);
nor U15874 (N_15874,N_10489,N_10983);
and U15875 (N_15875,N_9577,N_8433);
nand U15876 (N_15876,N_10922,N_10155);
nand U15877 (N_15877,N_11457,N_10537);
or U15878 (N_15878,N_10357,N_7516);
nand U15879 (N_15879,N_10371,N_11561);
xor U15880 (N_15880,N_7780,N_9428);
or U15881 (N_15881,N_6723,N_8764);
nand U15882 (N_15882,N_12116,N_8229);
nor U15883 (N_15883,N_7289,N_6774);
or U15884 (N_15884,N_10463,N_11665);
xnor U15885 (N_15885,N_7158,N_11598);
nor U15886 (N_15886,N_10774,N_9565);
and U15887 (N_15887,N_7952,N_8550);
or U15888 (N_15888,N_6689,N_10381);
nor U15889 (N_15889,N_12414,N_11331);
and U15890 (N_15890,N_11415,N_7448);
xor U15891 (N_15891,N_9190,N_9317);
or U15892 (N_15892,N_12117,N_7587);
nand U15893 (N_15893,N_8971,N_7586);
nor U15894 (N_15894,N_8876,N_8328);
nor U15895 (N_15895,N_7863,N_10433);
nor U15896 (N_15896,N_8567,N_11312);
or U15897 (N_15897,N_11621,N_7046);
nand U15898 (N_15898,N_7356,N_7657);
xor U15899 (N_15899,N_6927,N_7123);
xnor U15900 (N_15900,N_8161,N_9869);
nor U15901 (N_15901,N_6876,N_10844);
nor U15902 (N_15902,N_8095,N_9714);
and U15903 (N_15903,N_8995,N_12345);
nor U15904 (N_15904,N_8104,N_10833);
nor U15905 (N_15905,N_12334,N_8895);
nor U15906 (N_15906,N_7871,N_7753);
nor U15907 (N_15907,N_11458,N_6401);
or U15908 (N_15908,N_6754,N_6721);
nor U15909 (N_15909,N_6650,N_10170);
nor U15910 (N_15910,N_7745,N_11849);
xnor U15911 (N_15911,N_6346,N_8549);
and U15912 (N_15912,N_10332,N_11720);
nor U15913 (N_15913,N_8443,N_7811);
xor U15914 (N_15914,N_9974,N_11920);
or U15915 (N_15915,N_7230,N_10906);
xnor U15916 (N_15916,N_11285,N_8731);
nand U15917 (N_15917,N_6591,N_11726);
nor U15918 (N_15918,N_7923,N_8259);
and U15919 (N_15919,N_6981,N_6285);
or U15920 (N_15920,N_7158,N_11226);
or U15921 (N_15921,N_8027,N_10908);
and U15922 (N_15922,N_8063,N_10577);
nor U15923 (N_15923,N_8613,N_6310);
nand U15924 (N_15924,N_8046,N_8815);
and U15925 (N_15925,N_8067,N_11569);
and U15926 (N_15926,N_10248,N_8652);
or U15927 (N_15927,N_11460,N_6929);
and U15928 (N_15928,N_11601,N_7239);
nand U15929 (N_15929,N_12482,N_9800);
or U15930 (N_15930,N_6702,N_7271);
nor U15931 (N_15931,N_6741,N_7860);
nand U15932 (N_15932,N_6853,N_10775);
nand U15933 (N_15933,N_11774,N_11347);
nor U15934 (N_15934,N_11354,N_8640);
and U15935 (N_15935,N_10589,N_8219);
nand U15936 (N_15936,N_11147,N_6717);
nand U15937 (N_15937,N_12451,N_9576);
nand U15938 (N_15938,N_6640,N_9342);
nand U15939 (N_15939,N_8630,N_8004);
or U15940 (N_15940,N_8923,N_10119);
or U15941 (N_15941,N_6705,N_11953);
and U15942 (N_15942,N_12068,N_10211);
xnor U15943 (N_15943,N_8383,N_6390);
or U15944 (N_15944,N_6804,N_6351);
and U15945 (N_15945,N_8010,N_8203);
and U15946 (N_15946,N_12325,N_8702);
or U15947 (N_15947,N_11116,N_8143);
nand U15948 (N_15948,N_7411,N_8738);
or U15949 (N_15949,N_10145,N_8721);
and U15950 (N_15950,N_6634,N_11469);
and U15951 (N_15951,N_11123,N_8449);
nor U15952 (N_15952,N_8136,N_11967);
nor U15953 (N_15953,N_8589,N_10877);
or U15954 (N_15954,N_11621,N_7917);
or U15955 (N_15955,N_10779,N_9320);
nor U15956 (N_15956,N_11060,N_9913);
nor U15957 (N_15957,N_9942,N_12060);
nand U15958 (N_15958,N_9962,N_8781);
and U15959 (N_15959,N_7573,N_11810);
or U15960 (N_15960,N_7122,N_7934);
and U15961 (N_15961,N_7291,N_7716);
or U15962 (N_15962,N_6258,N_6295);
or U15963 (N_15963,N_12224,N_10271);
nor U15964 (N_15964,N_11835,N_6685);
or U15965 (N_15965,N_7644,N_12169);
nor U15966 (N_15966,N_9253,N_10174);
nand U15967 (N_15967,N_6865,N_7770);
nand U15968 (N_15968,N_7028,N_11306);
and U15969 (N_15969,N_9620,N_10364);
nand U15970 (N_15970,N_11748,N_7164);
and U15971 (N_15971,N_8110,N_7106);
and U15972 (N_15972,N_12254,N_7035);
nand U15973 (N_15973,N_7965,N_10203);
nand U15974 (N_15974,N_8957,N_9388);
xor U15975 (N_15975,N_6541,N_10253);
and U15976 (N_15976,N_10022,N_10460);
nor U15977 (N_15977,N_8290,N_7704);
and U15978 (N_15978,N_11653,N_6431);
or U15979 (N_15979,N_11474,N_9578);
and U15980 (N_15980,N_6747,N_10772);
nand U15981 (N_15981,N_9216,N_7436);
nand U15982 (N_15982,N_12345,N_9405);
xor U15983 (N_15983,N_9646,N_7112);
nor U15984 (N_15984,N_6466,N_9277);
or U15985 (N_15985,N_8302,N_11771);
or U15986 (N_15986,N_10978,N_7413);
nor U15987 (N_15987,N_11949,N_7371);
nor U15988 (N_15988,N_9761,N_12253);
nor U15989 (N_15989,N_8922,N_6832);
or U15990 (N_15990,N_8004,N_8755);
and U15991 (N_15991,N_6289,N_8044);
xnor U15992 (N_15992,N_8691,N_8036);
xnor U15993 (N_15993,N_11799,N_10969);
xnor U15994 (N_15994,N_7566,N_11372);
nand U15995 (N_15995,N_10368,N_11801);
nor U15996 (N_15996,N_12420,N_10721);
and U15997 (N_15997,N_9646,N_11641);
nor U15998 (N_15998,N_11869,N_7623);
and U15999 (N_15999,N_10705,N_7407);
and U16000 (N_16000,N_10443,N_10693);
nand U16001 (N_16001,N_11848,N_8835);
and U16002 (N_16002,N_8656,N_6250);
or U16003 (N_16003,N_7071,N_6656);
nor U16004 (N_16004,N_9331,N_8345);
nand U16005 (N_16005,N_6950,N_8594);
or U16006 (N_16006,N_6548,N_9568);
nand U16007 (N_16007,N_9448,N_7349);
nor U16008 (N_16008,N_6364,N_10221);
xor U16009 (N_16009,N_12334,N_8109);
nand U16010 (N_16010,N_8977,N_8964);
nor U16011 (N_16011,N_8271,N_6938);
nand U16012 (N_16012,N_8064,N_11190);
and U16013 (N_16013,N_9494,N_10820);
nor U16014 (N_16014,N_10269,N_11429);
nand U16015 (N_16015,N_10094,N_7007);
nor U16016 (N_16016,N_10160,N_11773);
and U16017 (N_16017,N_8206,N_7958);
nand U16018 (N_16018,N_10725,N_8035);
or U16019 (N_16019,N_8695,N_8968);
and U16020 (N_16020,N_8646,N_8296);
xnor U16021 (N_16021,N_7087,N_8004);
or U16022 (N_16022,N_9364,N_8216);
nor U16023 (N_16023,N_10673,N_12105);
or U16024 (N_16024,N_7383,N_9313);
xor U16025 (N_16025,N_7521,N_9154);
and U16026 (N_16026,N_9810,N_6334);
or U16027 (N_16027,N_7375,N_6888);
nor U16028 (N_16028,N_8813,N_12321);
nand U16029 (N_16029,N_7692,N_9964);
or U16030 (N_16030,N_8897,N_7991);
xor U16031 (N_16031,N_11531,N_8273);
and U16032 (N_16032,N_7257,N_8829);
nor U16033 (N_16033,N_6518,N_9495);
nor U16034 (N_16034,N_8640,N_10837);
nor U16035 (N_16035,N_11134,N_6820);
or U16036 (N_16036,N_6930,N_10970);
or U16037 (N_16037,N_8886,N_8906);
and U16038 (N_16038,N_9169,N_12313);
nor U16039 (N_16039,N_8183,N_10453);
and U16040 (N_16040,N_10034,N_11112);
and U16041 (N_16041,N_10257,N_10717);
or U16042 (N_16042,N_7547,N_10987);
nor U16043 (N_16043,N_9367,N_8101);
or U16044 (N_16044,N_12112,N_11546);
nor U16045 (N_16045,N_7889,N_10783);
nor U16046 (N_16046,N_6930,N_9782);
nand U16047 (N_16047,N_10615,N_8395);
nor U16048 (N_16048,N_12488,N_12342);
nand U16049 (N_16049,N_7573,N_7306);
nor U16050 (N_16050,N_8577,N_11707);
nor U16051 (N_16051,N_8957,N_8498);
xor U16052 (N_16052,N_12425,N_11304);
nor U16053 (N_16053,N_6547,N_9623);
nand U16054 (N_16054,N_8838,N_9543);
or U16055 (N_16055,N_6640,N_10359);
nand U16056 (N_16056,N_6292,N_6346);
nand U16057 (N_16057,N_11444,N_11808);
or U16058 (N_16058,N_10817,N_10812);
nor U16059 (N_16059,N_11925,N_6790);
xnor U16060 (N_16060,N_6598,N_7971);
and U16061 (N_16061,N_10078,N_8388);
and U16062 (N_16062,N_11514,N_9288);
nand U16063 (N_16063,N_9184,N_10691);
nor U16064 (N_16064,N_11237,N_8790);
nor U16065 (N_16065,N_9091,N_7936);
nor U16066 (N_16066,N_11652,N_11545);
and U16067 (N_16067,N_10087,N_11949);
nor U16068 (N_16068,N_11229,N_12336);
xnor U16069 (N_16069,N_7510,N_7149);
or U16070 (N_16070,N_12171,N_9890);
nor U16071 (N_16071,N_10699,N_6999);
nor U16072 (N_16072,N_10329,N_10726);
or U16073 (N_16073,N_7643,N_6854);
and U16074 (N_16074,N_11558,N_12325);
or U16075 (N_16075,N_8444,N_10148);
xnor U16076 (N_16076,N_9856,N_8022);
nand U16077 (N_16077,N_8634,N_7744);
nand U16078 (N_16078,N_7648,N_8949);
nor U16079 (N_16079,N_8494,N_7091);
nand U16080 (N_16080,N_8226,N_7279);
and U16081 (N_16081,N_11678,N_11889);
and U16082 (N_16082,N_12478,N_7505);
xor U16083 (N_16083,N_10819,N_11520);
or U16084 (N_16084,N_12049,N_9748);
or U16085 (N_16085,N_6583,N_7523);
xnor U16086 (N_16086,N_10614,N_6410);
or U16087 (N_16087,N_7080,N_6878);
and U16088 (N_16088,N_6436,N_7819);
or U16089 (N_16089,N_8398,N_8147);
nand U16090 (N_16090,N_8948,N_7050);
and U16091 (N_16091,N_9079,N_9366);
and U16092 (N_16092,N_11969,N_9873);
nor U16093 (N_16093,N_10284,N_10127);
nand U16094 (N_16094,N_11423,N_7813);
or U16095 (N_16095,N_10625,N_7027);
nor U16096 (N_16096,N_7136,N_11153);
nor U16097 (N_16097,N_8275,N_11034);
nand U16098 (N_16098,N_11564,N_10462);
and U16099 (N_16099,N_12182,N_7868);
xnor U16100 (N_16100,N_6397,N_11352);
or U16101 (N_16101,N_7684,N_8697);
nand U16102 (N_16102,N_8546,N_7359);
nand U16103 (N_16103,N_11891,N_7366);
nor U16104 (N_16104,N_9525,N_7372);
nand U16105 (N_16105,N_9979,N_12472);
nor U16106 (N_16106,N_11257,N_10487);
nand U16107 (N_16107,N_11739,N_11552);
nor U16108 (N_16108,N_10900,N_8557);
nand U16109 (N_16109,N_9196,N_10415);
or U16110 (N_16110,N_7699,N_9980);
xnor U16111 (N_16111,N_12265,N_8440);
and U16112 (N_16112,N_9098,N_11602);
nand U16113 (N_16113,N_8046,N_8086);
nor U16114 (N_16114,N_11697,N_7010);
and U16115 (N_16115,N_7771,N_12236);
nor U16116 (N_16116,N_12298,N_12223);
nand U16117 (N_16117,N_9777,N_10111);
or U16118 (N_16118,N_10039,N_8067);
xnor U16119 (N_16119,N_9544,N_7160);
nand U16120 (N_16120,N_8704,N_12055);
and U16121 (N_16121,N_8546,N_8589);
nand U16122 (N_16122,N_12030,N_10302);
or U16123 (N_16123,N_7247,N_9828);
xnor U16124 (N_16124,N_6745,N_7984);
and U16125 (N_16125,N_12479,N_8675);
nand U16126 (N_16126,N_12231,N_11599);
nand U16127 (N_16127,N_11693,N_8756);
nand U16128 (N_16128,N_6724,N_8422);
nand U16129 (N_16129,N_10319,N_10556);
and U16130 (N_16130,N_9103,N_9843);
or U16131 (N_16131,N_10645,N_10585);
nand U16132 (N_16132,N_9344,N_6485);
or U16133 (N_16133,N_9896,N_8595);
or U16134 (N_16134,N_10784,N_6767);
nand U16135 (N_16135,N_6612,N_12032);
or U16136 (N_16136,N_6893,N_9407);
or U16137 (N_16137,N_11949,N_10190);
and U16138 (N_16138,N_11808,N_6523);
and U16139 (N_16139,N_10180,N_12210);
nor U16140 (N_16140,N_11310,N_10174);
or U16141 (N_16141,N_7036,N_12097);
nor U16142 (N_16142,N_7141,N_9535);
nor U16143 (N_16143,N_6809,N_8304);
or U16144 (N_16144,N_11554,N_6747);
or U16145 (N_16145,N_7976,N_9379);
and U16146 (N_16146,N_11747,N_7617);
xor U16147 (N_16147,N_6535,N_7858);
nor U16148 (N_16148,N_7280,N_8225);
nor U16149 (N_16149,N_11151,N_9026);
xor U16150 (N_16150,N_7325,N_6438);
nand U16151 (N_16151,N_9139,N_7128);
nand U16152 (N_16152,N_7729,N_11731);
and U16153 (N_16153,N_7812,N_7764);
nor U16154 (N_16154,N_11396,N_12495);
xnor U16155 (N_16155,N_8708,N_10567);
nand U16156 (N_16156,N_8422,N_10860);
nor U16157 (N_16157,N_10054,N_9777);
nor U16158 (N_16158,N_6442,N_9227);
nor U16159 (N_16159,N_11780,N_10734);
or U16160 (N_16160,N_9758,N_8384);
and U16161 (N_16161,N_6833,N_12017);
nor U16162 (N_16162,N_6303,N_7647);
and U16163 (N_16163,N_10709,N_8837);
nor U16164 (N_16164,N_9660,N_8118);
nand U16165 (N_16165,N_10241,N_10540);
and U16166 (N_16166,N_7981,N_11228);
or U16167 (N_16167,N_6763,N_6992);
and U16168 (N_16168,N_7000,N_11707);
nor U16169 (N_16169,N_8095,N_11449);
and U16170 (N_16170,N_6936,N_8745);
xnor U16171 (N_16171,N_7062,N_6285);
and U16172 (N_16172,N_11960,N_10629);
nor U16173 (N_16173,N_11735,N_8694);
and U16174 (N_16174,N_6896,N_10621);
and U16175 (N_16175,N_9702,N_11406);
and U16176 (N_16176,N_6634,N_6271);
nor U16177 (N_16177,N_6579,N_7912);
and U16178 (N_16178,N_11098,N_8898);
and U16179 (N_16179,N_10895,N_6581);
nand U16180 (N_16180,N_9616,N_9258);
nand U16181 (N_16181,N_6378,N_7727);
and U16182 (N_16182,N_11967,N_8244);
and U16183 (N_16183,N_9343,N_7424);
nand U16184 (N_16184,N_6670,N_8901);
nor U16185 (N_16185,N_8412,N_7631);
and U16186 (N_16186,N_6571,N_11985);
nand U16187 (N_16187,N_7911,N_8376);
and U16188 (N_16188,N_9531,N_10907);
or U16189 (N_16189,N_12107,N_11429);
and U16190 (N_16190,N_10568,N_12012);
nand U16191 (N_16191,N_11423,N_8897);
nand U16192 (N_16192,N_8204,N_10177);
or U16193 (N_16193,N_6723,N_8276);
and U16194 (N_16194,N_7768,N_8602);
nand U16195 (N_16195,N_12321,N_11404);
xor U16196 (N_16196,N_12410,N_8673);
nor U16197 (N_16197,N_6583,N_9873);
or U16198 (N_16198,N_6285,N_10363);
and U16199 (N_16199,N_7736,N_8492);
or U16200 (N_16200,N_12131,N_6445);
and U16201 (N_16201,N_7314,N_8000);
nand U16202 (N_16202,N_6334,N_7041);
and U16203 (N_16203,N_9629,N_11866);
or U16204 (N_16204,N_8230,N_11964);
or U16205 (N_16205,N_10139,N_7190);
nand U16206 (N_16206,N_11715,N_12291);
nand U16207 (N_16207,N_10328,N_10790);
nand U16208 (N_16208,N_6662,N_9380);
and U16209 (N_16209,N_8711,N_10179);
xor U16210 (N_16210,N_12378,N_11415);
nand U16211 (N_16211,N_9033,N_12313);
nand U16212 (N_16212,N_9136,N_10362);
and U16213 (N_16213,N_10235,N_8882);
nand U16214 (N_16214,N_12301,N_10754);
or U16215 (N_16215,N_8448,N_11353);
nor U16216 (N_16216,N_6435,N_12053);
or U16217 (N_16217,N_6595,N_9749);
or U16218 (N_16218,N_11507,N_7482);
nand U16219 (N_16219,N_11624,N_10596);
nand U16220 (N_16220,N_10251,N_11369);
nand U16221 (N_16221,N_7273,N_11412);
and U16222 (N_16222,N_11735,N_9474);
xnor U16223 (N_16223,N_7033,N_12431);
and U16224 (N_16224,N_12044,N_10318);
or U16225 (N_16225,N_10785,N_11138);
or U16226 (N_16226,N_9201,N_7764);
or U16227 (N_16227,N_10333,N_11172);
and U16228 (N_16228,N_6278,N_6752);
nand U16229 (N_16229,N_11291,N_12409);
and U16230 (N_16230,N_12038,N_11191);
or U16231 (N_16231,N_9478,N_10438);
xnor U16232 (N_16232,N_6327,N_8223);
nor U16233 (N_16233,N_8859,N_8655);
and U16234 (N_16234,N_12268,N_9643);
nor U16235 (N_16235,N_9799,N_10107);
nand U16236 (N_16236,N_9490,N_11329);
nand U16237 (N_16237,N_12241,N_7758);
nand U16238 (N_16238,N_11846,N_6352);
nand U16239 (N_16239,N_11430,N_11483);
nor U16240 (N_16240,N_12180,N_6738);
xor U16241 (N_16241,N_8340,N_8370);
or U16242 (N_16242,N_8052,N_10502);
and U16243 (N_16243,N_10024,N_8673);
nor U16244 (N_16244,N_8167,N_8057);
xnor U16245 (N_16245,N_6713,N_10987);
nor U16246 (N_16246,N_9270,N_10325);
xnor U16247 (N_16247,N_9023,N_12198);
nor U16248 (N_16248,N_7057,N_8191);
nand U16249 (N_16249,N_8052,N_8950);
and U16250 (N_16250,N_8950,N_9332);
and U16251 (N_16251,N_11869,N_11185);
nor U16252 (N_16252,N_8389,N_12135);
nand U16253 (N_16253,N_7676,N_8950);
and U16254 (N_16254,N_8435,N_8844);
or U16255 (N_16255,N_11279,N_7572);
or U16256 (N_16256,N_7949,N_6907);
nor U16257 (N_16257,N_12074,N_11323);
nand U16258 (N_16258,N_8521,N_10767);
nand U16259 (N_16259,N_11339,N_9006);
xnor U16260 (N_16260,N_9576,N_7406);
nand U16261 (N_16261,N_8109,N_8053);
and U16262 (N_16262,N_6772,N_11524);
or U16263 (N_16263,N_9678,N_12344);
nand U16264 (N_16264,N_8562,N_12043);
nand U16265 (N_16265,N_10977,N_11398);
xor U16266 (N_16266,N_8907,N_8352);
nand U16267 (N_16267,N_8771,N_7610);
nor U16268 (N_16268,N_7580,N_6880);
nor U16269 (N_16269,N_11776,N_10362);
nand U16270 (N_16270,N_7539,N_10910);
and U16271 (N_16271,N_9455,N_11815);
and U16272 (N_16272,N_8762,N_12430);
nand U16273 (N_16273,N_7636,N_12425);
or U16274 (N_16274,N_10700,N_8557);
nand U16275 (N_16275,N_6362,N_6629);
xor U16276 (N_16276,N_6369,N_8754);
nor U16277 (N_16277,N_10633,N_12024);
or U16278 (N_16278,N_12428,N_11945);
nor U16279 (N_16279,N_9321,N_7224);
nor U16280 (N_16280,N_7563,N_8922);
and U16281 (N_16281,N_6765,N_11690);
nor U16282 (N_16282,N_11771,N_6844);
nor U16283 (N_16283,N_6570,N_6310);
xor U16284 (N_16284,N_7184,N_7206);
and U16285 (N_16285,N_12373,N_7821);
nand U16286 (N_16286,N_12235,N_12362);
and U16287 (N_16287,N_10754,N_10336);
xor U16288 (N_16288,N_9871,N_9683);
or U16289 (N_16289,N_8914,N_11936);
nor U16290 (N_16290,N_11120,N_11814);
nor U16291 (N_16291,N_10465,N_11246);
nor U16292 (N_16292,N_10619,N_10426);
nor U16293 (N_16293,N_6734,N_10880);
nor U16294 (N_16294,N_8369,N_7079);
or U16295 (N_16295,N_9375,N_11357);
nand U16296 (N_16296,N_6317,N_10393);
nand U16297 (N_16297,N_6902,N_11297);
nand U16298 (N_16298,N_12063,N_11317);
and U16299 (N_16299,N_12097,N_11113);
and U16300 (N_16300,N_7472,N_9470);
nor U16301 (N_16301,N_10340,N_8374);
nand U16302 (N_16302,N_6887,N_9883);
nand U16303 (N_16303,N_12038,N_12213);
or U16304 (N_16304,N_11049,N_11591);
or U16305 (N_16305,N_7837,N_8223);
or U16306 (N_16306,N_11128,N_11958);
xnor U16307 (N_16307,N_11942,N_10565);
and U16308 (N_16308,N_7501,N_9522);
or U16309 (N_16309,N_8737,N_11736);
or U16310 (N_16310,N_11682,N_7499);
xor U16311 (N_16311,N_8778,N_11061);
xor U16312 (N_16312,N_10766,N_11262);
nand U16313 (N_16313,N_11119,N_8253);
and U16314 (N_16314,N_11615,N_12297);
and U16315 (N_16315,N_8227,N_8797);
nor U16316 (N_16316,N_8710,N_11261);
nand U16317 (N_16317,N_8705,N_6429);
or U16318 (N_16318,N_6897,N_11254);
and U16319 (N_16319,N_10391,N_11838);
nand U16320 (N_16320,N_8783,N_11213);
and U16321 (N_16321,N_11596,N_8878);
nor U16322 (N_16322,N_9588,N_11288);
nor U16323 (N_16323,N_8752,N_10292);
or U16324 (N_16324,N_9392,N_11414);
nor U16325 (N_16325,N_8161,N_11198);
nor U16326 (N_16326,N_11454,N_8300);
and U16327 (N_16327,N_8659,N_7744);
nand U16328 (N_16328,N_8790,N_7112);
xnor U16329 (N_16329,N_11306,N_6926);
or U16330 (N_16330,N_12309,N_8455);
nor U16331 (N_16331,N_8544,N_7511);
nor U16332 (N_16332,N_8354,N_8898);
nand U16333 (N_16333,N_7428,N_6834);
xnor U16334 (N_16334,N_12381,N_12389);
and U16335 (N_16335,N_8752,N_7976);
nand U16336 (N_16336,N_8870,N_12383);
nand U16337 (N_16337,N_8779,N_9869);
or U16338 (N_16338,N_6496,N_11974);
nand U16339 (N_16339,N_8665,N_12004);
and U16340 (N_16340,N_10862,N_9310);
nor U16341 (N_16341,N_8772,N_10219);
and U16342 (N_16342,N_8063,N_10833);
nand U16343 (N_16343,N_6473,N_10111);
or U16344 (N_16344,N_8184,N_11505);
or U16345 (N_16345,N_7207,N_8165);
and U16346 (N_16346,N_6450,N_6791);
nand U16347 (N_16347,N_12226,N_11801);
nor U16348 (N_16348,N_11496,N_6701);
or U16349 (N_16349,N_10491,N_8301);
and U16350 (N_16350,N_11661,N_9436);
or U16351 (N_16351,N_10051,N_10275);
nor U16352 (N_16352,N_9366,N_7311);
and U16353 (N_16353,N_12407,N_9690);
or U16354 (N_16354,N_10311,N_10526);
nand U16355 (N_16355,N_7712,N_8515);
nand U16356 (N_16356,N_8503,N_11820);
nand U16357 (N_16357,N_9344,N_11107);
and U16358 (N_16358,N_9474,N_9466);
and U16359 (N_16359,N_11350,N_9825);
and U16360 (N_16360,N_9163,N_9018);
or U16361 (N_16361,N_8617,N_8801);
nor U16362 (N_16362,N_7558,N_12194);
and U16363 (N_16363,N_7744,N_9398);
nor U16364 (N_16364,N_6749,N_12495);
nor U16365 (N_16365,N_7998,N_11231);
or U16366 (N_16366,N_9810,N_12324);
and U16367 (N_16367,N_9429,N_6794);
nand U16368 (N_16368,N_7488,N_10565);
nand U16369 (N_16369,N_6814,N_10242);
and U16370 (N_16370,N_9386,N_6476);
and U16371 (N_16371,N_12374,N_9738);
nor U16372 (N_16372,N_9287,N_7928);
nand U16373 (N_16373,N_7753,N_10398);
or U16374 (N_16374,N_9290,N_9162);
xnor U16375 (N_16375,N_12282,N_8839);
nor U16376 (N_16376,N_9803,N_10725);
nand U16377 (N_16377,N_11806,N_10027);
xor U16378 (N_16378,N_11080,N_10181);
nand U16379 (N_16379,N_8179,N_11253);
nor U16380 (N_16380,N_7855,N_6605);
or U16381 (N_16381,N_10736,N_11537);
or U16382 (N_16382,N_10015,N_7155);
nor U16383 (N_16383,N_11990,N_9901);
and U16384 (N_16384,N_8477,N_12360);
or U16385 (N_16385,N_11791,N_9648);
nor U16386 (N_16386,N_10815,N_10508);
nand U16387 (N_16387,N_9199,N_8067);
nor U16388 (N_16388,N_8970,N_9809);
or U16389 (N_16389,N_9295,N_7879);
nand U16390 (N_16390,N_11057,N_7208);
nand U16391 (N_16391,N_6272,N_10121);
xor U16392 (N_16392,N_7072,N_11636);
xnor U16393 (N_16393,N_7430,N_11988);
xor U16394 (N_16394,N_6953,N_8570);
and U16395 (N_16395,N_8753,N_8491);
nor U16396 (N_16396,N_12402,N_10581);
nor U16397 (N_16397,N_10827,N_9680);
or U16398 (N_16398,N_7356,N_7733);
nor U16399 (N_16399,N_11589,N_9270);
nand U16400 (N_16400,N_10672,N_7549);
and U16401 (N_16401,N_12422,N_9131);
xor U16402 (N_16402,N_11072,N_8423);
nand U16403 (N_16403,N_12365,N_9113);
and U16404 (N_16404,N_11478,N_10066);
nand U16405 (N_16405,N_6467,N_11703);
nand U16406 (N_16406,N_7644,N_11253);
nand U16407 (N_16407,N_11486,N_8451);
nand U16408 (N_16408,N_6802,N_9397);
or U16409 (N_16409,N_9275,N_12307);
nor U16410 (N_16410,N_11676,N_8632);
or U16411 (N_16411,N_9583,N_9238);
nor U16412 (N_16412,N_11273,N_6991);
or U16413 (N_16413,N_7425,N_12324);
or U16414 (N_16414,N_11897,N_11654);
or U16415 (N_16415,N_9557,N_11592);
nand U16416 (N_16416,N_8531,N_10990);
or U16417 (N_16417,N_8641,N_11966);
nand U16418 (N_16418,N_6866,N_7508);
nand U16419 (N_16419,N_9892,N_9990);
and U16420 (N_16420,N_6661,N_9469);
nor U16421 (N_16421,N_10939,N_7397);
and U16422 (N_16422,N_6572,N_11840);
or U16423 (N_16423,N_9105,N_10491);
nor U16424 (N_16424,N_8180,N_8229);
xnor U16425 (N_16425,N_10684,N_6585);
nand U16426 (N_16426,N_9695,N_7199);
nand U16427 (N_16427,N_6311,N_7787);
and U16428 (N_16428,N_9718,N_12396);
nand U16429 (N_16429,N_11728,N_12331);
nand U16430 (N_16430,N_8837,N_10830);
or U16431 (N_16431,N_10906,N_9221);
nor U16432 (N_16432,N_7755,N_8112);
nor U16433 (N_16433,N_8535,N_12012);
nand U16434 (N_16434,N_9947,N_11646);
nand U16435 (N_16435,N_6835,N_9791);
and U16436 (N_16436,N_7588,N_6590);
and U16437 (N_16437,N_6564,N_9104);
or U16438 (N_16438,N_11868,N_12012);
and U16439 (N_16439,N_8610,N_6674);
and U16440 (N_16440,N_12117,N_11003);
or U16441 (N_16441,N_11767,N_8368);
nor U16442 (N_16442,N_7862,N_12449);
or U16443 (N_16443,N_7235,N_10058);
or U16444 (N_16444,N_8719,N_7654);
nand U16445 (N_16445,N_8227,N_8964);
nand U16446 (N_16446,N_11715,N_10565);
nand U16447 (N_16447,N_6296,N_11382);
nor U16448 (N_16448,N_12319,N_12033);
and U16449 (N_16449,N_7816,N_7558);
nor U16450 (N_16450,N_11808,N_9531);
or U16451 (N_16451,N_7696,N_8589);
nand U16452 (N_16452,N_10935,N_9213);
or U16453 (N_16453,N_11749,N_8549);
nor U16454 (N_16454,N_10546,N_6620);
nor U16455 (N_16455,N_10308,N_11999);
nor U16456 (N_16456,N_8560,N_8881);
nor U16457 (N_16457,N_11133,N_11316);
nor U16458 (N_16458,N_10040,N_7000);
xnor U16459 (N_16459,N_8849,N_6467);
nor U16460 (N_16460,N_8114,N_7998);
nand U16461 (N_16461,N_8881,N_8773);
nand U16462 (N_16462,N_11772,N_7773);
nand U16463 (N_16463,N_7509,N_7350);
nor U16464 (N_16464,N_10555,N_10098);
nand U16465 (N_16465,N_9125,N_12351);
nand U16466 (N_16466,N_12470,N_10549);
or U16467 (N_16467,N_10638,N_11294);
xnor U16468 (N_16468,N_8777,N_6622);
nor U16469 (N_16469,N_7626,N_7577);
nor U16470 (N_16470,N_10022,N_6385);
nor U16471 (N_16471,N_8381,N_11874);
nand U16472 (N_16472,N_11862,N_8946);
nand U16473 (N_16473,N_10682,N_10016);
nor U16474 (N_16474,N_10244,N_11165);
nor U16475 (N_16475,N_11441,N_11736);
and U16476 (N_16476,N_6580,N_10207);
or U16477 (N_16477,N_8583,N_10015);
or U16478 (N_16478,N_8409,N_9360);
nand U16479 (N_16479,N_8290,N_6319);
or U16480 (N_16480,N_8364,N_11513);
and U16481 (N_16481,N_10895,N_10047);
nor U16482 (N_16482,N_11152,N_12121);
and U16483 (N_16483,N_9003,N_11112);
and U16484 (N_16484,N_11738,N_9254);
nand U16485 (N_16485,N_10322,N_7663);
nand U16486 (N_16486,N_9655,N_8504);
nand U16487 (N_16487,N_9603,N_10277);
nand U16488 (N_16488,N_8154,N_10822);
or U16489 (N_16489,N_7759,N_9110);
nor U16490 (N_16490,N_9892,N_8637);
xor U16491 (N_16491,N_12179,N_6906);
nand U16492 (N_16492,N_7715,N_7099);
or U16493 (N_16493,N_10714,N_10040);
and U16494 (N_16494,N_10949,N_10208);
or U16495 (N_16495,N_10102,N_11585);
and U16496 (N_16496,N_6976,N_11392);
or U16497 (N_16497,N_7457,N_8344);
xnor U16498 (N_16498,N_10485,N_12012);
and U16499 (N_16499,N_11743,N_7120);
and U16500 (N_16500,N_7680,N_8329);
nand U16501 (N_16501,N_7822,N_9922);
or U16502 (N_16502,N_8960,N_8961);
and U16503 (N_16503,N_12322,N_7302);
or U16504 (N_16504,N_10934,N_7359);
xnor U16505 (N_16505,N_8144,N_9241);
nor U16506 (N_16506,N_12434,N_10623);
and U16507 (N_16507,N_7966,N_10706);
nor U16508 (N_16508,N_8120,N_7978);
nand U16509 (N_16509,N_8006,N_9881);
nor U16510 (N_16510,N_11430,N_9908);
and U16511 (N_16511,N_11348,N_11680);
nor U16512 (N_16512,N_11923,N_11059);
and U16513 (N_16513,N_6770,N_7450);
nor U16514 (N_16514,N_8267,N_11283);
nor U16515 (N_16515,N_6352,N_12069);
or U16516 (N_16516,N_9618,N_9303);
xnor U16517 (N_16517,N_10939,N_11995);
and U16518 (N_16518,N_11819,N_9827);
nor U16519 (N_16519,N_8387,N_9061);
xor U16520 (N_16520,N_9300,N_7035);
nand U16521 (N_16521,N_7831,N_12390);
nand U16522 (N_16522,N_10731,N_9790);
and U16523 (N_16523,N_7404,N_10547);
nor U16524 (N_16524,N_7221,N_6633);
nand U16525 (N_16525,N_7987,N_8920);
nor U16526 (N_16526,N_10877,N_9132);
nand U16527 (N_16527,N_6729,N_6786);
xnor U16528 (N_16528,N_11785,N_8696);
xnor U16529 (N_16529,N_7172,N_6668);
nand U16530 (N_16530,N_10507,N_11970);
xor U16531 (N_16531,N_7708,N_8394);
nand U16532 (N_16532,N_11685,N_8563);
and U16533 (N_16533,N_6659,N_12131);
or U16534 (N_16534,N_11279,N_6615);
nand U16535 (N_16535,N_7568,N_8726);
and U16536 (N_16536,N_10612,N_8818);
nor U16537 (N_16537,N_11084,N_7201);
or U16538 (N_16538,N_10744,N_8130);
xnor U16539 (N_16539,N_8622,N_11688);
nor U16540 (N_16540,N_8206,N_8002);
or U16541 (N_16541,N_10847,N_6882);
or U16542 (N_16542,N_8540,N_11212);
and U16543 (N_16543,N_11886,N_10246);
and U16544 (N_16544,N_10153,N_11806);
and U16545 (N_16545,N_6390,N_11690);
and U16546 (N_16546,N_8521,N_7247);
or U16547 (N_16547,N_11560,N_12414);
nor U16548 (N_16548,N_9299,N_11851);
nand U16549 (N_16549,N_8724,N_11478);
nand U16550 (N_16550,N_11776,N_6919);
nor U16551 (N_16551,N_6751,N_7257);
nand U16552 (N_16552,N_6953,N_7361);
nand U16553 (N_16553,N_6584,N_9579);
nor U16554 (N_16554,N_10381,N_6811);
nand U16555 (N_16555,N_6527,N_6808);
xor U16556 (N_16556,N_12217,N_9308);
or U16557 (N_16557,N_11658,N_7646);
or U16558 (N_16558,N_12244,N_9446);
and U16559 (N_16559,N_8831,N_10443);
or U16560 (N_16560,N_9228,N_8380);
nand U16561 (N_16561,N_9039,N_9508);
nand U16562 (N_16562,N_8587,N_7527);
xnor U16563 (N_16563,N_10492,N_11290);
nand U16564 (N_16564,N_8244,N_9958);
and U16565 (N_16565,N_6726,N_11800);
and U16566 (N_16566,N_11254,N_10059);
nand U16567 (N_16567,N_6914,N_8326);
xor U16568 (N_16568,N_7936,N_11865);
nor U16569 (N_16569,N_10837,N_10121);
nor U16570 (N_16570,N_12225,N_10819);
xor U16571 (N_16571,N_12026,N_7142);
nor U16572 (N_16572,N_6699,N_6827);
and U16573 (N_16573,N_7273,N_8482);
nand U16574 (N_16574,N_9876,N_6973);
nand U16575 (N_16575,N_11553,N_7961);
or U16576 (N_16576,N_10442,N_6672);
nand U16577 (N_16577,N_8193,N_8313);
nor U16578 (N_16578,N_12197,N_6767);
xnor U16579 (N_16579,N_11017,N_6681);
nand U16580 (N_16580,N_7854,N_10677);
or U16581 (N_16581,N_6253,N_8881);
xnor U16582 (N_16582,N_7223,N_6407);
and U16583 (N_16583,N_8961,N_11814);
nand U16584 (N_16584,N_9822,N_6513);
nand U16585 (N_16585,N_9636,N_12474);
or U16586 (N_16586,N_7432,N_9833);
nor U16587 (N_16587,N_11729,N_9960);
nor U16588 (N_16588,N_7353,N_8257);
nor U16589 (N_16589,N_6515,N_10864);
nor U16590 (N_16590,N_9897,N_10549);
nand U16591 (N_16591,N_11172,N_7324);
nand U16592 (N_16592,N_9937,N_10425);
xor U16593 (N_16593,N_6491,N_10787);
nand U16594 (N_16594,N_8868,N_8705);
and U16595 (N_16595,N_6441,N_10546);
nor U16596 (N_16596,N_10510,N_7561);
nand U16597 (N_16597,N_9855,N_11376);
or U16598 (N_16598,N_10205,N_10194);
xnor U16599 (N_16599,N_10525,N_6957);
or U16600 (N_16600,N_8465,N_9629);
and U16601 (N_16601,N_8816,N_11934);
nand U16602 (N_16602,N_11390,N_11176);
xor U16603 (N_16603,N_7408,N_6430);
nor U16604 (N_16604,N_7004,N_6781);
nand U16605 (N_16605,N_6283,N_7669);
or U16606 (N_16606,N_12486,N_8978);
nand U16607 (N_16607,N_11707,N_9994);
nand U16608 (N_16608,N_7250,N_6675);
nor U16609 (N_16609,N_9069,N_8334);
nor U16610 (N_16610,N_11024,N_9368);
nor U16611 (N_16611,N_6293,N_6967);
nor U16612 (N_16612,N_9065,N_11743);
and U16613 (N_16613,N_9775,N_9355);
or U16614 (N_16614,N_7488,N_9732);
nand U16615 (N_16615,N_11984,N_6485);
and U16616 (N_16616,N_8965,N_6964);
or U16617 (N_16617,N_7805,N_6396);
nor U16618 (N_16618,N_10585,N_7092);
or U16619 (N_16619,N_10199,N_6559);
or U16620 (N_16620,N_7332,N_8594);
nor U16621 (N_16621,N_9665,N_12149);
and U16622 (N_16622,N_6829,N_9546);
or U16623 (N_16623,N_11922,N_10178);
and U16624 (N_16624,N_11233,N_11459);
nor U16625 (N_16625,N_8173,N_6875);
nor U16626 (N_16626,N_12401,N_6745);
nor U16627 (N_16627,N_10837,N_7509);
or U16628 (N_16628,N_11099,N_12361);
and U16629 (N_16629,N_8276,N_10684);
nand U16630 (N_16630,N_7199,N_12358);
or U16631 (N_16631,N_8981,N_10334);
nand U16632 (N_16632,N_11309,N_8543);
nor U16633 (N_16633,N_7186,N_8637);
nor U16634 (N_16634,N_11928,N_6333);
nor U16635 (N_16635,N_7976,N_11118);
xor U16636 (N_16636,N_11254,N_9190);
nor U16637 (N_16637,N_8640,N_8350);
nor U16638 (N_16638,N_12238,N_8444);
nor U16639 (N_16639,N_9125,N_8086);
or U16640 (N_16640,N_6967,N_11802);
and U16641 (N_16641,N_7333,N_11278);
nor U16642 (N_16642,N_11123,N_6815);
and U16643 (N_16643,N_8339,N_11831);
nor U16644 (N_16644,N_11753,N_9548);
nand U16645 (N_16645,N_9169,N_6956);
nor U16646 (N_16646,N_6741,N_8290);
nand U16647 (N_16647,N_7124,N_11464);
nor U16648 (N_16648,N_7854,N_7961);
nor U16649 (N_16649,N_10161,N_10266);
and U16650 (N_16650,N_10040,N_12051);
or U16651 (N_16651,N_10497,N_11648);
xnor U16652 (N_16652,N_8667,N_12342);
nor U16653 (N_16653,N_10842,N_11902);
or U16654 (N_16654,N_7016,N_11991);
nand U16655 (N_16655,N_8201,N_6849);
or U16656 (N_16656,N_8175,N_8630);
nor U16657 (N_16657,N_7445,N_10022);
nor U16658 (N_16658,N_6567,N_10499);
nor U16659 (N_16659,N_7660,N_12126);
nand U16660 (N_16660,N_6808,N_12325);
nor U16661 (N_16661,N_9247,N_9417);
nand U16662 (N_16662,N_6671,N_11160);
nor U16663 (N_16663,N_11191,N_10595);
nand U16664 (N_16664,N_6779,N_7574);
nand U16665 (N_16665,N_8754,N_11556);
or U16666 (N_16666,N_8022,N_9204);
nand U16667 (N_16667,N_9044,N_7215);
or U16668 (N_16668,N_11641,N_6781);
and U16669 (N_16669,N_9407,N_11873);
nand U16670 (N_16670,N_7703,N_10311);
nand U16671 (N_16671,N_8330,N_9708);
nor U16672 (N_16672,N_7106,N_9958);
nor U16673 (N_16673,N_8537,N_9422);
nor U16674 (N_16674,N_7406,N_9060);
and U16675 (N_16675,N_9847,N_11436);
nor U16676 (N_16676,N_7206,N_9898);
or U16677 (N_16677,N_8212,N_10087);
or U16678 (N_16678,N_10714,N_7191);
or U16679 (N_16679,N_7503,N_8205);
and U16680 (N_16680,N_9645,N_8178);
nand U16681 (N_16681,N_8632,N_11704);
nand U16682 (N_16682,N_7014,N_10103);
or U16683 (N_16683,N_12155,N_7398);
nand U16684 (N_16684,N_11436,N_9468);
or U16685 (N_16685,N_8978,N_11689);
nor U16686 (N_16686,N_6747,N_6539);
nand U16687 (N_16687,N_6274,N_6636);
nor U16688 (N_16688,N_11475,N_8674);
nand U16689 (N_16689,N_12037,N_11416);
nor U16690 (N_16690,N_10443,N_11275);
and U16691 (N_16691,N_8418,N_11037);
or U16692 (N_16692,N_8936,N_12327);
nand U16693 (N_16693,N_10159,N_9157);
nand U16694 (N_16694,N_10091,N_6549);
or U16695 (N_16695,N_6346,N_9309);
or U16696 (N_16696,N_11952,N_6750);
nor U16697 (N_16697,N_7154,N_12403);
nand U16698 (N_16698,N_10712,N_7461);
or U16699 (N_16699,N_11712,N_6325);
nor U16700 (N_16700,N_6566,N_9164);
nor U16701 (N_16701,N_10979,N_6522);
or U16702 (N_16702,N_8070,N_7338);
and U16703 (N_16703,N_10569,N_10504);
nand U16704 (N_16704,N_8830,N_9195);
and U16705 (N_16705,N_7853,N_10543);
nor U16706 (N_16706,N_12442,N_10414);
nor U16707 (N_16707,N_9371,N_11796);
or U16708 (N_16708,N_10378,N_10418);
nor U16709 (N_16709,N_7444,N_6509);
and U16710 (N_16710,N_7190,N_11614);
nand U16711 (N_16711,N_9891,N_6864);
nor U16712 (N_16712,N_11512,N_7512);
nor U16713 (N_16713,N_7765,N_11094);
or U16714 (N_16714,N_7454,N_8220);
xor U16715 (N_16715,N_12000,N_10076);
nor U16716 (N_16716,N_10565,N_11257);
xor U16717 (N_16717,N_10572,N_10950);
or U16718 (N_16718,N_6750,N_8323);
or U16719 (N_16719,N_6252,N_11220);
nand U16720 (N_16720,N_7161,N_8372);
nor U16721 (N_16721,N_10003,N_10584);
nor U16722 (N_16722,N_10725,N_9974);
and U16723 (N_16723,N_10061,N_12361);
or U16724 (N_16724,N_9423,N_6455);
or U16725 (N_16725,N_9421,N_10417);
nand U16726 (N_16726,N_8354,N_7763);
nand U16727 (N_16727,N_6907,N_8614);
nor U16728 (N_16728,N_8601,N_9836);
xnor U16729 (N_16729,N_10590,N_12318);
and U16730 (N_16730,N_10954,N_7456);
nor U16731 (N_16731,N_12241,N_9501);
and U16732 (N_16732,N_8456,N_9855);
and U16733 (N_16733,N_6846,N_7768);
or U16734 (N_16734,N_8690,N_10368);
or U16735 (N_16735,N_11274,N_11128);
or U16736 (N_16736,N_7649,N_10210);
nor U16737 (N_16737,N_8413,N_10558);
and U16738 (N_16738,N_11438,N_6861);
and U16739 (N_16739,N_11666,N_9509);
nor U16740 (N_16740,N_11545,N_6603);
nand U16741 (N_16741,N_6369,N_12461);
and U16742 (N_16742,N_6393,N_11006);
nand U16743 (N_16743,N_11358,N_8003);
or U16744 (N_16744,N_6754,N_8763);
nand U16745 (N_16745,N_10298,N_12135);
xnor U16746 (N_16746,N_6269,N_6965);
nand U16747 (N_16747,N_7387,N_7564);
and U16748 (N_16748,N_12015,N_10961);
nand U16749 (N_16749,N_11876,N_9861);
and U16750 (N_16750,N_7495,N_7555);
nor U16751 (N_16751,N_10911,N_8414);
or U16752 (N_16752,N_12172,N_8799);
nor U16753 (N_16753,N_8282,N_10568);
nor U16754 (N_16754,N_12188,N_7649);
nor U16755 (N_16755,N_10737,N_11256);
or U16756 (N_16756,N_9324,N_11745);
nor U16757 (N_16757,N_10353,N_9752);
xnor U16758 (N_16758,N_11877,N_10277);
and U16759 (N_16759,N_9172,N_11242);
and U16760 (N_16760,N_7032,N_6715);
or U16761 (N_16761,N_9740,N_9374);
nand U16762 (N_16762,N_11566,N_7923);
or U16763 (N_16763,N_8587,N_10977);
or U16764 (N_16764,N_9975,N_10916);
and U16765 (N_16765,N_11775,N_8391);
or U16766 (N_16766,N_8423,N_12283);
or U16767 (N_16767,N_10305,N_8932);
nand U16768 (N_16768,N_11968,N_10636);
or U16769 (N_16769,N_10691,N_9646);
nor U16770 (N_16770,N_9056,N_9851);
and U16771 (N_16771,N_11830,N_6271);
or U16772 (N_16772,N_11239,N_12431);
and U16773 (N_16773,N_12023,N_8908);
and U16774 (N_16774,N_7638,N_12413);
nand U16775 (N_16775,N_7587,N_8233);
nand U16776 (N_16776,N_6759,N_8218);
nor U16777 (N_16777,N_8172,N_7536);
nand U16778 (N_16778,N_7326,N_10202);
and U16779 (N_16779,N_9919,N_8775);
or U16780 (N_16780,N_8954,N_6690);
nor U16781 (N_16781,N_6786,N_10146);
or U16782 (N_16782,N_9288,N_7304);
nor U16783 (N_16783,N_9387,N_8433);
nand U16784 (N_16784,N_9442,N_9836);
or U16785 (N_16785,N_7219,N_8230);
nor U16786 (N_16786,N_6768,N_8046);
or U16787 (N_16787,N_10081,N_10286);
nor U16788 (N_16788,N_11814,N_11988);
or U16789 (N_16789,N_9233,N_6893);
nand U16790 (N_16790,N_9963,N_9190);
nor U16791 (N_16791,N_6570,N_10095);
nor U16792 (N_16792,N_11538,N_7834);
and U16793 (N_16793,N_6530,N_10666);
nor U16794 (N_16794,N_9338,N_9085);
nand U16795 (N_16795,N_6470,N_7510);
nor U16796 (N_16796,N_8192,N_11967);
or U16797 (N_16797,N_6333,N_11079);
nor U16798 (N_16798,N_6789,N_12144);
nor U16799 (N_16799,N_11444,N_6494);
nand U16800 (N_16800,N_8072,N_11581);
nor U16801 (N_16801,N_7733,N_10445);
nand U16802 (N_16802,N_6415,N_11544);
or U16803 (N_16803,N_11756,N_9932);
nor U16804 (N_16804,N_8026,N_7757);
or U16805 (N_16805,N_9995,N_9366);
and U16806 (N_16806,N_10924,N_12475);
and U16807 (N_16807,N_10373,N_12183);
or U16808 (N_16808,N_11597,N_11540);
or U16809 (N_16809,N_11512,N_8257);
and U16810 (N_16810,N_9092,N_9908);
nor U16811 (N_16811,N_12173,N_9686);
nor U16812 (N_16812,N_8166,N_8862);
nand U16813 (N_16813,N_10220,N_8369);
nand U16814 (N_16814,N_7389,N_8480);
nor U16815 (N_16815,N_12156,N_8251);
nand U16816 (N_16816,N_7583,N_9915);
nor U16817 (N_16817,N_11335,N_11831);
and U16818 (N_16818,N_8867,N_6275);
nor U16819 (N_16819,N_6573,N_7037);
nor U16820 (N_16820,N_7157,N_11134);
or U16821 (N_16821,N_12080,N_8534);
xor U16822 (N_16822,N_7513,N_8707);
nor U16823 (N_16823,N_9673,N_9099);
and U16824 (N_16824,N_7299,N_7144);
nor U16825 (N_16825,N_11835,N_7873);
or U16826 (N_16826,N_9859,N_7912);
nor U16827 (N_16827,N_11870,N_7385);
nand U16828 (N_16828,N_6702,N_6736);
nand U16829 (N_16829,N_12354,N_12123);
nand U16830 (N_16830,N_12135,N_12168);
and U16831 (N_16831,N_7382,N_6749);
and U16832 (N_16832,N_10976,N_8337);
and U16833 (N_16833,N_8106,N_10990);
and U16834 (N_16834,N_11321,N_9804);
nand U16835 (N_16835,N_11849,N_9220);
nor U16836 (N_16836,N_7543,N_7280);
xnor U16837 (N_16837,N_11092,N_10350);
nor U16838 (N_16838,N_10451,N_6821);
nor U16839 (N_16839,N_8607,N_6745);
nor U16840 (N_16840,N_9923,N_6395);
nor U16841 (N_16841,N_8136,N_7876);
and U16842 (N_16842,N_10056,N_9884);
and U16843 (N_16843,N_10890,N_11317);
nand U16844 (N_16844,N_11635,N_10257);
or U16845 (N_16845,N_8079,N_8282);
nand U16846 (N_16846,N_10563,N_10717);
nor U16847 (N_16847,N_8929,N_12011);
and U16848 (N_16848,N_10991,N_12317);
nor U16849 (N_16849,N_11032,N_7269);
and U16850 (N_16850,N_10314,N_10984);
and U16851 (N_16851,N_8216,N_6991);
or U16852 (N_16852,N_11939,N_12397);
or U16853 (N_16853,N_9248,N_12333);
nor U16854 (N_16854,N_8425,N_9668);
or U16855 (N_16855,N_12056,N_8422);
nor U16856 (N_16856,N_10093,N_9257);
and U16857 (N_16857,N_9843,N_12001);
xor U16858 (N_16858,N_7318,N_8366);
or U16859 (N_16859,N_7191,N_10007);
nor U16860 (N_16860,N_6895,N_9429);
and U16861 (N_16861,N_10942,N_9033);
nand U16862 (N_16862,N_9148,N_9729);
nor U16863 (N_16863,N_9165,N_11808);
xor U16864 (N_16864,N_10420,N_10918);
and U16865 (N_16865,N_11314,N_9187);
xnor U16866 (N_16866,N_9862,N_10309);
nand U16867 (N_16867,N_7807,N_6830);
and U16868 (N_16868,N_12190,N_8761);
nor U16869 (N_16869,N_9296,N_10669);
nor U16870 (N_16870,N_6501,N_8588);
nor U16871 (N_16871,N_11440,N_7476);
and U16872 (N_16872,N_7404,N_7833);
nand U16873 (N_16873,N_11371,N_8958);
and U16874 (N_16874,N_6924,N_9849);
or U16875 (N_16875,N_8970,N_7482);
and U16876 (N_16876,N_10775,N_10246);
xnor U16877 (N_16877,N_8527,N_7490);
nand U16878 (N_16878,N_9914,N_10447);
and U16879 (N_16879,N_9698,N_8989);
or U16880 (N_16880,N_12254,N_8877);
nor U16881 (N_16881,N_11987,N_6921);
and U16882 (N_16882,N_11641,N_9766);
or U16883 (N_16883,N_8810,N_12149);
nand U16884 (N_16884,N_10272,N_11916);
nor U16885 (N_16885,N_11313,N_10033);
xor U16886 (N_16886,N_7630,N_10145);
nor U16887 (N_16887,N_8586,N_8470);
nand U16888 (N_16888,N_8719,N_8138);
or U16889 (N_16889,N_9186,N_8894);
or U16890 (N_16890,N_12339,N_10012);
and U16891 (N_16891,N_12149,N_8916);
or U16892 (N_16892,N_7528,N_6379);
or U16893 (N_16893,N_8347,N_9864);
and U16894 (N_16894,N_12190,N_8774);
nor U16895 (N_16895,N_8487,N_7450);
and U16896 (N_16896,N_10925,N_11492);
xor U16897 (N_16897,N_11405,N_10813);
xor U16898 (N_16898,N_8729,N_8716);
and U16899 (N_16899,N_10226,N_10247);
or U16900 (N_16900,N_11608,N_8870);
nor U16901 (N_16901,N_8895,N_10841);
nor U16902 (N_16902,N_7228,N_10245);
nand U16903 (N_16903,N_10023,N_9952);
and U16904 (N_16904,N_11864,N_11833);
and U16905 (N_16905,N_6535,N_6994);
and U16906 (N_16906,N_7075,N_9896);
nand U16907 (N_16907,N_8275,N_10580);
nor U16908 (N_16908,N_11932,N_10622);
or U16909 (N_16909,N_9096,N_10424);
nand U16910 (N_16910,N_11239,N_6441);
nand U16911 (N_16911,N_6869,N_9828);
nor U16912 (N_16912,N_9730,N_6322);
and U16913 (N_16913,N_8058,N_10204);
nand U16914 (N_16914,N_10913,N_9237);
nand U16915 (N_16915,N_8040,N_7688);
or U16916 (N_16916,N_8928,N_9454);
or U16917 (N_16917,N_9316,N_12223);
or U16918 (N_16918,N_7887,N_8293);
and U16919 (N_16919,N_9883,N_9819);
nand U16920 (N_16920,N_8356,N_8895);
nand U16921 (N_16921,N_9446,N_11498);
nor U16922 (N_16922,N_8662,N_7081);
nor U16923 (N_16923,N_8265,N_10301);
xor U16924 (N_16924,N_8101,N_7246);
nand U16925 (N_16925,N_7044,N_9776);
and U16926 (N_16926,N_6762,N_6865);
nand U16927 (N_16927,N_12495,N_8624);
xor U16928 (N_16928,N_12468,N_11482);
nor U16929 (N_16929,N_10628,N_6877);
nand U16930 (N_16930,N_10231,N_12085);
or U16931 (N_16931,N_8458,N_12009);
xor U16932 (N_16932,N_6401,N_10681);
and U16933 (N_16933,N_8994,N_11774);
nor U16934 (N_16934,N_11305,N_8851);
nor U16935 (N_16935,N_10461,N_9727);
nor U16936 (N_16936,N_7169,N_7068);
and U16937 (N_16937,N_6855,N_10471);
and U16938 (N_16938,N_7864,N_9017);
or U16939 (N_16939,N_6804,N_12285);
or U16940 (N_16940,N_9555,N_9038);
and U16941 (N_16941,N_10460,N_7482);
and U16942 (N_16942,N_11256,N_10079);
xor U16943 (N_16943,N_7955,N_8246);
nor U16944 (N_16944,N_9802,N_10000);
nand U16945 (N_16945,N_12051,N_7314);
xor U16946 (N_16946,N_10150,N_9570);
or U16947 (N_16947,N_8378,N_9418);
or U16948 (N_16948,N_7625,N_10481);
nor U16949 (N_16949,N_6331,N_6805);
or U16950 (N_16950,N_11384,N_7447);
and U16951 (N_16951,N_9941,N_11953);
nor U16952 (N_16952,N_12387,N_6922);
and U16953 (N_16953,N_11456,N_8300);
nand U16954 (N_16954,N_12089,N_7395);
or U16955 (N_16955,N_12120,N_10627);
and U16956 (N_16956,N_10262,N_11219);
nand U16957 (N_16957,N_9172,N_11628);
and U16958 (N_16958,N_10657,N_11003);
and U16959 (N_16959,N_6588,N_7935);
xnor U16960 (N_16960,N_8072,N_12228);
nor U16961 (N_16961,N_12445,N_8845);
and U16962 (N_16962,N_8480,N_10129);
or U16963 (N_16963,N_10268,N_6314);
and U16964 (N_16964,N_7255,N_6744);
nand U16965 (N_16965,N_10496,N_7143);
nand U16966 (N_16966,N_10252,N_10835);
nand U16967 (N_16967,N_10163,N_8240);
and U16968 (N_16968,N_11911,N_11355);
nand U16969 (N_16969,N_6677,N_9403);
and U16970 (N_16970,N_9781,N_10395);
or U16971 (N_16971,N_12439,N_7717);
or U16972 (N_16972,N_11190,N_9860);
nor U16973 (N_16973,N_12442,N_8353);
nand U16974 (N_16974,N_9274,N_11243);
nand U16975 (N_16975,N_9539,N_10126);
and U16976 (N_16976,N_12328,N_9118);
or U16977 (N_16977,N_11447,N_6781);
or U16978 (N_16978,N_8404,N_10396);
nor U16979 (N_16979,N_7036,N_11125);
and U16980 (N_16980,N_7114,N_11921);
nor U16981 (N_16981,N_7762,N_10700);
nor U16982 (N_16982,N_9446,N_9880);
and U16983 (N_16983,N_9749,N_6841);
xnor U16984 (N_16984,N_8178,N_8436);
or U16985 (N_16985,N_9149,N_7831);
and U16986 (N_16986,N_9248,N_7769);
nand U16987 (N_16987,N_6588,N_6636);
and U16988 (N_16988,N_10403,N_10294);
xnor U16989 (N_16989,N_10185,N_11110);
nor U16990 (N_16990,N_8696,N_10342);
and U16991 (N_16991,N_7650,N_8902);
or U16992 (N_16992,N_11640,N_10987);
xor U16993 (N_16993,N_6445,N_11374);
nor U16994 (N_16994,N_9036,N_6379);
or U16995 (N_16995,N_9104,N_8401);
nor U16996 (N_16996,N_7402,N_7135);
nor U16997 (N_16997,N_10380,N_12374);
xnor U16998 (N_16998,N_6558,N_8333);
or U16999 (N_16999,N_7634,N_12280);
and U17000 (N_17000,N_11480,N_12141);
nand U17001 (N_17001,N_7157,N_9419);
xnor U17002 (N_17002,N_11401,N_8189);
nor U17003 (N_17003,N_8347,N_8084);
or U17004 (N_17004,N_9429,N_10231);
and U17005 (N_17005,N_7667,N_12233);
and U17006 (N_17006,N_10088,N_6911);
or U17007 (N_17007,N_9059,N_8508);
nand U17008 (N_17008,N_8046,N_10775);
and U17009 (N_17009,N_9753,N_11625);
or U17010 (N_17010,N_8185,N_10767);
xnor U17011 (N_17011,N_8272,N_7790);
or U17012 (N_17012,N_9050,N_11321);
or U17013 (N_17013,N_8062,N_8445);
nor U17014 (N_17014,N_9166,N_7727);
and U17015 (N_17015,N_6808,N_12351);
or U17016 (N_17016,N_11464,N_7540);
and U17017 (N_17017,N_8515,N_7947);
or U17018 (N_17018,N_12274,N_8266);
or U17019 (N_17019,N_7164,N_10787);
and U17020 (N_17020,N_10722,N_10719);
nand U17021 (N_17021,N_11144,N_11992);
and U17022 (N_17022,N_8097,N_8598);
nand U17023 (N_17023,N_9165,N_10063);
and U17024 (N_17024,N_9328,N_10337);
xnor U17025 (N_17025,N_7839,N_8224);
nor U17026 (N_17026,N_7841,N_10095);
nor U17027 (N_17027,N_10006,N_11860);
nor U17028 (N_17028,N_7562,N_7948);
nor U17029 (N_17029,N_7000,N_11081);
and U17030 (N_17030,N_9503,N_9027);
xnor U17031 (N_17031,N_9212,N_7112);
nor U17032 (N_17032,N_12046,N_7851);
or U17033 (N_17033,N_7089,N_6991);
or U17034 (N_17034,N_11503,N_9191);
and U17035 (N_17035,N_10872,N_9571);
nand U17036 (N_17036,N_9716,N_6752);
nand U17037 (N_17037,N_7526,N_11119);
or U17038 (N_17038,N_10248,N_7719);
xnor U17039 (N_17039,N_11710,N_11568);
or U17040 (N_17040,N_10786,N_6493);
and U17041 (N_17041,N_7524,N_8743);
or U17042 (N_17042,N_8615,N_9482);
nand U17043 (N_17043,N_8517,N_9447);
nor U17044 (N_17044,N_8539,N_8607);
nor U17045 (N_17045,N_8737,N_8931);
nor U17046 (N_17046,N_7077,N_10381);
xnor U17047 (N_17047,N_7701,N_9859);
nor U17048 (N_17048,N_12318,N_12406);
or U17049 (N_17049,N_9268,N_10824);
nor U17050 (N_17050,N_9778,N_11373);
and U17051 (N_17051,N_12230,N_11802);
xnor U17052 (N_17052,N_11997,N_8715);
nor U17053 (N_17053,N_10226,N_9203);
xnor U17054 (N_17054,N_11843,N_11778);
nand U17055 (N_17055,N_7666,N_6938);
and U17056 (N_17056,N_7261,N_7313);
nor U17057 (N_17057,N_6474,N_9098);
xor U17058 (N_17058,N_12400,N_8706);
or U17059 (N_17059,N_10406,N_7459);
or U17060 (N_17060,N_7450,N_6765);
nor U17061 (N_17061,N_9006,N_7567);
and U17062 (N_17062,N_11185,N_7157);
or U17063 (N_17063,N_11312,N_6549);
nor U17064 (N_17064,N_6816,N_6286);
or U17065 (N_17065,N_11716,N_9310);
and U17066 (N_17066,N_11211,N_11322);
or U17067 (N_17067,N_10304,N_8791);
or U17068 (N_17068,N_8264,N_6406);
xnor U17069 (N_17069,N_8095,N_10411);
nor U17070 (N_17070,N_9826,N_11651);
or U17071 (N_17071,N_6930,N_9241);
nand U17072 (N_17072,N_9130,N_8007);
xnor U17073 (N_17073,N_10270,N_7801);
nor U17074 (N_17074,N_8831,N_6764);
or U17075 (N_17075,N_10342,N_10731);
and U17076 (N_17076,N_11115,N_8053);
nor U17077 (N_17077,N_9407,N_7194);
nand U17078 (N_17078,N_9359,N_9228);
and U17079 (N_17079,N_11584,N_7694);
or U17080 (N_17080,N_12154,N_12143);
nand U17081 (N_17081,N_9879,N_11248);
or U17082 (N_17082,N_10868,N_10174);
nand U17083 (N_17083,N_12410,N_8247);
or U17084 (N_17084,N_12160,N_6696);
xor U17085 (N_17085,N_9757,N_10576);
nand U17086 (N_17086,N_12418,N_11699);
or U17087 (N_17087,N_10107,N_12288);
nor U17088 (N_17088,N_11228,N_7888);
nor U17089 (N_17089,N_8784,N_10677);
nand U17090 (N_17090,N_7311,N_7596);
nor U17091 (N_17091,N_11941,N_7608);
nand U17092 (N_17092,N_7805,N_7346);
or U17093 (N_17093,N_8654,N_9527);
xnor U17094 (N_17094,N_9277,N_11965);
or U17095 (N_17095,N_8555,N_9675);
nor U17096 (N_17096,N_6685,N_9693);
nand U17097 (N_17097,N_11127,N_11742);
or U17098 (N_17098,N_9960,N_9004);
or U17099 (N_17099,N_9290,N_7128);
or U17100 (N_17100,N_6489,N_6698);
nor U17101 (N_17101,N_8016,N_9786);
nor U17102 (N_17102,N_8573,N_8227);
or U17103 (N_17103,N_11723,N_7137);
nor U17104 (N_17104,N_11435,N_12391);
nand U17105 (N_17105,N_6975,N_11928);
nor U17106 (N_17106,N_7973,N_7448);
and U17107 (N_17107,N_12467,N_8750);
and U17108 (N_17108,N_10095,N_11798);
nand U17109 (N_17109,N_9414,N_6791);
nand U17110 (N_17110,N_7475,N_6382);
or U17111 (N_17111,N_6600,N_12096);
or U17112 (N_17112,N_8011,N_8587);
nand U17113 (N_17113,N_10423,N_7559);
or U17114 (N_17114,N_7707,N_11750);
nor U17115 (N_17115,N_11891,N_9884);
or U17116 (N_17116,N_10343,N_6366);
nand U17117 (N_17117,N_7196,N_11708);
nand U17118 (N_17118,N_8552,N_7802);
nor U17119 (N_17119,N_9694,N_12099);
nand U17120 (N_17120,N_11602,N_8690);
xnor U17121 (N_17121,N_6628,N_11652);
and U17122 (N_17122,N_11783,N_8762);
nor U17123 (N_17123,N_8322,N_6528);
xnor U17124 (N_17124,N_9080,N_12480);
or U17125 (N_17125,N_7428,N_11358);
or U17126 (N_17126,N_12449,N_6880);
nor U17127 (N_17127,N_8563,N_10566);
or U17128 (N_17128,N_9507,N_10183);
nand U17129 (N_17129,N_10494,N_6456);
or U17130 (N_17130,N_6795,N_9640);
nor U17131 (N_17131,N_12270,N_9878);
nand U17132 (N_17132,N_11100,N_7980);
and U17133 (N_17133,N_7108,N_7982);
nand U17134 (N_17134,N_12145,N_11934);
nor U17135 (N_17135,N_9638,N_7619);
or U17136 (N_17136,N_8565,N_12064);
nand U17137 (N_17137,N_9070,N_10536);
nor U17138 (N_17138,N_10309,N_9245);
nor U17139 (N_17139,N_10017,N_6989);
nand U17140 (N_17140,N_10477,N_7123);
or U17141 (N_17141,N_8003,N_11181);
and U17142 (N_17142,N_8622,N_11282);
and U17143 (N_17143,N_7535,N_9772);
or U17144 (N_17144,N_7269,N_8413);
and U17145 (N_17145,N_8942,N_8066);
nor U17146 (N_17146,N_11836,N_8723);
or U17147 (N_17147,N_7135,N_12402);
nor U17148 (N_17148,N_7331,N_11592);
nor U17149 (N_17149,N_10037,N_10955);
and U17150 (N_17150,N_8706,N_7004);
nor U17151 (N_17151,N_9397,N_11584);
and U17152 (N_17152,N_11487,N_11590);
or U17153 (N_17153,N_10881,N_8578);
or U17154 (N_17154,N_6735,N_10384);
nor U17155 (N_17155,N_8037,N_12183);
or U17156 (N_17156,N_9586,N_11546);
nand U17157 (N_17157,N_6889,N_12313);
nor U17158 (N_17158,N_11218,N_6752);
nor U17159 (N_17159,N_9155,N_8215);
or U17160 (N_17160,N_8491,N_6857);
or U17161 (N_17161,N_11149,N_8069);
or U17162 (N_17162,N_10743,N_7939);
and U17163 (N_17163,N_12328,N_9266);
or U17164 (N_17164,N_8310,N_9962);
xnor U17165 (N_17165,N_9141,N_8076);
nor U17166 (N_17166,N_10461,N_8152);
and U17167 (N_17167,N_8083,N_11335);
and U17168 (N_17168,N_11888,N_10004);
nor U17169 (N_17169,N_8152,N_9146);
or U17170 (N_17170,N_11690,N_6609);
or U17171 (N_17171,N_10499,N_6868);
nor U17172 (N_17172,N_7476,N_8669);
nand U17173 (N_17173,N_6995,N_8988);
nand U17174 (N_17174,N_9142,N_8245);
nand U17175 (N_17175,N_12119,N_8135);
nor U17176 (N_17176,N_7989,N_12105);
or U17177 (N_17177,N_8095,N_8399);
or U17178 (N_17178,N_10377,N_7968);
xnor U17179 (N_17179,N_12345,N_11610);
nor U17180 (N_17180,N_10445,N_10051);
nor U17181 (N_17181,N_10453,N_10811);
xor U17182 (N_17182,N_9794,N_7710);
nand U17183 (N_17183,N_11975,N_10053);
or U17184 (N_17184,N_8834,N_10324);
or U17185 (N_17185,N_12208,N_9804);
nor U17186 (N_17186,N_10746,N_11106);
xnor U17187 (N_17187,N_9866,N_10365);
or U17188 (N_17188,N_12290,N_10125);
nand U17189 (N_17189,N_11015,N_10241);
or U17190 (N_17190,N_10240,N_8679);
nand U17191 (N_17191,N_10446,N_8243);
nor U17192 (N_17192,N_7620,N_11322);
or U17193 (N_17193,N_9951,N_11720);
or U17194 (N_17194,N_9394,N_9289);
xor U17195 (N_17195,N_6568,N_7541);
and U17196 (N_17196,N_9407,N_7287);
nand U17197 (N_17197,N_12177,N_9343);
and U17198 (N_17198,N_7090,N_10256);
or U17199 (N_17199,N_7635,N_8680);
nand U17200 (N_17200,N_12189,N_9638);
xor U17201 (N_17201,N_11925,N_11719);
nand U17202 (N_17202,N_10096,N_9198);
and U17203 (N_17203,N_11863,N_12124);
and U17204 (N_17204,N_6396,N_11695);
nand U17205 (N_17205,N_11937,N_9520);
xnor U17206 (N_17206,N_10591,N_7147);
or U17207 (N_17207,N_9170,N_6692);
or U17208 (N_17208,N_9967,N_7858);
or U17209 (N_17209,N_11521,N_10375);
or U17210 (N_17210,N_7037,N_6419);
or U17211 (N_17211,N_7160,N_11981);
or U17212 (N_17212,N_10042,N_9385);
nor U17213 (N_17213,N_11820,N_6421);
nand U17214 (N_17214,N_9537,N_10439);
nand U17215 (N_17215,N_9462,N_12194);
nor U17216 (N_17216,N_6784,N_10154);
nor U17217 (N_17217,N_11997,N_7903);
nand U17218 (N_17218,N_6555,N_7113);
and U17219 (N_17219,N_9308,N_10857);
or U17220 (N_17220,N_6610,N_9194);
nand U17221 (N_17221,N_10951,N_9774);
nor U17222 (N_17222,N_12401,N_10291);
or U17223 (N_17223,N_10648,N_7776);
nor U17224 (N_17224,N_6718,N_12438);
nand U17225 (N_17225,N_11236,N_10109);
nor U17226 (N_17226,N_8206,N_11034);
and U17227 (N_17227,N_7996,N_10486);
or U17228 (N_17228,N_9813,N_11689);
nand U17229 (N_17229,N_11673,N_7138);
or U17230 (N_17230,N_7781,N_7316);
nand U17231 (N_17231,N_11324,N_8002);
or U17232 (N_17232,N_8672,N_11520);
or U17233 (N_17233,N_6605,N_7839);
nand U17234 (N_17234,N_11544,N_11092);
or U17235 (N_17235,N_7437,N_9568);
nor U17236 (N_17236,N_6300,N_10616);
and U17237 (N_17237,N_9977,N_9615);
xor U17238 (N_17238,N_7634,N_8315);
nor U17239 (N_17239,N_8085,N_10179);
xnor U17240 (N_17240,N_11922,N_8472);
and U17241 (N_17241,N_10188,N_8562);
nor U17242 (N_17242,N_11165,N_10530);
nor U17243 (N_17243,N_10225,N_11443);
nand U17244 (N_17244,N_8285,N_11822);
nor U17245 (N_17245,N_7277,N_6541);
nand U17246 (N_17246,N_9811,N_8157);
nor U17247 (N_17247,N_6725,N_7686);
and U17248 (N_17248,N_9163,N_7974);
and U17249 (N_17249,N_6980,N_11808);
xnor U17250 (N_17250,N_11987,N_7059);
or U17251 (N_17251,N_9601,N_9633);
and U17252 (N_17252,N_12479,N_12480);
xor U17253 (N_17253,N_9403,N_6448);
nor U17254 (N_17254,N_10990,N_7355);
nor U17255 (N_17255,N_8751,N_11714);
nor U17256 (N_17256,N_8032,N_10161);
or U17257 (N_17257,N_11252,N_9315);
nand U17258 (N_17258,N_10657,N_8832);
xnor U17259 (N_17259,N_12234,N_6409);
or U17260 (N_17260,N_10103,N_11983);
and U17261 (N_17261,N_6322,N_7518);
or U17262 (N_17262,N_11963,N_9830);
or U17263 (N_17263,N_11247,N_6259);
xnor U17264 (N_17264,N_10646,N_8633);
or U17265 (N_17265,N_9858,N_7949);
and U17266 (N_17266,N_7892,N_9683);
nor U17267 (N_17267,N_7161,N_10099);
nor U17268 (N_17268,N_9219,N_7826);
and U17269 (N_17269,N_7065,N_8274);
and U17270 (N_17270,N_9701,N_9063);
and U17271 (N_17271,N_9242,N_10252);
nor U17272 (N_17272,N_7899,N_10006);
or U17273 (N_17273,N_7897,N_9235);
nor U17274 (N_17274,N_9064,N_10716);
nor U17275 (N_17275,N_10108,N_9533);
and U17276 (N_17276,N_7952,N_10323);
nor U17277 (N_17277,N_9989,N_11676);
nor U17278 (N_17278,N_12024,N_6308);
and U17279 (N_17279,N_8966,N_11605);
nand U17280 (N_17280,N_10329,N_9811);
and U17281 (N_17281,N_11034,N_12226);
nand U17282 (N_17282,N_8810,N_6972);
nor U17283 (N_17283,N_8407,N_7583);
nor U17284 (N_17284,N_7825,N_9759);
or U17285 (N_17285,N_8091,N_8019);
nand U17286 (N_17286,N_7367,N_6980);
and U17287 (N_17287,N_11414,N_10296);
or U17288 (N_17288,N_12370,N_8726);
nor U17289 (N_17289,N_9876,N_11594);
nor U17290 (N_17290,N_11542,N_11683);
xor U17291 (N_17291,N_8478,N_6802);
nand U17292 (N_17292,N_8663,N_9147);
and U17293 (N_17293,N_11556,N_8667);
nand U17294 (N_17294,N_11486,N_6452);
nor U17295 (N_17295,N_10873,N_11287);
or U17296 (N_17296,N_12138,N_12158);
nand U17297 (N_17297,N_9199,N_9878);
or U17298 (N_17298,N_8878,N_8625);
or U17299 (N_17299,N_12396,N_11805);
or U17300 (N_17300,N_10926,N_8469);
and U17301 (N_17301,N_11833,N_8990);
nand U17302 (N_17302,N_12038,N_12426);
nand U17303 (N_17303,N_7139,N_6328);
or U17304 (N_17304,N_12035,N_7373);
nor U17305 (N_17305,N_8036,N_8019);
nand U17306 (N_17306,N_8173,N_6729);
or U17307 (N_17307,N_12027,N_8130);
nand U17308 (N_17308,N_11216,N_6719);
and U17309 (N_17309,N_7312,N_7149);
nor U17310 (N_17310,N_11709,N_11258);
or U17311 (N_17311,N_11662,N_6633);
or U17312 (N_17312,N_6603,N_10750);
xnor U17313 (N_17313,N_7768,N_7049);
xor U17314 (N_17314,N_9810,N_8603);
and U17315 (N_17315,N_11147,N_10776);
nor U17316 (N_17316,N_8981,N_9004);
or U17317 (N_17317,N_9752,N_7006);
and U17318 (N_17318,N_7445,N_10631);
nand U17319 (N_17319,N_6258,N_11266);
nand U17320 (N_17320,N_12429,N_10324);
nor U17321 (N_17321,N_7728,N_12153);
nand U17322 (N_17322,N_6423,N_6400);
nand U17323 (N_17323,N_7721,N_6398);
xor U17324 (N_17324,N_9420,N_12068);
and U17325 (N_17325,N_10049,N_8521);
nand U17326 (N_17326,N_8003,N_7701);
nor U17327 (N_17327,N_7718,N_9279);
or U17328 (N_17328,N_9083,N_10591);
nor U17329 (N_17329,N_9470,N_9078);
and U17330 (N_17330,N_8748,N_11035);
and U17331 (N_17331,N_6994,N_9383);
or U17332 (N_17332,N_9244,N_10511);
nand U17333 (N_17333,N_9044,N_12392);
nand U17334 (N_17334,N_7454,N_11229);
nor U17335 (N_17335,N_7530,N_9178);
xor U17336 (N_17336,N_11602,N_6933);
nand U17337 (N_17337,N_12304,N_10484);
and U17338 (N_17338,N_7599,N_10577);
or U17339 (N_17339,N_12051,N_12156);
nor U17340 (N_17340,N_10268,N_9104);
xnor U17341 (N_17341,N_12142,N_10559);
or U17342 (N_17342,N_6752,N_9337);
or U17343 (N_17343,N_11295,N_8000);
nand U17344 (N_17344,N_10399,N_10686);
nor U17345 (N_17345,N_6871,N_8059);
xnor U17346 (N_17346,N_10464,N_7197);
nor U17347 (N_17347,N_8942,N_10275);
or U17348 (N_17348,N_9908,N_7942);
nand U17349 (N_17349,N_9515,N_6760);
nor U17350 (N_17350,N_9282,N_6271);
or U17351 (N_17351,N_9353,N_11981);
or U17352 (N_17352,N_7988,N_8726);
nand U17353 (N_17353,N_11971,N_8921);
nor U17354 (N_17354,N_9329,N_7474);
and U17355 (N_17355,N_11015,N_11604);
and U17356 (N_17356,N_11313,N_10938);
nor U17357 (N_17357,N_11964,N_7626);
nand U17358 (N_17358,N_11189,N_7570);
nand U17359 (N_17359,N_9170,N_10206);
xor U17360 (N_17360,N_9802,N_7984);
and U17361 (N_17361,N_9861,N_10597);
nor U17362 (N_17362,N_11467,N_12118);
or U17363 (N_17363,N_12312,N_10634);
nand U17364 (N_17364,N_10523,N_7695);
nand U17365 (N_17365,N_9145,N_10261);
nor U17366 (N_17366,N_6614,N_9026);
nand U17367 (N_17367,N_11485,N_7948);
nor U17368 (N_17368,N_10783,N_8454);
nand U17369 (N_17369,N_11541,N_10605);
nand U17370 (N_17370,N_6579,N_12241);
xnor U17371 (N_17371,N_11301,N_10701);
or U17372 (N_17372,N_12085,N_10690);
xor U17373 (N_17373,N_12142,N_12416);
nor U17374 (N_17374,N_11770,N_10443);
nor U17375 (N_17375,N_6337,N_9526);
or U17376 (N_17376,N_11862,N_7926);
xnor U17377 (N_17377,N_9560,N_7818);
and U17378 (N_17378,N_8084,N_6500);
and U17379 (N_17379,N_9930,N_11587);
or U17380 (N_17380,N_8608,N_7401);
and U17381 (N_17381,N_6693,N_9516);
nor U17382 (N_17382,N_11073,N_7096);
xor U17383 (N_17383,N_8878,N_7201);
or U17384 (N_17384,N_10955,N_7137);
nor U17385 (N_17385,N_6945,N_12066);
xor U17386 (N_17386,N_11571,N_10490);
and U17387 (N_17387,N_8037,N_6681);
and U17388 (N_17388,N_7534,N_11258);
and U17389 (N_17389,N_10459,N_6832);
xnor U17390 (N_17390,N_8301,N_6944);
xor U17391 (N_17391,N_10727,N_9316);
and U17392 (N_17392,N_9038,N_7406);
or U17393 (N_17393,N_7765,N_11921);
nor U17394 (N_17394,N_9948,N_10020);
and U17395 (N_17395,N_10450,N_11173);
nor U17396 (N_17396,N_10924,N_8969);
or U17397 (N_17397,N_11707,N_7603);
nor U17398 (N_17398,N_9632,N_6831);
or U17399 (N_17399,N_8875,N_9251);
and U17400 (N_17400,N_11134,N_8579);
and U17401 (N_17401,N_12399,N_8466);
xnor U17402 (N_17402,N_11790,N_6577);
and U17403 (N_17403,N_9174,N_11091);
nor U17404 (N_17404,N_12251,N_10812);
xor U17405 (N_17405,N_10511,N_10408);
nor U17406 (N_17406,N_10787,N_10943);
and U17407 (N_17407,N_7087,N_6929);
xor U17408 (N_17408,N_11529,N_12140);
or U17409 (N_17409,N_10369,N_8181);
xnor U17410 (N_17410,N_7034,N_11865);
nor U17411 (N_17411,N_11439,N_11116);
and U17412 (N_17412,N_12474,N_6807);
or U17413 (N_17413,N_7693,N_6749);
nand U17414 (N_17414,N_7743,N_11491);
nand U17415 (N_17415,N_9301,N_10772);
nor U17416 (N_17416,N_8242,N_11197);
or U17417 (N_17417,N_9546,N_9738);
nor U17418 (N_17418,N_7074,N_7829);
nand U17419 (N_17419,N_8081,N_7479);
nand U17420 (N_17420,N_11197,N_8155);
nor U17421 (N_17421,N_8039,N_7073);
xor U17422 (N_17422,N_11209,N_11984);
and U17423 (N_17423,N_6923,N_10048);
nor U17424 (N_17424,N_8309,N_10281);
or U17425 (N_17425,N_11424,N_10825);
and U17426 (N_17426,N_7189,N_11618);
and U17427 (N_17427,N_10747,N_11163);
nor U17428 (N_17428,N_7264,N_8801);
xor U17429 (N_17429,N_11413,N_6750);
or U17430 (N_17430,N_11390,N_8464);
and U17431 (N_17431,N_8100,N_10364);
nand U17432 (N_17432,N_9981,N_11095);
nand U17433 (N_17433,N_10184,N_11028);
xnor U17434 (N_17434,N_10474,N_11652);
and U17435 (N_17435,N_9398,N_11653);
and U17436 (N_17436,N_9348,N_11509);
nor U17437 (N_17437,N_7528,N_11832);
nand U17438 (N_17438,N_8710,N_10182);
nor U17439 (N_17439,N_11629,N_6798);
xnor U17440 (N_17440,N_11846,N_12185);
nor U17441 (N_17441,N_9891,N_11524);
nand U17442 (N_17442,N_9859,N_9829);
nor U17443 (N_17443,N_7870,N_9420);
xor U17444 (N_17444,N_6730,N_11219);
nand U17445 (N_17445,N_11760,N_10139);
xor U17446 (N_17446,N_6984,N_12473);
or U17447 (N_17447,N_12357,N_7779);
nor U17448 (N_17448,N_7345,N_11248);
or U17449 (N_17449,N_7034,N_8059);
nor U17450 (N_17450,N_10931,N_7928);
xor U17451 (N_17451,N_11459,N_9426);
nor U17452 (N_17452,N_10911,N_6909);
and U17453 (N_17453,N_7562,N_11744);
nand U17454 (N_17454,N_7150,N_8768);
or U17455 (N_17455,N_8427,N_10015);
nand U17456 (N_17456,N_7214,N_6621);
nand U17457 (N_17457,N_12057,N_10113);
or U17458 (N_17458,N_11405,N_7838);
or U17459 (N_17459,N_10193,N_9104);
and U17460 (N_17460,N_9384,N_7439);
nor U17461 (N_17461,N_7480,N_11053);
or U17462 (N_17462,N_6755,N_9913);
or U17463 (N_17463,N_9740,N_9234);
nand U17464 (N_17464,N_12379,N_8176);
and U17465 (N_17465,N_7533,N_9306);
nor U17466 (N_17466,N_8826,N_8105);
or U17467 (N_17467,N_9077,N_12012);
xnor U17468 (N_17468,N_10433,N_9524);
nor U17469 (N_17469,N_9369,N_7227);
or U17470 (N_17470,N_6281,N_11816);
nand U17471 (N_17471,N_9970,N_11381);
xnor U17472 (N_17472,N_7222,N_10310);
nor U17473 (N_17473,N_10359,N_9753);
nor U17474 (N_17474,N_11613,N_8781);
or U17475 (N_17475,N_9408,N_7470);
and U17476 (N_17476,N_6320,N_6968);
or U17477 (N_17477,N_11132,N_9900);
or U17478 (N_17478,N_10261,N_10760);
or U17479 (N_17479,N_9988,N_6590);
or U17480 (N_17480,N_8711,N_9754);
or U17481 (N_17481,N_10030,N_11369);
and U17482 (N_17482,N_11727,N_8959);
or U17483 (N_17483,N_9990,N_6927);
or U17484 (N_17484,N_11190,N_6672);
nand U17485 (N_17485,N_6991,N_11220);
and U17486 (N_17486,N_12158,N_9672);
or U17487 (N_17487,N_7459,N_9665);
nand U17488 (N_17488,N_6905,N_10742);
and U17489 (N_17489,N_8542,N_10455);
nand U17490 (N_17490,N_11971,N_10418);
nand U17491 (N_17491,N_9733,N_7289);
or U17492 (N_17492,N_10422,N_10526);
xor U17493 (N_17493,N_8087,N_10065);
xnor U17494 (N_17494,N_6403,N_8712);
and U17495 (N_17495,N_11735,N_9642);
nand U17496 (N_17496,N_8398,N_12316);
or U17497 (N_17497,N_11497,N_11937);
xor U17498 (N_17498,N_9923,N_11890);
and U17499 (N_17499,N_7255,N_12297);
nor U17500 (N_17500,N_7656,N_8250);
and U17501 (N_17501,N_8754,N_9907);
nand U17502 (N_17502,N_11477,N_8907);
and U17503 (N_17503,N_7480,N_9699);
nand U17504 (N_17504,N_8498,N_9338);
nand U17505 (N_17505,N_11618,N_8651);
nand U17506 (N_17506,N_10757,N_12480);
nand U17507 (N_17507,N_8376,N_9729);
or U17508 (N_17508,N_9732,N_11144);
or U17509 (N_17509,N_10116,N_9232);
nand U17510 (N_17510,N_11332,N_11968);
and U17511 (N_17511,N_10245,N_8698);
or U17512 (N_17512,N_7250,N_11303);
xnor U17513 (N_17513,N_9818,N_8681);
and U17514 (N_17514,N_7734,N_9952);
or U17515 (N_17515,N_6585,N_9838);
nand U17516 (N_17516,N_8601,N_9115);
nor U17517 (N_17517,N_8916,N_9132);
nor U17518 (N_17518,N_6509,N_12110);
nand U17519 (N_17519,N_11844,N_10673);
nor U17520 (N_17520,N_8471,N_11187);
and U17521 (N_17521,N_6486,N_6884);
and U17522 (N_17522,N_9956,N_6702);
nor U17523 (N_17523,N_12445,N_10014);
and U17524 (N_17524,N_10593,N_8595);
and U17525 (N_17525,N_9935,N_10685);
xnor U17526 (N_17526,N_10608,N_10851);
or U17527 (N_17527,N_11482,N_6994);
nand U17528 (N_17528,N_7569,N_8638);
or U17529 (N_17529,N_8489,N_9838);
and U17530 (N_17530,N_7734,N_9505);
and U17531 (N_17531,N_10496,N_10363);
or U17532 (N_17532,N_10708,N_10647);
nand U17533 (N_17533,N_6755,N_7586);
nand U17534 (N_17534,N_9009,N_10998);
or U17535 (N_17535,N_10712,N_8564);
xor U17536 (N_17536,N_6999,N_6631);
nand U17537 (N_17537,N_8723,N_8399);
nand U17538 (N_17538,N_8525,N_9090);
or U17539 (N_17539,N_7580,N_11348);
and U17540 (N_17540,N_11222,N_10242);
or U17541 (N_17541,N_8779,N_9192);
or U17542 (N_17542,N_11299,N_11969);
nor U17543 (N_17543,N_12338,N_9699);
nand U17544 (N_17544,N_8935,N_7183);
nor U17545 (N_17545,N_10571,N_9955);
xor U17546 (N_17546,N_11198,N_7567);
nand U17547 (N_17547,N_11382,N_9045);
and U17548 (N_17548,N_7200,N_7457);
nor U17549 (N_17549,N_8222,N_8166);
and U17550 (N_17550,N_7296,N_11713);
nor U17551 (N_17551,N_10492,N_11637);
or U17552 (N_17552,N_7515,N_7333);
and U17553 (N_17553,N_10331,N_7909);
nor U17554 (N_17554,N_11277,N_10087);
and U17555 (N_17555,N_9659,N_7980);
or U17556 (N_17556,N_10009,N_10787);
nand U17557 (N_17557,N_12142,N_12026);
nand U17558 (N_17558,N_9145,N_10913);
and U17559 (N_17559,N_11966,N_6774);
and U17560 (N_17560,N_11649,N_11154);
and U17561 (N_17561,N_11102,N_8956);
or U17562 (N_17562,N_6919,N_8298);
nand U17563 (N_17563,N_6539,N_9621);
nor U17564 (N_17564,N_6982,N_7910);
or U17565 (N_17565,N_7545,N_9969);
nand U17566 (N_17566,N_6963,N_10300);
nor U17567 (N_17567,N_7946,N_7963);
xnor U17568 (N_17568,N_11231,N_12092);
nor U17569 (N_17569,N_6959,N_6446);
or U17570 (N_17570,N_7707,N_12137);
nand U17571 (N_17571,N_6704,N_12193);
nor U17572 (N_17572,N_6314,N_6263);
xnor U17573 (N_17573,N_12124,N_9458);
nor U17574 (N_17574,N_7537,N_7289);
nor U17575 (N_17575,N_9762,N_9249);
xor U17576 (N_17576,N_12100,N_8083);
nand U17577 (N_17577,N_11968,N_6380);
nor U17578 (N_17578,N_8229,N_10463);
nand U17579 (N_17579,N_9813,N_12192);
xor U17580 (N_17580,N_6815,N_7835);
nor U17581 (N_17581,N_7097,N_12312);
nand U17582 (N_17582,N_12491,N_10968);
and U17583 (N_17583,N_9167,N_10261);
nand U17584 (N_17584,N_6777,N_7574);
nor U17585 (N_17585,N_6254,N_7619);
xor U17586 (N_17586,N_11573,N_9187);
and U17587 (N_17587,N_10329,N_10287);
or U17588 (N_17588,N_8391,N_9243);
and U17589 (N_17589,N_12258,N_6367);
xnor U17590 (N_17590,N_10103,N_12475);
or U17591 (N_17591,N_9500,N_7436);
nor U17592 (N_17592,N_9736,N_9581);
and U17593 (N_17593,N_12491,N_11565);
nor U17594 (N_17594,N_11609,N_11718);
nor U17595 (N_17595,N_11695,N_9711);
xor U17596 (N_17596,N_8879,N_10343);
nor U17597 (N_17597,N_9017,N_7603);
or U17598 (N_17598,N_9450,N_10155);
and U17599 (N_17599,N_11810,N_6365);
or U17600 (N_17600,N_7303,N_11974);
and U17601 (N_17601,N_8466,N_9797);
nand U17602 (N_17602,N_10335,N_9644);
nand U17603 (N_17603,N_10010,N_7754);
nand U17604 (N_17604,N_11378,N_10025);
nand U17605 (N_17605,N_9165,N_8636);
or U17606 (N_17606,N_9809,N_10321);
nand U17607 (N_17607,N_9723,N_7192);
nor U17608 (N_17608,N_10396,N_8724);
and U17609 (N_17609,N_9066,N_11718);
nand U17610 (N_17610,N_10742,N_6305);
xor U17611 (N_17611,N_6768,N_12426);
and U17612 (N_17612,N_8181,N_7632);
nand U17613 (N_17613,N_10624,N_10839);
or U17614 (N_17614,N_8026,N_7350);
and U17615 (N_17615,N_9403,N_7961);
xnor U17616 (N_17616,N_9956,N_9497);
xnor U17617 (N_17617,N_10785,N_11802);
nor U17618 (N_17618,N_10079,N_6862);
xor U17619 (N_17619,N_9305,N_7011);
nor U17620 (N_17620,N_10184,N_10850);
and U17621 (N_17621,N_6859,N_6583);
or U17622 (N_17622,N_10048,N_9534);
nand U17623 (N_17623,N_7334,N_11629);
nand U17624 (N_17624,N_10458,N_9456);
and U17625 (N_17625,N_8142,N_8224);
nor U17626 (N_17626,N_10307,N_9412);
or U17627 (N_17627,N_9028,N_6918);
and U17628 (N_17628,N_6270,N_7003);
and U17629 (N_17629,N_6709,N_6424);
and U17630 (N_17630,N_9543,N_6748);
nor U17631 (N_17631,N_12030,N_9736);
and U17632 (N_17632,N_6900,N_7851);
nand U17633 (N_17633,N_6643,N_9845);
xnor U17634 (N_17634,N_7593,N_11722);
or U17635 (N_17635,N_10685,N_11874);
nor U17636 (N_17636,N_9345,N_10111);
nor U17637 (N_17637,N_7222,N_11029);
xor U17638 (N_17638,N_6532,N_9732);
nor U17639 (N_17639,N_8630,N_9699);
and U17640 (N_17640,N_11679,N_11531);
nor U17641 (N_17641,N_7781,N_10923);
nand U17642 (N_17642,N_6771,N_11284);
or U17643 (N_17643,N_9617,N_12185);
nand U17644 (N_17644,N_6929,N_7002);
nor U17645 (N_17645,N_9595,N_9435);
nor U17646 (N_17646,N_10087,N_7634);
nand U17647 (N_17647,N_6934,N_12139);
nor U17648 (N_17648,N_9949,N_7936);
or U17649 (N_17649,N_10436,N_8798);
and U17650 (N_17650,N_7164,N_8702);
nor U17651 (N_17651,N_9613,N_7696);
nor U17652 (N_17652,N_10356,N_11535);
and U17653 (N_17653,N_11789,N_10623);
or U17654 (N_17654,N_11979,N_10289);
or U17655 (N_17655,N_6910,N_12464);
or U17656 (N_17656,N_10706,N_10599);
nor U17657 (N_17657,N_8133,N_8109);
or U17658 (N_17658,N_9811,N_7734);
or U17659 (N_17659,N_12430,N_9495);
nor U17660 (N_17660,N_6498,N_10634);
or U17661 (N_17661,N_9783,N_9201);
or U17662 (N_17662,N_6989,N_6661);
and U17663 (N_17663,N_12351,N_8065);
xor U17664 (N_17664,N_6669,N_11949);
nor U17665 (N_17665,N_6539,N_6711);
and U17666 (N_17666,N_8692,N_12097);
and U17667 (N_17667,N_12251,N_9002);
nand U17668 (N_17668,N_10978,N_6693);
or U17669 (N_17669,N_7105,N_11075);
nor U17670 (N_17670,N_11524,N_12338);
and U17671 (N_17671,N_9595,N_9135);
and U17672 (N_17672,N_7847,N_9783);
and U17673 (N_17673,N_8701,N_9109);
nand U17674 (N_17674,N_9606,N_12292);
and U17675 (N_17675,N_12169,N_11636);
nand U17676 (N_17676,N_8891,N_9947);
nor U17677 (N_17677,N_10470,N_7794);
nand U17678 (N_17678,N_10259,N_11498);
xor U17679 (N_17679,N_8765,N_9921);
nand U17680 (N_17680,N_8719,N_9713);
xor U17681 (N_17681,N_9326,N_9541);
and U17682 (N_17682,N_10590,N_10126);
nand U17683 (N_17683,N_12275,N_9375);
nand U17684 (N_17684,N_12294,N_12077);
xnor U17685 (N_17685,N_8560,N_9726);
and U17686 (N_17686,N_8099,N_9675);
nand U17687 (N_17687,N_6917,N_9829);
xor U17688 (N_17688,N_11395,N_12302);
nand U17689 (N_17689,N_12013,N_8690);
and U17690 (N_17690,N_6923,N_7993);
and U17691 (N_17691,N_7804,N_6466);
nand U17692 (N_17692,N_8070,N_8591);
or U17693 (N_17693,N_10278,N_6373);
or U17694 (N_17694,N_8753,N_7264);
and U17695 (N_17695,N_11978,N_7856);
or U17696 (N_17696,N_11354,N_7520);
xor U17697 (N_17697,N_7096,N_12094);
or U17698 (N_17698,N_8988,N_7520);
nand U17699 (N_17699,N_9227,N_7211);
nand U17700 (N_17700,N_11922,N_8916);
nand U17701 (N_17701,N_11057,N_9466);
and U17702 (N_17702,N_9022,N_6372);
and U17703 (N_17703,N_7375,N_12476);
or U17704 (N_17704,N_12258,N_10901);
nand U17705 (N_17705,N_10971,N_9283);
or U17706 (N_17706,N_9501,N_10294);
and U17707 (N_17707,N_8098,N_8325);
and U17708 (N_17708,N_7951,N_6310);
or U17709 (N_17709,N_10727,N_9971);
nor U17710 (N_17710,N_10157,N_12296);
and U17711 (N_17711,N_7112,N_10662);
xnor U17712 (N_17712,N_8347,N_11862);
xnor U17713 (N_17713,N_7545,N_9030);
xnor U17714 (N_17714,N_7444,N_7135);
or U17715 (N_17715,N_8729,N_10070);
or U17716 (N_17716,N_7184,N_8630);
or U17717 (N_17717,N_11109,N_9403);
nor U17718 (N_17718,N_12091,N_10428);
and U17719 (N_17719,N_7315,N_10446);
or U17720 (N_17720,N_6664,N_11999);
nor U17721 (N_17721,N_8388,N_8912);
nand U17722 (N_17722,N_7478,N_8467);
nand U17723 (N_17723,N_7653,N_7172);
or U17724 (N_17724,N_9883,N_7793);
xnor U17725 (N_17725,N_11928,N_11386);
or U17726 (N_17726,N_7116,N_8357);
and U17727 (N_17727,N_12499,N_12157);
nor U17728 (N_17728,N_11205,N_11172);
or U17729 (N_17729,N_9245,N_8749);
and U17730 (N_17730,N_8964,N_12008);
nor U17731 (N_17731,N_6646,N_11629);
nand U17732 (N_17732,N_7975,N_10673);
xnor U17733 (N_17733,N_11289,N_6600);
or U17734 (N_17734,N_7448,N_10981);
nand U17735 (N_17735,N_11119,N_9778);
nand U17736 (N_17736,N_12246,N_7908);
nand U17737 (N_17737,N_11070,N_11893);
and U17738 (N_17738,N_6547,N_9848);
nand U17739 (N_17739,N_6711,N_10393);
xnor U17740 (N_17740,N_11806,N_10594);
and U17741 (N_17741,N_10374,N_6700);
or U17742 (N_17742,N_10912,N_6666);
nor U17743 (N_17743,N_7713,N_6828);
nor U17744 (N_17744,N_8940,N_8547);
nand U17745 (N_17745,N_9703,N_7296);
nand U17746 (N_17746,N_8527,N_9911);
or U17747 (N_17747,N_6450,N_7186);
nand U17748 (N_17748,N_11413,N_6407);
nor U17749 (N_17749,N_8388,N_12096);
and U17750 (N_17750,N_8162,N_7930);
xor U17751 (N_17751,N_7339,N_9493);
nor U17752 (N_17752,N_12498,N_7645);
nand U17753 (N_17753,N_10496,N_7780);
and U17754 (N_17754,N_9919,N_8976);
and U17755 (N_17755,N_9495,N_7651);
and U17756 (N_17756,N_10217,N_11205);
or U17757 (N_17757,N_8060,N_12084);
nor U17758 (N_17758,N_7670,N_12441);
or U17759 (N_17759,N_8943,N_9897);
nor U17760 (N_17760,N_12025,N_11269);
or U17761 (N_17761,N_11275,N_9308);
or U17762 (N_17762,N_6756,N_7206);
xnor U17763 (N_17763,N_11262,N_6442);
and U17764 (N_17764,N_10807,N_7847);
and U17765 (N_17765,N_7224,N_10732);
and U17766 (N_17766,N_10384,N_9328);
nor U17767 (N_17767,N_10234,N_6502);
nor U17768 (N_17768,N_6646,N_7768);
nand U17769 (N_17769,N_6764,N_10290);
or U17770 (N_17770,N_6640,N_7828);
nor U17771 (N_17771,N_11668,N_11663);
or U17772 (N_17772,N_11076,N_9479);
xor U17773 (N_17773,N_7103,N_11692);
xnor U17774 (N_17774,N_11863,N_11179);
nand U17775 (N_17775,N_11556,N_9572);
nand U17776 (N_17776,N_10741,N_11875);
nor U17777 (N_17777,N_6768,N_9924);
or U17778 (N_17778,N_10739,N_11268);
nor U17779 (N_17779,N_7650,N_8140);
nor U17780 (N_17780,N_9283,N_8743);
and U17781 (N_17781,N_9956,N_8033);
and U17782 (N_17782,N_12136,N_7653);
or U17783 (N_17783,N_6646,N_12171);
and U17784 (N_17784,N_10758,N_7136);
xor U17785 (N_17785,N_7564,N_10779);
and U17786 (N_17786,N_10959,N_8019);
nor U17787 (N_17787,N_7287,N_8959);
and U17788 (N_17788,N_9674,N_9785);
and U17789 (N_17789,N_9675,N_12367);
and U17790 (N_17790,N_8564,N_6325);
nor U17791 (N_17791,N_6760,N_11693);
nor U17792 (N_17792,N_8668,N_6259);
and U17793 (N_17793,N_8511,N_7991);
nor U17794 (N_17794,N_9462,N_6922);
nor U17795 (N_17795,N_10114,N_7169);
or U17796 (N_17796,N_7152,N_9973);
or U17797 (N_17797,N_9600,N_10057);
and U17798 (N_17798,N_6918,N_6889);
or U17799 (N_17799,N_7461,N_9992);
nor U17800 (N_17800,N_9488,N_9277);
or U17801 (N_17801,N_6607,N_10188);
nand U17802 (N_17802,N_10468,N_7975);
or U17803 (N_17803,N_7268,N_11993);
nand U17804 (N_17804,N_10335,N_6716);
nand U17805 (N_17805,N_10182,N_9948);
xnor U17806 (N_17806,N_8753,N_7430);
nor U17807 (N_17807,N_9870,N_9153);
xnor U17808 (N_17808,N_10107,N_10904);
and U17809 (N_17809,N_10463,N_11132);
and U17810 (N_17810,N_6525,N_11097);
xor U17811 (N_17811,N_8140,N_7167);
nor U17812 (N_17812,N_6790,N_7148);
or U17813 (N_17813,N_12365,N_7078);
nand U17814 (N_17814,N_10458,N_10192);
and U17815 (N_17815,N_12239,N_7014);
xnor U17816 (N_17816,N_9124,N_7757);
or U17817 (N_17817,N_6636,N_10452);
or U17818 (N_17818,N_10894,N_6636);
nor U17819 (N_17819,N_11606,N_10546);
or U17820 (N_17820,N_10903,N_6290);
and U17821 (N_17821,N_6303,N_11055);
or U17822 (N_17822,N_10036,N_8487);
nor U17823 (N_17823,N_8215,N_11306);
nor U17824 (N_17824,N_10821,N_10653);
or U17825 (N_17825,N_9109,N_11972);
nor U17826 (N_17826,N_6491,N_11258);
nand U17827 (N_17827,N_11889,N_9545);
and U17828 (N_17828,N_12396,N_8382);
nor U17829 (N_17829,N_11004,N_6609);
nor U17830 (N_17830,N_12467,N_10461);
or U17831 (N_17831,N_10046,N_11682);
and U17832 (N_17832,N_10274,N_6970);
nor U17833 (N_17833,N_9893,N_7087);
nor U17834 (N_17834,N_11953,N_9190);
and U17835 (N_17835,N_12431,N_8398);
xor U17836 (N_17836,N_7448,N_10844);
and U17837 (N_17837,N_11001,N_10401);
or U17838 (N_17838,N_10176,N_8177);
nor U17839 (N_17839,N_6541,N_8738);
or U17840 (N_17840,N_7059,N_8794);
nand U17841 (N_17841,N_7749,N_9357);
nand U17842 (N_17842,N_7729,N_8295);
nor U17843 (N_17843,N_10333,N_8811);
or U17844 (N_17844,N_11217,N_6602);
and U17845 (N_17845,N_7970,N_9066);
and U17846 (N_17846,N_11010,N_9522);
or U17847 (N_17847,N_11841,N_7664);
nand U17848 (N_17848,N_6336,N_7802);
or U17849 (N_17849,N_11030,N_7177);
or U17850 (N_17850,N_7027,N_9224);
nor U17851 (N_17851,N_6611,N_10065);
and U17852 (N_17852,N_6949,N_8404);
and U17853 (N_17853,N_11135,N_8312);
or U17854 (N_17854,N_11633,N_10750);
or U17855 (N_17855,N_7192,N_11209);
and U17856 (N_17856,N_9319,N_6981);
xor U17857 (N_17857,N_9775,N_9793);
or U17858 (N_17858,N_8554,N_7929);
xor U17859 (N_17859,N_8460,N_11672);
nand U17860 (N_17860,N_7053,N_10409);
and U17861 (N_17861,N_10667,N_9726);
xnor U17862 (N_17862,N_9733,N_7238);
nand U17863 (N_17863,N_10221,N_7469);
nor U17864 (N_17864,N_10620,N_11351);
or U17865 (N_17865,N_11679,N_10537);
nand U17866 (N_17866,N_7433,N_6374);
nand U17867 (N_17867,N_8570,N_6854);
nand U17868 (N_17868,N_12094,N_10479);
nand U17869 (N_17869,N_11250,N_10907);
and U17870 (N_17870,N_7554,N_9242);
and U17871 (N_17871,N_10666,N_11640);
and U17872 (N_17872,N_6617,N_9051);
and U17873 (N_17873,N_11006,N_9367);
and U17874 (N_17874,N_7731,N_10033);
and U17875 (N_17875,N_7988,N_11519);
or U17876 (N_17876,N_8531,N_8022);
and U17877 (N_17877,N_7286,N_11188);
nand U17878 (N_17878,N_6402,N_7021);
and U17879 (N_17879,N_11300,N_12420);
nor U17880 (N_17880,N_8954,N_8499);
nand U17881 (N_17881,N_10103,N_6624);
nand U17882 (N_17882,N_9689,N_12023);
xor U17883 (N_17883,N_7493,N_11770);
nand U17884 (N_17884,N_12306,N_6494);
or U17885 (N_17885,N_11550,N_7972);
nor U17886 (N_17886,N_8702,N_8781);
nor U17887 (N_17887,N_7701,N_7175);
nor U17888 (N_17888,N_10286,N_7213);
xor U17889 (N_17889,N_9233,N_8757);
and U17890 (N_17890,N_6304,N_11304);
nand U17891 (N_17891,N_8758,N_10935);
nand U17892 (N_17892,N_8769,N_9922);
nand U17893 (N_17893,N_9934,N_9628);
xor U17894 (N_17894,N_7889,N_10308);
nor U17895 (N_17895,N_7196,N_9425);
nand U17896 (N_17896,N_10148,N_9233);
and U17897 (N_17897,N_10838,N_10325);
and U17898 (N_17898,N_11237,N_6929);
and U17899 (N_17899,N_10211,N_12248);
and U17900 (N_17900,N_10166,N_11476);
nor U17901 (N_17901,N_7528,N_8717);
and U17902 (N_17902,N_8015,N_12050);
nand U17903 (N_17903,N_11710,N_8786);
nand U17904 (N_17904,N_9871,N_7189);
nand U17905 (N_17905,N_6609,N_10658);
xnor U17906 (N_17906,N_11211,N_7857);
nand U17907 (N_17907,N_7385,N_10630);
nor U17908 (N_17908,N_8922,N_8307);
and U17909 (N_17909,N_11019,N_8309);
or U17910 (N_17910,N_11341,N_9971);
or U17911 (N_17911,N_10950,N_7615);
nor U17912 (N_17912,N_7540,N_9514);
nor U17913 (N_17913,N_11422,N_10822);
nor U17914 (N_17914,N_11631,N_11006);
or U17915 (N_17915,N_7831,N_10013);
nand U17916 (N_17916,N_11483,N_6558);
xnor U17917 (N_17917,N_10953,N_10821);
nor U17918 (N_17918,N_11720,N_10574);
xor U17919 (N_17919,N_11131,N_8161);
nor U17920 (N_17920,N_8437,N_6759);
nand U17921 (N_17921,N_10460,N_7182);
nor U17922 (N_17922,N_6661,N_10930);
and U17923 (N_17923,N_11517,N_11833);
nand U17924 (N_17924,N_11145,N_10995);
nor U17925 (N_17925,N_7187,N_12051);
nand U17926 (N_17926,N_10633,N_6565);
nor U17927 (N_17927,N_7344,N_11573);
xor U17928 (N_17928,N_9763,N_7781);
xor U17929 (N_17929,N_7661,N_10413);
nor U17930 (N_17930,N_6760,N_9629);
or U17931 (N_17931,N_8083,N_6285);
or U17932 (N_17932,N_12019,N_9133);
xnor U17933 (N_17933,N_9445,N_8328);
nand U17934 (N_17934,N_10202,N_11023);
nor U17935 (N_17935,N_10800,N_9496);
or U17936 (N_17936,N_6276,N_10880);
nand U17937 (N_17937,N_6386,N_8718);
nor U17938 (N_17938,N_10296,N_7204);
or U17939 (N_17939,N_9247,N_7907);
or U17940 (N_17940,N_7226,N_10660);
nand U17941 (N_17941,N_10689,N_6689);
nand U17942 (N_17942,N_10001,N_7951);
nor U17943 (N_17943,N_8267,N_11539);
nand U17944 (N_17944,N_11685,N_7847);
nand U17945 (N_17945,N_7764,N_10720);
xnor U17946 (N_17946,N_6893,N_7235);
nand U17947 (N_17947,N_11635,N_10261);
nand U17948 (N_17948,N_10500,N_8132);
or U17949 (N_17949,N_12415,N_9847);
or U17950 (N_17950,N_7341,N_6265);
nand U17951 (N_17951,N_9745,N_6701);
or U17952 (N_17952,N_11239,N_7089);
nand U17953 (N_17953,N_12418,N_8916);
nand U17954 (N_17954,N_7690,N_7404);
and U17955 (N_17955,N_8377,N_10146);
nand U17956 (N_17956,N_7181,N_7949);
nand U17957 (N_17957,N_6789,N_7593);
nor U17958 (N_17958,N_11593,N_7867);
or U17959 (N_17959,N_9857,N_8155);
xnor U17960 (N_17960,N_8431,N_11126);
nor U17961 (N_17961,N_9274,N_9862);
and U17962 (N_17962,N_7727,N_11423);
or U17963 (N_17963,N_6833,N_7436);
nor U17964 (N_17964,N_9258,N_11198);
or U17965 (N_17965,N_9684,N_11955);
nand U17966 (N_17966,N_7732,N_10722);
nor U17967 (N_17967,N_9033,N_9463);
nand U17968 (N_17968,N_12412,N_12036);
nand U17969 (N_17969,N_8872,N_9391);
nor U17970 (N_17970,N_6682,N_11306);
nor U17971 (N_17971,N_6760,N_8099);
or U17972 (N_17972,N_9068,N_6525);
nor U17973 (N_17973,N_11116,N_8968);
nand U17974 (N_17974,N_10621,N_9138);
nor U17975 (N_17975,N_11858,N_6419);
and U17976 (N_17976,N_11010,N_11415);
and U17977 (N_17977,N_6700,N_9782);
or U17978 (N_17978,N_9436,N_11940);
nand U17979 (N_17979,N_9600,N_9175);
or U17980 (N_17980,N_7921,N_10400);
and U17981 (N_17981,N_8101,N_9565);
xor U17982 (N_17982,N_11889,N_9743);
xor U17983 (N_17983,N_8108,N_12464);
nand U17984 (N_17984,N_8910,N_6750);
nand U17985 (N_17985,N_7649,N_11831);
and U17986 (N_17986,N_7254,N_8698);
nand U17987 (N_17987,N_6293,N_10310);
nand U17988 (N_17988,N_7160,N_12292);
or U17989 (N_17989,N_12483,N_7691);
nor U17990 (N_17990,N_9664,N_8367);
or U17991 (N_17991,N_7407,N_7506);
or U17992 (N_17992,N_7977,N_11039);
or U17993 (N_17993,N_10799,N_8913);
and U17994 (N_17994,N_9408,N_8121);
and U17995 (N_17995,N_9362,N_6951);
or U17996 (N_17996,N_8889,N_10093);
or U17997 (N_17997,N_12065,N_9948);
xor U17998 (N_17998,N_6470,N_10346);
nand U17999 (N_17999,N_7962,N_7321);
xnor U18000 (N_18000,N_7318,N_12476);
nand U18001 (N_18001,N_12233,N_11378);
and U18002 (N_18002,N_8675,N_7001);
and U18003 (N_18003,N_10258,N_6282);
xor U18004 (N_18004,N_8355,N_6622);
or U18005 (N_18005,N_9578,N_12131);
xnor U18006 (N_18006,N_7945,N_9776);
or U18007 (N_18007,N_8362,N_8335);
or U18008 (N_18008,N_7314,N_11806);
nor U18009 (N_18009,N_10269,N_9224);
nand U18010 (N_18010,N_6283,N_9301);
and U18011 (N_18011,N_9704,N_7235);
nor U18012 (N_18012,N_11987,N_12414);
or U18013 (N_18013,N_7354,N_9842);
or U18014 (N_18014,N_12476,N_8272);
and U18015 (N_18015,N_8683,N_11160);
and U18016 (N_18016,N_11910,N_12248);
and U18017 (N_18017,N_7516,N_7134);
nand U18018 (N_18018,N_12356,N_10676);
or U18019 (N_18019,N_10520,N_10224);
and U18020 (N_18020,N_7630,N_11054);
or U18021 (N_18021,N_9461,N_9607);
or U18022 (N_18022,N_10929,N_9818);
and U18023 (N_18023,N_7902,N_6730);
xnor U18024 (N_18024,N_12017,N_10083);
nand U18025 (N_18025,N_12198,N_11229);
nor U18026 (N_18026,N_10525,N_10124);
nand U18027 (N_18027,N_10834,N_11301);
and U18028 (N_18028,N_6631,N_6582);
nor U18029 (N_18029,N_7353,N_7965);
or U18030 (N_18030,N_8410,N_9115);
nand U18031 (N_18031,N_11971,N_8006);
xnor U18032 (N_18032,N_9563,N_10020);
nand U18033 (N_18033,N_11953,N_6959);
xnor U18034 (N_18034,N_6851,N_11667);
nand U18035 (N_18035,N_12181,N_11025);
nand U18036 (N_18036,N_10821,N_9327);
and U18037 (N_18037,N_11221,N_11303);
and U18038 (N_18038,N_7967,N_8354);
nor U18039 (N_18039,N_10849,N_12414);
nand U18040 (N_18040,N_8914,N_9576);
and U18041 (N_18041,N_9525,N_7326);
and U18042 (N_18042,N_10899,N_7110);
nor U18043 (N_18043,N_11997,N_6878);
and U18044 (N_18044,N_7072,N_6645);
and U18045 (N_18045,N_11097,N_6463);
or U18046 (N_18046,N_10370,N_9391);
nand U18047 (N_18047,N_9067,N_9120);
and U18048 (N_18048,N_8326,N_10096);
nand U18049 (N_18049,N_11414,N_10132);
or U18050 (N_18050,N_10748,N_11400);
and U18051 (N_18051,N_11423,N_6427);
nor U18052 (N_18052,N_10629,N_6793);
xor U18053 (N_18053,N_8719,N_9333);
nor U18054 (N_18054,N_9888,N_12183);
or U18055 (N_18055,N_10742,N_6572);
or U18056 (N_18056,N_11567,N_11674);
or U18057 (N_18057,N_11808,N_7573);
nand U18058 (N_18058,N_9960,N_6922);
xnor U18059 (N_18059,N_8220,N_7631);
nand U18060 (N_18060,N_7475,N_10169);
and U18061 (N_18061,N_11899,N_7096);
or U18062 (N_18062,N_10663,N_9364);
nor U18063 (N_18063,N_7607,N_6730);
nor U18064 (N_18064,N_8981,N_9806);
and U18065 (N_18065,N_8793,N_10845);
nor U18066 (N_18066,N_9345,N_9837);
and U18067 (N_18067,N_7533,N_10111);
or U18068 (N_18068,N_12239,N_7428);
and U18069 (N_18069,N_12415,N_11784);
nor U18070 (N_18070,N_6612,N_6335);
nor U18071 (N_18071,N_11559,N_8036);
nand U18072 (N_18072,N_11339,N_9036);
and U18073 (N_18073,N_6963,N_11135);
xnor U18074 (N_18074,N_8242,N_12492);
or U18075 (N_18075,N_8705,N_10908);
xnor U18076 (N_18076,N_11016,N_9722);
and U18077 (N_18077,N_11559,N_11476);
or U18078 (N_18078,N_9544,N_9305);
nor U18079 (N_18079,N_9900,N_6349);
and U18080 (N_18080,N_10399,N_7531);
nand U18081 (N_18081,N_9789,N_8007);
and U18082 (N_18082,N_8538,N_8469);
or U18083 (N_18083,N_6935,N_7343);
or U18084 (N_18084,N_9260,N_9704);
or U18085 (N_18085,N_9622,N_9706);
and U18086 (N_18086,N_10680,N_7087);
nand U18087 (N_18087,N_11702,N_7004);
nand U18088 (N_18088,N_12258,N_12123);
and U18089 (N_18089,N_10922,N_12487);
nor U18090 (N_18090,N_10851,N_8320);
nand U18091 (N_18091,N_9299,N_12165);
and U18092 (N_18092,N_7007,N_10057);
or U18093 (N_18093,N_8185,N_8277);
and U18094 (N_18094,N_8628,N_10048);
and U18095 (N_18095,N_7653,N_10574);
and U18096 (N_18096,N_9997,N_9811);
nand U18097 (N_18097,N_11305,N_9213);
nand U18098 (N_18098,N_11497,N_7672);
or U18099 (N_18099,N_7082,N_8629);
and U18100 (N_18100,N_8302,N_9860);
xnor U18101 (N_18101,N_10460,N_8634);
nor U18102 (N_18102,N_8904,N_8107);
nand U18103 (N_18103,N_11590,N_8282);
nand U18104 (N_18104,N_6695,N_8060);
or U18105 (N_18105,N_12145,N_10409);
xor U18106 (N_18106,N_12462,N_8667);
or U18107 (N_18107,N_9365,N_9162);
xnor U18108 (N_18108,N_6531,N_7283);
nand U18109 (N_18109,N_7879,N_7339);
and U18110 (N_18110,N_8811,N_6565);
nand U18111 (N_18111,N_7659,N_8615);
and U18112 (N_18112,N_11609,N_11817);
nand U18113 (N_18113,N_9418,N_10522);
nand U18114 (N_18114,N_7267,N_10345);
and U18115 (N_18115,N_11696,N_6332);
or U18116 (N_18116,N_6546,N_8340);
nand U18117 (N_18117,N_12375,N_9885);
or U18118 (N_18118,N_10305,N_8771);
nor U18119 (N_18119,N_8602,N_10032);
nor U18120 (N_18120,N_9648,N_11594);
nor U18121 (N_18121,N_8025,N_8468);
or U18122 (N_18122,N_10215,N_10780);
nor U18123 (N_18123,N_8700,N_10056);
or U18124 (N_18124,N_9817,N_7042);
or U18125 (N_18125,N_8872,N_8037);
or U18126 (N_18126,N_12054,N_9616);
xor U18127 (N_18127,N_10124,N_7738);
nand U18128 (N_18128,N_12156,N_11992);
nor U18129 (N_18129,N_10390,N_7832);
nand U18130 (N_18130,N_9983,N_8569);
and U18131 (N_18131,N_10463,N_11237);
nand U18132 (N_18132,N_7341,N_8188);
or U18133 (N_18133,N_8316,N_11170);
xor U18134 (N_18134,N_10027,N_10221);
xor U18135 (N_18135,N_9207,N_12108);
nand U18136 (N_18136,N_7994,N_11234);
nor U18137 (N_18137,N_6968,N_6711);
or U18138 (N_18138,N_8566,N_9099);
nand U18139 (N_18139,N_12075,N_10150);
nand U18140 (N_18140,N_9506,N_10192);
nand U18141 (N_18141,N_10916,N_9326);
nand U18142 (N_18142,N_9456,N_8108);
nand U18143 (N_18143,N_6867,N_11524);
xor U18144 (N_18144,N_7260,N_11718);
and U18145 (N_18145,N_7355,N_8231);
nand U18146 (N_18146,N_11233,N_8518);
or U18147 (N_18147,N_10486,N_6702);
or U18148 (N_18148,N_8088,N_7376);
nor U18149 (N_18149,N_11221,N_12330);
or U18150 (N_18150,N_11334,N_11191);
nand U18151 (N_18151,N_10425,N_8310);
nand U18152 (N_18152,N_9008,N_6375);
nor U18153 (N_18153,N_8484,N_10097);
xor U18154 (N_18154,N_11276,N_9141);
nor U18155 (N_18155,N_9189,N_7388);
or U18156 (N_18156,N_7183,N_7470);
nand U18157 (N_18157,N_7125,N_11287);
or U18158 (N_18158,N_8086,N_12457);
nand U18159 (N_18159,N_10211,N_11907);
and U18160 (N_18160,N_9362,N_8794);
nor U18161 (N_18161,N_9120,N_8206);
and U18162 (N_18162,N_7662,N_9564);
nand U18163 (N_18163,N_11253,N_6444);
or U18164 (N_18164,N_8884,N_6336);
xnor U18165 (N_18165,N_8728,N_6760);
nand U18166 (N_18166,N_11918,N_8930);
and U18167 (N_18167,N_8065,N_7774);
nor U18168 (N_18168,N_8959,N_10296);
and U18169 (N_18169,N_7234,N_9406);
nor U18170 (N_18170,N_8428,N_10617);
or U18171 (N_18171,N_9466,N_10015);
nand U18172 (N_18172,N_8374,N_10057);
nand U18173 (N_18173,N_9743,N_7719);
nor U18174 (N_18174,N_11552,N_7300);
nor U18175 (N_18175,N_8779,N_6562);
nor U18176 (N_18176,N_7081,N_10177);
nand U18177 (N_18177,N_11165,N_8910);
and U18178 (N_18178,N_7792,N_11079);
and U18179 (N_18179,N_7114,N_10337);
nand U18180 (N_18180,N_7391,N_9829);
nor U18181 (N_18181,N_10175,N_9758);
or U18182 (N_18182,N_9172,N_12309);
nor U18183 (N_18183,N_10462,N_9591);
and U18184 (N_18184,N_9886,N_11236);
and U18185 (N_18185,N_7744,N_11753);
nor U18186 (N_18186,N_6911,N_11288);
nor U18187 (N_18187,N_10146,N_10740);
or U18188 (N_18188,N_8698,N_8980);
nand U18189 (N_18189,N_8071,N_8735);
or U18190 (N_18190,N_9323,N_9448);
nand U18191 (N_18191,N_8002,N_7555);
nor U18192 (N_18192,N_10597,N_7196);
nor U18193 (N_18193,N_10336,N_7173);
nand U18194 (N_18194,N_6401,N_11875);
or U18195 (N_18195,N_6505,N_10656);
and U18196 (N_18196,N_7745,N_7154);
or U18197 (N_18197,N_6918,N_8459);
nand U18198 (N_18198,N_6283,N_7371);
nor U18199 (N_18199,N_6251,N_8950);
or U18200 (N_18200,N_7867,N_9112);
nor U18201 (N_18201,N_10854,N_9398);
nor U18202 (N_18202,N_6332,N_7434);
xnor U18203 (N_18203,N_10180,N_6843);
nor U18204 (N_18204,N_7084,N_8494);
or U18205 (N_18205,N_10003,N_11330);
or U18206 (N_18206,N_11982,N_8723);
nor U18207 (N_18207,N_12023,N_9710);
and U18208 (N_18208,N_10982,N_6474);
and U18209 (N_18209,N_12117,N_7288);
and U18210 (N_18210,N_10049,N_9026);
nand U18211 (N_18211,N_12298,N_8950);
and U18212 (N_18212,N_9163,N_6284);
and U18213 (N_18213,N_11027,N_10273);
nand U18214 (N_18214,N_7365,N_8587);
and U18215 (N_18215,N_11836,N_7150);
nand U18216 (N_18216,N_9154,N_12076);
nand U18217 (N_18217,N_12325,N_12170);
xor U18218 (N_18218,N_10717,N_11819);
nor U18219 (N_18219,N_7482,N_10997);
nand U18220 (N_18220,N_6599,N_11816);
or U18221 (N_18221,N_7671,N_9814);
and U18222 (N_18222,N_8649,N_10325);
or U18223 (N_18223,N_10164,N_8128);
nand U18224 (N_18224,N_7051,N_8186);
or U18225 (N_18225,N_8368,N_7361);
xor U18226 (N_18226,N_9657,N_11759);
nor U18227 (N_18227,N_11573,N_9580);
and U18228 (N_18228,N_7919,N_9745);
and U18229 (N_18229,N_10253,N_9104);
nor U18230 (N_18230,N_9977,N_8832);
or U18231 (N_18231,N_12143,N_10087);
nand U18232 (N_18232,N_11163,N_8535);
or U18233 (N_18233,N_12302,N_11502);
and U18234 (N_18234,N_12131,N_8637);
or U18235 (N_18235,N_8036,N_10307);
nand U18236 (N_18236,N_9181,N_7265);
nand U18237 (N_18237,N_6812,N_9343);
or U18238 (N_18238,N_11688,N_9815);
nand U18239 (N_18239,N_11356,N_9684);
or U18240 (N_18240,N_7030,N_12370);
or U18241 (N_18241,N_12469,N_11030);
nor U18242 (N_18242,N_11087,N_8771);
and U18243 (N_18243,N_12152,N_10887);
nand U18244 (N_18244,N_9602,N_7716);
or U18245 (N_18245,N_9257,N_7023);
nor U18246 (N_18246,N_6873,N_6607);
xor U18247 (N_18247,N_8979,N_7486);
xor U18248 (N_18248,N_9653,N_12481);
and U18249 (N_18249,N_8024,N_9778);
xnor U18250 (N_18250,N_8962,N_7421);
nor U18251 (N_18251,N_9915,N_6877);
nor U18252 (N_18252,N_10321,N_9417);
nand U18253 (N_18253,N_8475,N_7614);
nand U18254 (N_18254,N_7844,N_12060);
nor U18255 (N_18255,N_8416,N_9265);
nor U18256 (N_18256,N_12254,N_9987);
xnor U18257 (N_18257,N_10826,N_8976);
xnor U18258 (N_18258,N_11495,N_9056);
nand U18259 (N_18259,N_8545,N_10220);
xor U18260 (N_18260,N_6380,N_10066);
or U18261 (N_18261,N_12434,N_8459);
and U18262 (N_18262,N_7037,N_10233);
nor U18263 (N_18263,N_9073,N_6655);
nor U18264 (N_18264,N_6693,N_7855);
or U18265 (N_18265,N_7690,N_12246);
or U18266 (N_18266,N_7346,N_9369);
nor U18267 (N_18267,N_6967,N_7945);
xnor U18268 (N_18268,N_6807,N_11647);
nor U18269 (N_18269,N_10264,N_8518);
and U18270 (N_18270,N_11225,N_8537);
nor U18271 (N_18271,N_8655,N_10235);
and U18272 (N_18272,N_8988,N_12128);
and U18273 (N_18273,N_10301,N_11496);
nand U18274 (N_18274,N_6808,N_9769);
nor U18275 (N_18275,N_8599,N_10785);
and U18276 (N_18276,N_9027,N_7842);
and U18277 (N_18277,N_11290,N_10192);
nand U18278 (N_18278,N_6358,N_8394);
nand U18279 (N_18279,N_8834,N_8806);
nand U18280 (N_18280,N_6869,N_11028);
nand U18281 (N_18281,N_6867,N_9467);
and U18282 (N_18282,N_10764,N_7840);
and U18283 (N_18283,N_12487,N_12258);
nor U18284 (N_18284,N_7208,N_10305);
and U18285 (N_18285,N_10144,N_6782);
nor U18286 (N_18286,N_12451,N_7921);
nor U18287 (N_18287,N_10226,N_9577);
or U18288 (N_18288,N_11454,N_10176);
and U18289 (N_18289,N_6255,N_6457);
nand U18290 (N_18290,N_8640,N_6434);
nand U18291 (N_18291,N_9305,N_12045);
or U18292 (N_18292,N_9419,N_9525);
nor U18293 (N_18293,N_8903,N_9687);
nand U18294 (N_18294,N_10816,N_11974);
and U18295 (N_18295,N_9376,N_12398);
nor U18296 (N_18296,N_11685,N_10908);
or U18297 (N_18297,N_9309,N_9525);
nor U18298 (N_18298,N_8739,N_6593);
or U18299 (N_18299,N_11978,N_11785);
or U18300 (N_18300,N_7013,N_10932);
nor U18301 (N_18301,N_10755,N_7680);
xnor U18302 (N_18302,N_7868,N_11055);
and U18303 (N_18303,N_6910,N_12203);
and U18304 (N_18304,N_10702,N_7900);
nand U18305 (N_18305,N_8806,N_6852);
xnor U18306 (N_18306,N_9209,N_9210);
nor U18307 (N_18307,N_8575,N_8806);
or U18308 (N_18308,N_6314,N_8133);
nor U18309 (N_18309,N_6263,N_8339);
or U18310 (N_18310,N_9020,N_7908);
or U18311 (N_18311,N_8937,N_10164);
or U18312 (N_18312,N_7346,N_8386);
or U18313 (N_18313,N_10575,N_12169);
nand U18314 (N_18314,N_6934,N_9398);
nand U18315 (N_18315,N_12048,N_9883);
nor U18316 (N_18316,N_6871,N_9527);
xnor U18317 (N_18317,N_7646,N_7683);
or U18318 (N_18318,N_11710,N_6655);
and U18319 (N_18319,N_8853,N_6751);
and U18320 (N_18320,N_8615,N_9019);
nand U18321 (N_18321,N_7556,N_11015);
xnor U18322 (N_18322,N_6791,N_11326);
or U18323 (N_18323,N_6712,N_10118);
nor U18324 (N_18324,N_6585,N_10069);
or U18325 (N_18325,N_9959,N_8392);
nor U18326 (N_18326,N_10578,N_8813);
nand U18327 (N_18327,N_12153,N_8412);
nand U18328 (N_18328,N_10690,N_11546);
nor U18329 (N_18329,N_10186,N_8767);
nor U18330 (N_18330,N_9829,N_9486);
nor U18331 (N_18331,N_6627,N_8132);
nand U18332 (N_18332,N_7181,N_9496);
or U18333 (N_18333,N_6522,N_7286);
or U18334 (N_18334,N_8003,N_7544);
xnor U18335 (N_18335,N_8036,N_7134);
or U18336 (N_18336,N_12153,N_12241);
or U18337 (N_18337,N_11408,N_9215);
nand U18338 (N_18338,N_12065,N_7854);
or U18339 (N_18339,N_11343,N_11610);
nand U18340 (N_18340,N_9657,N_8219);
xnor U18341 (N_18341,N_6832,N_11579);
and U18342 (N_18342,N_6568,N_12225);
or U18343 (N_18343,N_8958,N_9225);
and U18344 (N_18344,N_8715,N_6995);
nor U18345 (N_18345,N_9065,N_8894);
or U18346 (N_18346,N_10106,N_11997);
and U18347 (N_18347,N_9952,N_9795);
nor U18348 (N_18348,N_9465,N_6822);
nand U18349 (N_18349,N_10252,N_8192);
nand U18350 (N_18350,N_9119,N_6616);
nor U18351 (N_18351,N_12148,N_9772);
or U18352 (N_18352,N_11156,N_9790);
and U18353 (N_18353,N_9703,N_8167);
or U18354 (N_18354,N_6665,N_7605);
or U18355 (N_18355,N_8362,N_9620);
or U18356 (N_18356,N_11853,N_7371);
nand U18357 (N_18357,N_8055,N_8024);
xnor U18358 (N_18358,N_8477,N_6666);
or U18359 (N_18359,N_9309,N_12339);
nand U18360 (N_18360,N_7986,N_8772);
xnor U18361 (N_18361,N_8356,N_8279);
nand U18362 (N_18362,N_8342,N_11733);
xnor U18363 (N_18363,N_12095,N_7340);
nand U18364 (N_18364,N_12389,N_12000);
nor U18365 (N_18365,N_6977,N_12189);
and U18366 (N_18366,N_8458,N_10727);
or U18367 (N_18367,N_10766,N_7376);
and U18368 (N_18368,N_12178,N_8940);
nor U18369 (N_18369,N_9981,N_8275);
and U18370 (N_18370,N_8983,N_12278);
nor U18371 (N_18371,N_8280,N_9388);
nor U18372 (N_18372,N_11814,N_7880);
and U18373 (N_18373,N_6455,N_6442);
xor U18374 (N_18374,N_9959,N_7715);
and U18375 (N_18375,N_10135,N_7496);
xnor U18376 (N_18376,N_10100,N_8103);
and U18377 (N_18377,N_7587,N_8650);
or U18378 (N_18378,N_11893,N_7153);
or U18379 (N_18379,N_10517,N_12190);
and U18380 (N_18380,N_7087,N_6501);
or U18381 (N_18381,N_9684,N_9853);
or U18382 (N_18382,N_7397,N_10233);
or U18383 (N_18383,N_9629,N_7141);
and U18384 (N_18384,N_9276,N_11605);
nor U18385 (N_18385,N_11315,N_8649);
or U18386 (N_18386,N_9072,N_6387);
xor U18387 (N_18387,N_8296,N_12284);
and U18388 (N_18388,N_9990,N_11105);
or U18389 (N_18389,N_8239,N_7135);
or U18390 (N_18390,N_8041,N_7609);
or U18391 (N_18391,N_10227,N_6630);
or U18392 (N_18392,N_11520,N_11863);
or U18393 (N_18393,N_11328,N_9500);
nand U18394 (N_18394,N_8801,N_10606);
nor U18395 (N_18395,N_9498,N_11124);
and U18396 (N_18396,N_8946,N_12343);
nand U18397 (N_18397,N_8697,N_10529);
nand U18398 (N_18398,N_9667,N_8711);
and U18399 (N_18399,N_7353,N_9341);
nand U18400 (N_18400,N_11771,N_9655);
nor U18401 (N_18401,N_12429,N_8747);
nor U18402 (N_18402,N_6719,N_7781);
xnor U18403 (N_18403,N_8787,N_8010);
nor U18404 (N_18404,N_12122,N_11509);
or U18405 (N_18405,N_6969,N_9209);
or U18406 (N_18406,N_10082,N_10569);
xor U18407 (N_18407,N_7129,N_12248);
and U18408 (N_18408,N_10316,N_10538);
or U18409 (N_18409,N_10552,N_10957);
nand U18410 (N_18410,N_8453,N_12361);
nor U18411 (N_18411,N_11560,N_9742);
and U18412 (N_18412,N_10867,N_11657);
and U18413 (N_18413,N_8137,N_12220);
or U18414 (N_18414,N_10650,N_12461);
and U18415 (N_18415,N_8976,N_11802);
and U18416 (N_18416,N_11839,N_12407);
and U18417 (N_18417,N_8036,N_10770);
and U18418 (N_18418,N_8123,N_10499);
nor U18419 (N_18419,N_10094,N_11857);
nor U18420 (N_18420,N_10787,N_9645);
or U18421 (N_18421,N_8638,N_7621);
and U18422 (N_18422,N_12179,N_12312);
nor U18423 (N_18423,N_9978,N_10997);
and U18424 (N_18424,N_11217,N_7928);
and U18425 (N_18425,N_8688,N_8441);
or U18426 (N_18426,N_11554,N_8541);
nand U18427 (N_18427,N_10107,N_8370);
and U18428 (N_18428,N_11098,N_6883);
nand U18429 (N_18429,N_9923,N_9530);
nor U18430 (N_18430,N_11090,N_9453);
nand U18431 (N_18431,N_11798,N_6965);
nand U18432 (N_18432,N_11900,N_10341);
nor U18433 (N_18433,N_11750,N_8793);
or U18434 (N_18434,N_9193,N_11645);
nand U18435 (N_18435,N_11089,N_9261);
and U18436 (N_18436,N_10918,N_12072);
nor U18437 (N_18437,N_8098,N_10108);
nand U18438 (N_18438,N_11835,N_8442);
and U18439 (N_18439,N_12321,N_9054);
and U18440 (N_18440,N_11970,N_8238);
nor U18441 (N_18441,N_12093,N_7885);
and U18442 (N_18442,N_8046,N_9119);
nor U18443 (N_18443,N_10152,N_12114);
nand U18444 (N_18444,N_11212,N_7545);
and U18445 (N_18445,N_8222,N_10702);
nand U18446 (N_18446,N_9966,N_6330);
nor U18447 (N_18447,N_8222,N_11566);
nor U18448 (N_18448,N_6659,N_6691);
nand U18449 (N_18449,N_7712,N_6875);
nand U18450 (N_18450,N_6489,N_8521);
and U18451 (N_18451,N_9950,N_7295);
nor U18452 (N_18452,N_10636,N_7269);
and U18453 (N_18453,N_11797,N_11586);
nand U18454 (N_18454,N_7277,N_10749);
nand U18455 (N_18455,N_9055,N_10405);
nand U18456 (N_18456,N_12089,N_6728);
nor U18457 (N_18457,N_7847,N_8561);
or U18458 (N_18458,N_10662,N_9735);
or U18459 (N_18459,N_9327,N_9845);
or U18460 (N_18460,N_6660,N_12411);
xor U18461 (N_18461,N_11193,N_12430);
nor U18462 (N_18462,N_8743,N_10248);
nand U18463 (N_18463,N_11608,N_11767);
nand U18464 (N_18464,N_6317,N_6879);
nand U18465 (N_18465,N_7523,N_9778);
or U18466 (N_18466,N_11572,N_12012);
or U18467 (N_18467,N_12499,N_8711);
xor U18468 (N_18468,N_8333,N_12372);
xor U18469 (N_18469,N_8139,N_11491);
xor U18470 (N_18470,N_10892,N_6550);
or U18471 (N_18471,N_11940,N_6619);
or U18472 (N_18472,N_11236,N_12315);
xnor U18473 (N_18473,N_7857,N_9006);
and U18474 (N_18474,N_9186,N_10841);
xor U18475 (N_18475,N_11949,N_8025);
nor U18476 (N_18476,N_8142,N_6810);
nand U18477 (N_18477,N_8588,N_7721);
nor U18478 (N_18478,N_9966,N_10086);
and U18479 (N_18479,N_9967,N_8948);
nor U18480 (N_18480,N_12252,N_6903);
and U18481 (N_18481,N_9835,N_11807);
or U18482 (N_18482,N_11400,N_12174);
nand U18483 (N_18483,N_8748,N_8050);
nand U18484 (N_18484,N_9214,N_9422);
nand U18485 (N_18485,N_8143,N_9630);
nor U18486 (N_18486,N_7782,N_10396);
nand U18487 (N_18487,N_8621,N_9285);
and U18488 (N_18488,N_12183,N_11843);
nand U18489 (N_18489,N_8653,N_12361);
and U18490 (N_18490,N_10253,N_6335);
nor U18491 (N_18491,N_8218,N_11339);
or U18492 (N_18492,N_8258,N_6982);
nor U18493 (N_18493,N_9043,N_6952);
nor U18494 (N_18494,N_8962,N_8264);
nor U18495 (N_18495,N_7034,N_7688);
and U18496 (N_18496,N_10804,N_10953);
and U18497 (N_18497,N_6908,N_9069);
or U18498 (N_18498,N_9958,N_8953);
or U18499 (N_18499,N_10859,N_6910);
nor U18500 (N_18500,N_11854,N_8650);
and U18501 (N_18501,N_12088,N_7263);
or U18502 (N_18502,N_11102,N_8323);
or U18503 (N_18503,N_12199,N_8075);
and U18504 (N_18504,N_11264,N_8621);
nand U18505 (N_18505,N_6697,N_10027);
or U18506 (N_18506,N_12242,N_12310);
nand U18507 (N_18507,N_10967,N_11178);
nor U18508 (N_18508,N_11060,N_9967);
nor U18509 (N_18509,N_8953,N_12471);
or U18510 (N_18510,N_9605,N_12184);
nand U18511 (N_18511,N_12068,N_6966);
or U18512 (N_18512,N_7510,N_7129);
xnor U18513 (N_18513,N_8436,N_11996);
and U18514 (N_18514,N_11244,N_12304);
and U18515 (N_18515,N_8685,N_8821);
nor U18516 (N_18516,N_10424,N_9798);
nor U18517 (N_18517,N_8842,N_11550);
or U18518 (N_18518,N_7038,N_6648);
nand U18519 (N_18519,N_10288,N_12259);
and U18520 (N_18520,N_6384,N_11653);
and U18521 (N_18521,N_9165,N_8699);
nand U18522 (N_18522,N_10860,N_11220);
or U18523 (N_18523,N_12396,N_9034);
and U18524 (N_18524,N_8013,N_11594);
xor U18525 (N_18525,N_6262,N_10942);
and U18526 (N_18526,N_11574,N_8884);
or U18527 (N_18527,N_11028,N_8916);
or U18528 (N_18528,N_9522,N_9735);
nand U18529 (N_18529,N_6460,N_10521);
nor U18530 (N_18530,N_6704,N_7731);
or U18531 (N_18531,N_9287,N_10276);
xnor U18532 (N_18532,N_10580,N_11190);
or U18533 (N_18533,N_8308,N_7382);
nor U18534 (N_18534,N_8888,N_11005);
nor U18535 (N_18535,N_8785,N_9451);
or U18536 (N_18536,N_10066,N_10470);
nand U18537 (N_18537,N_7256,N_10518);
nor U18538 (N_18538,N_7855,N_7861);
xor U18539 (N_18539,N_7865,N_11769);
or U18540 (N_18540,N_7572,N_7720);
nor U18541 (N_18541,N_6281,N_8030);
and U18542 (N_18542,N_9106,N_9778);
xnor U18543 (N_18543,N_11785,N_10589);
and U18544 (N_18544,N_8367,N_7439);
and U18545 (N_18545,N_9980,N_6297);
nor U18546 (N_18546,N_8510,N_10700);
nor U18547 (N_18547,N_8082,N_9773);
xnor U18548 (N_18548,N_7123,N_10194);
and U18549 (N_18549,N_7960,N_7246);
nor U18550 (N_18550,N_9411,N_11856);
nor U18551 (N_18551,N_6405,N_10027);
nor U18552 (N_18552,N_12018,N_6683);
or U18553 (N_18553,N_7484,N_9651);
xnor U18554 (N_18554,N_6640,N_12369);
nand U18555 (N_18555,N_8747,N_11608);
and U18556 (N_18556,N_6538,N_8179);
and U18557 (N_18557,N_11624,N_11778);
nor U18558 (N_18558,N_11556,N_10201);
nand U18559 (N_18559,N_6335,N_12432);
nor U18560 (N_18560,N_11482,N_9361);
and U18561 (N_18561,N_9892,N_11634);
nor U18562 (N_18562,N_8477,N_11550);
xor U18563 (N_18563,N_7059,N_12395);
or U18564 (N_18564,N_8152,N_10313);
or U18565 (N_18565,N_6813,N_6720);
nand U18566 (N_18566,N_6495,N_7835);
xor U18567 (N_18567,N_12402,N_10533);
or U18568 (N_18568,N_8906,N_7506);
nor U18569 (N_18569,N_7410,N_7717);
and U18570 (N_18570,N_11635,N_6458);
nand U18571 (N_18571,N_12059,N_6534);
xnor U18572 (N_18572,N_7675,N_8520);
xnor U18573 (N_18573,N_8213,N_9236);
nor U18574 (N_18574,N_11802,N_8494);
or U18575 (N_18575,N_7146,N_7636);
or U18576 (N_18576,N_9476,N_7716);
or U18577 (N_18577,N_10918,N_9564);
nor U18578 (N_18578,N_7336,N_7529);
or U18579 (N_18579,N_9587,N_8367);
nand U18580 (N_18580,N_8145,N_8804);
or U18581 (N_18581,N_8182,N_11047);
nor U18582 (N_18582,N_8760,N_12017);
nor U18583 (N_18583,N_6776,N_11583);
nand U18584 (N_18584,N_11826,N_7430);
xnor U18585 (N_18585,N_6719,N_6509);
and U18586 (N_18586,N_7694,N_12089);
and U18587 (N_18587,N_9429,N_8749);
nor U18588 (N_18588,N_7600,N_10482);
nand U18589 (N_18589,N_7146,N_11172);
nor U18590 (N_18590,N_12199,N_9703);
nand U18591 (N_18591,N_11223,N_8525);
nor U18592 (N_18592,N_7549,N_11730);
nand U18593 (N_18593,N_9660,N_7734);
nor U18594 (N_18594,N_10704,N_8556);
nand U18595 (N_18595,N_7417,N_8018);
xor U18596 (N_18596,N_9961,N_9505);
xnor U18597 (N_18597,N_10944,N_9407);
and U18598 (N_18598,N_9165,N_10829);
nor U18599 (N_18599,N_6526,N_6967);
and U18600 (N_18600,N_11145,N_12095);
and U18601 (N_18601,N_9246,N_9280);
xor U18602 (N_18602,N_11573,N_10070);
or U18603 (N_18603,N_11590,N_6719);
nand U18604 (N_18604,N_8999,N_10370);
or U18605 (N_18605,N_10047,N_9530);
xor U18606 (N_18606,N_12039,N_7960);
xor U18607 (N_18607,N_9119,N_6791);
or U18608 (N_18608,N_9803,N_9122);
nand U18609 (N_18609,N_11012,N_11024);
or U18610 (N_18610,N_7725,N_12045);
nand U18611 (N_18611,N_11927,N_9390);
nor U18612 (N_18612,N_9244,N_6843);
nor U18613 (N_18613,N_12436,N_8648);
nor U18614 (N_18614,N_9471,N_6419);
nand U18615 (N_18615,N_9543,N_12220);
or U18616 (N_18616,N_6349,N_11532);
nor U18617 (N_18617,N_10278,N_6942);
and U18618 (N_18618,N_9328,N_7173);
or U18619 (N_18619,N_11197,N_6583);
and U18620 (N_18620,N_12284,N_8769);
and U18621 (N_18621,N_8201,N_9020);
and U18622 (N_18622,N_12323,N_12488);
nor U18623 (N_18623,N_10955,N_6357);
nand U18624 (N_18624,N_7454,N_8733);
and U18625 (N_18625,N_10210,N_9898);
and U18626 (N_18626,N_6968,N_9856);
and U18627 (N_18627,N_6757,N_8809);
and U18628 (N_18628,N_9509,N_6420);
or U18629 (N_18629,N_9708,N_11601);
xnor U18630 (N_18630,N_6637,N_9263);
and U18631 (N_18631,N_11787,N_10578);
and U18632 (N_18632,N_12031,N_7066);
nand U18633 (N_18633,N_8455,N_10652);
and U18634 (N_18634,N_6519,N_10322);
nor U18635 (N_18635,N_9036,N_10780);
nor U18636 (N_18636,N_7071,N_12323);
and U18637 (N_18637,N_12392,N_7373);
and U18638 (N_18638,N_9113,N_11016);
nand U18639 (N_18639,N_7398,N_8518);
nor U18640 (N_18640,N_12114,N_7527);
and U18641 (N_18641,N_6574,N_7502);
nand U18642 (N_18642,N_6904,N_10055);
nand U18643 (N_18643,N_11158,N_8762);
and U18644 (N_18644,N_12197,N_6574);
or U18645 (N_18645,N_10098,N_8450);
nor U18646 (N_18646,N_8507,N_7655);
nor U18647 (N_18647,N_7247,N_10703);
or U18648 (N_18648,N_10867,N_11090);
nand U18649 (N_18649,N_7076,N_8812);
and U18650 (N_18650,N_12241,N_9085);
nand U18651 (N_18651,N_7612,N_11181);
nand U18652 (N_18652,N_10334,N_9519);
nor U18653 (N_18653,N_6860,N_9316);
nor U18654 (N_18654,N_6810,N_9804);
and U18655 (N_18655,N_7689,N_10436);
xor U18656 (N_18656,N_8559,N_6840);
or U18657 (N_18657,N_10591,N_8414);
or U18658 (N_18658,N_8640,N_10625);
nor U18659 (N_18659,N_11768,N_8419);
nor U18660 (N_18660,N_7069,N_8058);
nor U18661 (N_18661,N_9532,N_10286);
or U18662 (N_18662,N_9320,N_6656);
nand U18663 (N_18663,N_11950,N_8130);
and U18664 (N_18664,N_8446,N_9503);
or U18665 (N_18665,N_12483,N_8140);
or U18666 (N_18666,N_8752,N_10135);
nor U18667 (N_18667,N_7956,N_6251);
xor U18668 (N_18668,N_9543,N_11593);
nand U18669 (N_18669,N_10687,N_8472);
or U18670 (N_18670,N_9327,N_6447);
or U18671 (N_18671,N_8750,N_12459);
nand U18672 (N_18672,N_10356,N_7061);
nor U18673 (N_18673,N_7622,N_7085);
nor U18674 (N_18674,N_11304,N_11925);
and U18675 (N_18675,N_12389,N_8839);
xor U18676 (N_18676,N_8375,N_7130);
nand U18677 (N_18677,N_6715,N_9899);
or U18678 (N_18678,N_8515,N_10152);
nand U18679 (N_18679,N_12222,N_7816);
nand U18680 (N_18680,N_7507,N_8607);
and U18681 (N_18681,N_8866,N_9867);
or U18682 (N_18682,N_9900,N_7721);
nand U18683 (N_18683,N_10491,N_10385);
or U18684 (N_18684,N_6395,N_8144);
or U18685 (N_18685,N_7278,N_9204);
or U18686 (N_18686,N_11899,N_9382);
nor U18687 (N_18687,N_6605,N_12372);
and U18688 (N_18688,N_11337,N_8765);
and U18689 (N_18689,N_9966,N_6358);
xnor U18690 (N_18690,N_7178,N_11569);
nand U18691 (N_18691,N_8112,N_7660);
and U18692 (N_18692,N_11078,N_9852);
or U18693 (N_18693,N_11976,N_8637);
nand U18694 (N_18694,N_6969,N_10374);
nand U18695 (N_18695,N_6772,N_10829);
nor U18696 (N_18696,N_6587,N_9357);
nand U18697 (N_18697,N_6852,N_6797);
and U18698 (N_18698,N_11440,N_8875);
nor U18699 (N_18699,N_6633,N_11903);
nand U18700 (N_18700,N_8410,N_11535);
and U18701 (N_18701,N_9726,N_12302);
nand U18702 (N_18702,N_11707,N_6471);
nor U18703 (N_18703,N_8067,N_9635);
nor U18704 (N_18704,N_9115,N_10015);
nand U18705 (N_18705,N_6757,N_12170);
nor U18706 (N_18706,N_6953,N_10831);
nor U18707 (N_18707,N_8780,N_9679);
nor U18708 (N_18708,N_8923,N_9862);
or U18709 (N_18709,N_7208,N_11264);
and U18710 (N_18710,N_8495,N_11126);
nor U18711 (N_18711,N_10334,N_12415);
nand U18712 (N_18712,N_7296,N_11677);
xor U18713 (N_18713,N_6480,N_9745);
nand U18714 (N_18714,N_10656,N_10240);
nand U18715 (N_18715,N_12329,N_10670);
nor U18716 (N_18716,N_10334,N_11411);
nor U18717 (N_18717,N_12071,N_6452);
nor U18718 (N_18718,N_7310,N_10641);
nand U18719 (N_18719,N_6895,N_10030);
nand U18720 (N_18720,N_9362,N_12048);
nor U18721 (N_18721,N_7511,N_6718);
nor U18722 (N_18722,N_9569,N_8351);
nor U18723 (N_18723,N_8038,N_10833);
nor U18724 (N_18724,N_9911,N_9804);
and U18725 (N_18725,N_7695,N_6351);
nor U18726 (N_18726,N_11068,N_7695);
and U18727 (N_18727,N_9814,N_8255);
nand U18728 (N_18728,N_10857,N_11577);
xnor U18729 (N_18729,N_12399,N_8608);
nor U18730 (N_18730,N_10422,N_11588);
xor U18731 (N_18731,N_11843,N_11270);
nand U18732 (N_18732,N_12018,N_11683);
nor U18733 (N_18733,N_7314,N_10526);
nor U18734 (N_18734,N_10987,N_11245);
and U18735 (N_18735,N_9032,N_10019);
nor U18736 (N_18736,N_7450,N_11371);
xnor U18737 (N_18737,N_8603,N_11185);
or U18738 (N_18738,N_6961,N_8118);
nand U18739 (N_18739,N_9712,N_10896);
xor U18740 (N_18740,N_11742,N_11847);
nor U18741 (N_18741,N_10408,N_11031);
nor U18742 (N_18742,N_11552,N_12050);
xnor U18743 (N_18743,N_9564,N_9239);
nor U18744 (N_18744,N_10454,N_11396);
and U18745 (N_18745,N_8747,N_7177);
or U18746 (N_18746,N_6725,N_12431);
or U18747 (N_18747,N_9709,N_8111);
or U18748 (N_18748,N_8623,N_8195);
and U18749 (N_18749,N_10069,N_7036);
nor U18750 (N_18750,N_13870,N_16175);
nand U18751 (N_18751,N_15399,N_14077);
and U18752 (N_18752,N_14537,N_13733);
and U18753 (N_18753,N_14159,N_13620);
or U18754 (N_18754,N_13812,N_17960);
nand U18755 (N_18755,N_17321,N_18023);
nor U18756 (N_18756,N_18369,N_15508);
nand U18757 (N_18757,N_13234,N_17518);
xor U18758 (N_18758,N_15126,N_12916);
nor U18759 (N_18759,N_16650,N_13946);
nand U18760 (N_18760,N_16696,N_16584);
nand U18761 (N_18761,N_18375,N_15385);
nor U18762 (N_18762,N_17229,N_12649);
nor U18763 (N_18763,N_16321,N_13227);
xor U18764 (N_18764,N_18464,N_12630);
nor U18765 (N_18765,N_12516,N_15251);
nor U18766 (N_18766,N_17428,N_12781);
nand U18767 (N_18767,N_18113,N_16064);
nand U18768 (N_18768,N_16658,N_14706);
nor U18769 (N_18769,N_16425,N_15105);
and U18770 (N_18770,N_13862,N_14490);
nand U18771 (N_18771,N_13831,N_13873);
nand U18772 (N_18772,N_14853,N_15575);
nor U18773 (N_18773,N_14171,N_18471);
and U18774 (N_18774,N_14338,N_14111);
xnor U18775 (N_18775,N_17882,N_14367);
nand U18776 (N_18776,N_16940,N_16597);
nor U18777 (N_18777,N_12895,N_15987);
nor U18778 (N_18778,N_17963,N_12741);
nor U18779 (N_18779,N_18094,N_12521);
and U18780 (N_18780,N_17425,N_18565);
nor U18781 (N_18781,N_15965,N_15343);
nand U18782 (N_18782,N_16455,N_12519);
and U18783 (N_18783,N_17770,N_18497);
or U18784 (N_18784,N_12846,N_12711);
nand U18785 (N_18785,N_18727,N_17472);
nor U18786 (N_18786,N_12770,N_18641);
xnor U18787 (N_18787,N_13055,N_17607);
or U18788 (N_18788,N_14256,N_14481);
nand U18789 (N_18789,N_18746,N_14600);
nand U18790 (N_18790,N_13353,N_15020);
nand U18791 (N_18791,N_18311,N_18427);
nand U18792 (N_18792,N_15571,N_15631);
nand U18793 (N_18793,N_13629,N_15006);
nor U18794 (N_18794,N_16649,N_14483);
and U18795 (N_18795,N_13220,N_15321);
nand U18796 (N_18796,N_14654,N_12763);
or U18797 (N_18797,N_16486,N_13019);
xnor U18798 (N_18798,N_18568,N_16532);
or U18799 (N_18799,N_15143,N_14355);
and U18800 (N_18800,N_18037,N_12629);
and U18801 (N_18801,N_15540,N_16319);
nand U18802 (N_18802,N_16797,N_14923);
nand U18803 (N_18803,N_16416,N_17020);
and U18804 (N_18804,N_13002,N_12710);
or U18805 (N_18805,N_16182,N_15713);
and U18806 (N_18806,N_14788,N_16193);
or U18807 (N_18807,N_13962,N_17002);
nand U18808 (N_18808,N_14034,N_15400);
nand U18809 (N_18809,N_14060,N_14124);
and U18810 (N_18810,N_12607,N_12616);
nand U18811 (N_18811,N_14407,N_14979);
and U18812 (N_18812,N_14327,N_18609);
nand U18813 (N_18813,N_14083,N_13065);
nand U18814 (N_18814,N_18307,N_14402);
and U18815 (N_18815,N_12919,N_14296);
nor U18816 (N_18816,N_15795,N_15801);
nand U18817 (N_18817,N_16521,N_13726);
and U18818 (N_18818,N_17049,N_18473);
or U18819 (N_18819,N_18056,N_14874);
nand U18820 (N_18820,N_16169,N_13871);
and U18821 (N_18821,N_16531,N_17756);
nor U18822 (N_18822,N_15671,N_16502);
or U18823 (N_18823,N_15236,N_16747);
and U18824 (N_18824,N_16172,N_13079);
nand U18825 (N_18825,N_14522,N_15192);
nor U18826 (N_18826,N_15374,N_14168);
xnor U18827 (N_18827,N_14532,N_17189);
nand U18828 (N_18828,N_15428,N_15656);
and U18829 (N_18829,N_13463,N_16553);
nor U18830 (N_18830,N_18580,N_17719);
nand U18831 (N_18831,N_16731,N_12996);
or U18832 (N_18832,N_15879,N_15165);
nor U18833 (N_18833,N_14291,N_15083);
and U18834 (N_18834,N_16190,N_16652);
or U18835 (N_18835,N_16039,N_16832);
nor U18836 (N_18836,N_12853,N_15270);
xnor U18837 (N_18837,N_14378,N_16736);
nand U18838 (N_18838,N_17438,N_13829);
nand U18839 (N_18839,N_15181,N_14130);
and U18840 (N_18840,N_17737,N_13550);
or U18841 (N_18841,N_16110,N_18012);
and U18842 (N_18842,N_16807,N_17644);
and U18843 (N_18843,N_14737,N_15864);
nand U18844 (N_18844,N_12554,N_16329);
nor U18845 (N_18845,N_16285,N_17199);
nand U18846 (N_18846,N_16378,N_16314);
and U18847 (N_18847,N_13540,N_14386);
or U18848 (N_18848,N_18199,N_14004);
nor U18849 (N_18849,N_15767,N_18432);
or U18850 (N_18850,N_13299,N_12799);
and U18851 (N_18851,N_14696,N_13878);
and U18852 (N_18852,N_15634,N_14539);
and U18853 (N_18853,N_13247,N_17578);
and U18854 (N_18854,N_16888,N_15919);
nand U18855 (N_18855,N_18247,N_13290);
and U18856 (N_18856,N_13012,N_13251);
or U18857 (N_18857,N_17645,N_12686);
nand U18858 (N_18858,N_13628,N_13912);
nor U18859 (N_18859,N_16070,N_13884);
and U18860 (N_18860,N_14992,N_15233);
xor U18861 (N_18861,N_15498,N_16408);
and U18862 (N_18862,N_16345,N_16130);
or U18863 (N_18863,N_18670,N_17476);
nand U18864 (N_18864,N_12917,N_12700);
and U18865 (N_18865,N_17093,N_15413);
and U18866 (N_18866,N_16419,N_13898);
or U18867 (N_18867,N_18604,N_14844);
nor U18868 (N_18868,N_16199,N_13470);
xnor U18869 (N_18869,N_16377,N_12502);
xor U18870 (N_18870,N_13911,N_13376);
nand U18871 (N_18871,N_16376,N_18531);
or U18872 (N_18872,N_18010,N_18278);
nand U18873 (N_18873,N_15222,N_17484);
or U18874 (N_18874,N_13025,N_15053);
or U18875 (N_18875,N_15203,N_17186);
xor U18876 (N_18876,N_18384,N_16372);
nand U18877 (N_18877,N_13775,N_18650);
nand U18878 (N_18878,N_16886,N_16889);
and U18879 (N_18879,N_17279,N_13496);
nor U18880 (N_18880,N_14373,N_16457);
nand U18881 (N_18881,N_18550,N_13056);
nand U18882 (N_18882,N_12913,N_18409);
nand U18883 (N_18883,N_17102,N_12960);
or U18884 (N_18884,N_14703,N_16120);
and U18885 (N_18885,N_17608,N_16655);
nor U18886 (N_18886,N_15262,N_17012);
nand U18887 (N_18887,N_16897,N_12520);
nor U18888 (N_18888,N_13246,N_13634);
nand U18889 (N_18889,N_15673,N_17326);
xnor U18890 (N_18890,N_14792,N_13607);
and U18891 (N_18891,N_18257,N_17890);
nand U18892 (N_18892,N_15966,N_13805);
and U18893 (N_18893,N_18368,N_12619);
nor U18894 (N_18894,N_14070,N_17642);
xor U18895 (N_18895,N_14872,N_18057);
nand U18896 (N_18896,N_13180,N_13320);
and U18897 (N_18897,N_18380,N_18053);
nand U18898 (N_18898,N_14825,N_16327);
nor U18899 (N_18899,N_17195,N_13851);
nor U18900 (N_18900,N_14241,N_13771);
and U18901 (N_18901,N_14415,N_16435);
and U18902 (N_18902,N_16379,N_16047);
or U18903 (N_18903,N_17925,N_15948);
nor U18904 (N_18904,N_15587,N_16992);
or U18905 (N_18905,N_17896,N_13735);
and U18906 (N_18906,N_16214,N_17084);
and U18907 (N_18907,N_14847,N_13501);
and U18908 (N_18908,N_12721,N_18073);
and U18909 (N_18909,N_16100,N_16165);
or U18910 (N_18910,N_12728,N_17822);
nand U18911 (N_18911,N_16847,N_16443);
nand U18912 (N_18912,N_12576,N_18165);
and U18913 (N_18913,N_15846,N_15486);
nand U18914 (N_18914,N_12541,N_14993);
and U18915 (N_18915,N_13439,N_18514);
or U18916 (N_18916,N_13569,N_16777);
nor U18917 (N_18917,N_17872,N_15241);
or U18918 (N_18918,N_15788,N_13314);
or U18919 (N_18919,N_12581,N_14232);
and U18920 (N_18920,N_16499,N_16800);
nor U18921 (N_18921,N_17633,N_12790);
and U18922 (N_18922,N_14469,N_17436);
nand U18923 (N_18923,N_15902,N_16890);
nand U18924 (N_18924,N_15094,N_18396);
and U18925 (N_18925,N_15900,N_14337);
nand U18926 (N_18926,N_15534,N_18120);
or U18927 (N_18927,N_13276,N_15888);
nand U18928 (N_18928,N_17912,N_13259);
nand U18929 (N_18929,N_12839,N_16151);
xor U18930 (N_18930,N_13599,N_18239);
nor U18931 (N_18931,N_12510,N_12544);
and U18932 (N_18932,N_13457,N_13092);
and U18933 (N_18933,N_14117,N_15802);
and U18934 (N_18934,N_14828,N_17169);
xnor U18935 (N_18935,N_15347,N_16615);
nand U18936 (N_18936,N_18737,N_13033);
nand U18937 (N_18937,N_17674,N_16299);
nor U18938 (N_18938,N_18435,N_18534);
or U18939 (N_18939,N_16323,N_12538);
nor U18940 (N_18940,N_16243,N_15405);
or U18941 (N_18941,N_14743,N_14326);
nand U18942 (N_18942,N_16619,N_17036);
nor U18943 (N_18943,N_17687,N_13426);
and U18944 (N_18944,N_16679,N_14331);
or U18945 (N_18945,N_17840,N_12618);
xnor U18946 (N_18946,N_15050,N_18026);
or U18947 (N_18947,N_13603,N_14854);
nor U18948 (N_18948,N_17982,N_14862);
and U18949 (N_18949,N_16031,N_16637);
nor U18950 (N_18950,N_14697,N_17944);
and U18951 (N_18951,N_12725,N_15857);
or U18952 (N_18952,N_16928,N_14182);
and U18953 (N_18953,N_15354,N_12882);
or U18954 (N_18954,N_17748,N_16137);
nor U18955 (N_18955,N_13514,N_15430);
or U18956 (N_18956,N_18044,N_15353);
or U18957 (N_18957,N_16504,N_17570);
nand U18958 (N_18958,N_16582,N_17244);
nor U18959 (N_18959,N_12673,N_13799);
or U18960 (N_18960,N_17576,N_14271);
nand U18961 (N_18961,N_13355,N_16571);
and U18962 (N_18962,N_13380,N_18455);
xor U18963 (N_18963,N_17182,N_12946);
nand U18964 (N_18964,N_16469,N_13989);
xnor U18965 (N_18965,N_14592,N_16411);
or U18966 (N_18966,N_16648,N_16595);
nand U18967 (N_18967,N_16093,N_17345);
and U18968 (N_18968,N_13466,N_17233);
or U18969 (N_18969,N_14986,N_16335);
nor U18970 (N_18970,N_18575,N_16585);
nor U18971 (N_18971,N_14203,N_12636);
or U18972 (N_18972,N_13758,N_15359);
nand U18973 (N_18973,N_14863,N_14112);
nand U18974 (N_18974,N_16870,N_17395);
and U18975 (N_18975,N_12676,N_14651);
or U18976 (N_18976,N_13512,N_12614);
or U18977 (N_18977,N_13167,N_13529);
and U18978 (N_18978,N_13297,N_13631);
and U18979 (N_18979,N_15492,N_18137);
nor U18980 (N_18980,N_14739,N_15377);
xor U18981 (N_18981,N_13233,N_16694);
or U18982 (N_18982,N_13316,N_12995);
or U18983 (N_18983,N_18365,N_13235);
xnor U18984 (N_18984,N_14736,N_16248);
and U18985 (N_18985,N_17118,N_14621);
nor U18986 (N_18986,N_17902,N_14582);
nand U18987 (N_18987,N_12757,N_16393);
or U18988 (N_18988,N_14972,N_16467);
and U18989 (N_18989,N_12716,N_16882);
nor U18990 (N_18990,N_18089,N_15519);
nor U18991 (N_18991,N_13844,N_13972);
nor U18992 (N_18992,N_13654,N_16186);
nor U18993 (N_18993,N_14280,N_16105);
nor U18994 (N_18994,N_16007,N_17755);
nand U18995 (N_18995,N_16829,N_18009);
or U18996 (N_18996,N_14694,N_18379);
or U18997 (N_18997,N_14642,N_17273);
and U18998 (N_18998,N_13563,N_13018);
and U18999 (N_18999,N_15309,N_14200);
nor U19000 (N_19000,N_12517,N_18251);
or U19001 (N_19001,N_14687,N_18036);
and U19002 (N_19002,N_13123,N_15843);
nor U19003 (N_19003,N_16140,N_17723);
xor U19004 (N_19004,N_12971,N_18147);
nand U19005 (N_19005,N_14850,N_16758);
and U19006 (N_19006,N_18262,N_13876);
nand U19007 (N_19007,N_18295,N_17292);
or U19008 (N_19008,N_13286,N_17649);
nand U19009 (N_19009,N_16333,N_12966);
nand U19010 (N_19010,N_15162,N_17620);
or U19011 (N_19011,N_16177,N_17104);
or U19012 (N_19012,N_15939,N_15676);
xor U19013 (N_19013,N_18213,N_18242);
nand U19014 (N_19014,N_14523,N_16576);
or U19015 (N_19015,N_16464,N_14823);
and U19016 (N_19016,N_13717,N_17843);
or U19017 (N_19017,N_13084,N_17260);
nand U19018 (N_19018,N_15330,N_14977);
nor U19019 (N_19019,N_14812,N_15903);
or U19020 (N_19020,N_18013,N_15060);
nor U19021 (N_19021,N_13539,N_17775);
nor U19022 (N_19022,N_14753,N_12833);
nand U19023 (N_19023,N_12901,N_17178);
or U19024 (N_19024,N_16880,N_16164);
nand U19025 (N_19025,N_17482,N_14510);
xor U19026 (N_19026,N_17803,N_18709);
or U19027 (N_19027,N_15528,N_16304);
and U19028 (N_19028,N_14930,N_15882);
nand U19029 (N_19029,N_14136,N_16363);
or U19030 (N_19030,N_14251,N_16250);
nand U19031 (N_19031,N_14145,N_14772);
and U19032 (N_19032,N_17540,N_14842);
or U19033 (N_19033,N_15011,N_14606);
nor U19034 (N_19034,N_13298,N_18339);
nand U19035 (N_19035,N_13659,N_13900);
and U19036 (N_19036,N_15010,N_13986);
nor U19037 (N_19037,N_17796,N_16078);
or U19038 (N_19038,N_14486,N_12747);
or U19039 (N_19039,N_15117,N_16854);
and U19040 (N_19040,N_16723,N_15169);
and U19041 (N_19041,N_13778,N_18264);
and U19042 (N_19042,N_14775,N_16071);
nand U19043 (N_19043,N_13567,N_18639);
or U19044 (N_19044,N_13728,N_13164);
nand U19045 (N_19045,N_17252,N_12948);
nand U19046 (N_19046,N_18449,N_14127);
xnor U19047 (N_19047,N_13451,N_17485);
and U19048 (N_19048,N_12564,N_18499);
nor U19049 (N_19049,N_17416,N_14660);
or U19050 (N_19050,N_12631,N_12767);
nand U19051 (N_19051,N_13780,N_17010);
xor U19052 (N_19052,N_15581,N_18285);
and U19053 (N_19053,N_14673,N_15189);
or U19054 (N_19054,N_16505,N_18170);
or U19055 (N_19055,N_14829,N_18025);
and U19056 (N_19056,N_14951,N_17605);
and U19057 (N_19057,N_15810,N_17823);
or U19058 (N_19058,N_15123,N_15373);
or U19059 (N_19059,N_17079,N_14875);
or U19060 (N_19060,N_16225,N_17746);
nand U19061 (N_19061,N_14032,N_13330);
nand U19062 (N_19062,N_13042,N_15462);
nor U19063 (N_19063,N_16357,N_18007);
nand U19064 (N_19064,N_13379,N_18335);
or U19065 (N_19065,N_18500,N_15926);
and U19066 (N_19066,N_18667,N_16032);
nor U19067 (N_19067,N_18674,N_18062);
xnor U19068 (N_19068,N_18019,N_16642);
xor U19069 (N_19069,N_18530,N_16428);
and U19070 (N_19070,N_17710,N_16772);
nor U19071 (N_19071,N_14221,N_15897);
or U19072 (N_19072,N_16675,N_17015);
xnor U19073 (N_19073,N_15745,N_17088);
and U19074 (N_19074,N_12969,N_16010);
xnor U19075 (N_19075,N_17954,N_14672);
and U19076 (N_19076,N_16347,N_13504);
nor U19077 (N_19077,N_17977,N_15761);
and U19078 (N_19078,N_17489,N_16445);
or U19079 (N_19079,N_15455,N_16312);
nand U19080 (N_19080,N_17707,N_16232);
and U19081 (N_19081,N_14681,N_13337);
nor U19082 (N_19082,N_16485,N_18687);
or U19083 (N_19083,N_14547,N_13255);
and U19084 (N_19084,N_14234,N_18112);
nand U19085 (N_19085,N_18061,N_17386);
or U19086 (N_19086,N_16001,N_14458);
nor U19087 (N_19087,N_12678,N_12912);
or U19088 (N_19088,N_14509,N_16906);
nand U19089 (N_19089,N_18517,N_13060);
and U19090 (N_19090,N_15255,N_17767);
nor U19091 (N_19091,N_12536,N_15829);
or U19092 (N_19092,N_15063,N_13578);
and U19093 (N_19093,N_17166,N_14466);
nand U19094 (N_19094,N_13135,N_17711);
nor U19095 (N_19095,N_15837,N_12718);
xnor U19096 (N_19096,N_14639,N_12847);
nand U19097 (N_19097,N_16995,N_13821);
or U19098 (N_19098,N_13214,N_18128);
xor U19099 (N_19099,N_14525,N_18352);
nor U19100 (N_19100,N_15204,N_16222);
or U19101 (N_19101,N_18028,N_13681);
nor U19102 (N_19102,N_14099,N_13273);
nor U19103 (N_19103,N_16688,N_18282);
nor U19104 (N_19104,N_12652,N_13190);
nand U19105 (N_19105,N_13336,N_12598);
or U19106 (N_19106,N_16076,N_14389);
nand U19107 (N_19107,N_17883,N_14383);
and U19108 (N_19108,N_15844,N_16274);
or U19109 (N_19109,N_16835,N_16160);
or U19110 (N_19110,N_12923,N_17636);
nand U19111 (N_19111,N_16566,N_15084);
or U19112 (N_19112,N_15487,N_16048);
xor U19113 (N_19113,N_12865,N_17602);
and U19114 (N_19114,N_17493,N_18211);
or U19115 (N_19115,N_18031,N_17231);
nor U19116 (N_19116,N_17018,N_13108);
nor U19117 (N_19117,N_14158,N_16894);
or U19118 (N_19118,N_15834,N_15397);
nand U19119 (N_19119,N_17750,N_16237);
and U19120 (N_19120,N_14243,N_13346);
nand U19121 (N_19121,N_18344,N_13306);
nand U19122 (N_19122,N_17574,N_17417);
and U19123 (N_19123,N_14003,N_14713);
nor U19124 (N_19124,N_16872,N_13248);
nand U19125 (N_19125,N_14196,N_17217);
nor U19126 (N_19126,N_13444,N_17911);
nand U19127 (N_19127,N_15424,N_17647);
xor U19128 (N_19128,N_13809,N_16440);
nand U19129 (N_19129,N_17851,N_15022);
xor U19130 (N_19130,N_14170,N_13095);
nor U19131 (N_19131,N_16828,N_16982);
xor U19132 (N_19132,N_13267,N_15558);
or U19133 (N_19133,N_13687,N_18317);
or U19134 (N_19134,N_16706,N_12620);
nand U19135 (N_19135,N_15366,N_17390);
or U19136 (N_19136,N_12526,N_16359);
nand U19137 (N_19137,N_14485,N_14889);
nor U19138 (N_19138,N_17383,N_16107);
or U19139 (N_19139,N_15877,N_15536);
nand U19140 (N_19140,N_13016,N_14033);
nor U19141 (N_19141,N_16593,N_15614);
nor U19142 (N_19142,N_14315,N_14643);
and U19143 (N_19143,N_13342,N_13090);
or U19144 (N_19144,N_13264,N_15307);
and U19145 (N_19145,N_14177,N_13899);
nor U19146 (N_19146,N_13595,N_18040);
or U19147 (N_19147,N_17044,N_17011);
nand U19148 (N_19148,N_13043,N_16238);
nand U19149 (N_19149,N_17130,N_17192);
nor U19150 (N_19150,N_15098,N_18214);
nor U19151 (N_19151,N_14092,N_12759);
xor U19152 (N_19152,N_16824,N_13305);
nor U19153 (N_19153,N_18728,N_16041);
or U19154 (N_19154,N_16900,N_16602);
or U19155 (N_19155,N_15790,N_14341);
or U19156 (N_19156,N_17094,N_13404);
or U19157 (N_19157,N_15727,N_18561);
nor U19158 (N_19158,N_17239,N_17511);
nand U19159 (N_19159,N_16407,N_12706);
nor U19160 (N_19160,N_14143,N_12892);
and U19161 (N_19161,N_17487,N_18720);
and U19162 (N_19162,N_15086,N_14226);
and U19163 (N_19163,N_13335,N_18627);
nand U19164 (N_19164,N_13490,N_14231);
nand U19165 (N_19165,N_17632,N_17222);
xnor U19166 (N_19166,N_17988,N_12845);
nand U19167 (N_19167,N_16420,N_17028);
or U19168 (N_19168,N_16014,N_14279);
or U19169 (N_19169,N_13966,N_17156);
and U19170 (N_19170,N_17060,N_13614);
nand U19171 (N_19171,N_17396,N_18634);
nor U19172 (N_19172,N_15819,N_17995);
nand U19173 (N_19173,N_16068,N_15282);
nor U19174 (N_19174,N_14169,N_15346);
or U19175 (N_19175,N_12848,N_17308);
nor U19176 (N_19176,N_12965,N_14785);
nand U19177 (N_19177,N_16430,N_17136);
and U19178 (N_19178,N_16611,N_17564);
or U19179 (N_19179,N_16399,N_17786);
xor U19180 (N_19180,N_17779,N_15543);
nor U19181 (N_19181,N_15744,N_12730);
and U19182 (N_19182,N_18571,N_13324);
nand U19183 (N_19183,N_13369,N_17221);
and U19184 (N_19184,N_18260,N_13410);
xor U19185 (N_19185,N_12659,N_12881);
and U19186 (N_19186,N_17040,N_16843);
nand U19187 (N_19187,N_14504,N_13423);
nor U19188 (N_19188,N_18412,N_13644);
and U19189 (N_19189,N_16415,N_14885);
or U19190 (N_19190,N_13484,N_12866);
and U19191 (N_19191,N_13205,N_14649);
or U19192 (N_19192,N_18274,N_18419);
xnor U19193 (N_19193,N_16227,N_16353);
nor U19194 (N_19194,N_14095,N_16875);
nor U19195 (N_19195,N_16311,N_12774);
and U19196 (N_19196,N_16691,N_16301);
or U19197 (N_19197,N_14815,N_15751);
xnor U19198 (N_19198,N_15797,N_16862);
and U19199 (N_19199,N_15408,N_17834);
and U19200 (N_19200,N_16919,N_12590);
nor U19201 (N_19201,N_13474,N_18614);
nand U19202 (N_19202,N_12726,N_13702);
xor U19203 (N_19203,N_18310,N_13440);
nand U19204 (N_19204,N_12990,N_18281);
nand U19205 (N_19205,N_13743,N_14058);
xnor U19206 (N_19206,N_14856,N_16577);
nor U19207 (N_19207,N_16544,N_13250);
nor U19208 (N_19208,N_14173,N_13842);
nand U19209 (N_19209,N_12695,N_17149);
and U19210 (N_19210,N_12754,N_14559);
and U19211 (N_19211,N_15247,N_16475);
and U19212 (N_19212,N_13497,N_15707);
or U19213 (N_19213,N_15848,N_15785);
and U19214 (N_19214,N_15650,N_14988);
nor U19215 (N_19215,N_16432,N_18722);
nand U19216 (N_19216,N_13458,N_18498);
xnor U19217 (N_19217,N_15816,N_16173);
nand U19218 (N_19218,N_16664,N_14542);
or U19219 (N_19219,N_13333,N_13288);
or U19220 (N_19220,N_16871,N_18284);
nor U19221 (N_19221,N_15973,N_13610);
nor U19222 (N_19222,N_17857,N_15970);
and U19223 (N_19223,N_15317,N_12994);
nand U19224 (N_19224,N_13015,N_14354);
nor U19225 (N_19225,N_17521,N_18315);
and U19226 (N_19226,N_15553,N_15960);
or U19227 (N_19227,N_17754,N_13059);
and U19228 (N_19228,N_12569,N_18607);
and U19229 (N_19229,N_16119,N_15786);
nor U19230 (N_19230,N_17116,N_13063);
nor U19231 (N_19231,N_14098,N_12602);
nand U19232 (N_19232,N_16251,N_13481);
nand U19233 (N_19233,N_17979,N_18038);
nand U19234 (N_19234,N_13910,N_16195);
nor U19235 (N_19235,N_16258,N_15033);
nand U19236 (N_19236,N_13922,N_13198);
nand U19237 (N_19237,N_13798,N_14462);
or U19238 (N_19238,N_14357,N_12683);
nand U19239 (N_19239,N_13894,N_18093);
nand U19240 (N_19240,N_18731,N_13000);
and U19241 (N_19241,N_18657,N_16136);
nand U19242 (N_19242,N_14608,N_17641);
or U19243 (N_19243,N_16861,N_18489);
or U19244 (N_19244,N_16984,N_14190);
nand U19245 (N_19245,N_16022,N_18027);
and U19246 (N_19246,N_18668,N_18182);
or U19247 (N_19247,N_18480,N_17391);
nand U19248 (N_19248,N_13737,N_14768);
xnor U19249 (N_19249,N_17837,N_14056);
or U19250 (N_19250,N_14831,N_14472);
or U19251 (N_19251,N_13206,N_16059);
xnor U19252 (N_19252,N_14517,N_16074);
nor U19253 (N_19253,N_16262,N_16210);
or U19254 (N_19254,N_13516,N_17604);
nor U19255 (N_19255,N_12822,N_15286);
nand U19256 (N_19256,N_15590,N_16686);
or U19257 (N_19257,N_16384,N_14370);
and U19258 (N_19258,N_16033,N_13118);
nor U19259 (N_19259,N_13905,N_13925);
xnor U19260 (N_19260,N_15231,N_15694);
and U19261 (N_19261,N_17513,N_13408);
and U19262 (N_19262,N_15308,N_15196);
and U19263 (N_19263,N_15398,N_13772);
or U19264 (N_19264,N_17866,N_12670);
or U19265 (N_19265,N_14916,N_14162);
or U19266 (N_19266,N_16109,N_12762);
and U19267 (N_19267,N_12583,N_13616);
nor U19268 (N_19268,N_15439,N_17867);
nand U19269 (N_19269,N_16236,N_15578);
nor U19270 (N_19270,N_15260,N_16855);
or U19271 (N_19271,N_18159,N_18421);
or U19272 (N_19272,N_16020,N_17278);
nand U19273 (N_19273,N_15009,N_14771);
or U19274 (N_19274,N_15135,N_18689);
or U19275 (N_19275,N_18741,N_16484);
xor U19276 (N_19276,N_14922,N_17683);
xor U19277 (N_19277,N_15139,N_14894);
nor U19278 (N_19278,N_17583,N_14019);
xor U19279 (N_19279,N_17677,N_14715);
xor U19280 (N_19280,N_16337,N_15474);
nand U19281 (N_19281,N_15160,N_17606);
xor U19282 (N_19282,N_14108,N_17421);
and U19283 (N_19283,N_15026,N_15470);
nand U19284 (N_19284,N_15187,N_16623);
xor U19285 (N_19285,N_13176,N_17590);
nand U19286 (N_19286,N_16293,N_15344);
xnor U19287 (N_19287,N_13833,N_15429);
nor U19288 (N_19288,N_15557,N_16218);
nand U19289 (N_19289,N_13764,N_12751);
or U19290 (N_19290,N_14300,N_16999);
nand U19291 (N_19291,N_18393,N_13725);
nor U19292 (N_19292,N_18426,N_14845);
and U19293 (N_19293,N_14943,N_15716);
or U19294 (N_19294,N_18744,N_14489);
nand U19295 (N_19295,N_15597,N_14167);
nand U19296 (N_19296,N_16303,N_13104);
and U19297 (N_19297,N_12938,N_15747);
nand U19298 (N_19298,N_15318,N_15440);
or U19299 (N_19299,N_18154,N_13340);
nand U19300 (N_19300,N_12858,N_15272);
nand U19301 (N_19301,N_16755,N_15288);
xnor U19302 (N_19302,N_16034,N_13249);
or U19303 (N_19303,N_17628,N_14433);
xor U19304 (N_19304,N_13178,N_18646);
and U19305 (N_19305,N_16352,N_13525);
or U19306 (N_19306,N_14290,N_16763);
nor U19307 (N_19307,N_15770,N_13582);
nand U19308 (N_19308,N_18321,N_15618);
or U19309 (N_19309,N_15494,N_17942);
or U19310 (N_19310,N_16196,N_14858);
or U19311 (N_19311,N_14309,N_18133);
nand U19312 (N_19312,N_15212,N_16744);
or U19313 (N_19313,N_13593,N_13543);
nand U19314 (N_19314,N_13881,N_17893);
xnor U19315 (N_19315,N_17716,N_17885);
or U19316 (N_19316,N_16148,N_16698);
xor U19317 (N_19317,N_15205,N_18527);
or U19318 (N_19318,N_15001,N_13327);
or U19319 (N_19319,N_13957,N_13262);
nand U19320 (N_19320,N_13836,N_14135);
nand U19321 (N_19321,N_15443,N_17125);
and U19322 (N_19322,N_17934,N_16460);
or U19323 (N_19323,N_14554,N_17753);
nor U19324 (N_19324,N_14938,N_16525);
nor U19325 (N_19325,N_13742,N_15525);
and U19326 (N_19326,N_13933,N_15754);
nand U19327 (N_19327,N_14461,N_18475);
or U19328 (N_19328,N_14583,N_18659);
and U19329 (N_19329,N_17845,N_14852);
nand U19330 (N_19330,N_13338,N_12680);
nand U19331 (N_19331,N_16121,N_14959);
and U19332 (N_19332,N_15721,N_15945);
nand U19333 (N_19333,N_14456,N_18210);
xor U19334 (N_19334,N_17077,N_17939);
nand U19335 (N_19335,N_14543,N_15870);
or U19336 (N_19336,N_16398,N_18601);
nand U19337 (N_19337,N_18079,N_15000);
or U19338 (N_19338,N_14375,N_15103);
or U19339 (N_19339,N_18444,N_14619);
or U19340 (N_19340,N_17996,N_13506);
and U19341 (N_19341,N_16771,N_17200);
nand U19342 (N_19342,N_14482,N_14808);
xor U19343 (N_19343,N_13801,N_16437);
and U19344 (N_19344,N_13621,N_15549);
nand U19345 (N_19345,N_14371,N_17847);
nor U19346 (N_19346,N_17013,N_18395);
nand U19347 (N_19347,N_13661,N_14896);
xnor U19348 (N_19348,N_14799,N_13396);
nor U19349 (N_19349,N_15602,N_16656);
nor U19350 (N_19350,N_12795,N_18416);
nor U19351 (N_19351,N_16673,N_15736);
or U19352 (N_19352,N_17054,N_16780);
and U19353 (N_19353,N_16156,N_14069);
nor U19354 (N_19354,N_17005,N_18191);
and U19355 (N_19355,N_15048,N_14778);
nor U19356 (N_19356,N_15106,N_13994);
or U19357 (N_19357,N_13027,N_16994);
or U19358 (N_19358,N_18370,N_17071);
nor U19359 (N_19359,N_15244,N_17235);
nor U19360 (N_19360,N_17807,N_17863);
or U19361 (N_19361,N_12653,N_13706);
nand U19362 (N_19362,N_18174,N_18739);
or U19363 (N_19363,N_16268,N_13908);
or U19364 (N_19364,N_14460,N_13400);
or U19365 (N_19365,N_14857,N_18129);
nand U19366 (N_19366,N_13215,N_14683);
or U19367 (N_19367,N_13532,N_13106);
nor U19368 (N_19368,N_15221,N_17805);
nor U19369 (N_19369,N_12875,N_17219);
nor U19370 (N_19370,N_14635,N_16295);
nand U19371 (N_19371,N_15800,N_13162);
and U19372 (N_19372,N_18710,N_17547);
or U19373 (N_19373,N_15722,N_18467);
and U19374 (N_19374,N_14319,N_18020);
nand U19375 (N_19375,N_14962,N_14429);
xnor U19376 (N_19376,N_18114,N_12900);
and U19377 (N_19377,N_12985,N_18726);
and U19378 (N_19378,N_17500,N_15137);
nand U19379 (N_19379,N_13173,N_16027);
or U19380 (N_19380,N_13417,N_14627);
or U19381 (N_19381,N_14949,N_15659);
xor U19382 (N_19382,N_15168,N_14833);
and U19383 (N_19383,N_13843,N_13151);
or U19384 (N_19384,N_16123,N_13590);
and U19385 (N_19385,N_15274,N_15174);
and U19386 (N_19386,N_18567,N_15559);
or U19387 (N_19387,N_14134,N_17989);
and U19388 (N_19388,N_14605,N_13760);
xor U19389 (N_19389,N_13787,N_17133);
nor U19390 (N_19390,N_17281,N_14780);
nand U19391 (N_19391,N_15193,N_16725);
nor U19392 (N_19392,N_14237,N_17120);
xnor U19393 (N_19393,N_13662,N_13573);
and U19394 (N_19394,N_15544,N_15393);
and U19395 (N_19395,N_14822,N_15434);
and U19396 (N_19396,N_14645,N_16436);
nor U19397 (N_19397,N_18654,N_14950);
xnor U19398 (N_19398,N_12814,N_16804);
or U19399 (N_19399,N_17778,N_13145);
and U19400 (N_19400,N_15718,N_17266);
xnor U19401 (N_19401,N_14081,N_13152);
nor U19402 (N_19402,N_17978,N_17289);
nand U19403 (N_19403,N_13099,N_14185);
nand U19404 (N_19404,N_17594,N_13868);
nor U19405 (N_19405,N_13102,N_15155);
and U19406 (N_19406,N_13186,N_14041);
or U19407 (N_19407,N_15279,N_17975);
or U19408 (N_19408,N_17469,N_12920);
nor U19409 (N_19409,N_14029,N_13546);
nor U19410 (N_19410,N_17567,N_14811);
nand U19411 (N_19411,N_14154,N_16406);
xnor U19412 (N_19412,N_14484,N_15369);
nand U19413 (N_19413,N_14416,N_16966);
nand U19414 (N_19414,N_18616,N_17337);
or U19415 (N_19415,N_15641,N_17019);
and U19416 (N_19416,N_13988,N_14116);
and U19417 (N_19417,N_14216,N_16106);
nand U19418 (N_19418,N_15677,N_18006);
and U19419 (N_19419,N_13604,N_16760);
and U19420 (N_19420,N_12723,N_17410);
or U19421 (N_19421,N_14920,N_12964);
nand U19422 (N_19422,N_15904,N_17201);
and U19423 (N_19423,N_15969,N_16356);
and U19424 (N_19424,N_14946,N_16645);
or U19425 (N_19425,N_18067,N_14001);
or U19426 (N_19426,N_15059,N_14146);
xnor U19427 (N_19427,N_17413,N_13973);
nand U19428 (N_19428,N_15732,N_14115);
nand U19429 (N_19429,N_13656,N_15737);
or U19430 (N_19430,N_14679,N_16364);
nor U19431 (N_19431,N_14320,N_15396);
nand U19432 (N_19432,N_17399,N_18542);
or U19433 (N_19433,N_14316,N_16969);
and U19434 (N_19434,N_17232,N_17408);
and U19435 (N_19435,N_13011,N_17665);
and U19436 (N_19436,N_13195,N_12733);
nor U19437 (N_19437,N_17332,N_13425);
and U19438 (N_19438,N_15703,N_18502);
xor U19439 (N_19439,N_13997,N_13307);
nand U19440 (N_19440,N_16592,N_16003);
nand U19441 (N_19441,N_12760,N_18386);
nor U19442 (N_19442,N_15922,N_13916);
and U19443 (N_19443,N_15365,N_17196);
and U19444 (N_19444,N_16069,N_13549);
nor U19445 (N_19445,N_12931,N_17241);
nor U19446 (N_19446,N_15488,N_14101);
nor U19447 (N_19447,N_16371,N_12738);
nand U19448 (N_19448,N_16242,N_17021);
or U19449 (N_19449,N_18748,N_15824);
xnor U19450 (N_19450,N_16546,N_16957);
xnor U19451 (N_19451,N_16189,N_18729);
and U19452 (N_19452,N_15031,N_15665);
nand U19453 (N_19453,N_16503,N_18101);
or U19454 (N_19454,N_18385,N_15858);
nand U19455 (N_19455,N_13975,N_16178);
xnor U19456 (N_19456,N_14641,N_14045);
nand U19457 (N_19457,N_18458,N_14594);
xnor U19458 (N_19458,N_16491,N_15437);
and U19459 (N_19459,N_15018,N_15866);
nor U19460 (N_19460,N_12951,N_14376);
nor U19461 (N_19461,N_17446,N_16550);
or U19462 (N_19462,N_12891,N_14562);
nand U19463 (N_19463,N_13660,N_14107);
or U19464 (N_19464,N_17791,N_13397);
nand U19465 (N_19465,N_18183,N_17349);
nor U19466 (N_19466,N_13535,N_17941);
nand U19467 (N_19467,N_12842,N_13429);
nand U19468 (N_19468,N_15526,N_13153);
or U19469 (N_19469,N_15225,N_17833);
nor U19470 (N_19470,N_14334,N_16497);
nand U19471 (N_19471,N_12769,N_16476);
xnor U19472 (N_19472,N_18000,N_18232);
and U19473 (N_19473,N_16588,N_16851);
nor U19474 (N_19474,N_15450,N_15899);
nand U19475 (N_19475,N_14188,N_13472);
nor U19476 (N_19476,N_13740,N_13638);
or U19477 (N_19477,N_18619,N_15931);
nor U19478 (N_19478,N_13392,N_15297);
nor U19479 (N_19479,N_15340,N_17257);
xor U19480 (N_19480,N_18623,N_18597);
nor U19481 (N_19481,N_16930,N_17087);
nand U19482 (N_19482,N_14411,N_14071);
and U19483 (N_19483,N_18576,N_18066);
or U19484 (N_19484,N_13537,N_12883);
and U19485 (N_19485,N_18513,N_15072);
nand U19486 (N_19486,N_18536,N_17155);
and U19487 (N_19487,N_12955,N_18322);
nand U19488 (N_19488,N_16492,N_15503);
nand U19489 (N_19489,N_15489,N_13671);
and U19490 (N_19490,N_17198,N_14287);
nor U19491 (N_19491,N_12679,N_15218);
nand U19492 (N_19492,N_18190,N_15314);
or U19493 (N_19493,N_13360,N_18621);
or U19494 (N_19494,N_14018,N_18496);
and U19495 (N_19495,N_17690,N_17214);
and U19496 (N_19496,N_14878,N_17347);
or U19497 (N_19497,N_15932,N_16741);
or U19498 (N_19498,N_14749,N_13029);
nor U19499 (N_19499,N_14613,N_13160);
xor U19500 (N_19500,N_16768,N_14050);
nor U19501 (N_19501,N_13802,N_17427);
nand U19502 (N_19502,N_14571,N_15672);
nor U19503 (N_19503,N_16188,N_12840);
or U19504 (N_19504,N_15132,N_15976);
nor U19505 (N_19505,N_17717,N_15166);
or U19506 (N_19506,N_15892,N_16960);
nor U19507 (N_19507,N_14078,N_15772);
and U19508 (N_19508,N_15868,N_17855);
and U19509 (N_19509,N_14091,N_15159);
xnor U19510 (N_19510,N_15425,N_17901);
and U19511 (N_19511,N_18070,N_15108);
nand U19512 (N_19512,N_15925,N_12890);
or U19513 (N_19513,N_16471,N_15402);
nand U19514 (N_19514,N_13479,N_14339);
and U19515 (N_19515,N_18258,N_18539);
nor U19516 (N_19516,N_18745,N_13144);
nor U19517 (N_19517,N_15076,N_13804);
nand U19518 (N_19518,N_12504,N_14423);
nand U19519 (N_19519,N_14421,N_15871);
xnor U19520 (N_19520,N_17370,N_13865);
nand U19521 (N_19521,N_18685,N_13890);
or U19522 (N_19522,N_12761,N_17323);
and U19523 (N_19523,N_12688,N_17426);
and U19524 (N_19524,N_18336,N_15957);
xor U19525 (N_19525,N_16678,N_15841);
or U19526 (N_19526,N_16159,N_17918);
nand U19527 (N_19527,N_13332,N_17542);
and U19528 (N_19528,N_13154,N_16831);
nor U19529 (N_19529,N_16819,N_12756);
and U19530 (N_19530,N_16903,N_17573);
nand U19531 (N_19531,N_14549,N_17132);
or U19532 (N_19532,N_17110,N_18329);
and U19533 (N_19533,N_16836,N_15130);
and U19534 (N_19534,N_15860,N_18347);
or U19535 (N_19535,N_13284,N_13968);
xor U19536 (N_19536,N_17841,N_18390);
and U19537 (N_19537,N_16088,N_17204);
xnor U19538 (N_19538,N_15943,N_18446);
and U19539 (N_19539,N_13244,N_16448);
nand U19540 (N_19540,N_18606,N_17693);
and U19541 (N_19541,N_17218,N_12863);
xor U19542 (N_19542,N_16629,N_16454);
nor U19543 (N_19543,N_17220,N_15720);
or U19544 (N_19544,N_18562,N_17529);
or U19545 (N_19545,N_18389,N_18372);
xor U19546 (N_19546,N_14358,N_13503);
xnor U19547 (N_19547,N_13577,N_17137);
nand U19548 (N_19548,N_14026,N_14012);
or U19549 (N_19549,N_12609,N_14427);
or U19550 (N_19550,N_13896,N_14106);
and U19551 (N_19551,N_15110,N_14282);
or U19552 (N_19552,N_14211,N_16810);
and U19553 (N_19553,N_13230,N_12950);
and U19554 (N_19554,N_15420,N_17355);
and U19555 (N_19555,N_18050,N_13105);
nor U19556 (N_19556,N_13432,N_12798);
nand U19557 (N_19557,N_15074,N_17443);
and U19558 (N_19558,N_15234,N_18680);
nor U19559 (N_19559,N_16118,N_14385);
nor U19560 (N_19560,N_13931,N_13381);
and U19561 (N_19561,N_13793,N_18695);
xor U19562 (N_19562,N_16885,N_14392);
or U19563 (N_19563,N_13932,N_13762);
or U19564 (N_19564,N_17948,N_12930);
nand U19565 (N_19565,N_14400,N_12888);
nand U19566 (N_19566,N_14622,N_13623);
nand U19567 (N_19567,N_16235,N_15764);
or U19568 (N_19568,N_16842,N_16163);
or U19569 (N_19569,N_17634,N_18660);
or U19570 (N_19570,N_13915,N_15438);
and U19571 (N_19571,N_13731,N_13271);
or U19572 (N_19572,N_12647,N_14978);
or U19573 (N_19573,N_17935,N_18206);
and U19574 (N_19574,N_14834,N_15523);
and U19575 (N_19575,N_15651,N_17378);
xor U19576 (N_19576,N_12864,N_12784);
or U19577 (N_19577,N_17924,N_17291);
nor U19578 (N_19578,N_13182,N_16246);
nor U19579 (N_19579,N_17330,N_12874);
or U19580 (N_19580,N_16524,N_14747);
or U19581 (N_19581,N_17830,N_17735);
nor U19582 (N_19582,N_16480,N_16680);
xor U19583 (N_19583,N_16203,N_15457);
nand U19584 (N_19584,N_14928,N_12734);
or U19585 (N_19585,N_18333,N_13707);
nor U19586 (N_19586,N_13375,N_13570);
or U19587 (N_19587,N_17017,N_13129);
nand U19588 (N_19588,N_16180,N_17296);
nand U19589 (N_19589,N_12722,N_13611);
and U19590 (N_19590,N_13010,N_17029);
nor U19591 (N_19591,N_16300,N_16891);
nand U19592 (N_19592,N_17234,N_16887);
nor U19593 (N_19593,N_17304,N_16724);
and U19594 (N_19594,N_16072,N_14965);
or U19595 (N_19595,N_17790,N_15748);
nand U19596 (N_19596,N_13863,N_13938);
nand U19597 (N_19597,N_14565,N_18195);
nand U19598 (N_19598,N_13103,N_14960);
nor U19599 (N_19599,N_15603,N_17862);
nand U19600 (N_19600,N_14157,N_17471);
nor U19601 (N_19601,N_16143,N_17223);
and U19602 (N_19602,N_17887,N_14690);
nand U19603 (N_19603,N_17630,N_15327);
nor U19604 (N_19604,N_12635,N_16520);
or U19605 (N_19605,N_16738,N_16219);
and U19606 (N_19606,N_14496,N_14031);
or U19607 (N_19607,N_12775,N_18021);
nand U19608 (N_19608,N_16634,N_15004);
or U19609 (N_19609,N_14272,N_16877);
or U19610 (N_19610,N_16098,N_14556);
or U19611 (N_19611,N_17026,N_13642);
xnor U19612 (N_19612,N_16316,N_14848);
or U19613 (N_19613,N_14364,N_17303);
nand U19614 (N_19614,N_14105,N_13296);
and U19615 (N_19615,N_12530,N_15035);
or U19616 (N_19616,N_12608,N_15851);
or U19617 (N_19617,N_18243,N_17092);
nand U19618 (N_19618,N_16462,N_14588);
or U19619 (N_19619,N_17385,N_13482);
and U19620 (N_19620,N_17881,N_15555);
and U19621 (N_19621,N_17215,N_15728);
nor U19622 (N_19622,N_17302,N_15539);
or U19623 (N_19623,N_17468,N_14658);
or U19624 (N_19624,N_18361,N_13028);
nor U19625 (N_19625,N_15541,N_16456);
and U19626 (N_19626,N_16976,N_15556);
or U19627 (N_19627,N_16087,N_15312);
and U19628 (N_19628,N_15152,N_16548);
nand U19629 (N_19629,N_15652,N_17525);
nor U19630 (N_19630,N_15401,N_18624);
nand U19631 (N_19631,N_17256,N_18292);
nor U19632 (N_19632,N_17638,N_17148);
or U19633 (N_19633,N_13137,N_17366);
nand U19634 (N_19634,N_12694,N_18589);
xor U19635 (N_19635,N_16719,N_14294);
nor U19636 (N_19636,N_18742,N_14269);
nor U19637 (N_19637,N_18591,N_16988);
nor U19638 (N_19638,N_14728,N_17384);
nand U19639 (N_19639,N_15537,N_15980);
and U19640 (N_19640,N_15497,N_16641);
nand U19641 (N_19641,N_15423,N_13995);
nor U19642 (N_19642,N_18343,N_12899);
nor U19643 (N_19643,N_15202,N_18564);
or U19644 (N_19644,N_15276,N_13350);
or U19645 (N_19645,N_16095,N_17139);
and U19646 (N_19646,N_15512,N_12560);
and U19647 (N_19647,N_16948,N_17549);
xor U19648 (N_19648,N_16449,N_15092);
nand U19649 (N_19649,N_16253,N_15500);
nand U19650 (N_19650,N_15759,N_14935);
nand U19651 (N_19651,N_15830,N_15596);
or U19652 (N_19652,N_14830,N_16803);
and U19653 (N_19653,N_14035,N_18354);
and U19654 (N_19654,N_16614,N_18673);
and U19655 (N_19655,N_13174,N_14680);
nand U19656 (N_19656,N_13617,N_12982);
nor U19657 (N_19657,N_12924,N_17501);
or U19658 (N_19658,N_13581,N_16918);
xor U19659 (N_19659,N_13403,N_14498);
nor U19660 (N_19660,N_18192,N_18507);
or U19661 (N_19661,N_14214,N_18610);
or U19662 (N_19662,N_15037,N_17159);
or U19663 (N_19663,N_16863,N_16348);
xor U19664 (N_19664,N_14886,N_17361);
nand U19665 (N_19665,N_12727,N_16263);
nand U19666 (N_19666,N_16837,N_14374);
or U19667 (N_19667,N_18535,N_14205);
nand U19668 (N_19668,N_12625,N_16215);
xor U19669 (N_19669,N_18691,N_17559);
nand U19670 (N_19670,N_13089,N_14063);
and U19671 (N_19671,N_15073,N_12703);
nand U19672 (N_19672,N_14585,N_16971);
nor U19673 (N_19673,N_15079,N_17601);
or U19674 (N_19674,N_13258,N_15542);
or U19675 (N_19675,N_15412,N_14248);
nand U19676 (N_19676,N_12939,N_16815);
or U19677 (N_19677,N_12851,N_17510);
and U19678 (N_19678,N_13147,N_17499);
nor U19679 (N_19679,N_12797,N_15696);
or U19680 (N_19680,N_16474,N_16184);
and U19681 (N_19681,N_12988,N_18316);
nand U19682 (N_19682,N_16990,N_16360);
nand U19683 (N_19683,N_16493,N_13301);
nand U19684 (N_19684,N_18218,N_12952);
nor U19685 (N_19685,N_12777,N_14944);
or U19686 (N_19686,N_12947,N_14618);
nand U19687 (N_19687,N_17430,N_12937);
and U19688 (N_19688,N_13318,N_17411);
and U19689 (N_19689,N_18090,N_17504);
nor U19690 (N_19690,N_17362,N_13907);
and U19691 (N_19691,N_18472,N_13127);
or U19692 (N_19692,N_15207,N_14939);
nor U19693 (N_19693,N_14470,N_15357);
xnor U19694 (N_19694,N_15937,N_15679);
nand U19695 (N_19695,N_18410,N_14789);
and U19696 (N_19696,N_13653,N_18598);
nand U19697 (N_19697,N_16152,N_16556);
nand U19698 (N_19698,N_17508,N_14228);
nor U19699 (N_19699,N_18454,N_13005);
nor U19700 (N_19700,N_15323,N_16879);
or U19701 (N_19701,N_17062,N_16523);
or U19702 (N_19702,N_13952,N_18509);
and U19703 (N_19703,N_16036,N_18249);
xor U19704 (N_19704,N_14391,N_15678);
nand U19705 (N_19705,N_18436,N_15093);
nand U19706 (N_19706,N_17937,N_14054);
or U19707 (N_19707,N_16941,N_12508);
and U19708 (N_19708,N_14125,N_17098);
or U19709 (N_19709,N_14317,N_16774);
and U19710 (N_19710,N_12696,N_12992);
or U19711 (N_19711,N_16355,N_15121);
nand U19712 (N_19712,N_17392,N_18477);
nor U19713 (N_19713,N_15662,N_17131);
nor U19714 (N_19714,N_12668,N_13828);
or U19715 (N_19715,N_16949,N_18692);
nand U19716 (N_19716,N_15643,N_18701);
nand U19717 (N_19717,N_13368,N_14940);
nor U19718 (N_19718,N_18132,N_16640);
xor U19719 (N_19719,N_18248,N_18381);
or U19720 (N_19720,N_14994,N_18124);
or U19721 (N_19721,N_13112,N_15952);
and U19722 (N_19722,N_14138,N_12810);
xor U19723 (N_19723,N_13057,N_15621);
nand U19724 (N_19724,N_16973,N_17168);
and U19725 (N_19725,N_13732,N_18719);
or U19726 (N_19726,N_15704,N_12815);
nor U19727 (N_19727,N_12689,N_15509);
nand U19728 (N_19728,N_16325,N_18342);
nor U19729 (N_19729,N_14661,N_16987);
nand U19730 (N_19730,N_16846,N_15567);
nor U19731 (N_19731,N_15799,N_13117);
nand U19732 (N_19732,N_14688,N_12690);
or U19733 (N_19733,N_15856,N_17037);
nor U19734 (N_19734,N_13783,N_17860);
and U19735 (N_19735,N_17579,N_15082);
xnor U19736 (N_19736,N_14893,N_15502);
nor U19737 (N_19737,N_16767,N_17039);
nand U19738 (N_19738,N_14888,N_13378);
nor U19739 (N_19739,N_18611,N_15891);
nor U19740 (N_19740,N_15329,N_15052);
xor U19741 (N_19741,N_16625,N_14090);
nor U19742 (N_19742,N_12959,N_14900);
nor U19743 (N_19743,N_16850,N_17340);
and U19744 (N_19744,N_13776,N_15291);
nor U19745 (N_19745,N_17058,N_13468);
or U19746 (N_19746,N_13522,N_14620);
nand U19747 (N_19747,N_13213,N_13344);
or U19748 (N_19748,N_15226,N_15893);
or U19749 (N_19749,N_13365,N_13893);
or U19750 (N_19750,N_15607,N_17100);
nor U19751 (N_19751,N_17599,N_16834);
or U19752 (N_19752,N_15640,N_15811);
nor U19753 (N_19753,N_13211,N_18373);
and U19754 (N_19754,N_13991,N_16568);
nand U19755 (N_19755,N_15668,N_16788);
and U19756 (N_19756,N_15551,N_14626);
or U19757 (N_19757,N_12574,N_13701);
and U19758 (N_19758,N_16616,N_17839);
nand U19759 (N_19759,N_15254,N_12650);
or U19760 (N_19760,N_18459,N_16659);
nor U19761 (N_19761,N_16904,N_12500);
nand U19762 (N_19762,N_15660,N_16599);
nand U19763 (N_19763,N_16049,N_18125);
nor U19764 (N_19764,N_16590,N_18540);
or U19765 (N_19765,N_13697,N_18082);
or U19766 (N_19766,N_18633,N_16302);
nor U19767 (N_19767,N_13935,N_15635);
nor U19768 (N_19768,N_18338,N_16241);
and U19769 (N_19769,N_14087,N_18318);
nand U19770 (N_19770,N_18226,N_18510);
and U19771 (N_19771,N_15598,N_13982);
nand U19772 (N_19772,N_13814,N_15725);
nor U19773 (N_19773,N_14379,N_14131);
or U19774 (N_19774,N_13391,N_13231);
nand U19775 (N_19775,N_16962,N_18490);
nand U19776 (N_19776,N_13241,N_12787);
nand U19777 (N_19777,N_15206,N_14488);
or U19778 (N_19778,N_16939,N_17083);
and U19779 (N_19779,N_14584,N_15271);
nor U19780 (N_19780,N_17672,N_13334);
and U19781 (N_19781,N_18712,N_17439);
xor U19782 (N_19782,N_14516,N_14969);
or U19783 (N_19783,N_15699,N_15717);
nor U19784 (N_19784,N_17064,N_14085);
nand U19785 (N_19785,N_18577,N_17819);
and U19786 (N_19786,N_13052,N_16012);
xor U19787 (N_19787,N_15961,N_17889);
nand U19788 (N_19788,N_16785,N_12594);
nor U19789 (N_19789,N_18189,N_14245);
or U19790 (N_19790,N_12735,N_17353);
nor U19791 (N_19791,N_16722,N_16826);
nand U19792 (N_19792,N_13746,N_14446);
and U19793 (N_19793,N_16830,N_18220);
and U19794 (N_19794,N_16466,N_15421);
nand U19795 (N_19795,N_17776,N_12801);
and U19796 (N_19796,N_17808,N_13803);
and U19797 (N_19797,N_18296,N_15616);
xnor U19798 (N_19798,N_12984,N_16720);
nor U19799 (N_19799,N_15855,N_17263);
xnor U19800 (N_19800,N_16802,N_18223);
xnor U19801 (N_19801,N_13051,N_14727);
or U19802 (N_19802,N_14062,N_14239);
or U19803 (N_19803,N_17424,N_17708);
or U19804 (N_19804,N_13263,N_17874);
or U19805 (N_19805,N_13523,N_13054);
or U19806 (N_19806,N_14406,N_14369);
nor U19807 (N_19807,N_18557,N_16315);
nor U19808 (N_19808,N_13794,N_14432);
or U19809 (N_19809,N_16495,N_15017);
and U19810 (N_19810,N_13553,N_12586);
and U19811 (N_19811,N_17300,N_13752);
xor U19812 (N_19812,N_14192,N_17516);
or U19813 (N_19813,N_16766,N_17095);
or U19814 (N_19814,N_18059,N_18301);
and U19815 (N_19815,N_17817,N_15867);
nand U19816 (N_19816,N_18088,N_15043);
and U19817 (N_19817,N_16840,N_14434);
nand U19818 (N_19818,N_12621,N_13343);
or U19819 (N_19819,N_18245,N_18228);
and U19820 (N_19820,N_17915,N_16953);
nand U19821 (N_19821,N_14242,N_18241);
xnor U19822 (N_19822,N_18145,N_13411);
or U19823 (N_19823,N_17432,N_16533);
nor U19824 (N_19824,N_17990,N_18302);
nor U19825 (N_19825,N_14464,N_15391);
and U19826 (N_19826,N_17224,N_18403);
nor U19827 (N_19827,N_17356,N_16964);
and U19828 (N_19828,N_18618,N_12540);
nand U19829 (N_19829,N_16972,N_15852);
and U19830 (N_19830,N_12889,N_17964);
or U19831 (N_19831,N_17506,N_13088);
and U19832 (N_19832,N_17379,N_15927);
or U19833 (N_19833,N_16450,N_15708);
nor U19834 (N_19834,N_16983,N_14217);
nor U19835 (N_19835,N_17046,N_14677);
nand U19836 (N_19836,N_17643,N_15894);
nand U19837 (N_19837,N_17787,N_13944);
or U19838 (N_19838,N_17090,N_18463);
or U19839 (N_19839,N_14612,N_16701);
or U19840 (N_19840,N_17813,N_16276);
and U19841 (N_19841,N_17763,N_18476);
nor U19842 (N_19842,N_17794,N_16310);
or U19843 (N_19843,N_14568,N_16621);
nand U19844 (N_19844,N_17531,N_13488);
or U19845 (N_19845,N_16618,N_13555);
nand U19846 (N_19846,N_12615,N_15833);
or U19847 (N_19847,N_14072,N_16309);
nor U19848 (N_19848,N_16893,N_13518);
nand U19849 (N_19849,N_15150,N_14914);
nand U19850 (N_19850,N_12792,N_17368);
nand U19851 (N_19851,N_15884,N_14762);
and U19852 (N_19852,N_15422,N_15905);
nand U19853 (N_19853,N_15178,N_18596);
or U19854 (N_19854,N_16108,N_14698);
nand U19855 (N_19855,N_17953,N_17585);
nor U19856 (N_19856,N_14347,N_18267);
and U19857 (N_19857,N_15358,N_13283);
and U19858 (N_19858,N_14197,N_15638);
and U19859 (N_19859,N_18397,N_16647);
nand U19860 (N_19860,N_14791,N_15506);
nand U19861 (N_19861,N_14632,N_17434);
nand U19862 (N_19862,N_13853,N_13281);
nand U19863 (N_19863,N_16368,N_14352);
nor U19864 (N_19864,N_17429,N_17842);
nand U19865 (N_19865,N_16490,N_16991);
nand U19866 (N_19866,N_16090,N_15789);
or U19867 (N_19867,N_17589,N_14666);
and U19868 (N_19868,N_13487,N_16557);
and U19869 (N_19869,N_18749,N_12702);
or U19870 (N_19870,N_15724,N_17811);
nor U19871 (N_19871,N_14049,N_17346);
nand U19872 (N_19872,N_14546,N_12698);
nor U19873 (N_19873,N_18185,N_13309);
xor U19874 (N_19874,N_17553,N_14301);
and U19875 (N_19875,N_16955,N_13098);
xnor U19876 (N_19876,N_15955,N_16764);
and U19877 (N_19877,N_14793,N_14558);
nor U19878 (N_19878,N_15062,N_15697);
nand U19879 (N_19879,N_17544,N_16051);
nand U19880 (N_19880,N_16149,N_15776);
nor U19881 (N_19881,N_16438,N_17720);
nor U19882 (N_19882,N_18212,N_15974);
nand U19883 (N_19883,N_15805,N_15615);
nor U19884 (N_19884,N_14984,N_14137);
nor U19885 (N_19885,N_15281,N_14257);
and U19886 (N_19886,N_18603,N_16814);
or U19887 (N_19887,N_13370,N_18447);
xnor U19888 (N_19888,N_17809,N_14520);
nor U19889 (N_19889,N_16133,N_13067);
and U19890 (N_19890,N_16344,N_14961);
nor U19891 (N_19891,N_13797,N_13583);
xnor U19892 (N_19892,N_18201,N_14189);
or U19893 (N_19893,N_12719,N_14208);
and U19894 (N_19894,N_13024,N_12740);
nand U19895 (N_19895,N_13942,N_13605);
nand U19896 (N_19896,N_18219,N_18556);
and U19897 (N_19897,N_13830,N_17207);
nor U19898 (N_19898,N_17022,N_14636);
and U19899 (N_19899,N_14513,N_14079);
xor U19900 (N_19900,N_13131,N_17667);
nand U19901 (N_19901,N_14476,N_12925);
or U19902 (N_19902,N_18714,N_13664);
nand U19903 (N_19903,N_17327,N_17771);
nor U19904 (N_19904,N_15700,N_18612);
or U19905 (N_19905,N_14142,N_17453);
nand U19906 (N_19906,N_18631,N_17802);
and U19907 (N_19907,N_17966,N_14166);
and U19908 (N_19908,N_14030,N_13955);
nor U19909 (N_19909,N_12552,N_17534);
and U19910 (N_19910,N_13824,N_15138);
nor U19911 (N_19911,N_12566,N_16933);
or U19912 (N_19912,N_13615,N_13648);
and U19913 (N_19913,N_15845,N_15579);
and U19914 (N_19914,N_14380,N_16924);
and U19915 (N_19915,N_12861,N_18204);
nand U19916 (N_19916,N_14408,N_16779);
xor U19917 (N_19917,N_18270,N_16575);
or U19918 (N_19918,N_15781,N_14384);
and U19919 (N_19919,N_15872,N_18046);
nor U19920 (N_19920,N_16291,N_16282);
nor U19921 (N_19921,N_14240,N_15823);
xnor U19922 (N_19922,N_12522,N_18235);
and U19923 (N_19923,N_16008,N_15513);
xor U19924 (N_19924,N_16956,N_14052);
and U19925 (N_19925,N_16453,N_17749);
or U19926 (N_19926,N_14820,N_15689);
nand U19927 (N_19927,N_15757,N_13469);
and U19928 (N_19928,N_13534,N_14880);
and U19929 (N_19929,N_14597,N_14704);
nor U19930 (N_19930,N_18529,N_14952);
nand U19931 (N_19931,N_13609,N_17928);
and U19932 (N_19932,N_18665,N_14718);
nand U19933 (N_19933,N_13891,N_17376);
nor U19934 (N_19934,N_13507,N_15993);
nor U19935 (N_19935,N_16811,N_15723);
nand U19936 (N_19936,N_13700,N_15609);
and U19937 (N_19937,N_17917,N_12837);
nor U19938 (N_19938,N_15029,N_13785);
nand U19939 (N_19939,N_14399,N_12802);
or U19940 (N_19940,N_12821,N_14160);
nand U19941 (N_19941,N_17929,N_16598);
or U19942 (N_19942,N_15067,N_18425);
xor U19943 (N_19943,N_18080,N_12677);
or U19944 (N_19944,N_12511,N_13985);
nor U19945 (N_19945,N_18291,N_13530);
and U19946 (N_19946,N_13155,N_17497);
and U19947 (N_19947,N_13393,N_14452);
nand U19948 (N_19948,N_16292,N_16712);
or U19949 (N_19949,N_15047,N_15820);
xor U19950 (N_19950,N_13860,N_15403);
xnor U19951 (N_19951,N_17074,N_18506);
and U19952 (N_19952,N_17479,N_18083);
nand U19953 (N_19953,N_18197,N_14981);
or U19954 (N_19954,N_17581,N_12820);
nand U19955 (N_19955,N_13300,N_16463);
nor U19956 (N_19956,N_13691,N_16267);
nand U19957 (N_19957,N_13808,N_16265);
and U19958 (N_19958,N_14051,N_12632);
nand U19959 (N_19959,N_15355,N_15348);
or U19960 (N_19960,N_13187,N_16255);
or U19961 (N_19961,N_16058,N_14669);
nor U19962 (N_19962,N_12954,N_16750);
xnor U19963 (N_19963,N_14581,N_13680);
xor U19964 (N_19964,N_15873,N_15627);
nor U19965 (N_19965,N_16605,N_13242);
or U19966 (N_19966,N_13588,N_13502);
xor U19967 (N_19967,N_17768,N_13597);
xor U19968 (N_19968,N_15483,N_14699);
and U19969 (N_19969,N_12509,N_18394);
or U19970 (N_19970,N_13311,N_13374);
nor U19971 (N_19971,N_17853,N_15173);
and U19972 (N_19972,N_16439,N_13738);
and U19973 (N_19973,N_13165,N_17958);
or U19974 (N_19974,N_12871,N_15763);
and U19975 (N_19975,N_14449,N_17009);
or U19976 (N_19976,N_13272,N_15013);
nand U19977 (N_19977,N_13600,N_18187);
and U19978 (N_19978,N_12791,N_13721);
or U19979 (N_19979,N_14804,N_18356);
nor U19980 (N_19980,N_13325,N_13236);
nand U19981 (N_19981,N_16822,N_12804);
or U19982 (N_19982,N_17987,N_12572);
and U19983 (N_19983,N_12579,N_15547);
xnor U19984 (N_19984,N_13557,N_16442);
and U19985 (N_19985,N_14336,N_14926);
and U19986 (N_19986,N_16124,N_17420);
nor U19987 (N_19987,N_15865,N_14103);
or U19988 (N_19988,N_14451,N_17635);
or U19989 (N_19989,N_13696,N_13813);
nor U19990 (N_19990,N_13705,N_15381);
xnor U19991 (N_19991,N_18163,N_14121);
nand U19992 (N_19992,N_16468,N_13100);
nand U19993 (N_19993,N_12844,N_13533);
xnor U19994 (N_19994,N_18533,N_16805);
nor U19995 (N_19995,N_16587,N_13304);
nor U19996 (N_19996,N_14653,N_17514);
xnor U19997 (N_19997,N_14732,N_14273);
and U19998 (N_19998,N_13674,N_15296);
nand U19999 (N_19999,N_17126,N_13967);
xnor U20000 (N_20000,N_12968,N_18029);
or U20001 (N_20001,N_14264,N_13161);
and U20002 (N_20002,N_16294,N_17081);
and U20003 (N_20003,N_14531,N_14800);
or U20004 (N_20004,N_13969,N_18109);
and U20005 (N_20005,N_16980,N_14814);
or U20006 (N_20006,N_17827,N_16233);
and U20007 (N_20007,N_17625,N_14659);
nor U20008 (N_20008,N_14511,N_12637);
nor U20009 (N_20009,N_15490,N_12545);
and U20010 (N_20010,N_15572,N_17108);
nor U20011 (N_20011,N_13026,N_17736);
and U20012 (N_20012,N_16942,N_15482);
and U20013 (N_20013,N_16610,N_15529);
nor U20014 (N_20014,N_16739,N_15733);
nand U20015 (N_20015,N_14297,N_15250);
nand U20016 (N_20016,N_15743,N_13109);
or U20017 (N_20017,N_17998,N_16482);
or U20018 (N_20018,N_16998,N_14304);
nand U20019 (N_20019,N_15459,N_16287);
and U20020 (N_20020,N_18254,N_18401);
or U20021 (N_20021,N_13574,N_15667);
nor U20022 (N_20022,N_15702,N_13494);
nor U20023 (N_20023,N_18622,N_18328);
xor U20024 (N_20024,N_16996,N_18723);
and U20025 (N_20025,N_17766,N_15069);
or U20026 (N_20026,N_12681,N_14707);
xor U20027 (N_20027,N_12914,N_13430);
nand U20028 (N_20028,N_15682,N_15941);
and U20029 (N_20029,N_12867,N_18504);
and U20030 (N_20030,N_13280,N_18363);
or U20031 (N_20031,N_17191,N_15426);
nand U20032 (N_20032,N_13087,N_13319);
nor U20033 (N_20033,N_12870,N_16145);
and U20034 (N_20034,N_13556,N_17293);
or U20035 (N_20035,N_16365,N_16331);
or U20036 (N_20036,N_13139,N_15087);
nand U20037 (N_20037,N_17780,N_13521);
and U20038 (N_20038,N_15305,N_17433);
nor U20039 (N_20039,N_13115,N_18437);
xnor U20040 (N_20040,N_12897,N_16204);
nand U20041 (N_20041,N_13068,N_12634);
or U20042 (N_20042,N_16354,N_13519);
nor U20043 (N_20043,N_15316,N_16127);
and U20044 (N_20044,N_14150,N_15285);
nand U20045 (N_20045,N_15232,N_16369);
nor U20046 (N_20046,N_17374,N_18048);
xnor U20047 (N_20047,N_13886,N_12527);
nor U20048 (N_20048,N_17457,N_14302);
and U20049 (N_20049,N_16643,N_14144);
or U20050 (N_20050,N_16997,N_16806);
or U20051 (N_20051,N_13589,N_13257);
nand U20052 (N_20052,N_13974,N_15695);
nor U20053 (N_20053,N_15432,N_13489);
or U20054 (N_20054,N_15594,N_15167);
or U20055 (N_20055,N_15293,N_18320);
xor U20056 (N_20056,N_18519,N_12651);
and U20057 (N_20057,N_15452,N_15991);
nor U20058 (N_20058,N_16166,N_17299);
or U20059 (N_20059,N_18011,N_13275);
or U20060 (N_20060,N_14096,N_15986);
nand U20061 (N_20061,N_16689,N_14027);
or U20062 (N_20062,N_13351,N_16707);
and U20063 (N_20063,N_12878,N_18188);
and U20064 (N_20064,N_13657,N_17127);
and U20065 (N_20065,N_13348,N_13209);
or U20066 (N_20066,N_14414,N_16912);
xor U20067 (N_20067,N_15610,N_13384);
nand U20068 (N_20068,N_13823,N_13113);
and U20069 (N_20069,N_15775,N_17261);
nor U20070 (N_20070,N_17838,N_16296);
nor U20071 (N_20071,N_14860,N_13465);
or U20072 (N_20072,N_12737,N_15378);
and U20073 (N_20073,N_14398,N_18259);
xnor U20074 (N_20074,N_17101,N_15670);
or U20075 (N_20075,N_13928,N_17769);
nor U20076 (N_20076,N_12880,N_15024);
or U20077 (N_20077,N_14061,N_18377);
xnor U20078 (N_20078,N_16583,N_12832);
nor U20079 (N_20079,N_16527,N_13493);
xor U20080 (N_20080,N_13901,N_13405);
or U20081 (N_20081,N_15352,N_18462);
nor U20082 (N_20082,N_17097,N_13686);
nor U20083 (N_20083,N_17448,N_15576);
xnor U20084 (N_20084,N_17952,N_14046);
or U20085 (N_20085,N_14729,N_13767);
or U20086 (N_20086,N_18229,N_17367);
or U20087 (N_20087,N_13855,N_14638);
nor U20088 (N_20088,N_17030,N_12987);
nand U20089 (N_20089,N_13619,N_17048);
nand U20090 (N_20090,N_14515,N_14501);
and U20091 (N_20091,N_14430,N_15756);
or U20092 (N_20092,N_13636,N_13480);
and U20093 (N_20093,N_12834,N_16318);
nand U20094 (N_20094,N_12655,N_13630);
and U20095 (N_20095,N_14038,N_15779);
nand U20096 (N_20096,N_12692,N_14040);
xnor U20097 (N_20097,N_13239,N_17313);
or U20098 (N_20098,N_17078,N_15300);
nor U20099 (N_20099,N_13228,N_17255);
and U20100 (N_20100,N_18015,N_18645);
nor U20101 (N_20101,N_16488,N_14767);
and U20102 (N_20102,N_15601,N_18524);
or U20103 (N_20103,N_16498,N_14310);
and U20104 (N_20104,N_18289,N_15170);
nand U20105 (N_20105,N_16967,N_16374);
and U20106 (N_20106,N_12701,N_15817);
or U20107 (N_20107,N_18309,N_16373);
and U20108 (N_20108,N_13909,N_13323);
nand U20109 (N_20109,N_13562,N_16256);
nor U20110 (N_20110,N_16632,N_15075);
xor U20111 (N_20111,N_18334,N_16671);
xor U20112 (N_20112,N_13387,N_12578);
nor U20113 (N_20113,N_13172,N_14246);
xnor U20114 (N_20114,N_14705,N_12556);
and U20115 (N_20115,N_15220,N_14865);
nand U20116 (N_20116,N_17197,N_13677);
nand U20117 (N_20117,N_18538,N_17351);
or U20118 (N_20118,N_13394,N_15102);
nand U20119 (N_20119,N_12729,N_13531);
or U20120 (N_20120,N_17507,N_14995);
nor U20121 (N_20121,N_18097,N_13039);
or U20122 (N_20122,N_17107,N_16239);
or U20123 (N_20123,N_13157,N_12708);
nor U20124 (N_20124,N_18049,N_16349);
or U20125 (N_20125,N_13462,N_12973);
nand U20126 (N_20126,N_18294,N_17205);
or U20127 (N_20127,N_12902,N_17611);
and U20128 (N_20128,N_15068,N_15292);
nor U20129 (N_20129,N_14590,N_16563);
and U20130 (N_20130,N_17210,N_14794);
nor U20131 (N_20131,N_18378,N_16038);
nand U20132 (N_20132,N_14917,N_14420);
and U20133 (N_20133,N_15306,N_17157);
or U20134 (N_20134,N_15505,N_14437);
and U20135 (N_20135,N_15739,N_15175);
or U20136 (N_20136,N_12977,N_12953);
nor U20137 (N_20137,N_18288,N_18271);
or U20138 (N_20138,N_14964,N_16601);
or U20139 (N_20139,N_15471,N_12664);
nand U20140 (N_20140,N_13527,N_13826);
nand U20141 (N_20141,N_13193,N_15522);
xor U20142 (N_20142,N_13203,N_14564);
nand U20143 (N_20143,N_15501,N_17363);
and U20144 (N_20144,N_13341,N_15853);
nor U20145 (N_20145,N_14877,N_18268);
nand U20146 (N_20146,N_16066,N_16657);
or U20147 (N_20147,N_17179,N_18148);
and U20148 (N_20148,N_15983,N_18417);
nor U20149 (N_20149,N_13388,N_14866);
nor U20150 (N_20150,N_17732,N_13675);
nor U20151 (N_20151,N_15136,N_14890);
nand U20152 (N_20152,N_17618,N_18541);
and U20153 (N_20153,N_17899,N_16410);
nand U20154 (N_20154,N_18599,N_15371);
nand U20155 (N_20155,N_16977,N_17066);
nand U20156 (N_20156,N_13445,N_18703);
xnor U20157 (N_20157,N_18740,N_12506);
nand U20158 (N_20158,N_14909,N_14265);
nor U20159 (N_20159,N_16653,N_12944);
or U20160 (N_20160,N_15228,N_17976);
xnor U20161 (N_20161,N_16168,N_13270);
and U20162 (N_20162,N_16414,N_14207);
and U20163 (N_20163,N_14418,N_12505);
and U20164 (N_20164,N_17306,N_17593);
nor U20165 (N_20165,N_14507,N_14123);
or U20166 (N_20166,N_17460,N_16417);
nor U20167 (N_20167,N_13622,N_16336);
and U20168 (N_20168,N_12974,N_17631);
and U20169 (N_20169,N_15217,N_17043);
and U20170 (N_20170,N_17285,N_12648);
and U20171 (N_20171,N_14289,N_13872);
nor U20172 (N_20172,N_17145,N_15842);
nand U20173 (N_20173,N_13770,N_12557);
nand U20174 (N_20174,N_14365,N_12868);
or U20175 (N_20175,N_14544,N_16217);
or U20176 (N_20176,N_16244,N_15963);
nor U20177 (N_20177,N_16668,N_14013);
nand U20178 (N_20178,N_14723,N_13958);
or U20179 (N_20179,N_14075,N_13923);
nand U20180 (N_20180,N_14902,N_16951);
xor U20181 (N_20181,N_16528,N_18076);
nor U20182 (N_20182,N_14595,N_13282);
nor U20183 (N_20183,N_13149,N_13416);
or U20184 (N_20184,N_13168,N_12750);
nand U20185 (N_20185,N_12657,N_12823);
nor U20186 (N_20186,N_14419,N_16446);
nand U20187 (N_20187,N_15752,N_13449);
nor U20188 (N_20188,N_15269,N_15418);
and U20189 (N_20189,N_13339,N_14492);
or U20190 (N_20190,N_18563,N_17339);
nor U20191 (N_20191,N_13626,N_15416);
or U20192 (N_20192,N_13420,N_12755);
and U20193 (N_20193,N_16073,N_15661);
or U20194 (N_20194,N_14506,N_18222);
or U20195 (N_20195,N_12671,N_17068);
and U20196 (N_20196,N_16670,N_16633);
and U20197 (N_20197,N_14206,N_18068);
xnor U20198 (N_20198,N_13835,N_13071);
or U20199 (N_20199,N_15476,N_14132);
nor U20200 (N_20200,N_17318,N_15467);
or U20201 (N_20201,N_14181,N_16307);
and U20202 (N_20202,N_12639,N_15625);
nor U20203 (N_20203,N_17389,N_15326);
nor U20204 (N_20204,N_14502,N_13245);
or U20205 (N_20205,N_15027,N_14306);
or U20206 (N_20206,N_13328,N_17798);
or U20207 (N_20207,N_17124,N_16606);
xnor U20208 (N_20208,N_14343,N_15874);
nor U20209 (N_20209,N_16500,N_15277);
or U20210 (N_20210,N_14989,N_16104);
or U20211 (N_20211,N_15792,N_17898);
and U20212 (N_20212,N_13756,N_15624);
nand U20213 (N_20213,N_12515,N_12796);
or U20214 (N_20214,N_17075,N_17546);
nor U20215 (N_20215,N_13719,N_17397);
or U20216 (N_20216,N_17658,N_14321);
xnor U20217 (N_20217,N_17669,N_17951);
and U20218 (N_20218,N_14797,N_15990);
or U20219 (N_20219,N_13424,N_17173);
or U20220 (N_20220,N_14497,N_13856);
nand U20221 (N_20221,N_16094,N_17844);
or U20222 (N_20222,N_14766,N_16518);
and U20223 (N_20223,N_16362,N_13491);
or U20224 (N_20224,N_16639,N_15114);
and U20225 (N_20225,N_15738,N_13846);
nand U20226 (N_20226,N_15216,N_16697);
and U20227 (N_20227,N_12927,N_14734);
nor U20228 (N_20228,N_16554,N_14479);
nor U20229 (N_20229,N_12928,N_17591);
nand U20230 (N_20230,N_16340,N_17342);
nor U20231 (N_20231,N_17444,N_13709);
or U20232 (N_20232,N_15096,N_13357);
and U20233 (N_20233,N_13037,N_14634);
and U20234 (N_20234,N_14141,N_14500);
and U20235 (N_20235,N_14932,N_16479);
nand U20236 (N_20236,N_14104,N_17849);
nand U20237 (N_20237,N_13753,N_12546);
nor U20238 (N_20238,N_14541,N_15705);
nand U20239 (N_20239,N_14126,N_18230);
xor U20240 (N_20240,N_17905,N_13866);
and U20241 (N_20241,N_16794,N_17274);
nand U20242 (N_20242,N_13571,N_18482);
and U20243 (N_20243,N_12893,N_16084);
or U20244 (N_20244,N_16433,N_16043);
nand U20245 (N_20245,N_17056,N_15686);
or U20246 (N_20246,N_13062,N_15951);
nand U20247 (N_20247,N_18605,N_15840);
nor U20248 (N_20248,N_18662,N_18735);
nand U20249 (N_20249,N_12534,N_17946);
nand U20250 (N_20250,N_13796,N_18696);
nor U20251 (N_20251,N_18166,N_13960);
nand U20252 (N_20252,N_14937,N_17369);
nand U20253 (N_20253,N_13838,N_13240);
nand U20254 (N_20254,N_13204,N_16150);
xnor U20255 (N_20255,N_16220,N_15861);
nor U20256 (N_20256,N_14675,N_16740);
xnor U20257 (N_20257,N_15275,N_18130);
or U20258 (N_20258,N_16704,N_12585);
and U20259 (N_20259,N_16635,N_16429);
or U20260 (N_20260,N_13254,N_18392);
nand U20261 (N_20261,N_18391,N_16082);
nand U20262 (N_20262,N_12936,N_14435);
nand U20263 (N_20263,N_13580,N_18532);
and U20264 (N_20264,N_15639,N_15968);
or U20265 (N_20265,N_14308,N_13120);
or U20266 (N_20266,N_15657,N_16617);
or U20267 (N_20267,N_16350,N_17294);
or U20268 (N_20268,N_12976,N_12503);
nor U20269 (N_20269,N_16489,N_14426);
nand U20270 (N_20270,N_12999,N_17983);
or U20271 (N_20271,N_14572,N_15100);
or U20272 (N_20272,N_16447,N_17913);
xnor U20273 (N_20273,N_14227,N_14088);
or U20274 (N_20274,N_14332,N_17722);
nand U20275 (N_20275,N_18697,N_17637);
or U20276 (N_20276,N_13125,N_15835);
xor U20277 (N_20277,N_17828,N_18236);
or U20278 (N_20278,N_18173,N_13196);
nand U20279 (N_20279,N_16284,N_17527);
nor U20280 (N_20280,N_17810,N_16509);
nand U20281 (N_20281,N_18096,N_13038);
or U20282 (N_20282,N_18693,N_13407);
nor U20283 (N_20283,N_15433,N_14118);
and U20284 (N_20284,N_17121,N_17610);
and U20285 (N_20285,N_18408,N_15798);
nor U20286 (N_20286,N_15533,N_13150);
nor U20287 (N_20287,N_13030,N_18559);
xnor U20288 (N_20288,N_18460,N_16838);
or U20289 (N_20289,N_15118,N_12782);
nor U20290 (N_20290,N_17997,N_15342);
and U20291 (N_20291,N_18041,N_14201);
xor U20292 (N_20292,N_14249,N_17668);
nand U20293 (N_20293,N_14278,N_15783);
and U20294 (N_20294,N_16092,N_14781);
nand U20295 (N_20295,N_18225,N_16465);
and U20296 (N_20296,N_15954,N_12752);
and U20297 (N_20297,N_13857,N_15740);
or U20298 (N_20298,N_15180,N_17352);
nor U20299 (N_20299,N_18054,N_17614);
nor U20300 (N_20300,N_16351,N_15791);
xnor U20301 (N_20301,N_18578,N_14614);
nor U20302 (N_20302,N_17943,N_18179);
and U20303 (N_20303,N_17781,N_18052);
xor U20304 (N_20304,N_15479,N_17350);
nand U20305 (N_20305,N_14924,N_12809);
nor U20306 (N_20306,N_13889,N_13816);
nand U20307 (N_20307,N_18200,N_13852);
or U20308 (N_20308,N_17138,N_18240);
nand U20309 (N_20309,N_15235,N_17450);
xor U20310 (N_20310,N_17212,N_13013);
and U20311 (N_20311,N_16516,N_18115);
nand U20312 (N_20312,N_18521,N_13132);
nor U20313 (N_20313,N_14821,N_17561);
xor U20314 (N_20314,N_14260,N_15183);
or U20315 (N_20315,N_18244,N_13508);
nand U20316 (N_20316,N_17543,N_18277);
or U20317 (N_20317,N_16677,N_15909);
nand U20318 (N_20318,N_15809,N_14971);
and U20319 (N_20319,N_13639,N_15147);
and U20320 (N_20320,N_17400,N_17151);
and U20321 (N_20321,N_16978,N_16080);
nor U20322 (N_20322,N_14505,N_16075);
and U20323 (N_20323,N_12945,N_13467);
or U20324 (N_20324,N_18707,N_15574);
or U20325 (N_20325,N_13678,N_13473);
nor U20326 (N_20326,N_14575,N_15301);
nor U20327 (N_20327,N_16559,N_16114);
xnor U20328 (N_20328,N_13566,N_14955);
xnor U20329 (N_20329,N_15524,N_14463);
nor U20330 (N_20330,N_15854,N_17259);
or U20331 (N_20331,N_16860,N_17167);
and U20332 (N_20332,N_16390,N_16097);
and U20333 (N_20333,N_16782,N_15021);
nor U20334 (N_20334,N_16748,N_16902);
nand U20335 (N_20335,N_15364,N_12682);
or U20336 (N_20336,N_16099,N_17639);
nor U20337 (N_20337,N_15055,N_17973);
nor U20338 (N_20338,N_18142,N_18402);
nand U20339 (N_20339,N_13854,N_14948);
nand U20340 (N_20340,N_17654,N_18520);
nor U20341 (N_20341,N_17986,N_13252);
and U20342 (N_20342,N_18593,N_17577);
nor U20343 (N_20343,N_17275,N_14478);
nand U20344 (N_20344,N_17655,N_16873);
nor U20345 (N_20345,N_14395,N_17080);
or U20346 (N_20346,N_15427,N_15257);
nor U20347 (N_20347,N_14436,N_12697);
and U20348 (N_20348,N_16726,N_17563);
nand U20349 (N_20349,N_15674,N_16781);
or U20350 (N_20350,N_16692,N_15091);
or U20351 (N_20351,N_13795,N_14295);
nand U20352 (N_20352,N_17541,N_12523);
nor U20353 (N_20353,N_13310,N_16426);
nand U20354 (N_20354,N_16859,N_16839);
nand U20355 (N_20355,N_13363,N_17181);
nand U20356 (N_20356,N_16370,N_16260);
or U20357 (N_20357,N_17566,N_13171);
or U20358 (N_20358,N_17738,N_15372);
nand U20359 (N_20359,N_15535,N_18653);
nand U20360 (N_20360,N_18194,N_13859);
nand U20361 (N_20361,N_16547,N_15584);
nand U20362 (N_20362,N_14611,N_16091);
and U20363 (N_20363,N_17868,N_17052);
or U20364 (N_20364,N_14599,N_15246);
or U20365 (N_20365,N_18479,N_17269);
nand U20366 (N_20366,N_12613,N_17072);
and U20367 (N_20367,N_17684,N_17818);
nor U20368 (N_20368,N_16676,N_16289);
and U20369 (N_20369,N_17203,N_16663);
nand U20370 (N_20370,N_17135,N_13048);
and U20371 (N_20371,N_12906,N_15133);
nand U20372 (N_20372,N_16555,N_14037);
nor U20373 (N_20373,N_13049,N_12561);
xor U20374 (N_20374,N_17311,N_12666);
and U20375 (N_20375,N_18702,N_14721);
or U20376 (N_20376,N_15419,N_17908);
or U20377 (N_20377,N_12949,N_18323);
or U20378 (N_20378,N_18110,N_17617);
and U20379 (N_20379,N_17393,N_18637);
nand U20380 (N_20380,N_14760,N_18319);
nor U20381 (N_20381,N_15333,N_14417);
nor U20382 (N_20382,N_14754,N_14475);
and U20383 (N_20383,N_15568,N_12660);
and U20384 (N_20384,N_13007,N_15125);
nand U20385 (N_20385,N_14534,N_14667);
xnor U20386 (N_20386,N_13815,N_15999);
nand U20387 (N_20387,N_14255,N_14719);
and U20388 (N_20388,N_15289,N_14551);
nor U20389 (N_20389,N_16060,N_16844);
nand U20390 (N_20390,N_18092,N_15807);
and U20391 (N_20391,N_18265,N_15435);
nor U20392 (N_20392,N_16122,N_14524);
and U20393 (N_20393,N_16858,N_17251);
nand U20394 (N_20394,N_12876,N_13885);
and U20395 (N_20395,N_13367,N_17524);
or U20396 (N_20396,N_13956,N_18558);
and U20397 (N_20397,N_15604,N_15889);
or U20398 (N_20398,N_16923,N_18047);
nand U20399 (N_20399,N_14881,N_17027);
nor U20400 (N_20400,N_16683,N_14637);
nor U20401 (N_20401,N_14783,N_14656);
nor U20402 (N_20402,N_15916,N_16230);
or U20403 (N_20403,N_15158,N_13031);
and U20404 (N_20404,N_17059,N_18617);
and U20405 (N_20405,N_14676,N_16845);
xor U20406 (N_20406,N_13460,N_18583);
nand U20407 (N_20407,N_15461,N_17718);
xnor U20408 (N_20408,N_16025,N_17473);
or U20409 (N_20409,N_16773,N_14733);
nor U20410 (N_20410,N_12512,N_17086);
xnor U20411 (N_20411,N_15266,N_13422);
nand U20412 (N_20412,N_13294,N_17785);
and U20413 (N_20413,N_18203,N_15089);
nor U20414 (N_20414,N_16925,N_12513);
or U20415 (N_20415,N_14617,N_15363);
nor U20416 (N_20416,N_15622,N_17821);
nand U20417 (N_20417,N_12604,N_13021);
nor U20418 (N_20418,N_14533,N_13499);
or U20419 (N_20419,N_15685,N_13450);
nor U20420 (N_20420,N_12910,N_18252);
or U20421 (N_20421,N_18566,N_14329);
and U20422 (N_20422,N_15518,N_12753);
or U20423 (N_20423,N_17974,N_12884);
and U20424 (N_20424,N_13278,N_12597);
nand U20425 (N_20425,N_17307,N_14974);
and U20426 (N_20426,N_13714,N_15229);
and U20427 (N_20427,N_17209,N_13268);
nand U20428 (N_20428,N_14684,N_17431);
and U20429 (N_20429,N_15341,N_15995);
and U20430 (N_20430,N_18364,N_17442);
or U20431 (N_20431,N_18121,N_15200);
xnor U20432 (N_20432,N_13184,N_14252);
nand U20433 (N_20433,N_13232,N_18030);
nand U20434 (N_20434,N_13486,N_18543);
or U20435 (N_20435,N_15994,N_13673);
nor U20436 (N_20436,N_18677,N_15971);
nand U20437 (N_20437,N_18465,N_15066);
and U20438 (N_20438,N_14570,N_12788);
nand U20439 (N_20439,N_16139,N_16529);
nand U20440 (N_20440,N_14425,N_17725);
and U20441 (N_20441,N_13768,N_16699);
and U20442 (N_20442,N_13751,N_18105);
or U20443 (N_20443,N_13505,N_15097);
or U20444 (N_20444,N_17804,N_16494);
or U20445 (N_20445,N_14286,N_15876);
or U20446 (N_20446,N_16931,N_17406);
or U20447 (N_20447,N_16245,N_13864);
or U20448 (N_20448,N_14765,N_14363);
and U20449 (N_20449,N_17322,N_15356);
and U20450 (N_20450,N_15532,N_12573);
and U20451 (N_20451,N_13528,N_17538);
or U20452 (N_20452,N_13712,N_17295);
nor U20453 (N_20453,N_12633,N_16086);
and U20454 (N_20454,N_14663,N_13412);
nor U20455 (N_20455,N_18445,N_13749);
nand U20456 (N_20456,N_18686,N_18485);
nor U20457 (N_20457,N_17670,N_16401);
and U20458 (N_20458,N_13471,N_15436);
nor U20459 (N_20459,N_12601,N_16737);
or U20460 (N_20460,N_15687,N_16993);
and U20461 (N_20461,N_17782,N_14629);
nor U20462 (N_20462,N_13034,N_15901);
and U20463 (N_20463,N_13020,N_15554);
nand U20464 (N_20464,N_17008,N_13036);
nor U20465 (N_20465,N_17035,N_13256);
nor U20466 (N_20466,N_13841,N_15749);
or U20467 (N_20467,N_12638,N_13693);
nand U20468 (N_20468,N_16170,N_15654);
or U20469 (N_20469,N_13477,N_17282);
and U20470 (N_20470,N_12806,N_15959);
and U20471 (N_20471,N_17945,N_14445);
nand U20472 (N_20472,N_18738,N_14361);
or U20473 (N_20473,N_16029,N_17111);
nor U20474 (N_20474,N_18515,N_15057);
and U20475 (N_20475,N_18022,N_15755);
or U20476 (N_20476,N_16580,N_15095);
nand U20477 (N_20477,N_16264,N_17560);
nor U20478 (N_20478,N_13122,N_16270);
nor U20479 (N_20479,N_13663,N_17387);
nand U20480 (N_20480,N_15944,N_17926);
or U20481 (N_20481,N_16259,N_14976);
or U20482 (N_20482,N_15753,N_14155);
or U20483 (N_20483,N_17402,N_18579);
nand U20484 (N_20484,N_18582,N_13651);
or U20485 (N_20485,N_14757,N_18150);
and U20486 (N_20486,N_14005,N_16366);
nand U20487 (N_20487,N_14609,N_12855);
and U20488 (N_20488,N_14714,N_15263);
and U20489 (N_20489,N_14010,N_18299);
and U20490 (N_20490,N_12691,N_14867);
and U20491 (N_20491,N_15712,N_18615);
or U20492 (N_20492,N_13840,N_17788);
or U20493 (N_20493,N_13734,N_18161);
nand U20494 (N_20494,N_18481,N_16161);
and U20495 (N_20495,N_12819,N_18227);
xor U20496 (N_20496,N_13415,N_17452);
nor U20497 (N_20497,N_13431,N_13427);
and U20498 (N_20498,N_17211,N_17312);
nor U20499 (N_20499,N_17698,N_16714);
or U20500 (N_20500,N_15473,N_15099);
nor U20501 (N_20501,N_14024,N_17188);
nand U20502 (N_20502,N_14744,N_12528);
or U20503 (N_20503,N_13964,N_17712);
and U20504 (N_20504,N_16057,N_18304);
nand U20505 (N_20505,N_16730,N_14224);
nand U20506 (N_20506,N_17227,N_18308);
nor U20507 (N_20507,N_14021,N_18732);
nor U20508 (N_20508,N_15849,N_17694);
nor U20509 (N_20509,N_12705,N_17336);
nor U20510 (N_20510,N_13545,N_16534);
and U20511 (N_20511,N_17140,N_12593);
or U20512 (N_20512,N_13520,N_14616);
or U20513 (N_20513,N_15071,N_15040);
xor U20514 (N_20514,N_17873,N_17661);
and U20515 (N_20515,N_15746,N_14330);
nor U20516 (N_20516,N_17744,N_17236);
nor U20517 (N_20517,N_15481,N_18072);
or U20518 (N_20518,N_12672,N_12582);
and U20519 (N_20519,N_15214,N_15815);
or U20520 (N_20520,N_15046,N_18523);
nor U20521 (N_20521,N_12831,N_13295);
nand U20522 (N_20522,N_17646,N_13398);
and U20523 (N_20523,N_17588,N_16770);
nand U20524 (N_20524,N_14711,N_17171);
nand U20525 (N_20525,N_15546,N_15339);
nand U20526 (N_20526,N_12591,N_17242);
or U20527 (N_20527,N_16825,N_16249);
and U20528 (N_20528,N_15806,N_17091);
or U20529 (N_20529,N_13080,N_14746);
and U20530 (N_20530,N_15947,N_15784);
and U20531 (N_20531,N_15449,N_12612);
nand U20532 (N_20532,N_13875,N_18039);
xor U20533 (N_20533,N_17331,N_15949);
xnor U20534 (N_20534,N_15646,N_16702);
nor U20535 (N_20535,N_17980,N_16646);
nand U20536 (N_20536,N_15319,N_16981);
xor U20537 (N_20537,N_15383,N_15825);
and U20538 (N_20538,N_15962,N_17884);
nand U20539 (N_20539,N_18493,N_14284);
or U20540 (N_20540,N_18065,N_17459);
and U20541 (N_20541,N_18671,N_12507);
xnor U20542 (N_20542,N_16963,N_17969);
and U20543 (N_20543,N_16134,N_16685);
or U20544 (N_20544,N_13045,N_15881);
nand U20545 (N_20545,N_13091,N_18126);
nand U20546 (N_20546,N_16332,N_13819);
and U20547 (N_20547,N_16403,N_18552);
or U20548 (N_20548,N_17258,N_16809);
or U20549 (N_20549,N_16813,N_14275);
nand U20550 (N_20550,N_17920,N_14841);
nand U20551 (N_20551,N_14156,N_13633);
nand U20552 (N_20552,N_16932,N_13279);
nor U20553 (N_20553,N_13861,N_16413);
and U20554 (N_20554,N_12533,N_14905);
or U20555 (N_20555,N_17315,N_14368);
or U20556 (N_20556,N_15210,N_17310);
or U20557 (N_20557,N_13086,N_18005);
and U20558 (N_20558,N_16612,N_12859);
nor U20559 (N_20559,N_14394,N_18202);
nand U20560 (N_20560,N_14864,N_17051);
nand U20561 (N_20561,N_18452,N_16322);
and U20562 (N_20562,N_15163,N_16153);
xor U20563 (N_20563,N_17903,N_14163);
or U20564 (N_20564,N_17498,N_13613);
nand U20565 (N_20565,N_14958,N_12563);
nand U20566 (N_20566,N_14022,N_15765);
and U20567 (N_20567,N_15923,N_15249);
and U20568 (N_20568,N_18632,N_13708);
nand U20569 (N_20569,N_14055,N_17415);
nor U20570 (N_20570,N_13009,N_17153);
and U20571 (N_20571,N_14210,N_13747);
xor U20572 (N_20572,N_14720,N_15331);
or U20573 (N_20573,N_18131,N_14685);
nor U20574 (N_20574,N_15144,N_16627);
and U20575 (N_20575,N_17025,N_15349);
nor U20576 (N_20576,N_16841,N_14529);
nor U20577 (N_20577,N_16473,N_18069);
nand U20578 (N_20578,N_18164,N_18474);
nor U20579 (N_20579,N_17109,N_17283);
and U20580 (N_20580,N_15484,N_13452);
or U20581 (N_20581,N_13745,N_18300);
nor U20582 (N_20582,N_12603,N_12778);
or U20583 (N_20583,N_14186,N_16290);
or U20584 (N_20584,N_14148,N_13047);
xnor U20585 (N_20585,N_16624,N_16921);
nor U20586 (N_20586,N_15592,N_13903);
or U20587 (N_20587,N_18275,N_16387);
and U20588 (N_20588,N_15458,N_15088);
or U20589 (N_20589,N_14750,N_14816);
nor U20590 (N_20590,N_14346,N_16567);
xnor U20591 (N_20591,N_16926,N_17742);
nand U20592 (N_20592,N_13277,N_15886);
or U20593 (N_20593,N_17930,N_14849);
nand U20594 (N_20594,N_16085,N_17914);
and U20595 (N_20595,N_12606,N_16979);
or U20596 (N_20596,N_15766,N_15583);
xnor U20597 (N_20597,N_14219,N_16613);
nor U20598 (N_20598,N_12628,N_14139);
nand U20599 (N_20599,N_17923,N_14782);
or U20600 (N_20600,N_18743,N_14266);
nor U20601 (N_20601,N_18074,N_18424);
nand U20602 (N_20602,N_16141,N_18664);
nand U20603 (N_20603,N_18676,N_15256);
and U20604 (N_20604,N_18433,N_12780);
and U20605 (N_20605,N_16827,N_15605);
or U20606 (N_20606,N_18602,N_17202);
nor U20607 (N_20607,N_18032,N_17734);
nor U20608 (N_20608,N_14975,N_16742);
and U20609 (N_20609,N_17762,N_12811);
nor U20610 (N_20610,N_15979,N_16604);
nor U20611 (N_20611,N_16754,N_16784);
or U20612 (N_20612,N_18293,N_17398);
xor U20613 (N_20613,N_15407,N_17955);
nor U20614 (N_20614,N_15156,N_12739);
xor U20615 (N_20615,N_16950,N_18353);
nor U20616 (N_20616,N_15878,N_14183);
nand U20617 (N_20617,N_18374,N_12549);
nor U20618 (N_20618,N_15002,N_16402);
nand U20619 (N_20619,N_15345,N_18725);
and U20620 (N_20620,N_17904,N_12860);
xnor U20621 (N_20621,N_14824,N_17713);
nand U20622 (N_20622,N_14876,N_13107);
nand U20623 (N_20623,N_15003,N_17309);
xor U20624 (N_20624,N_15238,N_17680);
and U20625 (N_20625,N_16769,N_14861);
or U20626 (N_20626,N_13586,N_13612);
nor U20627 (N_20627,N_15360,N_16660);
nand U20628 (N_20628,N_17247,N_12908);
nand U20629 (N_20629,N_13070,N_13194);
or U20630 (N_20630,N_15227,N_17702);
nand U20631 (N_20631,N_16018,N_18253);
and U20632 (N_20632,N_15912,N_15008);
nor U20633 (N_20633,N_17031,N_12807);
nor U20634 (N_20634,N_18574,N_16380);
nand U20635 (N_20635,N_13766,N_13116);
and U20636 (N_20636,N_16202,N_17688);
or U20637 (N_20637,N_15762,N_16752);
and U20638 (N_20638,N_16911,N_16790);
or U20639 (N_20639,N_14644,N_16320);
or U20640 (N_20640,N_17112,N_13918);
and U20641 (N_20641,N_13200,N_15735);
nand U20642 (N_20642,N_12929,N_15929);
nand U20643 (N_20643,N_13926,N_16269);
nor U20644 (N_20644,N_14805,N_14165);
and U20645 (N_20645,N_13419,N_16389);
or U20646 (N_20646,N_13729,N_12785);
nor U20647 (N_20647,N_17262,N_14494);
or U20648 (N_20648,N_14774,N_18207);
and U20649 (N_20649,N_14396,N_17380);
and U20650 (N_20650,N_17403,N_13428);
nor U20651 (N_20651,N_18730,N_16916);
nand U20652 (N_20652,N_18217,N_14990);
or U20653 (N_20653,N_17906,N_14604);
nand U20654 (N_20654,N_14250,N_15185);
nand U20655 (N_20655,N_16223,N_17676);
nand U20656 (N_20656,N_17478,N_14270);
or U20657 (N_20657,N_17848,N_12887);
or U20658 (N_20658,N_12553,N_18383);
or U20659 (N_20659,N_17783,N_15019);
nand U20660 (N_20660,N_16895,N_13183);
and U20661 (N_20661,N_17409,N_15242);
xnor U20662 (N_20662,N_18547,N_15706);
nand U20663 (N_20663,N_14934,N_12600);
nor U20664 (N_20664,N_18077,N_13608);
nor U20665 (N_20665,N_12805,N_15208);
nand U20666 (N_20666,N_14283,N_14843);
or U20667 (N_20667,N_13552,N_17545);
and U20668 (N_20668,N_16441,N_16501);
nand U20669 (N_20669,N_17992,N_12712);
nand U20670 (N_20670,N_16016,N_14879);
or U20671 (N_20671,N_14837,N_13945);
xor U20672 (N_20672,N_13598,N_13443);
nor U20673 (N_20673,N_16111,N_18139);
and U20674 (N_20674,N_16083,N_15862);
nor U20675 (N_20675,N_18100,N_15273);
or U20676 (N_20676,N_17193,N_16006);
and U20677 (N_20677,N_18043,N_17032);
nand U20678 (N_20678,N_13158,N_15190);
nand U20679 (N_20679,N_14574,N_13274);
and U20680 (N_20680,N_17526,N_14474);
and U20681 (N_20681,N_17689,N_14796);
and U20682 (N_20682,N_17483,N_17595);
or U20683 (N_20683,N_14349,N_18713);
nand U20684 (N_20684,N_14887,N_15847);
and U20685 (N_20685,N_12568,N_15620);
and U20686 (N_20686,N_18233,N_17582);
nand U20687 (N_20687,N_17956,N_17709);
nor U20688 (N_20688,N_12997,N_16334);
xor U20689 (N_20689,N_17317,N_15917);
nand U20690 (N_20690,N_18255,N_17660);
and U20691 (N_20691,N_18628,N_14810);
and U20692 (N_20692,N_16945,N_15188);
and U20693 (N_20693,N_17280,N_17876);
and U20694 (N_20694,N_16192,N_14499);
nand U20695 (N_20695,N_15248,N_17864);
and U20696 (N_20696,N_14076,N_14591);
nand U20697 (N_20697,N_15107,N_14102);
nand U20698 (N_20698,N_15338,N_16056);
or U20699 (N_20699,N_18250,N_18018);
or U20700 (N_20700,N_17730,N_14963);
and U20701 (N_20701,N_18085,N_12922);
nor U20702 (N_20702,N_14726,N_15918);
nand U20703 (N_20703,N_15709,N_12661);
nor U20704 (N_20704,N_16630,N_12933);
nor U20705 (N_20705,N_15157,N_17697);
nor U20706 (N_20706,N_17623,N_16878);
or U20707 (N_20707,N_17401,N_16749);
nor U20708 (N_20708,N_17038,N_12869);
xnor U20709 (N_20709,N_17163,N_16216);
nor U20710 (N_20710,N_17629,N_17586);
or U20711 (N_20711,N_14468,N_16062);
and U20712 (N_20712,N_17328,N_15946);
or U20713 (N_20713,N_13541,N_15112);
nor U20714 (N_20714,N_16937,N_16009);
nand U20715 (N_20715,N_16853,N_13786);
nand U20716 (N_20716,N_14538,N_12957);
or U20717 (N_20717,N_15742,N_18675);
nand U20718 (N_20718,N_14011,N_17502);
nand U20719 (N_20719,N_16920,N_14598);
nor U20720 (N_20720,N_13003,N_14218);
xor U20721 (N_20721,N_15025,N_13495);
nand U20722 (N_20722,N_12818,N_15243);
and U20723 (N_20723,N_17612,N_15454);
or U20724 (N_20724,N_18064,N_18246);
xnor U20725 (N_20725,N_16669,N_15548);
or U20726 (N_20726,N_16917,N_15051);
and U20727 (N_20727,N_18405,N_18086);
nor U20728 (N_20728,N_14953,N_13453);
nand U20729 (N_20729,N_18099,N_17519);
nand U20730 (N_20730,N_14846,N_13181);
and U20731 (N_20731,N_15977,N_13044);
or U20732 (N_20732,N_14491,N_13321);
and U20733 (N_20733,N_16115,N_14563);
and U20734 (N_20734,N_16004,N_14911);
nand U20735 (N_20735,N_13981,N_15313);
nor U20736 (N_20736,N_17172,N_13163);
and U20737 (N_20737,N_18156,N_18171);
nand U20738 (N_20738,N_17932,N_17724);
and U20739 (N_20739,N_12524,N_18002);
and U20740 (N_20740,N_14209,N_15209);
xor U20741 (N_20741,N_18548,N_13716);
nor U20742 (N_20742,N_18638,N_15669);
nor U20743 (N_20743,N_18313,N_17208);
nand U20744 (N_20744,N_17799,N_16989);
and U20745 (N_20745,N_14756,N_13331);
xor U20746 (N_20746,N_12667,N_18208);
and U20747 (N_20747,N_13303,N_17147);
or U20748 (N_20748,N_14970,N_13748);
or U20749 (N_20749,N_17879,N_14229);
and U20750 (N_20750,N_18407,N_15191);
nand U20751 (N_20751,N_15154,N_16298);
nor U20752 (N_20752,N_12548,N_18205);
or U20753 (N_20753,N_12742,N_14057);
nor U20754 (N_20754,N_12558,N_17774);
xnor U20755 (N_20755,N_15267,N_15224);
nor U20756 (N_20756,N_15741,N_14633);
xnor U20757 (N_20757,N_13041,N_16028);
nand U20758 (N_20758,N_16560,N_12934);
or U20759 (N_20759,N_18438,N_16052);
nand U20760 (N_20760,N_12830,N_16735);
nor U20761 (N_20761,N_14212,N_15769);
nor U20762 (N_20762,N_18231,N_13624);
nand U20763 (N_20763,N_14745,N_18209);
nor U20764 (N_20764,N_12817,N_13515);
nor U20765 (N_20765,N_18682,N_17836);
or U20766 (N_20766,N_15938,N_15127);
xor U20767 (N_20767,N_13883,N_17237);
nand U20768 (N_20768,N_16513,N_16040);
or U20769 (N_20769,N_15409,N_15630);
and U20770 (N_20770,N_14868,N_16674);
nand U20771 (N_20771,N_17314,N_12808);
and U20772 (N_20772,N_13848,N_17271);
or U20773 (N_20773,N_15311,N_17245);
and U20774 (N_20774,N_15070,N_13822);
nand U20775 (N_20775,N_12854,N_12812);
xnor U20776 (N_20776,N_16631,N_14457);
nand U20777 (N_20777,N_14518,N_16535);
nor U20778 (N_20778,N_18584,N_18718);
xnor U20779 (N_20779,N_18717,N_17705);
or U20780 (N_20780,N_17967,N_18681);
and U20781 (N_20781,N_14576,N_12559);
xnor U20782 (N_20782,N_14855,N_17175);
nand U20783 (N_20783,N_17865,N_18573);
and U20784 (N_20784,N_12856,N_18095);
or U20785 (N_20785,N_18152,N_18661);
or U20786 (N_20786,N_16395,N_18175);
nand U20787 (N_20787,N_14247,N_15036);
or U20788 (N_20788,N_14233,N_12963);
xnor U20789 (N_20789,N_12943,N_15803);
and U20790 (N_20790,N_17824,N_15265);
and U20791 (N_20791,N_17572,N_15045);
nand U20792 (N_20792,N_17562,N_18640);
or U20793 (N_20793,N_18168,N_17861);
nor U20794 (N_20794,N_15448,N_16278);
nor U20795 (N_20795,N_15149,N_18279);
nor U20796 (N_20796,N_12501,N_14014);
or U20797 (N_20797,N_16570,N_12555);
nand U20798 (N_20798,N_12595,N_15034);
or U20799 (N_20799,N_14540,N_18699);
and U20800 (N_20800,N_16277,N_16710);
xnor U20801 (N_20801,N_15814,N_12849);
nor U20802 (N_20802,N_15054,N_18537);
nand U20803 (N_20803,N_13971,N_14527);
and U20804 (N_20804,N_14566,N_12993);
or U20805 (N_20805,N_15295,N_17703);
and U20806 (N_20806,N_15729,N_18704);
nand U20807 (N_20807,N_18371,N_14293);
and U20808 (N_20808,N_18590,N_14176);
nor U20809 (N_20809,N_14691,N_13834);
and U20810 (N_20810,N_13892,N_16280);
and U20811 (N_20811,N_16946,N_13456);
nor U20812 (N_20812,N_16281,N_14147);
or U20813 (N_20813,N_17152,N_12942);
and U20814 (N_20814,N_18071,N_16821);
xnor U20815 (N_20815,N_14372,N_13289);
nand U20816 (N_20816,N_17270,N_15832);
and U20817 (N_20817,N_17888,N_12879);
and U20818 (N_20818,N_14311,N_13655);
xnor U20819 (N_20819,N_18091,N_16341);
nor U20820 (N_20820,N_14991,N_15362);
and U20821 (N_20821,N_15992,N_18553);
nor U20822 (N_20822,N_18495,N_15507);
nand U20823 (N_20823,N_14094,N_18117);
or U20824 (N_20824,N_16154,N_13121);
or U20825 (N_20825,N_16708,N_15386);
nor U20826 (N_20826,N_15642,N_15368);
and U20827 (N_20827,N_13399,N_16743);
or U20828 (N_20828,N_16397,N_16187);
or U20829 (N_20829,N_17268,N_17539);
nand U20830 (N_20830,N_16117,N_13965);
nor U20831 (N_20831,N_16603,N_13072);
and U20832 (N_20832,N_13058,N_18186);
nor U20833 (N_20833,N_16751,N_13455);
nor U20834 (N_20834,N_17727,N_14674);
and U20835 (N_20835,N_16540,N_15219);
and U20836 (N_20836,N_17751,N_14528);
or U20837 (N_20837,N_13592,N_17826);
nor U20838 (N_20838,N_13053,N_14288);
xor U20839 (N_20839,N_13377,N_13761);
and U20840 (N_20840,N_12720,N_16024);
nor U20841 (N_20841,N_13526,N_15613);
or U20842 (N_20842,N_16665,N_17206);
or U20843 (N_20843,N_13817,N_14149);
or U20844 (N_20844,N_14503,N_13081);
nor U20845 (N_20845,N_16868,N_15593);
nor U20846 (N_20846,N_15655,N_18332);
and U20847 (N_20847,N_16798,N_14817);
and U20848 (N_20848,N_17801,N_15714);
or U20849 (N_20849,N_13114,N_18429);
nand U20850 (N_20850,N_16221,N_16211);
nand U20851 (N_20851,N_16113,N_15298);
and U20852 (N_20852,N_17076,N_13266);
nor U20853 (N_20853,N_12793,N_17354);
and U20854 (N_20854,N_16391,N_16054);
or U20855 (N_20855,N_16620,N_17870);
and U20856 (N_20856,N_16015,N_17793);
nor U20857 (N_20857,N_14390,N_14839);
or U20858 (N_20858,N_13548,N_14345);
nor U20859 (N_20859,N_15908,N_17480);
or U20860 (N_20860,N_16044,N_15141);
xor U20861 (N_20861,N_17523,N_16434);
and U20862 (N_20862,N_18155,N_14625);
nand U20863 (N_20863,N_16792,N_14140);
xnor U20864 (N_20864,N_16789,N_16522);
and U20865 (N_20865,N_15608,N_17897);
nand U20866 (N_20866,N_12918,N_16915);
xnor U20867 (N_20867,N_14404,N_12978);
nand U20868 (N_20868,N_16954,N_13554);
and U20869 (N_20869,N_14410,N_13315);
and U20870 (N_20870,N_15796,N_15294);
nand U20871 (N_20871,N_16721,N_18266);
xor U20872 (N_20872,N_15582,N_13635);
nor U20873 (N_20873,N_16142,N_13979);
nand U20874 (N_20874,N_14444,N_16023);
nor U20875 (N_20875,N_16820,N_16514);
nor U20876 (N_20876,N_17795,N_17675);
xor U20877 (N_20877,N_13478,N_17650);
and U20878 (N_20878,N_16537,N_18420);
nand U20879 (N_20879,N_15958,N_15447);
nand U20880 (N_20880,N_15451,N_17451);
and U20881 (N_20881,N_16313,N_17528);
and U20882 (N_20882,N_13763,N_17129);
nor U20883 (N_20883,N_14670,N_15446);
nand U20884 (N_20884,N_16013,N_13156);
or U20885 (N_20885,N_18158,N_13126);
nor U20886 (N_20886,N_13386,N_15895);
or U20887 (N_20887,N_13498,N_16938);
or U20888 (N_20888,N_13715,N_13695);
nor U20889 (N_20889,N_17358,N_13963);
nand U20890 (N_20890,N_18453,N_17991);
and U20891 (N_20891,N_12873,N_18700);
and U20892 (N_20892,N_17877,N_15701);
or U20893 (N_20893,N_14016,N_16899);
nand U20894 (N_20894,N_14891,N_18341);
nor U20895 (N_20895,N_15691,N_16733);
and U20896 (N_20896,N_16361,N_17743);
xnor U20897 (N_20897,N_15828,N_17014);
nand U20898 (N_20898,N_14724,N_18123);
and U20899 (N_20899,N_16412,N_18387);
and U20900 (N_20900,N_15675,N_15750);
nand U20901 (N_20901,N_14202,N_16452);
or U20902 (N_20902,N_16569,N_14080);
nand U20903 (N_20903,N_13575,N_18516);
and U20904 (N_20904,N_15491,N_16690);
and U20905 (N_20905,N_13839,N_17467);
and U20906 (N_20906,N_14987,N_14274);
or U20907 (N_20907,N_14550,N_12587);
nor U20908 (N_20908,N_16423,N_15758);
nand U20909 (N_20909,N_18492,N_13188);
and U20910 (N_20910,N_14761,N_17704);
nand U20911 (N_20911,N_16324,N_15930);
or U20912 (N_20912,N_15570,N_14580);
nor U20913 (N_20913,N_18443,N_13492);
nor U20914 (N_20914,N_18585,N_17143);
or U20915 (N_20915,N_16125,N_13094);
and U20916 (N_20916,N_13191,N_15466);
nor U20917 (N_20917,N_16539,N_16226);
xor U20918 (N_20918,N_14647,N_15920);
or U20919 (N_20919,N_17477,N_13692);
nand U20920 (N_20920,N_17238,N_17488);
xor U20921 (N_20921,N_14401,N_16734);
or U20922 (N_20922,N_18144,N_18428);
nor U20923 (N_20923,N_16574,N_15444);
and U20924 (N_20924,N_15080,N_16745);
or U20925 (N_20925,N_17910,N_16936);
xor U20926 (N_20926,N_13927,N_17419);
nand U20927 (N_20927,N_18694,N_18141);
nand U20928 (N_20928,N_15863,N_17160);
or U20929 (N_20929,N_14665,N_13832);
nand U20930 (N_20930,N_16778,N_15515);
nand U20931 (N_20931,N_13287,N_13083);
and U20932 (N_20932,N_13390,N_17180);
or U20933 (N_20933,N_14535,N_13265);
nand U20934 (N_20934,N_16103,N_16622);
nand U20935 (N_20935,N_18016,N_17659);
xor U20936 (N_20936,N_18721,N_16549);
and U20937 (N_20937,N_14453,N_12932);
nand U20938 (N_20938,N_17892,N_17815);
nand U20939 (N_20939,N_13632,N_12898);
or U20940 (N_20940,N_17757,N_17464);
and U20941 (N_20941,N_15493,N_17627);
nor U20942 (N_20942,N_17288,N_17301);
nor U20943 (N_20943,N_13285,N_16507);
nor U20944 (N_20944,N_13579,N_17134);
xor U20945 (N_20945,N_16695,N_14152);
and U20946 (N_20946,N_16343,N_13596);
or U20947 (N_20947,N_17537,N_18434);
xor U20948 (N_20948,N_18595,N_14519);
nor U20949 (N_20949,N_17949,N_17357);
or U20950 (N_20950,N_14512,N_15124);
xor U20951 (N_20951,N_17297,N_15197);
nand U20952 (N_20952,N_16753,N_16171);
and U20953 (N_20953,N_14682,N_14722);
nor U20954 (N_20954,N_15978,N_15485);
or U20955 (N_20955,N_18630,N_15933);
xnor U20956 (N_20956,N_16776,N_18478);
nor U20957 (N_20957,N_14114,N_17418);
nor U20958 (N_20958,N_13433,N_13322);
nand U20959 (N_20959,N_13179,N_15780);
or U20960 (N_20960,N_18648,N_17696);
nor U20961 (N_20961,N_16572,N_12758);
xor U20962 (N_20962,N_15875,N_16512);
nand U20963 (N_20963,N_17441,N_17850);
and U20964 (N_20964,N_18525,N_16818);
or U20965 (N_20965,N_15388,N_18358);
or U20966 (N_20966,N_17700,N_16065);
nor U20967 (N_20967,N_15310,N_16096);
or U20968 (N_20968,N_17869,N_17909);
or U20969 (N_20969,N_13953,N_14254);
nand U20970 (N_20970,N_14752,N_13097);
nor U20971 (N_20971,N_12611,N_15793);
or U20972 (N_20972,N_15914,N_16589);
and U20973 (N_20973,N_13777,N_13226);
and U20974 (N_20974,N_12981,N_14442);
xnor U20975 (N_20975,N_17971,N_13352);
and U20976 (N_20976,N_15804,N_15898);
and U20977 (N_20977,N_13185,N_14258);
and U20978 (N_20978,N_13877,N_12877);
nor U20979 (N_20979,N_17494,N_18678);
nor U20980 (N_20980,N_15989,N_16849);
nor U20981 (N_20981,N_14047,N_16651);
xor U20982 (N_20982,N_17533,N_17164);
or U20983 (N_20983,N_12567,N_14807);
xnor U20984 (N_20984,N_13703,N_13148);
xor U20985 (N_20985,N_14689,N_16155);
or U20986 (N_20986,N_13825,N_14708);
and U20987 (N_20987,N_14997,N_15410);
nand U20988 (N_20988,N_13146,N_14883);
xor U20989 (N_20989,N_14493,N_13913);
and U20990 (N_20990,N_18555,N_17492);
nand U20991 (N_20991,N_13741,N_15182);
nor U20992 (N_20992,N_17965,N_13961);
nand U20993 (N_20993,N_12904,N_12915);
or U20994 (N_20994,N_18587,N_15921);
nand U20995 (N_20995,N_13395,N_15252);
or U20996 (N_20996,N_14786,N_18087);
or U20997 (N_20997,N_16562,N_18683);
or U20998 (N_20998,N_15184,N_13513);
or U20999 (N_20999,N_17619,N_15586);
and U21000 (N_21000,N_14942,N_13670);
and U21001 (N_21001,N_15469,N_13544);
and U21002 (N_21002,N_17554,N_16002);
nor U21003 (N_21003,N_13136,N_18690);
xor U21004 (N_21004,N_15589,N_18003);
and U21005 (N_21005,N_14307,N_17972);
nand U21006 (N_21006,N_12623,N_12998);
and U21007 (N_21007,N_13383,N_17733);
xor U21008 (N_21008,N_18570,N_13317);
nand U21009 (N_21009,N_13313,N_15527);
nand U21010 (N_21010,N_17161,N_14941);
nor U21011 (N_21011,N_15924,N_17886);
and U21012 (N_21012,N_17657,N_14827);
xnor U21013 (N_21013,N_15336,N_13166);
and U21014 (N_21014,N_13897,N_14555);
or U21015 (N_21015,N_14000,N_13077);
nand U21016 (N_21016,N_18167,N_17846);
nor U21017 (N_21017,N_17162,N_15456);
nand U21018 (N_21018,N_13807,N_14652);
and U21019 (N_21019,N_14195,N_12736);
nor U21020 (N_21020,N_15395,N_18666);
nand U21021 (N_21021,N_14455,N_12550);
xnor U21022 (N_21022,N_15647,N_13646);
or U21023 (N_21023,N_15531,N_17761);
nand U21024 (N_21024,N_18501,N_15653);
nor U21025 (N_21025,N_17747,N_12903);
nand U21026 (N_21026,N_14678,N_13788);
xor U21027 (N_21027,N_14593,N_17777);
nand U21028 (N_21028,N_17752,N_17515);
or U21029 (N_21029,N_14603,N_18287);
or U21030 (N_21030,N_17552,N_16644);
nor U21031 (N_21031,N_15730,N_17532);
or U21032 (N_21032,N_14428,N_15633);
and U21033 (N_21033,N_14002,N_17338);
nor U21034 (N_21034,N_17115,N_15838);
nand U21035 (N_21035,N_14244,N_15325);
nor U21036 (N_21036,N_15475,N_14043);
or U21037 (N_21037,N_18237,N_16573);
or U21038 (N_21038,N_18747,N_18672);
nor U21039 (N_21039,N_18355,N_17715);
and U21040 (N_21040,N_13869,N_15078);
and U21041 (N_21041,N_13159,N_16459);
nor U21042 (N_21042,N_14740,N_15726);
or U21043 (N_21043,N_17816,N_14100);
and U21044 (N_21044,N_16564,N_17773);
and U21045 (N_21045,N_15361,N_14717);
nand U21046 (N_21046,N_17150,N_14313);
nand U21047 (N_21047,N_14779,N_16703);
nor U21048 (N_21048,N_17466,N_18505);
nand U21049 (N_21049,N_14465,N_16306);
nand U21050 (N_21050,N_14832,N_13601);
xor U21051 (N_21051,N_17016,N_13576);
nor U21052 (N_21052,N_17170,N_14459);
xnor U21053 (N_21053,N_17344,N_16558);
or U21054 (N_21054,N_16596,N_12979);
or U21055 (N_21055,N_13906,N_15906);
nand U21056 (N_21056,N_17985,N_15109);
and U21057 (N_21057,N_13684,N_15573);
or U21058 (N_21058,N_16179,N_14657);
nand U21059 (N_21059,N_14646,N_16958);
and U21060 (N_21060,N_15302,N_15760);
nand U21061 (N_21061,N_16252,N_13561);
nand U21062 (N_21062,N_12684,N_12656);
and U21063 (N_21063,N_17287,N_13676);
nor U21064 (N_21064,N_14773,N_18014);
nand U21065 (N_21065,N_18184,N_18103);
or U21066 (N_21066,N_13110,N_14120);
and U21067 (N_21067,N_15411,N_14223);
and U21068 (N_21068,N_16793,N_15186);
nor U21069 (N_21069,N_15517,N_12531);
xor U21070 (N_21070,N_17176,N_13565);
nand U21071 (N_21071,N_18151,N_15771);
or U21072 (N_21072,N_18084,N_14602);
xor U21073 (N_21073,N_14362,N_17023);
or U21074 (N_21074,N_17797,N_12575);
and U21075 (N_21075,N_15606,N_14892);
nand U21076 (N_21076,N_14381,N_15778);
and U21077 (N_21077,N_17584,N_15911);
nand U21078 (N_21078,N_12571,N_16382);
and U21079 (N_21079,N_14322,N_18196);
nor U21080 (N_21080,N_14235,N_17695);
and U21081 (N_21081,N_13625,N_14204);
nand U21082 (N_21082,N_17082,N_12713);
nor U21083 (N_21083,N_15612,N_16026);
and U21084 (N_21084,N_13511,N_17394);
nand U21085 (N_21085,N_12654,N_17950);
or U21086 (N_21086,N_12622,N_13744);
and U21087 (N_21087,N_18303,N_14314);
nand U21088 (N_21088,N_18546,N_17034);
nand U21089 (N_21089,N_16530,N_17832);
nand U21090 (N_21090,N_17907,N_12624);
nor U21091 (N_21091,N_14851,N_15375);
xnor U21092 (N_21092,N_14956,N_15711);
xnor U21093 (N_21093,N_13362,N_14927);
nor U21094 (N_21094,N_12825,N_13500);
or U21095 (N_21095,N_15140,N_14835);
and U21096 (N_21096,N_13845,N_15151);
and U21097 (N_21097,N_14175,N_12744);
nand U21098 (N_21098,N_13142,N_12627);
nor U21099 (N_21099,N_15562,N_15564);
xnor U21100 (N_21100,N_15896,N_18122);
nand U21101 (N_21101,N_15514,N_15384);
or U21102 (N_21102,N_18116,N_15111);
nand U21103 (N_21103,N_14487,N_17320);
nand U21104 (N_21104,N_16131,N_12617);
nand U21105 (N_21105,N_16541,N_12896);
nor U21106 (N_21106,N_12529,N_16396);
nor U21107 (N_21107,N_18314,N_13914);
and U21108 (N_21108,N_15552,N_16869);
and U21109 (N_21109,N_17343,N_17699);
and U21110 (N_21110,N_17377,N_18001);
or U21111 (N_21111,N_17509,N_17931);
and U21112 (N_21112,N_16705,N_14725);
and U21113 (N_21113,N_15915,N_14610);
or U21114 (N_21114,N_17253,N_17142);
or U21115 (N_21115,N_15268,N_14702);
nand U21116 (N_21116,N_15380,N_18724);
nand U21117 (N_21117,N_14838,N_15176);
nand U21118 (N_21118,N_16138,N_13645);
or U21119 (N_21119,N_12662,N_16667);
xnor U21120 (N_21120,N_13361,N_16959);
nand U21121 (N_21121,N_12962,N_13199);
or U21122 (N_21122,N_12813,N_17921);
and U21123 (N_21123,N_16952,N_14873);
or U21124 (N_21124,N_18119,N_18177);
nor U21125 (N_21125,N_13101,N_18431);
or U21126 (N_21126,N_14225,N_14471);
and U21127 (N_21127,N_16197,N_17739);
nand U21128 (N_21128,N_14915,N_17006);
and U21129 (N_21129,N_13658,N_16077);
and U21130 (N_21130,N_13459,N_14999);
nor U21131 (N_21131,N_13882,N_12885);
nand U21132 (N_21132,N_15056,N_12537);
and U21133 (N_21133,N_16208,N_16472);
or U21134 (N_21134,N_16693,N_14454);
nor U21135 (N_21135,N_15623,N_13627);
nor U21136 (N_21136,N_14589,N_18652);
nand U21137 (N_21137,N_17565,N_14579);
nor U21138 (N_21138,N_15648,N_13939);
nor U21139 (N_21139,N_17254,N_13096);
nor U21140 (N_21140,N_16254,N_16922);
and U21141 (N_21141,N_13637,N_15812);
or U21142 (N_21142,N_16586,N_14467);
nand U21143 (N_21143,N_14982,N_13669);
or U21144 (N_21144,N_18698,N_15128);
xnor U21145 (N_21145,N_16947,N_16037);
nor U21146 (N_21146,N_13345,N_13757);
nor U21147 (N_21147,N_15808,N_14303);
nand U21148 (N_21148,N_14015,N_13389);
and U21149 (N_21149,N_18224,N_18440);
or U21150 (N_21150,N_14180,N_14601);
nor U21151 (N_21151,N_15164,N_18468);
and U21152 (N_21152,N_15664,N_12843);
nor U21153 (N_21153,N_15910,N_13774);
nand U21154 (N_21154,N_15984,N_13510);
or U21155 (N_21155,N_17225,N_18518);
and U21156 (N_21156,N_15521,N_13739);
or U21157 (N_21157,N_14526,N_18414);
nand U21158 (N_21158,N_17568,N_16757);
or U21159 (N_21159,N_18143,N_16717);
nand U21160 (N_21160,N_17728,N_17440);
and U21161 (N_21161,N_16283,N_18172);
or U21162 (N_21162,N_13292,N_12967);
xnor U21163 (N_21163,N_17277,N_17154);
or U21164 (N_21164,N_15710,N_16985);
nor U21165 (N_21165,N_17458,N_17267);
nor U21166 (N_21166,N_14686,N_16326);
and U21167 (N_21167,N_12970,N_14230);
nor U21168 (N_21168,N_16011,N_14191);
xor U21169 (N_21169,N_14344,N_13713);
nor U21170 (N_21170,N_17609,N_18198);
xnor U21171 (N_21171,N_14017,N_13587);
and U21172 (N_21172,N_14133,N_12779);
nor U21173 (N_21173,N_15585,N_17731);
nor U21174 (N_21174,N_18484,N_13560);
nand U21175 (N_21175,N_14764,N_14966);
nor U21176 (N_21176,N_16542,N_13649);
xor U21177 (N_21177,N_18008,N_14009);
and U21178 (N_21178,N_14912,N_17333);
xnor U21179 (N_21179,N_17622,N_17067);
nand U21180 (N_21180,N_15101,N_14065);
xnor U21181 (N_21181,N_17128,N_18488);
and U21182 (N_21182,N_17447,N_15666);
nor U21183 (N_21183,N_14236,N_14193);
and U21184 (N_21184,N_16628,N_14759);
nor U21185 (N_21185,N_17858,N_15478);
nand U21186 (N_21186,N_14763,N_12803);
and U21187 (N_21187,N_14153,N_18511);
nor U21188 (N_21188,N_16607,N_18655);
or U21189 (N_21189,N_18560,N_18146);
xnor U21190 (N_21190,N_14073,N_12645);
nor U21191 (N_21191,N_12599,N_14801);
xnor U21192 (N_21192,N_16005,N_14813);
nand U21193 (N_21193,N_15463,N_18215);
nand U21194 (N_21194,N_17536,N_12675);
nand U21195 (N_21195,N_16308,N_18442);
or U21196 (N_21196,N_16483,N_16965);
or U21197 (N_21197,N_15081,N_12640);
or U21198 (N_21198,N_17264,N_18404);
nand U21199 (N_21199,N_13781,N_14353);
nand U21200 (N_21200,N_16799,N_18625);
nor U21201 (N_21201,N_13371,N_13517);
or U21202 (N_21202,N_15698,N_18551);
or U21203 (N_21203,N_14238,N_12986);
nor U21204 (N_21204,N_18060,N_16470);
nand U21205 (N_21205,N_13987,N_18330);
xnor U21206 (N_21206,N_18503,N_18111);
nand U21207 (N_21207,N_12850,N_14161);
xnor U21208 (N_21208,N_18643,N_13169);
or U21209 (N_21209,N_15415,N_17240);
or U21210 (N_21210,N_14870,N_15090);
nor U21211 (N_21211,N_17792,N_13711);
nor U21212 (N_21212,N_17475,N_15030);
or U21213 (N_21213,N_13373,N_14447);
or U21214 (N_21214,N_13666,N_14586);
or U21215 (N_21215,N_18024,N_12768);
or U21216 (N_21216,N_18162,N_15215);
nand U21217 (N_21217,N_17663,N_17615);
nand U21218 (N_21218,N_17613,N_17423);
nand U21219 (N_21219,N_13483,N_14008);
nand U21220 (N_21220,N_15223,N_12983);
and U21221 (N_21221,N_18411,N_18221);
or U21222 (N_21222,N_16212,N_17571);
or U21223 (N_21223,N_17900,N_17174);
nand U21224 (N_21224,N_13448,N_17470);
xnor U21225 (N_21225,N_16913,N_15632);
nand U21226 (N_21226,N_14122,N_14044);
and U21227 (N_21227,N_13647,N_16375);
or U21228 (N_21228,N_12646,N_15240);
nand U21229 (N_21229,N_16728,N_16102);
xor U21230 (N_21230,N_17671,N_13421);
nand U21231 (N_21231,N_16608,N_16551);
nor U21232 (N_21232,N_15821,N_14954);
nand U21233 (N_21233,N_17691,N_15787);
and U21234 (N_21234,N_17250,N_15085);
and U21235 (N_21235,N_17437,N_17760);
nor U21236 (N_21236,N_13064,N_12975);
and U21237 (N_21237,N_14028,N_16207);
xnor U21238 (N_21238,N_14731,N_14596);
and U21239 (N_21239,N_13919,N_15511);
or U21240 (N_21240,N_14086,N_13990);
nand U21241 (N_21241,N_15334,N_15394);
and U21242 (N_21242,N_13970,N_15988);
nand U21243 (N_21243,N_18098,N_14776);
nand U21244 (N_21244,N_17106,N_12543);
and U21245 (N_21245,N_14553,N_17600);
and U21246 (N_21246,N_16812,N_16030);
and U21247 (N_21247,N_18140,N_13689);
or U21248 (N_21248,N_17063,N_14607);
and U21249 (N_21249,N_15370,N_18413);
and U21250 (N_21250,N_15404,N_17265);
nor U21251 (N_21251,N_16796,N_13329);
nand U21252 (N_21252,N_14784,N_17569);
or U21253 (N_21253,N_13406,N_15322);
nand U21254 (N_21254,N_13874,N_17765);
and U21255 (N_21255,N_16561,N_17024);
or U21256 (N_21256,N_15376,N_13992);
or U21257 (N_21257,N_14573,N_15530);
or U21258 (N_21258,N_12714,N_16682);
and U21259 (N_21259,N_15328,N_17359);
nor U21260 (N_21260,N_18658,N_16626);
or U21261 (N_21261,N_16519,N_16409);
xor U21262 (N_21262,N_15975,N_18042);
and U21263 (N_21263,N_13849,N_14477);
nand U21264 (N_21264,N_12685,N_17970);
or U21265 (N_21265,N_12940,N_13082);
or U21266 (N_21266,N_13454,N_16716);
or U21267 (N_21267,N_16272,N_14403);
and U21268 (N_21268,N_15077,N_13218);
and U21269 (N_21269,N_13806,N_16046);
nor U21270 (N_21270,N_16101,N_14215);
nor U21271 (N_21271,N_15658,N_15038);
nand U21272 (N_21272,N_13291,N_15550);
or U21273 (N_21273,N_17624,N_17530);
or U21274 (N_21274,N_15777,N_18331);
xor U21275 (N_21275,N_16191,N_14906);
nor U21276 (N_21276,N_18388,N_13050);
nor U21277 (N_21277,N_16816,N_13683);
or U21278 (N_21278,N_13006,N_15153);
or U21279 (N_21279,N_15194,N_16385);
nor U21280 (N_21280,N_16852,N_16461);
and U21281 (N_21281,N_14480,N_14569);
and U21282 (N_21282,N_18290,N_16775);
nor U21283 (N_21283,N_15332,N_14348);
or U21284 (N_21284,N_17922,N_16715);
or U21285 (N_21285,N_13418,N_15171);
or U21286 (N_21286,N_17603,N_16594);
nand U21287 (N_21287,N_13001,N_12935);
and U21288 (N_21288,N_15591,N_15942);
nor U21289 (N_21289,N_14220,N_12596);
nor U21290 (N_21290,N_18360,N_12589);
nand U21291 (N_21291,N_17596,N_13308);
and U21292 (N_21292,N_15042,N_18102);
and U21293 (N_21293,N_14409,N_15239);
nand U21294 (N_21294,N_15794,N_14819);
xor U21295 (N_21295,N_18157,N_17548);
nand U21296 (N_21296,N_18273,N_13867);
or U21297 (N_21297,N_15122,N_15611);
xor U21298 (N_21298,N_13441,N_15116);
nor U21299 (N_21299,N_12765,N_12577);
nand U21300 (N_21300,N_12731,N_14587);
or U21301 (N_21301,N_14770,N_18107);
nand U21302 (N_21302,N_16795,N_16328);
nand U21303 (N_21303,N_13134,N_12961);
nand U21304 (N_21304,N_13302,N_15350);
nor U21305 (N_21305,N_13685,N_17404);
nand U21306 (N_21306,N_16896,N_18035);
nand U21307 (N_21307,N_15859,N_13414);
nand U21308 (N_21308,N_16907,N_13640);
nand U21309 (N_21309,N_18512,N_13827);
xor U21310 (N_21310,N_17947,N_14268);
nor U21311 (N_21311,N_17033,N_15516);
and U21312 (N_21312,N_13950,N_12584);
and U21313 (N_21313,N_16132,N_14172);
and U21314 (N_21314,N_16881,N_13850);
nor U21315 (N_21315,N_17616,N_15887);
nand U21316 (N_21316,N_18451,N_15441);
or U21317 (N_21317,N_15684,N_13949);
nand U21318 (N_21318,N_15510,N_15148);
nand U21319 (N_21319,N_15996,N_17981);
and U21320 (N_21320,N_15414,N_14259);
nor U21321 (N_21321,N_15290,N_15113);
or U21322 (N_21322,N_18734,N_13606);
and U21323 (N_21323,N_14448,N_13442);
nor U21324 (N_21324,N_16901,N_12972);
or U21325 (N_21325,N_12764,N_15134);
and U21326 (N_21326,N_17463,N_18134);
nor U21327 (N_21327,N_16864,N_17626);
nand U21328 (N_21328,N_18644,N_13547);
nor U21329 (N_21329,N_15934,N_13192);
nand U21330 (N_21330,N_18636,N_13730);
or U21331 (N_21331,N_15626,N_17640);
nor U21332 (N_21332,N_16986,N_18439);
and U21333 (N_21333,N_15179,N_16909);
and U21334 (N_21334,N_14194,N_17550);
nor U21335 (N_21335,N_16135,N_16867);
nand U21336 (N_21336,N_15417,N_13888);
nor U21337 (N_21337,N_12989,N_17050);
nand U21338 (N_21338,N_12644,N_13253);
or U21339 (N_21339,N_16338,N_14084);
nor U21340 (N_21340,N_15813,N_15468);
and U21341 (N_21341,N_17276,N_15161);
and U21342 (N_21342,N_15956,N_17190);
nor U21343 (N_21343,N_13464,N_14921);
xor U21344 (N_21344,N_16021,N_14066);
nand U21345 (N_21345,N_17891,N_14967);
and U21346 (N_21346,N_13920,N_18075);
or U21347 (N_21347,N_18350,N_17382);
or U21348 (N_21348,N_18545,N_14023);
or U21349 (N_21349,N_13435,N_15284);
nand U21350 (N_21350,N_13810,N_18136);
nor U21351 (N_21351,N_14298,N_15283);
nor U21352 (N_21352,N_16146,N_13032);
and U21353 (N_21353,N_14179,N_14925);
nand U21354 (N_21354,N_12605,N_13170);
xnor U21355 (N_21355,N_14933,N_16833);
and U21356 (N_21356,N_14097,N_17555);
nor U21357 (N_21357,N_13237,N_16330);
nand U21358 (N_21358,N_15831,N_13141);
and U21359 (N_21359,N_13672,N_14439);
nand U21360 (N_21360,N_15201,N_13996);
nand U21361 (N_21361,N_18181,N_13929);
or U21362 (N_21362,N_14836,N_14495);
and U21363 (N_21363,N_18706,N_15883);
or U21364 (N_21364,N_17919,N_18366);
or U21365 (N_21365,N_18528,N_17146);
nand U21366 (N_21366,N_12921,N_17365);
nor U21367 (N_21367,N_18592,N_16883);
or U21368 (N_21368,N_13035,N_17284);
xor U21369 (N_21369,N_15198,N_13217);
nor U21370 (N_21370,N_17042,N_14716);
nand U21371 (N_21371,N_16404,N_14806);
or U21372 (N_21372,N_12724,N_14910);
or U21373 (N_21373,N_13447,N_16961);
nand U21374 (N_21374,N_18326,N_18422);
nor U21375 (N_21375,N_13075,N_18684);
nand U21376 (N_21376,N_14742,N_14898);
nor U21377 (N_21377,N_15940,N_13699);
nand U21378 (N_21378,N_15195,N_15997);
nor U21379 (N_21379,N_16206,N_13437);
and U21380 (N_21380,N_16271,N_15628);
and U21381 (N_21381,N_14059,N_16848);
or U21382 (N_21382,N_16517,N_16508);
nand U21383 (N_21383,N_17726,N_17825);
nor U21384 (N_21384,N_16910,N_15773);
nand U21385 (N_21385,N_12838,N_15041);
nor U21386 (N_21386,N_16874,N_16157);
and U21387 (N_21387,N_12525,N_13078);
nand U21388 (N_21388,N_17933,N_17800);
and U21389 (N_21389,N_18382,N_12776);
nor U21390 (N_21390,N_15644,N_14440);
or U21391 (N_21391,N_16167,N_17491);
and U21392 (N_21392,N_14473,N_18635);
xnor U21393 (N_21393,N_14318,N_14628);
nand U21394 (N_21394,N_12794,N_14068);
or U21395 (N_21395,N_13568,N_13980);
nand U21396 (N_21396,N_16394,N_17692);
or U21397 (N_21397,N_17319,N_16876);
or U21398 (N_21398,N_12852,N_16661);
xnor U21399 (N_21399,N_18216,N_13773);
nand U21400 (N_21400,N_13943,N_16279);
nand U21401 (N_21401,N_14285,N_12911);
and U21402 (N_21402,N_16672,N_15131);
xor U21403 (N_21403,N_18483,N_17829);
nor U21404 (N_21404,N_15953,N_16209);
nand U21405 (N_21405,N_15836,N_12547);
nand U21406 (N_21406,N_17454,N_16388);
or U21407 (N_21407,N_13858,N_14709);
or U21408 (N_21408,N_14536,N_18715);
xnor U21409 (N_21409,N_18613,N_16205);
or U21410 (N_21410,N_16711,N_17503);
and U21411 (N_21411,N_18263,N_14178);
and U21412 (N_21412,N_18153,N_17371);
or U21413 (N_21413,N_13902,N_14818);
and U21414 (N_21414,N_18549,N_17117);
and U21415 (N_21415,N_15104,N_15304);
nand U21416 (N_21416,N_15390,N_13880);
nand U21417 (N_21417,N_17859,N_16381);
or U21418 (N_21418,N_15580,N_16063);
nand U21419 (N_21419,N_14648,N_18306);
and U21420 (N_21420,N_13924,N_14128);
and U21421 (N_21421,N_18337,N_13364);
xor U21422 (N_21422,N_13222,N_15049);
nor U21423 (N_21423,N_12699,N_13572);
nor U21424 (N_21424,N_14968,N_15913);
or U21425 (N_21425,N_15693,N_13941);
and U21426 (N_21426,N_14020,N_18359);
or U21427 (N_21427,N_17481,N_18305);
and U21428 (N_21428,N_17745,N_14693);
or U21429 (N_21429,N_14277,N_18572);
or U21430 (N_21430,N_16421,N_14110);
nand U21431 (N_21431,N_16128,N_18679);
or U21432 (N_21432,N_14664,N_13143);
or U21433 (N_21433,N_17878,N_15563);
nand U21434 (N_21434,N_13008,N_16081);
and U21435 (N_21435,N_13820,N_13366);
and U21436 (N_21436,N_13710,N_15177);
nand U21437 (N_21437,N_13224,N_14751);
and U21438 (N_21438,N_17556,N_15032);
or U21439 (N_21439,N_17141,N_17666);
nand U21440 (N_21440,N_14884,N_13436);
nor U21441 (N_21441,N_18135,N_13837);
and U21442 (N_21442,N_18450,N_13014);
nand U21443 (N_21443,N_15315,N_18406);
nand U21444 (N_21444,N_16158,N_17938);
nor U21445 (N_21445,N_12766,N_14907);
or U21446 (N_21446,N_14738,N_13073);
and U21447 (N_21447,N_16727,N_16273);
or U21448 (N_21448,N_12542,N_14802);
or U21449 (N_21449,N_18415,N_15826);
nor U21450 (N_21450,N_13076,N_17789);
nand U21451 (N_21451,N_15064,N_14650);
and U21452 (N_21452,N_14198,N_18362);
nor U21453 (N_21453,N_17678,N_18193);
nand U21454 (N_21454,N_12926,N_17216);
nand U21455 (N_21455,N_17373,N_16079);
nor U21456 (N_21456,N_15012,N_12704);
xnor U21457 (N_21457,N_12872,N_13347);
and U21458 (N_21458,N_18081,N_17962);
nor U21459 (N_21459,N_16067,N_17065);
or U21460 (N_21460,N_13385,N_16229);
nand U21461 (N_21461,N_13269,N_16761);
xnor U21462 (N_21462,N_14281,N_16927);
nand U21463 (N_21463,N_17741,N_13225);
or U21464 (N_21464,N_16943,N_17598);
or U21465 (N_21465,N_13954,N_13947);
xor U21466 (N_21466,N_12786,N_13641);
nand U21467 (N_21467,N_16536,N_15230);
nand U21468 (N_21468,N_13201,N_13999);
xnor U21469 (N_21469,N_14382,N_12674);
and U21470 (N_21470,N_18647,N_17073);
or U21471 (N_21471,N_17652,N_17053);
nand U21472 (N_21472,N_15538,N_17405);
and U21473 (N_21473,N_13769,N_17852);
nor U21474 (N_21474,N_15379,N_14692);
nand U21475 (N_21475,N_12841,N_14957);
and U21476 (N_21476,N_15782,N_14119);
or U21477 (N_21477,N_15320,N_14640);
and U21478 (N_21478,N_13718,N_16581);
nor U21479 (N_21479,N_16786,N_14795);
and U21480 (N_21480,N_16481,N_16458);
nor U21481 (N_21481,N_16636,N_14082);
xor U21482 (N_21482,N_18456,N_15253);
and U21483 (N_21483,N_15014,N_15649);
or U21484 (N_21484,N_17123,N_14053);
nor U21485 (N_21485,N_18017,N_16578);
nor U21486 (N_21486,N_14514,N_15981);
nand U21487 (N_21487,N_17089,N_18351);
or U21488 (N_21488,N_14424,N_17522);
nor U21489 (N_21489,N_14267,N_16801);
or U21490 (N_21490,N_12732,N_13847);
and U21491 (N_21491,N_14325,N_16305);
nor U21492 (N_21492,N_14936,N_17961);
nand U21493 (N_21493,N_13895,N_13524);
xor U21494 (N_21494,N_15387,N_15465);
nand U21495 (N_21495,N_15039,N_14840);
or U21496 (N_21496,N_15237,N_14809);
nand U21497 (N_21497,N_18286,N_18127);
and U21498 (N_21498,N_13779,N_15768);
xor U21499 (N_21499,N_18269,N_17047);
or U21500 (N_21500,N_14798,N_18469);
nand U21501 (N_21501,N_13789,N_17664);
and U21502 (N_21502,N_13177,N_13212);
and U21503 (N_21503,N_17194,N_14859);
or U21504 (N_21504,N_12828,N_17103);
nand U21505 (N_21505,N_14422,N_13372);
and U21506 (N_21506,N_16654,N_16732);
and U21507 (N_21507,N_17372,N_15636);
and U21508 (N_21508,N_15335,N_15058);
or U21509 (N_21509,N_18441,N_16392);
nor U21510 (N_21510,N_16478,N_17226);
nor U21511 (N_21511,N_17854,N_15496);
or U21512 (N_21512,N_15023,N_14388);
nor U21513 (N_21513,N_16783,N_17806);
nand U21514 (N_21514,N_16162,N_12687);
nor U21515 (N_21515,N_18357,N_17041);
nor U21516 (N_21516,N_17286,N_16506);
or U21517 (N_21517,N_15472,N_13017);
or U21518 (N_21518,N_17070,N_18108);
nand U21519 (N_21519,N_16194,N_15839);
nor U21520 (N_21520,N_14074,N_14351);
nor U21521 (N_21521,N_12715,N_16405);
or U21522 (N_21522,N_13765,N_14089);
nand U21523 (N_21523,N_13066,N_17003);
xnor U21524 (N_21524,N_18063,N_15692);
nor U21525 (N_21525,N_15015,N_14356);
nor U21526 (N_21526,N_13260,N_14323);
and U21527 (N_21527,N_13238,N_16729);
xor U21528 (N_21528,N_13594,N_16213);
xor U21529 (N_21529,N_12749,N_14741);
nand U21530 (N_21530,N_14222,N_17772);
nand U21531 (N_21531,N_18058,N_14443);
and U21532 (N_21532,N_13536,N_16718);
nand U21533 (N_21533,N_17558,N_16201);
nor U21534 (N_21534,N_14093,N_17597);
nand U21535 (N_21535,N_18733,N_14557);
or U21536 (N_21536,N_13665,N_16358);
and U21537 (N_21537,N_15600,N_13879);
and U21538 (N_21538,N_12693,N_13736);
or U21539 (N_21539,N_18138,N_14187);
nor U21540 (N_21540,N_14048,N_17681);
nor U21541 (N_21541,N_15061,N_13983);
nor U21542 (N_21542,N_14929,N_17414);
nor U21543 (N_21543,N_16666,N_15690);
and U21544 (N_21544,N_13219,N_14561);
and U21545 (N_21545,N_17375,N_12824);
nor U21546 (N_21546,N_16865,N_16817);
xor U21547 (N_21547,N_15560,N_16823);
nor U21548 (N_21548,N_15565,N_17993);
or U21549 (N_21549,N_16116,N_14397);
nor U21550 (N_21550,N_15504,N_17894);
nand U21551 (N_21551,N_15985,N_13358);
and U21552 (N_21552,N_12641,N_14996);
and U21553 (N_21553,N_17449,N_13130);
nand U21554 (N_21554,N_13790,N_15028);
and U21555 (N_21555,N_13585,N_16662);
or U21556 (N_21556,N_12886,N_15119);
nand U21557 (N_21557,N_16147,N_17495);
nand U21558 (N_21558,N_15261,N_16856);
or U21559 (N_21559,N_15890,N_15172);
xnor U21560 (N_21560,N_17045,N_14007);
nor U21561 (N_21561,N_13207,N_16600);
nand U21562 (N_21562,N_12551,N_17099);
nor U21563 (N_21563,N_14548,N_12789);
or U21564 (N_21564,N_15967,N_17706);
nor U21565 (N_21565,N_13978,N_13818);
and U21566 (N_21566,N_13904,N_16342);
or U21567 (N_21567,N_16934,N_13951);
and U21568 (N_21568,N_17000,N_15044);
and U21569 (N_21569,N_17461,N_13791);
nand U21570 (N_21570,N_13643,N_14901);
xor U21571 (N_21571,N_14006,N_14710);
nor U21572 (N_21572,N_15477,N_16681);
nor U21573 (N_21573,N_12642,N_15007);
nand U21574 (N_21574,N_15545,N_16297);
nand U21575 (N_21575,N_14350,N_17721);
nand U21576 (N_21576,N_12980,N_17324);
nor U21577 (N_21577,N_13921,N_17096);
and U21578 (N_21578,N_17968,N_17122);
nand U21579 (N_21579,N_14701,N_18367);
xor U21580 (N_21580,N_13694,N_13223);
and U21581 (N_21581,N_13558,N_14312);
and U21582 (N_21582,N_14042,N_16791);
xor U21583 (N_21583,N_17085,N_16444);
and U21584 (N_21584,N_15442,N_16234);
or U21585 (N_21585,N_12570,N_17455);
nand U21586 (N_21586,N_17113,N_13682);
nor U21587 (N_21587,N_18457,N_15599);
or U21588 (N_21588,N_16112,N_17158);
and U21589 (N_21589,N_13959,N_15637);
and U21590 (N_21590,N_17758,N_14630);
nand U21591 (N_21591,N_13476,N_16174);
or U21592 (N_21592,N_13784,N_16687);
nand U21593 (N_21593,N_15715,N_13750);
nand U21594 (N_21594,N_17381,N_17055);
nand U21595 (N_21595,N_14560,N_15734);
or U21596 (N_21596,N_15460,N_13382);
nor U21597 (N_21597,N_13312,N_14253);
or U21598 (N_21598,N_16808,N_14913);
or U21599 (N_21599,N_13652,N_12800);
nand U21600 (N_21600,N_17114,N_18554);
nor U21601 (N_21601,N_12862,N_12836);
xnor U21602 (N_21602,N_16089,N_15595);
and U21603 (N_21603,N_14869,N_12773);
xor U21604 (N_21604,N_14671,N_17936);
nor U21605 (N_21605,N_18276,N_13202);
nor U21606 (N_21606,N_15617,N_17812);
nand U21607 (N_21607,N_15199,N_17871);
xnor U21608 (N_21608,N_16431,N_13124);
and U21609 (N_21609,N_15561,N_17831);
and U21610 (N_21610,N_13216,N_16427);
nor U21611 (N_21611,N_13917,N_12658);
nor U21612 (N_21612,N_14945,N_17685);
or U21613 (N_21613,N_17551,N_13618);
and U21614 (N_21614,N_18663,N_16126);
nand U21615 (N_21615,N_16526,N_14755);
nand U21616 (N_21616,N_13722,N_16035);
nor U21617 (N_21617,N_12771,N_16709);
nor U21618 (N_21618,N_18376,N_16418);
nand U21619 (N_21619,N_17673,N_14261);
xor U21620 (N_21620,N_13208,N_18234);
nand U21621 (N_21621,N_13679,N_16884);
nor U21622 (N_21622,N_12909,N_18104);
or U21623 (N_21623,N_17069,N_16055);
nor U21624 (N_21624,N_13584,N_15499);
nand U21625 (N_21625,N_18586,N_13800);
nor U21626 (N_21626,N_13690,N_15569);
or U21627 (N_21627,N_18688,N_13413);
xnor U21628 (N_21628,N_14998,N_18508);
nor U21629 (N_21629,N_14899,N_16968);
nand U21630 (N_21630,N_13140,N_17587);
nand U21631 (N_21631,N_17248,N_14359);
nor U21632 (N_21632,N_18261,N_18708);
nand U21633 (N_21633,N_14039,N_16261);
or U21634 (N_21634,N_14366,N_17959);
nor U21635 (N_21635,N_16935,N_13119);
or U21636 (N_21636,N_14790,N_15445);
nand U21637 (N_21637,N_18588,N_14213);
or U21638 (N_21638,N_18055,N_14405);
and U21639 (N_21639,N_18600,N_13792);
nand U21640 (N_21640,N_14064,N_15146);
nand U21641 (N_21641,N_18325,N_15115);
and U21642 (N_21642,N_13261,N_13727);
or U21643 (N_21643,N_16756,N_17957);
nor U21644 (N_21644,N_17456,N_16759);
and U21645 (N_21645,N_15869,N_18629);
nand U21646 (N_21646,N_13998,N_18345);
nand U21647 (N_21647,N_12745,N_16129);
and U21648 (N_21648,N_13650,N_16275);
and U21649 (N_21649,N_17334,N_17187);
nor U21650 (N_21650,N_18160,N_14897);
nor U21651 (N_21651,N_15287,N_18340);
nand U21652 (N_21652,N_18608,N_16240);
nand U21653 (N_21653,N_15719,N_14521);
nor U21654 (N_21654,N_17729,N_17230);
nor U21655 (N_21655,N_17505,N_16866);
and U21656 (N_21656,N_15588,N_17298);
or U21657 (N_21657,N_18051,N_16787);
and U21658 (N_21658,N_12746,N_17435);
xor U21659 (N_21659,N_13128,N_15453);
or U21660 (N_21660,N_15818,N_18238);
nor U21661 (N_21661,N_14441,N_13602);
and U21662 (N_21662,N_12816,N_18669);
and U21663 (N_21663,N_15392,N_13133);
and U21664 (N_21664,N_16929,N_13976);
or U21665 (N_21665,N_13409,N_16970);
nor U21666 (N_21666,N_18298,N_16017);
nor U21667 (N_21667,N_12991,N_12743);
nand U21668 (N_21668,N_14552,N_13349);
and U21669 (N_21669,N_16638,N_13040);
nor U21670 (N_21670,N_15129,N_18169);
and U21671 (N_21671,N_17895,N_15005);
nor U21672 (N_21672,N_18526,N_18398);
and U21673 (N_21673,N_16053,N_17535);
or U21674 (N_21674,N_18711,N_15645);
nor U21675 (N_21675,N_15065,N_17316);
and U21676 (N_21676,N_16451,N_18312);
nand U21677 (N_21677,N_17940,N_12663);
and U21678 (N_21678,N_16383,N_16400);
nand U21679 (N_21679,N_15964,N_14980);
nor U21680 (N_21680,N_16257,N_14758);
nand U21681 (N_21681,N_14335,N_18487);
xnor U21682 (N_21682,N_13046,N_15324);
nor U21683 (N_21683,N_12783,N_13085);
nand U21684 (N_21684,N_16609,N_16200);
and U21685 (N_21685,N_16579,N_17246);
or U21686 (N_21686,N_17875,N_15520);
and U21687 (N_21687,N_16892,N_16386);
or U21688 (N_21688,N_16898,N_12592);
or U21689 (N_21689,N_18033,N_13221);
nor U21690 (N_21690,N_16545,N_15337);
nor U21691 (N_21691,N_14393,N_12827);
nand U21692 (N_21692,N_13591,N_13948);
and U21693 (N_21693,N_13667,N_14748);
nand U21694 (N_21694,N_17759,N_14324);
and U21695 (N_21695,N_15688,N_17662);
and U21696 (N_21696,N_14164,N_14730);
nor U21697 (N_21697,N_18297,N_13542);
and U21698 (N_21698,N_13704,N_15577);
nor U21699 (N_21699,N_12643,N_17474);
or U21700 (N_21700,N_17213,N_18656);
nor U21701 (N_21701,N_18544,N_13023);
nand U21702 (N_21702,N_14624,N_14895);
and U21703 (N_21703,N_13074,N_17184);
or U21704 (N_21704,N_18176,N_16019);
nand U21705 (N_21705,N_13936,N_17422);
nand U21706 (N_21706,N_15822,N_15389);
and U21707 (N_21707,N_15880,N_18004);
or U21708 (N_21708,N_16183,N_13438);
or U21709 (N_21709,N_18399,N_14129);
nand U21710 (N_21710,N_16975,N_18491);
nor U21711 (N_21711,N_14567,N_12665);
and U21712 (N_21712,N_17004,N_18522);
and U21713 (N_21713,N_15935,N_14904);
and U21714 (N_21714,N_14199,N_16424);
nor U21715 (N_21715,N_12532,N_14662);
and U21716 (N_21716,N_13551,N_18034);
nor U21717 (N_21717,N_13022,N_16288);
or U21718 (N_21718,N_17364,N_17820);
and U21719 (N_21719,N_13293,N_17557);
nor U21720 (N_21720,N_13446,N_17740);
nand U21721 (N_21721,N_14360,N_15406);
nor U21722 (N_21722,N_14151,N_14787);
and U21723 (N_21723,N_15680,N_13461);
and U21724 (N_21724,N_12835,N_15629);
nor U21725 (N_21725,N_14655,N_13937);
xnor U21726 (N_21726,N_12707,N_14387);
and U21727 (N_21727,N_13326,N_13111);
nor U21728 (N_21728,N_12535,N_14931);
nor U21729 (N_21729,N_14545,N_17653);
or U21730 (N_21730,N_15731,N_17185);
nand U21731 (N_21731,N_14508,N_15016);
nand U21732 (N_21732,N_16061,N_17999);
nand U21733 (N_21733,N_17412,N_16176);
and U21734 (N_21734,N_18626,N_17348);
and U21735 (N_21735,N_16765,N_18620);
nand U21736 (N_21736,N_17105,N_18423);
nand U21737 (N_21737,N_16339,N_16552);
xnor U21738 (N_21738,N_17329,N_13755);
xor U21739 (N_21739,N_17648,N_15303);
nor U21740 (N_21740,N_16944,N_18448);
or U21741 (N_21741,N_18327,N_15280);
xnor U21742 (N_21742,N_14413,N_17465);
nor U21743 (N_21743,N_15950,N_15259);
and U21744 (N_21744,N_15145,N_12717);
and U21745 (N_21745,N_13354,N_17243);
nand U21746 (N_21746,N_13004,N_18400);
nor U21747 (N_21747,N_17445,N_14615);
nand U21748 (N_21748,N_12907,N_17290);
and U21749 (N_21749,N_18348,N_17007);
or U21750 (N_21750,N_17249,N_16857);
nand U21751 (N_21751,N_17228,N_17462);
or U21752 (N_21752,N_12709,N_12956);
nand U21753 (N_21753,N_18470,N_17341);
and U21754 (N_21754,N_15982,N_13175);
nor U21755 (N_21755,N_14276,N_14450);
and U21756 (N_21756,N_14174,N_15213);
and U21757 (N_21757,N_12562,N_18494);
or U21758 (N_21758,N_14577,N_12669);
or U21759 (N_21759,N_12518,N_14918);
or U21760 (N_21760,N_17177,N_16181);
nor U21761 (N_21761,N_13887,N_13069);
or U21762 (N_21762,N_18581,N_16144);
nor U21763 (N_21763,N_17575,N_16914);
or U21764 (N_21764,N_12565,N_17814);
nor U21765 (N_21765,N_13723,N_15827);
nor U21766 (N_21766,N_17784,N_18461);
and U21767 (N_21767,N_16185,N_17682);
nor U21768 (N_21768,N_18430,N_18324);
and U21769 (N_21769,N_15566,N_17994);
and U21770 (N_21770,N_13564,N_14973);
nand U21771 (N_21771,N_13759,N_17880);
and U21772 (N_21772,N_12894,N_14578);
nand U21773 (N_21773,N_17701,N_15142);
nand U21774 (N_21774,N_15998,N_15972);
and U21775 (N_21775,N_16266,N_16538);
or U21776 (N_21776,N_18118,N_17580);
nor U21777 (N_21777,N_17651,N_15431);
nor U21778 (N_21778,N_15907,N_15619);
nand U21779 (N_21779,N_13434,N_13229);
and U21780 (N_21780,N_15683,N_18466);
nor U21781 (N_21781,N_17517,N_16713);
and U21782 (N_21782,N_17388,N_17144);
nor U21783 (N_21783,N_18642,N_16286);
nand U21784 (N_21784,N_13754,N_14769);
nand U21785 (N_21785,N_14903,N_16000);
nand U21786 (N_21786,N_16224,N_13356);
or U21787 (N_21787,N_15774,N_13402);
nor U21788 (N_21788,N_17305,N_13984);
nand U21789 (N_21789,N_17165,N_12905);
nor U21790 (N_21790,N_12539,N_18486);
nand U21791 (N_21791,N_13559,N_13720);
and U21792 (N_21792,N_14695,N_17490);
nor U21793 (N_21793,N_14530,N_17984);
or U21794 (N_21794,N_14262,N_16700);
nor U21795 (N_21795,N_18716,N_14113);
nand U21796 (N_21796,N_13509,N_14184);
and U21797 (N_21797,N_16746,N_14803);
nand U21798 (N_21798,N_18649,N_17764);
and U21799 (N_21799,N_18180,N_13993);
or U21800 (N_21800,N_15382,N_17520);
or U21801 (N_21801,N_14340,N_15120);
nand U21802 (N_21802,N_16496,N_16228);
nand U21803 (N_21803,N_16591,N_17714);
nor U21804 (N_21804,N_12588,N_17057);
nand U21805 (N_21805,N_18149,N_14333);
nor U21806 (N_21806,N_16247,N_18736);
and U21807 (N_21807,N_17119,N_18256);
nand U21808 (N_21808,N_13061,N_17061);
nand U21809 (N_21809,N_16422,N_14438);
or U21810 (N_21810,N_16543,N_13724);
and U21811 (N_21811,N_18346,N_14431);
xor U21812 (N_21812,N_18569,N_17272);
nand U21813 (N_21813,N_17856,N_17325);
nor U21814 (N_21814,N_13189,N_13359);
or U21815 (N_21815,N_12610,N_16231);
nor U21816 (N_21816,N_14919,N_18106);
and U21817 (N_21817,N_15885,N_12772);
or U21818 (N_21818,N_14377,N_13977);
or U21819 (N_21819,N_13093,N_15299);
nand U21820 (N_21820,N_16565,N_17001);
and U21821 (N_21821,N_17360,N_14908);
nor U21822 (N_21822,N_13934,N_16684);
or U21823 (N_21823,N_15681,N_16515);
nand U21824 (N_21824,N_18283,N_13210);
nor U21825 (N_21825,N_13485,N_17679);
and U21826 (N_21826,N_15351,N_14947);
or U21827 (N_21827,N_16510,N_16045);
and U21828 (N_21828,N_15928,N_17183);
nand U21829 (N_21829,N_14983,N_14328);
nand U21830 (N_21830,N_14299,N_17335);
nand U21831 (N_21831,N_13811,N_16511);
nor U21832 (N_21832,N_16050,N_12748);
xor U21833 (N_21833,N_13538,N_18280);
nand U21834 (N_21834,N_16367,N_17407);
xnor U21835 (N_21835,N_14263,N_14700);
or U21836 (N_21836,N_13688,N_14292);
or U21837 (N_21837,N_16908,N_16346);
nor U21838 (N_21838,N_15495,N_15264);
or U21839 (N_21839,N_14036,N_17621);
nand U21840 (N_21840,N_14735,N_13782);
nor U21841 (N_21841,N_14623,N_14712);
or U21842 (N_21842,N_13930,N_15850);
and U21843 (N_21843,N_16477,N_17835);
nor U21844 (N_21844,N_15936,N_15278);
nand U21845 (N_21845,N_12958,N_15258);
or U21846 (N_21846,N_14342,N_13138);
nand U21847 (N_21847,N_12826,N_16974);
nor U21848 (N_21848,N_18078,N_13401);
nor U21849 (N_21849,N_18178,N_17686);
or U21850 (N_21850,N_14305,N_18705);
nor U21851 (N_21851,N_18045,N_18349);
nand U21852 (N_21852,N_17656,N_15480);
or U21853 (N_21853,N_16762,N_14777);
and U21854 (N_21854,N_15367,N_16198);
xor U21855 (N_21855,N_18418,N_12941);
or U21856 (N_21856,N_15211,N_13475);
and U21857 (N_21857,N_13698,N_17512);
nor U21858 (N_21858,N_13668,N_12857);
xnor U21859 (N_21859,N_14412,N_14668);
nand U21860 (N_21860,N_16905,N_14025);
nor U21861 (N_21861,N_17927,N_12580);
and U21862 (N_21862,N_12514,N_16487);
xnor U21863 (N_21863,N_17496,N_15663);
nand U21864 (N_21864,N_14109,N_14871);
or U21865 (N_21865,N_14985,N_14882);
nand U21866 (N_21866,N_18272,N_18651);
and U21867 (N_21867,N_17916,N_13243);
or U21868 (N_21868,N_16042,N_16317);
or U21869 (N_21869,N_15245,N_14067);
and U21870 (N_21870,N_12829,N_14631);
nor U21871 (N_21871,N_13197,N_14826);
nand U21872 (N_21872,N_15464,N_13940);
or U21873 (N_21873,N_17592,N_12626);
and U21874 (N_21874,N_17486,N_18594);
nor U21875 (N_21875,N_16764,N_13635);
xor U21876 (N_21876,N_18121,N_18074);
nand U21877 (N_21877,N_15463,N_17624);
nor U21878 (N_21878,N_18243,N_17504);
and U21879 (N_21879,N_15078,N_16496);
nor U21880 (N_21880,N_18674,N_16290);
and U21881 (N_21881,N_13156,N_16776);
nand U21882 (N_21882,N_12730,N_17215);
or U21883 (N_21883,N_13110,N_15837);
xor U21884 (N_21884,N_17129,N_14494);
xor U21885 (N_21885,N_15164,N_17421);
and U21886 (N_21886,N_16356,N_15019);
xnor U21887 (N_21887,N_17891,N_12621);
nand U21888 (N_21888,N_15756,N_15589);
or U21889 (N_21889,N_18432,N_15291);
nand U21890 (N_21890,N_18545,N_14751);
nor U21891 (N_21891,N_14874,N_16694);
xor U21892 (N_21892,N_14087,N_13994);
or U21893 (N_21893,N_16213,N_13710);
nor U21894 (N_21894,N_18333,N_16623);
nand U21895 (N_21895,N_17892,N_16736);
nor U21896 (N_21896,N_18436,N_14506);
nor U21897 (N_21897,N_17888,N_14087);
or U21898 (N_21898,N_16003,N_13349);
and U21899 (N_21899,N_17089,N_13682);
and U21900 (N_21900,N_15898,N_13825);
nor U21901 (N_21901,N_13404,N_16802);
nor U21902 (N_21902,N_16596,N_13886);
nor U21903 (N_21903,N_13078,N_16033);
and U21904 (N_21904,N_16847,N_17788);
and U21905 (N_21905,N_13848,N_15829);
nand U21906 (N_21906,N_16667,N_14344);
or U21907 (N_21907,N_17893,N_16123);
xnor U21908 (N_21908,N_15338,N_15977);
or U21909 (N_21909,N_16120,N_18521);
nand U21910 (N_21910,N_18130,N_17222);
and U21911 (N_21911,N_15684,N_14006);
nor U21912 (N_21912,N_12578,N_15365);
or U21913 (N_21913,N_14097,N_14449);
nand U21914 (N_21914,N_16223,N_13907);
nand U21915 (N_21915,N_18355,N_16066);
and U21916 (N_21916,N_17347,N_17269);
nand U21917 (N_21917,N_15505,N_18491);
xnor U21918 (N_21918,N_15892,N_18635);
nor U21919 (N_21919,N_16498,N_15210);
or U21920 (N_21920,N_14948,N_17621);
and U21921 (N_21921,N_16219,N_17719);
nor U21922 (N_21922,N_17635,N_16756);
nor U21923 (N_21923,N_13924,N_15869);
nor U21924 (N_21924,N_18186,N_13504);
nand U21925 (N_21925,N_16490,N_13812);
nand U21926 (N_21926,N_14419,N_14047);
nand U21927 (N_21927,N_13448,N_13096);
nor U21928 (N_21928,N_13345,N_13897);
nand U21929 (N_21929,N_18529,N_13676);
nor U21930 (N_21930,N_12865,N_15220);
and U21931 (N_21931,N_12809,N_13730);
nor U21932 (N_21932,N_16783,N_13146);
or U21933 (N_21933,N_13131,N_14790);
xor U21934 (N_21934,N_15814,N_18478);
nor U21935 (N_21935,N_15189,N_17359);
and U21936 (N_21936,N_15454,N_13103);
or U21937 (N_21937,N_16305,N_16672);
or U21938 (N_21938,N_14644,N_17984);
nand U21939 (N_21939,N_14554,N_16474);
nand U21940 (N_21940,N_17952,N_13477);
nor U21941 (N_21941,N_13718,N_16635);
or U21942 (N_21942,N_14302,N_12655);
nand U21943 (N_21943,N_14185,N_12945);
nor U21944 (N_21944,N_14733,N_17430);
nor U21945 (N_21945,N_16647,N_12748);
and U21946 (N_21946,N_17262,N_17506);
xnor U21947 (N_21947,N_15756,N_18124);
or U21948 (N_21948,N_13456,N_16633);
or U21949 (N_21949,N_16905,N_13206);
and U21950 (N_21950,N_16437,N_17731);
nand U21951 (N_21951,N_15753,N_16148);
nand U21952 (N_21952,N_17918,N_15071);
and U21953 (N_21953,N_18090,N_17432);
and U21954 (N_21954,N_17932,N_12872);
xor U21955 (N_21955,N_13711,N_17296);
nor U21956 (N_21956,N_16847,N_13033);
or U21957 (N_21957,N_17612,N_18650);
or U21958 (N_21958,N_14020,N_13086);
and U21959 (N_21959,N_17702,N_14053);
or U21960 (N_21960,N_16050,N_18393);
nand U21961 (N_21961,N_15333,N_14462);
nand U21962 (N_21962,N_12642,N_17615);
xor U21963 (N_21963,N_17792,N_17432);
and U21964 (N_21964,N_15744,N_15987);
nor U21965 (N_21965,N_14306,N_18330);
nand U21966 (N_21966,N_17712,N_17752);
or U21967 (N_21967,N_15857,N_17919);
and U21968 (N_21968,N_16772,N_14002);
and U21969 (N_21969,N_14200,N_13779);
and U21970 (N_21970,N_18309,N_18485);
or U21971 (N_21971,N_17216,N_14326);
and U21972 (N_21972,N_14506,N_16322);
xnor U21973 (N_21973,N_15195,N_17847);
and U21974 (N_21974,N_15905,N_13927);
and U21975 (N_21975,N_15415,N_15108);
and U21976 (N_21976,N_17227,N_18602);
or U21977 (N_21977,N_17541,N_14777);
xor U21978 (N_21978,N_13455,N_18260);
or U21979 (N_21979,N_17265,N_17638);
nand U21980 (N_21980,N_16607,N_16405);
xor U21981 (N_21981,N_15917,N_14132);
nand U21982 (N_21982,N_18532,N_13763);
or U21983 (N_21983,N_12558,N_18694);
or U21984 (N_21984,N_12853,N_17056);
nor U21985 (N_21985,N_14273,N_17008);
nand U21986 (N_21986,N_17696,N_16939);
or U21987 (N_21987,N_17216,N_15193);
and U21988 (N_21988,N_15902,N_13146);
nand U21989 (N_21989,N_17798,N_13554);
nor U21990 (N_21990,N_15735,N_17811);
xnor U21991 (N_21991,N_16577,N_16363);
xnor U21992 (N_21992,N_17216,N_17755);
and U21993 (N_21993,N_16842,N_13916);
or U21994 (N_21994,N_14820,N_16723);
nor U21995 (N_21995,N_17338,N_16908);
nand U21996 (N_21996,N_18669,N_16095);
nand U21997 (N_21997,N_17402,N_15664);
or U21998 (N_21998,N_16650,N_12708);
nor U21999 (N_21999,N_14775,N_14810);
nor U22000 (N_22000,N_13668,N_18090);
nor U22001 (N_22001,N_17545,N_15151);
nand U22002 (N_22002,N_18508,N_17612);
or U22003 (N_22003,N_14542,N_15341);
or U22004 (N_22004,N_18313,N_17838);
or U22005 (N_22005,N_13103,N_16200);
xnor U22006 (N_22006,N_18314,N_12596);
and U22007 (N_22007,N_12580,N_14184);
and U22008 (N_22008,N_13617,N_16642);
nand U22009 (N_22009,N_13963,N_13559);
or U22010 (N_22010,N_13788,N_14564);
or U22011 (N_22011,N_14000,N_18464);
nor U22012 (N_22012,N_17669,N_15662);
nand U22013 (N_22013,N_18239,N_15806);
nor U22014 (N_22014,N_18672,N_16827);
xor U22015 (N_22015,N_15692,N_12617);
and U22016 (N_22016,N_16279,N_17001);
and U22017 (N_22017,N_14411,N_17854);
or U22018 (N_22018,N_15781,N_17197);
nor U22019 (N_22019,N_14827,N_17662);
nand U22020 (N_22020,N_14159,N_13398);
or U22021 (N_22021,N_14686,N_15166);
nand U22022 (N_22022,N_16888,N_15264);
and U22023 (N_22023,N_17182,N_14120);
and U22024 (N_22024,N_13586,N_14379);
or U22025 (N_22025,N_14539,N_13961);
or U22026 (N_22026,N_16793,N_14013);
or U22027 (N_22027,N_13527,N_17728);
and U22028 (N_22028,N_13476,N_13650);
nand U22029 (N_22029,N_17853,N_17456);
nor U22030 (N_22030,N_16765,N_16501);
nand U22031 (N_22031,N_14927,N_15047);
nor U22032 (N_22032,N_14884,N_12855);
and U22033 (N_22033,N_14922,N_17113);
nor U22034 (N_22034,N_14765,N_17059);
nor U22035 (N_22035,N_14040,N_12882);
or U22036 (N_22036,N_16170,N_12820);
or U22037 (N_22037,N_16097,N_15986);
and U22038 (N_22038,N_16117,N_17880);
nor U22039 (N_22039,N_17056,N_13203);
nor U22040 (N_22040,N_18728,N_14042);
and U22041 (N_22041,N_17432,N_16414);
and U22042 (N_22042,N_16669,N_14291);
and U22043 (N_22043,N_12650,N_17223);
nand U22044 (N_22044,N_14126,N_12687);
and U22045 (N_22045,N_15135,N_18242);
and U22046 (N_22046,N_12578,N_18122);
nor U22047 (N_22047,N_18340,N_16888);
and U22048 (N_22048,N_14787,N_16066);
nand U22049 (N_22049,N_18281,N_17246);
or U22050 (N_22050,N_17706,N_17960);
nand U22051 (N_22051,N_18492,N_14415);
or U22052 (N_22052,N_13140,N_17911);
or U22053 (N_22053,N_13644,N_13923);
nor U22054 (N_22054,N_16116,N_18460);
and U22055 (N_22055,N_13310,N_16865);
nor U22056 (N_22056,N_17303,N_16813);
nand U22057 (N_22057,N_14443,N_13270);
or U22058 (N_22058,N_16721,N_13683);
nor U22059 (N_22059,N_15055,N_17870);
or U22060 (N_22060,N_12760,N_16151);
nand U22061 (N_22061,N_14214,N_15074);
xnor U22062 (N_22062,N_17775,N_16621);
nand U22063 (N_22063,N_14156,N_13222);
and U22064 (N_22064,N_13458,N_18744);
nand U22065 (N_22065,N_16556,N_12555);
or U22066 (N_22066,N_15858,N_14078);
or U22067 (N_22067,N_18264,N_18360);
and U22068 (N_22068,N_13780,N_14101);
and U22069 (N_22069,N_15469,N_13124);
and U22070 (N_22070,N_14121,N_18476);
nor U22071 (N_22071,N_16878,N_14213);
or U22072 (N_22072,N_13956,N_13951);
or U22073 (N_22073,N_18583,N_17058);
or U22074 (N_22074,N_13190,N_15826);
or U22075 (N_22075,N_17027,N_13666);
nand U22076 (N_22076,N_14132,N_14420);
nor U22077 (N_22077,N_15640,N_13857);
and U22078 (N_22078,N_14991,N_17159);
nor U22079 (N_22079,N_14514,N_16909);
nor U22080 (N_22080,N_14439,N_17490);
or U22081 (N_22081,N_14425,N_13302);
or U22082 (N_22082,N_16397,N_16466);
nor U22083 (N_22083,N_12598,N_15148);
nor U22084 (N_22084,N_15619,N_17960);
nand U22085 (N_22085,N_15009,N_14643);
or U22086 (N_22086,N_15179,N_13731);
and U22087 (N_22087,N_14967,N_16657);
or U22088 (N_22088,N_15998,N_12942);
nor U22089 (N_22089,N_14602,N_15952);
or U22090 (N_22090,N_12586,N_13551);
or U22091 (N_22091,N_14662,N_14325);
or U22092 (N_22092,N_17472,N_15652);
and U22093 (N_22093,N_15502,N_12945);
nor U22094 (N_22094,N_12917,N_18412);
xnor U22095 (N_22095,N_17456,N_15438);
and U22096 (N_22096,N_13185,N_15489);
nand U22097 (N_22097,N_17194,N_16297);
nor U22098 (N_22098,N_16466,N_18550);
nand U22099 (N_22099,N_18685,N_14197);
or U22100 (N_22100,N_15924,N_17148);
nand U22101 (N_22101,N_13677,N_16074);
or U22102 (N_22102,N_12785,N_16588);
or U22103 (N_22103,N_18619,N_14945);
and U22104 (N_22104,N_18717,N_15339);
or U22105 (N_22105,N_15543,N_13803);
nand U22106 (N_22106,N_16905,N_16314);
and U22107 (N_22107,N_18033,N_13421);
nand U22108 (N_22108,N_14310,N_18492);
or U22109 (N_22109,N_15628,N_15900);
nor U22110 (N_22110,N_17035,N_15155);
or U22111 (N_22111,N_18282,N_13336);
nor U22112 (N_22112,N_15849,N_16239);
or U22113 (N_22113,N_15237,N_16793);
or U22114 (N_22114,N_16043,N_17589);
nor U22115 (N_22115,N_13607,N_16793);
xnor U22116 (N_22116,N_15544,N_18477);
nor U22117 (N_22117,N_17307,N_14088);
nor U22118 (N_22118,N_12759,N_16680);
nand U22119 (N_22119,N_15911,N_17291);
and U22120 (N_22120,N_14622,N_15659);
xnor U22121 (N_22121,N_15870,N_17557);
nor U22122 (N_22122,N_12525,N_18576);
and U22123 (N_22123,N_13412,N_16983);
or U22124 (N_22124,N_16705,N_15271);
nand U22125 (N_22125,N_16587,N_13271);
xnor U22126 (N_22126,N_14601,N_18456);
nand U22127 (N_22127,N_14675,N_16360);
or U22128 (N_22128,N_16276,N_13363);
nor U22129 (N_22129,N_15939,N_18463);
and U22130 (N_22130,N_16649,N_16937);
xnor U22131 (N_22131,N_13369,N_18008);
xor U22132 (N_22132,N_13036,N_18411);
or U22133 (N_22133,N_16877,N_12657);
nor U22134 (N_22134,N_15441,N_18530);
and U22135 (N_22135,N_18410,N_16572);
nor U22136 (N_22136,N_16694,N_13258);
nor U22137 (N_22137,N_18347,N_14845);
xnor U22138 (N_22138,N_13518,N_15176);
or U22139 (N_22139,N_13778,N_17865);
and U22140 (N_22140,N_18313,N_13787);
and U22141 (N_22141,N_14363,N_13868);
nand U22142 (N_22142,N_14098,N_16201);
nor U22143 (N_22143,N_15548,N_15951);
or U22144 (N_22144,N_14390,N_14856);
xor U22145 (N_22145,N_18404,N_16511);
and U22146 (N_22146,N_12677,N_16650);
nand U22147 (N_22147,N_14341,N_16086);
or U22148 (N_22148,N_17203,N_13609);
xnor U22149 (N_22149,N_15752,N_13555);
nor U22150 (N_22150,N_18413,N_14534);
nand U22151 (N_22151,N_16061,N_17649);
nand U22152 (N_22152,N_14048,N_12734);
xor U22153 (N_22153,N_17244,N_14899);
nor U22154 (N_22154,N_15288,N_17728);
or U22155 (N_22155,N_12813,N_14387);
nand U22156 (N_22156,N_14209,N_17943);
nor U22157 (N_22157,N_17443,N_17189);
xor U22158 (N_22158,N_18426,N_13345);
nand U22159 (N_22159,N_16165,N_13730);
nor U22160 (N_22160,N_16658,N_16233);
or U22161 (N_22161,N_18325,N_13196);
and U22162 (N_22162,N_14187,N_16798);
or U22163 (N_22163,N_14322,N_16312);
and U22164 (N_22164,N_15816,N_17211);
or U22165 (N_22165,N_18026,N_13863);
or U22166 (N_22166,N_13556,N_13784);
nor U22167 (N_22167,N_14711,N_12678);
and U22168 (N_22168,N_18061,N_13518);
or U22169 (N_22169,N_15313,N_12854);
xor U22170 (N_22170,N_16395,N_16834);
or U22171 (N_22171,N_17046,N_13589);
and U22172 (N_22172,N_13454,N_18437);
or U22173 (N_22173,N_14090,N_16577);
and U22174 (N_22174,N_14108,N_16996);
nor U22175 (N_22175,N_13386,N_14332);
nand U22176 (N_22176,N_16844,N_16058);
nor U22177 (N_22177,N_16087,N_14160);
or U22178 (N_22178,N_14291,N_18585);
and U22179 (N_22179,N_17436,N_14563);
nor U22180 (N_22180,N_17453,N_15845);
and U22181 (N_22181,N_17393,N_12947);
nor U22182 (N_22182,N_18635,N_14163);
nor U22183 (N_22183,N_13154,N_17499);
xor U22184 (N_22184,N_17566,N_18218);
nand U22185 (N_22185,N_13191,N_15847);
and U22186 (N_22186,N_14029,N_15197);
nand U22187 (N_22187,N_13629,N_17846);
nor U22188 (N_22188,N_15244,N_17093);
nand U22189 (N_22189,N_17983,N_13331);
nand U22190 (N_22190,N_13087,N_18028);
or U22191 (N_22191,N_12686,N_17376);
nand U22192 (N_22192,N_12823,N_14982);
nor U22193 (N_22193,N_14895,N_16674);
nand U22194 (N_22194,N_13214,N_16248);
or U22195 (N_22195,N_14201,N_17658);
and U22196 (N_22196,N_13711,N_13054);
nand U22197 (N_22197,N_17298,N_18659);
and U22198 (N_22198,N_13952,N_12555);
and U22199 (N_22199,N_13885,N_13468);
nand U22200 (N_22200,N_16373,N_17085);
nor U22201 (N_22201,N_17808,N_14984);
or U22202 (N_22202,N_13331,N_12573);
or U22203 (N_22203,N_18221,N_14633);
nor U22204 (N_22204,N_16330,N_17328);
or U22205 (N_22205,N_12533,N_17485);
nand U22206 (N_22206,N_16542,N_15472);
nor U22207 (N_22207,N_16378,N_18466);
and U22208 (N_22208,N_13491,N_13035);
nor U22209 (N_22209,N_16670,N_13622);
and U22210 (N_22210,N_13842,N_14168);
nand U22211 (N_22211,N_13077,N_18296);
nand U22212 (N_22212,N_17165,N_16276);
nor U22213 (N_22213,N_13461,N_17600);
nor U22214 (N_22214,N_14890,N_15195);
and U22215 (N_22215,N_14827,N_16567);
nand U22216 (N_22216,N_12553,N_13923);
nor U22217 (N_22217,N_13528,N_13374);
and U22218 (N_22218,N_18706,N_13033);
and U22219 (N_22219,N_17465,N_18636);
and U22220 (N_22220,N_12520,N_15096);
and U22221 (N_22221,N_14595,N_14360);
or U22222 (N_22222,N_15108,N_14705);
nor U22223 (N_22223,N_16484,N_12844);
and U22224 (N_22224,N_12728,N_13984);
nor U22225 (N_22225,N_12503,N_12874);
nand U22226 (N_22226,N_15550,N_15328);
xor U22227 (N_22227,N_15557,N_17728);
and U22228 (N_22228,N_13571,N_16291);
nand U22229 (N_22229,N_18398,N_14833);
and U22230 (N_22230,N_13267,N_13125);
and U22231 (N_22231,N_14832,N_14417);
or U22232 (N_22232,N_12992,N_15963);
xor U22233 (N_22233,N_16935,N_17065);
nand U22234 (N_22234,N_13538,N_15920);
and U22235 (N_22235,N_14964,N_14695);
nor U22236 (N_22236,N_17086,N_18232);
nor U22237 (N_22237,N_13341,N_17060);
and U22238 (N_22238,N_14986,N_12792);
xor U22239 (N_22239,N_16501,N_16298);
or U22240 (N_22240,N_14370,N_14849);
nand U22241 (N_22241,N_14482,N_17773);
nand U22242 (N_22242,N_12796,N_14080);
or U22243 (N_22243,N_14761,N_13039);
and U22244 (N_22244,N_15400,N_14499);
or U22245 (N_22245,N_18641,N_13511);
and U22246 (N_22246,N_16703,N_17111);
nor U22247 (N_22247,N_18583,N_13418);
nor U22248 (N_22248,N_13788,N_17580);
or U22249 (N_22249,N_16128,N_12644);
nor U22250 (N_22250,N_12760,N_16987);
nand U22251 (N_22251,N_16621,N_17291);
or U22252 (N_22252,N_18705,N_15378);
xnor U22253 (N_22253,N_13284,N_17860);
xnor U22254 (N_22254,N_14859,N_18449);
nor U22255 (N_22255,N_12944,N_17239);
nand U22256 (N_22256,N_13099,N_18148);
xnor U22257 (N_22257,N_14919,N_14615);
nor U22258 (N_22258,N_15699,N_13157);
or U22259 (N_22259,N_12724,N_13835);
nand U22260 (N_22260,N_14484,N_14514);
nor U22261 (N_22261,N_16707,N_17911);
nand U22262 (N_22262,N_16440,N_14473);
and U22263 (N_22263,N_13228,N_16623);
nor U22264 (N_22264,N_17125,N_15739);
and U22265 (N_22265,N_14923,N_14558);
nor U22266 (N_22266,N_16670,N_14653);
and U22267 (N_22267,N_17900,N_16836);
or U22268 (N_22268,N_13449,N_13028);
and U22269 (N_22269,N_14588,N_15134);
xor U22270 (N_22270,N_14702,N_14778);
or U22271 (N_22271,N_17285,N_16146);
and U22272 (N_22272,N_18440,N_14986);
or U22273 (N_22273,N_13609,N_16495);
nand U22274 (N_22274,N_14664,N_13038);
nor U22275 (N_22275,N_13876,N_16303);
or U22276 (N_22276,N_17120,N_17674);
or U22277 (N_22277,N_14056,N_14076);
nand U22278 (N_22278,N_16069,N_13122);
and U22279 (N_22279,N_17899,N_16741);
nand U22280 (N_22280,N_14306,N_12816);
and U22281 (N_22281,N_16087,N_14116);
and U22282 (N_22282,N_17441,N_15980);
nor U22283 (N_22283,N_12551,N_12814);
xnor U22284 (N_22284,N_16516,N_15921);
and U22285 (N_22285,N_16688,N_17286);
and U22286 (N_22286,N_17100,N_18062);
and U22287 (N_22287,N_18090,N_14458);
and U22288 (N_22288,N_16717,N_15850);
or U22289 (N_22289,N_18695,N_15221);
nor U22290 (N_22290,N_15611,N_13587);
or U22291 (N_22291,N_15582,N_15543);
nand U22292 (N_22292,N_16366,N_18346);
nor U22293 (N_22293,N_14469,N_16186);
nand U22294 (N_22294,N_16914,N_14849);
and U22295 (N_22295,N_16723,N_16445);
or U22296 (N_22296,N_17807,N_15267);
nor U22297 (N_22297,N_18384,N_14230);
or U22298 (N_22298,N_16850,N_16475);
nand U22299 (N_22299,N_13376,N_17502);
or U22300 (N_22300,N_15778,N_16579);
xor U22301 (N_22301,N_13857,N_14302);
and U22302 (N_22302,N_18523,N_17116);
nand U22303 (N_22303,N_14072,N_17711);
and U22304 (N_22304,N_14135,N_17017);
nand U22305 (N_22305,N_18355,N_15815);
and U22306 (N_22306,N_17575,N_15727);
and U22307 (N_22307,N_13911,N_18746);
and U22308 (N_22308,N_16424,N_17337);
nand U22309 (N_22309,N_14671,N_13058);
or U22310 (N_22310,N_13202,N_16038);
or U22311 (N_22311,N_14359,N_16394);
nor U22312 (N_22312,N_16932,N_15425);
nand U22313 (N_22313,N_17002,N_15708);
and U22314 (N_22314,N_14596,N_13174);
or U22315 (N_22315,N_16475,N_15463);
and U22316 (N_22316,N_18163,N_16219);
nand U22317 (N_22317,N_18358,N_18716);
and U22318 (N_22318,N_15841,N_15281);
nor U22319 (N_22319,N_15357,N_15984);
xor U22320 (N_22320,N_12944,N_15530);
nand U22321 (N_22321,N_13510,N_13832);
and U22322 (N_22322,N_18392,N_13096);
and U22323 (N_22323,N_18668,N_17238);
or U22324 (N_22324,N_18395,N_15205);
nor U22325 (N_22325,N_15829,N_15635);
nor U22326 (N_22326,N_15786,N_17932);
or U22327 (N_22327,N_16986,N_15108);
xnor U22328 (N_22328,N_17694,N_16908);
nor U22329 (N_22329,N_14647,N_18105);
and U22330 (N_22330,N_13392,N_16486);
nand U22331 (N_22331,N_18064,N_18438);
nand U22332 (N_22332,N_14997,N_18536);
nor U22333 (N_22333,N_14848,N_14585);
and U22334 (N_22334,N_14985,N_16685);
and U22335 (N_22335,N_14551,N_13817);
or U22336 (N_22336,N_15036,N_17347);
nand U22337 (N_22337,N_16901,N_12696);
and U22338 (N_22338,N_14807,N_12627);
nor U22339 (N_22339,N_14173,N_15155);
xnor U22340 (N_22340,N_15393,N_14233);
and U22341 (N_22341,N_18618,N_16390);
nor U22342 (N_22342,N_16769,N_12916);
nor U22343 (N_22343,N_15971,N_13765);
nor U22344 (N_22344,N_14017,N_14397);
and U22345 (N_22345,N_15498,N_17013);
and U22346 (N_22346,N_13399,N_16791);
nor U22347 (N_22347,N_15931,N_14664);
nor U22348 (N_22348,N_14106,N_14762);
nor U22349 (N_22349,N_14513,N_14714);
or U22350 (N_22350,N_13450,N_15838);
nand U22351 (N_22351,N_17481,N_14400);
nand U22352 (N_22352,N_15453,N_16011);
and U22353 (N_22353,N_16878,N_12736);
nor U22354 (N_22354,N_18179,N_17654);
or U22355 (N_22355,N_17901,N_16773);
or U22356 (N_22356,N_17892,N_18042);
xnor U22357 (N_22357,N_17999,N_17962);
and U22358 (N_22358,N_16309,N_15680);
nand U22359 (N_22359,N_15138,N_16478);
nor U22360 (N_22360,N_12892,N_18748);
nand U22361 (N_22361,N_12888,N_13446);
nor U22362 (N_22362,N_18459,N_13927);
nand U22363 (N_22363,N_15898,N_15764);
and U22364 (N_22364,N_16727,N_13169);
and U22365 (N_22365,N_16435,N_16715);
nor U22366 (N_22366,N_17554,N_18435);
and U22367 (N_22367,N_14657,N_16342);
nor U22368 (N_22368,N_16144,N_15673);
xor U22369 (N_22369,N_16033,N_15532);
and U22370 (N_22370,N_14915,N_14887);
or U22371 (N_22371,N_12747,N_16416);
xnor U22372 (N_22372,N_12811,N_13316);
nor U22373 (N_22373,N_15542,N_13136);
or U22374 (N_22374,N_17260,N_16455);
nand U22375 (N_22375,N_17386,N_18568);
and U22376 (N_22376,N_12877,N_14175);
and U22377 (N_22377,N_14282,N_13035);
and U22378 (N_22378,N_13051,N_14134);
or U22379 (N_22379,N_17971,N_18613);
nor U22380 (N_22380,N_15351,N_13932);
or U22381 (N_22381,N_15266,N_14117);
nand U22382 (N_22382,N_13435,N_16856);
nand U22383 (N_22383,N_14731,N_16113);
nand U22384 (N_22384,N_15952,N_17166);
and U22385 (N_22385,N_14275,N_13677);
or U22386 (N_22386,N_18711,N_14903);
and U22387 (N_22387,N_16027,N_13017);
nand U22388 (N_22388,N_13231,N_17227);
nand U22389 (N_22389,N_17164,N_14307);
or U22390 (N_22390,N_15548,N_18455);
or U22391 (N_22391,N_15078,N_15275);
or U22392 (N_22392,N_17238,N_13983);
nor U22393 (N_22393,N_12845,N_14093);
or U22394 (N_22394,N_13042,N_17159);
nand U22395 (N_22395,N_17648,N_15593);
nor U22396 (N_22396,N_18372,N_14091);
or U22397 (N_22397,N_17142,N_16233);
nand U22398 (N_22398,N_17128,N_18565);
and U22399 (N_22399,N_16777,N_14745);
nor U22400 (N_22400,N_13741,N_13920);
nand U22401 (N_22401,N_13079,N_17679);
xnor U22402 (N_22402,N_13526,N_16606);
or U22403 (N_22403,N_15057,N_13378);
xor U22404 (N_22404,N_17402,N_14946);
nor U22405 (N_22405,N_17379,N_18066);
nor U22406 (N_22406,N_18341,N_15683);
or U22407 (N_22407,N_16081,N_14308);
or U22408 (N_22408,N_17645,N_18612);
nand U22409 (N_22409,N_13677,N_17988);
or U22410 (N_22410,N_13191,N_13344);
or U22411 (N_22411,N_13974,N_14737);
and U22412 (N_22412,N_13540,N_16623);
nand U22413 (N_22413,N_14447,N_16781);
and U22414 (N_22414,N_14960,N_17756);
nand U22415 (N_22415,N_16433,N_17200);
and U22416 (N_22416,N_13695,N_15998);
nand U22417 (N_22417,N_14073,N_13891);
or U22418 (N_22418,N_14396,N_15986);
nand U22419 (N_22419,N_15510,N_17309);
nor U22420 (N_22420,N_12716,N_15824);
and U22421 (N_22421,N_13985,N_14905);
and U22422 (N_22422,N_12670,N_12920);
nor U22423 (N_22423,N_15724,N_16720);
xor U22424 (N_22424,N_15775,N_17049);
nor U22425 (N_22425,N_12900,N_12606);
and U22426 (N_22426,N_13070,N_17814);
nand U22427 (N_22427,N_13618,N_15448);
and U22428 (N_22428,N_13789,N_18056);
and U22429 (N_22429,N_13116,N_14057);
and U22430 (N_22430,N_16352,N_16181);
nand U22431 (N_22431,N_15823,N_12710);
nor U22432 (N_22432,N_16277,N_17304);
nor U22433 (N_22433,N_18190,N_16109);
and U22434 (N_22434,N_13665,N_16967);
or U22435 (N_22435,N_14588,N_18654);
or U22436 (N_22436,N_14493,N_17001);
or U22437 (N_22437,N_18038,N_14054);
nand U22438 (N_22438,N_14763,N_17303);
nand U22439 (N_22439,N_16306,N_17113);
and U22440 (N_22440,N_14259,N_18052);
and U22441 (N_22441,N_17579,N_17983);
and U22442 (N_22442,N_14571,N_17824);
nand U22443 (N_22443,N_18171,N_13484);
nand U22444 (N_22444,N_18194,N_14014);
nand U22445 (N_22445,N_14760,N_16287);
nor U22446 (N_22446,N_12803,N_15730);
nand U22447 (N_22447,N_15594,N_14195);
nor U22448 (N_22448,N_12625,N_17124);
nand U22449 (N_22449,N_15136,N_13371);
nor U22450 (N_22450,N_15855,N_15395);
nand U22451 (N_22451,N_16832,N_15609);
or U22452 (N_22452,N_18472,N_18340);
and U22453 (N_22453,N_15625,N_13433);
nand U22454 (N_22454,N_14754,N_14610);
nor U22455 (N_22455,N_14691,N_14553);
xnor U22456 (N_22456,N_17570,N_16321);
or U22457 (N_22457,N_16843,N_15020);
or U22458 (N_22458,N_13535,N_18648);
nor U22459 (N_22459,N_16845,N_17002);
xor U22460 (N_22460,N_16800,N_18719);
nand U22461 (N_22461,N_14000,N_14940);
nand U22462 (N_22462,N_18689,N_17601);
and U22463 (N_22463,N_14837,N_13859);
nor U22464 (N_22464,N_18018,N_15611);
or U22465 (N_22465,N_14832,N_16191);
and U22466 (N_22466,N_16165,N_17359);
or U22467 (N_22467,N_14783,N_17798);
or U22468 (N_22468,N_12929,N_15464);
or U22469 (N_22469,N_14276,N_13893);
and U22470 (N_22470,N_12544,N_18378);
and U22471 (N_22471,N_16517,N_16840);
nand U22472 (N_22472,N_16707,N_14258);
nor U22473 (N_22473,N_13085,N_15112);
and U22474 (N_22474,N_14912,N_16482);
nand U22475 (N_22475,N_18368,N_14949);
nand U22476 (N_22476,N_17540,N_16567);
nand U22477 (N_22477,N_12730,N_16474);
or U22478 (N_22478,N_15507,N_15792);
and U22479 (N_22479,N_16961,N_13404);
nor U22480 (N_22480,N_12866,N_18503);
nand U22481 (N_22481,N_14821,N_15405);
nand U22482 (N_22482,N_16465,N_13090);
nor U22483 (N_22483,N_15054,N_17617);
nand U22484 (N_22484,N_13661,N_16587);
and U22485 (N_22485,N_17674,N_12908);
and U22486 (N_22486,N_13364,N_15962);
nand U22487 (N_22487,N_16868,N_14443);
nor U22488 (N_22488,N_15199,N_16518);
xor U22489 (N_22489,N_17014,N_15625);
nor U22490 (N_22490,N_17587,N_13424);
nand U22491 (N_22491,N_15432,N_15537);
or U22492 (N_22492,N_12920,N_13838);
nor U22493 (N_22493,N_13463,N_16614);
nor U22494 (N_22494,N_12539,N_14421);
nor U22495 (N_22495,N_17945,N_14458);
nand U22496 (N_22496,N_16138,N_13520);
and U22497 (N_22497,N_13466,N_13881);
and U22498 (N_22498,N_17252,N_15510);
nand U22499 (N_22499,N_17378,N_17991);
nor U22500 (N_22500,N_12746,N_12513);
and U22501 (N_22501,N_15077,N_16111);
nand U22502 (N_22502,N_14245,N_12623);
nand U22503 (N_22503,N_16472,N_17767);
and U22504 (N_22504,N_15321,N_17078);
or U22505 (N_22505,N_18284,N_15811);
nor U22506 (N_22506,N_13510,N_16043);
or U22507 (N_22507,N_16852,N_16144);
or U22508 (N_22508,N_16786,N_17991);
and U22509 (N_22509,N_16417,N_12521);
and U22510 (N_22510,N_18675,N_15656);
nand U22511 (N_22511,N_16581,N_17061);
and U22512 (N_22512,N_16492,N_15686);
nor U22513 (N_22513,N_12689,N_15446);
or U22514 (N_22514,N_13168,N_12968);
nand U22515 (N_22515,N_12779,N_13283);
or U22516 (N_22516,N_18391,N_13872);
xnor U22517 (N_22517,N_17702,N_17880);
nand U22518 (N_22518,N_17673,N_14262);
nand U22519 (N_22519,N_18614,N_12683);
and U22520 (N_22520,N_16498,N_16147);
nor U22521 (N_22521,N_16766,N_16960);
nand U22522 (N_22522,N_17494,N_16210);
nand U22523 (N_22523,N_13184,N_12636);
nand U22524 (N_22524,N_15861,N_15120);
nand U22525 (N_22525,N_14596,N_12790);
nand U22526 (N_22526,N_13588,N_17665);
and U22527 (N_22527,N_17450,N_18176);
xor U22528 (N_22528,N_12990,N_13616);
and U22529 (N_22529,N_17087,N_17975);
nor U22530 (N_22530,N_15330,N_15275);
and U22531 (N_22531,N_18483,N_15973);
nand U22532 (N_22532,N_16199,N_12904);
or U22533 (N_22533,N_14444,N_17585);
nor U22534 (N_22534,N_14796,N_18489);
nand U22535 (N_22535,N_15053,N_17844);
nor U22536 (N_22536,N_14252,N_14639);
nor U22537 (N_22537,N_13738,N_14677);
or U22538 (N_22538,N_16963,N_14534);
nand U22539 (N_22539,N_13169,N_15238);
nand U22540 (N_22540,N_17522,N_17833);
nor U22541 (N_22541,N_17502,N_13892);
nand U22542 (N_22542,N_17096,N_12993);
nor U22543 (N_22543,N_15167,N_13469);
and U22544 (N_22544,N_17990,N_16303);
nor U22545 (N_22545,N_14384,N_15995);
nand U22546 (N_22546,N_16746,N_14091);
nand U22547 (N_22547,N_12523,N_12761);
and U22548 (N_22548,N_16868,N_16929);
or U22549 (N_22549,N_14891,N_18373);
or U22550 (N_22550,N_14930,N_13702);
nor U22551 (N_22551,N_14962,N_15335);
or U22552 (N_22552,N_14315,N_15818);
nor U22553 (N_22553,N_14363,N_16402);
nor U22554 (N_22554,N_12704,N_13078);
or U22555 (N_22555,N_17977,N_16413);
nor U22556 (N_22556,N_13503,N_14204);
nand U22557 (N_22557,N_15521,N_14643);
or U22558 (N_22558,N_13918,N_13348);
or U22559 (N_22559,N_17657,N_12653);
xnor U22560 (N_22560,N_17267,N_17308);
nor U22561 (N_22561,N_14968,N_17454);
xnor U22562 (N_22562,N_16599,N_13863);
xor U22563 (N_22563,N_16976,N_17460);
nand U22564 (N_22564,N_14357,N_17233);
nor U22565 (N_22565,N_13837,N_14716);
and U22566 (N_22566,N_12920,N_18312);
and U22567 (N_22567,N_13685,N_13246);
and U22568 (N_22568,N_14941,N_14322);
or U22569 (N_22569,N_14121,N_16170);
or U22570 (N_22570,N_14067,N_13105);
nand U22571 (N_22571,N_16434,N_13820);
and U22572 (N_22572,N_16384,N_14092);
and U22573 (N_22573,N_16522,N_14022);
or U22574 (N_22574,N_14526,N_18654);
nand U22575 (N_22575,N_15910,N_18039);
nand U22576 (N_22576,N_15158,N_15359);
nor U22577 (N_22577,N_14028,N_13323);
nand U22578 (N_22578,N_13633,N_18356);
nor U22579 (N_22579,N_16662,N_15801);
nand U22580 (N_22580,N_13408,N_16693);
nor U22581 (N_22581,N_18682,N_14574);
xor U22582 (N_22582,N_16591,N_18347);
or U22583 (N_22583,N_14440,N_15646);
or U22584 (N_22584,N_15866,N_14892);
or U22585 (N_22585,N_18299,N_18175);
xor U22586 (N_22586,N_13301,N_16131);
and U22587 (N_22587,N_13024,N_14215);
and U22588 (N_22588,N_16217,N_18053);
and U22589 (N_22589,N_14117,N_15221);
or U22590 (N_22590,N_13790,N_13474);
or U22591 (N_22591,N_14304,N_14632);
and U22592 (N_22592,N_14297,N_14571);
and U22593 (N_22593,N_18549,N_13494);
nor U22594 (N_22594,N_14784,N_14352);
nor U22595 (N_22595,N_14493,N_16970);
and U22596 (N_22596,N_16473,N_16553);
or U22597 (N_22597,N_14399,N_14944);
and U22598 (N_22598,N_16597,N_13213);
xor U22599 (N_22599,N_14626,N_17441);
and U22600 (N_22600,N_17240,N_18123);
nor U22601 (N_22601,N_17895,N_15589);
nor U22602 (N_22602,N_13900,N_12933);
and U22603 (N_22603,N_16133,N_14481);
nor U22604 (N_22604,N_12925,N_14530);
or U22605 (N_22605,N_15528,N_13512);
nor U22606 (N_22606,N_16984,N_16621);
and U22607 (N_22607,N_16338,N_13190);
or U22608 (N_22608,N_13833,N_14546);
or U22609 (N_22609,N_16026,N_17477);
or U22610 (N_22610,N_13049,N_16178);
or U22611 (N_22611,N_14884,N_16237);
nor U22612 (N_22612,N_16980,N_13972);
and U22613 (N_22613,N_18322,N_18329);
nor U22614 (N_22614,N_13258,N_16193);
nand U22615 (N_22615,N_14709,N_13195);
nand U22616 (N_22616,N_13269,N_16194);
or U22617 (N_22617,N_13896,N_15916);
or U22618 (N_22618,N_16629,N_15395);
nand U22619 (N_22619,N_17165,N_15646);
nand U22620 (N_22620,N_14386,N_15574);
nand U22621 (N_22621,N_17150,N_14772);
and U22622 (N_22622,N_13525,N_17260);
and U22623 (N_22623,N_13165,N_12538);
nand U22624 (N_22624,N_18471,N_13326);
or U22625 (N_22625,N_17356,N_13761);
nor U22626 (N_22626,N_13855,N_14367);
nor U22627 (N_22627,N_13227,N_17578);
nand U22628 (N_22628,N_13379,N_18114);
nor U22629 (N_22629,N_15373,N_13323);
and U22630 (N_22630,N_17753,N_15948);
nand U22631 (N_22631,N_14100,N_14474);
nor U22632 (N_22632,N_14954,N_13381);
xnor U22633 (N_22633,N_14346,N_15061);
nor U22634 (N_22634,N_15498,N_14990);
or U22635 (N_22635,N_15404,N_16691);
xor U22636 (N_22636,N_15545,N_15165);
nand U22637 (N_22637,N_12504,N_14392);
and U22638 (N_22638,N_14790,N_12762);
nor U22639 (N_22639,N_13859,N_13188);
nand U22640 (N_22640,N_15814,N_18262);
nor U22641 (N_22641,N_16816,N_14209);
or U22642 (N_22642,N_17399,N_18188);
nand U22643 (N_22643,N_16838,N_13452);
nor U22644 (N_22644,N_14607,N_13881);
nand U22645 (N_22645,N_13289,N_15715);
xor U22646 (N_22646,N_18082,N_15985);
nand U22647 (N_22647,N_14346,N_17400);
and U22648 (N_22648,N_17532,N_15125);
and U22649 (N_22649,N_15743,N_12768);
and U22650 (N_22650,N_17686,N_16702);
nand U22651 (N_22651,N_15822,N_16526);
nor U22652 (N_22652,N_18568,N_13579);
nand U22653 (N_22653,N_16083,N_13456);
or U22654 (N_22654,N_14547,N_15445);
nand U22655 (N_22655,N_14985,N_17307);
or U22656 (N_22656,N_16542,N_15938);
nand U22657 (N_22657,N_12828,N_16725);
nand U22658 (N_22658,N_18578,N_17738);
or U22659 (N_22659,N_14925,N_17491);
or U22660 (N_22660,N_16917,N_12793);
or U22661 (N_22661,N_14530,N_13419);
nand U22662 (N_22662,N_13848,N_12870);
or U22663 (N_22663,N_16290,N_16451);
nand U22664 (N_22664,N_12934,N_12887);
and U22665 (N_22665,N_14717,N_18295);
nand U22666 (N_22666,N_12682,N_14499);
or U22667 (N_22667,N_16866,N_17083);
nor U22668 (N_22668,N_15444,N_13403);
or U22669 (N_22669,N_12779,N_18315);
and U22670 (N_22670,N_18725,N_18027);
xor U22671 (N_22671,N_17868,N_14766);
or U22672 (N_22672,N_14197,N_18312);
nor U22673 (N_22673,N_16211,N_13529);
and U22674 (N_22674,N_16172,N_17384);
and U22675 (N_22675,N_16332,N_15443);
and U22676 (N_22676,N_12809,N_17118);
and U22677 (N_22677,N_14846,N_17581);
and U22678 (N_22678,N_16333,N_14163);
or U22679 (N_22679,N_15303,N_18341);
and U22680 (N_22680,N_12912,N_14427);
or U22681 (N_22681,N_13961,N_15458);
and U22682 (N_22682,N_18048,N_15769);
and U22683 (N_22683,N_16455,N_14338);
xnor U22684 (N_22684,N_16614,N_14368);
or U22685 (N_22685,N_16163,N_18575);
nand U22686 (N_22686,N_15427,N_15967);
nor U22687 (N_22687,N_18260,N_15265);
nor U22688 (N_22688,N_18178,N_15325);
nand U22689 (N_22689,N_12664,N_16887);
and U22690 (N_22690,N_16899,N_15156);
xnor U22691 (N_22691,N_13225,N_16643);
nand U22692 (N_22692,N_15493,N_14891);
and U22693 (N_22693,N_15836,N_16574);
nand U22694 (N_22694,N_15280,N_13106);
nor U22695 (N_22695,N_18029,N_12888);
nor U22696 (N_22696,N_14225,N_13911);
and U22697 (N_22697,N_16466,N_18224);
nor U22698 (N_22698,N_16833,N_17903);
nor U22699 (N_22699,N_16543,N_13063);
or U22700 (N_22700,N_16366,N_12820);
nor U22701 (N_22701,N_18248,N_14372);
and U22702 (N_22702,N_18372,N_15427);
and U22703 (N_22703,N_13229,N_13859);
nand U22704 (N_22704,N_14307,N_17201);
nor U22705 (N_22705,N_14774,N_15070);
nand U22706 (N_22706,N_16305,N_14415);
nand U22707 (N_22707,N_13293,N_14312);
xor U22708 (N_22708,N_13682,N_18101);
or U22709 (N_22709,N_15428,N_16324);
or U22710 (N_22710,N_15254,N_15423);
xnor U22711 (N_22711,N_15274,N_14052);
xnor U22712 (N_22712,N_17992,N_17789);
nand U22713 (N_22713,N_17954,N_15438);
and U22714 (N_22714,N_13668,N_18363);
nand U22715 (N_22715,N_16325,N_18572);
and U22716 (N_22716,N_16294,N_12585);
nor U22717 (N_22717,N_16760,N_13996);
nand U22718 (N_22718,N_13056,N_17787);
or U22719 (N_22719,N_16731,N_17775);
xor U22720 (N_22720,N_15216,N_13090);
and U22721 (N_22721,N_16175,N_14707);
nor U22722 (N_22722,N_16208,N_17338);
nor U22723 (N_22723,N_15992,N_15298);
nand U22724 (N_22724,N_14398,N_13809);
xnor U22725 (N_22725,N_16109,N_14393);
and U22726 (N_22726,N_15653,N_16430);
and U22727 (N_22727,N_14417,N_17370);
or U22728 (N_22728,N_18060,N_17479);
nand U22729 (N_22729,N_12814,N_15146);
or U22730 (N_22730,N_16301,N_17109);
xor U22731 (N_22731,N_18138,N_17379);
and U22732 (N_22732,N_18325,N_13595);
and U22733 (N_22733,N_14555,N_16176);
nor U22734 (N_22734,N_16803,N_14588);
and U22735 (N_22735,N_15165,N_16461);
or U22736 (N_22736,N_14209,N_15540);
and U22737 (N_22737,N_13166,N_16420);
or U22738 (N_22738,N_18141,N_13526);
nor U22739 (N_22739,N_16985,N_13285);
or U22740 (N_22740,N_12917,N_15758);
and U22741 (N_22741,N_12566,N_14285);
and U22742 (N_22742,N_16497,N_13316);
or U22743 (N_22743,N_16722,N_14454);
nor U22744 (N_22744,N_13234,N_16678);
or U22745 (N_22745,N_17994,N_18267);
or U22746 (N_22746,N_16892,N_14420);
xor U22747 (N_22747,N_14863,N_17993);
nor U22748 (N_22748,N_12790,N_15292);
or U22749 (N_22749,N_18417,N_14263);
nand U22750 (N_22750,N_18542,N_12806);
and U22751 (N_22751,N_14787,N_16876);
and U22752 (N_22752,N_14458,N_13881);
and U22753 (N_22753,N_15809,N_12979);
and U22754 (N_22754,N_15149,N_16156);
nor U22755 (N_22755,N_17920,N_15209);
nor U22756 (N_22756,N_17875,N_12805);
nor U22757 (N_22757,N_12985,N_17674);
nor U22758 (N_22758,N_13380,N_13297);
nand U22759 (N_22759,N_18020,N_13490);
nand U22760 (N_22760,N_16565,N_16554);
or U22761 (N_22761,N_15706,N_15177);
xnor U22762 (N_22762,N_13587,N_15825);
and U22763 (N_22763,N_18189,N_17698);
or U22764 (N_22764,N_18442,N_18618);
and U22765 (N_22765,N_17121,N_16798);
nand U22766 (N_22766,N_13246,N_15650);
or U22767 (N_22767,N_12739,N_18420);
or U22768 (N_22768,N_17880,N_16712);
or U22769 (N_22769,N_14359,N_12928);
nand U22770 (N_22770,N_16376,N_15029);
nand U22771 (N_22771,N_12835,N_15196);
and U22772 (N_22772,N_16332,N_18211);
and U22773 (N_22773,N_14168,N_13506);
or U22774 (N_22774,N_13599,N_17004);
nor U22775 (N_22775,N_18647,N_15184);
or U22776 (N_22776,N_16184,N_16536);
xor U22777 (N_22777,N_12711,N_17261);
nor U22778 (N_22778,N_17113,N_15357);
nand U22779 (N_22779,N_15691,N_18201);
or U22780 (N_22780,N_15655,N_16324);
nor U22781 (N_22781,N_16088,N_14433);
nand U22782 (N_22782,N_18132,N_15632);
nand U22783 (N_22783,N_16426,N_18639);
and U22784 (N_22784,N_18211,N_15845);
or U22785 (N_22785,N_15844,N_17629);
nand U22786 (N_22786,N_13257,N_15245);
and U22787 (N_22787,N_12592,N_17863);
xnor U22788 (N_22788,N_14525,N_14651);
nor U22789 (N_22789,N_12764,N_16104);
nand U22790 (N_22790,N_14312,N_16548);
or U22791 (N_22791,N_17102,N_17598);
and U22792 (N_22792,N_16109,N_14501);
nor U22793 (N_22793,N_17528,N_17047);
nor U22794 (N_22794,N_16389,N_16484);
nor U22795 (N_22795,N_15446,N_18646);
or U22796 (N_22796,N_17807,N_15817);
or U22797 (N_22797,N_15649,N_18675);
and U22798 (N_22798,N_13532,N_15372);
and U22799 (N_22799,N_17888,N_17398);
and U22800 (N_22800,N_13127,N_18025);
and U22801 (N_22801,N_13966,N_13478);
and U22802 (N_22802,N_13698,N_17423);
nand U22803 (N_22803,N_13803,N_18056);
nor U22804 (N_22804,N_13761,N_12999);
nand U22805 (N_22805,N_18311,N_16616);
or U22806 (N_22806,N_14919,N_12841);
or U22807 (N_22807,N_13507,N_13112);
nor U22808 (N_22808,N_15089,N_15495);
or U22809 (N_22809,N_14748,N_18411);
nor U22810 (N_22810,N_14829,N_17563);
nor U22811 (N_22811,N_17130,N_14949);
and U22812 (N_22812,N_14010,N_14107);
nand U22813 (N_22813,N_17398,N_13879);
or U22814 (N_22814,N_15963,N_12944);
and U22815 (N_22815,N_13700,N_15430);
or U22816 (N_22816,N_16275,N_14237);
nand U22817 (N_22817,N_12811,N_14031);
and U22818 (N_22818,N_14368,N_16341);
or U22819 (N_22819,N_15646,N_15857);
nand U22820 (N_22820,N_17011,N_16750);
nor U22821 (N_22821,N_18322,N_18195);
nand U22822 (N_22822,N_16369,N_16381);
and U22823 (N_22823,N_14871,N_16502);
or U22824 (N_22824,N_15024,N_18319);
nand U22825 (N_22825,N_14737,N_13248);
nand U22826 (N_22826,N_17250,N_17447);
or U22827 (N_22827,N_15708,N_16566);
and U22828 (N_22828,N_18129,N_18739);
nand U22829 (N_22829,N_17265,N_13279);
and U22830 (N_22830,N_13687,N_12689);
or U22831 (N_22831,N_12809,N_15927);
and U22832 (N_22832,N_15016,N_16242);
nand U22833 (N_22833,N_13568,N_14470);
and U22834 (N_22834,N_15651,N_16410);
nand U22835 (N_22835,N_15434,N_12828);
and U22836 (N_22836,N_16838,N_13838);
xnor U22837 (N_22837,N_12957,N_16770);
and U22838 (N_22838,N_18447,N_13952);
and U22839 (N_22839,N_16560,N_16575);
and U22840 (N_22840,N_15209,N_16256);
or U22841 (N_22841,N_14678,N_15943);
nor U22842 (N_22842,N_18664,N_18515);
or U22843 (N_22843,N_14347,N_16834);
xor U22844 (N_22844,N_12941,N_12571);
or U22845 (N_22845,N_14888,N_17318);
nor U22846 (N_22846,N_14133,N_13268);
or U22847 (N_22847,N_13345,N_16120);
nor U22848 (N_22848,N_17831,N_18264);
nand U22849 (N_22849,N_17587,N_17138);
or U22850 (N_22850,N_13018,N_14291);
or U22851 (N_22851,N_14850,N_17690);
or U22852 (N_22852,N_18687,N_17336);
nor U22853 (N_22853,N_15163,N_14917);
or U22854 (N_22854,N_15482,N_16002);
xnor U22855 (N_22855,N_17145,N_18697);
nand U22856 (N_22856,N_12927,N_12605);
and U22857 (N_22857,N_16851,N_14340);
nor U22858 (N_22858,N_14888,N_13255);
or U22859 (N_22859,N_13817,N_12603);
nor U22860 (N_22860,N_13488,N_15782);
nand U22861 (N_22861,N_15374,N_17394);
or U22862 (N_22862,N_15296,N_15394);
nor U22863 (N_22863,N_12614,N_13977);
nor U22864 (N_22864,N_12639,N_17942);
or U22865 (N_22865,N_15962,N_14725);
and U22866 (N_22866,N_12672,N_13640);
nand U22867 (N_22867,N_17345,N_16443);
or U22868 (N_22868,N_14952,N_14615);
nor U22869 (N_22869,N_17024,N_14466);
nand U22870 (N_22870,N_15559,N_16674);
nor U22871 (N_22871,N_15500,N_16803);
or U22872 (N_22872,N_15566,N_18479);
nor U22873 (N_22873,N_14518,N_16174);
and U22874 (N_22874,N_18341,N_14275);
or U22875 (N_22875,N_16675,N_17200);
xor U22876 (N_22876,N_16919,N_12852);
and U22877 (N_22877,N_18652,N_16181);
or U22878 (N_22878,N_16469,N_18158);
nand U22879 (N_22879,N_18635,N_14644);
and U22880 (N_22880,N_17364,N_14798);
or U22881 (N_22881,N_13843,N_18168);
xor U22882 (N_22882,N_17223,N_13080);
and U22883 (N_22883,N_12502,N_16600);
nor U22884 (N_22884,N_17484,N_12754);
and U22885 (N_22885,N_18574,N_13229);
and U22886 (N_22886,N_14598,N_15866);
or U22887 (N_22887,N_18011,N_15254);
and U22888 (N_22888,N_16709,N_15865);
and U22889 (N_22889,N_13647,N_12836);
xnor U22890 (N_22890,N_13499,N_18632);
nand U22891 (N_22891,N_16389,N_15870);
and U22892 (N_22892,N_17917,N_16907);
and U22893 (N_22893,N_17875,N_13237);
xnor U22894 (N_22894,N_15814,N_13389);
or U22895 (N_22895,N_13690,N_13350);
or U22896 (N_22896,N_17822,N_13812);
and U22897 (N_22897,N_15251,N_13107);
nand U22898 (N_22898,N_13713,N_18183);
xor U22899 (N_22899,N_15034,N_14599);
nand U22900 (N_22900,N_13698,N_12528);
nand U22901 (N_22901,N_15842,N_16911);
and U22902 (N_22902,N_17475,N_16225);
or U22903 (N_22903,N_15074,N_17089);
or U22904 (N_22904,N_18252,N_14558);
and U22905 (N_22905,N_17476,N_14356);
nor U22906 (N_22906,N_17135,N_16317);
or U22907 (N_22907,N_13825,N_16626);
nand U22908 (N_22908,N_17675,N_14020);
or U22909 (N_22909,N_14161,N_16225);
and U22910 (N_22910,N_13634,N_15988);
nand U22911 (N_22911,N_15490,N_13214);
nor U22912 (N_22912,N_18744,N_16827);
nand U22913 (N_22913,N_17851,N_13286);
or U22914 (N_22914,N_15205,N_14465);
nand U22915 (N_22915,N_17103,N_15749);
or U22916 (N_22916,N_18110,N_13044);
and U22917 (N_22917,N_13830,N_12993);
or U22918 (N_22918,N_17098,N_15364);
nand U22919 (N_22919,N_16425,N_17248);
or U22920 (N_22920,N_14746,N_15394);
and U22921 (N_22921,N_18725,N_13966);
or U22922 (N_22922,N_15843,N_14995);
and U22923 (N_22923,N_18436,N_13493);
or U22924 (N_22924,N_12983,N_16898);
and U22925 (N_22925,N_13277,N_13384);
nor U22926 (N_22926,N_16139,N_13163);
xnor U22927 (N_22927,N_15960,N_15209);
nor U22928 (N_22928,N_13856,N_17622);
and U22929 (N_22929,N_12778,N_15705);
nor U22930 (N_22930,N_12905,N_14048);
xnor U22931 (N_22931,N_17194,N_16063);
nand U22932 (N_22932,N_17829,N_17581);
nor U22933 (N_22933,N_15243,N_16852);
nor U22934 (N_22934,N_13497,N_13484);
nand U22935 (N_22935,N_17920,N_18466);
nor U22936 (N_22936,N_14903,N_16778);
and U22937 (N_22937,N_16026,N_18618);
and U22938 (N_22938,N_14517,N_15823);
and U22939 (N_22939,N_17789,N_14594);
nand U22940 (N_22940,N_17806,N_15719);
or U22941 (N_22941,N_18540,N_17238);
nand U22942 (N_22942,N_17834,N_16516);
nor U22943 (N_22943,N_17887,N_18161);
or U22944 (N_22944,N_17607,N_13795);
nand U22945 (N_22945,N_14847,N_15230);
nor U22946 (N_22946,N_12510,N_15769);
xor U22947 (N_22947,N_15541,N_18512);
nor U22948 (N_22948,N_18580,N_13273);
nand U22949 (N_22949,N_16565,N_17632);
nor U22950 (N_22950,N_18707,N_18709);
xnor U22951 (N_22951,N_16326,N_12954);
and U22952 (N_22952,N_17445,N_13651);
nand U22953 (N_22953,N_15132,N_15087);
and U22954 (N_22954,N_15592,N_16452);
nand U22955 (N_22955,N_18406,N_14444);
or U22956 (N_22956,N_15730,N_13533);
and U22957 (N_22957,N_17961,N_13923);
and U22958 (N_22958,N_13476,N_14537);
xnor U22959 (N_22959,N_12833,N_18073);
nor U22960 (N_22960,N_17730,N_16585);
nor U22961 (N_22961,N_15587,N_14594);
and U22962 (N_22962,N_17532,N_17331);
and U22963 (N_22963,N_17171,N_13179);
or U22964 (N_22964,N_17458,N_16230);
and U22965 (N_22965,N_16920,N_15161);
xnor U22966 (N_22966,N_16612,N_13674);
and U22967 (N_22967,N_14704,N_16244);
nand U22968 (N_22968,N_14535,N_16426);
nand U22969 (N_22969,N_12857,N_15943);
nand U22970 (N_22970,N_18180,N_17997);
nand U22971 (N_22971,N_17620,N_18521);
and U22972 (N_22972,N_17540,N_14457);
nor U22973 (N_22973,N_16340,N_15152);
xnor U22974 (N_22974,N_16824,N_15697);
and U22975 (N_22975,N_17236,N_16438);
nand U22976 (N_22976,N_13535,N_14343);
nor U22977 (N_22977,N_16131,N_18080);
nor U22978 (N_22978,N_13855,N_13495);
nor U22979 (N_22979,N_12743,N_17772);
and U22980 (N_22980,N_16945,N_18157);
or U22981 (N_22981,N_18019,N_16745);
or U22982 (N_22982,N_18735,N_13087);
and U22983 (N_22983,N_14469,N_14018);
and U22984 (N_22984,N_16969,N_13172);
and U22985 (N_22985,N_18038,N_16943);
nor U22986 (N_22986,N_15914,N_16615);
and U22987 (N_22987,N_14385,N_12708);
or U22988 (N_22988,N_15455,N_13124);
nand U22989 (N_22989,N_14167,N_17280);
nor U22990 (N_22990,N_12606,N_16183);
nor U22991 (N_22991,N_15270,N_13901);
nor U22992 (N_22992,N_15895,N_13524);
nor U22993 (N_22993,N_16334,N_15304);
nand U22994 (N_22994,N_17607,N_16420);
nor U22995 (N_22995,N_12541,N_14342);
nand U22996 (N_22996,N_14766,N_17650);
and U22997 (N_22997,N_16800,N_17791);
nor U22998 (N_22998,N_15534,N_15983);
nor U22999 (N_22999,N_15861,N_14693);
and U23000 (N_23000,N_16085,N_14980);
or U23001 (N_23001,N_14941,N_13300);
nand U23002 (N_23002,N_16988,N_15722);
or U23003 (N_23003,N_13549,N_16445);
nor U23004 (N_23004,N_17938,N_17144);
or U23005 (N_23005,N_15484,N_13715);
nand U23006 (N_23006,N_15916,N_12709);
nand U23007 (N_23007,N_12558,N_15234);
nand U23008 (N_23008,N_14833,N_18067);
nand U23009 (N_23009,N_14320,N_16250);
nand U23010 (N_23010,N_12949,N_18630);
nand U23011 (N_23011,N_17520,N_17414);
nand U23012 (N_23012,N_16823,N_16560);
nand U23013 (N_23013,N_12769,N_17385);
nor U23014 (N_23014,N_17865,N_14214);
and U23015 (N_23015,N_16214,N_17373);
and U23016 (N_23016,N_18242,N_16943);
and U23017 (N_23017,N_16893,N_18042);
nor U23018 (N_23018,N_13225,N_15731);
nor U23019 (N_23019,N_17545,N_13437);
xnor U23020 (N_23020,N_15595,N_17690);
nor U23021 (N_23021,N_14540,N_17559);
nand U23022 (N_23022,N_17534,N_18314);
nand U23023 (N_23023,N_16924,N_14747);
nor U23024 (N_23024,N_15279,N_16753);
or U23025 (N_23025,N_12530,N_17073);
nor U23026 (N_23026,N_14556,N_15060);
nor U23027 (N_23027,N_12515,N_18619);
nor U23028 (N_23028,N_16199,N_16703);
or U23029 (N_23029,N_17219,N_13676);
nand U23030 (N_23030,N_14098,N_18302);
or U23031 (N_23031,N_15316,N_14289);
or U23032 (N_23032,N_15823,N_14650);
and U23033 (N_23033,N_17000,N_16897);
nor U23034 (N_23034,N_16828,N_18306);
nor U23035 (N_23035,N_17915,N_15941);
or U23036 (N_23036,N_17125,N_12543);
or U23037 (N_23037,N_15378,N_18618);
nand U23038 (N_23038,N_15516,N_16993);
nor U23039 (N_23039,N_17979,N_18091);
xnor U23040 (N_23040,N_14300,N_14856);
nor U23041 (N_23041,N_14337,N_14231);
nor U23042 (N_23042,N_14763,N_15399);
and U23043 (N_23043,N_16637,N_14686);
and U23044 (N_23044,N_14894,N_16789);
nor U23045 (N_23045,N_12879,N_15238);
nor U23046 (N_23046,N_14836,N_14692);
and U23047 (N_23047,N_15297,N_16686);
xnor U23048 (N_23048,N_14690,N_13102);
nor U23049 (N_23049,N_14447,N_13234);
and U23050 (N_23050,N_15690,N_15302);
xor U23051 (N_23051,N_16847,N_17969);
nand U23052 (N_23052,N_12523,N_16940);
nand U23053 (N_23053,N_13361,N_13469);
or U23054 (N_23054,N_18170,N_12796);
nand U23055 (N_23055,N_17917,N_18577);
xnor U23056 (N_23056,N_18714,N_16858);
or U23057 (N_23057,N_16336,N_16834);
nor U23058 (N_23058,N_15943,N_12781);
nand U23059 (N_23059,N_18505,N_15535);
nand U23060 (N_23060,N_14716,N_17920);
or U23061 (N_23061,N_13843,N_14424);
nor U23062 (N_23062,N_14667,N_17775);
nor U23063 (N_23063,N_12632,N_16391);
nor U23064 (N_23064,N_17832,N_12598);
or U23065 (N_23065,N_15438,N_14110);
and U23066 (N_23066,N_13931,N_17203);
or U23067 (N_23067,N_14617,N_13817);
nor U23068 (N_23068,N_15330,N_18175);
nand U23069 (N_23069,N_13595,N_12789);
nand U23070 (N_23070,N_18065,N_15285);
and U23071 (N_23071,N_18329,N_12538);
or U23072 (N_23072,N_18230,N_14498);
nand U23073 (N_23073,N_15515,N_12674);
or U23074 (N_23074,N_16072,N_17850);
and U23075 (N_23075,N_14357,N_15114);
nor U23076 (N_23076,N_16869,N_15918);
xnor U23077 (N_23077,N_16657,N_14009);
nand U23078 (N_23078,N_15037,N_15978);
or U23079 (N_23079,N_12665,N_14472);
nand U23080 (N_23080,N_14123,N_16201);
xnor U23081 (N_23081,N_12865,N_15133);
xor U23082 (N_23082,N_18172,N_18747);
and U23083 (N_23083,N_16889,N_16527);
and U23084 (N_23084,N_17450,N_16491);
nor U23085 (N_23085,N_18350,N_14335);
nor U23086 (N_23086,N_16396,N_15013);
nand U23087 (N_23087,N_18534,N_18180);
or U23088 (N_23088,N_15369,N_14632);
nand U23089 (N_23089,N_12908,N_17445);
and U23090 (N_23090,N_15999,N_16587);
xnor U23091 (N_23091,N_18676,N_15307);
nand U23092 (N_23092,N_17763,N_13296);
xnor U23093 (N_23093,N_14448,N_15865);
or U23094 (N_23094,N_16851,N_17153);
and U23095 (N_23095,N_14070,N_17058);
and U23096 (N_23096,N_18393,N_13313);
nand U23097 (N_23097,N_15373,N_14647);
nand U23098 (N_23098,N_17879,N_16739);
xnor U23099 (N_23099,N_15335,N_16135);
or U23100 (N_23100,N_13739,N_16904);
or U23101 (N_23101,N_12815,N_13769);
nand U23102 (N_23102,N_18558,N_16954);
nor U23103 (N_23103,N_15551,N_15643);
nor U23104 (N_23104,N_13639,N_16727);
and U23105 (N_23105,N_18055,N_13124);
nand U23106 (N_23106,N_16476,N_15525);
nand U23107 (N_23107,N_14997,N_16327);
nor U23108 (N_23108,N_16780,N_13833);
nor U23109 (N_23109,N_12878,N_17708);
nor U23110 (N_23110,N_17613,N_17058);
and U23111 (N_23111,N_17412,N_14728);
and U23112 (N_23112,N_12979,N_18391);
xnor U23113 (N_23113,N_16036,N_17620);
or U23114 (N_23114,N_17723,N_14382);
nor U23115 (N_23115,N_17011,N_15068);
or U23116 (N_23116,N_18065,N_13113);
nor U23117 (N_23117,N_14324,N_13622);
and U23118 (N_23118,N_17276,N_17515);
nand U23119 (N_23119,N_14102,N_18289);
nor U23120 (N_23120,N_13411,N_14430);
xor U23121 (N_23121,N_12916,N_15748);
nor U23122 (N_23122,N_18119,N_18443);
or U23123 (N_23123,N_12715,N_15839);
and U23124 (N_23124,N_17562,N_12963);
or U23125 (N_23125,N_15702,N_18305);
nand U23126 (N_23126,N_13524,N_17128);
nor U23127 (N_23127,N_13006,N_18253);
and U23128 (N_23128,N_14205,N_14537);
or U23129 (N_23129,N_12567,N_14493);
xnor U23130 (N_23130,N_17851,N_16033);
nor U23131 (N_23131,N_14874,N_13560);
and U23132 (N_23132,N_14857,N_18684);
or U23133 (N_23133,N_14067,N_14032);
and U23134 (N_23134,N_13093,N_14056);
or U23135 (N_23135,N_13777,N_17033);
and U23136 (N_23136,N_14579,N_17338);
or U23137 (N_23137,N_17914,N_12701);
and U23138 (N_23138,N_16674,N_17103);
nor U23139 (N_23139,N_12864,N_17350);
nand U23140 (N_23140,N_18240,N_14859);
and U23141 (N_23141,N_15237,N_16186);
nand U23142 (N_23142,N_15739,N_16237);
and U23143 (N_23143,N_15201,N_15244);
xor U23144 (N_23144,N_14274,N_15557);
nor U23145 (N_23145,N_18431,N_14620);
xnor U23146 (N_23146,N_15327,N_16982);
or U23147 (N_23147,N_12881,N_18200);
nor U23148 (N_23148,N_17121,N_13348);
nand U23149 (N_23149,N_12939,N_17115);
nor U23150 (N_23150,N_14936,N_12673);
nor U23151 (N_23151,N_14350,N_12779);
or U23152 (N_23152,N_18600,N_17561);
nand U23153 (N_23153,N_17045,N_17396);
xor U23154 (N_23154,N_16118,N_13990);
or U23155 (N_23155,N_13767,N_13373);
xor U23156 (N_23156,N_14944,N_15824);
or U23157 (N_23157,N_18546,N_18198);
or U23158 (N_23158,N_16434,N_13006);
and U23159 (N_23159,N_15326,N_15588);
nand U23160 (N_23160,N_17511,N_18652);
nand U23161 (N_23161,N_17053,N_13020);
nor U23162 (N_23162,N_15684,N_16273);
nor U23163 (N_23163,N_13994,N_14505);
and U23164 (N_23164,N_15141,N_13682);
or U23165 (N_23165,N_17992,N_15212);
xor U23166 (N_23166,N_12502,N_12744);
nand U23167 (N_23167,N_15181,N_15841);
or U23168 (N_23168,N_18093,N_16771);
and U23169 (N_23169,N_13007,N_17089);
or U23170 (N_23170,N_17791,N_15744);
nor U23171 (N_23171,N_13170,N_12745);
nand U23172 (N_23172,N_15146,N_13888);
or U23173 (N_23173,N_14131,N_15800);
nor U23174 (N_23174,N_16459,N_14123);
or U23175 (N_23175,N_12914,N_17927);
nand U23176 (N_23176,N_15388,N_18479);
or U23177 (N_23177,N_15220,N_13746);
nand U23178 (N_23178,N_15636,N_16861);
and U23179 (N_23179,N_18249,N_12665);
or U23180 (N_23180,N_17799,N_16613);
or U23181 (N_23181,N_13301,N_14107);
nor U23182 (N_23182,N_13571,N_12819);
nor U23183 (N_23183,N_14749,N_14471);
or U23184 (N_23184,N_15250,N_15061);
or U23185 (N_23185,N_15411,N_15976);
xor U23186 (N_23186,N_17115,N_13696);
or U23187 (N_23187,N_18639,N_16398);
nor U23188 (N_23188,N_13350,N_17820);
or U23189 (N_23189,N_17916,N_17922);
and U23190 (N_23190,N_16562,N_12989);
or U23191 (N_23191,N_13924,N_14207);
nand U23192 (N_23192,N_17180,N_12879);
or U23193 (N_23193,N_13441,N_13752);
nor U23194 (N_23194,N_14158,N_13403);
xnor U23195 (N_23195,N_18625,N_14007);
and U23196 (N_23196,N_13959,N_16085);
nor U23197 (N_23197,N_15866,N_16847);
nand U23198 (N_23198,N_18541,N_13961);
xnor U23199 (N_23199,N_16378,N_16906);
nand U23200 (N_23200,N_12748,N_15854);
nand U23201 (N_23201,N_18735,N_16546);
xnor U23202 (N_23202,N_16253,N_14617);
nand U23203 (N_23203,N_15020,N_12525);
nor U23204 (N_23204,N_17708,N_17746);
nand U23205 (N_23205,N_17212,N_13129);
or U23206 (N_23206,N_14743,N_14347);
nor U23207 (N_23207,N_15818,N_13357);
nor U23208 (N_23208,N_15640,N_16294);
nor U23209 (N_23209,N_12819,N_18102);
nor U23210 (N_23210,N_16601,N_14977);
and U23211 (N_23211,N_13353,N_18286);
and U23212 (N_23212,N_18440,N_12986);
nor U23213 (N_23213,N_14401,N_18675);
nand U23214 (N_23214,N_17280,N_15083);
and U23215 (N_23215,N_12933,N_18051);
and U23216 (N_23216,N_14322,N_14683);
nand U23217 (N_23217,N_16365,N_15532);
and U23218 (N_23218,N_14347,N_15038);
and U23219 (N_23219,N_12842,N_14891);
nand U23220 (N_23220,N_13795,N_15733);
or U23221 (N_23221,N_12959,N_17137);
or U23222 (N_23222,N_15433,N_16031);
or U23223 (N_23223,N_14039,N_17890);
nand U23224 (N_23224,N_15968,N_14224);
nand U23225 (N_23225,N_14290,N_18564);
nand U23226 (N_23226,N_12674,N_18309);
nand U23227 (N_23227,N_14389,N_17991);
or U23228 (N_23228,N_15296,N_16701);
xor U23229 (N_23229,N_18374,N_17946);
nor U23230 (N_23230,N_16341,N_17637);
and U23231 (N_23231,N_15323,N_18549);
nor U23232 (N_23232,N_14055,N_17576);
or U23233 (N_23233,N_15295,N_13257);
and U23234 (N_23234,N_14144,N_15464);
xor U23235 (N_23235,N_17672,N_15667);
nand U23236 (N_23236,N_15904,N_16566);
nor U23237 (N_23237,N_14936,N_18197);
xor U23238 (N_23238,N_15743,N_14560);
nor U23239 (N_23239,N_13694,N_16026);
nor U23240 (N_23240,N_15520,N_17253);
or U23241 (N_23241,N_16463,N_15915);
and U23242 (N_23242,N_13244,N_17043);
and U23243 (N_23243,N_12522,N_14269);
and U23244 (N_23244,N_16499,N_16006);
nand U23245 (N_23245,N_15953,N_17862);
nor U23246 (N_23246,N_13863,N_13952);
or U23247 (N_23247,N_14836,N_14069);
or U23248 (N_23248,N_13774,N_17772);
and U23249 (N_23249,N_13530,N_18740);
and U23250 (N_23250,N_16875,N_13113);
nor U23251 (N_23251,N_18074,N_16768);
nor U23252 (N_23252,N_12737,N_16015);
and U23253 (N_23253,N_16535,N_17619);
nand U23254 (N_23254,N_17939,N_13892);
nand U23255 (N_23255,N_16432,N_17051);
and U23256 (N_23256,N_12977,N_18549);
xor U23257 (N_23257,N_15556,N_15991);
and U23258 (N_23258,N_13978,N_16022);
nand U23259 (N_23259,N_15597,N_16825);
and U23260 (N_23260,N_17115,N_18366);
and U23261 (N_23261,N_17490,N_15308);
or U23262 (N_23262,N_17751,N_16248);
nand U23263 (N_23263,N_17998,N_15061);
nand U23264 (N_23264,N_14745,N_13004);
nor U23265 (N_23265,N_17308,N_16220);
nor U23266 (N_23266,N_14624,N_13385);
or U23267 (N_23267,N_14890,N_13356);
or U23268 (N_23268,N_14443,N_16593);
nand U23269 (N_23269,N_17463,N_13098);
nor U23270 (N_23270,N_16323,N_13699);
nand U23271 (N_23271,N_13767,N_12931);
and U23272 (N_23272,N_17907,N_17623);
nor U23273 (N_23273,N_15141,N_16192);
or U23274 (N_23274,N_14670,N_14843);
or U23275 (N_23275,N_12786,N_13356);
xor U23276 (N_23276,N_15818,N_17053);
or U23277 (N_23277,N_12784,N_15004);
nand U23278 (N_23278,N_16780,N_12928);
and U23279 (N_23279,N_14675,N_16868);
nor U23280 (N_23280,N_15068,N_13315);
nand U23281 (N_23281,N_18505,N_16855);
or U23282 (N_23282,N_14670,N_17301);
and U23283 (N_23283,N_17182,N_14369);
nand U23284 (N_23284,N_18133,N_13561);
nor U23285 (N_23285,N_16824,N_17643);
or U23286 (N_23286,N_14006,N_15489);
or U23287 (N_23287,N_16826,N_13817);
or U23288 (N_23288,N_18739,N_15873);
or U23289 (N_23289,N_14669,N_14541);
nand U23290 (N_23290,N_18141,N_13470);
nor U23291 (N_23291,N_14353,N_17074);
xnor U23292 (N_23292,N_16004,N_14413);
and U23293 (N_23293,N_17281,N_17733);
and U23294 (N_23294,N_17037,N_14834);
xor U23295 (N_23295,N_18565,N_18366);
xnor U23296 (N_23296,N_14642,N_15571);
and U23297 (N_23297,N_17468,N_15120);
nand U23298 (N_23298,N_12933,N_13091);
and U23299 (N_23299,N_18170,N_13702);
nor U23300 (N_23300,N_14424,N_18630);
and U23301 (N_23301,N_15086,N_16036);
or U23302 (N_23302,N_15269,N_15967);
nand U23303 (N_23303,N_13886,N_15147);
nand U23304 (N_23304,N_12941,N_18399);
nand U23305 (N_23305,N_14665,N_13437);
nand U23306 (N_23306,N_16552,N_13457);
or U23307 (N_23307,N_13459,N_16526);
and U23308 (N_23308,N_15078,N_15069);
and U23309 (N_23309,N_16344,N_15435);
xnor U23310 (N_23310,N_17659,N_13938);
xnor U23311 (N_23311,N_18168,N_14029);
nand U23312 (N_23312,N_15202,N_15957);
nor U23313 (N_23313,N_18742,N_13177);
nor U23314 (N_23314,N_16211,N_18515);
and U23315 (N_23315,N_15938,N_13610);
nand U23316 (N_23316,N_14624,N_16352);
and U23317 (N_23317,N_18438,N_17632);
or U23318 (N_23318,N_13280,N_18030);
and U23319 (N_23319,N_15228,N_13569);
xnor U23320 (N_23320,N_14489,N_13673);
and U23321 (N_23321,N_17786,N_15697);
or U23322 (N_23322,N_14820,N_15723);
xor U23323 (N_23323,N_14928,N_15751);
nand U23324 (N_23324,N_17393,N_12593);
nor U23325 (N_23325,N_18397,N_14852);
nand U23326 (N_23326,N_15655,N_17431);
or U23327 (N_23327,N_18505,N_15207);
or U23328 (N_23328,N_16614,N_13586);
or U23329 (N_23329,N_15703,N_13614);
and U23330 (N_23330,N_13362,N_12794);
nand U23331 (N_23331,N_17489,N_17495);
and U23332 (N_23332,N_14322,N_12576);
or U23333 (N_23333,N_13273,N_13682);
or U23334 (N_23334,N_18496,N_15898);
nand U23335 (N_23335,N_12631,N_14019);
xnor U23336 (N_23336,N_18040,N_15272);
nor U23337 (N_23337,N_14370,N_17536);
nor U23338 (N_23338,N_17262,N_12934);
nand U23339 (N_23339,N_16538,N_15432);
or U23340 (N_23340,N_12685,N_14522);
nand U23341 (N_23341,N_17483,N_18408);
nor U23342 (N_23342,N_17087,N_15672);
and U23343 (N_23343,N_14209,N_16821);
and U23344 (N_23344,N_14549,N_17696);
or U23345 (N_23345,N_14738,N_17927);
nand U23346 (N_23346,N_17993,N_17174);
nand U23347 (N_23347,N_16309,N_15825);
and U23348 (N_23348,N_17624,N_18292);
xor U23349 (N_23349,N_15486,N_14985);
and U23350 (N_23350,N_14667,N_12624);
and U23351 (N_23351,N_14132,N_14601);
nor U23352 (N_23352,N_13932,N_16299);
and U23353 (N_23353,N_14116,N_18743);
and U23354 (N_23354,N_16147,N_17667);
xnor U23355 (N_23355,N_13159,N_14774);
or U23356 (N_23356,N_17184,N_15037);
nor U23357 (N_23357,N_17502,N_18228);
nor U23358 (N_23358,N_14537,N_17847);
nor U23359 (N_23359,N_14990,N_16191);
nor U23360 (N_23360,N_14379,N_15667);
xor U23361 (N_23361,N_14890,N_16899);
and U23362 (N_23362,N_17750,N_16436);
xor U23363 (N_23363,N_15582,N_13156);
or U23364 (N_23364,N_15535,N_16154);
nor U23365 (N_23365,N_18493,N_13986);
nor U23366 (N_23366,N_15153,N_16025);
nand U23367 (N_23367,N_14246,N_14443);
and U23368 (N_23368,N_16755,N_13966);
or U23369 (N_23369,N_15169,N_13436);
or U23370 (N_23370,N_12607,N_16643);
nor U23371 (N_23371,N_15132,N_17288);
or U23372 (N_23372,N_16320,N_17410);
and U23373 (N_23373,N_14129,N_14495);
xor U23374 (N_23374,N_16925,N_13063);
or U23375 (N_23375,N_13352,N_16734);
or U23376 (N_23376,N_16116,N_18042);
nand U23377 (N_23377,N_18656,N_18164);
or U23378 (N_23378,N_16535,N_17738);
or U23379 (N_23379,N_16700,N_14458);
and U23380 (N_23380,N_17303,N_12685);
nand U23381 (N_23381,N_18194,N_17214);
nand U23382 (N_23382,N_14607,N_13681);
or U23383 (N_23383,N_15207,N_15123);
nand U23384 (N_23384,N_18599,N_14088);
and U23385 (N_23385,N_14225,N_16878);
nand U23386 (N_23386,N_13756,N_13425);
nand U23387 (N_23387,N_16691,N_18300);
nand U23388 (N_23388,N_15220,N_18365);
and U23389 (N_23389,N_17701,N_13378);
nor U23390 (N_23390,N_15264,N_17598);
nand U23391 (N_23391,N_17396,N_14936);
nor U23392 (N_23392,N_14817,N_14121);
and U23393 (N_23393,N_18113,N_15063);
or U23394 (N_23394,N_17414,N_14753);
nor U23395 (N_23395,N_15667,N_13387);
and U23396 (N_23396,N_13045,N_14097);
or U23397 (N_23397,N_14049,N_18420);
or U23398 (N_23398,N_18192,N_15467);
or U23399 (N_23399,N_16828,N_18013);
nor U23400 (N_23400,N_16978,N_14361);
or U23401 (N_23401,N_12875,N_17316);
nand U23402 (N_23402,N_17796,N_14298);
and U23403 (N_23403,N_13970,N_16958);
and U23404 (N_23404,N_12785,N_15903);
or U23405 (N_23405,N_12675,N_18315);
or U23406 (N_23406,N_15926,N_14756);
xor U23407 (N_23407,N_18318,N_14971);
xor U23408 (N_23408,N_17494,N_12996);
nor U23409 (N_23409,N_16556,N_13807);
or U23410 (N_23410,N_17426,N_17593);
and U23411 (N_23411,N_17424,N_13995);
or U23412 (N_23412,N_17274,N_18631);
or U23413 (N_23413,N_13439,N_14020);
nor U23414 (N_23414,N_16847,N_18664);
nand U23415 (N_23415,N_17662,N_18221);
nand U23416 (N_23416,N_14699,N_17110);
nor U23417 (N_23417,N_13288,N_18094);
or U23418 (N_23418,N_15678,N_12927);
nor U23419 (N_23419,N_18152,N_16120);
xor U23420 (N_23420,N_17492,N_13333);
nand U23421 (N_23421,N_12635,N_18710);
nor U23422 (N_23422,N_16279,N_14567);
nand U23423 (N_23423,N_12558,N_13916);
and U23424 (N_23424,N_13615,N_15073);
or U23425 (N_23425,N_14679,N_17157);
nor U23426 (N_23426,N_15104,N_17700);
or U23427 (N_23427,N_13987,N_17636);
or U23428 (N_23428,N_13881,N_15071);
or U23429 (N_23429,N_12554,N_16375);
xor U23430 (N_23430,N_13801,N_16862);
nor U23431 (N_23431,N_12998,N_15079);
or U23432 (N_23432,N_16314,N_15862);
and U23433 (N_23433,N_18377,N_17576);
and U23434 (N_23434,N_16717,N_13405);
or U23435 (N_23435,N_12708,N_13652);
or U23436 (N_23436,N_13564,N_14762);
and U23437 (N_23437,N_15648,N_15900);
and U23438 (N_23438,N_13920,N_17469);
or U23439 (N_23439,N_13868,N_15520);
or U23440 (N_23440,N_12557,N_13512);
nor U23441 (N_23441,N_17816,N_16872);
nor U23442 (N_23442,N_15425,N_16535);
or U23443 (N_23443,N_16117,N_16401);
and U23444 (N_23444,N_16183,N_12836);
and U23445 (N_23445,N_14285,N_16472);
or U23446 (N_23446,N_15637,N_16895);
xnor U23447 (N_23447,N_14922,N_15912);
or U23448 (N_23448,N_17510,N_17532);
nor U23449 (N_23449,N_17471,N_16809);
or U23450 (N_23450,N_13849,N_15211);
or U23451 (N_23451,N_18035,N_17067);
and U23452 (N_23452,N_16457,N_13813);
nand U23453 (N_23453,N_16363,N_13910);
or U23454 (N_23454,N_14101,N_12837);
nor U23455 (N_23455,N_13114,N_12547);
and U23456 (N_23456,N_15539,N_18562);
and U23457 (N_23457,N_13158,N_14099);
xnor U23458 (N_23458,N_13462,N_13529);
nand U23459 (N_23459,N_15969,N_13235);
nand U23460 (N_23460,N_14214,N_17459);
or U23461 (N_23461,N_13598,N_16152);
or U23462 (N_23462,N_17246,N_16184);
nor U23463 (N_23463,N_15937,N_15463);
or U23464 (N_23464,N_16361,N_18439);
nand U23465 (N_23465,N_12538,N_15857);
nand U23466 (N_23466,N_14374,N_16114);
xnor U23467 (N_23467,N_16512,N_13844);
nor U23468 (N_23468,N_16697,N_17657);
nand U23469 (N_23469,N_14431,N_17599);
or U23470 (N_23470,N_15102,N_17897);
nand U23471 (N_23471,N_14935,N_14798);
and U23472 (N_23472,N_13592,N_14719);
and U23473 (N_23473,N_13814,N_18493);
or U23474 (N_23474,N_15522,N_12950);
and U23475 (N_23475,N_13224,N_18011);
and U23476 (N_23476,N_14475,N_15606);
nand U23477 (N_23477,N_12792,N_16797);
nand U23478 (N_23478,N_14594,N_15644);
or U23479 (N_23479,N_13142,N_16488);
nor U23480 (N_23480,N_12747,N_15030);
nand U23481 (N_23481,N_15580,N_14290);
nor U23482 (N_23482,N_14775,N_18040);
and U23483 (N_23483,N_16564,N_16741);
nor U23484 (N_23484,N_14016,N_17559);
nor U23485 (N_23485,N_14274,N_12694);
and U23486 (N_23486,N_18498,N_16659);
or U23487 (N_23487,N_17417,N_16917);
nand U23488 (N_23488,N_13625,N_12914);
nand U23489 (N_23489,N_15635,N_13193);
or U23490 (N_23490,N_17841,N_12801);
and U23491 (N_23491,N_16450,N_13462);
and U23492 (N_23492,N_12986,N_14619);
nor U23493 (N_23493,N_18326,N_16627);
and U23494 (N_23494,N_17886,N_17081);
nand U23495 (N_23495,N_12517,N_16310);
and U23496 (N_23496,N_12861,N_15096);
and U23497 (N_23497,N_14185,N_14183);
xnor U23498 (N_23498,N_13370,N_14825);
nor U23499 (N_23499,N_18240,N_15999);
nand U23500 (N_23500,N_14582,N_13896);
nand U23501 (N_23501,N_18451,N_16049);
nand U23502 (N_23502,N_14707,N_16766);
nor U23503 (N_23503,N_15327,N_16410);
and U23504 (N_23504,N_16343,N_13714);
nor U23505 (N_23505,N_15380,N_17257);
nand U23506 (N_23506,N_15112,N_12756);
or U23507 (N_23507,N_18359,N_17307);
xor U23508 (N_23508,N_17667,N_13017);
or U23509 (N_23509,N_16562,N_12595);
nand U23510 (N_23510,N_13160,N_15293);
nand U23511 (N_23511,N_16888,N_17766);
or U23512 (N_23512,N_15074,N_13637);
nor U23513 (N_23513,N_13222,N_13425);
nand U23514 (N_23514,N_17434,N_12756);
or U23515 (N_23515,N_14055,N_14659);
xnor U23516 (N_23516,N_15223,N_13858);
xnor U23517 (N_23517,N_16663,N_13637);
or U23518 (N_23518,N_15973,N_17403);
nand U23519 (N_23519,N_16266,N_18420);
and U23520 (N_23520,N_12696,N_13545);
nor U23521 (N_23521,N_13873,N_17315);
nor U23522 (N_23522,N_13146,N_13623);
nand U23523 (N_23523,N_16217,N_18366);
xor U23524 (N_23524,N_15553,N_12880);
xor U23525 (N_23525,N_14179,N_16421);
nor U23526 (N_23526,N_18566,N_17560);
or U23527 (N_23527,N_18463,N_18628);
and U23528 (N_23528,N_17013,N_16389);
nor U23529 (N_23529,N_13796,N_18055);
nor U23530 (N_23530,N_13175,N_17791);
or U23531 (N_23531,N_14486,N_13410);
nand U23532 (N_23532,N_16777,N_15350);
or U23533 (N_23533,N_18273,N_12996);
or U23534 (N_23534,N_12794,N_15703);
and U23535 (N_23535,N_15544,N_18289);
and U23536 (N_23536,N_12800,N_18200);
and U23537 (N_23537,N_14456,N_17158);
nand U23538 (N_23538,N_13718,N_18732);
nor U23539 (N_23539,N_18426,N_17134);
and U23540 (N_23540,N_13634,N_12649);
nor U23541 (N_23541,N_16418,N_12832);
or U23542 (N_23542,N_13533,N_16914);
or U23543 (N_23543,N_12923,N_16559);
and U23544 (N_23544,N_15870,N_12914);
nand U23545 (N_23545,N_17992,N_17912);
and U23546 (N_23546,N_12866,N_16230);
nor U23547 (N_23547,N_18749,N_16079);
xnor U23548 (N_23548,N_14061,N_13103);
nor U23549 (N_23549,N_16278,N_17279);
nor U23550 (N_23550,N_18416,N_13493);
and U23551 (N_23551,N_16379,N_18007);
and U23552 (N_23552,N_14715,N_14322);
xnor U23553 (N_23553,N_12700,N_12689);
or U23554 (N_23554,N_17338,N_16441);
nand U23555 (N_23555,N_17060,N_12991);
or U23556 (N_23556,N_18303,N_14422);
xnor U23557 (N_23557,N_17832,N_14182);
nor U23558 (N_23558,N_18375,N_16626);
nand U23559 (N_23559,N_16118,N_16320);
and U23560 (N_23560,N_14452,N_18021);
and U23561 (N_23561,N_17374,N_13870);
nand U23562 (N_23562,N_13896,N_13543);
nand U23563 (N_23563,N_13069,N_15902);
and U23564 (N_23564,N_13739,N_17803);
and U23565 (N_23565,N_17879,N_14007);
nand U23566 (N_23566,N_16777,N_17980);
and U23567 (N_23567,N_15350,N_18160);
nand U23568 (N_23568,N_13302,N_18727);
xnor U23569 (N_23569,N_17950,N_17426);
or U23570 (N_23570,N_13111,N_17805);
or U23571 (N_23571,N_13919,N_18176);
or U23572 (N_23572,N_15123,N_16461);
xnor U23573 (N_23573,N_18473,N_16724);
xnor U23574 (N_23574,N_13614,N_16806);
nand U23575 (N_23575,N_13604,N_12677);
and U23576 (N_23576,N_14639,N_13021);
nand U23577 (N_23577,N_14062,N_13657);
nor U23578 (N_23578,N_13935,N_18027);
or U23579 (N_23579,N_12872,N_18231);
and U23580 (N_23580,N_14919,N_13793);
nand U23581 (N_23581,N_14180,N_17055);
or U23582 (N_23582,N_18419,N_17933);
or U23583 (N_23583,N_13067,N_18442);
and U23584 (N_23584,N_14404,N_18728);
and U23585 (N_23585,N_16890,N_14106);
nand U23586 (N_23586,N_18179,N_17411);
nand U23587 (N_23587,N_17828,N_16151);
or U23588 (N_23588,N_16741,N_13689);
or U23589 (N_23589,N_13253,N_17386);
nand U23590 (N_23590,N_18693,N_17101);
nor U23591 (N_23591,N_14832,N_16958);
or U23592 (N_23592,N_15731,N_12703);
or U23593 (N_23593,N_14370,N_13980);
or U23594 (N_23594,N_18587,N_13561);
nand U23595 (N_23595,N_17034,N_16200);
or U23596 (N_23596,N_16761,N_15062);
xor U23597 (N_23597,N_14826,N_17849);
and U23598 (N_23598,N_17408,N_17136);
nand U23599 (N_23599,N_18127,N_15172);
and U23600 (N_23600,N_15698,N_14946);
and U23601 (N_23601,N_13784,N_14341);
nand U23602 (N_23602,N_12871,N_17700);
or U23603 (N_23603,N_14524,N_18495);
xnor U23604 (N_23604,N_16904,N_16330);
nor U23605 (N_23605,N_14099,N_17466);
or U23606 (N_23606,N_18204,N_14215);
or U23607 (N_23607,N_14587,N_14755);
nand U23608 (N_23608,N_17261,N_13815);
nor U23609 (N_23609,N_13114,N_14592);
or U23610 (N_23610,N_18094,N_14798);
or U23611 (N_23611,N_15756,N_16365);
nand U23612 (N_23612,N_17664,N_18494);
nor U23613 (N_23613,N_14691,N_14174);
nand U23614 (N_23614,N_15693,N_16823);
and U23615 (N_23615,N_14523,N_17166);
and U23616 (N_23616,N_16329,N_15070);
xnor U23617 (N_23617,N_14974,N_14593);
or U23618 (N_23618,N_17647,N_16603);
nand U23619 (N_23619,N_14333,N_17809);
nor U23620 (N_23620,N_17297,N_17765);
or U23621 (N_23621,N_16257,N_12538);
xor U23622 (N_23622,N_14754,N_17530);
nand U23623 (N_23623,N_13374,N_16673);
nor U23624 (N_23624,N_16806,N_13110);
or U23625 (N_23625,N_13475,N_13491);
nor U23626 (N_23626,N_14912,N_13784);
or U23627 (N_23627,N_13928,N_17711);
nand U23628 (N_23628,N_13952,N_14746);
or U23629 (N_23629,N_14185,N_15519);
nor U23630 (N_23630,N_15439,N_15754);
and U23631 (N_23631,N_14568,N_17417);
and U23632 (N_23632,N_12971,N_13787);
nand U23633 (N_23633,N_14886,N_15355);
nand U23634 (N_23634,N_18294,N_14665);
nor U23635 (N_23635,N_14547,N_12861);
nor U23636 (N_23636,N_14114,N_18048);
xor U23637 (N_23637,N_18640,N_17310);
nor U23638 (N_23638,N_13679,N_13891);
and U23639 (N_23639,N_16793,N_17176);
or U23640 (N_23640,N_12733,N_14972);
or U23641 (N_23641,N_13348,N_12764);
or U23642 (N_23642,N_14041,N_16929);
nand U23643 (N_23643,N_15053,N_16103);
and U23644 (N_23644,N_13543,N_16992);
nor U23645 (N_23645,N_18407,N_12747);
nand U23646 (N_23646,N_18261,N_12933);
and U23647 (N_23647,N_16120,N_18529);
and U23648 (N_23648,N_17779,N_16359);
or U23649 (N_23649,N_16536,N_12748);
and U23650 (N_23650,N_13539,N_18553);
or U23651 (N_23651,N_15937,N_15324);
xor U23652 (N_23652,N_17360,N_16686);
xor U23653 (N_23653,N_18234,N_17389);
nand U23654 (N_23654,N_13525,N_18540);
xnor U23655 (N_23655,N_14641,N_17312);
nand U23656 (N_23656,N_15237,N_14085);
or U23657 (N_23657,N_15420,N_17897);
nor U23658 (N_23658,N_13440,N_14470);
nor U23659 (N_23659,N_15223,N_12627);
xnor U23660 (N_23660,N_13140,N_13914);
nor U23661 (N_23661,N_13011,N_15224);
nand U23662 (N_23662,N_17006,N_15884);
nor U23663 (N_23663,N_16274,N_15041);
xor U23664 (N_23664,N_18394,N_14035);
or U23665 (N_23665,N_14069,N_16551);
nor U23666 (N_23666,N_15913,N_14071);
or U23667 (N_23667,N_18628,N_15096);
nor U23668 (N_23668,N_14351,N_13741);
nor U23669 (N_23669,N_17675,N_15350);
nor U23670 (N_23670,N_16369,N_16561);
nor U23671 (N_23671,N_17098,N_15714);
nand U23672 (N_23672,N_16221,N_16462);
or U23673 (N_23673,N_17470,N_15864);
or U23674 (N_23674,N_18582,N_16309);
nor U23675 (N_23675,N_14654,N_17265);
nand U23676 (N_23676,N_17770,N_13906);
nor U23677 (N_23677,N_12956,N_16665);
nand U23678 (N_23678,N_13312,N_14948);
xor U23679 (N_23679,N_18168,N_17018);
and U23680 (N_23680,N_15840,N_16188);
and U23681 (N_23681,N_13065,N_17945);
xor U23682 (N_23682,N_16281,N_17196);
nor U23683 (N_23683,N_13611,N_13636);
or U23684 (N_23684,N_18029,N_13375);
nand U23685 (N_23685,N_16973,N_14668);
and U23686 (N_23686,N_18675,N_17381);
xor U23687 (N_23687,N_17323,N_14292);
or U23688 (N_23688,N_13286,N_17166);
nor U23689 (N_23689,N_15049,N_16566);
nand U23690 (N_23690,N_13244,N_17311);
xor U23691 (N_23691,N_16589,N_13457);
nand U23692 (N_23692,N_15024,N_15451);
or U23693 (N_23693,N_17053,N_13743);
or U23694 (N_23694,N_15665,N_15327);
and U23695 (N_23695,N_16942,N_13360);
nor U23696 (N_23696,N_15173,N_12807);
xor U23697 (N_23697,N_18167,N_12717);
or U23698 (N_23698,N_14483,N_12952);
and U23699 (N_23699,N_12959,N_16111);
or U23700 (N_23700,N_13527,N_16406);
xnor U23701 (N_23701,N_16835,N_16549);
nor U23702 (N_23702,N_13629,N_12829);
and U23703 (N_23703,N_17892,N_17962);
nand U23704 (N_23704,N_14275,N_17399);
nand U23705 (N_23705,N_15926,N_18597);
nor U23706 (N_23706,N_14994,N_14130);
and U23707 (N_23707,N_16049,N_17666);
xnor U23708 (N_23708,N_14031,N_13254);
nand U23709 (N_23709,N_18337,N_16987);
nor U23710 (N_23710,N_14032,N_16325);
nand U23711 (N_23711,N_15137,N_14908);
nor U23712 (N_23712,N_16484,N_15278);
nor U23713 (N_23713,N_13005,N_12819);
or U23714 (N_23714,N_14420,N_13406);
nor U23715 (N_23715,N_16865,N_13327);
nand U23716 (N_23716,N_13041,N_14593);
and U23717 (N_23717,N_14723,N_13658);
or U23718 (N_23718,N_17754,N_18333);
nor U23719 (N_23719,N_17261,N_12919);
or U23720 (N_23720,N_13734,N_16764);
or U23721 (N_23721,N_14436,N_14637);
or U23722 (N_23722,N_17296,N_17373);
nand U23723 (N_23723,N_16981,N_16374);
or U23724 (N_23724,N_17609,N_17595);
and U23725 (N_23725,N_14652,N_13269);
and U23726 (N_23726,N_13626,N_12713);
or U23727 (N_23727,N_16995,N_14637);
xor U23728 (N_23728,N_18285,N_18634);
and U23729 (N_23729,N_16237,N_15499);
nand U23730 (N_23730,N_15794,N_14924);
nand U23731 (N_23731,N_14902,N_15399);
xor U23732 (N_23732,N_18486,N_14231);
nor U23733 (N_23733,N_15797,N_15408);
nand U23734 (N_23734,N_14705,N_15885);
nand U23735 (N_23735,N_14065,N_16833);
nor U23736 (N_23736,N_15578,N_16106);
and U23737 (N_23737,N_17902,N_17023);
and U23738 (N_23738,N_16228,N_18281);
or U23739 (N_23739,N_16011,N_15753);
xnor U23740 (N_23740,N_17629,N_13510);
or U23741 (N_23741,N_17832,N_14617);
and U23742 (N_23742,N_16064,N_17234);
or U23743 (N_23743,N_16166,N_13329);
or U23744 (N_23744,N_15617,N_13444);
or U23745 (N_23745,N_14855,N_15150);
and U23746 (N_23746,N_17509,N_14497);
nand U23747 (N_23747,N_13906,N_15897);
and U23748 (N_23748,N_14068,N_17893);
nor U23749 (N_23749,N_14103,N_16677);
or U23750 (N_23750,N_14609,N_12734);
or U23751 (N_23751,N_14904,N_17972);
nand U23752 (N_23752,N_18624,N_14000);
nor U23753 (N_23753,N_13056,N_15119);
and U23754 (N_23754,N_13541,N_17842);
or U23755 (N_23755,N_15726,N_17160);
xnor U23756 (N_23756,N_14455,N_13725);
nand U23757 (N_23757,N_15533,N_17903);
and U23758 (N_23758,N_12687,N_16843);
and U23759 (N_23759,N_16232,N_16834);
or U23760 (N_23760,N_13803,N_13345);
and U23761 (N_23761,N_15837,N_13244);
nor U23762 (N_23762,N_13559,N_14893);
and U23763 (N_23763,N_13039,N_15594);
nand U23764 (N_23764,N_15028,N_17592);
and U23765 (N_23765,N_13814,N_18139);
and U23766 (N_23766,N_14176,N_12504);
or U23767 (N_23767,N_17281,N_16976);
nand U23768 (N_23768,N_16902,N_16642);
nor U23769 (N_23769,N_16504,N_17308);
and U23770 (N_23770,N_14903,N_13859);
nor U23771 (N_23771,N_14087,N_14526);
or U23772 (N_23772,N_15144,N_18168);
nand U23773 (N_23773,N_14399,N_13018);
nor U23774 (N_23774,N_16721,N_15443);
and U23775 (N_23775,N_16097,N_16114);
or U23776 (N_23776,N_13343,N_16086);
nor U23777 (N_23777,N_16931,N_12605);
and U23778 (N_23778,N_17339,N_15909);
xor U23779 (N_23779,N_14587,N_16550);
nand U23780 (N_23780,N_13927,N_13144);
nand U23781 (N_23781,N_17073,N_13243);
and U23782 (N_23782,N_15197,N_13407);
nor U23783 (N_23783,N_17965,N_18077);
nand U23784 (N_23784,N_14539,N_18370);
or U23785 (N_23785,N_16060,N_12792);
nor U23786 (N_23786,N_12650,N_14427);
nand U23787 (N_23787,N_15595,N_13796);
and U23788 (N_23788,N_13219,N_16688);
and U23789 (N_23789,N_13607,N_13232);
nand U23790 (N_23790,N_18618,N_14350);
and U23791 (N_23791,N_14628,N_13988);
or U23792 (N_23792,N_14504,N_16768);
and U23793 (N_23793,N_14374,N_15257);
nand U23794 (N_23794,N_17144,N_16170);
or U23795 (N_23795,N_13940,N_14133);
nor U23796 (N_23796,N_15009,N_16179);
nor U23797 (N_23797,N_14131,N_12671);
nand U23798 (N_23798,N_15825,N_18053);
and U23799 (N_23799,N_15701,N_13941);
or U23800 (N_23800,N_13244,N_18709);
or U23801 (N_23801,N_15122,N_17151);
nand U23802 (N_23802,N_12584,N_13659);
nand U23803 (N_23803,N_15671,N_18511);
xnor U23804 (N_23804,N_16818,N_15493);
and U23805 (N_23805,N_16873,N_16071);
or U23806 (N_23806,N_13310,N_16448);
nand U23807 (N_23807,N_18635,N_15617);
and U23808 (N_23808,N_14759,N_18655);
nand U23809 (N_23809,N_16274,N_18069);
nand U23810 (N_23810,N_16796,N_12992);
or U23811 (N_23811,N_15410,N_15910);
nor U23812 (N_23812,N_17154,N_16705);
or U23813 (N_23813,N_15323,N_18296);
nand U23814 (N_23814,N_18286,N_17999);
or U23815 (N_23815,N_16154,N_13193);
or U23816 (N_23816,N_16342,N_12606);
nor U23817 (N_23817,N_14445,N_13276);
or U23818 (N_23818,N_15846,N_17832);
nor U23819 (N_23819,N_18176,N_13137);
xor U23820 (N_23820,N_16649,N_18289);
nand U23821 (N_23821,N_16456,N_14933);
nand U23822 (N_23822,N_14524,N_14655);
and U23823 (N_23823,N_13413,N_17051);
and U23824 (N_23824,N_15067,N_13283);
and U23825 (N_23825,N_15558,N_15785);
nand U23826 (N_23826,N_13712,N_16573);
nand U23827 (N_23827,N_13219,N_14993);
or U23828 (N_23828,N_14286,N_17069);
nand U23829 (N_23829,N_15776,N_18546);
and U23830 (N_23830,N_15467,N_14300);
or U23831 (N_23831,N_17213,N_14999);
and U23832 (N_23832,N_14414,N_16940);
and U23833 (N_23833,N_13256,N_17058);
or U23834 (N_23834,N_14294,N_13142);
xnor U23835 (N_23835,N_14558,N_17677);
or U23836 (N_23836,N_15724,N_18716);
nand U23837 (N_23837,N_12651,N_18446);
or U23838 (N_23838,N_15907,N_12868);
nor U23839 (N_23839,N_13761,N_12621);
or U23840 (N_23840,N_14195,N_17628);
nand U23841 (N_23841,N_13574,N_13440);
and U23842 (N_23842,N_14937,N_15069);
nand U23843 (N_23843,N_13787,N_14810);
and U23844 (N_23844,N_18114,N_12869);
or U23845 (N_23845,N_16544,N_17070);
nor U23846 (N_23846,N_14816,N_16922);
and U23847 (N_23847,N_13241,N_13464);
nand U23848 (N_23848,N_16095,N_13944);
or U23849 (N_23849,N_15227,N_14815);
or U23850 (N_23850,N_14276,N_17933);
nor U23851 (N_23851,N_16216,N_12505);
nand U23852 (N_23852,N_15702,N_15120);
and U23853 (N_23853,N_12730,N_14867);
nor U23854 (N_23854,N_14926,N_17073);
nor U23855 (N_23855,N_17171,N_15676);
or U23856 (N_23856,N_17753,N_14720);
or U23857 (N_23857,N_12850,N_16104);
xnor U23858 (N_23858,N_14735,N_13070);
xnor U23859 (N_23859,N_15674,N_12755);
nor U23860 (N_23860,N_16942,N_14078);
and U23861 (N_23861,N_12853,N_16725);
nand U23862 (N_23862,N_16373,N_12838);
xnor U23863 (N_23863,N_13443,N_17226);
or U23864 (N_23864,N_17001,N_15037);
nor U23865 (N_23865,N_14666,N_18032);
and U23866 (N_23866,N_14486,N_15411);
nor U23867 (N_23867,N_16523,N_17507);
nor U23868 (N_23868,N_17711,N_18684);
and U23869 (N_23869,N_17832,N_13908);
nor U23870 (N_23870,N_16997,N_15360);
nor U23871 (N_23871,N_15824,N_16198);
nor U23872 (N_23872,N_14968,N_14974);
nor U23873 (N_23873,N_13230,N_18488);
nand U23874 (N_23874,N_15257,N_12980);
or U23875 (N_23875,N_13945,N_15374);
nor U23876 (N_23876,N_14465,N_15657);
nand U23877 (N_23877,N_18161,N_15163);
nand U23878 (N_23878,N_14413,N_15948);
or U23879 (N_23879,N_18421,N_14962);
nor U23880 (N_23880,N_12901,N_12981);
or U23881 (N_23881,N_14005,N_16592);
xor U23882 (N_23882,N_14201,N_13513);
or U23883 (N_23883,N_13135,N_17908);
and U23884 (N_23884,N_18732,N_14539);
xor U23885 (N_23885,N_12722,N_18310);
or U23886 (N_23886,N_16052,N_15906);
nand U23887 (N_23887,N_12815,N_15737);
or U23888 (N_23888,N_18674,N_15187);
and U23889 (N_23889,N_13235,N_14588);
nand U23890 (N_23890,N_15506,N_13679);
xnor U23891 (N_23891,N_15805,N_13955);
nor U23892 (N_23892,N_13775,N_18268);
and U23893 (N_23893,N_16267,N_12710);
or U23894 (N_23894,N_14758,N_16106);
xnor U23895 (N_23895,N_13495,N_17062);
and U23896 (N_23896,N_14355,N_18542);
nor U23897 (N_23897,N_12881,N_15107);
nand U23898 (N_23898,N_17218,N_15248);
and U23899 (N_23899,N_18388,N_13329);
and U23900 (N_23900,N_17959,N_16582);
nand U23901 (N_23901,N_15120,N_14803);
and U23902 (N_23902,N_17427,N_13552);
nor U23903 (N_23903,N_13653,N_18185);
xor U23904 (N_23904,N_16339,N_18194);
nand U23905 (N_23905,N_17456,N_17390);
nand U23906 (N_23906,N_17785,N_14974);
nor U23907 (N_23907,N_13386,N_13862);
nor U23908 (N_23908,N_17991,N_14785);
xor U23909 (N_23909,N_17413,N_16058);
nor U23910 (N_23910,N_14953,N_13192);
or U23911 (N_23911,N_16016,N_16036);
xnor U23912 (N_23912,N_15032,N_16972);
nor U23913 (N_23913,N_18155,N_17026);
nor U23914 (N_23914,N_16486,N_14889);
or U23915 (N_23915,N_17882,N_18312);
and U23916 (N_23916,N_12787,N_14055);
xnor U23917 (N_23917,N_13942,N_15037);
nor U23918 (N_23918,N_17162,N_18358);
and U23919 (N_23919,N_17501,N_15461);
nand U23920 (N_23920,N_14727,N_18009);
or U23921 (N_23921,N_13463,N_17064);
and U23922 (N_23922,N_13915,N_14636);
xor U23923 (N_23923,N_14792,N_15143);
and U23924 (N_23924,N_16341,N_13822);
or U23925 (N_23925,N_16644,N_12662);
and U23926 (N_23926,N_18023,N_17263);
nand U23927 (N_23927,N_16462,N_17311);
or U23928 (N_23928,N_17173,N_15827);
nand U23929 (N_23929,N_17888,N_15470);
nor U23930 (N_23930,N_16976,N_15453);
nand U23931 (N_23931,N_14780,N_16579);
nand U23932 (N_23932,N_12939,N_16031);
and U23933 (N_23933,N_17005,N_15269);
nor U23934 (N_23934,N_15216,N_18159);
and U23935 (N_23935,N_12910,N_16003);
or U23936 (N_23936,N_16042,N_15299);
nor U23937 (N_23937,N_18406,N_13176);
nor U23938 (N_23938,N_14002,N_18275);
and U23939 (N_23939,N_15359,N_14358);
xnor U23940 (N_23940,N_18112,N_13252);
or U23941 (N_23941,N_13421,N_14807);
nand U23942 (N_23942,N_16961,N_17200);
nor U23943 (N_23943,N_14698,N_12654);
nor U23944 (N_23944,N_13918,N_13616);
and U23945 (N_23945,N_12870,N_17364);
and U23946 (N_23946,N_17082,N_17827);
nor U23947 (N_23947,N_14002,N_16144);
and U23948 (N_23948,N_17810,N_17123);
nor U23949 (N_23949,N_15491,N_18387);
or U23950 (N_23950,N_14166,N_15988);
or U23951 (N_23951,N_18681,N_15943);
or U23952 (N_23952,N_13521,N_16951);
or U23953 (N_23953,N_14541,N_13004);
nor U23954 (N_23954,N_14515,N_12755);
nand U23955 (N_23955,N_15586,N_17603);
or U23956 (N_23956,N_12597,N_16461);
nand U23957 (N_23957,N_17595,N_17927);
or U23958 (N_23958,N_13231,N_12579);
or U23959 (N_23959,N_14178,N_17576);
or U23960 (N_23960,N_14640,N_17699);
or U23961 (N_23961,N_16025,N_17187);
nor U23962 (N_23962,N_13068,N_13816);
or U23963 (N_23963,N_13857,N_14233);
or U23964 (N_23964,N_15081,N_14749);
and U23965 (N_23965,N_13612,N_12611);
nand U23966 (N_23966,N_14409,N_15933);
and U23967 (N_23967,N_18323,N_15380);
nor U23968 (N_23968,N_18697,N_16844);
xor U23969 (N_23969,N_15229,N_15950);
xnor U23970 (N_23970,N_13536,N_13124);
or U23971 (N_23971,N_14232,N_17728);
and U23972 (N_23972,N_15892,N_16549);
nand U23973 (N_23973,N_15747,N_17769);
nand U23974 (N_23974,N_17287,N_14150);
nor U23975 (N_23975,N_16830,N_12817);
xnor U23976 (N_23976,N_12612,N_14269);
nand U23977 (N_23977,N_17608,N_13838);
and U23978 (N_23978,N_12576,N_17080);
xor U23979 (N_23979,N_16047,N_17779);
nand U23980 (N_23980,N_15881,N_17857);
and U23981 (N_23981,N_16175,N_14536);
nand U23982 (N_23982,N_17098,N_17250);
and U23983 (N_23983,N_15374,N_16178);
and U23984 (N_23984,N_16019,N_12900);
nor U23985 (N_23985,N_16273,N_15094);
and U23986 (N_23986,N_17554,N_15300);
nand U23987 (N_23987,N_13399,N_16024);
nor U23988 (N_23988,N_17124,N_15137);
xnor U23989 (N_23989,N_13761,N_18705);
or U23990 (N_23990,N_18575,N_12961);
nand U23991 (N_23991,N_17343,N_12952);
or U23992 (N_23992,N_14635,N_17912);
nand U23993 (N_23993,N_17837,N_13118);
nand U23994 (N_23994,N_17552,N_13383);
nor U23995 (N_23995,N_16019,N_18561);
or U23996 (N_23996,N_15694,N_13967);
nor U23997 (N_23997,N_17856,N_14519);
or U23998 (N_23998,N_16947,N_15101);
xnor U23999 (N_23999,N_17494,N_12962);
nand U24000 (N_24000,N_14896,N_12544);
nand U24001 (N_24001,N_12590,N_18485);
nor U24002 (N_24002,N_13228,N_17470);
nand U24003 (N_24003,N_14516,N_17263);
nand U24004 (N_24004,N_14261,N_14844);
or U24005 (N_24005,N_17115,N_18072);
nand U24006 (N_24006,N_14397,N_12789);
nand U24007 (N_24007,N_17010,N_16215);
or U24008 (N_24008,N_18471,N_14122);
nor U24009 (N_24009,N_13883,N_14625);
and U24010 (N_24010,N_17235,N_16695);
and U24011 (N_24011,N_14738,N_18295);
xnor U24012 (N_24012,N_17950,N_15947);
nor U24013 (N_24013,N_15882,N_16585);
nand U24014 (N_24014,N_15038,N_13485);
nor U24015 (N_24015,N_13077,N_16692);
xnor U24016 (N_24016,N_16167,N_12894);
nand U24017 (N_24017,N_16525,N_13657);
and U24018 (N_24018,N_14912,N_16701);
or U24019 (N_24019,N_14597,N_16731);
or U24020 (N_24020,N_16393,N_15516);
and U24021 (N_24021,N_14865,N_18153);
xor U24022 (N_24022,N_12506,N_14383);
and U24023 (N_24023,N_18132,N_14810);
and U24024 (N_24024,N_15917,N_14609);
or U24025 (N_24025,N_13806,N_16655);
and U24026 (N_24026,N_16437,N_17559);
or U24027 (N_24027,N_17108,N_16640);
nand U24028 (N_24028,N_17260,N_16947);
nor U24029 (N_24029,N_15026,N_12901);
nor U24030 (N_24030,N_15588,N_13913);
and U24031 (N_24031,N_12959,N_16722);
nand U24032 (N_24032,N_16753,N_18266);
nor U24033 (N_24033,N_17333,N_18268);
xnor U24034 (N_24034,N_16037,N_16297);
xnor U24035 (N_24035,N_17171,N_16664);
nor U24036 (N_24036,N_13896,N_12922);
nand U24037 (N_24037,N_12590,N_13833);
nand U24038 (N_24038,N_18406,N_17267);
and U24039 (N_24039,N_15907,N_16201);
and U24040 (N_24040,N_17424,N_17062);
or U24041 (N_24041,N_13864,N_14269);
and U24042 (N_24042,N_13262,N_13461);
or U24043 (N_24043,N_18080,N_13048);
and U24044 (N_24044,N_13302,N_13236);
nor U24045 (N_24045,N_14513,N_15224);
and U24046 (N_24046,N_14811,N_17485);
or U24047 (N_24047,N_15254,N_13802);
nand U24048 (N_24048,N_16181,N_13571);
nor U24049 (N_24049,N_14760,N_17238);
and U24050 (N_24050,N_17452,N_12531);
and U24051 (N_24051,N_16896,N_17718);
xnor U24052 (N_24052,N_13980,N_13039);
nand U24053 (N_24053,N_13834,N_15433);
or U24054 (N_24054,N_16998,N_13818);
or U24055 (N_24055,N_17706,N_15992);
and U24056 (N_24056,N_13719,N_17030);
nor U24057 (N_24057,N_13238,N_12925);
or U24058 (N_24058,N_13571,N_17786);
nand U24059 (N_24059,N_18264,N_18599);
or U24060 (N_24060,N_13224,N_14432);
and U24061 (N_24061,N_16809,N_13284);
xnor U24062 (N_24062,N_17709,N_16625);
nand U24063 (N_24063,N_16697,N_14896);
nor U24064 (N_24064,N_12555,N_12620);
and U24065 (N_24065,N_15300,N_17415);
nor U24066 (N_24066,N_17761,N_13487);
nor U24067 (N_24067,N_14347,N_18317);
xor U24068 (N_24068,N_16637,N_16817);
nand U24069 (N_24069,N_16951,N_17965);
nand U24070 (N_24070,N_13626,N_12756);
nor U24071 (N_24071,N_13862,N_15218);
nor U24072 (N_24072,N_12867,N_17558);
or U24073 (N_24073,N_18037,N_16495);
or U24074 (N_24074,N_14631,N_14778);
nor U24075 (N_24075,N_12589,N_12879);
nor U24076 (N_24076,N_16490,N_14995);
nand U24077 (N_24077,N_16445,N_17511);
nand U24078 (N_24078,N_15850,N_18204);
nor U24079 (N_24079,N_17613,N_16712);
nor U24080 (N_24080,N_12545,N_18381);
or U24081 (N_24081,N_16285,N_13010);
nor U24082 (N_24082,N_18180,N_13601);
nand U24083 (N_24083,N_12557,N_15200);
and U24084 (N_24084,N_15060,N_13641);
nand U24085 (N_24085,N_14304,N_12906);
and U24086 (N_24086,N_15570,N_13845);
or U24087 (N_24087,N_17820,N_15759);
and U24088 (N_24088,N_16364,N_16575);
xor U24089 (N_24089,N_13079,N_16788);
and U24090 (N_24090,N_18395,N_16517);
and U24091 (N_24091,N_14183,N_13025);
nand U24092 (N_24092,N_16543,N_14013);
nand U24093 (N_24093,N_16461,N_13156);
and U24094 (N_24094,N_18157,N_18271);
or U24095 (N_24095,N_13157,N_15319);
and U24096 (N_24096,N_17360,N_15425);
nand U24097 (N_24097,N_16529,N_12919);
nor U24098 (N_24098,N_14226,N_13254);
nor U24099 (N_24099,N_15351,N_13342);
and U24100 (N_24100,N_17542,N_17061);
nor U24101 (N_24101,N_14968,N_14547);
nand U24102 (N_24102,N_14290,N_17252);
nand U24103 (N_24103,N_18571,N_13522);
or U24104 (N_24104,N_14526,N_17155);
nand U24105 (N_24105,N_15075,N_18528);
and U24106 (N_24106,N_16092,N_15507);
and U24107 (N_24107,N_16983,N_16607);
nand U24108 (N_24108,N_14960,N_17043);
or U24109 (N_24109,N_18221,N_14270);
nor U24110 (N_24110,N_12645,N_15898);
nor U24111 (N_24111,N_14908,N_12635);
nand U24112 (N_24112,N_17982,N_14292);
nor U24113 (N_24113,N_16677,N_16329);
nand U24114 (N_24114,N_13160,N_14636);
nand U24115 (N_24115,N_15918,N_14991);
or U24116 (N_24116,N_16080,N_15286);
and U24117 (N_24117,N_16088,N_13806);
and U24118 (N_24118,N_13669,N_12512);
nor U24119 (N_24119,N_16808,N_18427);
and U24120 (N_24120,N_17875,N_17080);
and U24121 (N_24121,N_18701,N_17137);
or U24122 (N_24122,N_13532,N_15635);
nand U24123 (N_24123,N_18236,N_15984);
xnor U24124 (N_24124,N_17936,N_13817);
nor U24125 (N_24125,N_14463,N_18313);
or U24126 (N_24126,N_12880,N_14334);
or U24127 (N_24127,N_14572,N_15460);
nand U24128 (N_24128,N_13413,N_17910);
or U24129 (N_24129,N_13090,N_16731);
or U24130 (N_24130,N_17194,N_17562);
nor U24131 (N_24131,N_18602,N_18262);
xor U24132 (N_24132,N_13769,N_15811);
nor U24133 (N_24133,N_16210,N_14116);
or U24134 (N_24134,N_17331,N_12670);
xnor U24135 (N_24135,N_13730,N_18693);
and U24136 (N_24136,N_16545,N_17476);
and U24137 (N_24137,N_14472,N_16032);
nand U24138 (N_24138,N_14983,N_18369);
xnor U24139 (N_24139,N_17927,N_15618);
or U24140 (N_24140,N_18677,N_18293);
and U24141 (N_24141,N_16042,N_13879);
nand U24142 (N_24142,N_16438,N_12582);
or U24143 (N_24143,N_12522,N_17349);
nor U24144 (N_24144,N_14115,N_17185);
nor U24145 (N_24145,N_18532,N_13019);
or U24146 (N_24146,N_17981,N_14274);
xor U24147 (N_24147,N_15112,N_14806);
or U24148 (N_24148,N_13948,N_15572);
xor U24149 (N_24149,N_18647,N_17866);
or U24150 (N_24150,N_12666,N_13315);
and U24151 (N_24151,N_14570,N_17970);
and U24152 (N_24152,N_12973,N_15880);
and U24153 (N_24153,N_14945,N_17106);
nor U24154 (N_24154,N_18617,N_18573);
or U24155 (N_24155,N_16941,N_18747);
xnor U24156 (N_24156,N_14109,N_16552);
nor U24157 (N_24157,N_18086,N_12899);
and U24158 (N_24158,N_14244,N_14283);
or U24159 (N_24159,N_17123,N_14221);
xor U24160 (N_24160,N_16845,N_17089);
nand U24161 (N_24161,N_16633,N_13989);
nor U24162 (N_24162,N_17644,N_14203);
or U24163 (N_24163,N_15428,N_15409);
nor U24164 (N_24164,N_16890,N_12556);
nor U24165 (N_24165,N_13428,N_17846);
nand U24166 (N_24166,N_14047,N_16148);
nand U24167 (N_24167,N_13990,N_12763);
nor U24168 (N_24168,N_16392,N_15121);
nand U24169 (N_24169,N_17032,N_15657);
or U24170 (N_24170,N_12590,N_13598);
or U24171 (N_24171,N_13907,N_17577);
and U24172 (N_24172,N_16054,N_18038);
nand U24173 (N_24173,N_18520,N_13507);
or U24174 (N_24174,N_13922,N_17915);
nand U24175 (N_24175,N_12799,N_15431);
xor U24176 (N_24176,N_18362,N_16414);
or U24177 (N_24177,N_16254,N_17878);
nand U24178 (N_24178,N_16808,N_16495);
nand U24179 (N_24179,N_16955,N_17722);
or U24180 (N_24180,N_14767,N_18344);
or U24181 (N_24181,N_18455,N_13978);
xor U24182 (N_24182,N_14330,N_13223);
and U24183 (N_24183,N_15090,N_13705);
or U24184 (N_24184,N_13011,N_16425);
nor U24185 (N_24185,N_16623,N_14337);
nand U24186 (N_24186,N_16198,N_17879);
and U24187 (N_24187,N_13886,N_17764);
nand U24188 (N_24188,N_16188,N_15900);
xor U24189 (N_24189,N_14055,N_12907);
nand U24190 (N_24190,N_12536,N_18577);
nor U24191 (N_24191,N_17688,N_15806);
xor U24192 (N_24192,N_15684,N_16706);
nand U24193 (N_24193,N_18464,N_17411);
or U24194 (N_24194,N_17492,N_14764);
or U24195 (N_24195,N_12804,N_14052);
and U24196 (N_24196,N_16354,N_17923);
or U24197 (N_24197,N_17638,N_15533);
or U24198 (N_24198,N_12604,N_17654);
xor U24199 (N_24199,N_12631,N_13773);
nand U24200 (N_24200,N_13712,N_16275);
and U24201 (N_24201,N_17039,N_14756);
nand U24202 (N_24202,N_17691,N_18274);
nand U24203 (N_24203,N_18303,N_14622);
and U24204 (N_24204,N_15407,N_13528);
and U24205 (N_24205,N_18103,N_18650);
xor U24206 (N_24206,N_13236,N_12780);
nand U24207 (N_24207,N_15400,N_12611);
and U24208 (N_24208,N_17967,N_18453);
and U24209 (N_24209,N_14270,N_18533);
or U24210 (N_24210,N_13525,N_13848);
xnor U24211 (N_24211,N_16971,N_12794);
and U24212 (N_24212,N_16959,N_14458);
or U24213 (N_24213,N_12635,N_17227);
or U24214 (N_24214,N_17494,N_16603);
nand U24215 (N_24215,N_16160,N_15877);
xor U24216 (N_24216,N_13033,N_14600);
nand U24217 (N_24217,N_18375,N_17099);
and U24218 (N_24218,N_16047,N_12526);
nor U24219 (N_24219,N_13873,N_12569);
xnor U24220 (N_24220,N_13644,N_17337);
and U24221 (N_24221,N_12906,N_18501);
xor U24222 (N_24222,N_12671,N_16914);
or U24223 (N_24223,N_17927,N_15372);
nor U24224 (N_24224,N_15127,N_17429);
nor U24225 (N_24225,N_17806,N_16807);
and U24226 (N_24226,N_17471,N_16719);
nor U24227 (N_24227,N_16444,N_16793);
or U24228 (N_24228,N_14879,N_18257);
and U24229 (N_24229,N_15490,N_12551);
nor U24230 (N_24230,N_15673,N_13384);
nand U24231 (N_24231,N_16269,N_15945);
nor U24232 (N_24232,N_12731,N_18152);
or U24233 (N_24233,N_14927,N_15541);
nand U24234 (N_24234,N_17672,N_15013);
and U24235 (N_24235,N_16139,N_17769);
or U24236 (N_24236,N_17456,N_17141);
xor U24237 (N_24237,N_13627,N_18015);
and U24238 (N_24238,N_17601,N_17155);
and U24239 (N_24239,N_15135,N_16441);
and U24240 (N_24240,N_14044,N_17342);
nand U24241 (N_24241,N_17303,N_15525);
and U24242 (N_24242,N_17642,N_16393);
nand U24243 (N_24243,N_17008,N_12928);
nand U24244 (N_24244,N_12836,N_16739);
nor U24245 (N_24245,N_12761,N_18009);
nor U24246 (N_24246,N_15340,N_17329);
or U24247 (N_24247,N_18249,N_14063);
or U24248 (N_24248,N_13524,N_14869);
and U24249 (N_24249,N_13467,N_17752);
nor U24250 (N_24250,N_16370,N_17580);
nor U24251 (N_24251,N_15557,N_18242);
or U24252 (N_24252,N_17347,N_17648);
nand U24253 (N_24253,N_18697,N_16818);
xor U24254 (N_24254,N_17478,N_14804);
nor U24255 (N_24255,N_17997,N_15860);
xnor U24256 (N_24256,N_17547,N_14137);
or U24257 (N_24257,N_14800,N_18505);
or U24258 (N_24258,N_17859,N_15640);
nand U24259 (N_24259,N_15969,N_16108);
xor U24260 (N_24260,N_18279,N_16556);
xor U24261 (N_24261,N_16336,N_18715);
nand U24262 (N_24262,N_13721,N_17737);
and U24263 (N_24263,N_13945,N_13574);
nand U24264 (N_24264,N_16424,N_18098);
nand U24265 (N_24265,N_16355,N_13434);
nor U24266 (N_24266,N_14757,N_16706);
nor U24267 (N_24267,N_12587,N_12570);
nand U24268 (N_24268,N_15362,N_14315);
or U24269 (N_24269,N_17396,N_15091);
or U24270 (N_24270,N_16357,N_13773);
nor U24271 (N_24271,N_18007,N_13461);
nor U24272 (N_24272,N_15700,N_18535);
and U24273 (N_24273,N_14033,N_13460);
nor U24274 (N_24274,N_18719,N_13615);
and U24275 (N_24275,N_17934,N_15594);
or U24276 (N_24276,N_18499,N_18070);
nor U24277 (N_24277,N_14853,N_18127);
nand U24278 (N_24278,N_12523,N_14365);
nor U24279 (N_24279,N_13279,N_15746);
or U24280 (N_24280,N_14538,N_17446);
xnor U24281 (N_24281,N_17893,N_15420);
xnor U24282 (N_24282,N_13909,N_12707);
nand U24283 (N_24283,N_17976,N_17172);
nand U24284 (N_24284,N_16629,N_15998);
nand U24285 (N_24285,N_14206,N_18401);
or U24286 (N_24286,N_18407,N_18509);
and U24287 (N_24287,N_15454,N_16072);
nor U24288 (N_24288,N_15162,N_17038);
or U24289 (N_24289,N_17760,N_18391);
nand U24290 (N_24290,N_12595,N_17047);
nor U24291 (N_24291,N_15738,N_18068);
or U24292 (N_24292,N_13853,N_18363);
or U24293 (N_24293,N_13342,N_16405);
and U24294 (N_24294,N_16460,N_17960);
nor U24295 (N_24295,N_17866,N_14945);
xnor U24296 (N_24296,N_18458,N_15056);
nand U24297 (N_24297,N_15983,N_17158);
xnor U24298 (N_24298,N_17702,N_18718);
and U24299 (N_24299,N_18038,N_13569);
or U24300 (N_24300,N_18413,N_14739);
nand U24301 (N_24301,N_13172,N_12653);
xnor U24302 (N_24302,N_14838,N_15012);
xor U24303 (N_24303,N_13929,N_16212);
or U24304 (N_24304,N_17180,N_18021);
and U24305 (N_24305,N_18560,N_16466);
xor U24306 (N_24306,N_14768,N_18261);
xnor U24307 (N_24307,N_15311,N_18029);
nor U24308 (N_24308,N_14217,N_16746);
nand U24309 (N_24309,N_17679,N_17091);
xor U24310 (N_24310,N_15434,N_15701);
nor U24311 (N_24311,N_17028,N_16685);
nand U24312 (N_24312,N_13032,N_14442);
xor U24313 (N_24313,N_14476,N_14920);
nor U24314 (N_24314,N_17075,N_15972);
nand U24315 (N_24315,N_14234,N_16531);
nor U24316 (N_24316,N_18469,N_14928);
nor U24317 (N_24317,N_14077,N_17548);
nor U24318 (N_24318,N_17625,N_18483);
nand U24319 (N_24319,N_18640,N_16089);
nand U24320 (N_24320,N_18364,N_12676);
and U24321 (N_24321,N_14017,N_14219);
and U24322 (N_24322,N_16907,N_13549);
or U24323 (N_24323,N_15056,N_14687);
or U24324 (N_24324,N_15709,N_17403);
and U24325 (N_24325,N_17955,N_13476);
or U24326 (N_24326,N_17936,N_16858);
xor U24327 (N_24327,N_15883,N_12726);
and U24328 (N_24328,N_15493,N_13983);
nor U24329 (N_24329,N_13845,N_16815);
nor U24330 (N_24330,N_17051,N_16178);
and U24331 (N_24331,N_17252,N_13652);
or U24332 (N_24332,N_13558,N_13437);
nor U24333 (N_24333,N_16839,N_14278);
nor U24334 (N_24334,N_14726,N_16382);
nand U24335 (N_24335,N_12808,N_15423);
or U24336 (N_24336,N_17277,N_18450);
or U24337 (N_24337,N_17302,N_16746);
or U24338 (N_24338,N_17035,N_18232);
nor U24339 (N_24339,N_15330,N_16683);
nor U24340 (N_24340,N_18367,N_17039);
nor U24341 (N_24341,N_17439,N_18402);
nand U24342 (N_24342,N_17991,N_14384);
and U24343 (N_24343,N_12853,N_15244);
nand U24344 (N_24344,N_13020,N_13230);
and U24345 (N_24345,N_18630,N_13007);
or U24346 (N_24346,N_16529,N_15635);
nand U24347 (N_24347,N_14901,N_14955);
nand U24348 (N_24348,N_15439,N_16757);
nor U24349 (N_24349,N_18263,N_14784);
or U24350 (N_24350,N_16024,N_17212);
nand U24351 (N_24351,N_16119,N_18467);
and U24352 (N_24352,N_13481,N_13263);
or U24353 (N_24353,N_17160,N_17211);
and U24354 (N_24354,N_15913,N_17760);
xnor U24355 (N_24355,N_12690,N_15679);
or U24356 (N_24356,N_13664,N_18483);
nor U24357 (N_24357,N_12790,N_18625);
nor U24358 (N_24358,N_17195,N_15744);
nand U24359 (N_24359,N_13580,N_13608);
nand U24360 (N_24360,N_14712,N_16387);
xor U24361 (N_24361,N_16757,N_13533);
or U24362 (N_24362,N_15414,N_16868);
nor U24363 (N_24363,N_14022,N_14908);
nor U24364 (N_24364,N_15016,N_14886);
nand U24365 (N_24365,N_12829,N_14849);
xor U24366 (N_24366,N_15389,N_16916);
nand U24367 (N_24367,N_16701,N_17873);
nand U24368 (N_24368,N_15406,N_17518);
nor U24369 (N_24369,N_17060,N_15570);
or U24370 (N_24370,N_14896,N_17419);
or U24371 (N_24371,N_14040,N_17536);
or U24372 (N_24372,N_17282,N_13144);
xnor U24373 (N_24373,N_16107,N_12934);
xor U24374 (N_24374,N_14849,N_18387);
nor U24375 (N_24375,N_16509,N_15982);
or U24376 (N_24376,N_17732,N_13701);
or U24377 (N_24377,N_14186,N_16060);
xnor U24378 (N_24378,N_14705,N_18380);
or U24379 (N_24379,N_15521,N_15288);
or U24380 (N_24380,N_16347,N_16206);
and U24381 (N_24381,N_12503,N_12866);
nor U24382 (N_24382,N_17698,N_16314);
nand U24383 (N_24383,N_17191,N_13165);
or U24384 (N_24384,N_14526,N_18333);
xnor U24385 (N_24385,N_18428,N_16272);
nor U24386 (N_24386,N_13122,N_13443);
or U24387 (N_24387,N_16705,N_15089);
nor U24388 (N_24388,N_13870,N_13810);
and U24389 (N_24389,N_15668,N_15772);
and U24390 (N_24390,N_17410,N_17451);
nor U24391 (N_24391,N_16308,N_17229);
nand U24392 (N_24392,N_16907,N_13113);
nor U24393 (N_24393,N_16957,N_15851);
and U24394 (N_24394,N_18074,N_14461);
and U24395 (N_24395,N_13226,N_12951);
or U24396 (N_24396,N_12638,N_15538);
or U24397 (N_24397,N_18502,N_14442);
nand U24398 (N_24398,N_12537,N_16874);
xnor U24399 (N_24399,N_13145,N_16054);
or U24400 (N_24400,N_16915,N_18568);
and U24401 (N_24401,N_14449,N_12933);
and U24402 (N_24402,N_14874,N_14694);
or U24403 (N_24403,N_18102,N_17963);
nand U24404 (N_24404,N_14246,N_17211);
or U24405 (N_24405,N_16549,N_12753);
nor U24406 (N_24406,N_15921,N_15486);
nand U24407 (N_24407,N_13492,N_18093);
nor U24408 (N_24408,N_17879,N_13928);
and U24409 (N_24409,N_15163,N_17085);
and U24410 (N_24410,N_16526,N_17430);
xnor U24411 (N_24411,N_17415,N_17929);
nand U24412 (N_24412,N_17729,N_16670);
nor U24413 (N_24413,N_16819,N_13264);
nor U24414 (N_24414,N_12910,N_18691);
and U24415 (N_24415,N_12505,N_14845);
and U24416 (N_24416,N_16487,N_14382);
or U24417 (N_24417,N_13872,N_14816);
nand U24418 (N_24418,N_18729,N_13353);
and U24419 (N_24419,N_12500,N_12801);
or U24420 (N_24420,N_13138,N_16829);
and U24421 (N_24421,N_15783,N_15454);
nor U24422 (N_24422,N_18251,N_18064);
or U24423 (N_24423,N_13269,N_18707);
or U24424 (N_24424,N_17666,N_18075);
nand U24425 (N_24425,N_14620,N_16173);
or U24426 (N_24426,N_14732,N_14828);
and U24427 (N_24427,N_12885,N_15497);
or U24428 (N_24428,N_15310,N_17624);
nor U24429 (N_24429,N_14864,N_14789);
and U24430 (N_24430,N_18361,N_13724);
nand U24431 (N_24431,N_15538,N_13723);
nor U24432 (N_24432,N_13831,N_18094);
nor U24433 (N_24433,N_12560,N_14363);
nand U24434 (N_24434,N_12612,N_12936);
nor U24435 (N_24435,N_14266,N_13121);
xor U24436 (N_24436,N_15468,N_13007);
and U24437 (N_24437,N_15040,N_13775);
nand U24438 (N_24438,N_14157,N_18423);
and U24439 (N_24439,N_18478,N_14547);
or U24440 (N_24440,N_15181,N_12878);
nor U24441 (N_24441,N_14388,N_16074);
or U24442 (N_24442,N_15334,N_17718);
nand U24443 (N_24443,N_15407,N_13963);
nand U24444 (N_24444,N_17218,N_16080);
nand U24445 (N_24445,N_12819,N_17758);
nor U24446 (N_24446,N_17186,N_16575);
nand U24447 (N_24447,N_14086,N_18465);
nor U24448 (N_24448,N_13432,N_13874);
xor U24449 (N_24449,N_14920,N_12914);
nand U24450 (N_24450,N_16608,N_18456);
or U24451 (N_24451,N_14215,N_16995);
nand U24452 (N_24452,N_17749,N_15609);
nor U24453 (N_24453,N_18597,N_15182);
nand U24454 (N_24454,N_13606,N_13881);
xnor U24455 (N_24455,N_14358,N_14676);
nor U24456 (N_24456,N_13559,N_12775);
and U24457 (N_24457,N_16858,N_15497);
nand U24458 (N_24458,N_13692,N_17646);
or U24459 (N_24459,N_17018,N_17711);
or U24460 (N_24460,N_18251,N_14606);
xnor U24461 (N_24461,N_17857,N_15556);
or U24462 (N_24462,N_13315,N_13080);
nor U24463 (N_24463,N_13999,N_16308);
nor U24464 (N_24464,N_17803,N_18413);
and U24465 (N_24465,N_12503,N_17560);
nand U24466 (N_24466,N_17546,N_14650);
nor U24467 (N_24467,N_13709,N_13885);
nand U24468 (N_24468,N_15750,N_14576);
or U24469 (N_24469,N_16351,N_17636);
or U24470 (N_24470,N_12694,N_16522);
nand U24471 (N_24471,N_16233,N_13604);
and U24472 (N_24472,N_15757,N_17488);
nor U24473 (N_24473,N_16771,N_12683);
xor U24474 (N_24474,N_18450,N_18741);
nand U24475 (N_24475,N_14300,N_16599);
or U24476 (N_24476,N_14023,N_15804);
nand U24477 (N_24477,N_12692,N_15237);
or U24478 (N_24478,N_12572,N_13896);
xor U24479 (N_24479,N_12778,N_16917);
nand U24480 (N_24480,N_16881,N_18207);
and U24481 (N_24481,N_13050,N_13789);
or U24482 (N_24482,N_15397,N_16123);
xnor U24483 (N_24483,N_14883,N_13575);
nor U24484 (N_24484,N_17941,N_13131);
or U24485 (N_24485,N_13059,N_12581);
xor U24486 (N_24486,N_18419,N_14023);
or U24487 (N_24487,N_15267,N_15941);
or U24488 (N_24488,N_15506,N_16905);
and U24489 (N_24489,N_14033,N_16718);
and U24490 (N_24490,N_16386,N_16407);
and U24491 (N_24491,N_13516,N_16467);
or U24492 (N_24492,N_13515,N_15739);
or U24493 (N_24493,N_16596,N_17046);
nand U24494 (N_24494,N_18587,N_13193);
nand U24495 (N_24495,N_16728,N_16080);
or U24496 (N_24496,N_14950,N_13732);
nor U24497 (N_24497,N_12593,N_13621);
nand U24498 (N_24498,N_13585,N_15920);
nor U24499 (N_24499,N_13580,N_12931);
or U24500 (N_24500,N_13564,N_17347);
or U24501 (N_24501,N_16144,N_16131);
nor U24502 (N_24502,N_18543,N_15249);
nand U24503 (N_24503,N_17646,N_16503);
nand U24504 (N_24504,N_12515,N_18705);
nor U24505 (N_24505,N_13928,N_13318);
nor U24506 (N_24506,N_15469,N_14389);
or U24507 (N_24507,N_16753,N_17911);
or U24508 (N_24508,N_17416,N_13213);
nor U24509 (N_24509,N_15224,N_18119);
nand U24510 (N_24510,N_13371,N_15133);
nor U24511 (N_24511,N_14861,N_15345);
nor U24512 (N_24512,N_13355,N_16049);
and U24513 (N_24513,N_18425,N_15204);
and U24514 (N_24514,N_15641,N_13159);
nand U24515 (N_24515,N_16207,N_13067);
nand U24516 (N_24516,N_15187,N_16519);
or U24517 (N_24517,N_17356,N_16213);
and U24518 (N_24518,N_13169,N_15360);
xnor U24519 (N_24519,N_15841,N_17648);
nor U24520 (N_24520,N_16933,N_14295);
and U24521 (N_24521,N_16843,N_17840);
or U24522 (N_24522,N_16133,N_18183);
or U24523 (N_24523,N_14220,N_13741);
and U24524 (N_24524,N_15487,N_15635);
nor U24525 (N_24525,N_14183,N_13389);
xor U24526 (N_24526,N_14667,N_12852);
xnor U24527 (N_24527,N_13820,N_16006);
or U24528 (N_24528,N_15689,N_18654);
nor U24529 (N_24529,N_16699,N_15226);
or U24530 (N_24530,N_13691,N_18339);
xor U24531 (N_24531,N_14672,N_14684);
xor U24532 (N_24532,N_14138,N_14303);
and U24533 (N_24533,N_17521,N_15562);
nor U24534 (N_24534,N_16510,N_17690);
nor U24535 (N_24535,N_16037,N_13066);
nand U24536 (N_24536,N_15878,N_15460);
nor U24537 (N_24537,N_13022,N_15067);
nor U24538 (N_24538,N_13155,N_18381);
or U24539 (N_24539,N_13688,N_14747);
nand U24540 (N_24540,N_17582,N_12759);
and U24541 (N_24541,N_15325,N_14020);
nor U24542 (N_24542,N_14755,N_13835);
nand U24543 (N_24543,N_18589,N_18662);
nor U24544 (N_24544,N_13750,N_13070);
and U24545 (N_24545,N_16540,N_17112);
and U24546 (N_24546,N_16539,N_17289);
nor U24547 (N_24547,N_18251,N_17560);
nor U24548 (N_24548,N_13132,N_17293);
and U24549 (N_24549,N_17977,N_13083);
nand U24550 (N_24550,N_14304,N_15477);
and U24551 (N_24551,N_15692,N_16730);
and U24552 (N_24552,N_18088,N_16107);
and U24553 (N_24553,N_13897,N_16722);
or U24554 (N_24554,N_18197,N_13556);
xnor U24555 (N_24555,N_16456,N_13780);
or U24556 (N_24556,N_17020,N_18217);
nor U24557 (N_24557,N_18026,N_16969);
and U24558 (N_24558,N_15538,N_17210);
and U24559 (N_24559,N_15662,N_13399);
xnor U24560 (N_24560,N_15868,N_14669);
and U24561 (N_24561,N_17820,N_13238);
or U24562 (N_24562,N_17256,N_18597);
xnor U24563 (N_24563,N_14521,N_17996);
or U24564 (N_24564,N_16266,N_15061);
nor U24565 (N_24565,N_17750,N_17770);
nor U24566 (N_24566,N_15256,N_15637);
xnor U24567 (N_24567,N_17480,N_16471);
xor U24568 (N_24568,N_13975,N_17224);
nand U24569 (N_24569,N_17882,N_15747);
nor U24570 (N_24570,N_18362,N_15617);
nor U24571 (N_24571,N_14837,N_13182);
and U24572 (N_24572,N_13209,N_13640);
and U24573 (N_24573,N_14907,N_16335);
or U24574 (N_24574,N_14445,N_13938);
and U24575 (N_24575,N_17036,N_17517);
or U24576 (N_24576,N_16932,N_13286);
or U24577 (N_24577,N_12841,N_13143);
or U24578 (N_24578,N_18158,N_15692);
nor U24579 (N_24579,N_16421,N_17106);
nor U24580 (N_24580,N_12825,N_14872);
or U24581 (N_24581,N_17281,N_16249);
nor U24582 (N_24582,N_13583,N_17017);
or U24583 (N_24583,N_16979,N_15341);
nand U24584 (N_24584,N_14051,N_12656);
nand U24585 (N_24585,N_13292,N_16884);
nor U24586 (N_24586,N_13960,N_17999);
xnor U24587 (N_24587,N_18084,N_13471);
nor U24588 (N_24588,N_17669,N_14333);
nand U24589 (N_24589,N_13799,N_18692);
or U24590 (N_24590,N_15042,N_13739);
or U24591 (N_24591,N_13678,N_12554);
and U24592 (N_24592,N_12634,N_14869);
or U24593 (N_24593,N_18496,N_15896);
and U24594 (N_24594,N_13296,N_18121);
or U24595 (N_24595,N_13399,N_17343);
or U24596 (N_24596,N_12728,N_17471);
nor U24597 (N_24597,N_17781,N_14730);
nand U24598 (N_24598,N_18470,N_15143);
and U24599 (N_24599,N_14522,N_12736);
or U24600 (N_24600,N_13557,N_17429);
nand U24601 (N_24601,N_15800,N_13566);
or U24602 (N_24602,N_14240,N_18205);
or U24603 (N_24603,N_17716,N_17091);
nand U24604 (N_24604,N_12905,N_15357);
or U24605 (N_24605,N_16101,N_16312);
and U24606 (N_24606,N_16125,N_18445);
or U24607 (N_24607,N_17915,N_16521);
and U24608 (N_24608,N_17815,N_17990);
and U24609 (N_24609,N_12504,N_15144);
nand U24610 (N_24610,N_15617,N_13303);
xor U24611 (N_24611,N_17983,N_14285);
nor U24612 (N_24612,N_15992,N_13995);
xor U24613 (N_24613,N_15613,N_16344);
or U24614 (N_24614,N_15300,N_14880);
or U24615 (N_24615,N_17413,N_17414);
xnor U24616 (N_24616,N_17733,N_18714);
nand U24617 (N_24617,N_15751,N_18339);
and U24618 (N_24618,N_14050,N_15541);
nor U24619 (N_24619,N_14749,N_13203);
nor U24620 (N_24620,N_13413,N_17255);
and U24621 (N_24621,N_18352,N_18278);
nand U24622 (N_24622,N_14899,N_15679);
or U24623 (N_24623,N_17999,N_18710);
or U24624 (N_24624,N_15007,N_18332);
and U24625 (N_24625,N_17767,N_17018);
and U24626 (N_24626,N_16418,N_17855);
nor U24627 (N_24627,N_12800,N_16239);
nand U24628 (N_24628,N_13813,N_17857);
and U24629 (N_24629,N_14706,N_17743);
nand U24630 (N_24630,N_14189,N_15122);
xnor U24631 (N_24631,N_15317,N_17730);
nand U24632 (N_24632,N_13277,N_17946);
nand U24633 (N_24633,N_15613,N_15778);
nor U24634 (N_24634,N_16891,N_18729);
nand U24635 (N_24635,N_14110,N_16287);
nor U24636 (N_24636,N_12867,N_17799);
or U24637 (N_24637,N_18100,N_18199);
and U24638 (N_24638,N_17986,N_18676);
and U24639 (N_24639,N_13866,N_15263);
nor U24640 (N_24640,N_15039,N_16839);
and U24641 (N_24641,N_16633,N_13257);
nor U24642 (N_24642,N_12922,N_18710);
xor U24643 (N_24643,N_18291,N_17157);
or U24644 (N_24644,N_16377,N_14014);
nor U24645 (N_24645,N_13062,N_13557);
nand U24646 (N_24646,N_12725,N_15736);
or U24647 (N_24647,N_15602,N_13128);
or U24648 (N_24648,N_14938,N_16328);
nor U24649 (N_24649,N_15432,N_16697);
nor U24650 (N_24650,N_12653,N_17641);
nand U24651 (N_24651,N_14096,N_12805);
xnor U24652 (N_24652,N_14860,N_15618);
nor U24653 (N_24653,N_12880,N_15552);
nor U24654 (N_24654,N_18281,N_16607);
and U24655 (N_24655,N_15188,N_12980);
and U24656 (N_24656,N_18247,N_12970);
nor U24657 (N_24657,N_18107,N_14920);
or U24658 (N_24658,N_12784,N_17263);
nor U24659 (N_24659,N_16351,N_13700);
nand U24660 (N_24660,N_14179,N_15506);
xor U24661 (N_24661,N_12981,N_12638);
and U24662 (N_24662,N_15066,N_15010);
nor U24663 (N_24663,N_17472,N_14345);
xnor U24664 (N_24664,N_13767,N_15540);
nand U24665 (N_24665,N_16996,N_16673);
nand U24666 (N_24666,N_16378,N_16458);
nand U24667 (N_24667,N_14249,N_17727);
and U24668 (N_24668,N_12939,N_16328);
nor U24669 (N_24669,N_16384,N_13193);
xnor U24670 (N_24670,N_18382,N_13855);
xnor U24671 (N_24671,N_15883,N_17821);
and U24672 (N_24672,N_16752,N_13354);
and U24673 (N_24673,N_12604,N_13175);
or U24674 (N_24674,N_17795,N_13652);
nand U24675 (N_24675,N_15753,N_12756);
and U24676 (N_24676,N_13957,N_15812);
or U24677 (N_24677,N_15223,N_12767);
nand U24678 (N_24678,N_15420,N_12743);
or U24679 (N_24679,N_17391,N_12913);
and U24680 (N_24680,N_14594,N_12699);
nand U24681 (N_24681,N_17408,N_15528);
or U24682 (N_24682,N_14763,N_14529);
or U24683 (N_24683,N_12960,N_15242);
nand U24684 (N_24684,N_14256,N_13874);
and U24685 (N_24685,N_14160,N_17573);
or U24686 (N_24686,N_15155,N_16221);
xnor U24687 (N_24687,N_13890,N_14327);
or U24688 (N_24688,N_13284,N_12919);
xnor U24689 (N_24689,N_16326,N_12828);
and U24690 (N_24690,N_16365,N_17084);
nand U24691 (N_24691,N_16367,N_17846);
or U24692 (N_24692,N_15618,N_12971);
or U24693 (N_24693,N_13910,N_13822);
xnor U24694 (N_24694,N_13873,N_12545);
and U24695 (N_24695,N_13312,N_14657);
and U24696 (N_24696,N_18633,N_16952);
and U24697 (N_24697,N_18640,N_13786);
nor U24698 (N_24698,N_13221,N_16553);
nand U24699 (N_24699,N_16599,N_14069);
nand U24700 (N_24700,N_13677,N_18186);
nor U24701 (N_24701,N_15628,N_15526);
nor U24702 (N_24702,N_15496,N_17002);
or U24703 (N_24703,N_18432,N_17362);
and U24704 (N_24704,N_16192,N_14983);
nor U24705 (N_24705,N_13823,N_13572);
and U24706 (N_24706,N_14654,N_18012);
nor U24707 (N_24707,N_13312,N_14695);
or U24708 (N_24708,N_16974,N_14321);
or U24709 (N_24709,N_18639,N_13671);
and U24710 (N_24710,N_18608,N_15174);
nand U24711 (N_24711,N_13066,N_18383);
and U24712 (N_24712,N_17368,N_14697);
nand U24713 (N_24713,N_12513,N_16792);
nor U24714 (N_24714,N_18511,N_13317);
nand U24715 (N_24715,N_17868,N_12865);
and U24716 (N_24716,N_13407,N_17175);
or U24717 (N_24717,N_17192,N_16403);
nand U24718 (N_24718,N_17087,N_16229);
nand U24719 (N_24719,N_16480,N_16670);
nand U24720 (N_24720,N_13223,N_14706);
or U24721 (N_24721,N_12658,N_17366);
nand U24722 (N_24722,N_13758,N_16902);
nand U24723 (N_24723,N_13811,N_14927);
nand U24724 (N_24724,N_18308,N_12571);
and U24725 (N_24725,N_17692,N_17799);
nand U24726 (N_24726,N_14869,N_17656);
nand U24727 (N_24727,N_13011,N_15378);
nor U24728 (N_24728,N_16194,N_14283);
and U24729 (N_24729,N_15989,N_18417);
xor U24730 (N_24730,N_15905,N_12939);
nand U24731 (N_24731,N_17185,N_12604);
or U24732 (N_24732,N_13457,N_14877);
and U24733 (N_24733,N_18660,N_16334);
and U24734 (N_24734,N_17091,N_12786);
and U24735 (N_24735,N_17493,N_15138);
or U24736 (N_24736,N_18328,N_12849);
and U24737 (N_24737,N_14417,N_13768);
nand U24738 (N_24738,N_14026,N_13613);
nor U24739 (N_24739,N_12862,N_15482);
nand U24740 (N_24740,N_15866,N_13698);
and U24741 (N_24741,N_18298,N_17490);
nand U24742 (N_24742,N_13917,N_13478);
nor U24743 (N_24743,N_16106,N_13067);
and U24744 (N_24744,N_15953,N_13884);
xnor U24745 (N_24745,N_15638,N_13500);
nor U24746 (N_24746,N_15771,N_14864);
xnor U24747 (N_24747,N_18122,N_16742);
or U24748 (N_24748,N_17251,N_16071);
xor U24749 (N_24749,N_14763,N_16902);
xnor U24750 (N_24750,N_16019,N_17477);
or U24751 (N_24751,N_12635,N_16603);
nand U24752 (N_24752,N_15563,N_12720);
nor U24753 (N_24753,N_15486,N_18057);
nor U24754 (N_24754,N_15117,N_13131);
xor U24755 (N_24755,N_12595,N_17095);
nand U24756 (N_24756,N_13964,N_13010);
nand U24757 (N_24757,N_14086,N_16494);
xnor U24758 (N_24758,N_16759,N_12521);
and U24759 (N_24759,N_14842,N_12947);
nand U24760 (N_24760,N_16649,N_13904);
xnor U24761 (N_24761,N_17790,N_17762);
or U24762 (N_24762,N_17214,N_13694);
xnor U24763 (N_24763,N_16185,N_12834);
nor U24764 (N_24764,N_14263,N_15808);
nand U24765 (N_24765,N_17043,N_17969);
nand U24766 (N_24766,N_13679,N_17113);
nand U24767 (N_24767,N_14420,N_13716);
nand U24768 (N_24768,N_16143,N_17563);
nor U24769 (N_24769,N_15966,N_13025);
or U24770 (N_24770,N_14745,N_16488);
nand U24771 (N_24771,N_13554,N_17103);
or U24772 (N_24772,N_13562,N_13436);
nor U24773 (N_24773,N_17829,N_13058);
nand U24774 (N_24774,N_18327,N_15653);
and U24775 (N_24775,N_12830,N_13505);
nand U24776 (N_24776,N_16726,N_14366);
nor U24777 (N_24777,N_13536,N_12635);
nor U24778 (N_24778,N_14765,N_13569);
nor U24779 (N_24779,N_18010,N_16386);
nand U24780 (N_24780,N_13007,N_14052);
nor U24781 (N_24781,N_13408,N_12774);
or U24782 (N_24782,N_17607,N_17316);
or U24783 (N_24783,N_13174,N_13190);
nand U24784 (N_24784,N_13077,N_15010);
nand U24785 (N_24785,N_18161,N_16510);
and U24786 (N_24786,N_13031,N_15381);
or U24787 (N_24787,N_13497,N_18556);
and U24788 (N_24788,N_12543,N_18039);
or U24789 (N_24789,N_16575,N_15200);
and U24790 (N_24790,N_16272,N_17700);
or U24791 (N_24791,N_13980,N_16627);
xor U24792 (N_24792,N_17592,N_15698);
nand U24793 (N_24793,N_15517,N_18317);
xnor U24794 (N_24794,N_17081,N_17612);
or U24795 (N_24795,N_15609,N_14139);
xor U24796 (N_24796,N_14485,N_17411);
or U24797 (N_24797,N_14752,N_15146);
or U24798 (N_24798,N_17934,N_13232);
nor U24799 (N_24799,N_14239,N_16011);
nand U24800 (N_24800,N_17135,N_14811);
and U24801 (N_24801,N_17938,N_14300);
nand U24802 (N_24802,N_12658,N_15802);
or U24803 (N_24803,N_18475,N_16960);
nor U24804 (N_24804,N_18272,N_15720);
or U24805 (N_24805,N_14986,N_18139);
or U24806 (N_24806,N_14044,N_13911);
nor U24807 (N_24807,N_16768,N_14044);
or U24808 (N_24808,N_13631,N_16526);
and U24809 (N_24809,N_12677,N_12627);
or U24810 (N_24810,N_16610,N_16903);
nand U24811 (N_24811,N_18326,N_13816);
nand U24812 (N_24812,N_15784,N_16763);
nor U24813 (N_24813,N_14787,N_12915);
nand U24814 (N_24814,N_15468,N_15772);
and U24815 (N_24815,N_15959,N_16824);
or U24816 (N_24816,N_13127,N_16230);
nor U24817 (N_24817,N_15143,N_15466);
nor U24818 (N_24818,N_12751,N_17652);
and U24819 (N_24819,N_13008,N_12655);
nand U24820 (N_24820,N_16434,N_15694);
nor U24821 (N_24821,N_17949,N_14319);
or U24822 (N_24822,N_18564,N_17327);
nand U24823 (N_24823,N_14952,N_14716);
and U24824 (N_24824,N_17378,N_16196);
nor U24825 (N_24825,N_13284,N_17585);
or U24826 (N_24826,N_12688,N_12756);
or U24827 (N_24827,N_14528,N_15205);
nor U24828 (N_24828,N_13144,N_15678);
nand U24829 (N_24829,N_15274,N_15911);
nor U24830 (N_24830,N_14523,N_15648);
nor U24831 (N_24831,N_17118,N_13428);
nand U24832 (N_24832,N_12917,N_16706);
nor U24833 (N_24833,N_14612,N_17008);
nand U24834 (N_24834,N_16214,N_17937);
and U24835 (N_24835,N_16446,N_14864);
or U24836 (N_24836,N_13853,N_15158);
and U24837 (N_24837,N_12992,N_13036);
nand U24838 (N_24838,N_17452,N_16252);
and U24839 (N_24839,N_17952,N_15063);
nor U24840 (N_24840,N_16682,N_16458);
xnor U24841 (N_24841,N_18102,N_13512);
nand U24842 (N_24842,N_13435,N_13172);
nand U24843 (N_24843,N_16273,N_18188);
nor U24844 (N_24844,N_12632,N_13220);
nand U24845 (N_24845,N_18526,N_15162);
nor U24846 (N_24846,N_15485,N_18497);
xnor U24847 (N_24847,N_15749,N_14442);
nand U24848 (N_24848,N_17032,N_16221);
or U24849 (N_24849,N_16319,N_16701);
and U24850 (N_24850,N_15858,N_13691);
or U24851 (N_24851,N_16976,N_16654);
nor U24852 (N_24852,N_14274,N_14489);
nor U24853 (N_24853,N_18235,N_18459);
or U24854 (N_24854,N_16728,N_17374);
nand U24855 (N_24855,N_14532,N_17359);
nand U24856 (N_24856,N_15403,N_14139);
or U24857 (N_24857,N_15949,N_12854);
and U24858 (N_24858,N_15096,N_13487);
nor U24859 (N_24859,N_18442,N_17443);
or U24860 (N_24860,N_14303,N_16991);
and U24861 (N_24861,N_17915,N_13472);
nand U24862 (N_24862,N_16133,N_18122);
or U24863 (N_24863,N_13243,N_18607);
or U24864 (N_24864,N_17548,N_13560);
nor U24865 (N_24865,N_18120,N_15953);
or U24866 (N_24866,N_13649,N_13520);
nand U24867 (N_24867,N_16945,N_14256);
nor U24868 (N_24868,N_16167,N_13544);
nand U24869 (N_24869,N_15168,N_18665);
nand U24870 (N_24870,N_14678,N_16469);
and U24871 (N_24871,N_13484,N_17252);
nor U24872 (N_24872,N_13431,N_14175);
nand U24873 (N_24873,N_13475,N_15365);
or U24874 (N_24874,N_18584,N_15768);
and U24875 (N_24875,N_14526,N_14141);
and U24876 (N_24876,N_13117,N_16221);
or U24877 (N_24877,N_17126,N_15687);
nor U24878 (N_24878,N_15776,N_15920);
or U24879 (N_24879,N_12806,N_18533);
and U24880 (N_24880,N_16986,N_16395);
nor U24881 (N_24881,N_16207,N_13119);
or U24882 (N_24882,N_12686,N_15569);
nand U24883 (N_24883,N_14127,N_14865);
nand U24884 (N_24884,N_16433,N_14286);
or U24885 (N_24885,N_15802,N_17558);
nor U24886 (N_24886,N_16587,N_17159);
or U24887 (N_24887,N_16421,N_14415);
and U24888 (N_24888,N_16705,N_15195);
and U24889 (N_24889,N_13679,N_13332);
nand U24890 (N_24890,N_16960,N_15657);
or U24891 (N_24891,N_18480,N_16010);
nor U24892 (N_24892,N_15536,N_14489);
or U24893 (N_24893,N_14088,N_17819);
and U24894 (N_24894,N_17938,N_14346);
or U24895 (N_24895,N_17808,N_13215);
xnor U24896 (N_24896,N_16044,N_14867);
nor U24897 (N_24897,N_14576,N_14998);
and U24898 (N_24898,N_16581,N_18126);
or U24899 (N_24899,N_15494,N_17842);
nor U24900 (N_24900,N_18633,N_15243);
nor U24901 (N_24901,N_17947,N_17339);
xor U24902 (N_24902,N_18188,N_12822);
nand U24903 (N_24903,N_12533,N_14940);
and U24904 (N_24904,N_18520,N_12909);
nor U24905 (N_24905,N_14029,N_18169);
nand U24906 (N_24906,N_17671,N_13417);
or U24907 (N_24907,N_16044,N_16450);
xor U24908 (N_24908,N_16777,N_14078);
or U24909 (N_24909,N_15002,N_12901);
nand U24910 (N_24910,N_14136,N_16820);
or U24911 (N_24911,N_15536,N_16253);
nor U24912 (N_24912,N_15779,N_13295);
and U24913 (N_24913,N_17817,N_17409);
and U24914 (N_24914,N_14391,N_12526);
or U24915 (N_24915,N_15979,N_16611);
or U24916 (N_24916,N_18514,N_16559);
or U24917 (N_24917,N_14050,N_14892);
nor U24918 (N_24918,N_13741,N_14143);
nand U24919 (N_24919,N_18196,N_15945);
nor U24920 (N_24920,N_13187,N_15692);
and U24921 (N_24921,N_13421,N_13218);
nand U24922 (N_24922,N_16996,N_14995);
or U24923 (N_24923,N_16275,N_12725);
nor U24924 (N_24924,N_16536,N_15972);
or U24925 (N_24925,N_13185,N_16854);
or U24926 (N_24926,N_17970,N_13269);
nand U24927 (N_24927,N_12940,N_16087);
nand U24928 (N_24928,N_17084,N_13977);
or U24929 (N_24929,N_17512,N_15814);
nand U24930 (N_24930,N_13599,N_17862);
nor U24931 (N_24931,N_14128,N_16208);
and U24932 (N_24932,N_18709,N_14373);
or U24933 (N_24933,N_16914,N_14537);
xnor U24934 (N_24934,N_14216,N_17929);
nor U24935 (N_24935,N_13859,N_14390);
nand U24936 (N_24936,N_18461,N_15934);
or U24937 (N_24937,N_14069,N_15354);
and U24938 (N_24938,N_13711,N_17009);
and U24939 (N_24939,N_18572,N_13327);
nand U24940 (N_24940,N_14376,N_13676);
xnor U24941 (N_24941,N_13508,N_12999);
nor U24942 (N_24942,N_17212,N_16472);
or U24943 (N_24943,N_14726,N_18494);
nand U24944 (N_24944,N_13101,N_13380);
nor U24945 (N_24945,N_18727,N_15299);
nand U24946 (N_24946,N_18371,N_17158);
nand U24947 (N_24947,N_14483,N_17041);
nor U24948 (N_24948,N_16015,N_16211);
nand U24949 (N_24949,N_14308,N_17968);
or U24950 (N_24950,N_13022,N_14497);
and U24951 (N_24951,N_14345,N_17616);
or U24952 (N_24952,N_15398,N_16936);
and U24953 (N_24953,N_17374,N_17588);
nor U24954 (N_24954,N_13366,N_15087);
nand U24955 (N_24955,N_17572,N_15016);
nand U24956 (N_24956,N_16501,N_17488);
nor U24957 (N_24957,N_17508,N_14748);
nor U24958 (N_24958,N_13456,N_12564);
nor U24959 (N_24959,N_17664,N_16653);
xor U24960 (N_24960,N_17362,N_13763);
and U24961 (N_24961,N_14302,N_15185);
nor U24962 (N_24962,N_14479,N_18192);
nand U24963 (N_24963,N_14103,N_12763);
or U24964 (N_24964,N_18544,N_17729);
nand U24965 (N_24965,N_18190,N_14282);
or U24966 (N_24966,N_15802,N_13054);
or U24967 (N_24967,N_17108,N_14298);
or U24968 (N_24968,N_13909,N_16570);
and U24969 (N_24969,N_13679,N_17036);
nand U24970 (N_24970,N_15638,N_15964);
and U24971 (N_24971,N_18614,N_18415);
nor U24972 (N_24972,N_17421,N_17162);
or U24973 (N_24973,N_18098,N_16797);
or U24974 (N_24974,N_12986,N_13082);
or U24975 (N_24975,N_17514,N_12500);
nor U24976 (N_24976,N_14011,N_15467);
and U24977 (N_24977,N_16507,N_15429);
nand U24978 (N_24978,N_14190,N_14306);
and U24979 (N_24979,N_18647,N_13055);
nor U24980 (N_24980,N_17562,N_14746);
or U24981 (N_24981,N_14529,N_15089);
or U24982 (N_24982,N_16181,N_16195);
nand U24983 (N_24983,N_17205,N_15237);
or U24984 (N_24984,N_17800,N_13354);
or U24985 (N_24985,N_15246,N_15768);
and U24986 (N_24986,N_18447,N_18296);
nor U24987 (N_24987,N_13345,N_13805);
xor U24988 (N_24988,N_15033,N_15243);
nor U24989 (N_24989,N_16106,N_12709);
nand U24990 (N_24990,N_16269,N_18540);
nor U24991 (N_24991,N_16351,N_17999);
nand U24992 (N_24992,N_14930,N_16200);
or U24993 (N_24993,N_17029,N_12746);
nand U24994 (N_24994,N_18038,N_13683);
nor U24995 (N_24995,N_18376,N_18343);
nand U24996 (N_24996,N_16145,N_16513);
and U24997 (N_24997,N_17393,N_16528);
or U24998 (N_24998,N_12618,N_15709);
or U24999 (N_24999,N_14153,N_18144);
and UO_0 (O_0,N_20528,N_24098);
nand UO_1 (O_1,N_19109,N_21819);
nor UO_2 (O_2,N_21988,N_18750);
nor UO_3 (O_3,N_21298,N_22689);
or UO_4 (O_4,N_20179,N_22001);
nor UO_5 (O_5,N_24428,N_24571);
nor UO_6 (O_6,N_23568,N_22993);
nor UO_7 (O_7,N_20084,N_21323);
or UO_8 (O_8,N_21110,N_22629);
nor UO_9 (O_9,N_21620,N_19511);
nand UO_10 (O_10,N_24598,N_19492);
or UO_11 (O_11,N_20908,N_19522);
or UO_12 (O_12,N_24321,N_23804);
and UO_13 (O_13,N_19456,N_22023);
nor UO_14 (O_14,N_20951,N_24707);
or UO_15 (O_15,N_22029,N_24672);
and UO_16 (O_16,N_20129,N_22936);
or UO_17 (O_17,N_23551,N_20101);
nand UO_18 (O_18,N_22058,N_20656);
or UO_19 (O_19,N_22800,N_20978);
and UO_20 (O_20,N_23164,N_22495);
and UO_21 (O_21,N_24867,N_22753);
nand UO_22 (O_22,N_21136,N_21230);
nor UO_23 (O_23,N_21144,N_20533);
or UO_24 (O_24,N_21077,N_24331);
and UO_25 (O_25,N_21129,N_19494);
nand UO_26 (O_26,N_18939,N_23962);
nand UO_27 (O_27,N_20677,N_22918);
nor UO_28 (O_28,N_22873,N_18827);
and UO_29 (O_29,N_21092,N_20395);
xor UO_30 (O_30,N_21366,N_18821);
and UO_31 (O_31,N_21378,N_20505);
and UO_32 (O_32,N_24775,N_24225);
or UO_33 (O_33,N_22383,N_19729);
or UO_34 (O_34,N_23717,N_22087);
xnor UO_35 (O_35,N_19948,N_24100);
and UO_36 (O_36,N_21722,N_23990);
and UO_37 (O_37,N_23739,N_18925);
or UO_38 (O_38,N_21813,N_21425);
nand UO_39 (O_39,N_24372,N_24697);
xor UO_40 (O_40,N_23214,N_23132);
nand UO_41 (O_41,N_21654,N_24378);
nor UO_42 (O_42,N_23583,N_24963);
nand UO_43 (O_43,N_23511,N_19556);
and UO_44 (O_44,N_23417,N_24642);
nand UO_45 (O_45,N_22210,N_23951);
nand UO_46 (O_46,N_22217,N_19223);
nor UO_47 (O_47,N_23917,N_19629);
nor UO_48 (O_48,N_19785,N_20018);
nand UO_49 (O_49,N_22507,N_20137);
nor UO_50 (O_50,N_18849,N_20565);
and UO_51 (O_51,N_22005,N_24234);
and UO_52 (O_52,N_23737,N_22372);
and UO_53 (O_53,N_24858,N_22461);
or UO_54 (O_54,N_21244,N_21507);
or UO_55 (O_55,N_20948,N_23764);
or UO_56 (O_56,N_21339,N_24316);
or UO_57 (O_57,N_19475,N_24210);
or UO_58 (O_58,N_20039,N_22437);
and UO_59 (O_59,N_20351,N_20864);
nor UO_60 (O_60,N_21325,N_19217);
nor UO_61 (O_61,N_22342,N_23019);
nor UO_62 (O_62,N_21393,N_20597);
or UO_63 (O_63,N_21274,N_21733);
and UO_64 (O_64,N_24186,N_19411);
or UO_65 (O_65,N_20176,N_20110);
and UO_66 (O_66,N_18907,N_19014);
and UO_67 (O_67,N_22769,N_23237);
or UO_68 (O_68,N_19910,N_21334);
and UO_69 (O_69,N_22442,N_22581);
xor UO_70 (O_70,N_23674,N_20027);
and UO_71 (O_71,N_23660,N_19008);
xor UO_72 (O_72,N_18798,N_22790);
and UO_73 (O_73,N_24142,N_21044);
xor UO_74 (O_74,N_20240,N_22482);
and UO_75 (O_75,N_23597,N_24533);
nand UO_76 (O_76,N_20476,N_19968);
or UO_77 (O_77,N_21481,N_19627);
or UO_78 (O_78,N_20836,N_24441);
xnor UO_79 (O_79,N_22156,N_23032);
xor UO_80 (O_80,N_19613,N_24118);
and UO_81 (O_81,N_23817,N_20471);
or UO_82 (O_82,N_24468,N_20235);
or UO_83 (O_83,N_23454,N_24214);
or UO_84 (O_84,N_22522,N_24201);
or UO_85 (O_85,N_24952,N_21256);
and UO_86 (O_86,N_20103,N_24906);
nand UO_87 (O_87,N_24226,N_23490);
nor UO_88 (O_88,N_18890,N_20975);
nand UO_89 (O_89,N_18893,N_20197);
nand UO_90 (O_90,N_22018,N_18788);
nor UO_91 (O_91,N_22424,N_24427);
nand UO_92 (O_92,N_24156,N_19604);
nand UO_93 (O_93,N_21780,N_20093);
or UO_94 (O_94,N_22472,N_22140);
and UO_95 (O_95,N_21952,N_22226);
nor UO_96 (O_96,N_24285,N_21105);
xor UO_97 (O_97,N_24147,N_24423);
nand UO_98 (O_98,N_21829,N_19433);
or UO_99 (O_99,N_21789,N_20209);
and UO_100 (O_100,N_19210,N_23519);
nand UO_101 (O_101,N_24038,N_19835);
nand UO_102 (O_102,N_23964,N_19128);
and UO_103 (O_103,N_23312,N_20270);
or UO_104 (O_104,N_23120,N_21193);
nand UO_105 (O_105,N_18872,N_19010);
nor UO_106 (O_106,N_22544,N_19382);
or UO_107 (O_107,N_22542,N_24259);
nor UO_108 (O_108,N_19147,N_24635);
or UO_109 (O_109,N_21627,N_21709);
nand UO_110 (O_110,N_21958,N_20159);
nor UO_111 (O_111,N_21773,N_20357);
nand UO_112 (O_112,N_20259,N_24604);
or UO_113 (O_113,N_20051,N_22902);
nor UO_114 (O_114,N_22426,N_20319);
or UO_115 (O_115,N_24817,N_24460);
or UO_116 (O_116,N_21540,N_23382);
nand UO_117 (O_117,N_19046,N_22113);
and UO_118 (O_118,N_19247,N_21902);
nand UO_119 (O_119,N_20760,N_20313);
nor UO_120 (O_120,N_23628,N_24405);
nor UO_121 (O_121,N_21943,N_23751);
and UO_122 (O_122,N_20797,N_21258);
and UO_123 (O_123,N_24138,N_21447);
nor UO_124 (O_124,N_23246,N_19236);
nand UO_125 (O_125,N_20717,N_24242);
nand UO_126 (O_126,N_20839,N_22767);
nand UO_127 (O_127,N_24010,N_21974);
xor UO_128 (O_128,N_19279,N_21072);
nor UO_129 (O_129,N_24729,N_19328);
xnor UO_130 (O_130,N_21273,N_20338);
or UO_131 (O_131,N_23325,N_19523);
nand UO_132 (O_132,N_24475,N_22758);
nor UO_133 (O_133,N_20489,N_22419);
xor UO_134 (O_134,N_21957,N_20897);
or UO_135 (O_135,N_19882,N_24905);
nand UO_136 (O_136,N_23997,N_20635);
nand UO_137 (O_137,N_23979,N_24872);
and UO_138 (O_138,N_22157,N_23870);
or UO_139 (O_139,N_21655,N_23153);
and UO_140 (O_140,N_20526,N_23476);
and UO_141 (O_141,N_20355,N_20546);
or UO_142 (O_142,N_24292,N_23556);
nand UO_143 (O_143,N_22407,N_24746);
nand UO_144 (O_144,N_24245,N_22405);
nand UO_145 (O_145,N_24901,N_20377);
nand UO_146 (O_146,N_20178,N_20666);
or UO_147 (O_147,N_21584,N_21309);
nand UO_148 (O_148,N_22571,N_22613);
nor UO_149 (O_149,N_23850,N_22489);
nand UO_150 (O_150,N_24120,N_20363);
nand UO_151 (O_151,N_20157,N_22717);
or UO_152 (O_152,N_22905,N_22840);
nand UO_153 (O_153,N_22933,N_19198);
nand UO_154 (O_154,N_23031,N_20428);
nor UO_155 (O_155,N_22051,N_20906);
or UO_156 (O_156,N_19311,N_22885);
or UO_157 (O_157,N_24713,N_19656);
nor UO_158 (O_158,N_24046,N_22016);
and UO_159 (O_159,N_20964,N_24566);
and UO_160 (O_160,N_19533,N_20070);
nand UO_161 (O_161,N_23912,N_22517);
nor UO_162 (O_162,N_24854,N_21804);
and UO_163 (O_163,N_22180,N_23770);
nand UO_164 (O_164,N_24451,N_22708);
and UO_165 (O_165,N_24273,N_19354);
or UO_166 (O_166,N_21248,N_24485);
or UO_167 (O_167,N_18812,N_24415);
nor UO_168 (O_168,N_24197,N_24094);
nor UO_169 (O_169,N_23387,N_20261);
nand UO_170 (O_170,N_24923,N_24004);
nor UO_171 (O_171,N_23543,N_19645);
and UO_172 (O_172,N_21630,N_21420);
xor UO_173 (O_173,N_24258,N_22651);
or UO_174 (O_174,N_19989,N_22211);
nor UO_175 (O_175,N_24082,N_20433);
and UO_176 (O_176,N_22375,N_22720);
or UO_177 (O_177,N_23500,N_20506);
nor UO_178 (O_178,N_20005,N_24266);
and UO_179 (O_179,N_20558,N_23247);
or UO_180 (O_180,N_20116,N_19049);
and UO_181 (O_181,N_21293,N_24904);
xnor UO_182 (O_182,N_19111,N_24932);
or UO_183 (O_183,N_21717,N_23527);
and UO_184 (O_184,N_22484,N_19712);
or UO_185 (O_185,N_22501,N_22220);
nand UO_186 (O_186,N_21411,N_18958);
nand UO_187 (O_187,N_20837,N_24974);
nand UO_188 (O_188,N_20081,N_24787);
nor UO_189 (O_189,N_22052,N_23895);
nand UO_190 (O_190,N_20435,N_20090);
and UO_191 (O_191,N_21856,N_22197);
xor UO_192 (O_192,N_19927,N_24850);
nand UO_193 (O_193,N_22692,N_24329);
or UO_194 (O_194,N_24852,N_21900);
nand UO_195 (O_195,N_20577,N_19415);
or UO_196 (O_196,N_24101,N_24907);
xnor UO_197 (O_197,N_20622,N_21538);
xor UO_198 (O_198,N_20193,N_24339);
xor UO_199 (O_199,N_22115,N_23687);
nand UO_200 (O_200,N_21923,N_18998);
nand UO_201 (O_201,N_23627,N_20617);
nor UO_202 (O_202,N_19563,N_19956);
and UO_203 (O_203,N_19545,N_21840);
nand UO_204 (O_204,N_24039,N_21180);
and UO_205 (O_205,N_24471,N_23983);
or UO_206 (O_206,N_24174,N_19895);
nand UO_207 (O_207,N_24014,N_20379);
or UO_208 (O_208,N_24778,N_18799);
and UO_209 (O_209,N_22283,N_19634);
xnor UO_210 (O_210,N_24392,N_22703);
nor UO_211 (O_211,N_23505,N_19591);
or UO_212 (O_212,N_21675,N_20352);
or UO_213 (O_213,N_24359,N_20973);
and UO_214 (O_214,N_19325,N_24074);
or UO_215 (O_215,N_21250,N_23212);
nor UO_216 (O_216,N_23923,N_22365);
nor UO_217 (O_217,N_24452,N_22002);
and UO_218 (O_218,N_20469,N_22969);
or UO_219 (O_219,N_19313,N_22027);
or UO_220 (O_220,N_22626,N_21915);
and UO_221 (O_221,N_20960,N_22582);
nor UO_222 (O_222,N_19250,N_23093);
xor UO_223 (O_223,N_19174,N_24883);
and UO_224 (O_224,N_18791,N_23281);
or UO_225 (O_225,N_24232,N_21758);
xor UO_226 (O_226,N_22463,N_24551);
or UO_227 (O_227,N_22543,N_21471);
xor UO_228 (O_228,N_22731,N_22775);
and UO_229 (O_229,N_23196,N_24346);
nor UO_230 (O_230,N_22187,N_19639);
and UO_231 (O_231,N_23774,N_19443);
nand UO_232 (O_232,N_22218,N_21567);
and UO_233 (O_233,N_23516,N_21174);
and UO_234 (O_234,N_18778,N_21009);
nor UO_235 (O_235,N_21604,N_24785);
nand UO_236 (O_236,N_21629,N_21254);
or UO_237 (O_237,N_20241,N_23677);
or UO_238 (O_238,N_22153,N_19098);
nand UO_239 (O_239,N_19536,N_20638);
nor UO_240 (O_240,N_20641,N_19896);
and UO_241 (O_241,N_19142,N_23297);
nor UO_242 (O_242,N_19846,N_21704);
nand UO_243 (O_243,N_20606,N_22768);
and UO_244 (O_244,N_24811,N_21084);
nand UO_245 (O_245,N_22538,N_20397);
and UO_246 (O_246,N_22329,N_21417);
or UO_247 (O_247,N_23190,N_22229);
nand UO_248 (O_248,N_20867,N_21997);
and UO_249 (O_249,N_21187,N_21166);
nor UO_250 (O_250,N_22385,N_24224);
or UO_251 (O_251,N_24588,N_21211);
or UO_252 (O_252,N_18824,N_21795);
nand UO_253 (O_253,N_22341,N_23856);
nor UO_254 (O_254,N_23711,N_24354);
nand UO_255 (O_255,N_19625,N_19268);
nand UO_256 (O_256,N_19954,N_22549);
nand UO_257 (O_257,N_23113,N_20072);
or UO_258 (O_258,N_24334,N_21150);
nor UO_259 (O_259,N_20750,N_20424);
or UO_260 (O_260,N_24721,N_18926);
nor UO_261 (O_261,N_22949,N_21666);
nor UO_262 (O_262,N_19949,N_18963);
nand UO_263 (O_263,N_21463,N_18904);
and UO_264 (O_264,N_20410,N_19466);
nor UO_265 (O_265,N_23054,N_20955);
or UO_266 (O_266,N_21610,N_21590);
and UO_267 (O_267,N_23580,N_20722);
xnor UO_268 (O_268,N_18768,N_21458);
nand UO_269 (O_269,N_23258,N_19992);
or UO_270 (O_270,N_22687,N_23594);
or UO_271 (O_271,N_21059,N_21632);
and UO_272 (O_272,N_22836,N_24646);
and UO_273 (O_273,N_21470,N_19449);
and UO_274 (O_274,N_20822,N_24580);
nand UO_275 (O_275,N_23086,N_19859);
nand UO_276 (O_276,N_21576,N_23986);
xor UO_277 (O_277,N_21993,N_19692);
and UO_278 (O_278,N_19442,N_20670);
or UO_279 (O_279,N_23096,N_21938);
or UO_280 (O_280,N_20277,N_23844);
nand UO_281 (O_281,N_22853,N_19241);
nor UO_282 (O_282,N_22095,N_21455);
nand UO_283 (O_283,N_19737,N_22006);
nor UO_284 (O_284,N_22599,N_21769);
and UO_285 (O_285,N_19769,N_22702);
or UO_286 (O_286,N_22275,N_23940);
and UO_287 (O_287,N_21271,N_18805);
nor UO_288 (O_288,N_24639,N_22718);
nor UO_289 (O_289,N_22286,N_23443);
nand UO_290 (O_290,N_22468,N_21452);
xnor UO_291 (O_291,N_19359,N_23431);
and UO_292 (O_292,N_23754,N_20772);
and UO_293 (O_293,N_19974,N_24215);
nand UO_294 (O_294,N_19810,N_22362);
nand UO_295 (O_295,N_23935,N_23253);
and UO_296 (O_296,N_20658,N_23077);
or UO_297 (O_297,N_19051,N_20782);
nand UO_298 (O_298,N_22530,N_21644);
nand UO_299 (O_299,N_20588,N_22915);
nand UO_300 (O_300,N_23938,N_24200);
or UO_301 (O_301,N_21793,N_24298);
and UO_302 (O_302,N_20390,N_19923);
or UO_303 (O_303,N_23915,N_22805);
and UO_304 (O_304,N_24466,N_24500);
or UO_305 (O_305,N_21219,N_20556);
or UO_306 (O_306,N_20801,N_23016);
or UO_307 (O_307,N_21402,N_22097);
nand UO_308 (O_308,N_20814,N_19681);
nand UO_309 (O_309,N_20762,N_20511);
or UO_310 (O_310,N_20199,N_23503);
xnor UO_311 (O_311,N_20632,N_20102);
and UO_312 (O_312,N_21579,N_24599);
nor UO_313 (O_313,N_22457,N_22883);
or UO_314 (O_314,N_22306,N_19614);
nor UO_315 (O_315,N_19920,N_24047);
nor UO_316 (O_316,N_22627,N_23578);
and UO_317 (O_317,N_19277,N_20162);
or UO_318 (O_318,N_19933,N_19275);
and UO_319 (O_319,N_22054,N_20712);
xnor UO_320 (O_320,N_20296,N_20630);
and UO_321 (O_321,N_20984,N_20727);
and UO_322 (O_322,N_19966,N_18949);
nand UO_323 (O_323,N_20215,N_21689);
nand UO_324 (O_324,N_23814,N_22182);
nand UO_325 (O_325,N_22589,N_21866);
nor UO_326 (O_326,N_19249,N_21825);
nor UO_327 (O_327,N_23868,N_23510);
or UO_328 (O_328,N_22194,N_24706);
and UO_329 (O_329,N_23478,N_22988);
or UO_330 (O_330,N_19716,N_20777);
nand UO_331 (O_331,N_21637,N_23030);
nor UO_332 (O_332,N_19461,N_22019);
or UO_333 (O_333,N_18980,N_20521);
xor UO_334 (O_334,N_20312,N_19877);
nand UO_335 (O_335,N_19999,N_24964);
nand UO_336 (O_336,N_23173,N_23396);
and UO_337 (O_337,N_18990,N_19368);
nor UO_338 (O_338,N_23330,N_19738);
nor UO_339 (O_339,N_24037,N_20965);
nor UO_340 (O_340,N_19588,N_19905);
nor UO_341 (O_341,N_20494,N_20128);
nor UO_342 (O_342,N_21653,N_22535);
and UO_343 (O_343,N_23879,N_23048);
or UO_344 (O_344,N_24132,N_19472);
or UO_345 (O_345,N_22366,N_24476);
nor UO_346 (O_346,N_23522,N_20720);
and UO_347 (O_347,N_21714,N_22200);
nor UO_348 (O_348,N_20966,N_22819);
and UO_349 (O_349,N_23299,N_23474);
nor UO_350 (O_350,N_23352,N_21983);
or UO_351 (O_351,N_22181,N_21748);
or UO_352 (O_352,N_23683,N_20492);
nand UO_353 (O_353,N_22914,N_21034);
or UO_354 (O_354,N_23900,N_21218);
and UO_355 (O_355,N_23833,N_20148);
nor UO_356 (O_356,N_23009,N_23904);
xnor UO_357 (O_357,N_19931,N_24136);
xor UO_358 (O_358,N_21330,N_20592);
and UO_359 (O_359,N_20980,N_24712);
nand UO_360 (O_360,N_20219,N_22455);
nand UO_361 (O_361,N_21349,N_22267);
nand UO_362 (O_362,N_21217,N_20019);
nand UO_363 (O_363,N_24828,N_19139);
or UO_364 (O_364,N_21645,N_22945);
and UO_365 (O_365,N_19932,N_23996);
or UO_366 (O_366,N_19520,N_19836);
and UO_367 (O_367,N_18928,N_22655);
nand UO_368 (O_368,N_19670,N_22374);
nand UO_369 (O_369,N_23262,N_22351);
or UO_370 (O_370,N_23180,N_20725);
xnor UO_371 (O_371,N_24115,N_20675);
nor UO_372 (O_372,N_19900,N_22304);
nand UO_373 (O_373,N_22825,N_23094);
or UO_374 (O_374,N_23818,N_23105);
and UO_375 (O_375,N_21986,N_24893);
nand UO_376 (O_376,N_23139,N_21797);
nor UO_377 (O_377,N_19374,N_23995);
nand UO_378 (O_378,N_21283,N_21888);
and UO_379 (O_379,N_20374,N_22886);
nor UO_380 (O_380,N_22952,N_22765);
nand UO_381 (O_381,N_19011,N_21305);
nand UO_382 (O_382,N_24650,N_22297);
and UO_383 (O_383,N_20429,N_24560);
or UO_384 (O_384,N_24129,N_19326);
nand UO_385 (O_385,N_20171,N_24950);
and UO_386 (O_386,N_23480,N_24430);
nand UO_387 (O_387,N_23198,N_20545);
and UO_388 (O_388,N_21991,N_20316);
or UO_389 (O_389,N_20502,N_23141);
or UO_390 (O_390,N_19087,N_20651);
xnor UO_391 (O_391,N_24124,N_20123);
nand UO_392 (O_392,N_21033,N_23898);
nand UO_393 (O_393,N_19379,N_19420);
and UO_394 (O_394,N_22956,N_19435);
xnor UO_395 (O_395,N_24583,N_23432);
nand UO_396 (O_396,N_21251,N_22307);
nand UO_397 (O_397,N_21560,N_19793);
or UO_398 (O_398,N_20944,N_20117);
nor UO_399 (O_399,N_24634,N_22046);
and UO_400 (O_400,N_19193,N_23462);
or UO_401 (O_401,N_20522,N_18770);
nor UO_402 (O_402,N_21683,N_22563);
nand UO_403 (O_403,N_21635,N_19144);
or UO_404 (O_404,N_23709,N_20647);
nor UO_405 (O_405,N_19784,N_21281);
xor UO_406 (O_406,N_19207,N_19151);
xor UO_407 (O_407,N_23600,N_20213);
or UO_408 (O_408,N_23378,N_18915);
or UO_409 (O_409,N_24790,N_19172);
and UO_410 (O_410,N_21336,N_24264);
or UO_411 (O_411,N_18976,N_21679);
and UO_412 (O_412,N_18996,N_22788);
or UO_413 (O_413,N_20917,N_24664);
nand UO_414 (O_414,N_24554,N_19641);
nor UO_415 (O_415,N_19127,N_19222);
nor UO_416 (O_416,N_20341,N_20284);
and UO_417 (O_417,N_24312,N_24976);
nor UO_418 (O_418,N_20350,N_23082);
nand UO_419 (O_419,N_20267,N_20667);
nand UO_420 (O_420,N_24892,N_19718);
nand UO_421 (O_421,N_22831,N_19584);
nand UO_422 (O_422,N_21743,N_24418);
or UO_423 (O_423,N_24735,N_24962);
nand UO_424 (O_424,N_20495,N_21356);
xnor UO_425 (O_425,N_23045,N_21143);
nor UO_426 (O_426,N_18782,N_19482);
or UO_427 (O_427,N_19367,N_23947);
nor UO_428 (O_428,N_24897,N_22268);
or UO_429 (O_429,N_21864,N_24945);
nor UO_430 (O_430,N_19802,N_23599);
nand UO_431 (O_431,N_22201,N_22178);
or UO_432 (O_432,N_22043,N_19342);
nand UO_433 (O_433,N_20816,N_19348);
nor UO_434 (O_434,N_23468,N_24421);
nand UO_435 (O_435,N_20683,N_21849);
and UO_436 (O_436,N_20943,N_19568);
nor UO_437 (O_437,N_19610,N_21661);
and UO_438 (O_438,N_21133,N_23670);
or UO_439 (O_439,N_20770,N_24806);
nand UO_440 (O_440,N_19636,N_18841);
nand UO_441 (O_441,N_20611,N_19765);
nand UO_442 (O_442,N_23664,N_19547);
or UO_443 (O_443,N_21746,N_24192);
nand UO_444 (O_444,N_21581,N_23361);
nand UO_445 (O_445,N_21301,N_22077);
nor UO_446 (O_446,N_19682,N_23213);
or UO_447 (O_447,N_22179,N_23059);
nor UO_448 (O_448,N_23274,N_22849);
and UO_449 (O_449,N_19617,N_19294);
nand UO_450 (O_450,N_21784,N_24400);
or UO_451 (O_451,N_24462,N_24975);
and UO_452 (O_452,N_19253,N_21000);
nor UO_453 (O_453,N_22161,N_24908);
nor UO_454 (O_454,N_19265,N_21857);
nand UO_455 (O_455,N_18950,N_20470);
nand UO_456 (O_456,N_23326,N_19768);
or UO_457 (O_457,N_18829,N_21592);
and UO_458 (O_458,N_23722,N_22704);
or UO_459 (O_459,N_19271,N_22889);
nor UO_460 (O_460,N_24766,N_24891);
nand UO_461 (O_461,N_19709,N_24877);
xnor UO_462 (O_462,N_20245,N_21222);
nor UO_463 (O_463,N_19830,N_21115);
nor UO_464 (O_464,N_20690,N_19936);
nand UO_465 (O_465,N_20464,N_22408);
xor UO_466 (O_466,N_19478,N_23830);
and UO_467 (O_467,N_20515,N_20210);
nand UO_468 (O_468,N_21541,N_21762);
nand UO_469 (O_469,N_24618,N_20281);
nand UO_470 (O_470,N_20280,N_24957);
nor UO_471 (O_471,N_24845,N_24969);
nor UO_472 (O_472,N_21613,N_24573);
nor UO_473 (O_473,N_24154,N_20188);
xnor UO_474 (O_474,N_22661,N_21240);
and UO_475 (O_475,N_23292,N_24515);
xor UO_476 (O_476,N_21961,N_19499);
nor UO_477 (O_477,N_19660,N_21944);
and UO_478 (O_478,N_23100,N_21729);
nor UO_479 (O_479,N_24608,N_24060);
and UO_480 (O_480,N_24102,N_19609);
and UO_481 (O_481,N_23867,N_22590);
or UO_482 (O_482,N_23542,N_18945);
nand UO_483 (O_483,N_23199,N_21459);
xor UO_484 (O_484,N_21288,N_21977);
xnor UO_485 (O_485,N_20878,N_21872);
xor UO_486 (O_486,N_20961,N_24875);
nor UO_487 (O_487,N_21842,N_19928);
or UO_488 (O_488,N_20499,N_23554);
xor UO_489 (O_489,N_20979,N_24472);
and UO_490 (O_490,N_20255,N_23347);
and UO_491 (O_491,N_22036,N_21435);
nand UO_492 (O_492,N_20330,N_22621);
nor UO_493 (O_493,N_21817,N_22233);
nand UO_494 (O_494,N_21060,N_24925);
or UO_495 (O_495,N_23821,N_20924);
and UO_496 (O_496,N_19592,N_19881);
or UO_497 (O_497,N_20449,N_24196);
and UO_498 (O_498,N_19848,N_22376);
nor UO_499 (O_499,N_22913,N_20548);
or UO_500 (O_500,N_23678,N_21778);
or UO_501 (O_501,N_21368,N_23486);
nor UO_502 (O_502,N_22884,N_23760);
and UO_503 (O_503,N_21238,N_22101);
and UO_504 (O_504,N_24457,N_21224);
or UO_505 (O_505,N_22526,N_21677);
or UO_506 (O_506,N_22724,N_20151);
nand UO_507 (O_507,N_23875,N_19616);
nand UO_508 (O_508,N_19377,N_21557);
nor UO_509 (O_509,N_21533,N_22057);
nand UO_510 (O_510,N_20028,N_19904);
and UO_511 (O_511,N_20655,N_22235);
or UO_512 (O_512,N_18809,N_19912);
and UO_513 (O_513,N_23092,N_19230);
nand UO_514 (O_514,N_23943,N_23106);
nand UO_515 (O_515,N_24390,N_23634);
or UO_516 (O_516,N_22996,N_19873);
nor UO_517 (O_517,N_19403,N_18792);
nor UO_518 (O_518,N_23571,N_20400);
and UO_519 (O_519,N_22262,N_19080);
nand UO_520 (O_520,N_21725,N_21934);
xor UO_521 (O_521,N_24403,N_18923);
or UO_522 (O_522,N_23216,N_24253);
nor UO_523 (O_523,N_20305,N_22428);
nand UO_524 (O_524,N_24998,N_22158);
nor UO_525 (O_525,N_22285,N_21351);
or UO_526 (O_526,N_24203,N_21354);
or UO_527 (O_527,N_20068,N_23968);
or UO_528 (O_528,N_19842,N_20477);
nor UO_529 (O_529,N_21467,N_19345);
xor UO_530 (O_530,N_23147,N_19378);
nor UO_531 (O_531,N_18956,N_20855);
and UO_532 (O_532,N_24365,N_21488);
and UO_533 (O_533,N_21882,N_24960);
or UO_534 (O_534,N_20404,N_23372);
nand UO_535 (O_535,N_23411,N_21408);
nor UO_536 (O_536,N_23383,N_19680);
and UO_537 (O_537,N_19451,N_23589);
nor UO_538 (O_538,N_21652,N_21041);
nor UO_539 (O_539,N_20744,N_24789);
nand UO_540 (O_540,N_20756,N_24172);
nand UO_541 (O_541,N_20608,N_19474);
or UO_542 (O_542,N_22470,N_20554);
xnor UO_543 (O_543,N_21523,N_20012);
nor UO_544 (O_544,N_23593,N_24161);
or UO_545 (O_545,N_20015,N_20799);
xor UO_546 (O_546,N_22104,N_19788);
nand UO_547 (O_547,N_21727,N_19984);
nand UO_548 (O_548,N_22425,N_20161);
or UO_549 (O_549,N_19107,N_24984);
xnor UO_550 (O_550,N_22799,N_22771);
nor UO_551 (O_551,N_20835,N_24473);
and UO_552 (O_552,N_19512,N_23303);
or UO_553 (O_553,N_23663,N_24271);
and UO_554 (O_554,N_22536,N_19229);
nor UO_555 (O_555,N_20002,N_22208);
nand UO_556 (O_556,N_22995,N_24399);
nor UO_557 (O_557,N_20881,N_23977);
or UO_558 (O_558,N_21770,N_22524);
nor UO_559 (O_559,N_23076,N_24183);
or UO_560 (O_560,N_19383,N_23766);
nor UO_561 (O_561,N_20249,N_20687);
nor UO_562 (O_562,N_19668,N_22477);
and UO_563 (O_563,N_23430,N_19962);
or UO_564 (O_564,N_20856,N_19957);
nor UO_565 (O_565,N_22516,N_19622);
nor UO_566 (O_566,N_21113,N_21345);
or UO_567 (O_567,N_19458,N_22764);
xor UO_568 (O_568,N_19820,N_23366);
nand UO_569 (O_569,N_20517,N_22594);
and UO_570 (O_570,N_23323,N_24176);
and UO_571 (O_571,N_22481,N_22124);
and UO_572 (O_572,N_22322,N_23063);
or UO_573 (O_573,N_20576,N_21448);
nor UO_574 (O_574,N_20686,N_21303);
nor UO_575 (O_575,N_23643,N_21569);
and UO_576 (O_576,N_21834,N_24249);
and UO_577 (O_577,N_20551,N_19524);
nor UO_578 (O_578,N_24239,N_20500);
nor UO_579 (O_579,N_24188,N_21577);
and UO_580 (O_580,N_21011,N_23479);
nor UO_581 (O_581,N_19364,N_20463);
nor UO_582 (O_582,N_24376,N_23718);
nor UO_583 (O_583,N_20992,N_23103);
nor UO_584 (O_584,N_20009,N_18816);
and UO_585 (O_585,N_19187,N_22637);
nor UO_586 (O_586,N_21236,N_21416);
xor UO_587 (O_587,N_19647,N_18762);
and UO_588 (O_588,N_22712,N_20033);
and UO_589 (O_589,N_24968,N_20870);
nand UO_590 (O_590,N_19502,N_22628);
or UO_591 (O_591,N_20125,N_24871);
or UO_592 (O_592,N_23874,N_19292);
or UO_593 (O_593,N_24576,N_24042);
nand UO_594 (O_594,N_22438,N_18804);
and UO_595 (O_595,N_24866,N_24080);
or UO_596 (O_596,N_22830,N_22392);
and UO_597 (O_597,N_22142,N_23062);
or UO_598 (O_598,N_24035,N_22160);
xor UO_599 (O_599,N_22204,N_23209);
or UO_600 (O_600,N_22337,N_19689);
xor UO_601 (O_601,N_22984,N_21255);
nor UO_602 (O_602,N_19837,N_21572);
xor UO_603 (O_603,N_24282,N_24869);
or UO_604 (O_604,N_23371,N_20396);
nand UO_605 (O_605,N_22387,N_24049);
nand UO_606 (O_606,N_21525,N_24611);
nor UO_607 (O_607,N_19710,N_20890);
and UO_608 (O_608,N_18819,N_21980);
and UO_609 (O_609,N_18790,N_20386);
nand UO_610 (O_610,N_22977,N_20322);
nand UO_611 (O_611,N_19398,N_18847);
nand UO_612 (O_612,N_20573,N_23458);
or UO_613 (O_613,N_24636,N_24758);
xnor UO_614 (O_614,N_21949,N_20347);
nor UO_615 (O_615,N_22975,N_22386);
or UO_616 (O_616,N_19394,N_20328);
nand UO_617 (O_617,N_22154,N_24517);
nor UO_618 (O_618,N_20361,N_23654);
and UO_619 (O_619,N_23743,N_19597);
or UO_620 (O_620,N_21814,N_19704);
nand UO_621 (O_621,N_19037,N_19714);
and UO_622 (O_622,N_22904,N_19698);
or UO_623 (O_623,N_19365,N_20803);
or UO_624 (O_624,N_19486,N_24570);
nand UO_625 (O_625,N_21464,N_22658);
nand UO_626 (O_626,N_23883,N_23226);
nor UO_627 (O_627,N_24884,N_18814);
or UO_628 (O_628,N_21671,N_18869);
and UO_629 (O_629,N_21445,N_20336);
nand UO_630 (O_630,N_21845,N_18826);
nand UO_631 (O_631,N_24288,N_22280);
xnor UO_632 (O_632,N_22305,N_19436);
nor UO_633 (O_633,N_21877,N_20854);
and UO_634 (O_634,N_23261,N_24375);
or UO_635 (O_635,N_22967,N_19314);
and UO_636 (O_636,N_18978,N_21879);
nor UO_637 (O_637,N_24480,N_23146);
nand UO_638 (O_638,N_24007,N_18981);
nor UO_639 (O_639,N_18766,N_20938);
or UO_640 (O_640,N_20244,N_19498);
and UO_641 (O_641,N_23370,N_23823);
or UO_642 (O_642,N_22301,N_24043);
or UO_643 (O_643,N_23957,N_23338);
or UO_644 (O_644,N_19238,N_23428);
and UO_645 (O_645,N_20740,N_24678);
and UO_646 (O_646,N_19947,N_24396);
and UO_647 (O_647,N_24052,N_19686);
nor UO_648 (O_648,N_20531,N_23350);
and UO_649 (O_649,N_22887,N_22130);
nand UO_650 (O_650,N_20454,N_19291);
and UO_651 (O_651,N_22748,N_22697);
nand UO_652 (O_652,N_19876,N_23099);
nand UO_653 (O_653,N_19891,N_20668);
nor UO_654 (O_654,N_20031,N_19262);
nor UO_655 (O_655,N_20243,N_24304);
or UO_656 (O_656,N_24028,N_22102);
and UO_657 (O_657,N_24767,N_22378);
nand UO_658 (O_658,N_24296,N_22611);
and UO_659 (O_659,N_19796,N_22107);
or UO_660 (O_660,N_19826,N_23949);
nor UO_661 (O_661,N_22569,N_24607);
or UO_662 (O_662,N_24416,N_24406);
and UO_663 (O_663,N_19535,N_22309);
and UO_664 (O_664,N_23914,N_20536);
nor UO_665 (O_665,N_19684,N_19462);
and UO_666 (O_666,N_19118,N_22228);
or UO_667 (O_667,N_23606,N_19340);
xor UO_668 (O_668,N_19245,N_23410);
and UO_669 (O_669,N_23267,N_22614);
and UO_670 (O_670,N_20607,N_24336);
or UO_671 (O_671,N_21532,N_22827);
or UO_672 (O_672,N_20331,N_21156);
and UO_673 (O_673,N_22175,N_19117);
or UO_674 (O_674,N_24177,N_24720);
xnor UO_675 (O_675,N_22694,N_21479);
or UO_676 (O_676,N_20602,N_19105);
nand UO_677 (O_677,N_23565,N_22333);
nand UO_678 (O_678,N_20865,N_20614);
nor UO_679 (O_679,N_23026,N_23893);
and UO_680 (O_680,N_21973,N_19880);
xnor UO_681 (O_681,N_23269,N_21205);
or UO_682 (O_682,N_24303,N_24005);
and UO_683 (O_683,N_19421,N_23994);
nand UO_684 (O_684,N_24584,N_24013);
or UO_685 (O_685,N_24738,N_22931);
and UO_686 (O_686,N_20950,N_20247);
nor UO_687 (O_687,N_21322,N_24095);
or UO_688 (O_688,N_20307,N_24841);
nand UO_689 (O_689,N_19950,N_22238);
and UO_690 (O_690,N_20513,N_19542);
and UO_691 (O_691,N_19958,N_21706);
xnor UO_692 (O_692,N_23742,N_20061);
xor UO_693 (O_693,N_24328,N_19565);
nor UO_694 (O_694,N_19648,N_24637);
nor UO_695 (O_695,N_24483,N_19606);
nor UO_696 (O_696,N_22777,N_22796);
nand UO_697 (O_697,N_19997,N_23456);
or UO_698 (O_698,N_19150,N_19149);
nand UO_699 (O_699,N_23197,N_20566);
xnor UO_700 (O_700,N_19446,N_19336);
nand UO_701 (O_701,N_23037,N_23793);
or UO_702 (O_702,N_23934,N_19518);
or UO_703 (O_703,N_19863,N_20315);
xnor UO_704 (O_704,N_18918,N_22837);
xnor UO_705 (O_705,N_21487,N_20375);
and UO_706 (O_706,N_21003,N_19575);
or UO_707 (O_707,N_21894,N_21418);
or UO_708 (O_708,N_24807,N_22413);
or UO_709 (O_709,N_22266,N_21966);
xnor UO_710 (O_710,N_22642,N_23924);
and UO_711 (O_711,N_20143,N_19805);
nand UO_712 (O_712,N_22440,N_19349);
and UO_713 (O_713,N_24626,N_21233);
or UO_714 (O_714,N_18962,N_20729);
nor UO_715 (O_715,N_20300,N_21215);
or UO_716 (O_716,N_22741,N_23203);
or UO_717 (O_717,N_22039,N_20055);
and UO_718 (O_718,N_22462,N_22259);
xnor UO_719 (O_719,N_20971,N_24824);
nor UO_720 (O_720,N_21633,N_18897);
nand UO_721 (O_721,N_24338,N_23002);
or UO_722 (O_722,N_19308,N_21761);
nand UO_723 (O_723,N_23158,N_22649);
or UO_724 (O_724,N_19943,N_21615);
nand UO_725 (O_725,N_19633,N_24189);
or UO_726 (O_726,N_23688,N_21895);
or UO_727 (O_727,N_21951,N_24695);
and UO_728 (O_728,N_20618,N_19607);
nand UO_729 (O_729,N_21766,N_19827);
nor UO_730 (O_730,N_21266,N_23332);
and UO_731 (O_731,N_19600,N_24740);
and UO_732 (O_732,N_19334,N_21809);
or UO_733 (O_733,N_22331,N_24838);
xor UO_734 (O_734,N_19497,N_18917);
nand UO_735 (O_735,N_21792,N_21710);
nor UO_736 (O_736,N_19567,N_22959);
xor UO_737 (O_737,N_21659,N_20832);
or UO_738 (O_738,N_24973,N_22049);
nand UO_739 (O_739,N_22033,N_21663);
nor UO_740 (O_740,N_24477,N_18946);
xor UO_741 (O_741,N_20399,N_24941);
and UO_742 (O_742,N_22150,N_18794);
nor UO_743 (O_743,N_22723,N_21674);
nand UO_744 (O_744,N_24757,N_23950);
nor UO_745 (O_745,N_24278,N_22469);
and UO_746 (O_746,N_19792,N_22384);
and UO_747 (O_747,N_20807,N_24502);
nand UO_748 (O_748,N_24055,N_21209);
and UO_749 (O_749,N_21494,N_21558);
and UO_750 (O_750,N_19199,N_18931);
nand UO_751 (O_751,N_23319,N_24204);
nand UO_752 (O_752,N_19677,N_20022);
nor UO_753 (O_753,N_22615,N_20298);
and UO_754 (O_754,N_23367,N_18943);
nor UO_755 (O_755,N_21607,N_18851);
nand UO_756 (O_756,N_18898,N_21695);
nor UO_757 (O_757,N_24107,N_20701);
nand UO_758 (O_758,N_22693,N_24062);
nand UO_759 (O_759,N_19231,N_18781);
and UO_760 (O_760,N_24936,N_23576);
or UO_761 (O_761,N_19386,N_18825);
and UO_762 (O_762,N_19893,N_23148);
and UO_763 (O_763,N_19832,N_22512);
or UO_764 (O_764,N_19173,N_19527);
or UO_765 (O_765,N_20892,N_21697);
nor UO_766 (O_766,N_24725,N_20177);
or UO_767 (O_767,N_19194,N_19740);
or UO_768 (O_768,N_24104,N_24185);
nor UO_769 (O_769,N_22165,N_23324);
and UO_770 (O_770,N_23901,N_20831);
and UO_771 (O_771,N_21718,N_20574);
nand UO_772 (O_772,N_22804,N_23541);
nand UO_773 (O_773,N_19828,N_23284);
or UO_774 (O_774,N_22088,N_21984);
or UO_775 (O_775,N_23257,N_22382);
and UO_776 (O_776,N_21053,N_24800);
xor UO_777 (O_777,N_22193,N_23730);
or UO_778 (O_778,N_19990,N_22456);
nor UO_779 (O_779,N_24317,N_23925);
nand UO_780 (O_780,N_22937,N_19307);
nor UO_781 (O_781,N_21061,N_24810);
and UO_782 (O_782,N_20840,N_24315);
nor UO_783 (O_783,N_22292,N_19120);
nand UO_784 (O_784,N_22066,N_23178);
and UO_785 (O_785,N_23976,N_23909);
and UO_786 (O_786,N_23162,N_20082);
nor UO_787 (O_787,N_21898,N_21277);
nand UO_788 (O_788,N_21002,N_19746);
nor UO_789 (O_789,N_21624,N_18861);
nand UO_790 (O_790,N_21332,N_19175);
nor UO_791 (O_791,N_21911,N_20437);
nor UO_792 (O_792,N_21182,N_24981);
or UO_793 (O_793,N_22505,N_19883);
nor UO_794 (O_794,N_22816,N_23613);
nand UO_795 (O_795,N_22675,N_23467);
or UO_796 (O_796,N_23716,N_21955);
nor UO_797 (O_797,N_23321,N_20644);
and UO_798 (O_798,N_20590,N_21646);
nand UO_799 (O_799,N_23958,N_23888);
and UO_800 (O_800,N_19515,N_22155);
xor UO_801 (O_801,N_22448,N_23574);
nor UO_802 (O_802,N_20853,N_23789);
and UO_803 (O_803,N_21519,N_24613);
or UO_804 (O_804,N_19021,N_20032);
or UO_805 (O_805,N_24822,N_22899);
and UO_806 (O_806,N_18758,N_19059);
nor UO_807 (O_807,N_19060,N_20422);
xnor UO_808 (O_808,N_24744,N_23618);
and UO_809 (O_809,N_22953,N_22325);
nand UO_810 (O_810,N_24956,N_23605);
or UO_811 (O_811,N_20568,N_22747);
nand UO_812 (O_812,N_19296,N_22295);
or UO_813 (O_813,N_20194,N_19531);
nor UO_814 (O_814,N_24847,N_19082);
and UO_815 (O_815,N_21948,N_22011);
and UO_816 (O_816,N_20990,N_19352);
xnor UO_817 (O_817,N_19347,N_22416);
nor UO_818 (O_818,N_22490,N_24763);
and UO_819 (O_819,N_23217,N_23587);
nor UO_820 (O_820,N_20182,N_22263);
and UO_821 (O_821,N_21127,N_21880);
nor UO_822 (O_822,N_21412,N_24325);
nor UO_823 (O_823,N_22906,N_21771);
xnor UO_824 (O_824,N_24493,N_20127);
nand UO_825 (O_825,N_23822,N_20848);
xor UO_826 (O_826,N_20077,N_20583);
or UO_827 (O_827,N_18883,N_24750);
nand UO_828 (O_828,N_24680,N_23886);
nor UO_829 (O_829,N_22667,N_21422);
nand UO_830 (O_830,N_19985,N_22688);
nand UO_831 (O_831,N_23160,N_23154);
xnor UO_832 (O_832,N_23005,N_21153);
and UO_833 (O_833,N_21424,N_20265);
or UO_834 (O_834,N_24277,N_20473);
nand UO_835 (O_835,N_18909,N_22149);
xor UO_836 (O_836,N_18818,N_23193);
or UO_837 (O_837,N_21039,N_22300);
nor UO_838 (O_838,N_22186,N_22811);
or UO_839 (O_839,N_24887,N_19350);
or UO_840 (O_840,N_19412,N_23757);
or UO_841 (O_841,N_20595,N_20349);
or UO_842 (O_842,N_20451,N_19743);
nor UO_843 (O_843,N_20098,N_21014);
nand UO_844 (O_844,N_18902,N_23307);
nand UO_845 (O_845,N_24970,N_19766);
nand UO_846 (O_846,N_23225,N_20444);
nor UO_847 (O_847,N_19373,N_24402);
nor UO_848 (O_848,N_24935,N_24110);
nand UO_849 (O_849,N_20017,N_23369);
xor UO_850 (O_850,N_24447,N_19829);
or UO_851 (O_851,N_22531,N_21589);
or UO_852 (O_852,N_19935,N_24267);
or UO_853 (O_853,N_24550,N_22147);
nor UO_854 (O_854,N_24422,N_23465);
nor UO_855 (O_855,N_23992,N_21862);
nor UO_856 (O_856,N_19281,N_18927);
nor UO_857 (O_857,N_20327,N_21314);
nor UO_858 (O_858,N_20343,N_24227);
or UO_859 (O_859,N_20652,N_23966);
xor UO_860 (O_860,N_23930,N_24532);
or UO_861 (O_861,N_20947,N_20126);
nor UO_862 (O_862,N_20509,N_20879);
nor UO_863 (O_863,N_23521,N_19131);
and UO_864 (O_864,N_19753,N_20752);
nor UO_865 (O_865,N_18880,N_24381);
nor UO_866 (O_866,N_20735,N_21469);
xor UO_867 (O_867,N_22047,N_22880);
nor UO_868 (O_868,N_19384,N_24445);
and UO_869 (O_869,N_19981,N_19919);
nand UO_870 (O_870,N_19137,N_22562);
nor UO_871 (O_871,N_21386,N_24190);
or UO_872 (O_872,N_20672,N_23128);
nand UO_873 (O_873,N_19095,N_24048);
or UO_874 (O_874,N_22042,N_24131);
nand UO_875 (O_875,N_20158,N_19263);
nand UO_876 (O_876,N_23713,N_19665);
and UO_877 (O_877,N_24353,N_18891);
and UO_878 (O_878,N_21138,N_18752);
nor UO_879 (O_879,N_24498,N_22460);
nand UO_880 (O_880,N_23546,N_23745);
and UO_881 (O_881,N_19408,N_24689);
and UO_882 (O_882,N_23720,N_19288);
or UO_883 (O_883,N_22103,N_22578);
or UO_884 (O_884,N_19503,N_21295);
or UO_885 (O_885,N_21234,N_24512);
and UO_886 (O_886,N_24965,N_23945);
and UO_887 (O_887,N_21313,N_24289);
and UO_888 (O_888,N_24463,N_18922);
and UO_889 (O_889,N_21350,N_22809);
nand UO_890 (O_890,N_22532,N_19067);
nor UO_891 (O_891,N_23499,N_24439);
and UO_892 (O_892,N_18901,N_20728);
and UO_893 (O_893,N_21601,N_21715);
or UO_894 (O_894,N_20639,N_23941);
nand UO_895 (O_895,N_24793,N_23008);
or UO_896 (O_896,N_24876,N_20414);
nand UO_897 (O_897,N_23386,N_20180);
or UO_898 (O_898,N_19177,N_19221);
and UO_899 (O_899,N_22145,N_20730);
and UO_900 (O_900,N_22466,N_21148);
nand UO_901 (O_901,N_21937,N_19521);
and UO_902 (O_902,N_24572,N_19867);
nor UO_903 (O_903,N_24917,N_20604);
nor UO_904 (O_904,N_21331,N_22326);
nor UO_905 (O_905,N_18942,N_21050);
nand UO_906 (O_906,N_22606,N_24307);
nor UO_907 (O_907,N_23315,N_19064);
nand UO_908 (O_908,N_21520,N_21865);
nor UO_909 (O_909,N_23134,N_24099);
and UO_910 (O_910,N_20282,N_22017);
nand UO_911 (O_911,N_19537,N_24078);
nor UO_912 (O_912,N_21466,N_22414);
nand UO_913 (O_913,N_21787,N_24330);
and UO_914 (O_914,N_19180,N_19539);
and UO_915 (O_915,N_24765,N_19298);
and UO_916 (O_916,N_20800,N_24986);
nor UO_917 (O_917,N_24061,N_23022);
nor UO_918 (O_918,N_23459,N_24276);
nor UO_919 (O_919,N_19023,N_23359);
and UO_920 (O_920,N_24603,N_21565);
nor UO_921 (O_921,N_24090,N_22350);
nor UO_922 (O_922,N_23637,N_19110);
or UO_923 (O_923,N_24844,N_22068);
or UO_924 (O_924,N_19017,N_22698);
and UO_925 (O_925,N_24309,N_24546);
nand UO_926 (O_926,N_19959,N_21383);
or UO_927 (O_927,N_19721,N_22979);
nand UO_928 (O_928,N_23288,N_18896);
nor UO_929 (O_929,N_19982,N_20834);
and UO_930 (O_930,N_22854,N_23775);
and UO_931 (O_931,N_20860,N_21312);
nor UO_932 (O_932,N_23487,N_21324);
nor UO_933 (O_933,N_24362,N_24579);
and UO_934 (O_934,N_21286,N_18779);
or UO_935 (O_935,N_20323,N_22605);
and UO_936 (O_936,N_20207,N_18879);
or UO_937 (O_937,N_23518,N_19644);
and UO_938 (O_938,N_21527,N_22409);
nand UO_939 (O_939,N_20121,N_24444);
or UO_940 (O_940,N_23653,N_23699);
nor UO_941 (O_941,N_22985,N_20203);
and UO_942 (O_942,N_21165,N_20381);
and UO_943 (O_943,N_24531,N_20187);
and UO_944 (O_944,N_21736,N_20220);
nand UO_945 (O_945,N_20609,N_22746);
nor UO_946 (O_946,N_23890,N_23065);
and UO_947 (O_947,N_19302,N_21836);
and UO_948 (O_948,N_20657,N_24541);
or UO_949 (O_949,N_22779,N_20996);
nand UO_950 (O_950,N_19058,N_20589);
and UO_951 (O_951,N_24256,N_24130);
or UO_952 (O_952,N_22665,N_22992);
xor UO_953 (O_953,N_22498,N_21502);
nand UO_954 (O_954,N_22349,N_19429);
nor UO_955 (O_955,N_22445,N_19165);
or UO_956 (O_956,N_19921,N_22290);
and UO_957 (O_957,N_24220,N_24503);
and UO_958 (O_958,N_18803,N_22841);
nor UO_959 (O_959,N_20578,N_20224);
xnor UO_960 (O_960,N_22683,N_24692);
and UO_961 (O_961,N_21178,N_23693);
and UO_962 (O_962,N_22454,N_22393);
nor UO_963 (O_963,N_24640,N_22946);
nor UO_964 (O_964,N_21381,N_19577);
and UO_965 (O_965,N_19084,N_22221);
nand UO_966 (O_966,N_20529,N_21423);
nand UO_967 (O_967,N_23413,N_23873);
and UO_968 (O_968,N_24333,N_21892);
or UO_969 (O_969,N_20096,N_19838);
or UO_970 (O_970,N_22877,N_21344);
and UO_971 (O_971,N_23696,N_19141);
nand UO_972 (O_972,N_23007,N_21184);
or UO_973 (O_973,N_23528,N_24357);
nand UO_974 (O_974,N_19467,N_24609);
and UO_975 (O_975,N_21800,N_24233);
or UO_976 (O_976,N_24861,N_20935);
nor UO_977 (O_977,N_23283,N_19282);
or UO_978 (O_978,N_20314,N_20535);
nor UO_979 (O_979,N_21055,N_18914);
nor UO_980 (O_980,N_22846,N_19169);
nand UO_981 (O_981,N_20631,N_24212);
and UO_982 (O_982,N_19004,N_20508);
nor UO_983 (O_983,N_20047,N_23090);
xor UO_984 (O_984,N_19944,N_23922);
nor UO_985 (O_985,N_24464,N_19413);
and UO_986 (O_986,N_19728,N_19079);
nand UO_987 (O_987,N_22040,N_24388);
or UO_988 (O_988,N_20789,N_23374);
nor UO_989 (O_989,N_23234,N_21082);
nand UO_990 (O_990,N_23506,N_23609);
nand UO_991 (O_991,N_22663,N_19203);
xor UO_992 (O_992,N_20173,N_24855);
nand UO_993 (O_993,N_19602,N_23919);
and UO_994 (O_994,N_20001,N_22900);
nand UO_995 (O_995,N_21711,N_18846);
nor UO_996 (O_996,N_21020,N_20929);
or UO_997 (O_997,N_20423,N_20997);
and UO_998 (O_998,N_24761,N_22183);
nor UO_999 (O_999,N_23552,N_20468);
and UO_1000 (O_1000,N_21774,N_19605);
or UO_1001 (O_1001,N_24363,N_22310);
and UO_1002 (O_1002,N_20046,N_19126);
xor UO_1003 (O_1003,N_24287,N_24469);
xnor UO_1004 (O_1004,N_23039,N_19078);
nor UO_1005 (O_1005,N_20903,N_21320);
nor UO_1006 (O_1006,N_21401,N_20185);
nand UO_1007 (O_1007,N_22974,N_21702);
and UO_1008 (O_1008,N_22941,N_20024);
nor UO_1009 (O_1009,N_21669,N_20060);
nor UO_1010 (O_1010,N_20448,N_24219);
nand UO_1011 (O_1011,N_24459,N_23024);
and UO_1012 (O_1012,N_23238,N_23166);
or UO_1013 (O_1013,N_23156,N_23525);
and UO_1014 (O_1014,N_20273,N_20886);
or UO_1015 (O_1015,N_22989,N_19991);
nor UO_1016 (O_1016,N_19564,N_23135);
and UO_1017 (O_1017,N_22978,N_24139);
nand UO_1018 (O_1018,N_19154,N_21811);
nor UO_1019 (O_1019,N_18913,N_23972);
or UO_1020 (O_1020,N_21641,N_23066);
and UO_1021 (O_1021,N_24308,N_19794);
or UO_1022 (O_1022,N_19164,N_23665);
or UO_1023 (O_1023,N_20516,N_21563);
and UO_1024 (O_1024,N_19745,N_22381);
xor UO_1025 (O_1025,N_21530,N_22955);
nand UO_1026 (O_1026,N_22935,N_24567);
nand UO_1027 (O_1027,N_19234,N_23707);
nor UO_1028 (O_1028,N_20914,N_22099);
nor UO_1029 (O_1029,N_22302,N_20438);
and UO_1030 (O_1030,N_21071,N_24041);
nand UO_1031 (O_1031,N_22856,N_19155);
or UO_1032 (O_1032,N_24864,N_20056);
nor UO_1033 (O_1033,N_18754,N_21206);
nand UO_1034 (O_1034,N_21098,N_19642);
xor UO_1035 (O_1035,N_21756,N_19857);
nand UO_1036 (O_1036,N_21022,N_22789);
nand UO_1037 (O_1037,N_19161,N_21728);
or UO_1038 (O_1038,N_20326,N_20716);
xor UO_1039 (O_1039,N_21434,N_19760);
nor UO_1040 (O_1040,N_20896,N_18985);
xor UO_1041 (O_1041,N_23001,N_24319);
nor UO_1042 (O_1042,N_22389,N_19732);
nand UO_1043 (O_1043,N_20420,N_21228);
nand UO_1044 (O_1044,N_22670,N_22176);
nand UO_1045 (O_1045,N_21651,N_22592);
or UO_1046 (O_1046,N_20324,N_20006);
and UO_1047 (O_1047,N_23548,N_22745);
xnor UO_1048 (O_1048,N_22868,N_24073);
or UO_1049 (O_1049,N_23177,N_20804);
nor UO_1050 (O_1050,N_20926,N_19970);
nor UO_1051 (O_1051,N_19752,N_20000);
or UO_1052 (O_1052,N_22277,N_21611);
or UO_1053 (O_1053,N_19918,N_18970);
nor UO_1054 (O_1054,N_23905,N_22420);
and UO_1055 (O_1055,N_23884,N_22855);
nor UO_1056 (O_1056,N_21798,N_20353);
nor UO_1057 (O_1057,N_20385,N_20105);
nor UO_1058 (O_1058,N_20190,N_23682);
or UO_1059 (O_1059,N_22948,N_23956);
and UO_1060 (O_1060,N_22539,N_22196);
nor UO_1061 (O_1061,N_22546,N_23863);
nand UO_1062 (O_1062,N_21642,N_24324);
nor UO_1063 (O_1063,N_23851,N_19332);
and UO_1064 (O_1064,N_23866,N_21738);
nor UO_1065 (O_1065,N_22232,N_21846);
and UO_1066 (O_1066,N_23960,N_19346);
or UO_1067 (O_1067,N_19685,N_18789);
nand UO_1068 (O_1068,N_19585,N_20539);
or UO_1069 (O_1069,N_20628,N_20785);
nand UO_1070 (O_1070,N_23591,N_20332);
nand UO_1071 (O_1071,N_22499,N_19940);
nand UO_1072 (O_1072,N_23205,N_24732);
xor UO_1073 (O_1073,N_21476,N_23470);
nand UO_1074 (O_1074,N_24175,N_23107);
nand UO_1075 (O_1075,N_18845,N_19581);
or UO_1076 (O_1076,N_19967,N_24122);
and UO_1077 (O_1077,N_24167,N_20297);
nor UO_1078 (O_1078,N_21496,N_21149);
or UO_1079 (O_1079,N_19700,N_18764);
and UO_1080 (O_1080,N_19650,N_19507);
and UO_1081 (O_1081,N_18777,N_23971);
and UO_1082 (O_1082,N_23186,N_22994);
xor UO_1083 (O_1083,N_22063,N_24837);
or UO_1084 (O_1084,N_19994,N_24257);
nand UO_1085 (O_1085,N_24492,N_24829);
xnor UO_1086 (O_1086,N_24377,N_19840);
nor UO_1087 (O_1087,N_21026,N_22822);
or UO_1088 (O_1088,N_21667,N_18759);
xnor UO_1089 (O_1089,N_24369,N_18870);
or UO_1090 (O_1090,N_21907,N_20100);
nand UO_1091 (O_1091,N_20139,N_20251);
nand UO_1092 (O_1092,N_20764,N_24023);
nor UO_1093 (O_1093,N_19573,N_23590);
or UO_1094 (O_1094,N_22380,N_21981);
nor UO_1095 (O_1095,N_21310,N_22358);
nor UO_1096 (O_1096,N_22835,N_22639);
xor UO_1097 (O_1097,N_21382,N_19476);
and UO_1098 (O_1098,N_23439,N_20694);
nand UO_1099 (O_1099,N_20598,N_24556);
nand UO_1100 (O_1100,N_24745,N_21985);
or UO_1101 (O_1101,N_18989,N_18934);
nand UO_1102 (O_1102,N_23630,N_20078);
xnor UO_1103 (O_1103,N_23782,N_23690);
nand UO_1104 (O_1104,N_19817,N_23349);
and UO_1105 (O_1105,N_24280,N_19038);
nor UO_1106 (O_1106,N_22079,N_19321);
nand UO_1107 (O_1107,N_19274,N_18857);
and UO_1108 (O_1108,N_24163,N_22510);
and UO_1109 (O_1109,N_23507,N_20174);
and UO_1110 (O_1110,N_23604,N_21586);
nand UO_1111 (O_1111,N_24108,N_19351);
or UO_1112 (O_1112,N_23429,N_23512);
or UO_1113 (O_1113,N_24591,N_19258);
xor UO_1114 (O_1114,N_20048,N_24739);
xnor UO_1115 (O_1115,N_24195,N_23978);
nand UO_1116 (O_1116,N_22399,N_19303);
nand UO_1117 (O_1117,N_23881,N_24146);
xnor UO_1118 (O_1118,N_23820,N_20877);
or UO_1119 (O_1119,N_24805,N_24719);
or UO_1120 (O_1120,N_20678,N_23662);
nand UO_1121 (O_1121,N_21707,N_22299);
and UO_1122 (O_1122,N_24535,N_19306);
nor UO_1123 (O_1123,N_24568,N_23526);
nor UO_1124 (O_1124,N_21259,N_23187);
nand UO_1125 (O_1125,N_24857,N_24592);
xnor UO_1126 (O_1126,N_24170,N_22603);
or UO_1127 (O_1127,N_21384,N_22369);
nand UO_1128 (O_1128,N_23981,N_23734);
or UO_1129 (O_1129,N_20311,N_21186);
nor UO_1130 (O_1130,N_22537,N_19615);
and UO_1131 (O_1131,N_22534,N_20474);
nor UO_1132 (O_1132,N_24865,N_20387);
and UO_1133 (O_1133,N_23143,N_19691);
nand UO_1134 (O_1134,N_20680,N_21429);
and UO_1135 (O_1135,N_20767,N_22207);
nand UO_1136 (O_1136,N_19034,N_22736);
nand UO_1137 (O_1137,N_24987,N_21587);
nand UO_1138 (O_1138,N_21299,N_22276);
or UO_1139 (O_1139,N_24915,N_20862);
nand UO_1140 (O_1140,N_22737,N_20858);
xor UO_1141 (O_1141,N_21906,N_23118);
xor UO_1142 (O_1142,N_23698,N_19062);
or UO_1143 (O_1143,N_18813,N_24628);
nand UO_1144 (O_1144,N_24539,N_21554);
or UO_1145 (O_1145,N_19490,N_21696);
and UO_1146 (O_1146,N_22987,N_19094);
or UO_1147 (O_1147,N_23876,N_22164);
nor UO_1148 (O_1148,N_22070,N_21874);
or UO_1149 (O_1149,N_22269,N_18852);
nand UO_1150 (O_1150,N_19260,N_22441);
and UO_1151 (O_1151,N_20654,N_21426);
or UO_1152 (O_1152,N_20932,N_23249);
nor UO_1153 (O_1153,N_21886,N_21767);
xnor UO_1154 (O_1154,N_24386,N_22942);
nor UO_1155 (O_1155,N_22826,N_22360);
nor UO_1156 (O_1156,N_21861,N_22635);
nor UO_1157 (O_1157,N_22355,N_21117);
nor UO_1158 (O_1158,N_23471,N_24809);
nand UO_1159 (O_1159,N_23270,N_24490);
or UO_1160 (O_1160,N_22806,N_24614);
nand UO_1161 (O_1161,N_22272,N_21164);
and UO_1162 (O_1162,N_22735,N_24653);
or UO_1163 (O_1163,N_20356,N_22230);
nor UO_1164 (O_1164,N_20755,N_21431);
xor UO_1165 (O_1165,N_24702,N_19839);
nand UO_1166 (O_1166,N_20525,N_20401);
and UO_1167 (O_1167,N_22726,N_23227);
or UO_1168 (O_1168,N_23948,N_19643);
nor UO_1169 (O_1169,N_19240,N_18850);
nor UO_1170 (O_1170,N_24083,N_22520);
and UO_1171 (O_1171,N_24479,N_20898);
nand UO_1172 (O_1172,N_19445,N_20023);
or UO_1173 (O_1173,N_23502,N_20620);
and UO_1174 (O_1174,N_24294,N_20748);
and UO_1175 (O_1175,N_23491,N_21111);
xor UO_1176 (O_1176,N_20993,N_20792);
nor UO_1177 (O_1177,N_23404,N_22890);
and UO_1178 (O_1178,N_24971,N_19108);
nand UO_1179 (O_1179,N_22169,N_18979);
xor UO_1180 (O_1180,N_24522,N_19439);
or UO_1181 (O_1181,N_22427,N_24559);
and UO_1182 (O_1182,N_22552,N_21070);
and UO_1183 (O_1183,N_21147,N_19965);
nor UO_1184 (O_1184,N_20587,N_20671);
nand UO_1185 (O_1185,N_22215,N_22185);
nand UO_1186 (O_1186,N_24616,N_22999);
xnor UO_1187 (O_1187,N_21449,N_21231);
xnor UO_1188 (O_1188,N_22254,N_22247);
nor UO_1189 (O_1189,N_24569,N_23836);
and UO_1190 (O_1190,N_21747,N_19619);
nand UO_1191 (O_1191,N_19256,N_20114);
or UO_1192 (O_1192,N_24863,N_20780);
or UO_1193 (O_1193,N_22513,N_21173);
and UO_1194 (O_1194,N_23140,N_19596);
nor UO_1195 (O_1195,N_21462,N_23582);
nor UO_1196 (O_1196,N_21123,N_20043);
nand UO_1197 (O_1197,N_21032,N_19875);
nand UO_1198 (O_1198,N_18910,N_24240);
and UO_1199 (O_1199,N_23791,N_22696);
or UO_1200 (O_1200,N_19834,N_24769);
and UO_1201 (O_1201,N_24951,N_22734);
nor UO_1202 (O_1202,N_22901,N_22450);
xnor UO_1203 (O_1203,N_20378,N_23612);
nor UO_1204 (O_1204,N_18973,N_19952);
and UO_1205 (O_1205,N_21755,N_24030);
nand UO_1206 (O_1206,N_21608,N_22722);
or UO_1207 (O_1207,N_19808,N_22315);
and UO_1208 (O_1208,N_19658,N_18971);
xnor UO_1209 (O_1209,N_21873,N_20884);
nand UO_1210 (O_1210,N_19076,N_24839);
nand UO_1211 (O_1211,N_24379,N_22264);
nand UO_1212 (O_1212,N_20811,N_20812);
or UO_1213 (O_1213,N_22545,N_18892);
nor UO_1214 (O_1214,N_21260,N_24283);
nor UO_1215 (O_1215,N_18780,N_23602);
nand UO_1216 (O_1216,N_24458,N_20817);
nand UO_1217 (O_1217,N_19724,N_19595);
and UO_1218 (O_1218,N_24275,N_21982);
and UO_1219 (O_1219,N_22069,N_20673);
nor UO_1220 (O_1220,N_22727,N_19006);
nand UO_1221 (O_1221,N_20646,N_20768);
xor UO_1222 (O_1222,N_24340,N_23955);
and UO_1223 (O_1223,N_20821,N_22246);
nor UO_1224 (O_1224,N_24989,N_23539);
or UO_1225 (O_1225,N_19986,N_19072);
and UO_1226 (O_1226,N_18796,N_23072);
xnor UO_1227 (O_1227,N_22607,N_19434);
and UO_1228 (O_1228,N_22007,N_22523);
or UO_1229 (O_1229,N_20124,N_18855);
xor UO_1230 (O_1230,N_19042,N_19483);
and UO_1231 (O_1231,N_22620,N_22561);
nand UO_1232 (O_1232,N_21506,N_21788);
xnor UO_1233 (O_1233,N_22625,N_21045);
or UO_1234 (O_1234,N_21764,N_24424);
or UO_1235 (O_1235,N_20237,N_23295);
nor UO_1236 (O_1236,N_21457,N_24751);
and UO_1237 (O_1237,N_22676,N_20702);
or UO_1238 (O_1238,N_19179,N_22998);
nor UO_1239 (O_1239,N_22814,N_24155);
nor UO_1240 (O_1240,N_20563,N_19695);
nand UO_1241 (O_1241,N_24297,N_18835);
nand UO_1242 (O_1242,N_21621,N_21617);
and UO_1243 (O_1243,N_24772,N_19343);
or UO_1244 (O_1244,N_21501,N_22679);
nor UO_1245 (O_1245,N_20108,N_19338);
xor UO_1246 (O_1246,N_20236,N_22298);
and UO_1247 (O_1247,N_21392,N_23125);
or UO_1248 (O_1248,N_19868,N_22258);
xor UO_1249 (O_1249,N_23616,N_18930);
nor UO_1250 (O_1250,N_21037,N_24698);
and UO_1251 (O_1251,N_24373,N_21177);
xnor UO_1252 (O_1252,N_18806,N_20044);
or UO_1253 (O_1253,N_19166,N_24181);
nand UO_1254 (O_1254,N_23078,N_23741);
and UO_1255 (O_1255,N_18984,N_20283);
xor UO_1256 (O_1256,N_19866,N_19376);
nand UO_1257 (O_1257,N_19027,N_21614);
and UO_1258 (O_1258,N_22109,N_20407);
nand UO_1259 (O_1259,N_22636,N_22110);
nor UO_1260 (O_1260,N_18769,N_21939);
xnor UO_1261 (O_1261,N_19419,N_20714);
xor UO_1262 (O_1262,N_21801,N_19951);
nor UO_1263 (O_1263,N_19455,N_20514);
xnor UO_1264 (O_1264,N_20596,N_24849);
xnor UO_1265 (O_1265,N_24794,N_23569);
nor UO_1266 (O_1266,N_20802,N_19869);
and UO_1267 (O_1267,N_23381,N_19942);
nor UO_1268 (O_1268,N_22346,N_23412);
or UO_1269 (O_1269,N_19676,N_24437);
nor UO_1270 (O_1270,N_20488,N_20291);
nand UO_1271 (O_1271,N_24658,N_22601);
xor UO_1272 (O_1272,N_23807,N_19742);
nor UO_1273 (O_1273,N_24620,N_23728);
and UO_1274 (O_1274,N_21552,N_23219);
or UO_1275 (O_1275,N_21600,N_21088);
nand UO_1276 (O_1276,N_21509,N_23027);
nand UO_1277 (O_1277,N_24450,N_21419);
nand UO_1278 (O_1278,N_24773,N_21514);
and UO_1279 (O_1279,N_22766,N_20164);
nand UO_1280 (O_1280,N_23746,N_22080);
or UO_1281 (O_1281,N_24545,N_21460);
nor UO_1282 (O_1282,N_20254,N_20537);
or UO_1283 (O_1283,N_22398,N_24578);
or UO_1284 (O_1284,N_22014,N_23980);
or UO_1285 (O_1285,N_20527,N_20181);
nand UO_1286 (O_1286,N_24641,N_18834);
and UO_1287 (O_1287,N_18854,N_18757);
xnor UO_1288 (O_1288,N_24433,N_21896);
nand UO_1289 (O_1289,N_24438,N_23254);
nor UO_1290 (O_1290,N_19319,N_19115);
and UO_1291 (O_1291,N_22293,N_24831);
and UO_1292 (O_1292,N_23138,N_24250);
or UO_1293 (O_1293,N_19312,N_19257);
nand UO_1294 (O_1294,N_19337,N_21075);
or UO_1295 (O_1295,N_21720,N_22423);
nand UO_1296 (O_1296,N_19504,N_24979);
nand UO_1297 (O_1297,N_19558,N_19135);
nand UO_1298 (O_1298,N_23691,N_19460);
or UO_1299 (O_1299,N_21357,N_18840);
nand UO_1300 (O_1300,N_22136,N_21210);
nor UO_1301 (O_1301,N_21490,N_21678);
and UO_1302 (O_1302,N_20593,N_20869);
nand UO_1303 (O_1303,N_22202,N_19106);
nor UO_1304 (O_1304,N_20798,N_24456);
nand UO_1305 (O_1305,N_20569,N_21759);
or UO_1306 (O_1306,N_23038,N_23149);
or UO_1307 (O_1307,N_23829,N_22981);
or UO_1308 (O_1308,N_21242,N_19039);
xnor UO_1309 (O_1309,N_22662,N_20806);
nor UO_1310 (O_1310,N_24305,N_22528);
and UO_1311 (O_1311,N_20119,N_21932);
nand UO_1312 (O_1312,N_20930,N_19329);
or UO_1313 (O_1313,N_21086,N_19033);
and UO_1314 (O_1314,N_23131,N_23018);
nand UO_1315 (O_1315,N_24704,N_21216);
nor UO_1316 (O_1316,N_22114,N_23397);
nand UO_1317 (O_1317,N_20662,N_23860);
nand UO_1318 (O_1318,N_22744,N_21820);
or UO_1319 (O_1319,N_21772,N_23137);
nor UO_1320 (O_1320,N_24663,N_19874);
nand UO_1321 (O_1321,N_22072,N_22654);
or UO_1322 (O_1322,N_20663,N_20403);
or UO_1323 (O_1323,N_21183,N_24085);
nand UO_1324 (O_1324,N_19781,N_24953);
nand UO_1325 (O_1325,N_20510,N_23017);
or UO_1326 (O_1326,N_23339,N_24434);
nand UO_1327 (O_1327,N_20676,N_19651);
nor UO_1328 (O_1328,N_20786,N_24961);
nor UO_1329 (O_1329,N_24449,N_22131);
xor UO_1330 (O_1330,N_23706,N_23749);
nor UO_1331 (O_1331,N_19315,N_23335);
or UO_1332 (O_1332,N_20995,N_21158);
or UO_1333 (O_1333,N_24966,N_23765);
nor UO_1334 (O_1334,N_24878,N_22558);
and UO_1335 (O_1335,N_23161,N_21684);
nor UO_1336 (O_1336,N_22755,N_24027);
or UO_1337 (O_1337,N_19430,N_21292);
nor UO_1338 (O_1338,N_21482,N_19657);
or UO_1339 (O_1339,N_23055,N_22397);
or UO_1340 (O_1340,N_20773,N_21142);
or UO_1341 (O_1341,N_23658,N_22340);
nor UO_1342 (O_1342,N_21151,N_19213);
xor UO_1343 (O_1343,N_23788,N_19018);
and UO_1344 (O_1344,N_24255,N_23684);
nand UO_1345 (O_1345,N_24284,N_20827);
and UO_1346 (O_1346,N_19623,N_22927);
and UO_1347 (O_1347,N_20693,N_21638);
nor UO_1348 (O_1348,N_21371,N_20586);
and UO_1349 (O_1349,N_20025,N_21421);
nand UO_1350 (O_1350,N_23639,N_21130);
nor UO_1351 (O_1351,N_23864,N_23920);
nand UO_1352 (O_1352,N_18975,N_20561);
nor UO_1353 (O_1353,N_20383,N_22458);
nand UO_1354 (O_1354,N_24109,N_24216);
nor UO_1355 (O_1355,N_19410,N_19783);
nor UO_1356 (O_1356,N_21047,N_21574);
nor UO_1357 (O_1357,N_20112,N_22818);
and UO_1358 (O_1358,N_23296,N_23398);
nand UO_1359 (O_1359,N_23114,N_24919);
nand UO_1360 (O_1360,N_19701,N_21226);
and UO_1361 (O_1361,N_24978,N_22801);
xor UO_1362 (O_1362,N_22851,N_21107);
nor UO_1363 (O_1363,N_21844,N_24260);
nor UO_1364 (O_1364,N_22056,N_21257);
or UO_1365 (O_1365,N_21941,N_19181);
nor UO_1366 (O_1366,N_20842,N_20062);
and UO_1367 (O_1367,N_23501,N_20907);
nand UO_1368 (O_1368,N_21734,N_23337);
or UO_1369 (O_1369,N_18972,N_24235);
and UO_1370 (O_1370,N_23123,N_22912);
xnor UO_1371 (O_1371,N_23598,N_23418);
nand UO_1372 (O_1372,N_20705,N_20572);
or UO_1373 (O_1373,N_19370,N_23360);
nor UO_1374 (O_1374,N_21400,N_24587);
nand UO_1375 (O_1375,N_19450,N_23845);
or UO_1376 (O_1376,N_21785,N_24696);
and UO_1377 (O_1377,N_18884,N_19395);
nor UO_1378 (O_1378,N_22443,N_20726);
or UO_1379 (O_1379,N_19441,N_20260);
nor UO_1380 (O_1380,N_20682,N_21369);
xnor UO_1381 (O_1381,N_23640,N_22911);
or UO_1382 (O_1382,N_18924,N_24018);
or UO_1383 (O_1383,N_19540,N_22009);
nand UO_1384 (O_1384,N_20624,N_21212);
and UO_1385 (O_1385,N_21304,N_24318);
and UO_1386 (O_1386,N_19821,N_23259);
nand UO_1387 (O_1387,N_24868,N_19590);
and UO_1388 (O_1388,N_23786,N_23340);
or UO_1389 (O_1389,N_24633,N_24446);
and UO_1390 (O_1390,N_23222,N_20757);
nor UO_1391 (O_1391,N_23824,N_20696);
nand UO_1392 (O_1392,N_22112,N_23172);
nand UO_1393 (O_1393,N_23029,N_22893);
nand UO_1394 (O_1394,N_19103,N_21647);
or UO_1395 (O_1395,N_21917,N_23515);
nand UO_1396 (O_1396,N_24705,N_19550);
nand UO_1397 (O_1397,N_22844,N_23825);
nor UO_1398 (O_1398,N_20418,N_23080);
or UO_1399 (O_1399,N_24853,N_24916);
or UO_1400 (O_1400,N_19849,N_21081);
and UO_1401 (O_1401,N_19833,N_20703);
and UO_1402 (O_1402,N_24801,N_24407);
nand UO_1403 (O_1403,N_24977,N_20458);
and UO_1404 (O_1404,N_19133,N_20645);
and UO_1405 (O_1405,N_22584,N_21112);
xnor UO_1406 (O_1406,N_18920,N_22842);
nor UO_1407 (O_1407,N_24946,N_19086);
or UO_1408 (O_1408,N_19454,N_21595);
and UO_1409 (O_1409,N_23896,N_21536);
or UO_1410 (O_1410,N_20795,N_22700);
xnor UO_1411 (O_1411,N_24749,N_23641);
or UO_1412 (O_1412,N_20949,N_20099);
or UO_1413 (O_1413,N_23837,N_21703);
nand UO_1414 (O_1414,N_22451,N_21916);
nor UO_1415 (O_1415,N_19286,N_23619);
or UO_1416 (O_1416,N_24796,N_20409);
nand UO_1417 (O_1417,N_18995,N_23549);
nand UO_1418 (O_1418,N_23617,N_19693);
xnor UO_1419 (O_1419,N_20954,N_20783);
nand UO_1420 (O_1420,N_20183,N_19929);
nand UO_1421 (O_1421,N_23129,N_23268);
nand UO_1422 (O_1422,N_24677,N_20934);
and UO_1423 (O_1423,N_24327,N_23014);
xnor UO_1424 (O_1424,N_21097,N_20184);
nor UO_1425 (O_1425,N_23241,N_20707);
nor UO_1426 (O_1426,N_21499,N_19671);
and UO_1427 (O_1427,N_21201,N_20562);
or UO_1428 (O_1428,N_19853,N_24371);
and UO_1429 (O_1429,N_19100,N_20138);
xnor UO_1430 (O_1430,N_24669,N_23363);
nand UO_1431 (O_1431,N_21656,N_21352);
or UO_1432 (O_1432,N_21279,N_20079);
nand UO_1433 (O_1433,N_18787,N_23621);
and UO_1434 (O_1434,N_24619,N_24223);
nand UO_1435 (O_1435,N_19063,N_23097);
nor UO_1436 (O_1436,N_20758,N_22467);
or UO_1437 (O_1437,N_22205,N_22249);
nor UO_1438 (O_1438,N_20968,N_23838);
or UO_1439 (O_1439,N_22432,N_23320);
nand UO_1440 (O_1440,N_20321,N_21340);
or UO_1441 (O_1441,N_23533,N_20111);
or UO_1442 (O_1442,N_23704,N_19649);
and UO_1443 (O_1443,N_23392,N_24565);
nand UO_1444 (O_1444,N_22646,N_20946);
nand UO_1445 (O_1445,N_19603,N_23406);
and UO_1446 (O_1446,N_23840,N_20432);
nand UO_1447 (O_1447,N_19293,N_20459);
and UO_1448 (O_1448,N_21394,N_22435);
nand UO_1449 (O_1449,N_21282,N_22038);
xor UO_1450 (O_1450,N_20749,N_19731);
xnor UO_1451 (O_1451,N_19735,N_23811);
or UO_1452 (O_1452,N_24488,N_20491);
and UO_1453 (O_1453,N_24105,N_23603);
xnor UO_1454 (O_1454,N_22222,N_19831);
and UO_1455 (O_1455,N_24389,N_23006);
nand UO_1456 (O_1456,N_23069,N_19757);
and UO_1457 (O_1457,N_19469,N_18888);
xor UO_1458 (O_1458,N_20442,N_24690);
xor UO_1459 (O_1459,N_19136,N_21294);
nand UO_1460 (O_1460,N_20957,N_22035);
and UO_1461 (O_1461,N_20075,N_22572);
or UO_1462 (O_1462,N_20358,N_21493);
or UO_1463 (O_1463,N_24934,N_22476);
xnor UO_1464 (O_1464,N_24632,N_24000);
and UO_1465 (O_1465,N_20922,N_22903);
and UO_1466 (O_1466,N_24836,N_24741);
or UO_1467 (O_1467,N_19500,N_23021);
nand UO_1468 (O_1468,N_20279,N_22919);
nor UO_1469 (O_1469,N_19116,N_21511);
or UO_1470 (O_1470,N_19206,N_21739);
or UO_1471 (O_1471,N_23409,N_20104);
nand UO_1472 (O_1472,N_22503,N_21548);
nor UO_1473 (O_1473,N_20091,N_19586);
or UO_1474 (O_1474,N_22129,N_23189);
nand UO_1475 (O_1475,N_23991,N_24151);
or UO_1476 (O_1476,N_23828,N_19516);
and UO_1477 (O_1477,N_23278,N_18969);
or UO_1478 (O_1478,N_22859,N_20895);
nor UO_1479 (O_1479,N_20512,N_21194);
and UO_1480 (O_1480,N_24349,N_21508);
xnor UO_1481 (O_1481,N_24675,N_21040);
and UO_1482 (O_1482,N_24021,N_24771);
nor UO_1483 (O_1483,N_19572,N_22506);
nand UO_1484 (O_1484,N_20195,N_22486);
or UO_1485 (O_1485,N_24681,N_24499);
xor UO_1486 (O_1486,N_21492,N_24024);
xnor UO_1487 (O_1487,N_23799,N_22116);
nand UO_1488 (O_1488,N_22950,N_18988);
and UO_1489 (O_1489,N_24383,N_22195);
and UO_1490 (O_1490,N_20719,N_20486);
or UO_1491 (O_1491,N_22074,N_19055);
and UO_1492 (O_1492,N_19162,N_21253);
or UO_1493 (O_1493,N_22970,N_20582);
xor UO_1494 (O_1494,N_24506,N_21118);
nor UO_1495 (O_1495,N_19397,N_24059);
nand UO_1496 (O_1496,N_23290,N_18982);
nor UO_1497 (O_1497,N_18774,N_19316);
nor UO_1498 (O_1498,N_19153,N_19361);
and UO_1499 (O_1499,N_24091,N_21327);
or UO_1500 (O_1500,N_20376,N_23744);
or UO_1501 (O_1501,N_22583,N_23738);
or UO_1502 (O_1502,N_23885,N_21454);
nand UO_1503 (O_1503,N_19385,N_20170);
nand UO_1504 (O_1504,N_24113,N_24848);
nand UO_1505 (O_1505,N_23608,N_20542);
nor UO_1506 (O_1506,N_23601,N_23041);
nand UO_1507 (O_1507,N_21940,N_21609);
and UO_1508 (O_1508,N_22320,N_24217);
and UO_1509 (O_1509,N_18954,N_19513);
nand UO_1510 (O_1510,N_24056,N_22808);
nand UO_1511 (O_1511,N_20269,N_22845);
nand UO_1512 (O_1512,N_22664,N_21757);
xor UO_1513 (O_1513,N_22706,N_22402);
and UO_1514 (O_1514,N_20708,N_22431);
nor UO_1515 (O_1515,N_24688,N_24299);
or UO_1516 (O_1516,N_19661,N_21261);
and UO_1517 (O_1517,N_23859,N_21765);
and UO_1518 (O_1518,N_21284,N_20909);
and UO_1519 (O_1519,N_24926,N_23144);
nand UO_1520 (O_1520,N_21329,N_19114);
or UO_1521 (O_1521,N_20570,N_19580);
nand UO_1522 (O_1522,N_22519,N_21619);
nand UO_1523 (O_1523,N_21321,N_22244);
nand UO_1524 (O_1524,N_22652,N_23921);
and UO_1525 (O_1525,N_20796,N_19797);
and UO_1526 (O_1526,N_23083,N_24182);
or UO_1527 (O_1527,N_21791,N_19734);
nor UO_1528 (O_1528,N_19758,N_23540);
or UO_1529 (O_1529,N_24279,N_24443);
or UO_1530 (O_1530,N_24135,N_20753);
nand UO_1531 (O_1531,N_20156,N_21694);
xor UO_1532 (O_1532,N_22715,N_19123);
xnor UO_1533 (O_1533,N_22446,N_19779);
and UO_1534 (O_1534,N_19749,N_23869);
and UO_1535 (O_1535,N_18968,N_21119);
nor UO_1536 (O_1536,N_19777,N_19005);
xor UO_1537 (O_1537,N_22106,N_22478);
or UO_1538 (O_1538,N_24631,N_21837);
xnor UO_1539 (O_1539,N_22371,N_19819);
nand UO_1540 (O_1540,N_23455,N_21054);
and UO_1541 (O_1541,N_24676,N_22647);
nand UO_1542 (O_1542,N_21338,N_20292);
nor UO_1543 (O_1543,N_23620,N_22772);
and UO_1544 (O_1544,N_23133,N_23661);
nand UO_1545 (O_1545,N_19678,N_18765);
or UO_1546 (O_1546,N_23343,N_20905);
nor UO_1547 (O_1547,N_21875,N_19917);
nor UO_1548 (O_1548,N_21987,N_19775);
or UO_1549 (O_1549,N_24519,N_24655);
nand UO_1550 (O_1550,N_22281,N_23889);
or UO_1551 (O_1551,N_21237,N_20918);
nor UO_1552 (O_1552,N_23656,N_21512);
or UO_1553 (O_1553,N_23776,N_22279);
nand UO_1554 (O_1554,N_24207,N_21893);
nor UO_1555 (O_1555,N_24070,N_22225);
nor UO_1556 (O_1556,N_22990,N_20035);
nor UO_1557 (O_1557,N_24621,N_20212);
nor UO_1558 (O_1558,N_21959,N_24589);
or UO_1559 (O_1559,N_23579,N_20605);
or UO_1560 (O_1560,N_23091,N_19344);
nor UO_1561 (O_1561,N_20257,N_22958);
nand UO_1562 (O_1562,N_23056,N_23806);
nor UO_1563 (O_1563,N_24454,N_21539);
xor UO_1564 (O_1564,N_23903,N_20010);
and UO_1565 (O_1565,N_24367,N_21017);
or UO_1566 (O_1566,N_23136,N_23607);
nand UO_1567 (O_1567,N_20230,N_20828);
xor UO_1568 (O_1568,N_22618,N_24344);
nor UO_1569 (O_1569,N_19428,N_19003);
and UO_1570 (O_1570,N_24542,N_19969);
xor UO_1571 (O_1571,N_23365,N_24687);
or UO_1572 (O_1572,N_23402,N_21625);
xor UO_1573 (O_1573,N_23880,N_23424);
and UO_1574 (O_1574,N_24518,N_18830);
or UO_1575 (O_1575,N_19019,N_19251);
xor UO_1576 (O_1576,N_23260,N_23794);
nand UO_1577 (O_1577,N_21036,N_24899);
nand UO_1578 (O_1578,N_23702,N_24051);
xnor UO_1579 (O_1579,N_21498,N_23555);
nor UO_1580 (O_1580,N_19897,N_19447);
and UO_1581 (O_1581,N_19736,N_19519);
nand UO_1582 (O_1582,N_21316,N_22216);
nor UO_1583 (O_1583,N_21198,N_21404);
nand UO_1584 (O_1584,N_19574,N_21134);
xnor UO_1585 (O_1585,N_24075,N_20766);
nor UO_1586 (O_1586,N_19192,N_20097);
nand UO_1587 (O_1587,N_22270,N_20642);
nand UO_1588 (O_1588,N_19372,N_19560);
nor UO_1589 (O_1589,N_22415,N_24411);
nor UO_1590 (O_1590,N_24202,N_24679);
nand UO_1591 (O_1591,N_21227,N_23795);
or UO_1592 (O_1592,N_23484,N_20389);
and UO_1593 (O_1593,N_22751,N_19012);
nor UO_1594 (O_1594,N_24602,N_19669);
or UO_1595 (O_1595,N_21179,N_21947);
nand UO_1596 (O_1596,N_23625,N_20880);
and UO_1597 (O_1597,N_21716,N_22166);
nand UO_1598 (O_1598,N_20490,N_19002);
and UO_1599 (O_1599,N_24461,N_18878);
xor UO_1600 (O_1600,N_20440,N_21942);
and UO_1601 (O_1601,N_21073,N_22608);
or UO_1602 (O_1602,N_21751,N_22824);
or UO_1603 (O_1603,N_19976,N_19485);
and UO_1604 (O_1604,N_24764,N_23116);
or UO_1605 (O_1605,N_20692,N_20074);
nand UO_1606 (O_1606,N_19888,N_20591);
or UO_1607 (O_1607,N_19800,N_23070);
xor UO_1608 (O_1608,N_23553,N_23623);
nor UO_1609 (O_1609,N_19284,N_22963);
nand UO_1610 (O_1610,N_23483,N_24881);
nand UO_1611 (O_1611,N_24314,N_20889);
or UO_1612 (O_1612,N_21928,N_21247);
and UO_1613 (O_1613,N_22634,N_21395);
and UO_1614 (O_1614,N_21839,N_19029);
nor UO_1615 (O_1615,N_23287,N_21007);
and UO_1616 (O_1616,N_19487,N_21171);
or UO_1617 (O_1617,N_22593,N_22896);
and UO_1618 (O_1618,N_20461,N_23251);
nor UO_1619 (O_1619,N_21542,N_21963);
nor UO_1620 (O_1620,N_21950,N_24173);
or UO_1621 (O_1621,N_22630,N_22598);
or UO_1622 (O_1622,N_22865,N_20008);
nor UO_1623 (O_1623,N_24709,N_24191);
nor UO_1624 (O_1624,N_22274,N_21145);
nor UO_1625 (O_1625,N_19914,N_23040);
or UO_1626 (O_1626,N_23179,N_20398);
and UO_1627 (O_1627,N_19851,N_21409);
nor UO_1628 (O_1628,N_19327,N_19824);
or UO_1629 (O_1629,N_20923,N_20434);
nor UO_1630 (O_1630,N_22316,N_21899);
xor UO_1631 (O_1631,N_20419,N_20094);
nor UO_1632 (O_1632,N_21491,N_22078);
and UO_1633 (O_1633,N_21478,N_20092);
nand UO_1634 (O_1634,N_24335,N_23858);
or UO_1635 (O_1635,N_22504,N_20784);
nand UO_1636 (O_1636,N_21367,N_24409);
and UO_1637 (O_1637,N_20226,N_19501);
xor UO_1638 (O_1638,N_19856,N_23003);
nor UO_1639 (O_1639,N_20710,N_23207);
and UO_1640 (O_1640,N_20846,N_23473);
and UO_1641 (O_1641,N_18775,N_21891);
xor UO_1642 (O_1642,N_21370,N_20928);
and UO_1643 (O_1643,N_24726,N_23545);
nand UO_1644 (O_1644,N_22502,N_24322);
nor UO_1645 (O_1645,N_24753,N_23289);
or UO_1646 (O_1646,N_24320,N_18948);
or UO_1647 (O_1647,N_21526,N_21505);
xnor UO_1648 (O_1648,N_23117,N_20931);
nor UO_1649 (O_1649,N_24718,N_21657);
nor UO_1650 (O_1650,N_24586,N_23067);
nor UO_1651 (O_1651,N_21048,N_20134);
and UO_1652 (O_1652,N_21239,N_23802);
nand UO_1653 (O_1653,N_19582,N_24003);
xnor UO_1654 (O_1654,N_19683,N_23482);
nor UO_1655 (O_1655,N_21779,N_19228);
or UO_1656 (O_1656,N_24011,N_22240);
nor UO_1657 (O_1657,N_20135,N_20446);
or UO_1658 (O_1658,N_20736,N_24507);
nand UO_1659 (O_1659,N_21768,N_23047);
nand UO_1660 (O_1660,N_24724,N_22003);
nand UO_1661 (O_1661,N_24606,N_23301);
nor UO_1662 (O_1662,N_23463,N_20603);
nor UO_1663 (O_1663,N_21672,N_19778);
nor UO_1664 (O_1664,N_23852,N_22947);
nand UO_1665 (O_1665,N_21019,N_21978);
and UO_1666 (O_1666,N_19964,N_24165);
or UO_1667 (O_1667,N_21835,N_21794);
nor UO_1668 (O_1668,N_23586,N_24818);
nor UO_1669 (O_1669,N_18916,N_21790);
nor UO_1670 (O_1670,N_19823,N_22926);
or UO_1671 (O_1671,N_22749,N_20450);
or UO_1672 (O_1672,N_23813,N_24164);
nand UO_1673 (O_1673,N_19406,N_19541);
xor UO_1674 (O_1674,N_20794,N_19070);
nor UO_1675 (O_1675,N_20985,N_20689);
or UO_1676 (O_1676,N_20732,N_22595);
and UO_1677 (O_1677,N_22710,N_20198);
nand UO_1678 (O_1678,N_22245,N_21333);
or UO_1679 (O_1679,N_22488,N_21265);
and UO_1680 (O_1680,N_24412,N_23705);
nor UO_1681 (O_1681,N_22224,N_20040);
nor UO_1682 (O_1682,N_23354,N_18994);
nand UO_1683 (O_1683,N_19170,N_22379);
and UO_1684 (O_1684,N_19579,N_19239);
nand UO_1685 (O_1685,N_23236,N_22795);
or UO_1686 (O_1686,N_22312,N_18800);
nand UO_1687 (O_1687,N_23975,N_22048);
nand UO_1688 (O_1688,N_22743,N_22847);
nor UO_1689 (O_1689,N_22660,N_20541);
and UO_1690 (O_1690,N_23157,N_18895);
nor UO_1691 (O_1691,N_19031,N_20544);
or UO_1692 (O_1692,N_21848,N_21912);
nor UO_1693 (O_1693,N_23053,N_22802);
and UO_1694 (O_1694,N_19459,N_18865);
nand UO_1695 (O_1695,N_20823,N_18986);
and UO_1696 (O_1696,N_21585,N_23489);
or UO_1697 (O_1697,N_21631,N_23932);
or UO_1698 (O_1698,N_20263,N_23020);
xnor UO_1699 (O_1699,N_24274,N_23735);
or UO_1700 (O_1700,N_19993,N_22004);
nand UO_1701 (O_1701,N_22168,N_21867);
or UO_1702 (O_1702,N_24528,N_24524);
nor UO_1703 (O_1703,N_22473,N_19587);
or UO_1704 (O_1704,N_20504,N_22568);
nor UO_1705 (O_1705,N_19593,N_21518);
and UO_1706 (O_1706,N_23679,N_23959);
xnor UO_1707 (O_1707,N_23750,N_23228);
nand UO_1708 (O_1708,N_21909,N_19035);
or UO_1709 (O_1709,N_21863,N_24781);
nand UO_1710 (O_1710,N_19916,N_24384);
nor UO_1711 (O_1711,N_23493,N_22821);
nor UO_1712 (O_1712,N_23088,N_19953);
or UO_1713 (O_1713,N_23785,N_23942);
or UO_1714 (O_1714,N_20933,N_23808);
or UO_1715 (O_1715,N_19674,N_18966);
and UO_1716 (O_1716,N_20421,N_24994);
and UO_1717 (O_1717,N_20619,N_22943);
or UO_1718 (O_1718,N_18828,N_19091);
or UO_1719 (O_1719,N_23918,N_20553);
or UO_1720 (O_1720,N_20761,N_24674);
nor UO_1721 (O_1721,N_18936,N_23233);
or UO_1722 (O_1722,N_18815,N_22612);
or UO_1723 (O_1723,N_20160,N_22924);
and UO_1724 (O_1724,N_22367,N_20754);
nand UO_1725 (O_1725,N_24874,N_21262);
and UO_1726 (O_1726,N_23827,N_20165);
and UO_1727 (O_1727,N_21185,N_20354);
and UO_1728 (O_1728,N_23231,N_19679);
nor UO_1729 (O_1729,N_23376,N_21500);
xnor UO_1730 (O_1730,N_20981,N_24103);
or UO_1731 (O_1731,N_24722,N_23275);
and UO_1732 (O_1732,N_24326,N_23475);
and UO_1733 (O_1733,N_21658,N_23508);
or UO_1734 (O_1734,N_22954,N_21406);
and UO_1735 (O_1735,N_24097,N_23902);
nor UO_1736 (O_1736,N_21302,N_19632);
and UO_1737 (O_1737,N_20465,N_21280);
or UO_1738 (O_1738,N_22565,N_23999);
nand UO_1739 (O_1739,N_21214,N_23544);
nand UO_1740 (O_1740,N_21721,N_22678);
or UO_1741 (O_1741,N_23650,N_21109);
nand UO_1742 (O_1742,N_22055,N_24067);
nor UO_1743 (O_1743,N_22553,N_21030);
and UO_1744 (O_1744,N_22410,N_18784);
nand UO_1745 (O_1745,N_22422,N_19477);
and UO_1746 (O_1746,N_22780,N_21531);
nand UO_1747 (O_1747,N_20988,N_22081);
nand UO_1748 (O_1748,N_22430,N_23181);
and UO_1749 (O_1749,N_22492,N_20408);
and UO_1750 (O_1750,N_19267,N_23910);
and UO_1751 (O_1751,N_21564,N_23636);
nor UO_1752 (O_1752,N_21808,N_24622);
and UO_1753 (O_1753,N_18889,N_22792);
or UO_1754 (O_1754,N_20859,N_19381);
and UO_1755 (O_1755,N_23174,N_24927);
and UO_1756 (O_1756,N_23481,N_21593);
nand UO_1757 (O_1757,N_20147,N_21626);
nor UO_1758 (O_1758,N_19405,N_23244);
nor UO_1759 (O_1759,N_20623,N_18761);
or UO_1760 (O_1760,N_21810,N_21513);
and UO_1761 (O_1761,N_23263,N_23151);
nand UO_1762 (O_1762,N_19069,N_20293);
or UO_1763 (O_1763,N_22570,N_20080);
nor UO_1764 (O_1764,N_22784,N_20248);
nand UO_1765 (O_1765,N_18860,N_21159);
nor UO_1766 (O_1766,N_19243,N_20660);
nor UO_1767 (O_1767,N_22089,N_21065);
nor UO_1768 (O_1768,N_20613,N_19898);
xnor UO_1769 (O_1769,N_24045,N_22493);
nor UO_1770 (O_1770,N_22564,N_24352);
nand UO_1771 (O_1771,N_22576,N_22964);
nor UO_1772 (O_1772,N_20841,N_20372);
nand UO_1773 (O_1773,N_20857,N_23035);
nor UO_1774 (O_1774,N_23215,N_23388);
xor UO_1775 (O_1775,N_20599,N_24799);
nor UO_1776 (O_1776,N_22910,N_19626);
and UO_1777 (O_1777,N_23184,N_20192);
nor UO_1778 (O_1778,N_20086,N_23000);
and UO_1779 (O_1779,N_18783,N_20329);
or UO_1780 (O_1780,N_21999,N_20234);
and UO_1781 (O_1781,N_19862,N_22050);
nand UO_1782 (O_1782,N_20063,N_20290);
nor UO_1783 (O_1783,N_19930,N_24830);
nor UO_1784 (O_1784,N_21015,N_20579);
or UO_1785 (O_1785,N_23721,N_18863);
or UO_1786 (O_1786,N_21841,N_22757);
nor UO_1787 (O_1787,N_21365,N_21235);
xnor UO_1788 (O_1788,N_21189,N_19555);
nor UO_1789 (O_1789,N_24069,N_20141);
nor UO_1790 (O_1790,N_22496,N_22773);
xor UO_1791 (O_1791,N_24262,N_22962);
nor UO_1792 (O_1792,N_19858,N_20058);
nor UO_1793 (O_1793,N_22065,N_20665);
and UO_1794 (O_1794,N_20069,N_24595);
and UO_1795 (O_1795,N_22256,N_22596);
and UO_1796 (O_1796,N_22920,N_20231);
nand UO_1797 (O_1797,N_24237,N_19902);
nor UO_1798 (O_1798,N_20876,N_21094);
nand UO_1799 (O_1799,N_20167,N_24002);
nand UO_1800 (O_1800,N_20373,N_24481);
nor UO_1801 (O_1801,N_21930,N_24997);
nor UO_1802 (O_1802,N_22923,N_20972);
nor UO_1803 (O_1803,N_19184,N_21699);
or UO_1804 (O_1804,N_20480,N_20066);
and UO_1805 (O_1805,N_21724,N_19673);
nor UO_1806 (O_1806,N_19841,N_24050);
and UO_1807 (O_1807,N_20524,N_22622);
and UO_1808 (O_1808,N_23075,N_22082);
or UO_1809 (O_1809,N_18838,N_22786);
xnor UO_1810 (O_1810,N_24660,N_22541);
nor UO_1811 (O_1811,N_18983,N_24691);
nor UO_1812 (O_1812,N_24194,N_19915);
nor UO_1813 (O_1813,N_23109,N_24728);
nor UO_1814 (O_1814,N_20394,N_20659);
or UO_1815 (O_1815,N_23373,N_19409);
nand UO_1816 (O_1816,N_20155,N_23944);
and UO_1817 (O_1817,N_24665,N_21596);
nand UO_1818 (O_1818,N_19687,N_19546);
nand UO_1819 (O_1819,N_22500,N_21946);
nand UO_1820 (O_1820,N_19767,N_22098);
xnor UO_1821 (O_1821,N_18961,N_24025);
and UO_1822 (O_1822,N_20640,N_19631);
and UO_1823 (O_1823,N_19360,N_21241);
xor UO_1824 (O_1824,N_24395,N_22791);
nand UO_1825 (O_1825,N_19369,N_24630);
and UO_1826 (O_1826,N_21665,N_23726);
or UO_1827 (O_1827,N_24652,N_24153);
and UO_1828 (O_1828,N_20217,N_24835);
and UO_1829 (O_1829,N_19362,N_19713);
and UO_1830 (O_1830,N_20721,N_23119);
nor UO_1831 (O_1831,N_19801,N_21093);
and UO_1832 (O_1832,N_24703,N_22406);
or UO_1833 (O_1833,N_20472,N_21013);
or UO_1834 (O_1834,N_21883,N_18876);
nand UO_1835 (O_1835,N_20252,N_22674);
nand UO_1836 (O_1836,N_18837,N_20967);
or UO_1837 (O_1837,N_19036,N_18953);
nand UO_1838 (O_1838,N_23689,N_20087);
or UO_1839 (O_1839,N_24980,N_20919);
and UO_1840 (O_1840,N_23563,N_22348);
nor UO_1841 (O_1841,N_21783,N_21200);
nor UO_1842 (O_1842,N_21547,N_24033);
and UO_1843 (O_1843,N_21475,N_23566);
xnor UO_1844 (O_1844,N_21871,N_19052);
nor UO_1845 (O_1845,N_22403,N_19101);
nand UO_1846 (O_1846,N_21085,N_20253);
xor UO_1847 (O_1847,N_19425,N_19104);
and UO_1848 (O_1848,N_20900,N_22091);
and UO_1849 (O_1849,N_20737,N_22864);
or UO_1850 (O_1850,N_20715,N_21372);
or UO_1851 (O_1851,N_19664,N_20643);
or UO_1852 (O_1852,N_24350,N_20775);
nor UO_1853 (O_1853,N_19216,N_21598);
nand UO_1854 (O_1854,N_21562,N_23671);
and UO_1855 (O_1855,N_18887,N_19945);
or UO_1856 (O_1856,N_19787,N_21919);
nand UO_1857 (O_1857,N_23779,N_21827);
nand UO_1858 (O_1858,N_23449,N_22108);
or UO_1859 (O_1859,N_24076,N_21664);
nand UO_1860 (O_1860,N_19811,N_20747);
nor UO_1861 (O_1861,N_24019,N_20650);
xor UO_1862 (O_1862,N_24034,N_18801);
or UO_1863 (O_1863,N_20288,N_19053);
nand UO_1864 (O_1864,N_21838,N_21524);
or UO_1865 (O_1865,N_23988,N_19554);
nand UO_1866 (O_1866,N_23495,N_19825);
nor UO_1867 (O_1867,N_23529,N_18873);
or UO_1868 (O_1868,N_18839,N_22347);
or UO_1869 (O_1869,N_19083,N_22327);
and UO_1870 (O_1870,N_24928,N_20916);
or UO_1871 (O_1871,N_20304,N_23509);
and UO_1872 (O_1872,N_22681,N_20538);
nand UO_1873 (O_1873,N_24693,N_24804);
and UO_1874 (O_1874,N_22092,N_23165);
and UO_1875 (O_1875,N_23723,N_23142);
and UO_1876 (O_1876,N_23453,N_23498);
nor UO_1877 (O_1877,N_22586,N_21451);
or UO_1878 (O_1878,N_22152,N_19269);
nand UO_1879 (O_1879,N_21146,N_23042);
or UO_1880 (O_1880,N_22265,N_21023);
and UO_1881 (O_1881,N_24734,N_21990);
xnor UO_1882 (O_1882,N_23989,N_24054);
and UO_1883 (O_1883,N_24886,N_24802);
nand UO_1884 (O_1884,N_21575,N_23341);
nand UO_1885 (O_1885,N_20053,N_20584);
or UO_1886 (O_1886,N_22022,N_24840);
and UO_1887 (O_1887,N_22863,N_23294);
and UO_1888 (O_1888,N_22480,N_19703);
xnor UO_1889 (O_1889,N_23344,N_21308);
xor UO_1890 (O_1890,N_24053,N_24006);
or UO_1891 (O_1891,N_21137,N_23464);
nor UO_1892 (O_1892,N_19906,N_23538);
nor UO_1893 (O_1893,N_19202,N_19934);
nand UO_1894 (O_1894,N_19717,N_21343);
nor UO_1895 (O_1895,N_21693,N_22862);
and UO_1896 (O_1896,N_19601,N_21605);
nor UO_1897 (O_1897,N_20885,N_24128);
xor UO_1898 (O_1898,N_21068,N_19892);
nor UO_1899 (O_1899,N_23849,N_22787);
or UO_1900 (O_1900,N_20168,N_20497);
or UO_1901 (O_1901,N_20120,N_23450);
nand UO_1902 (O_1902,N_21126,N_19791);
and UO_1903 (O_1903,N_22738,N_21199);
nor UO_1904 (O_1904,N_23792,N_20580);
or UO_1905 (O_1905,N_22774,N_22567);
and UO_1906 (O_1906,N_22060,N_24537);
and UO_1907 (O_1907,N_21246,N_22701);
or UO_1908 (O_1908,N_19730,N_24114);
nand UO_1909 (O_1909,N_23034,N_24548);
nor UO_1910 (O_1910,N_24063,N_21347);
nand UO_1911 (O_1911,N_22973,N_22982);
nand UO_1912 (O_1912,N_21510,N_24137);
or UO_1913 (O_1913,N_24149,N_23271);
and UO_1914 (O_1914,N_23466,N_20113);
nor UO_1915 (O_1915,N_24272,N_19299);
nor UO_1916 (O_1916,N_24360,N_21042);
xnor UO_1917 (O_1917,N_23862,N_20287);
or UO_1918 (O_1918,N_24954,N_18912);
nor UO_1919 (O_1919,N_24356,N_19961);
and UO_1920 (O_1920,N_24610,N_19739);
nand UO_1921 (O_1921,N_18955,N_23375);
xor UO_1922 (O_1922,N_20132,N_19225);
or UO_1923 (O_1923,N_19751,N_22061);
nand UO_1924 (O_1924,N_22404,N_20172);
nor UO_1925 (O_1925,N_22857,N_24860);
nor UO_1926 (O_1926,N_21682,N_22939);
nand UO_1927 (O_1927,N_23342,N_24211);
or UO_1928 (O_1928,N_22330,N_19423);
or UO_1929 (O_1929,N_21361,N_24180);
and UO_1930 (O_1930,N_20674,N_24600);
or UO_1931 (O_1931,N_24776,N_20873);
nor UO_1932 (O_1932,N_24662,N_23285);
and UO_1933 (O_1933,N_24015,N_22515);
nand UO_1934 (O_1934,N_24601,N_22465);
nand UO_1935 (O_1935,N_23736,N_23438);
nand UO_1936 (O_1936,N_22361,N_24931);
and UO_1937 (O_1937,N_23242,N_21528);
or UO_1938 (O_1938,N_24813,N_23169);
and UO_1939 (O_1939,N_24491,N_24140);
nor UO_1940 (O_1940,N_22026,N_24236);
nand UO_1941 (O_1941,N_19771,N_19089);
nand UO_1942 (O_1942,N_19152,N_23675);
nor UO_1943 (O_1943,N_22739,N_24762);
nand UO_1944 (O_1944,N_21385,N_19733);
xor UO_1945 (O_1945,N_22585,N_23631);
or UO_1946 (O_1946,N_19894,N_21992);
or UO_1947 (O_1947,N_24440,N_22494);
or UO_1948 (O_1948,N_24909,N_23703);
xor UO_1949 (O_1949,N_21816,N_18842);
nand UO_1950 (O_1950,N_20991,N_20830);
nand UO_1951 (O_1951,N_24302,N_19186);
and UO_1952 (O_1952,N_19903,N_18965);
and UO_1953 (O_1953,N_24612,N_19244);
and UO_1954 (O_1954,N_20733,N_19215);
and UO_1955 (O_1955,N_21995,N_19569);
nor UO_1956 (O_1956,N_20201,N_21049);
nand UO_1957 (O_1957,N_19333,N_20225);
nor UO_1958 (O_1958,N_23355,N_20238);
xnor UO_1959 (O_1959,N_21970,N_21456);
nand UO_1960 (O_1960,N_20787,N_22356);
nand UO_1961 (O_1961,N_22713,N_21057);
xnor UO_1962 (O_1962,N_23891,N_19879);
or UO_1963 (O_1963,N_24547,N_21688);
xnor UO_1964 (O_1964,N_19764,N_23200);
nor UO_1965 (O_1965,N_19755,N_22657);
nor UO_1966 (O_1966,N_21358,N_23442);
nor UO_1967 (O_1967,N_21818,N_20223);
xor UO_1968 (O_1968,N_24596,N_21578);
nor UO_1969 (O_1969,N_19232,N_20360);
nor UO_1970 (O_1970,N_21362,N_23592);
and UO_1971 (O_1971,N_18937,N_20970);
nand UO_1972 (O_1972,N_20633,N_23204);
nand UO_1973 (O_1973,N_20038,N_24644);
nand UO_1974 (O_1974,N_22721,N_24141);
and UO_1975 (O_1975,N_22071,N_21662);
and UO_1976 (O_1976,N_23304,N_21202);
nand UO_1977 (O_1977,N_23666,N_22223);
xnor UO_1978 (O_1978,N_24208,N_24756);
nand UO_1979 (O_1979,N_23784,N_21561);
or UO_1980 (O_1980,N_23894,N_21052);
or UO_1981 (O_1981,N_24967,N_20050);
or UO_1982 (O_1982,N_20340,N_21341);
nor UO_1983 (O_1983,N_19608,N_22823);
nand UO_1984 (O_1984,N_21066,N_24187);
or UO_1985 (O_1985,N_21363,N_21921);
and UO_1986 (O_1986,N_19119,N_21154);
nor UO_1987 (O_1987,N_24231,N_20863);
and UO_1988 (O_1988,N_24585,N_22960);
nor UO_1989 (O_1989,N_22076,N_24597);
or UO_1990 (O_1990,N_23025,N_22690);
nand UO_1991 (O_1991,N_23202,N_23812);
nand UO_1992 (O_1992,N_19534,N_23993);
or UO_1993 (O_1993,N_22760,N_23145);
xnor UO_1994 (O_1994,N_19937,N_21858);
nand UO_1995 (O_1995,N_24527,N_23302);
and UO_1996 (O_1996,N_22588,N_20983);
and UO_1997 (O_1997,N_22659,N_19417);
nor UO_1998 (O_1998,N_24774,N_24816);
nand UO_1999 (O_1999,N_21924,N_18786);
nor UO_2000 (O_2000,N_23577,N_21700);
or UO_2001 (O_2001,N_22411,N_21826);
xor UO_2002 (O_2002,N_23408,N_20411);
nand UO_2003 (O_2003,N_22479,N_21847);
xnor UO_2004 (O_2004,N_19026,N_22695);
or UO_2005 (O_2005,N_24470,N_20286);
and UO_2006 (O_2006,N_19301,N_23472);
nand UO_2007 (O_2007,N_20519,N_22135);
xor UO_2008 (O_2008,N_21495,N_18903);
and UO_2009 (O_2009,N_23316,N_21390);
nor UO_2010 (O_2010,N_22944,N_21796);
nor UO_2011 (O_2011,N_18987,N_19148);
nand UO_2012 (O_2012,N_21935,N_23652);
xnor UO_2013 (O_2013,N_19889,N_21701);
or UO_2014 (O_2014,N_22871,N_19310);
nor UO_2015 (O_2015,N_24008,N_19861);
or UO_2016 (O_2016,N_23206,N_19789);
and UO_2017 (O_2017,N_20348,N_20958);
and UO_2018 (O_2018,N_23672,N_22640);
or UO_2019 (O_2019,N_19470,N_23405);
nor UO_2020 (O_2020,N_20852,N_22643);
nor UO_2021 (O_2021,N_23087,N_23329);
nand UO_2022 (O_2022,N_20014,N_21535);
nand UO_2023 (O_2023,N_21685,N_23399);
nand UO_2024 (O_2024,N_19043,N_21028);
or UO_2025 (O_2025,N_21996,N_22527);
xor UO_2026 (O_2026,N_21890,N_19770);
or UO_2027 (O_2027,N_18843,N_19054);
xor UO_2028 (O_2028,N_24649,N_18858);
and UO_2029 (O_2029,N_23649,N_21360);
and UO_2030 (O_2030,N_24221,N_22368);
or UO_2031 (O_2031,N_24834,N_22332);
xnor UO_2032 (O_2032,N_22776,N_19697);
or UO_2033 (O_2033,N_24821,N_23073);
xnor UO_2034 (O_2034,N_21264,N_22171);
nand UO_2035 (O_2035,N_20883,N_20912);
nor UO_2036 (O_2036,N_19393,N_19621);
nand UO_2037 (O_2037,N_23878,N_19570);
nand UO_2038 (O_2038,N_24116,N_20875);
and UO_2039 (O_2039,N_24982,N_19309);
or UO_2040 (O_2040,N_22728,N_19795);
nor UO_2041 (O_2041,N_23266,N_19220);
or UO_2042 (O_2042,N_23965,N_24243);
nand UO_2043 (O_2043,N_20211,N_22010);
nor UO_2044 (O_2044,N_21965,N_24684);
or UO_2045 (O_2045,N_21897,N_22357);
and UO_2046 (O_2046,N_22373,N_21018);
nor UO_2047 (O_2047,N_23897,N_24920);
nor UO_2048 (O_2048,N_22241,N_24482);
nand UO_2049 (O_2049,N_22459,N_22449);
and UO_2050 (O_2050,N_20149,N_23327);
and UO_2051 (O_2051,N_21005,N_22334);
or UO_2052 (O_2052,N_23974,N_19013);
or UO_2053 (O_2053,N_22212,N_19090);
and UO_2054 (O_2054,N_22609,N_19093);
or UO_2055 (O_2055,N_24193,N_22756);
and UO_2056 (O_2056,N_21125,N_22094);
or UO_2057 (O_2057,N_19045,N_20808);
xor UO_2058 (O_2058,N_22096,N_22138);
nand UO_2059 (O_2059,N_22686,N_19488);
nor UO_2060 (O_2060,N_20320,N_21833);
or UO_2061 (O_2061,N_19287,N_22257);
and UO_2062 (O_2062,N_22291,N_20974);
nor UO_2063 (O_2063,N_23632,N_20136);
nor UO_2064 (O_2064,N_22707,N_24484);
and UO_2065 (O_2065,N_22209,N_23570);
nand UO_2066 (O_2066,N_23819,N_23485);
nand UO_2067 (O_2067,N_23071,N_24577);
nor UO_2068 (O_2068,N_18921,N_22879);
nor UO_2069 (O_2069,N_23931,N_22248);
xnor UO_2070 (O_2070,N_19878,N_23255);
or UO_2071 (O_2071,N_23229,N_20518);
nand UO_2072 (O_2072,N_22032,N_24581);
or UO_2073 (O_2073,N_22991,N_22271);
xnor UO_2074 (O_2074,N_23331,N_20559);
nor UO_2075 (O_2075,N_23061,N_19705);
nor UO_2076 (O_2076,N_22118,N_21058);
and UO_2077 (O_2077,N_19525,N_21582);
nor UO_2078 (O_2078,N_21364,N_23046);
nand UO_2079 (O_2079,N_18974,N_23892);
or UO_2080 (O_2080,N_24694,N_24992);
or UO_2081 (O_2081,N_24290,N_22617);
or UO_2082 (O_2082,N_23668,N_23595);
nor UO_2083 (O_2083,N_21191,N_24410);
and UO_2084 (O_2084,N_20901,N_18772);
and UO_2085 (O_2085,N_22997,N_19138);
and UO_2086 (O_2086,N_20555,N_24247);
and UO_2087 (O_2087,N_19653,N_19355);
nand UO_2088 (O_2088,N_20976,N_19356);
and UO_2089 (O_2089,N_22203,N_23725);
and UO_2090 (O_2090,N_22025,N_21824);
or UO_2091 (O_2091,N_20872,N_19182);
xor UO_2092 (O_2092,N_22188,N_23732);
or UO_2093 (O_2093,N_23115,N_20301);
or UO_2094 (O_2094,N_20560,N_24179);
nor UO_2095 (O_2095,N_22648,N_24058);
nor UO_2096 (O_2096,N_19544,N_24723);
nor UO_2097 (O_2097,N_19762,N_24393);
nor UO_2098 (O_2098,N_20003,N_20661);
or UO_2099 (O_2099,N_24826,N_23276);
or UO_2100 (O_2100,N_20370,N_20805);
or UO_2101 (O_2101,N_22464,N_24540);
nor UO_2102 (O_2102,N_24244,N_22971);
and UO_2103 (O_2103,N_23855,N_21480);
xnor UO_2104 (O_2104,N_19559,N_24516);
or UO_2105 (O_2105,N_22184,N_22554);
and UO_2106 (O_2106,N_19387,N_23051);
xor UO_2107 (O_2107,N_24823,N_19208);
nor UO_2108 (O_2108,N_22673,N_19130);
nor UO_2109 (O_2109,N_20679,N_23012);
and UO_2110 (O_2110,N_24133,N_21497);
and UO_2111 (O_2111,N_22134,N_18807);
nor UO_2112 (O_2112,N_19426,N_21232);
nand UO_2113 (O_2113,N_20904,N_22921);
nor UO_2114 (O_2114,N_19032,N_20140);
nor UO_2115 (O_2115,N_24206,N_20359);
nor UO_2116 (O_2116,N_23280,N_22013);
nor UO_2117 (O_2117,N_19071,N_23122);
nand UO_2118 (O_2118,N_23524,N_20478);
and UO_2119 (O_2119,N_20850,N_22214);
nor UO_2120 (O_2120,N_19431,N_22888);
nand UO_2121 (O_2121,N_22874,N_19509);
or UO_2122 (O_2122,N_22377,N_23740);
nand UO_2123 (O_2123,N_23861,N_20738);
and UO_2124 (O_2124,N_23719,N_21979);
xnor UO_2125 (O_2125,N_24448,N_21690);
and UO_2126 (O_2126,N_23633,N_19242);
nand UO_2127 (O_2127,N_22965,N_21616);
nor UO_2128 (O_2128,N_22296,N_20649);
nor UO_2129 (O_2129,N_22390,N_23753);
and UO_2130 (O_2130,N_19009,N_21223);
nor UO_2131 (O_2131,N_24825,N_21885);
nand UO_2132 (O_2132,N_18867,N_19188);
nand UO_2133 (O_2133,N_23084,N_24711);
nand UO_2134 (O_2134,N_19759,N_18871);
and UO_2135 (O_2135,N_23547,N_23998);
nand UO_2136 (O_2136,N_23384,N_21453);
or UO_2137 (O_2137,N_24843,N_22192);
nand UO_2138 (O_2138,N_20364,N_18908);
and UO_2139 (O_2139,N_19776,N_19391);
nand UO_2140 (O_2140,N_19099,N_24429);
nand UO_2141 (O_2141,N_20153,N_21936);
nor UO_2142 (O_2142,N_24169,N_24937);
nand UO_2143 (O_2143,N_20089,N_19655);
xnor UO_2144 (O_2144,N_18941,N_19448);
nor UO_2145 (O_2145,N_22691,N_21069);
and UO_2146 (O_2146,N_21878,N_24903);
and UO_2147 (O_2147,N_21731,N_20818);
and UO_2148 (O_2148,N_21606,N_22127);
or UO_2149 (O_2149,N_20365,N_23469);
or UO_2150 (O_2150,N_24117,N_19884);
or UO_2151 (O_2151,N_22289,N_22672);
or UO_2152 (O_2152,N_19804,N_20073);
or UO_2153 (O_2153,N_24536,N_21083);
or UO_2154 (O_2154,N_20085,N_19295);
and UO_2155 (O_2155,N_20718,N_24111);
or UO_2156 (O_2156,N_21021,N_22861);
nor UO_2157 (O_2157,N_20585,N_20547);
nor UO_2158 (O_2158,N_23358,N_18894);
and UO_2159 (O_2159,N_21484,N_21546);
or UO_2160 (O_2160,N_24152,N_20893);
nand UO_2161 (O_2161,N_23310,N_21297);
and UO_2162 (O_2162,N_21398,N_20962);
nand UO_2163 (O_2163,N_20221,N_23300);
nor UO_2164 (O_2164,N_23872,N_20218);
and UO_2165 (O_2165,N_23839,N_19987);
and UO_2166 (O_2166,N_23068,N_24552);
or UO_2167 (O_2167,N_19371,N_18952);
nand UO_2168 (O_2168,N_21976,N_23224);
and UO_2169 (O_2169,N_21643,N_18756);
nor UO_2170 (O_2170,N_24889,N_23264);
nand UO_2171 (O_2171,N_21969,N_22763);
nor UO_2172 (O_2172,N_22122,N_23159);
nor UO_2173 (O_2173,N_23700,N_24983);
xor UO_2174 (O_2174,N_19813,N_19464);
and UO_2175 (O_2175,N_22951,N_22881);
or UO_2176 (O_2176,N_19444,N_24347);
and UO_2177 (O_2177,N_22716,N_19073);
or UO_2178 (O_2178,N_22932,N_20041);
and UO_2179 (O_2179,N_23049,N_19178);
or UO_2180 (O_2180,N_20067,N_23611);
nor UO_2181 (O_2181,N_22870,N_24730);
and UO_2182 (O_2182,N_19322,N_19300);
xor UO_2183 (O_2183,N_21650,N_22294);
nor UO_2184 (O_2184,N_19261,N_24310);
and UO_2185 (O_2185,N_20131,N_22680);
and UO_2186 (O_2186,N_19085,N_24404);
nand UO_2187 (O_2187,N_22034,N_20697);
nor UO_2188 (O_2188,N_22447,N_22191);
xnor UO_2189 (O_2189,N_18900,N_21249);
xor UO_2190 (O_2190,N_20891,N_24341);
nand UO_2191 (O_2191,N_19975,N_24914);
nand UO_2192 (O_2192,N_23727,N_23079);
and UO_2193 (O_2193,N_21326,N_23778);
or UO_2194 (O_2194,N_23155,N_24425);
nor UO_2195 (O_2195,N_23701,N_20826);
and UO_2196 (O_2196,N_24009,N_23562);
nor UO_2197 (O_2197,N_18964,N_23013);
and UO_2198 (O_2198,N_19814,N_21698);
or UO_2199 (O_2199,N_22288,N_21124);
or UO_2200 (O_2200,N_23407,N_24654);
nor UO_2201 (O_2201,N_21195,N_22251);
nor UO_2202 (O_2202,N_23208,N_23043);
nand UO_2203 (O_2203,N_19479,N_20523);
or UO_2204 (O_2204,N_19666,N_20052);
xnor UO_2205 (O_2205,N_19741,N_21925);
xor UO_2206 (O_2206,N_21161,N_23520);
nand UO_2207 (O_2207,N_20612,N_19938);
nor UO_2208 (O_2208,N_22059,N_23761);
or UO_2209 (O_2209,N_18944,N_23314);
nand UO_2210 (O_2210,N_21432,N_22714);
or UO_2211 (O_2211,N_19158,N_21594);
or UO_2212 (O_2212,N_21504,N_19246);
nand UO_2213 (O_2213,N_19782,N_24755);
and UO_2214 (O_2214,N_19214,N_20847);
or UO_2215 (O_2215,N_19722,N_24311);
or UO_2216 (O_2216,N_24394,N_24391);
and UO_2217 (O_2217,N_21732,N_21376);
and UO_2218 (O_2218,N_22236,N_20610);
and UO_2219 (O_2219,N_23421,N_19885);
or UO_2220 (O_2220,N_21687,N_23801);
or UO_2221 (O_2221,N_21067,N_23210);
nand UO_2222 (O_2222,N_18836,N_21860);
or UO_2223 (O_2223,N_24803,N_22394);
nand UO_2224 (O_2224,N_18763,N_22781);
xor UO_2225 (O_2225,N_24478,N_23714);
or UO_2226 (O_2226,N_21931,N_21397);
or UO_2227 (O_2227,N_24910,N_24768);
or UO_2228 (O_2228,N_23239,N_24241);
nand UO_2229 (O_2229,N_21851,N_21649);
or UO_2230 (O_2230,N_19978,N_24022);
nand UO_2231 (O_2231,N_23023,N_19323);
nor UO_2232 (O_2232,N_21691,N_24996);
and UO_2233 (O_2233,N_21413,N_21103);
nor UO_2234 (O_2234,N_20550,N_23567);
and UO_2235 (O_2235,N_20302,N_21870);
nand UO_2236 (O_2236,N_19517,N_22418);
and UO_2237 (O_2237,N_22551,N_23756);
and UO_2238 (O_2238,N_21213,N_19505);
nor UO_2239 (O_2239,N_23345,N_21328);
and UO_2240 (O_2240,N_21603,N_21822);
nor UO_2241 (O_2241,N_24040,N_22353);
nand UO_2242 (O_2242,N_23531,N_20724);
and UO_2243 (O_2243,N_20496,N_22529);
and UO_2244 (O_2244,N_20868,N_23758);
and UO_2245 (O_2245,N_22318,N_23104);
xor UO_2246 (O_2246,N_24900,N_20482);
or UO_2247 (O_2247,N_22159,N_23098);
and UO_2248 (O_2248,N_21516,N_20325);
or UO_2249 (O_2249,N_23973,N_21132);
nand UO_2250 (O_2250,N_23426,N_23906);
or UO_2251 (O_2251,N_19583,N_22752);
or UO_2252 (O_2252,N_21024,N_20704);
or UO_2253 (O_2253,N_23393,N_24792);
and UO_2254 (O_2254,N_20258,N_23939);
or UO_2255 (O_2255,N_21745,N_22833);
and UO_2256 (O_2256,N_24166,N_19113);
nor UO_2257 (O_2257,N_20625,N_20130);
nor UO_2258 (O_2258,N_19922,N_19772);
nand UO_2259 (O_2259,N_20436,N_21095);
nand UO_2260 (O_2260,N_19847,N_24938);
and UO_2261 (O_2261,N_21135,N_23536);
and UO_2262 (O_2262,N_20335,N_23692);
nor UO_2263 (O_2263,N_22090,N_20342);
and UO_2264 (O_2264,N_22031,N_20266);
nand UO_2265 (O_2265,N_24625,N_21181);
nand UO_2266 (O_2266,N_21583,N_20272);
or UO_2267 (O_2267,N_21444,N_23089);
nand UO_2268 (O_2268,N_20759,N_24894);
nor UO_2269 (O_2269,N_21116,N_21120);
and UO_2270 (O_2270,N_21188,N_24555);
nand UO_2271 (O_2271,N_21489,N_24066);
nand UO_2272 (O_2272,N_20415,N_20146);
or UO_2273 (O_2273,N_23532,N_19200);
or UO_2274 (O_2274,N_23686,N_20122);
xor UO_2275 (O_2275,N_23353,N_22815);
nor UO_2276 (O_2276,N_22219,N_21852);
xnor UO_2277 (O_2277,N_18959,N_24715);
or UO_2278 (O_2278,N_22008,N_23357);
nand UO_2279 (O_2279,N_23771,N_24590);
nor UO_2280 (O_2280,N_24435,N_21550);
and UO_2281 (O_2281,N_20189,N_19706);
or UO_2282 (O_2282,N_22983,N_19635);
nor UO_2283 (O_2283,N_20152,N_21537);
and UO_2284 (O_2284,N_22866,N_22287);
nor UO_2285 (O_2285,N_19913,N_19201);
xnor UO_2286 (O_2286,N_22227,N_21926);
or UO_2287 (O_2287,N_20700,N_19553);
xnor UO_2288 (O_2288,N_21670,N_23984);
nand UO_2289 (O_2289,N_21389,N_23394);
nand UO_2290 (O_2290,N_20851,N_23916);
and UO_2291 (O_2291,N_24770,N_20742);
or UO_2292 (O_2292,N_22668,N_23648);
and UO_2293 (O_2293,N_19662,N_21307);
nand UO_2294 (O_2294,N_19401,N_19190);
nor UO_2295 (O_2295,N_23415,N_23803);
and UO_2296 (O_2296,N_20998,N_23220);
nor UO_2297 (O_2297,N_19481,N_22412);
nor UO_2298 (O_2298,N_22189,N_21922);
nor UO_2299 (O_2299,N_23644,N_21960);
and UO_2300 (O_2300,N_22968,N_21207);
and UO_2301 (O_2301,N_19424,N_23191);
nor UO_2302 (O_2302,N_20163,N_23328);
nand UO_2303 (O_2303,N_20278,N_19339);
or UO_2304 (O_2304,N_22126,N_24561);
or UO_2305 (O_2305,N_24358,N_24420);
and UO_2306 (O_2306,N_21064,N_22125);
nand UO_2307 (O_2307,N_23659,N_19756);
xor UO_2308 (O_2308,N_24922,N_18823);
and UO_2309 (O_2309,N_21275,N_20594);
and UO_2310 (O_2310,N_22085,N_23240);
nor UO_2311 (O_2311,N_23348,N_19971);
or UO_2312 (O_2312,N_22907,N_19865);
and UO_2313 (O_2313,N_22867,N_21648);
nor UO_2314 (O_2314,N_23052,N_18885);
and UO_2315 (O_2315,N_19266,N_23899);
and UO_2316 (O_2316,N_20268,N_21080);
or UO_2317 (O_2317,N_20337,N_18929);
and UO_2318 (O_2318,N_19780,N_24659);
nor UO_2319 (O_2319,N_24544,N_19145);
or UO_2320 (O_2320,N_24737,N_20925);
and UO_2321 (O_2321,N_21243,N_19276);
or UO_2322 (O_2322,N_24016,N_22167);
nand UO_2323 (O_2323,N_22916,N_20987);
or UO_2324 (O_2324,N_22810,N_21337);
or UO_2325 (O_2325,N_20939,N_24064);
nand UO_2326 (O_2326,N_21602,N_19189);
and UO_2327 (O_2327,N_21396,N_20498);
and UO_2328 (O_2328,N_20540,N_20994);
and UO_2329 (O_2329,N_19748,N_24134);
or UO_2330 (O_2330,N_23667,N_19972);
and UO_2331 (O_2331,N_24543,N_20911);
or UO_2332 (O_2332,N_21074,N_22421);
nor UO_2333 (O_2333,N_19719,N_23946);
or UO_2334 (O_2334,N_22314,N_19911);
nand UO_2335 (O_2335,N_22151,N_20479);
or UO_2336 (O_2336,N_20942,N_23182);
or UO_2337 (O_2337,N_23523,N_21570);
and UO_2338 (O_2338,N_24783,N_23192);
or UO_2339 (O_2339,N_23334,N_21549);
or UO_2340 (O_2340,N_20064,N_22252);
nand UO_2341 (O_2341,N_22163,N_23108);
nand UO_2342 (O_2342,N_23010,N_19248);
and UO_2343 (O_2343,N_20637,N_21442);
nor UO_2344 (O_2344,N_21744,N_21913);
nor UO_2345 (O_2345,N_20057,N_20664);
nand UO_2346 (O_2346,N_19432,N_22170);
nor UO_2347 (O_2347,N_20076,N_24281);
nor UO_2348 (O_2348,N_22525,N_24671);
nand UO_2349 (O_2349,N_23112,N_19418);
xor UO_2350 (O_2350,N_20443,N_23530);
nor UO_2351 (O_2351,N_24269,N_24198);
xor UO_2352 (O_2352,N_18767,N_23657);
or UO_2353 (O_2353,N_21051,N_24218);
nor UO_2354 (O_2354,N_24748,N_21388);
xnor UO_2355 (O_2355,N_23581,N_20953);
and UO_2356 (O_2356,N_23390,N_19465);
xnor UO_2357 (O_2357,N_19850,N_23982);
nand UO_2358 (O_2358,N_24985,N_22439);
xnor UO_2359 (O_2359,N_19056,N_24530);
and UO_2360 (O_2360,N_19925,N_21342);
nor UO_2361 (O_2361,N_23232,N_22839);
nand UO_2362 (O_2362,N_22719,N_24001);
nor UO_2363 (O_2363,N_24343,N_19273);
nand UO_2364 (O_2364,N_21910,N_20021);
xor UO_2365 (O_2365,N_23492,N_24882);
xor UO_2366 (O_2366,N_21433,N_24918);
nand UO_2367 (O_2367,N_24651,N_19806);
and UO_2368 (O_2368,N_23211,N_22759);
or UO_2369 (O_2369,N_23908,N_23585);
xnor UO_2370 (O_2370,N_18862,N_19380);
nand UO_2371 (O_2371,N_21713,N_24345);
or UO_2372 (O_2372,N_19548,N_23537);
xnor UO_2373 (O_2373,N_22370,N_19774);
nor UO_2374 (O_2374,N_24160,N_19798);
xor UO_2375 (O_2375,N_19040,N_21692);
nand UO_2376 (O_2376,N_19066,N_22709);
and UO_2377 (O_2377,N_24121,N_19807);
or UO_2378 (O_2378,N_23322,N_23847);
nor UO_2379 (O_2379,N_21450,N_24731);
nand UO_2380 (O_2380,N_21723,N_23558);
and UO_2381 (O_2381,N_24084,N_18795);
nand UO_2382 (O_2382,N_21543,N_20054);
nor UO_2383 (O_2383,N_21884,N_24072);
and UO_2384 (O_2384,N_23195,N_19654);
xnor UO_2385 (O_2385,N_20769,N_22313);
nor UO_2386 (O_2386,N_23152,N_22891);
and UO_2387 (O_2387,N_21091,N_23130);
nor UO_2388 (O_2388,N_24668,N_24777);
nand UO_2389 (O_2389,N_20384,N_24398);
and UO_2390 (O_2390,N_18833,N_22750);
nand UO_2391 (O_2391,N_23110,N_19844);
nor UO_2392 (O_2392,N_20007,N_19640);
or UO_2393 (O_2393,N_21348,N_22682);
xnor UO_2394 (O_2394,N_24514,N_20037);
and UO_2395 (O_2395,N_18957,N_18906);
nand UO_2396 (O_2396,N_23126,N_21903);
or UO_2397 (O_2397,N_22671,N_21998);
nor UO_2398 (O_2398,N_21823,N_24397);
xnor UO_2399 (O_2399,N_23176,N_22509);
nand UO_2400 (O_2400,N_21106,N_23235);
nor UO_2401 (O_2401,N_23256,N_19102);
and UO_2402 (O_2402,N_19578,N_22321);
nor UO_2403 (O_2403,N_19694,N_19707);
nor UO_2404 (O_2404,N_21869,N_21483);
nor UO_2405 (O_2405,N_22485,N_18881);
or UO_2406 (O_2406,N_22199,N_22793);
and UO_2407 (O_2407,N_24940,N_23494);
xnor UO_2408 (O_2408,N_19163,N_20763);
nand UO_2409 (O_2409,N_22015,N_21750);
or UO_2410 (O_2410,N_23433,N_22666);
or UO_2411 (O_2411,N_22677,N_22336);
xor UO_2412 (O_2412,N_24788,N_24261);
or UO_2413 (O_2413,N_24178,N_23929);
and UO_2414 (O_2414,N_22798,N_19016);
or UO_2415 (O_2415,N_24096,N_20142);
nand UO_2416 (O_2416,N_21046,N_23313);
or UO_2417 (O_2417,N_20899,N_23781);
nor UO_2418 (O_2418,N_21521,N_19075);
nor UO_2419 (O_2419,N_24199,N_21591);
or UO_2420 (O_2420,N_19440,N_23970);
and UO_2421 (O_2421,N_21719,N_24623);
nand UO_2422 (O_2422,N_19125,N_21087);
nor UO_2423 (O_2423,N_20262,N_22239);
or UO_2424 (O_2424,N_20982,N_24645);
xor UO_2425 (O_2425,N_22323,N_22782);
or UO_2426 (O_2426,N_20299,N_24184);
nor UO_2427 (O_2427,N_20034,N_21599);
nor UO_2428 (O_2428,N_24087,N_23293);
and UO_2429 (O_2429,N_21290,N_19543);
nand UO_2430 (O_2430,N_19815,N_21225);
and UO_2431 (O_2431,N_23127,N_20106);
nor UO_2432 (O_2432,N_19065,N_24990);
or UO_2433 (O_2433,N_22255,N_19484);
and UO_2434 (O_2434,N_23967,N_20275);
and UO_2435 (O_2435,N_23747,N_24413);
or UO_2436 (O_2436,N_19007,N_24291);
and UO_2437 (O_2437,N_20552,N_22328);
nand UO_2438 (O_2438,N_24029,N_19996);
nor UO_2439 (O_2439,N_22024,N_21473);
nand UO_2440 (O_2440,N_18760,N_21176);
and UO_2441 (O_2441,N_18832,N_21929);
or UO_2442 (O_2442,N_22311,N_18771);
nand UO_2443 (O_2443,N_23250,N_24251);
nand UO_2444 (O_2444,N_24902,N_23400);
or UO_2445 (O_2445,N_22317,N_20543);
and UO_2446 (O_2446,N_24348,N_23588);
xnor UO_2447 (O_2447,N_20118,N_24077);
and UO_2448 (O_2448,N_20216,N_19320);
nand UO_2449 (O_2449,N_24870,N_23715);
nand UO_2450 (O_2450,N_23626,N_19803);
and UO_2451 (O_2451,N_20844,N_22237);
nor UO_2452 (O_2452,N_20416,N_19050);
and UO_2453 (O_2453,N_20264,N_24254);
nor UO_2454 (O_2454,N_20601,N_22120);
or UO_2455 (O_2455,N_20481,N_24743);
nand UO_2456 (O_2456,N_18932,N_22875);
xor UO_2457 (O_2457,N_19715,N_24943);
and UO_2458 (O_2458,N_20963,N_19708);
nor UO_2459 (O_2459,N_20016,N_23057);
or UO_2460 (O_2460,N_24988,N_23419);
xor UO_2461 (O_2461,N_24248,N_21904);
or UO_2462 (O_2462,N_21220,N_22483);
nor UO_2463 (O_2463,N_23298,N_21730);
nand UO_2464 (O_2464,N_24355,N_20309);
or UO_2465 (O_2465,N_23831,N_24230);
and UO_2466 (O_2466,N_24594,N_21441);
and UO_2467 (O_2467,N_18874,N_19414);
and UO_2468 (O_2468,N_19318,N_24921);
nand UO_2469 (O_2469,N_21415,N_24670);
nor UO_2470 (O_2470,N_21477,N_24385);
or UO_2471 (O_2471,N_20653,N_24081);
nand UO_2472 (O_2472,N_24453,N_23252);
nor UO_2473 (O_2473,N_22100,N_24808);
nand UO_2474 (O_2474,N_23911,N_19167);
and UO_2475 (O_2475,N_24717,N_19864);
nor UO_2476 (O_2476,N_23748,N_24760);
xor UO_2477 (O_2477,N_20271,N_20020);
or UO_2478 (O_2478,N_21319,N_21566);
and UO_2479 (O_2479,N_20485,N_23936);
and UO_2480 (O_2480,N_21821,N_18977);
and UO_2481 (O_2481,N_19437,N_20371);
nand UO_2482 (O_2482,N_23273,N_23015);
and UO_2483 (O_2483,N_24092,N_24497);
nor UO_2484 (O_2484,N_24939,N_24012);
nor UO_2485 (O_2485,N_21208,N_21270);
and UO_2486 (O_2486,N_22872,N_18822);
xnor UO_2487 (O_2487,N_20431,N_21668);
and UO_2488 (O_2488,N_22619,N_21076);
nor UO_2489 (O_2489,N_23857,N_22783);
nand UO_2490 (O_2490,N_23933,N_24784);
nand UO_2491 (O_2491,N_22105,N_19886);
nor UO_2492 (O_2492,N_24145,N_21962);
nand UO_2493 (O_2493,N_24710,N_23422);
nor UO_2494 (O_2494,N_22566,N_23937);
nand UO_2495 (O_2495,N_24991,N_23535);
and UO_2496 (O_2496,N_23797,N_20843);
nand UO_2497 (O_2497,N_21742,N_24168);
nor UO_2498 (O_2498,N_24733,N_19156);
nand UO_2499 (O_2499,N_19552,N_23854);
nor UO_2500 (O_2500,N_23175,N_24089);
and UO_2501 (O_2501,N_21278,N_21157);
or UO_2502 (O_2502,N_20274,N_19068);
or UO_2503 (O_2503,N_20695,N_19363);
or UO_2504 (O_2504,N_18831,N_20466);
xor UO_2505 (O_2505,N_24511,N_24127);
nand UO_2506 (O_2506,N_23248,N_20413);
and UO_2507 (O_2507,N_24895,N_21346);
nor UO_2508 (O_2508,N_18802,N_21972);
nand UO_2509 (O_2509,N_23694,N_21391);
and UO_2510 (O_2510,N_21618,N_19871);
nor UO_2511 (O_2511,N_22600,N_21859);
and UO_2512 (O_2512,N_22273,N_24366);
xnor UO_2513 (O_2513,N_21006,N_21465);
or UO_2514 (O_2514,N_21169,N_22132);
xor UO_2515 (O_2515,N_22850,N_18853);
nand UO_2516 (O_2516,N_18933,N_20388);
xor UO_2517 (O_2517,N_21681,N_20731);
nand UO_2518 (O_2518,N_22834,N_22645);
and UO_2519 (O_2519,N_24106,N_20681);
or UO_2520 (O_2520,N_22733,N_24313);
or UO_2521 (O_2521,N_24238,N_22119);
and UO_2522 (O_2522,N_19924,N_19209);
xnor UO_2523 (O_2523,N_19988,N_21568);
and UO_2524 (O_2524,N_22560,N_19205);
and UO_2525 (O_2525,N_19528,N_23385);
nand UO_2526 (O_2526,N_24071,N_22986);
xnor UO_2527 (O_2527,N_24342,N_23420);
or UO_2528 (O_2528,N_21901,N_20166);
or UO_2529 (O_2529,N_21440,N_24574);
nand UO_2530 (O_2530,N_21597,N_22282);
nand UO_2531 (O_2531,N_22364,N_19112);
nor UO_2532 (O_2532,N_21229,N_20874);
and UO_2533 (O_2533,N_22429,N_20191);
nand UO_2534 (O_2534,N_24123,N_18797);
and UO_2535 (O_2535,N_21439,N_23926);
nor UO_2536 (O_2536,N_22344,N_20295);
nor UO_2537 (O_2537,N_19124,N_22794);
or UO_2538 (O_2538,N_18940,N_21559);
and UO_2539 (O_2539,N_22574,N_24332);
nor UO_2540 (O_2540,N_23095,N_23277);
and UO_2541 (O_2541,N_19353,N_23201);
or UO_2542 (O_2542,N_23642,N_21089);
and UO_2543 (O_2543,N_24119,N_24442);
nand UO_2544 (O_2544,N_21680,N_22961);
and UO_2545 (O_2545,N_21252,N_24213);
and UO_2546 (O_2546,N_22400,N_18773);
xnor UO_2547 (O_2547,N_21102,N_20915);
xnor UO_2548 (O_2548,N_19020,N_23752);
or UO_2549 (O_2549,N_19270,N_24795);
nand UO_2550 (O_2550,N_19725,N_22820);
or UO_2551 (O_2551,N_21221,N_22497);
or UO_2552 (O_2552,N_22632,N_21131);
or UO_2553 (O_2553,N_22641,N_23311);
or UO_2554 (O_2554,N_24754,N_22391);
nand UO_2555 (O_2555,N_19939,N_24782);
nand UO_2556 (O_2556,N_20751,N_23575);
nor UO_2557 (O_2557,N_20741,N_18844);
nor UO_2558 (O_2558,N_21803,N_21914);
or UO_2559 (O_2559,N_18776,N_19129);
nand UO_2560 (O_2560,N_18875,N_19285);
nand UO_2561 (O_2561,N_19618,N_22878);
or UO_2562 (O_2562,N_22624,N_19224);
nor UO_2563 (O_2563,N_23221,N_23291);
or UO_2564 (O_2564,N_21141,N_23452);
or UO_2565 (O_2565,N_22550,N_24624);
or UO_2566 (O_2566,N_22540,N_20615);
nand UO_2567 (O_2567,N_22308,N_20564);
nor UO_2568 (O_2568,N_24426,N_22514);
nand UO_2569 (O_2569,N_24667,N_21268);
nand UO_2570 (O_2570,N_21437,N_19427);
and UO_2571 (O_2571,N_24564,N_19233);
and UO_2572 (O_2572,N_22705,N_19854);
and UO_2573 (O_2573,N_23441,N_19061);
nor UO_2574 (O_2574,N_21989,N_24159);
and UO_2575 (O_2575,N_24832,N_20815);
or UO_2576 (O_2576,N_19675,N_21775);
and UO_2577 (O_2577,N_21485,N_21843);
nand UO_2578 (O_2578,N_24538,N_19237);
or UO_2579 (O_2579,N_19727,N_19754);
or UO_2580 (O_2580,N_19122,N_19526);
xor UO_2581 (O_2581,N_21096,N_19612);
nor UO_2582 (O_2582,N_20339,N_22401);
nand UO_2583 (O_2583,N_20318,N_20036);
nor UO_2584 (O_2584,N_23461,N_21287);
nand UO_2585 (O_2585,N_22338,N_23777);
nand UO_2586 (O_2586,N_21373,N_22143);
nand UO_2587 (O_2587,N_21004,N_23913);
or UO_2588 (O_2588,N_21399,N_21545);
xnor UO_2589 (O_2589,N_24419,N_20169);
or UO_2590 (O_2590,N_24648,N_21140);
nor UO_2591 (O_2591,N_20317,N_20392);
nor UO_2592 (O_2592,N_23517,N_20503);
and UO_2593 (O_2593,N_24563,N_23064);
nand UO_2594 (O_2594,N_19074,N_22354);
nand UO_2595 (O_2595,N_19809,N_19140);
or UO_2596 (O_2596,N_20600,N_23279);
nor UO_2597 (O_2597,N_23669,N_21197);
or UO_2598 (O_2598,N_19097,N_24820);
or UO_2599 (O_2599,N_24736,N_24913);
xnor UO_2600 (O_2600,N_22511,N_24617);
and UO_2601 (O_2601,N_24959,N_23680);
nor UO_2602 (O_2602,N_22117,N_20616);
and UO_2603 (O_2603,N_23477,N_24529);
xor UO_2604 (O_2604,N_19375,N_24401);
and UO_2605 (O_2605,N_20334,N_21035);
nor UO_2606 (O_2606,N_22699,N_19196);
nor UO_2607 (O_2607,N_19495,N_19025);
xnor UO_2608 (O_2608,N_20581,N_19404);
nor UO_2609 (O_2609,N_21407,N_22146);
nor UO_2610 (O_2610,N_22174,N_21267);
or UO_2611 (O_2611,N_19183,N_18817);
nor UO_2612 (O_2612,N_19529,N_24431);
or UO_2613 (O_2613,N_21777,N_23011);
xor UO_2614 (O_2614,N_21887,N_24747);
and UO_2615 (O_2615,N_19491,N_21474);
and UO_2616 (O_2616,N_21063,N_19890);
and UO_2617 (O_2617,N_19204,N_21468);
nand UO_2618 (O_2618,N_24955,N_21889);
and UO_2619 (O_2619,N_19628,N_20790);
and UO_2620 (O_2620,N_18947,N_23401);
and UO_2621 (O_2621,N_23379,N_23843);
xnor UO_2622 (O_2622,N_22242,N_21612);
xnor UO_2623 (O_2623,N_20095,N_21099);
xor UO_2624 (O_2624,N_22075,N_24526);
nor UO_2625 (O_2625,N_19134,N_18911);
nor UO_2626 (O_2626,N_23150,N_24246);
nor UO_2627 (O_2627,N_24686,N_23309);
nor UO_2628 (O_2628,N_21101,N_20691);
xor UO_2629 (O_2629,N_18886,N_18820);
and UO_2630 (O_2630,N_20941,N_22335);
nand UO_2631 (O_2631,N_20246,N_22144);
or UO_2632 (O_2632,N_19390,N_22250);
or UO_2633 (O_2633,N_19816,N_24368);
nor UO_2634 (O_2634,N_20439,N_20688);
nand UO_2635 (O_2635,N_24031,N_20045);
or UO_2636 (O_2636,N_19637,N_20029);
and UO_2637 (O_2637,N_22093,N_20888);
nand UO_2638 (O_2638,N_21175,N_22644);
nand UO_2639 (O_2639,N_24414,N_23317);
or UO_2640 (O_2640,N_20743,N_21754);
or UO_2641 (O_2641,N_22894,N_20186);
nor UO_2642 (O_2642,N_23651,N_23496);
nand UO_2643 (O_2643,N_21104,N_21090);
nor UO_2644 (O_2644,N_19973,N_22471);
and UO_2645 (O_2645,N_19290,N_20959);
and UO_2646 (O_2646,N_20723,N_19855);
or UO_2647 (O_2647,N_22121,N_20530);
nor UO_2648 (O_2648,N_19407,N_23356);
or UO_2649 (O_2649,N_19688,N_23425);
or UO_2650 (O_2650,N_24791,N_21812);
nor UO_2651 (O_2651,N_22917,N_19297);
and UO_2652 (O_2652,N_19422,N_24780);
or UO_2653 (O_2653,N_22729,N_24627);
nand UO_2654 (O_2654,N_22869,N_20920);
or UO_2655 (O_2655,N_22972,N_21908);
or UO_2656 (O_2656,N_23769,N_24295);
nand UO_2657 (O_2657,N_23351,N_20745);
nand UO_2658 (O_2658,N_23712,N_20829);
and UO_2659 (O_2659,N_21038,N_24814);
nor UO_2660 (O_2660,N_22908,N_24958);
nand UO_2661 (O_2661,N_20989,N_23655);
nand UO_2662 (O_2662,N_23168,N_23783);
and UO_2663 (O_2663,N_19589,N_24361);
and UO_2664 (O_2664,N_23646,N_19702);
or UO_2665 (O_2665,N_21918,N_22084);
and UO_2666 (O_2666,N_20936,N_20952);
or UO_2667 (O_2667,N_22898,N_23380);
nor UO_2668 (O_2668,N_22111,N_20011);
nand UO_2669 (O_2669,N_20345,N_23183);
or UO_2670 (O_2670,N_24812,N_20065);
nor UO_2671 (O_2671,N_20467,N_19551);
or UO_2672 (O_2672,N_20819,N_20937);
and UO_2673 (O_2673,N_21272,N_19452);
or UO_2674 (O_2674,N_22922,N_22453);
and UO_2675 (O_2675,N_19227,N_24467);
nand UO_2676 (O_2676,N_18938,N_22828);
and UO_2677 (O_2677,N_22137,N_24752);
or UO_2678 (O_2678,N_23364,N_20405);
xor UO_2679 (O_2679,N_21956,N_23573);
xor UO_2680 (O_2680,N_21008,N_22602);
and UO_2681 (O_2681,N_22012,N_23848);
or UO_2682 (O_2682,N_19496,N_21571);
xor UO_2683 (O_2683,N_22030,N_19576);
and UO_2684 (O_2684,N_21786,N_20669);
nand UO_2685 (O_2685,N_19646,N_23218);
nor UO_2686 (O_2686,N_23389,N_24999);
nor UO_2687 (O_2687,N_23724,N_20866);
xnor UO_2688 (O_2688,N_19599,N_19887);
nand UO_2689 (O_2689,N_24562,N_23810);
xor UO_2690 (O_2690,N_24125,N_22067);
xor UO_2691 (O_2691,N_20774,N_21203);
or UO_2692 (O_2692,N_23985,N_23286);
and UO_2693 (O_2693,N_19305,N_21580);
or UO_2694 (O_2694,N_20256,N_20402);
nor UO_2695 (O_2695,N_21139,N_20634);
nor UO_2696 (O_2696,N_19663,N_20453);
xor UO_2697 (O_2697,N_21318,N_23403);
nor UO_2698 (O_2698,N_24949,N_22754);
and UO_2699 (O_2699,N_22518,N_19843);
or UO_2700 (O_2700,N_21062,N_23036);
and UO_2701 (O_2701,N_19254,N_22177);
and UO_2702 (O_2702,N_19219,N_22817);
nand UO_2703 (O_2703,N_21016,N_23928);
and UO_2704 (O_2704,N_19366,N_20734);
or UO_2705 (O_2705,N_19845,N_19941);
nor UO_2706 (O_2706,N_23446,N_20232);
and UO_2707 (O_2707,N_20557,N_23610);
nand UO_2708 (O_2708,N_21544,N_23809);
or UO_2709 (O_2709,N_23028,N_21517);
and UO_2710 (O_2710,N_22128,N_19598);
nor UO_2711 (O_2711,N_22685,N_24582);
xor UO_2712 (O_2712,N_19143,N_22897);
nor UO_2713 (O_2713,N_19400,N_23044);
nand UO_2714 (O_2714,N_19121,N_24509);
and UO_2715 (O_2715,N_21975,N_21515);
nor UO_2716 (O_2716,N_24661,N_21551);
nor UO_2717 (O_2717,N_24638,N_22303);
and UO_2718 (O_2718,N_21269,N_19720);
and UO_2719 (O_2719,N_23377,N_19453);
and UO_2720 (O_2720,N_20447,N_22123);
nor UO_2721 (O_2721,N_21853,N_19197);
xor UO_2722 (O_2722,N_20913,N_24819);
or UO_2723 (O_2723,N_20894,N_20621);
nor UO_2724 (O_2724,N_19980,N_22141);
and UO_2725 (O_2725,N_22785,N_21405);
nor UO_2726 (O_2726,N_20427,N_22928);
nor UO_2727 (O_2727,N_24911,N_23800);
xor UO_2728 (O_2728,N_20115,N_20778);
xnor UO_2729 (O_2729,N_19358,N_21529);
nand UO_2730 (O_2730,N_21428,N_22555);
nand UO_2731 (O_2731,N_21306,N_20306);
and UO_2732 (O_2732,N_23437,N_20845);
nor UO_2733 (O_2733,N_20154,N_23572);
or UO_2734 (O_2734,N_21335,N_23121);
nor UO_2735 (O_2735,N_23245,N_19750);
or UO_2736 (O_2736,N_24436,N_21522);
xor UO_2737 (O_2737,N_24032,N_21726);
nand UO_2738 (O_2738,N_22807,N_19146);
nand UO_2739 (O_2739,N_20228,N_23058);
and UO_2740 (O_2740,N_22852,N_24890);
nor UO_2741 (O_2741,N_21503,N_20940);
xor UO_2742 (O_2742,N_23865,N_22573);
nand UO_2743 (O_2743,N_21122,N_19438);
nand UO_2744 (O_2744,N_23561,N_24685);
nand UO_2745 (O_2745,N_20956,N_23846);
nand UO_2746 (O_2746,N_19471,N_18856);
and UO_2747 (O_2747,N_24144,N_24112);
and UO_2748 (O_2748,N_20452,N_19630);
or UO_2749 (O_2749,N_20426,N_22653);
nor UO_2750 (O_2750,N_20871,N_24673);
and UO_2751 (O_2751,N_23834,N_24508);
nand UO_2752 (O_2752,N_19289,N_21162);
and UO_2753 (O_2753,N_23767,N_19799);
nor UO_2754 (O_2754,N_22491,N_19699);
nand UO_2755 (O_2755,N_21414,N_20781);
xnor UO_2756 (O_2756,N_19015,N_18866);
and UO_2757 (O_2757,N_21994,N_21708);
nor UO_2758 (O_2758,N_19331,N_23952);
nor UO_2759 (O_2759,N_21170,N_22591);
or UO_2760 (O_2760,N_20969,N_20289);
xor UO_2761 (O_2761,N_20629,N_18755);
xor UO_2762 (O_2762,N_22206,N_24300);
nand UO_2763 (O_2763,N_21741,N_21712);
nand UO_2764 (O_2764,N_23557,N_23954);
and UO_2765 (O_2765,N_21168,N_18877);
and UO_2766 (O_2766,N_21355,N_23243);
or UO_2767 (O_2767,N_24944,N_20250);
nor UO_2768 (O_2768,N_21079,N_24912);
or UO_2769 (O_2769,N_22533,N_19357);
xnor UO_2770 (O_2770,N_21031,N_23835);
or UO_2771 (O_2771,N_22083,N_23050);
nor UO_2772 (O_2772,N_23445,N_19744);
nor UO_2773 (O_2773,N_20026,N_19264);
nand UO_2774 (O_2774,N_20369,N_21192);
nand UO_2775 (O_2775,N_24162,N_21686);
and UO_2776 (O_2776,N_19022,N_19786);
and UO_2777 (O_2777,N_18997,N_23060);
nor UO_2778 (O_2778,N_21737,N_19304);
nor UO_2779 (O_2779,N_24972,N_24158);
nand UO_2780 (O_2780,N_22742,N_23708);
nand UO_2781 (O_2781,N_21100,N_23444);
xor UO_2782 (O_2782,N_22343,N_21311);
nor UO_2783 (O_2783,N_23853,N_20809);
nand UO_2784 (O_2784,N_22633,N_21263);
nand UO_2785 (O_2785,N_19272,N_21920);
or UO_2786 (O_2786,N_19335,N_22487);
and UO_2787 (O_2787,N_23681,N_23624);
or UO_2788 (O_2788,N_21155,N_24885);
nand UO_2789 (O_2789,N_22062,N_21108);
and UO_2790 (O_2790,N_20771,N_22086);
nand UO_2791 (O_2791,N_20746,N_19672);
xnor UO_2792 (O_2792,N_24827,N_23796);
xor UO_2793 (O_2793,N_18751,N_20887);
and UO_2794 (O_2794,N_19171,N_24026);
nand UO_2795 (O_2795,N_18811,N_22339);
nand UO_2796 (O_2796,N_21828,N_22073);
nand UO_2797 (O_2797,N_20927,N_24682);
nand UO_2798 (O_2798,N_21291,N_21964);
and UO_2799 (O_2799,N_24948,N_24888);
or UO_2800 (O_2800,N_19028,N_21805);
nand UO_2801 (O_2801,N_19195,N_24862);
or UO_2802 (O_2802,N_23448,N_24995);
nand UO_2803 (O_2803,N_21622,N_19489);
and UO_2804 (O_2804,N_19723,N_24815);
and UO_2805 (O_2805,N_19041,N_23188);
nand UO_2806 (O_2806,N_24465,N_22730);
nand UO_2807 (O_2807,N_18919,N_21640);
nor UO_2808 (O_2808,N_23710,N_20838);
or UO_2809 (O_2809,N_24486,N_19899);
and UO_2810 (O_2810,N_20083,N_21749);
nor UO_2811 (O_2811,N_19667,N_22521);
or UO_2812 (O_2812,N_22474,N_22139);
nand UO_2813 (O_2813,N_20825,N_20793);
or UO_2814 (O_2814,N_23963,N_19690);
nor UO_2815 (O_2815,N_19392,N_20575);
nor UO_2816 (O_2816,N_20636,N_23451);
nor UO_2817 (O_2817,N_19211,N_19000);
and UO_2818 (O_2818,N_19773,N_23763);
and UO_2819 (O_2819,N_22976,N_23124);
or UO_2820 (O_2820,N_19057,N_23460);
and UO_2821 (O_2821,N_20833,N_19624);
nor UO_2822 (O_2822,N_19611,N_19132);
and UO_2823 (O_2823,N_21012,N_22559);
and UO_2824 (O_2824,N_21799,N_19044);
nand UO_2825 (O_2825,N_24513,N_20333);
and UO_2826 (O_2826,N_22231,N_22803);
and UO_2827 (O_2827,N_20222,N_20204);
or UO_2828 (O_2828,N_21025,N_24699);
or UO_2829 (O_2829,N_20430,N_18793);
nor UO_2830 (O_2830,N_18960,N_20820);
nor UO_2831 (O_2831,N_22579,N_19530);
and UO_2832 (O_2832,N_19048,N_18999);
nand UO_2833 (O_2833,N_19396,N_20133);
and UO_2834 (O_2834,N_22650,N_22452);
nor UO_2835 (O_2835,N_23333,N_21927);
or UO_2836 (O_2836,N_21472,N_23832);
xnor UO_2837 (O_2837,N_23790,N_23414);
and UO_2838 (O_2838,N_20206,N_19092);
nand UO_2839 (O_2839,N_19212,N_24229);
nor UO_2840 (O_2840,N_19955,N_24044);
or UO_2841 (O_2841,N_21285,N_22684);
nand UO_2842 (O_2842,N_23102,N_22604);
nand UO_2843 (O_2843,N_23841,N_22064);
and UO_2844 (O_2844,N_22190,N_24643);
nor UO_2845 (O_2845,N_21359,N_24846);
nand UO_2846 (O_2846,N_18991,N_21967);
nor UO_2847 (O_2847,N_22548,N_19566);
xnor UO_2848 (O_2848,N_23423,N_21673);
nor UO_2849 (O_2849,N_24148,N_20713);
or UO_2850 (O_2850,N_20648,N_22980);
xor UO_2851 (O_2851,N_21078,N_22876);
nor UO_2852 (O_2852,N_20791,N_22930);
or UO_2853 (O_2853,N_19283,N_21196);
and UO_2854 (O_2854,N_20406,N_21167);
nand UO_2855 (O_2855,N_20107,N_19711);
and UO_2856 (O_2856,N_19259,N_24521);
xor UO_2857 (O_2857,N_21623,N_20049);
nand UO_2858 (O_2858,N_22812,N_24263);
nand UO_2859 (O_2859,N_21427,N_23416);
nor UO_2860 (O_2860,N_24408,N_23815);
or UO_2861 (O_2861,N_23768,N_23961);
and UO_2862 (O_2862,N_23762,N_20626);
xnor UO_2863 (O_2863,N_22345,N_20276);
nor UO_2864 (O_2864,N_23336,N_24534);
nor UO_2865 (O_2865,N_23194,N_20571);
nor UO_2866 (O_2866,N_24380,N_24727);
nand UO_2867 (O_2867,N_19907,N_21868);
or UO_2868 (O_2868,N_24549,N_23504);
nor UO_2869 (O_2869,N_19818,N_19081);
nand UO_2870 (O_2870,N_23457,N_19812);
or UO_2871 (O_2871,N_24387,N_24593);
and UO_2872 (O_2872,N_20861,N_24020);
nand UO_2873 (O_2873,N_23638,N_23362);
and UO_2874 (O_2874,N_19659,N_23907);
nor UO_2875 (O_2875,N_22173,N_19860);
xor UO_2876 (O_2876,N_19652,N_22260);
xor UO_2877 (O_2877,N_21128,N_24228);
nor UO_2878 (O_2878,N_24879,N_21114);
nand UO_2879 (O_2879,N_24017,N_21588);
nor UO_2880 (O_2880,N_21781,N_21436);
nand UO_2881 (O_2881,N_19510,N_18859);
nand UO_2882 (O_2882,N_19508,N_21276);
and UO_2883 (O_2883,N_21854,N_21555);
and UO_2884 (O_2884,N_24143,N_24797);
and UO_2885 (O_2885,N_21628,N_21933);
nand UO_2886 (O_2886,N_23887,N_23436);
nand UO_2887 (O_2887,N_24553,N_21438);
nor UO_2888 (O_2888,N_23629,N_23676);
and UO_2889 (O_2889,N_21056,N_19983);
and UO_2890 (O_2890,N_21968,N_20462);
and UO_2891 (O_2891,N_18810,N_22045);
and UO_2892 (O_2892,N_23695,N_18951);
nand UO_2893 (O_2893,N_20227,N_20425);
xor UO_2894 (O_2894,N_20456,N_22832);
xnor UO_2895 (O_2895,N_23488,N_21410);
nor UO_2896 (O_2896,N_20382,N_24293);
or UO_2897 (O_2897,N_23497,N_19514);
or UO_2898 (O_2898,N_20391,N_24557);
nor UO_2899 (O_2899,N_24370,N_19160);
and UO_2900 (O_2900,N_20977,N_20475);
nor UO_2901 (O_2901,N_23882,N_24859);
nand UO_2902 (O_2902,N_18868,N_23805);
or UO_2903 (O_2903,N_22547,N_19088);
nor UO_2904 (O_2904,N_20813,N_21815);
nor UO_2905 (O_2905,N_24501,N_20308);
and UO_2906 (O_2906,N_24947,N_21315);
nand UO_2907 (O_2907,N_19226,N_22587);
and UO_2908 (O_2908,N_21043,N_19594);
or UO_2909 (O_2909,N_24930,N_23697);
or UO_2910 (O_2910,N_23230,N_20627);
or UO_2911 (O_2911,N_23434,N_19901);
or UO_2912 (O_2912,N_19747,N_20776);
nor UO_2913 (O_2913,N_24942,N_23265);
or UO_2914 (O_2914,N_23440,N_19620);
nor UO_2915 (O_2915,N_18905,N_23391);
or UO_2916 (O_2916,N_20484,N_20071);
or UO_2917 (O_2917,N_24432,N_19696);
nor UO_2918 (O_2918,N_22557,N_22957);
nand UO_2919 (O_2919,N_21832,N_20711);
or UO_2920 (O_2920,N_19946,N_23559);
xor UO_2921 (O_2921,N_22243,N_21556);
nand UO_2922 (O_2922,N_22797,N_21876);
xnor UO_2923 (O_2923,N_21172,N_23435);
nand UO_2924 (O_2924,N_20739,N_22000);
nor UO_2925 (O_2925,N_21010,N_19557);
or UO_2926 (O_2926,N_19963,N_24666);
and UO_2927 (O_2927,N_19077,N_24505);
nor UO_2928 (O_2928,N_22610,N_20393);
nand UO_2929 (O_2929,N_21029,N_22044);
or UO_2930 (O_2930,N_20344,N_20088);
nand UO_2931 (O_2931,N_21300,N_20175);
nand UO_2932 (O_2932,N_20200,N_18864);
xnor UO_2933 (O_2933,N_21760,N_23635);
nor UO_2934 (O_2934,N_22929,N_18899);
xor UO_2935 (O_2935,N_24657,N_23773);
nor UO_2936 (O_2936,N_21204,N_19278);
nor UO_2937 (O_2937,N_23305,N_21446);
and UO_2938 (O_2938,N_22433,N_23163);
nor UO_2939 (O_2939,N_23081,N_22278);
and UO_2940 (O_2940,N_24057,N_19908);
or UO_2941 (O_2941,N_21850,N_24873);
nand UO_2942 (O_2942,N_24701,N_23395);
nand UO_2943 (O_2943,N_24933,N_19159);
or UO_2944 (O_2944,N_19761,N_20202);
or UO_2945 (O_2945,N_24898,N_23647);
nor UO_2946 (O_2946,N_21317,N_22770);
nand UO_2947 (O_2947,N_23111,N_21443);
or UO_2948 (O_2948,N_21534,N_23842);
or UO_2949 (O_2949,N_22966,N_22162);
nor UO_2950 (O_2950,N_24504,N_19388);
and UO_2951 (O_2951,N_21486,N_21776);
nand UO_2952 (O_2952,N_22732,N_24205);
and UO_2953 (O_2953,N_22711,N_22925);
or UO_2954 (O_2954,N_23272,N_22938);
and UO_2955 (O_2955,N_22395,N_21753);
and UO_2956 (O_2956,N_22892,N_21945);
and UO_2957 (O_2957,N_23514,N_23171);
xnor UO_2958 (O_2958,N_24525,N_20849);
nand UO_2959 (O_2959,N_22053,N_23953);
and UO_2960 (O_2960,N_23645,N_23306);
and UO_2961 (O_2961,N_24455,N_21636);
xor UO_2962 (O_2962,N_19457,N_19852);
and UO_2963 (O_2963,N_24222,N_19960);
nand UO_2964 (O_2964,N_20902,N_23729);
nand UO_2965 (O_2965,N_21676,N_21387);
or UO_2966 (O_2966,N_23318,N_21881);
nand UO_2967 (O_2967,N_20549,N_22575);
xnor UO_2968 (O_2968,N_21802,N_24700);
xor UO_2969 (O_2969,N_22762,N_19389);
or UO_2970 (O_2970,N_24036,N_19341);
or UO_2971 (O_2971,N_21573,N_20684);
and UO_2972 (O_2972,N_23513,N_22669);
and UO_2973 (O_2973,N_23085,N_24896);
and UO_2974 (O_2974,N_24615,N_20441);
nor UO_2975 (O_2975,N_19561,N_19506);
or UO_2976 (O_2976,N_24856,N_22556);
nor UO_2977 (O_2977,N_24929,N_23074);
and UO_2978 (O_2978,N_20042,N_21855);
xnor UO_2979 (O_2979,N_23223,N_22133);
xor UO_2980 (O_2980,N_21152,N_20380);
xnor UO_2981 (O_2981,N_24374,N_22895);
or UO_2982 (O_2982,N_20367,N_24647);
nand UO_2983 (O_2983,N_22631,N_18882);
nand UO_2984 (O_2984,N_24683,N_18935);
nor UO_2985 (O_2985,N_20520,N_22623);
or UO_2986 (O_2986,N_22363,N_20709);
or UO_2987 (O_2987,N_21160,N_22616);
xor UO_2988 (O_2988,N_20242,N_20699);
nand UO_2989 (O_2989,N_23615,N_19001);
and UO_2990 (O_2990,N_20501,N_21660);
and UO_2991 (O_2991,N_22656,N_20455);
nor UO_2992 (O_2992,N_20765,N_20196);
or UO_2993 (O_2993,N_23755,N_22388);
and UO_2994 (O_2994,N_21461,N_20150);
and UO_2995 (O_2995,N_21954,N_22436);
nand UO_2996 (O_2996,N_22577,N_23673);
xnor UO_2997 (O_2997,N_23185,N_22148);
and UO_2998 (O_2998,N_20487,N_22597);
and UO_2999 (O_2999,N_24157,N_20824);
endmodule