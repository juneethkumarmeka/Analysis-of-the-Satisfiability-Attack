module basic_2000_20000_2500_10_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
xor U0 (N_0,In_1803,In_165);
and U1 (N_1,In_1213,In_968);
nor U2 (N_2,In_1795,In_1839);
nand U3 (N_3,In_1021,In_738);
or U4 (N_4,In_112,In_660);
nand U5 (N_5,In_78,In_1154);
nor U6 (N_6,In_1541,In_847);
xor U7 (N_7,In_1333,In_1511);
and U8 (N_8,In_525,In_1435);
and U9 (N_9,In_640,In_1480);
nor U10 (N_10,In_923,In_1892);
nand U11 (N_11,In_54,In_7);
and U12 (N_12,In_1761,In_1450);
nor U13 (N_13,In_427,In_1764);
nor U14 (N_14,In_59,In_792);
and U15 (N_15,In_79,In_1935);
nand U16 (N_16,In_388,In_1703);
and U17 (N_17,In_672,In_295);
and U18 (N_18,In_906,In_551);
nor U19 (N_19,In_948,In_69);
nand U20 (N_20,In_304,In_440);
nor U21 (N_21,In_908,In_210);
xor U22 (N_22,In_93,In_396);
nor U23 (N_23,In_1594,In_721);
and U24 (N_24,In_285,In_1693);
or U25 (N_25,In_580,In_29);
xnor U26 (N_26,In_113,In_1147);
xor U27 (N_27,In_24,In_674);
and U28 (N_28,In_174,In_1269);
or U29 (N_29,In_1775,In_586);
nor U30 (N_30,In_1349,In_1714);
nor U31 (N_31,In_911,In_357);
and U32 (N_32,In_1730,In_1842);
or U33 (N_33,In_279,In_1262);
xnor U34 (N_34,In_1891,In_766);
xnor U35 (N_35,In_1265,In_1477);
xor U36 (N_36,In_362,In_412);
nor U37 (N_37,In_498,In_1978);
or U38 (N_38,In_882,In_1276);
nand U39 (N_39,In_497,In_1448);
or U40 (N_40,In_1157,In_1417);
nand U41 (N_41,In_269,In_1883);
or U42 (N_42,In_550,In_1385);
nand U43 (N_43,In_1325,In_306);
nand U44 (N_44,In_715,In_592);
nand U45 (N_45,In_869,In_1034);
nor U46 (N_46,In_596,In_1672);
xor U47 (N_47,In_1826,In_316);
nand U48 (N_48,In_978,In_938);
nor U49 (N_49,In_1521,In_961);
nand U50 (N_50,In_934,In_1704);
and U51 (N_51,In_1944,In_56);
or U52 (N_52,In_670,In_191);
xor U53 (N_53,In_562,In_940);
or U54 (N_54,In_1994,In_1425);
and U55 (N_55,In_1355,In_103);
nand U56 (N_56,In_53,In_1732);
or U57 (N_57,In_1872,In_237);
or U58 (N_58,In_259,In_1763);
or U59 (N_59,In_98,In_1148);
xnor U60 (N_60,In_1811,In_1231);
nor U61 (N_61,In_927,In_1837);
nor U62 (N_62,In_99,In_190);
nand U63 (N_63,In_1848,In_1382);
xnor U64 (N_64,In_599,In_251);
xor U65 (N_65,In_1913,In_514);
and U66 (N_66,In_1652,In_1311);
or U67 (N_67,In_778,In_1131);
xnor U68 (N_68,In_1018,In_1838);
or U69 (N_69,In_1215,In_390);
or U70 (N_70,In_1182,In_662);
xnor U71 (N_71,In_1739,In_1694);
nand U72 (N_72,In_233,In_104);
nor U73 (N_73,In_181,In_1044);
nor U74 (N_74,In_1907,In_506);
or U75 (N_75,In_1785,In_816);
or U76 (N_76,In_1023,In_166);
nand U77 (N_77,In_1248,In_613);
nand U78 (N_78,In_432,In_39);
nand U79 (N_79,In_1646,In_762);
nor U80 (N_80,In_408,In_384);
and U81 (N_81,In_128,In_712);
nor U82 (N_82,In_1643,In_1045);
and U83 (N_83,In_1183,In_1239);
and U84 (N_84,In_101,In_433);
or U85 (N_85,In_773,In_1705);
or U86 (N_86,In_1595,In_1356);
nand U87 (N_87,In_1606,In_1484);
and U88 (N_88,In_323,In_667);
nor U89 (N_89,In_783,In_1386);
xor U90 (N_90,In_548,In_1257);
or U91 (N_91,In_569,In_235);
or U92 (N_92,In_1960,In_561);
xnor U93 (N_93,In_1936,In_929);
nand U94 (N_94,In_280,In_1568);
nor U95 (N_95,In_240,In_1315);
and U96 (N_96,In_468,In_1323);
xor U97 (N_97,In_294,In_266);
nand U98 (N_98,In_1874,In_886);
xnor U99 (N_99,In_921,In_1189);
and U100 (N_100,In_1106,In_1104);
nor U101 (N_101,In_1982,In_1895);
or U102 (N_102,In_696,In_168);
nand U103 (N_103,In_889,In_593);
xor U104 (N_104,In_1490,In_8);
or U105 (N_105,In_770,In_695);
and U106 (N_106,In_189,In_392);
nand U107 (N_107,In_1716,In_1937);
and U108 (N_108,In_977,In_1181);
nand U109 (N_109,In_1979,In_275);
nor U110 (N_110,In_92,In_589);
nand U111 (N_111,In_1039,In_1105);
xor U112 (N_112,In_1669,In_22);
nor U113 (N_113,In_154,In_1140);
nor U114 (N_114,In_1667,In_1992);
nor U115 (N_115,In_1436,In_239);
nor U116 (N_116,In_804,In_1923);
xor U117 (N_117,In_1125,In_1049);
nand U118 (N_118,In_900,In_60);
xor U119 (N_119,In_1778,In_661);
nor U120 (N_120,In_1861,In_305);
and U121 (N_121,In_499,In_1514);
or U122 (N_122,In_677,In_1787);
nor U123 (N_123,In_1799,In_1458);
or U124 (N_124,In_182,In_504);
or U125 (N_125,In_1564,In_126);
nor U126 (N_126,In_606,In_187);
xnor U127 (N_127,In_833,In_1136);
nor U128 (N_128,In_331,In_322);
and U129 (N_129,In_1881,In_332);
and U130 (N_130,In_1101,In_1073);
nand U131 (N_131,In_105,In_997);
nor U132 (N_132,In_834,In_1142);
nor U133 (N_133,In_710,In_1614);
or U134 (N_134,In_884,In_1590);
or U135 (N_135,In_650,In_207);
or U136 (N_136,In_693,In_1917);
nand U137 (N_137,In_1472,In_625);
xor U138 (N_138,In_1567,In_1440);
and U139 (N_139,In_1378,In_1958);
xor U140 (N_140,In_1933,In_1320);
or U141 (N_141,In_480,In_1807);
nand U142 (N_142,In_888,In_1699);
and U143 (N_143,In_1988,In_519);
and U144 (N_144,In_576,In_1242);
xnor U145 (N_145,In_733,In_1662);
nor U146 (N_146,In_857,In_1321);
xnor U147 (N_147,In_754,In_27);
or U148 (N_148,In_1855,In_784);
xnor U149 (N_149,In_986,In_1942);
or U150 (N_150,In_1274,In_974);
nor U151 (N_151,In_102,In_996);
nand U152 (N_152,In_799,In_526);
nand U153 (N_153,In_198,In_1095);
xnor U154 (N_154,In_35,In_345);
nor U155 (N_155,In_355,In_1768);
nand U156 (N_156,In_871,In_1893);
xor U157 (N_157,In_86,In_1814);
nor U158 (N_158,In_1038,In_585);
or U159 (N_159,In_564,In_813);
nor U160 (N_160,In_1040,In_1439);
nand U161 (N_161,In_1746,In_1585);
or U162 (N_162,In_1919,In_1530);
and U163 (N_163,In_641,In_646);
xor U164 (N_164,In_363,In_750);
xor U165 (N_165,In_1240,In_1486);
nor U166 (N_166,In_1586,In_1075);
nand U167 (N_167,In_920,In_1433);
nand U168 (N_168,In_907,In_1540);
nand U169 (N_169,In_591,In_638);
and U170 (N_170,In_1020,In_1451);
nand U171 (N_171,In_971,In_916);
and U172 (N_172,In_1901,In_607);
nor U173 (N_173,In_1307,In_462);
nor U174 (N_174,In_1805,In_767);
or U175 (N_175,In_628,In_1343);
nor U176 (N_176,In_310,In_10);
or U177 (N_177,In_829,In_1178);
xor U178 (N_178,In_1835,In_698);
xnor U179 (N_179,In_1275,In_314);
xor U180 (N_180,In_1870,In_1903);
and U181 (N_181,In_1267,In_1229);
xor U182 (N_182,In_1012,In_897);
or U183 (N_183,In_1492,In_666);
nand U184 (N_184,In_1645,In_1670);
or U185 (N_185,In_1469,In_990);
or U186 (N_186,In_220,In_885);
nor U187 (N_187,In_846,In_481);
nand U188 (N_188,In_966,In_1843);
or U189 (N_189,In_287,In_425);
nand U190 (N_190,In_219,In_1666);
nand U191 (N_191,In_116,In_124);
and U192 (N_192,In_1200,In_48);
and U193 (N_193,In_547,In_64);
xor U194 (N_194,In_361,In_1909);
xor U195 (N_195,In_236,In_1352);
or U196 (N_196,In_1818,In_450);
nand U197 (N_197,In_1427,In_1447);
nor U198 (N_198,In_1896,In_1951);
or U199 (N_199,In_1299,In_901);
and U200 (N_200,In_111,In_0);
nand U201 (N_201,In_1060,In_1547);
xnor U202 (N_202,In_680,In_1802);
xnor U203 (N_203,In_204,In_16);
xnor U204 (N_204,In_577,In_1186);
nor U205 (N_205,In_457,In_837);
xnor U206 (N_206,In_1711,In_1364);
nand U207 (N_207,In_1798,In_341);
xor U208 (N_208,In_1428,In_1264);
nand U209 (N_209,In_87,In_651);
nor U210 (N_210,In_820,In_1007);
or U211 (N_211,In_228,In_1583);
and U212 (N_212,In_300,In_1792);
nand U213 (N_213,In_1036,In_171);
or U214 (N_214,In_1285,In_609);
nand U215 (N_215,In_398,In_373);
and U216 (N_216,In_617,In_702);
or U217 (N_217,In_213,In_1770);
nand U218 (N_218,In_484,In_271);
nor U219 (N_219,In_23,In_129);
and U220 (N_220,In_1324,In_1389);
nor U221 (N_221,In_1615,In_226);
or U222 (N_222,In_1487,In_937);
xnor U223 (N_223,In_1150,In_511);
xnor U224 (N_224,In_470,In_153);
or U225 (N_225,In_368,In_1420);
nand U226 (N_226,In_426,In_394);
and U227 (N_227,In_309,In_1756);
and U228 (N_228,In_1121,In_1680);
xor U229 (N_229,In_528,In_467);
nor U230 (N_230,In_708,In_512);
xnor U231 (N_231,In_824,In_1743);
nand U232 (N_232,In_659,In_386);
and U233 (N_233,In_1434,In_1537);
and U234 (N_234,In_771,In_735);
or U235 (N_235,In_616,In_299);
or U236 (N_236,In_1237,In_1931);
or U237 (N_237,In_896,In_1661);
xnor U238 (N_238,In_337,In_1969);
xnor U239 (N_239,In_1072,In_1123);
xnor U240 (N_240,In_270,In_1441);
nor U241 (N_241,In_701,In_1784);
or U242 (N_242,In_556,In_1097);
nor U243 (N_243,In_730,In_1681);
xnor U244 (N_244,In_546,In_1216);
or U245 (N_245,In_380,In_1372);
and U246 (N_246,In_434,In_1501);
nor U247 (N_247,In_1862,In_1729);
or U248 (N_248,In_1185,In_1735);
and U249 (N_249,In_687,In_803);
xor U250 (N_250,In_438,In_1491);
or U251 (N_251,In_873,In_472);
nor U252 (N_252,In_1526,In_1688);
nand U253 (N_253,In_186,In_21);
xor U254 (N_254,In_568,In_620);
nand U255 (N_255,In_465,In_1042);
xor U256 (N_256,In_1461,In_1227);
nand U257 (N_257,In_72,In_673);
and U258 (N_258,In_1103,In_37);
and U259 (N_259,In_1980,In_1793);
xnor U260 (N_260,In_830,In_981);
nor U261 (N_261,In_1945,In_1630);
nor U262 (N_262,In_1513,In_1574);
nand U263 (N_263,In_1999,In_880);
nor U264 (N_264,In_1347,In_953);
or U265 (N_265,In_1952,In_1745);
or U266 (N_266,In_178,In_1579);
and U267 (N_267,In_1241,In_1391);
xor U268 (N_268,In_571,In_789);
nand U269 (N_269,In_1809,In_892);
and U270 (N_270,In_1011,In_303);
xnor U271 (N_271,In_1317,In_1889);
xnor U272 (N_272,In_1297,In_1258);
nand U273 (N_273,In_1119,In_1555);
xor U274 (N_274,In_1904,In_570);
xor U275 (N_275,In_150,In_283);
xnor U276 (N_276,In_1359,In_1174);
xnor U277 (N_277,In_274,In_273);
xnor U278 (N_278,In_1902,In_52);
xor U279 (N_279,In_1731,In_755);
nand U280 (N_280,In_1354,In_1210);
and U281 (N_281,In_1986,In_243);
nand U282 (N_282,In_893,In_486);
and U283 (N_283,In_1709,In_567);
xnor U284 (N_284,In_1550,In_898);
nand U285 (N_285,In_419,In_841);
nand U286 (N_286,In_1518,In_1362);
xnor U287 (N_287,In_878,In_1760);
nand U288 (N_288,In_1642,In_594);
nor U289 (N_289,In_1723,In_1528);
nor U290 (N_290,In_531,In_1462);
nand U291 (N_291,In_6,In_939);
nor U292 (N_292,In_1525,In_1207);
xor U293 (N_293,In_1871,In_1532);
xnor U294 (N_294,In_130,In_336);
nand U295 (N_295,In_402,In_1908);
xnor U296 (N_296,In_1975,In_925);
nor U297 (N_297,In_214,In_679);
or U298 (N_298,In_1673,In_705);
nor U299 (N_299,In_552,In_1520);
and U300 (N_300,In_1411,In_1758);
nor U301 (N_301,In_1742,In_1399);
nor U302 (N_302,In_1914,In_1940);
nor U303 (N_303,In_1538,In_955);
nand U304 (N_304,In_964,In_119);
or U305 (N_305,In_579,In_1234);
nand U306 (N_306,In_876,In_1067);
and U307 (N_307,In_1054,In_1092);
xnor U308 (N_308,In_395,In_658);
and U309 (N_309,In_1946,In_216);
or U310 (N_310,In_933,In_38);
and U311 (N_311,In_618,In_1310);
and U312 (N_312,In_464,In_1845);
or U313 (N_313,In_1636,In_706);
xnor U314 (N_314,In_867,In_1022);
xor U315 (N_315,In_232,In_1668);
nand U316 (N_316,In_572,In_418);
nor U317 (N_317,In_1406,In_265);
and U318 (N_318,In_1519,In_1050);
xor U319 (N_319,In_615,In_1863);
and U320 (N_320,In_167,In_1651);
nand U321 (N_321,In_994,In_671);
xnor U322 (N_322,In_769,In_1459);
and U323 (N_323,In_1465,In_1719);
xor U324 (N_324,In_941,In_1212);
or U325 (N_325,In_1198,In_1118);
xnor U326 (N_326,In_447,In_1345);
nor U327 (N_327,In_263,In_1314);
or U328 (N_328,In_1612,In_1812);
and U329 (N_329,In_951,In_1443);
and U330 (N_330,In_991,In_1222);
or U331 (N_331,In_1987,In_713);
xnor U332 (N_332,In_611,In_491);
and U333 (N_333,In_110,In_1383);
and U334 (N_334,In_522,In_381);
and U335 (N_335,In_1013,In_1397);
and U336 (N_336,In_1085,In_1536);
and U337 (N_337,In_714,In_1808);
and U338 (N_338,In_918,In_1404);
nor U339 (N_339,In_808,In_560);
and U340 (N_340,In_652,In_1145);
and U341 (N_341,In_980,In_121);
or U342 (N_342,In_1989,In_183);
xor U343 (N_343,In_453,In_172);
or U344 (N_344,In_1094,In_1588);
or U345 (N_345,In_1569,In_377);
nand U346 (N_346,In_500,In_1962);
nand U347 (N_347,In_765,In_151);
or U348 (N_348,In_970,In_1079);
nand U349 (N_349,In_746,In_318);
nor U350 (N_350,In_844,In_1081);
xor U351 (N_351,In_1272,In_1801);
or U352 (N_352,In_1153,In_812);
nor U353 (N_353,In_1164,In_372);
nor U354 (N_354,In_1080,In_642);
or U355 (N_355,In_744,In_145);
nand U356 (N_356,In_1332,In_209);
nand U357 (N_357,In_517,In_1852);
nand U358 (N_358,In_791,In_1063);
nor U359 (N_359,In_1571,In_1941);
or U360 (N_360,In_1375,In_1309);
xnor U361 (N_361,In_647,In_452);
and U362 (N_362,In_643,In_819);
or U363 (N_363,In_975,In_1707);
and U364 (N_364,In_421,In_1995);
or U365 (N_365,In_1771,In_62);
xnor U366 (N_366,In_148,In_1246);
nor U367 (N_367,In_720,In_65);
or U368 (N_368,In_946,In_1306);
or U369 (N_369,In_262,In_523);
or U370 (N_370,In_1794,In_1850);
xor U371 (N_371,In_1266,In_1713);
nor U372 (N_372,In_930,In_320);
xor U373 (N_373,In_875,In_903);
xor U374 (N_374,In_170,In_1090);
xor U375 (N_375,In_1622,In_1948);
nand U376 (N_376,In_1757,In_1985);
nor U377 (N_377,In_890,In_790);
and U378 (N_378,In_222,In_751);
and U379 (N_379,In_1625,In_854);
nor U380 (N_380,In_383,In_482);
nor U381 (N_381,In_1584,In_1312);
nand U382 (N_382,In_33,In_193);
xnor U383 (N_383,In_1689,In_1899);
nor U384 (N_384,In_1506,In_1128);
xnor U385 (N_385,In_1194,In_1083);
nor U386 (N_386,In_760,In_1875);
and U387 (N_387,In_1500,In_1750);
xnor U388 (N_388,In_774,In_489);
nand U389 (N_389,In_327,In_1495);
or U390 (N_390,In_297,In_249);
and U391 (N_391,In_1344,In_158);
and U392 (N_392,In_1048,In_1452);
nand U393 (N_393,In_1602,In_135);
or U394 (N_394,In_1442,In_725);
nor U395 (N_395,In_107,In_1419);
xnor U396 (N_396,In_1720,In_218);
nor U397 (N_397,In_1014,In_1331);
nand U398 (N_398,In_95,In_1533);
nor U399 (N_399,In_1170,In_728);
nand U400 (N_400,In_308,In_43);
xnor U401 (N_401,In_1296,In_973);
xnor U402 (N_402,In_1172,In_1833);
nand U403 (N_403,In_2,In_1762);
nand U404 (N_404,In_1357,In_328);
or U405 (N_405,In_818,In_1912);
nor U406 (N_406,In_379,In_1927);
xor U407 (N_407,In_1984,In_224);
nor U408 (N_408,In_1570,In_1557);
nor U409 (N_409,In_1456,In_1820);
xnor U410 (N_410,In_1139,In_775);
and U411 (N_411,In_399,In_1086);
and U412 (N_412,In_284,In_215);
nor U413 (N_413,In_635,In_741);
or U414 (N_414,In_1233,In_1592);
xor U415 (N_415,In_753,In_413);
nand U416 (N_416,In_723,In_238);
or U417 (N_417,In_339,In_370);
and U418 (N_418,In_1336,In_1607);
or U419 (N_419,In_1634,In_1910);
xnor U420 (N_420,In_205,In_1744);
or U421 (N_421,In_45,In_1846);
nor U422 (N_422,In_1407,In_1560);
or U423 (N_423,In_1016,In_1259);
nand U424 (N_424,In_208,In_1414);
and U425 (N_425,In_1611,In_1836);
and U426 (N_426,In_1395,In_147);
and U427 (N_427,In_922,In_231);
nor U428 (N_428,In_1410,In_144);
nor U429 (N_429,In_1777,In_473);
and U430 (N_430,In_1639,In_632);
nor U431 (N_431,In_1260,In_1544);
nor U432 (N_432,In_1496,In_836);
xor U433 (N_433,In_1074,In_724);
and U434 (N_434,In_1658,In_123);
nor U435 (N_435,In_88,In_315);
and U436 (N_436,In_338,In_66);
xnor U437 (N_437,In_1619,In_1939);
nor U438 (N_438,In_949,In_477);
nand U439 (N_439,In_805,In_1387);
nor U440 (N_440,In_1865,In_1091);
nand U441 (N_441,In_1338,In_405);
or U442 (N_442,In_1499,In_324);
xnor U443 (N_443,In_1059,In_127);
or U444 (N_444,In_1632,In_230);
nor U445 (N_445,In_669,In_505);
xnor U446 (N_446,In_1286,In_1159);
xor U447 (N_447,In_956,In_1244);
and U448 (N_448,In_1392,In_1817);
nand U449 (N_449,In_689,In_1654);
nor U450 (N_450,In_1149,In_538);
nand U451 (N_451,In_1078,In_827);
nand U452 (N_452,In_764,In_1202);
nor U453 (N_453,In_623,In_1726);
nor U454 (N_454,In_347,In_629);
and U455 (N_455,In_1868,In_1379);
xnor U456 (N_456,In_106,In_801);
nand U457 (N_457,In_325,In_456);
nor U458 (N_458,In_335,In_832);
xnor U459 (N_459,In_1279,In_1460);
nand U460 (N_460,In_1796,In_759);
and U461 (N_461,In_1656,In_727);
nor U462 (N_462,In_581,In_268);
xor U463 (N_463,In_1476,In_518);
xor U464 (N_464,In_329,In_802);
nand U465 (N_465,In_1273,In_437);
nand U466 (N_466,In_1466,In_1653);
and U467 (N_467,In_601,In_861);
or U468 (N_468,In_1116,In_1997);
xor U469 (N_469,In_1640,In_36);
or U470 (N_470,In_967,In_192);
nand U471 (N_471,In_358,In_1717);
xnor U472 (N_472,In_863,In_301);
or U473 (N_473,In_1188,In_1618);
xnor U474 (N_474,In_1193,In_1566);
nor U475 (N_475,In_637,In_296);
nor U476 (N_476,In_1915,In_959);
and U477 (N_477,In_1000,In_1576);
or U478 (N_478,In_1373,In_400);
xnor U479 (N_479,In_1291,In_699);
nand U480 (N_480,In_1886,In_1696);
and U481 (N_481,In_602,In_1381);
nand U482 (N_482,In_47,In_619);
nand U483 (N_483,In_1367,In_902);
nand U484 (N_484,In_343,In_866);
xor U485 (N_485,In_1337,In_449);
or U486 (N_486,In_359,In_1334);
xor U487 (N_487,In_777,In_469);
nor U488 (N_488,In_267,In_555);
and U489 (N_489,In_1629,In_1575);
xnor U490 (N_490,In_1829,In_1813);
or U491 (N_491,In_80,In_747);
xor U492 (N_492,In_1449,In_82);
nand U493 (N_493,In_1675,In_1431);
nor U494 (N_494,In_1191,In_354);
nor U495 (N_495,In_681,In_429);
and U496 (N_496,In_688,In_1374);
and U497 (N_497,In_1089,In_1024);
xor U498 (N_498,In_826,In_371);
xnor U499 (N_499,In_411,In_1691);
nor U500 (N_500,In_18,In_71);
xor U501 (N_501,In_1099,In_726);
nor U502 (N_502,In_155,In_1204);
and U503 (N_503,In_256,In_1162);
nand U504 (N_504,In_845,In_1884);
and U505 (N_505,In_1287,In_391);
nand U506 (N_506,In_794,In_1218);
nand U507 (N_507,In_1376,In_1676);
nor U508 (N_508,In_1252,In_57);
or U509 (N_509,In_1955,In_965);
xnor U510 (N_510,In_255,In_118);
or U511 (N_511,In_534,In_1076);
and U512 (N_512,In_626,In_1593);
nor U513 (N_513,In_133,In_1815);
or U514 (N_514,In_1069,In_1350);
or U515 (N_515,In_1028,In_731);
or U516 (N_516,In_485,In_333);
xor U517 (N_517,In_156,In_1553);
and U518 (N_518,In_554,In_1082);
nor U519 (N_519,In_874,In_1957);
or U520 (N_520,In_1482,In_954);
nor U521 (N_521,In_958,In_1608);
xnor U522 (N_522,In_1780,In_645);
or U523 (N_523,In_446,In_1192);
nor U524 (N_524,In_159,In_1300);
nand U525 (N_525,In_634,In_1277);
and U526 (N_526,In_1905,In_1328);
xnor U527 (N_527,In_1316,In_272);
nor U528 (N_528,In_188,In_758);
nor U529 (N_529,In_474,In_1245);
and U530 (N_530,In_950,In_1424);
nor U531 (N_531,In_1545,In_1747);
xnor U532 (N_532,In_1208,In_1464);
nor U533 (N_533,In_1722,In_1064);
nor U534 (N_534,In_840,In_756);
or U535 (N_535,In_807,In_1686);
nor U536 (N_536,In_1885,In_657);
nor U537 (N_537,In_1413,In_860);
and U538 (N_538,In_545,In_140);
nor U539 (N_539,In_1779,In_229);
nand U540 (N_540,In_120,In_1130);
nand U541 (N_541,In_1924,In_385);
and U542 (N_542,In_584,In_50);
nor U543 (N_543,In_1152,In_73);
or U544 (N_544,In_169,In_743);
or U545 (N_545,In_1515,In_463);
and U546 (N_546,In_1236,In_1494);
nor U547 (N_547,In_1834,In_1644);
or U548 (N_548,In_1765,In_1998);
or U549 (N_549,In_1173,In_1769);
xnor U550 (N_550,In_1341,In_459);
xnor U551 (N_551,In_1479,In_828);
nor U552 (N_552,In_67,In_1754);
or U553 (N_553,In_1598,In_4);
xnor U554 (N_554,In_422,In_1037);
or U555 (N_555,In_1683,In_839);
xnor U556 (N_556,In_1114,In_122);
xor U557 (N_557,In_31,In_1353);
or U558 (N_558,In_1056,In_1580);
nand U559 (N_559,In_404,In_565);
nand U560 (N_560,In_1554,In_895);
nand U561 (N_561,In_1888,In_524);
and U562 (N_562,In_353,In_984);
or U563 (N_563,In_1171,In_1217);
or U564 (N_564,In_821,In_352);
xnor U565 (N_565,In_1841,In_369);
and U566 (N_566,In_654,In_1562);
nor U567 (N_567,In_443,In_417);
and U568 (N_568,In_772,In_800);
and U569 (N_569,In_1953,In_1284);
nand U570 (N_570,In_1361,In_389);
nand U571 (N_571,In_1363,In_1168);
or U572 (N_572,In_1949,In_1702);
nor U573 (N_573,In_58,In_117);
nor U574 (N_574,In_879,In_703);
or U575 (N_575,In_1721,In_1096);
nand U576 (N_576,In_988,In_1209);
and U577 (N_577,In_557,In_831);
xor U578 (N_578,In_864,In_1358);
nor U579 (N_579,In_1512,In_1457);
and U580 (N_580,In_732,In_1620);
or U581 (N_581,In_1062,In_1423);
nor U582 (N_582,In_1788,In_1638);
xor U583 (N_583,In_1977,In_1041);
or U584 (N_584,In_1393,In_1858);
xor U585 (N_585,In_700,In_1684);
nand U586 (N_586,In_1250,In_675);
or U587 (N_587,In_1577,In_225);
or U588 (N_588,In_1070,In_1351);
nor U589 (N_589,In_1887,In_1766);
xor U590 (N_590,In_734,In_1032);
or U591 (N_591,In_1549,In_1290);
nor U592 (N_592,In_360,In_1624);
or U593 (N_593,In_1524,In_558);
xor U594 (N_594,In_521,In_455);
or U595 (N_595,In_1700,In_364);
nand U596 (N_596,In_1582,In_1828);
or U597 (N_597,In_290,In_842);
nor U598 (N_598,In_1184,In_678);
nand U599 (N_599,In_1559,In_1228);
nor U600 (N_600,In_1853,In_1974);
nand U601 (N_601,In_288,In_1281);
or U602 (N_602,In_676,In_97);
nor U603 (N_603,In_1539,In_149);
nor U604 (N_604,In_138,In_1005);
or U605 (N_605,In_960,In_206);
and U606 (N_606,In_1254,In_1710);
nand U607 (N_607,In_291,In_311);
xor U608 (N_608,In_532,In_1621);
and U609 (N_609,In_245,In_1563);
and U610 (N_610,In_109,In_1631);
or U611 (N_611,In_835,In_697);
and U612 (N_612,In_779,In_1109);
nor U613 (N_613,In_1800,In_1791);
or U614 (N_614,In_1517,In_1973);
nand U615 (N_615,In_1956,In_1230);
xor U616 (N_616,In_330,In_1415);
xor U617 (N_617,In_28,In_1776);
and U618 (N_618,In_248,In_1860);
xnor U619 (N_619,In_1627,In_1503);
nand U620 (N_620,In_1223,In_716);
nor U621 (N_621,In_690,In_877);
and U622 (N_622,In_1695,In_162);
nor U623 (N_623,In_20,In_899);
or U624 (N_624,In_1255,In_987);
xor U625 (N_625,In_709,In_1535);
nor U626 (N_626,In_96,In_1647);
nand U627 (N_627,In_859,In_1972);
xor U628 (N_628,In_1493,In_478);
and U629 (N_629,In_683,In_742);
xor U630 (N_630,In_539,In_1180);
nand U631 (N_631,In_1115,In_1507);
nor U632 (N_632,In_1825,In_1508);
and U633 (N_633,In_321,In_260);
nor U634 (N_634,In_366,In_1534);
nand U635 (N_635,In_1292,In_1271);
and U636 (N_636,In_496,In_76);
nand U637 (N_637,In_1816,In_1029);
or U638 (N_638,In_1922,In_566);
and U639 (N_639,In_614,In_1368);
and U640 (N_640,In_439,In_63);
nor U641 (N_641,In_1400,In_1752);
xnor U642 (N_642,In_1278,In_1203);
or U643 (N_643,In_1616,In_1918);
or U644 (N_644,In_631,In_1879);
and U645 (N_645,In_1268,In_513);
nand U646 (N_646,In_483,In_196);
xor U647 (N_647,In_729,In_376);
nand U648 (N_648,In_1677,In_1065);
and U649 (N_649,In_1117,In_293);
xor U650 (N_650,In_1068,In_544);
nand U651 (N_651,In_1637,In_136);
or U652 (N_652,In_1623,In_1134);
and U653 (N_653,In_663,In_823);
nor U654 (N_654,In_1195,In_132);
nand U655 (N_655,In_910,In_51);
nor U656 (N_656,In_479,In_258);
and U657 (N_657,In_559,In_582);
nor U658 (N_658,In_542,In_1371);
nor U659 (N_659,In_1489,In_1628);
or U660 (N_660,In_1295,In_1061);
and U661 (N_661,In_1605,In_42);
and U662 (N_662,In_814,In_1548);
and U663 (N_663,In_1898,In_490);
nor U664 (N_664,In_1531,In_644);
or U665 (N_665,In_1558,In_1052);
nor U666 (N_666,In_292,In_1043);
or U667 (N_667,In_1990,In_1516);
xnor U668 (N_668,In_247,In_1432);
or U669 (N_669,In_993,In_1522);
nor U670 (N_670,In_257,In_1685);
xor U671 (N_671,In_403,In_969);
or U672 (N_672,In_817,In_1755);
xnor U673 (N_673,In_983,In_718);
or U674 (N_674,In_282,In_227);
nand U675 (N_675,In_91,In_1253);
xnor U676 (N_676,In_1734,In_1326);
or U677 (N_677,In_587,In_1403);
nand U678 (N_678,In_424,In_1697);
xnor U679 (N_679,In_1418,In_985);
and U680 (N_680,In_1057,In_1950);
nand U681 (N_681,In_858,In_1727);
and U682 (N_682,In_935,In_1179);
xor U683 (N_683,In_55,In_134);
or U684 (N_684,In_1304,In_1015);
nor U685 (N_685,In_998,In_298);
xnor U686 (N_686,In_143,In_161);
and U687 (N_687,In_1819,In_1087);
and U688 (N_688,In_1728,In_711);
nor U689 (N_689,In_1650,In_664);
or U690 (N_690,In_1221,In_868);
nor U691 (N_691,In_41,In_1071);
xnor U692 (N_692,In_1313,In_1243);
and U693 (N_693,In_1107,In_211);
and U694 (N_694,In_748,In_1961);
or U695 (N_695,In_1738,In_501);
and U696 (N_696,In_1740,In_583);
xnor U697 (N_697,In_972,In_5);
nand U698 (N_698,In_1649,In_1690);
nor U699 (N_699,In_319,In_515);
or U700 (N_700,In_199,In_493);
nand U701 (N_701,In_1641,In_194);
and U702 (N_702,In_1565,In_1167);
or U703 (N_703,In_1679,In_393);
and U704 (N_704,In_203,In_83);
nand U705 (N_705,In_1335,In_1046);
or U706 (N_706,In_1422,In_1963);
nor U707 (N_707,In_1169,In_822);
xnor U708 (N_708,In_1055,In_1416);
nor U709 (N_709,In_995,In_1505);
and U710 (N_710,In_1687,In_653);
and U711 (N_711,In_722,In_454);
and U712 (N_712,In_806,In_1206);
nor U713 (N_713,In_668,In_853);
or U714 (N_714,In_32,In_197);
nor U715 (N_715,In_1002,In_1098);
xor U716 (N_716,In_1635,In_1454);
nor U717 (N_717,In_241,In_999);
nand U718 (N_718,In_979,In_414);
xor U719 (N_719,In_1214,In_1475);
and U720 (N_720,In_410,In_1444);
or U721 (N_721,In_409,In_1882);
and U722 (N_722,In_12,In_1981);
xnor U723 (N_723,In_573,In_1366);
nand U724 (N_724,In_1398,In_992);
xor U725 (N_725,In_1289,In_1733);
and U726 (N_726,In_1671,In_1010);
or U727 (N_727,In_276,In_1348);
nor U728 (N_728,In_77,In_852);
or U729 (N_729,In_1293,In_1968);
xnor U730 (N_730,In_1856,In_786);
xnor U731 (N_731,In_1190,In_252);
nor U732 (N_732,In_1305,In_334);
or U733 (N_733,In_201,In_1821);
nand U734 (N_734,In_1866,In_780);
nand U735 (N_735,In_15,In_1201);
or U736 (N_736,In_401,In_704);
nand U737 (N_737,In_849,In_1294);
nand U738 (N_738,In_340,In_1126);
xor U739 (N_739,In_26,In_152);
or U740 (N_740,In_1084,In_253);
xnor U741 (N_741,In_1108,In_1426);
xor U742 (N_742,In_1161,In_1077);
and U743 (N_743,In_1394,In_1327);
nand U744 (N_744,In_1030,In_34);
nor U745 (N_745,In_894,In_1405);
xor U746 (N_746,In_317,In_1601);
nand U747 (N_747,In_1430,In_1135);
nor U748 (N_748,In_740,In_1712);
nand U749 (N_749,In_1429,In_163);
and U750 (N_750,In_963,In_1934);
xnor U751 (N_751,In_745,In_796);
xnor U752 (N_752,In_451,In_70);
nor U753 (N_753,In_1996,In_768);
and U754 (N_754,In_749,In_535);
and U755 (N_755,In_471,In_936);
nor U756 (N_756,In_1659,In_1288);
nor U757 (N_757,In_1663,In_1017);
or U758 (N_758,In_752,In_1749);
and U759 (N_759,In_904,In_448);
nand U760 (N_760,In_250,In_1370);
nand U761 (N_761,In_1485,In_1847);
or U762 (N_762,In_1346,In_466);
or U763 (N_763,In_1551,In_461);
xnor U764 (N_764,In_367,In_1589);
nor U765 (N_765,In_1587,In_810);
xor U766 (N_766,In_75,In_1112);
or U767 (N_767,In_1876,In_1412);
nand U768 (N_768,In_639,In_1552);
and U769 (N_769,In_1725,In_887);
nand U770 (N_770,In_1572,In_349);
nand U771 (N_771,In_1133,In_85);
nand U772 (N_772,In_1388,In_1748);
and U773 (N_773,In_1205,In_115);
xor U774 (N_774,In_553,In_1527);
and U775 (N_775,In_1781,In_202);
or U776 (N_776,In_1911,In_1783);
nand U777 (N_777,In_1026,In_549);
nor U778 (N_778,In_881,In_788);
nor U779 (N_779,In_883,In_114);
and U780 (N_780,In_1543,In_782);
nor U781 (N_781,In_1226,In_346);
xor U782 (N_782,In_811,In_1759);
nand U783 (N_783,In_344,In_540);
nor U784 (N_784,In_1058,In_416);
and U785 (N_785,In_1122,In_1991);
and U786 (N_786,In_350,In_1377);
xor U787 (N_787,In_707,In_415);
xor U788 (N_788,In_1003,In_1235);
xor U789 (N_789,In_1497,In_1120);
or U790 (N_790,In_1706,In_1100);
xnor U791 (N_791,In_428,In_1561);
nor U792 (N_792,In_761,In_89);
nor U793 (N_793,In_365,In_141);
nor U794 (N_794,In_856,In_234);
nor U795 (N_795,In_1308,In_870);
nor U796 (N_796,In_68,In_1384);
nand U797 (N_797,In_1573,In_1983);
xnor U798 (N_798,In_1138,In_1736);
or U799 (N_799,In_1609,In_1938);
nor U800 (N_800,In_574,In_1916);
xor U801 (N_801,In_855,In_146);
and U802 (N_802,In_656,In_502);
nand U803 (N_803,In_1330,In_1869);
nand U804 (N_804,In_1810,In_781);
nor U805 (N_805,In_1822,In_1926);
nor U806 (N_806,In_223,In_692);
and U807 (N_807,In_1965,In_1971);
nand U808 (N_808,In_1851,In_928);
or U809 (N_809,In_137,In_610);
nor U810 (N_810,In_633,In_1603);
and U811 (N_811,In_40,In_608);
or U812 (N_812,In_600,In_179);
or U813 (N_813,In_905,In_838);
nor U814 (N_814,In_797,In_139);
nand U815 (N_815,In_1144,In_686);
xor U816 (N_816,In_1322,In_1256);
and U817 (N_817,In_1473,In_436);
xnor U818 (N_818,In_1737,In_1166);
xor U819 (N_819,In_1342,In_264);
nand U820 (N_820,In_603,In_108);
xor U821 (N_821,In_25,In_442);
nand U822 (N_822,In_431,In_81);
xnor U823 (N_823,In_1751,In_1025);
nor U824 (N_824,In_289,In_848);
or U825 (N_825,In_685,In_94);
nand U826 (N_826,In_1626,In_509);
xor U827 (N_827,In_1283,In_520);
nor U828 (N_828,In_217,In_1156);
nand U829 (N_829,In_397,In_1340);
nor U830 (N_830,In_717,In_1947);
nand U831 (N_831,In_1225,In_503);
xor U832 (N_832,In_342,In_184);
xnor U833 (N_833,In_976,In_100);
or U834 (N_834,In_1066,In_1445);
nand U835 (N_835,In_1282,In_1867);
nor U836 (N_836,In_1546,In_648);
xor U837 (N_837,In_1102,In_649);
nor U838 (N_838,In_1674,In_1806);
and U839 (N_839,In_1088,In_1009);
and U840 (N_840,In_407,In_1318);
xnor U841 (N_841,In_809,In_942);
or U842 (N_842,In_1529,In_1471);
or U843 (N_843,In_1657,In_476);
xor U844 (N_844,In_597,In_1789);
nor U845 (N_845,In_1797,In_1993);
xor U846 (N_846,In_1474,In_488);
or U847 (N_847,In_212,In_1302);
or U848 (N_848,In_1093,In_1111);
or U849 (N_849,In_49,In_180);
nand U850 (N_850,In_665,In_598);
or U851 (N_851,In_1921,In_1175);
nand U852 (N_852,In_795,In_1581);
or U853 (N_853,In_420,In_865);
nor U854 (N_854,In_913,In_516);
nand U855 (N_855,In_1832,In_1964);
nand U856 (N_856,In_636,In_378);
nor U857 (N_857,In_286,In_1249);
or U858 (N_858,In_1610,In_909);
nand U859 (N_859,In_1648,In_1840);
and U860 (N_860,In_200,In_1591);
or U861 (N_861,In_1664,In_757);
xnor U862 (N_862,In_1849,In_1510);
and U863 (N_863,In_1633,In_9);
xor U864 (N_864,In_1823,In_1197);
and U865 (N_865,In_595,In_1483);
xnor U866 (N_866,In_1959,In_736);
or U867 (N_867,In_1655,In_195);
and U868 (N_868,In_1844,In_1790);
nor U869 (N_869,In_694,In_1365);
and U870 (N_870,In_1455,In_989);
nor U871 (N_871,In_1006,In_1187);
nor U872 (N_872,In_1008,In_1151);
or U873 (N_873,In_621,In_1301);
xor U874 (N_874,In_261,In_1857);
nor U875 (N_875,In_1504,In_787);
xnor U876 (N_876,In_931,In_312);
and U877 (N_877,In_1773,In_1141);
and U878 (N_878,In_1329,In_1599);
xnor U879 (N_879,In_541,In_1617);
or U880 (N_880,In_125,In_1438);
and U881 (N_881,In_1270,In_13);
nor U882 (N_882,In_1137,In_815);
nor U883 (N_883,In_1053,In_1360);
nand U884 (N_884,In_492,In_1827);
or U885 (N_885,In_1767,In_1880);
nand U886 (N_886,In_1224,In_1930);
xnor U887 (N_887,In_157,In_1051);
and U888 (N_888,In_926,In_1409);
nor U889 (N_889,In_495,In_375);
and U890 (N_890,In_441,In_1019);
and U891 (N_891,In_19,In_1954);
xnor U892 (N_892,In_1782,In_1196);
nand U893 (N_893,In_1238,In_1027);
nand U894 (N_894,In_61,In_1);
xnor U895 (N_895,In_246,In_1890);
xnor U896 (N_896,In_175,In_445);
nand U897 (N_897,In_1211,In_17);
or U898 (N_898,In_1753,In_947);
and U899 (N_899,In_655,In_1708);
nand U900 (N_900,In_590,In_604);
nor U901 (N_901,In_891,In_494);
and U902 (N_902,In_944,In_1741);
nor U903 (N_903,In_374,In_1127);
nor U904 (N_904,In_1600,In_1402);
nor U905 (N_905,In_444,In_1220);
and U906 (N_906,In_277,In_1897);
xnor U907 (N_907,In_1698,In_588);
xnor U908 (N_908,In_1110,In_458);
xor U909 (N_909,In_957,In_44);
and U910 (N_910,In_1804,In_1047);
xnor U911 (N_911,In_14,In_527);
xor U912 (N_912,In_382,In_737);
and U913 (N_913,In_313,In_850);
nor U914 (N_914,In_1900,In_507);
nor U915 (N_915,In_30,In_1421);
or U916 (N_916,In_624,In_605);
nor U917 (N_917,In_1468,In_563);
xnor U918 (N_918,In_1303,In_510);
nand U919 (N_919,In_46,In_843);
nor U920 (N_920,In_508,In_90);
or U921 (N_921,In_278,In_1132);
nand U922 (N_922,In_962,In_1597);
and U923 (N_923,In_1463,In_1718);
xnor U924 (N_924,In_924,In_164);
xnor U925 (N_925,In_1143,In_952);
xor U926 (N_926,In_1578,In_1408);
xor U927 (N_927,In_945,In_1824);
and U928 (N_928,In_430,In_1920);
and U929 (N_929,In_1446,In_1163);
xor U930 (N_930,In_684,In_1001);
nor U931 (N_931,In_1943,In_1113);
nand U932 (N_932,In_1298,In_1509);
or U933 (N_933,In_460,In_1498);
xor U934 (N_934,In_912,In_1724);
or U935 (N_935,In_1453,In_1390);
xor U936 (N_936,In_543,In_914);
xnor U937 (N_937,In_1219,In_1369);
xor U938 (N_938,In_1854,In_423);
xor U939 (N_939,In_242,In_1396);
nor U940 (N_940,In_1967,In_326);
nor U941 (N_941,In_1976,In_1280);
nor U942 (N_942,In_131,In_1682);
xor U943 (N_943,In_1261,In_872);
and U944 (N_944,In_351,In_1556);
xor U945 (N_945,In_622,In_1467);
xnor U946 (N_946,In_185,In_691);
xor U947 (N_947,In_435,In_1251);
nand U948 (N_948,In_1319,In_1165);
xnor U949 (N_949,In_1488,In_1772);
xor U950 (N_950,In_254,In_682);
or U951 (N_951,In_1701,In_1146);
xor U952 (N_952,In_387,In_1604);
and U953 (N_953,In_537,In_530);
and U954 (N_954,In_1523,In_74);
nor U955 (N_955,In_1124,In_719);
nand U956 (N_956,In_1678,In_1906);
nand U957 (N_957,In_785,In_862);
and U958 (N_958,In_1859,In_1158);
and U959 (N_959,In_1177,In_919);
and U960 (N_960,In_1247,In_1774);
xnor U961 (N_961,In_487,In_1715);
nor U962 (N_962,In_142,In_575);
nor U963 (N_963,In_84,In_1502);
nand U964 (N_964,In_793,In_533);
or U965 (N_965,In_1878,In_1786);
xor U966 (N_966,In_917,In_1692);
and U967 (N_967,In_763,In_1004);
xor U968 (N_968,In_1877,In_1966);
nor U969 (N_969,In_776,In_348);
or U970 (N_970,In_739,In_1929);
xnor U971 (N_971,In_302,In_1613);
or U972 (N_972,In_1830,In_851);
or U973 (N_973,In_1199,In_1596);
or U974 (N_974,In_1925,In_1401);
xnor U975 (N_975,In_177,In_1176);
nor U976 (N_976,In_536,In_160);
xor U977 (N_977,In_475,In_1129);
nor U978 (N_978,In_1932,In_406);
xor U979 (N_979,In_244,In_1831);
xnor U980 (N_980,In_630,In_798);
and U981 (N_981,In_173,In_1873);
and U982 (N_982,In_281,In_1380);
nand U983 (N_983,In_1894,In_1160);
or U984 (N_984,In_825,In_1864);
and U985 (N_985,In_1155,In_11);
nor U986 (N_986,In_943,In_3);
and U987 (N_987,In_356,In_1660);
or U988 (N_988,In_1339,In_1470);
or U989 (N_989,In_1031,In_1232);
nand U990 (N_990,In_578,In_529);
xnor U991 (N_991,In_627,In_1481);
xor U992 (N_992,In_1665,In_1437);
nand U993 (N_993,In_1970,In_1263);
or U994 (N_994,In_915,In_307);
or U995 (N_995,In_1478,In_176);
and U996 (N_996,In_982,In_1035);
and U997 (N_997,In_932,In_1542);
or U998 (N_998,In_1033,In_1928);
nor U999 (N_999,In_612,In_221);
or U1000 (N_1000,In_124,In_358);
and U1001 (N_1001,In_664,In_1109);
xnor U1002 (N_1002,In_1976,In_439);
xnor U1003 (N_1003,In_1789,In_205);
nand U1004 (N_1004,In_1570,In_63);
and U1005 (N_1005,In_1418,In_579);
and U1006 (N_1006,In_1595,In_908);
or U1007 (N_1007,In_1983,In_740);
nand U1008 (N_1008,In_579,In_978);
nand U1009 (N_1009,In_712,In_572);
and U1010 (N_1010,In_1804,In_201);
nand U1011 (N_1011,In_1854,In_1070);
or U1012 (N_1012,In_1750,In_1297);
nand U1013 (N_1013,In_1551,In_146);
and U1014 (N_1014,In_1111,In_1739);
nor U1015 (N_1015,In_1702,In_271);
nand U1016 (N_1016,In_386,In_534);
and U1017 (N_1017,In_695,In_1939);
or U1018 (N_1018,In_1392,In_855);
nor U1019 (N_1019,In_658,In_927);
xor U1020 (N_1020,In_486,In_1877);
nand U1021 (N_1021,In_689,In_109);
nand U1022 (N_1022,In_323,In_766);
or U1023 (N_1023,In_1372,In_1022);
xnor U1024 (N_1024,In_146,In_130);
xnor U1025 (N_1025,In_1825,In_1712);
xnor U1026 (N_1026,In_1721,In_1393);
and U1027 (N_1027,In_82,In_819);
xnor U1028 (N_1028,In_838,In_532);
nand U1029 (N_1029,In_726,In_1605);
and U1030 (N_1030,In_630,In_1324);
and U1031 (N_1031,In_1407,In_1164);
nor U1032 (N_1032,In_30,In_890);
xnor U1033 (N_1033,In_694,In_1739);
or U1034 (N_1034,In_1338,In_1298);
and U1035 (N_1035,In_1977,In_1010);
nand U1036 (N_1036,In_1294,In_1920);
xnor U1037 (N_1037,In_203,In_1034);
nor U1038 (N_1038,In_10,In_930);
nor U1039 (N_1039,In_177,In_367);
nor U1040 (N_1040,In_969,In_472);
nand U1041 (N_1041,In_845,In_1261);
nor U1042 (N_1042,In_1403,In_52);
xnor U1043 (N_1043,In_1485,In_1813);
xnor U1044 (N_1044,In_1772,In_620);
nand U1045 (N_1045,In_327,In_391);
nor U1046 (N_1046,In_1285,In_381);
xor U1047 (N_1047,In_1487,In_754);
and U1048 (N_1048,In_902,In_128);
or U1049 (N_1049,In_1478,In_122);
nand U1050 (N_1050,In_806,In_39);
and U1051 (N_1051,In_366,In_859);
nand U1052 (N_1052,In_1406,In_1748);
and U1053 (N_1053,In_1616,In_481);
nor U1054 (N_1054,In_846,In_343);
and U1055 (N_1055,In_1261,In_1818);
nand U1056 (N_1056,In_1184,In_1992);
xor U1057 (N_1057,In_110,In_1953);
xor U1058 (N_1058,In_320,In_1315);
nor U1059 (N_1059,In_1564,In_434);
xor U1060 (N_1060,In_11,In_1281);
nand U1061 (N_1061,In_1781,In_537);
or U1062 (N_1062,In_1474,In_18);
nor U1063 (N_1063,In_947,In_334);
and U1064 (N_1064,In_1226,In_813);
nand U1065 (N_1065,In_185,In_1936);
or U1066 (N_1066,In_1908,In_1181);
and U1067 (N_1067,In_1344,In_1738);
or U1068 (N_1068,In_1122,In_915);
xor U1069 (N_1069,In_407,In_660);
and U1070 (N_1070,In_703,In_1366);
or U1071 (N_1071,In_857,In_1138);
xor U1072 (N_1072,In_1005,In_1211);
nor U1073 (N_1073,In_486,In_1336);
and U1074 (N_1074,In_1152,In_1042);
xor U1075 (N_1075,In_902,In_143);
nor U1076 (N_1076,In_1934,In_1012);
nor U1077 (N_1077,In_567,In_1826);
xor U1078 (N_1078,In_1712,In_342);
nor U1079 (N_1079,In_460,In_834);
nor U1080 (N_1080,In_723,In_975);
xnor U1081 (N_1081,In_472,In_1881);
nor U1082 (N_1082,In_1127,In_357);
xnor U1083 (N_1083,In_683,In_22);
xnor U1084 (N_1084,In_1013,In_277);
and U1085 (N_1085,In_351,In_1216);
nand U1086 (N_1086,In_214,In_1910);
and U1087 (N_1087,In_1079,In_1225);
nand U1088 (N_1088,In_935,In_351);
nor U1089 (N_1089,In_408,In_1535);
and U1090 (N_1090,In_1712,In_1919);
nand U1091 (N_1091,In_1353,In_709);
or U1092 (N_1092,In_1415,In_1707);
xor U1093 (N_1093,In_1049,In_1355);
and U1094 (N_1094,In_917,In_588);
and U1095 (N_1095,In_53,In_28);
or U1096 (N_1096,In_276,In_1316);
and U1097 (N_1097,In_711,In_507);
and U1098 (N_1098,In_1714,In_1258);
nor U1099 (N_1099,In_144,In_1544);
or U1100 (N_1100,In_1551,In_1626);
nand U1101 (N_1101,In_296,In_1167);
nor U1102 (N_1102,In_1441,In_790);
and U1103 (N_1103,In_1224,In_182);
or U1104 (N_1104,In_212,In_1756);
nor U1105 (N_1105,In_1550,In_768);
and U1106 (N_1106,In_1165,In_1919);
or U1107 (N_1107,In_1430,In_1378);
xnor U1108 (N_1108,In_200,In_433);
and U1109 (N_1109,In_1586,In_956);
nand U1110 (N_1110,In_1167,In_1355);
nand U1111 (N_1111,In_505,In_307);
and U1112 (N_1112,In_1477,In_1923);
or U1113 (N_1113,In_1014,In_1548);
or U1114 (N_1114,In_385,In_828);
nor U1115 (N_1115,In_85,In_1155);
nor U1116 (N_1116,In_351,In_724);
nor U1117 (N_1117,In_606,In_851);
and U1118 (N_1118,In_155,In_1673);
nand U1119 (N_1119,In_134,In_1518);
nand U1120 (N_1120,In_1503,In_1775);
nand U1121 (N_1121,In_743,In_633);
nor U1122 (N_1122,In_1031,In_1948);
and U1123 (N_1123,In_1176,In_414);
nand U1124 (N_1124,In_146,In_1306);
or U1125 (N_1125,In_850,In_604);
xor U1126 (N_1126,In_893,In_927);
or U1127 (N_1127,In_1578,In_1458);
or U1128 (N_1128,In_1825,In_1215);
xnor U1129 (N_1129,In_736,In_412);
nand U1130 (N_1130,In_807,In_1383);
and U1131 (N_1131,In_825,In_712);
nand U1132 (N_1132,In_656,In_332);
nand U1133 (N_1133,In_178,In_816);
xor U1134 (N_1134,In_1677,In_1824);
or U1135 (N_1135,In_1721,In_491);
or U1136 (N_1136,In_1992,In_1226);
nor U1137 (N_1137,In_18,In_493);
nor U1138 (N_1138,In_1669,In_851);
or U1139 (N_1139,In_1124,In_452);
nor U1140 (N_1140,In_1434,In_624);
and U1141 (N_1141,In_318,In_706);
xor U1142 (N_1142,In_244,In_1353);
nor U1143 (N_1143,In_1556,In_463);
and U1144 (N_1144,In_172,In_99);
xor U1145 (N_1145,In_782,In_1098);
nand U1146 (N_1146,In_570,In_863);
xor U1147 (N_1147,In_896,In_996);
nor U1148 (N_1148,In_1753,In_297);
xor U1149 (N_1149,In_856,In_297);
or U1150 (N_1150,In_336,In_21);
nor U1151 (N_1151,In_516,In_1537);
xnor U1152 (N_1152,In_831,In_643);
or U1153 (N_1153,In_1770,In_1200);
or U1154 (N_1154,In_1815,In_852);
or U1155 (N_1155,In_750,In_560);
and U1156 (N_1156,In_1282,In_1209);
or U1157 (N_1157,In_498,In_1032);
and U1158 (N_1158,In_1183,In_1342);
or U1159 (N_1159,In_1279,In_670);
nor U1160 (N_1160,In_760,In_271);
nand U1161 (N_1161,In_1719,In_665);
nand U1162 (N_1162,In_1091,In_167);
nor U1163 (N_1163,In_534,In_1468);
nor U1164 (N_1164,In_1978,In_1162);
nor U1165 (N_1165,In_582,In_1752);
xnor U1166 (N_1166,In_945,In_1505);
nor U1167 (N_1167,In_72,In_935);
or U1168 (N_1168,In_725,In_1967);
nand U1169 (N_1169,In_1133,In_726);
and U1170 (N_1170,In_427,In_1415);
nor U1171 (N_1171,In_1158,In_548);
xor U1172 (N_1172,In_216,In_1930);
xnor U1173 (N_1173,In_738,In_497);
nand U1174 (N_1174,In_1687,In_1229);
nand U1175 (N_1175,In_342,In_1000);
nand U1176 (N_1176,In_1412,In_1712);
nor U1177 (N_1177,In_645,In_1096);
xnor U1178 (N_1178,In_815,In_468);
nand U1179 (N_1179,In_197,In_1637);
nand U1180 (N_1180,In_329,In_1162);
or U1181 (N_1181,In_1675,In_1414);
nor U1182 (N_1182,In_650,In_823);
xor U1183 (N_1183,In_1678,In_399);
nor U1184 (N_1184,In_848,In_1727);
xor U1185 (N_1185,In_1085,In_1641);
nand U1186 (N_1186,In_541,In_1883);
nand U1187 (N_1187,In_388,In_1208);
or U1188 (N_1188,In_159,In_332);
nor U1189 (N_1189,In_1777,In_699);
and U1190 (N_1190,In_725,In_1196);
xnor U1191 (N_1191,In_275,In_1774);
nor U1192 (N_1192,In_1863,In_619);
nor U1193 (N_1193,In_1487,In_59);
and U1194 (N_1194,In_908,In_1781);
xnor U1195 (N_1195,In_260,In_236);
and U1196 (N_1196,In_727,In_618);
xnor U1197 (N_1197,In_1184,In_1030);
xnor U1198 (N_1198,In_1643,In_20);
nor U1199 (N_1199,In_1770,In_1442);
nand U1200 (N_1200,In_1136,In_1890);
xnor U1201 (N_1201,In_886,In_795);
nand U1202 (N_1202,In_842,In_920);
and U1203 (N_1203,In_1690,In_435);
nor U1204 (N_1204,In_1163,In_671);
nor U1205 (N_1205,In_1754,In_1923);
nand U1206 (N_1206,In_528,In_1992);
xnor U1207 (N_1207,In_435,In_1467);
and U1208 (N_1208,In_504,In_257);
and U1209 (N_1209,In_739,In_849);
xor U1210 (N_1210,In_122,In_108);
nand U1211 (N_1211,In_1895,In_846);
or U1212 (N_1212,In_384,In_482);
or U1213 (N_1213,In_939,In_229);
nor U1214 (N_1214,In_1300,In_1034);
nand U1215 (N_1215,In_1843,In_813);
xnor U1216 (N_1216,In_1237,In_1184);
and U1217 (N_1217,In_1394,In_719);
or U1218 (N_1218,In_959,In_236);
and U1219 (N_1219,In_1983,In_200);
and U1220 (N_1220,In_87,In_1742);
and U1221 (N_1221,In_1186,In_278);
xnor U1222 (N_1222,In_1157,In_1309);
xor U1223 (N_1223,In_1471,In_852);
and U1224 (N_1224,In_243,In_1541);
xnor U1225 (N_1225,In_1750,In_233);
and U1226 (N_1226,In_982,In_471);
nor U1227 (N_1227,In_1386,In_527);
or U1228 (N_1228,In_367,In_1705);
nand U1229 (N_1229,In_105,In_1185);
or U1230 (N_1230,In_1307,In_312);
xnor U1231 (N_1231,In_1751,In_360);
nand U1232 (N_1232,In_103,In_647);
xnor U1233 (N_1233,In_193,In_558);
xnor U1234 (N_1234,In_390,In_1245);
or U1235 (N_1235,In_1450,In_1652);
nand U1236 (N_1236,In_739,In_787);
or U1237 (N_1237,In_931,In_9);
or U1238 (N_1238,In_708,In_296);
nand U1239 (N_1239,In_488,In_1850);
and U1240 (N_1240,In_1911,In_937);
or U1241 (N_1241,In_743,In_1593);
or U1242 (N_1242,In_663,In_1032);
and U1243 (N_1243,In_1402,In_1472);
nor U1244 (N_1244,In_1385,In_1554);
and U1245 (N_1245,In_1581,In_1742);
xnor U1246 (N_1246,In_1140,In_1949);
or U1247 (N_1247,In_382,In_1474);
or U1248 (N_1248,In_1529,In_822);
nor U1249 (N_1249,In_466,In_1641);
and U1250 (N_1250,In_1803,In_1586);
and U1251 (N_1251,In_1045,In_1373);
and U1252 (N_1252,In_1004,In_1552);
xor U1253 (N_1253,In_1462,In_834);
or U1254 (N_1254,In_1524,In_1015);
xnor U1255 (N_1255,In_865,In_764);
nor U1256 (N_1256,In_54,In_916);
nand U1257 (N_1257,In_1955,In_1545);
nor U1258 (N_1258,In_1709,In_219);
and U1259 (N_1259,In_1607,In_355);
and U1260 (N_1260,In_290,In_1550);
and U1261 (N_1261,In_1637,In_1322);
or U1262 (N_1262,In_1828,In_118);
and U1263 (N_1263,In_183,In_1587);
nor U1264 (N_1264,In_155,In_1640);
xnor U1265 (N_1265,In_1540,In_634);
or U1266 (N_1266,In_1269,In_1193);
or U1267 (N_1267,In_510,In_230);
and U1268 (N_1268,In_309,In_836);
and U1269 (N_1269,In_1750,In_1171);
nand U1270 (N_1270,In_1606,In_1633);
and U1271 (N_1271,In_302,In_93);
or U1272 (N_1272,In_388,In_1559);
and U1273 (N_1273,In_1385,In_1722);
nand U1274 (N_1274,In_1363,In_1169);
nor U1275 (N_1275,In_1963,In_1900);
or U1276 (N_1276,In_1436,In_198);
or U1277 (N_1277,In_1836,In_1824);
and U1278 (N_1278,In_941,In_609);
xor U1279 (N_1279,In_341,In_1097);
and U1280 (N_1280,In_681,In_159);
xnor U1281 (N_1281,In_181,In_1436);
or U1282 (N_1282,In_1247,In_733);
or U1283 (N_1283,In_551,In_613);
xor U1284 (N_1284,In_634,In_214);
or U1285 (N_1285,In_1655,In_681);
nand U1286 (N_1286,In_193,In_883);
or U1287 (N_1287,In_735,In_110);
or U1288 (N_1288,In_1140,In_1674);
xnor U1289 (N_1289,In_1585,In_1527);
xnor U1290 (N_1290,In_1739,In_1090);
and U1291 (N_1291,In_1048,In_540);
nand U1292 (N_1292,In_380,In_1889);
nand U1293 (N_1293,In_894,In_1742);
xnor U1294 (N_1294,In_1793,In_1638);
and U1295 (N_1295,In_525,In_827);
and U1296 (N_1296,In_808,In_1555);
nor U1297 (N_1297,In_1514,In_1005);
nor U1298 (N_1298,In_56,In_1838);
or U1299 (N_1299,In_1388,In_1281);
and U1300 (N_1300,In_731,In_1981);
xnor U1301 (N_1301,In_1979,In_640);
and U1302 (N_1302,In_1611,In_1003);
or U1303 (N_1303,In_1485,In_1734);
and U1304 (N_1304,In_1847,In_359);
xor U1305 (N_1305,In_1751,In_238);
xor U1306 (N_1306,In_1211,In_1586);
xor U1307 (N_1307,In_225,In_1915);
xnor U1308 (N_1308,In_1816,In_794);
and U1309 (N_1309,In_1134,In_1052);
xor U1310 (N_1310,In_1205,In_1474);
or U1311 (N_1311,In_1711,In_721);
xor U1312 (N_1312,In_1113,In_1737);
and U1313 (N_1313,In_25,In_1427);
xnor U1314 (N_1314,In_1253,In_1969);
nor U1315 (N_1315,In_54,In_1185);
xor U1316 (N_1316,In_689,In_981);
xnor U1317 (N_1317,In_1953,In_727);
or U1318 (N_1318,In_1315,In_490);
or U1319 (N_1319,In_856,In_1242);
and U1320 (N_1320,In_755,In_1111);
nor U1321 (N_1321,In_726,In_659);
nand U1322 (N_1322,In_1009,In_1833);
or U1323 (N_1323,In_537,In_23);
xor U1324 (N_1324,In_684,In_505);
nand U1325 (N_1325,In_1025,In_1052);
and U1326 (N_1326,In_52,In_11);
nor U1327 (N_1327,In_1560,In_1562);
nand U1328 (N_1328,In_1890,In_1285);
nor U1329 (N_1329,In_1036,In_1363);
and U1330 (N_1330,In_1407,In_344);
xnor U1331 (N_1331,In_490,In_1003);
and U1332 (N_1332,In_761,In_622);
or U1333 (N_1333,In_1238,In_298);
and U1334 (N_1334,In_1388,In_1994);
nor U1335 (N_1335,In_1170,In_294);
and U1336 (N_1336,In_1741,In_1286);
or U1337 (N_1337,In_628,In_1977);
nand U1338 (N_1338,In_104,In_243);
xor U1339 (N_1339,In_1185,In_1288);
and U1340 (N_1340,In_1348,In_1653);
nand U1341 (N_1341,In_1296,In_864);
nand U1342 (N_1342,In_691,In_1027);
nor U1343 (N_1343,In_234,In_1265);
and U1344 (N_1344,In_1607,In_1891);
or U1345 (N_1345,In_1805,In_1934);
or U1346 (N_1346,In_1797,In_1508);
xnor U1347 (N_1347,In_1890,In_1785);
nand U1348 (N_1348,In_1852,In_146);
xnor U1349 (N_1349,In_1096,In_1565);
nand U1350 (N_1350,In_401,In_1025);
nand U1351 (N_1351,In_349,In_1339);
or U1352 (N_1352,In_535,In_1089);
nor U1353 (N_1353,In_362,In_1734);
and U1354 (N_1354,In_541,In_581);
and U1355 (N_1355,In_1136,In_314);
nor U1356 (N_1356,In_1246,In_1436);
and U1357 (N_1357,In_749,In_424);
or U1358 (N_1358,In_1862,In_208);
and U1359 (N_1359,In_541,In_1238);
xor U1360 (N_1360,In_264,In_1261);
nor U1361 (N_1361,In_470,In_449);
nand U1362 (N_1362,In_1682,In_741);
or U1363 (N_1363,In_1270,In_1364);
nor U1364 (N_1364,In_187,In_106);
or U1365 (N_1365,In_1834,In_1102);
nand U1366 (N_1366,In_493,In_651);
or U1367 (N_1367,In_1860,In_865);
nand U1368 (N_1368,In_591,In_263);
and U1369 (N_1369,In_1590,In_307);
xor U1370 (N_1370,In_267,In_68);
and U1371 (N_1371,In_957,In_1957);
and U1372 (N_1372,In_1153,In_189);
and U1373 (N_1373,In_1436,In_1179);
nand U1374 (N_1374,In_179,In_1323);
and U1375 (N_1375,In_1421,In_206);
or U1376 (N_1376,In_1372,In_620);
nand U1377 (N_1377,In_1670,In_1200);
nor U1378 (N_1378,In_590,In_1168);
or U1379 (N_1379,In_1126,In_1922);
xor U1380 (N_1380,In_490,In_1525);
or U1381 (N_1381,In_1198,In_1942);
nand U1382 (N_1382,In_1697,In_1217);
nor U1383 (N_1383,In_612,In_554);
nand U1384 (N_1384,In_1024,In_190);
and U1385 (N_1385,In_1357,In_180);
nor U1386 (N_1386,In_941,In_1453);
xnor U1387 (N_1387,In_307,In_954);
nor U1388 (N_1388,In_1869,In_1049);
or U1389 (N_1389,In_302,In_1482);
or U1390 (N_1390,In_702,In_1670);
xnor U1391 (N_1391,In_511,In_462);
nor U1392 (N_1392,In_604,In_989);
and U1393 (N_1393,In_625,In_1671);
or U1394 (N_1394,In_686,In_1542);
nand U1395 (N_1395,In_1157,In_966);
nor U1396 (N_1396,In_499,In_809);
xor U1397 (N_1397,In_824,In_1740);
or U1398 (N_1398,In_529,In_2);
nand U1399 (N_1399,In_1186,In_1825);
or U1400 (N_1400,In_888,In_781);
nand U1401 (N_1401,In_1527,In_1257);
or U1402 (N_1402,In_384,In_959);
nor U1403 (N_1403,In_1082,In_334);
nor U1404 (N_1404,In_281,In_1322);
xnor U1405 (N_1405,In_1650,In_1715);
nand U1406 (N_1406,In_361,In_230);
xor U1407 (N_1407,In_1154,In_1541);
and U1408 (N_1408,In_964,In_1604);
nor U1409 (N_1409,In_442,In_902);
or U1410 (N_1410,In_443,In_171);
nor U1411 (N_1411,In_740,In_1563);
or U1412 (N_1412,In_1271,In_566);
and U1413 (N_1413,In_1918,In_210);
and U1414 (N_1414,In_1515,In_1523);
nor U1415 (N_1415,In_1160,In_1986);
nor U1416 (N_1416,In_72,In_451);
or U1417 (N_1417,In_1434,In_1810);
and U1418 (N_1418,In_1597,In_1474);
nand U1419 (N_1419,In_514,In_455);
xnor U1420 (N_1420,In_458,In_806);
nor U1421 (N_1421,In_884,In_1720);
nand U1422 (N_1422,In_978,In_85);
or U1423 (N_1423,In_1680,In_1613);
xor U1424 (N_1424,In_99,In_1234);
xnor U1425 (N_1425,In_1473,In_1557);
xor U1426 (N_1426,In_343,In_1968);
nor U1427 (N_1427,In_747,In_1801);
nand U1428 (N_1428,In_981,In_615);
nor U1429 (N_1429,In_1301,In_927);
or U1430 (N_1430,In_713,In_1662);
or U1431 (N_1431,In_309,In_965);
or U1432 (N_1432,In_1078,In_192);
or U1433 (N_1433,In_945,In_380);
nand U1434 (N_1434,In_637,In_1723);
nand U1435 (N_1435,In_1943,In_1909);
xnor U1436 (N_1436,In_1027,In_1779);
or U1437 (N_1437,In_1789,In_1297);
and U1438 (N_1438,In_792,In_439);
nor U1439 (N_1439,In_910,In_474);
and U1440 (N_1440,In_904,In_169);
nor U1441 (N_1441,In_955,In_852);
and U1442 (N_1442,In_1172,In_1903);
nor U1443 (N_1443,In_598,In_1342);
nand U1444 (N_1444,In_81,In_1084);
xor U1445 (N_1445,In_1871,In_507);
xor U1446 (N_1446,In_1933,In_1680);
and U1447 (N_1447,In_619,In_1030);
and U1448 (N_1448,In_312,In_350);
nand U1449 (N_1449,In_1551,In_1758);
and U1450 (N_1450,In_770,In_1214);
xnor U1451 (N_1451,In_260,In_332);
nor U1452 (N_1452,In_529,In_1255);
and U1453 (N_1453,In_1571,In_1367);
or U1454 (N_1454,In_199,In_605);
and U1455 (N_1455,In_445,In_1967);
or U1456 (N_1456,In_625,In_342);
nor U1457 (N_1457,In_1296,In_794);
nor U1458 (N_1458,In_973,In_1868);
and U1459 (N_1459,In_794,In_1799);
nor U1460 (N_1460,In_1477,In_922);
or U1461 (N_1461,In_1285,In_765);
or U1462 (N_1462,In_179,In_1981);
xor U1463 (N_1463,In_1257,In_1224);
nor U1464 (N_1464,In_1043,In_1907);
nand U1465 (N_1465,In_1523,In_1019);
xor U1466 (N_1466,In_1520,In_1692);
nand U1467 (N_1467,In_422,In_1458);
xor U1468 (N_1468,In_1533,In_160);
nand U1469 (N_1469,In_52,In_788);
nand U1470 (N_1470,In_562,In_649);
nand U1471 (N_1471,In_1661,In_761);
xor U1472 (N_1472,In_1622,In_338);
or U1473 (N_1473,In_1606,In_778);
nor U1474 (N_1474,In_1416,In_950);
nand U1475 (N_1475,In_1625,In_1606);
and U1476 (N_1476,In_1890,In_1278);
nor U1477 (N_1477,In_946,In_1421);
and U1478 (N_1478,In_174,In_1280);
and U1479 (N_1479,In_542,In_893);
and U1480 (N_1480,In_560,In_1841);
xnor U1481 (N_1481,In_1574,In_744);
xor U1482 (N_1482,In_1223,In_1336);
nand U1483 (N_1483,In_670,In_282);
xnor U1484 (N_1484,In_728,In_571);
xor U1485 (N_1485,In_1598,In_1975);
or U1486 (N_1486,In_1656,In_248);
nor U1487 (N_1487,In_818,In_1506);
nand U1488 (N_1488,In_809,In_1126);
nor U1489 (N_1489,In_241,In_671);
or U1490 (N_1490,In_713,In_1608);
or U1491 (N_1491,In_182,In_1358);
and U1492 (N_1492,In_1559,In_799);
nor U1493 (N_1493,In_1664,In_1569);
and U1494 (N_1494,In_850,In_955);
and U1495 (N_1495,In_1810,In_905);
xnor U1496 (N_1496,In_1440,In_670);
and U1497 (N_1497,In_150,In_5);
nand U1498 (N_1498,In_146,In_1053);
and U1499 (N_1499,In_1030,In_280);
nand U1500 (N_1500,In_799,In_38);
nor U1501 (N_1501,In_222,In_1597);
nand U1502 (N_1502,In_1545,In_1063);
and U1503 (N_1503,In_327,In_192);
or U1504 (N_1504,In_1606,In_1929);
or U1505 (N_1505,In_1585,In_765);
or U1506 (N_1506,In_1691,In_48);
nor U1507 (N_1507,In_1156,In_1670);
or U1508 (N_1508,In_1510,In_184);
and U1509 (N_1509,In_831,In_1300);
and U1510 (N_1510,In_396,In_1570);
and U1511 (N_1511,In_1946,In_1791);
or U1512 (N_1512,In_1799,In_43);
or U1513 (N_1513,In_1418,In_1400);
or U1514 (N_1514,In_816,In_1385);
and U1515 (N_1515,In_892,In_125);
or U1516 (N_1516,In_1629,In_683);
xnor U1517 (N_1517,In_1314,In_598);
xnor U1518 (N_1518,In_352,In_1440);
nor U1519 (N_1519,In_1250,In_1811);
xnor U1520 (N_1520,In_910,In_403);
and U1521 (N_1521,In_1313,In_439);
xnor U1522 (N_1522,In_54,In_1576);
xnor U1523 (N_1523,In_118,In_1045);
xnor U1524 (N_1524,In_371,In_141);
or U1525 (N_1525,In_1653,In_1174);
and U1526 (N_1526,In_491,In_1960);
xnor U1527 (N_1527,In_1599,In_1390);
xnor U1528 (N_1528,In_795,In_1267);
xor U1529 (N_1529,In_792,In_421);
xor U1530 (N_1530,In_1688,In_62);
nor U1531 (N_1531,In_438,In_1280);
xnor U1532 (N_1532,In_1708,In_1185);
nand U1533 (N_1533,In_51,In_1288);
or U1534 (N_1534,In_526,In_811);
nor U1535 (N_1535,In_757,In_1081);
nand U1536 (N_1536,In_1159,In_497);
and U1537 (N_1537,In_1650,In_1952);
or U1538 (N_1538,In_483,In_708);
and U1539 (N_1539,In_1267,In_624);
xnor U1540 (N_1540,In_617,In_71);
nand U1541 (N_1541,In_691,In_1609);
nor U1542 (N_1542,In_1365,In_914);
xor U1543 (N_1543,In_1386,In_822);
and U1544 (N_1544,In_592,In_963);
nand U1545 (N_1545,In_933,In_1825);
and U1546 (N_1546,In_732,In_449);
or U1547 (N_1547,In_1727,In_504);
xnor U1548 (N_1548,In_1094,In_649);
xor U1549 (N_1549,In_1951,In_1348);
xor U1550 (N_1550,In_255,In_917);
or U1551 (N_1551,In_1245,In_741);
nand U1552 (N_1552,In_1821,In_601);
xnor U1553 (N_1553,In_422,In_1848);
xnor U1554 (N_1554,In_989,In_912);
xor U1555 (N_1555,In_46,In_966);
xor U1556 (N_1556,In_658,In_1717);
or U1557 (N_1557,In_1230,In_639);
or U1558 (N_1558,In_1364,In_1242);
nand U1559 (N_1559,In_1046,In_1760);
or U1560 (N_1560,In_668,In_1448);
nand U1561 (N_1561,In_1602,In_1623);
and U1562 (N_1562,In_1325,In_22);
nand U1563 (N_1563,In_1772,In_1903);
nand U1564 (N_1564,In_1942,In_1422);
and U1565 (N_1565,In_475,In_1098);
and U1566 (N_1566,In_1664,In_1050);
xnor U1567 (N_1567,In_1412,In_601);
and U1568 (N_1568,In_1426,In_1026);
or U1569 (N_1569,In_1631,In_624);
and U1570 (N_1570,In_1600,In_831);
nand U1571 (N_1571,In_1650,In_1176);
or U1572 (N_1572,In_39,In_1019);
xnor U1573 (N_1573,In_638,In_527);
nand U1574 (N_1574,In_655,In_1229);
or U1575 (N_1575,In_830,In_222);
nand U1576 (N_1576,In_642,In_1821);
nand U1577 (N_1577,In_1221,In_581);
xor U1578 (N_1578,In_911,In_727);
nor U1579 (N_1579,In_1851,In_1133);
nand U1580 (N_1580,In_1360,In_872);
nand U1581 (N_1581,In_523,In_1869);
nor U1582 (N_1582,In_208,In_757);
xor U1583 (N_1583,In_771,In_664);
nand U1584 (N_1584,In_158,In_1175);
xor U1585 (N_1585,In_1255,In_275);
nor U1586 (N_1586,In_312,In_1180);
and U1587 (N_1587,In_672,In_338);
nor U1588 (N_1588,In_1888,In_1626);
nor U1589 (N_1589,In_1701,In_342);
nand U1590 (N_1590,In_1369,In_1133);
nor U1591 (N_1591,In_457,In_198);
and U1592 (N_1592,In_315,In_782);
nand U1593 (N_1593,In_467,In_923);
or U1594 (N_1594,In_942,In_517);
and U1595 (N_1595,In_1557,In_1573);
and U1596 (N_1596,In_257,In_298);
or U1597 (N_1597,In_1491,In_1100);
xor U1598 (N_1598,In_695,In_1391);
and U1599 (N_1599,In_1747,In_268);
and U1600 (N_1600,In_850,In_470);
nor U1601 (N_1601,In_947,In_613);
xnor U1602 (N_1602,In_1104,In_760);
nand U1603 (N_1603,In_1190,In_782);
or U1604 (N_1604,In_939,In_1911);
nand U1605 (N_1605,In_1574,In_1162);
xor U1606 (N_1606,In_32,In_1104);
nand U1607 (N_1607,In_884,In_317);
xnor U1608 (N_1608,In_834,In_823);
xnor U1609 (N_1609,In_311,In_702);
or U1610 (N_1610,In_542,In_656);
or U1611 (N_1611,In_1235,In_996);
xnor U1612 (N_1612,In_1948,In_1107);
xor U1613 (N_1613,In_1703,In_991);
or U1614 (N_1614,In_428,In_1817);
or U1615 (N_1615,In_468,In_1347);
nand U1616 (N_1616,In_975,In_865);
or U1617 (N_1617,In_801,In_394);
or U1618 (N_1618,In_928,In_1529);
nand U1619 (N_1619,In_714,In_379);
and U1620 (N_1620,In_1991,In_386);
nand U1621 (N_1621,In_1181,In_1193);
nor U1622 (N_1622,In_1384,In_256);
nand U1623 (N_1623,In_196,In_395);
xor U1624 (N_1624,In_1539,In_846);
and U1625 (N_1625,In_1184,In_42);
nand U1626 (N_1626,In_648,In_161);
or U1627 (N_1627,In_1587,In_11);
or U1628 (N_1628,In_1499,In_1838);
nand U1629 (N_1629,In_4,In_1008);
and U1630 (N_1630,In_106,In_1123);
xor U1631 (N_1631,In_269,In_176);
nand U1632 (N_1632,In_471,In_1109);
or U1633 (N_1633,In_1785,In_844);
xnor U1634 (N_1634,In_1706,In_1927);
xor U1635 (N_1635,In_955,In_1952);
nand U1636 (N_1636,In_937,In_1835);
and U1637 (N_1637,In_1649,In_392);
nor U1638 (N_1638,In_373,In_867);
nor U1639 (N_1639,In_692,In_1209);
nor U1640 (N_1640,In_1920,In_1622);
nor U1641 (N_1641,In_1212,In_1226);
and U1642 (N_1642,In_635,In_1676);
nand U1643 (N_1643,In_601,In_1983);
nand U1644 (N_1644,In_106,In_1293);
and U1645 (N_1645,In_216,In_362);
or U1646 (N_1646,In_116,In_416);
or U1647 (N_1647,In_777,In_772);
or U1648 (N_1648,In_373,In_1057);
nand U1649 (N_1649,In_1229,In_495);
nor U1650 (N_1650,In_722,In_1380);
nand U1651 (N_1651,In_1194,In_768);
nor U1652 (N_1652,In_1169,In_1655);
nand U1653 (N_1653,In_942,In_687);
xnor U1654 (N_1654,In_1287,In_117);
and U1655 (N_1655,In_713,In_1487);
xor U1656 (N_1656,In_1903,In_1217);
and U1657 (N_1657,In_1943,In_298);
and U1658 (N_1658,In_302,In_468);
nor U1659 (N_1659,In_238,In_1530);
nand U1660 (N_1660,In_1880,In_551);
and U1661 (N_1661,In_1943,In_446);
nor U1662 (N_1662,In_1841,In_1919);
or U1663 (N_1663,In_1136,In_1258);
xor U1664 (N_1664,In_1182,In_1077);
nand U1665 (N_1665,In_837,In_185);
nor U1666 (N_1666,In_448,In_1052);
xor U1667 (N_1667,In_731,In_1490);
or U1668 (N_1668,In_1432,In_772);
xor U1669 (N_1669,In_1389,In_195);
xor U1670 (N_1670,In_1760,In_4);
xor U1671 (N_1671,In_1728,In_779);
nand U1672 (N_1672,In_1537,In_1512);
xor U1673 (N_1673,In_1622,In_1839);
or U1674 (N_1674,In_132,In_1183);
xor U1675 (N_1675,In_1098,In_871);
or U1676 (N_1676,In_1051,In_945);
xor U1677 (N_1677,In_625,In_1169);
nand U1678 (N_1678,In_1261,In_979);
xor U1679 (N_1679,In_768,In_913);
or U1680 (N_1680,In_768,In_1355);
nor U1681 (N_1681,In_952,In_1222);
xor U1682 (N_1682,In_105,In_423);
xnor U1683 (N_1683,In_844,In_1400);
xnor U1684 (N_1684,In_135,In_4);
and U1685 (N_1685,In_1454,In_1936);
or U1686 (N_1686,In_855,In_12);
or U1687 (N_1687,In_143,In_170);
nor U1688 (N_1688,In_787,In_1389);
xnor U1689 (N_1689,In_590,In_14);
and U1690 (N_1690,In_1419,In_378);
nor U1691 (N_1691,In_158,In_1885);
and U1692 (N_1692,In_1620,In_1067);
nor U1693 (N_1693,In_1168,In_54);
and U1694 (N_1694,In_458,In_147);
or U1695 (N_1695,In_132,In_1839);
nand U1696 (N_1696,In_1357,In_1530);
or U1697 (N_1697,In_1000,In_946);
nor U1698 (N_1698,In_623,In_1916);
xnor U1699 (N_1699,In_982,In_871);
nand U1700 (N_1700,In_844,In_531);
and U1701 (N_1701,In_873,In_1700);
nor U1702 (N_1702,In_1692,In_944);
xor U1703 (N_1703,In_179,In_276);
nor U1704 (N_1704,In_1873,In_1321);
nand U1705 (N_1705,In_1407,In_1162);
nand U1706 (N_1706,In_1908,In_465);
nor U1707 (N_1707,In_1706,In_884);
and U1708 (N_1708,In_567,In_729);
nor U1709 (N_1709,In_1500,In_1950);
nand U1710 (N_1710,In_1453,In_1510);
xor U1711 (N_1711,In_1918,In_1750);
xor U1712 (N_1712,In_110,In_1045);
or U1713 (N_1713,In_332,In_1410);
nand U1714 (N_1714,In_1455,In_307);
nor U1715 (N_1715,In_971,In_1844);
nand U1716 (N_1716,In_1113,In_484);
and U1717 (N_1717,In_1473,In_1361);
nand U1718 (N_1718,In_477,In_688);
xnor U1719 (N_1719,In_1331,In_1339);
or U1720 (N_1720,In_1955,In_896);
and U1721 (N_1721,In_1900,In_1015);
or U1722 (N_1722,In_1302,In_1162);
or U1723 (N_1723,In_1184,In_481);
or U1724 (N_1724,In_1691,In_188);
nor U1725 (N_1725,In_1317,In_1633);
or U1726 (N_1726,In_920,In_1201);
nand U1727 (N_1727,In_926,In_1983);
and U1728 (N_1728,In_1493,In_1408);
xor U1729 (N_1729,In_309,In_544);
nor U1730 (N_1730,In_1407,In_293);
or U1731 (N_1731,In_1054,In_671);
or U1732 (N_1732,In_1913,In_1336);
or U1733 (N_1733,In_1266,In_76);
xor U1734 (N_1734,In_1643,In_1639);
and U1735 (N_1735,In_681,In_400);
or U1736 (N_1736,In_1567,In_258);
or U1737 (N_1737,In_677,In_846);
and U1738 (N_1738,In_485,In_1231);
and U1739 (N_1739,In_706,In_112);
nor U1740 (N_1740,In_304,In_856);
nor U1741 (N_1741,In_605,In_461);
or U1742 (N_1742,In_1579,In_572);
or U1743 (N_1743,In_1122,In_1329);
or U1744 (N_1744,In_552,In_1273);
xor U1745 (N_1745,In_1105,In_1979);
xor U1746 (N_1746,In_1317,In_245);
nand U1747 (N_1747,In_1352,In_1126);
xnor U1748 (N_1748,In_1230,In_280);
nor U1749 (N_1749,In_701,In_1871);
and U1750 (N_1750,In_482,In_1361);
or U1751 (N_1751,In_326,In_1485);
xor U1752 (N_1752,In_932,In_1019);
nand U1753 (N_1753,In_1449,In_1793);
nor U1754 (N_1754,In_1005,In_1314);
and U1755 (N_1755,In_1671,In_1230);
nand U1756 (N_1756,In_1072,In_322);
or U1757 (N_1757,In_1833,In_1685);
or U1758 (N_1758,In_1983,In_1802);
nor U1759 (N_1759,In_1767,In_633);
nand U1760 (N_1760,In_772,In_359);
and U1761 (N_1761,In_210,In_1251);
or U1762 (N_1762,In_302,In_1229);
xnor U1763 (N_1763,In_477,In_1918);
nor U1764 (N_1764,In_1182,In_924);
nand U1765 (N_1765,In_1829,In_601);
and U1766 (N_1766,In_1968,In_143);
or U1767 (N_1767,In_1784,In_1775);
nor U1768 (N_1768,In_1897,In_1505);
xor U1769 (N_1769,In_1807,In_1112);
xnor U1770 (N_1770,In_823,In_1654);
nor U1771 (N_1771,In_369,In_126);
and U1772 (N_1772,In_1762,In_1186);
xnor U1773 (N_1773,In_345,In_1460);
xnor U1774 (N_1774,In_1741,In_128);
nand U1775 (N_1775,In_456,In_1383);
nor U1776 (N_1776,In_1944,In_637);
or U1777 (N_1777,In_782,In_1827);
nand U1778 (N_1778,In_1954,In_1111);
and U1779 (N_1779,In_716,In_776);
xor U1780 (N_1780,In_874,In_866);
xnor U1781 (N_1781,In_416,In_1932);
and U1782 (N_1782,In_330,In_278);
or U1783 (N_1783,In_1884,In_1789);
and U1784 (N_1784,In_81,In_1515);
nor U1785 (N_1785,In_904,In_1873);
nand U1786 (N_1786,In_301,In_374);
or U1787 (N_1787,In_869,In_1917);
xor U1788 (N_1788,In_1938,In_1936);
nand U1789 (N_1789,In_1540,In_61);
or U1790 (N_1790,In_1026,In_287);
nand U1791 (N_1791,In_221,In_500);
or U1792 (N_1792,In_1200,In_580);
xor U1793 (N_1793,In_1638,In_867);
nor U1794 (N_1794,In_541,In_1987);
and U1795 (N_1795,In_113,In_250);
nor U1796 (N_1796,In_670,In_1171);
xor U1797 (N_1797,In_471,In_1382);
or U1798 (N_1798,In_684,In_44);
or U1799 (N_1799,In_1863,In_682);
or U1800 (N_1800,In_1267,In_687);
or U1801 (N_1801,In_1897,In_226);
nor U1802 (N_1802,In_984,In_1930);
or U1803 (N_1803,In_691,In_534);
and U1804 (N_1804,In_1286,In_1547);
xor U1805 (N_1805,In_1724,In_510);
xor U1806 (N_1806,In_523,In_183);
nand U1807 (N_1807,In_388,In_1511);
and U1808 (N_1808,In_963,In_1589);
and U1809 (N_1809,In_755,In_1118);
nand U1810 (N_1810,In_970,In_1975);
or U1811 (N_1811,In_308,In_1314);
and U1812 (N_1812,In_218,In_925);
or U1813 (N_1813,In_1164,In_1562);
nor U1814 (N_1814,In_1608,In_1129);
or U1815 (N_1815,In_1867,In_100);
nor U1816 (N_1816,In_1132,In_1767);
xor U1817 (N_1817,In_1573,In_1244);
nand U1818 (N_1818,In_370,In_336);
nor U1819 (N_1819,In_1782,In_964);
nand U1820 (N_1820,In_334,In_805);
and U1821 (N_1821,In_617,In_892);
nor U1822 (N_1822,In_1478,In_1173);
nor U1823 (N_1823,In_713,In_581);
nand U1824 (N_1824,In_464,In_617);
and U1825 (N_1825,In_1019,In_319);
xor U1826 (N_1826,In_1786,In_1962);
nand U1827 (N_1827,In_1640,In_1514);
nand U1828 (N_1828,In_1965,In_214);
and U1829 (N_1829,In_1245,In_1740);
and U1830 (N_1830,In_555,In_1503);
nand U1831 (N_1831,In_1687,In_507);
nor U1832 (N_1832,In_1776,In_1934);
and U1833 (N_1833,In_1949,In_1449);
nand U1834 (N_1834,In_1990,In_1218);
nand U1835 (N_1835,In_1556,In_443);
nor U1836 (N_1836,In_422,In_391);
or U1837 (N_1837,In_1182,In_372);
and U1838 (N_1838,In_312,In_213);
or U1839 (N_1839,In_1465,In_42);
nand U1840 (N_1840,In_646,In_274);
or U1841 (N_1841,In_1410,In_563);
or U1842 (N_1842,In_1594,In_622);
and U1843 (N_1843,In_1281,In_633);
or U1844 (N_1844,In_643,In_1546);
or U1845 (N_1845,In_1921,In_1267);
nand U1846 (N_1846,In_768,In_58);
nand U1847 (N_1847,In_1993,In_670);
xor U1848 (N_1848,In_138,In_1611);
and U1849 (N_1849,In_242,In_1183);
nand U1850 (N_1850,In_453,In_1031);
nor U1851 (N_1851,In_1316,In_650);
nor U1852 (N_1852,In_1825,In_406);
nand U1853 (N_1853,In_179,In_671);
or U1854 (N_1854,In_1701,In_1655);
xor U1855 (N_1855,In_261,In_1112);
or U1856 (N_1856,In_1030,In_1731);
or U1857 (N_1857,In_980,In_495);
xor U1858 (N_1858,In_1309,In_1529);
xor U1859 (N_1859,In_749,In_30);
xor U1860 (N_1860,In_1897,In_139);
or U1861 (N_1861,In_1671,In_1533);
and U1862 (N_1862,In_929,In_1636);
nor U1863 (N_1863,In_783,In_121);
nor U1864 (N_1864,In_991,In_1297);
nor U1865 (N_1865,In_6,In_751);
xnor U1866 (N_1866,In_153,In_583);
nand U1867 (N_1867,In_1238,In_339);
xnor U1868 (N_1868,In_547,In_842);
xor U1869 (N_1869,In_646,In_1017);
xor U1870 (N_1870,In_443,In_61);
or U1871 (N_1871,In_989,In_1535);
and U1872 (N_1872,In_754,In_409);
and U1873 (N_1873,In_1722,In_1223);
nor U1874 (N_1874,In_1107,In_371);
or U1875 (N_1875,In_1851,In_1308);
nor U1876 (N_1876,In_1337,In_775);
nand U1877 (N_1877,In_1375,In_1925);
nor U1878 (N_1878,In_1121,In_1418);
or U1879 (N_1879,In_1910,In_46);
nand U1880 (N_1880,In_397,In_774);
nand U1881 (N_1881,In_850,In_649);
xnor U1882 (N_1882,In_1312,In_1607);
or U1883 (N_1883,In_542,In_1996);
xnor U1884 (N_1884,In_194,In_1392);
or U1885 (N_1885,In_1684,In_687);
or U1886 (N_1886,In_1763,In_1523);
and U1887 (N_1887,In_1405,In_7);
xor U1888 (N_1888,In_882,In_1219);
or U1889 (N_1889,In_1224,In_1487);
or U1890 (N_1890,In_1290,In_1790);
or U1891 (N_1891,In_1379,In_1700);
nand U1892 (N_1892,In_1817,In_1544);
nor U1893 (N_1893,In_1670,In_1118);
or U1894 (N_1894,In_733,In_1079);
or U1895 (N_1895,In_1923,In_1372);
nand U1896 (N_1896,In_69,In_702);
nand U1897 (N_1897,In_1709,In_597);
nand U1898 (N_1898,In_725,In_425);
nor U1899 (N_1899,In_1794,In_1773);
xnor U1900 (N_1900,In_1878,In_1512);
or U1901 (N_1901,In_1932,In_63);
or U1902 (N_1902,In_498,In_1697);
nand U1903 (N_1903,In_1238,In_160);
nand U1904 (N_1904,In_1632,In_1053);
nand U1905 (N_1905,In_1893,In_276);
xor U1906 (N_1906,In_962,In_106);
nand U1907 (N_1907,In_1485,In_607);
or U1908 (N_1908,In_1197,In_405);
xnor U1909 (N_1909,In_47,In_1722);
nor U1910 (N_1910,In_937,In_32);
nand U1911 (N_1911,In_1469,In_183);
xor U1912 (N_1912,In_229,In_372);
xnor U1913 (N_1913,In_1582,In_129);
xor U1914 (N_1914,In_97,In_787);
and U1915 (N_1915,In_1297,In_179);
and U1916 (N_1916,In_692,In_1320);
xnor U1917 (N_1917,In_1142,In_346);
nand U1918 (N_1918,In_1037,In_1333);
and U1919 (N_1919,In_1340,In_1911);
and U1920 (N_1920,In_135,In_1051);
nor U1921 (N_1921,In_1641,In_1718);
and U1922 (N_1922,In_1460,In_1559);
xnor U1923 (N_1923,In_1611,In_1005);
nor U1924 (N_1924,In_159,In_346);
xnor U1925 (N_1925,In_1991,In_692);
nor U1926 (N_1926,In_1995,In_588);
xor U1927 (N_1927,In_1208,In_91);
xor U1928 (N_1928,In_88,In_1853);
nor U1929 (N_1929,In_27,In_167);
xnor U1930 (N_1930,In_623,In_1743);
xor U1931 (N_1931,In_93,In_1226);
nand U1932 (N_1932,In_246,In_892);
xnor U1933 (N_1933,In_588,In_358);
nor U1934 (N_1934,In_1039,In_751);
or U1935 (N_1935,In_28,In_20);
nand U1936 (N_1936,In_590,In_1443);
or U1937 (N_1937,In_974,In_1923);
xnor U1938 (N_1938,In_343,In_1273);
nor U1939 (N_1939,In_1047,In_259);
or U1940 (N_1940,In_1417,In_349);
and U1941 (N_1941,In_425,In_1392);
and U1942 (N_1942,In_123,In_1966);
xor U1943 (N_1943,In_595,In_855);
nor U1944 (N_1944,In_1428,In_861);
nor U1945 (N_1945,In_1674,In_409);
and U1946 (N_1946,In_197,In_560);
or U1947 (N_1947,In_1378,In_631);
nand U1948 (N_1948,In_1575,In_1590);
and U1949 (N_1949,In_748,In_827);
xor U1950 (N_1950,In_1393,In_1567);
xnor U1951 (N_1951,In_670,In_744);
xor U1952 (N_1952,In_673,In_1933);
nand U1953 (N_1953,In_315,In_597);
nand U1954 (N_1954,In_110,In_464);
nand U1955 (N_1955,In_1632,In_1220);
xor U1956 (N_1956,In_75,In_280);
xor U1957 (N_1957,In_1222,In_520);
and U1958 (N_1958,In_1798,In_1309);
xor U1959 (N_1959,In_1320,In_1489);
or U1960 (N_1960,In_363,In_1148);
or U1961 (N_1961,In_1385,In_1638);
or U1962 (N_1962,In_598,In_1483);
nor U1963 (N_1963,In_1830,In_254);
nand U1964 (N_1964,In_374,In_1630);
xnor U1965 (N_1965,In_1825,In_1125);
and U1966 (N_1966,In_1424,In_1053);
or U1967 (N_1967,In_1381,In_487);
xnor U1968 (N_1968,In_1679,In_1657);
nor U1969 (N_1969,In_1750,In_1518);
and U1970 (N_1970,In_622,In_1995);
xnor U1971 (N_1971,In_1040,In_907);
xnor U1972 (N_1972,In_730,In_1717);
nand U1973 (N_1973,In_999,In_1028);
and U1974 (N_1974,In_1943,In_875);
and U1975 (N_1975,In_428,In_316);
nand U1976 (N_1976,In_1506,In_1236);
nor U1977 (N_1977,In_517,In_792);
nand U1978 (N_1978,In_17,In_1798);
and U1979 (N_1979,In_1207,In_167);
or U1980 (N_1980,In_138,In_1325);
nor U1981 (N_1981,In_2,In_80);
nand U1982 (N_1982,In_1058,In_1382);
nor U1983 (N_1983,In_486,In_1062);
and U1984 (N_1984,In_1943,In_114);
nand U1985 (N_1985,In_864,In_1171);
nor U1986 (N_1986,In_1767,In_1393);
and U1987 (N_1987,In_1340,In_103);
nand U1988 (N_1988,In_1230,In_710);
nor U1989 (N_1989,In_1301,In_178);
nor U1990 (N_1990,In_1198,In_225);
nand U1991 (N_1991,In_1215,In_135);
xnor U1992 (N_1992,In_1546,In_1214);
and U1993 (N_1993,In_287,In_1808);
nor U1994 (N_1994,In_1428,In_1282);
nor U1995 (N_1995,In_148,In_198);
nand U1996 (N_1996,In_1537,In_57);
and U1997 (N_1997,In_1904,In_162);
nand U1998 (N_1998,In_1779,In_1103);
or U1999 (N_1999,In_1375,In_341);
xnor U2000 (N_2000,N_501,N_1691);
nor U2001 (N_2001,N_1121,N_413);
and U2002 (N_2002,N_85,N_546);
nor U2003 (N_2003,N_1950,N_252);
xor U2004 (N_2004,N_1737,N_1171);
nand U2005 (N_2005,N_1647,N_536);
or U2006 (N_2006,N_830,N_207);
nand U2007 (N_2007,N_581,N_1142);
or U2008 (N_2008,N_677,N_1956);
xor U2009 (N_2009,N_353,N_1236);
nor U2010 (N_2010,N_580,N_1626);
or U2011 (N_2011,N_1746,N_1185);
nor U2012 (N_2012,N_1936,N_600);
xnor U2013 (N_2013,N_796,N_1814);
and U2014 (N_2014,N_720,N_807);
nand U2015 (N_2015,N_1187,N_545);
and U2016 (N_2016,N_1207,N_1643);
nand U2017 (N_2017,N_1095,N_1711);
and U2018 (N_2018,N_1369,N_923);
nand U2019 (N_2019,N_1281,N_1082);
nand U2020 (N_2020,N_103,N_1728);
xor U2021 (N_2021,N_524,N_775);
and U2022 (N_2022,N_575,N_648);
and U2023 (N_2023,N_907,N_1701);
nor U2024 (N_2024,N_506,N_1484);
and U2025 (N_2025,N_1973,N_334);
nor U2026 (N_2026,N_742,N_1926);
nand U2027 (N_2027,N_1325,N_1278);
and U2028 (N_2028,N_1940,N_990);
and U2029 (N_2029,N_1147,N_289);
xor U2030 (N_2030,N_1288,N_1388);
and U2031 (N_2031,N_1470,N_672);
or U2032 (N_2032,N_735,N_687);
nand U2033 (N_2033,N_1404,N_539);
nand U2034 (N_2034,N_1159,N_1262);
xnor U2035 (N_2035,N_588,N_1290);
nor U2036 (N_2036,N_194,N_29);
nand U2037 (N_2037,N_1745,N_1579);
and U2038 (N_2038,N_949,N_1552);
xor U2039 (N_2039,N_630,N_594);
and U2040 (N_2040,N_1461,N_351);
nor U2041 (N_2041,N_1893,N_1487);
and U2042 (N_2042,N_45,N_1047);
or U2043 (N_2043,N_809,N_920);
or U2044 (N_2044,N_360,N_939);
or U2045 (N_2045,N_1546,N_603);
nor U2046 (N_2046,N_248,N_965);
and U2047 (N_2047,N_265,N_1900);
nor U2048 (N_2048,N_340,N_1889);
and U2049 (N_2049,N_123,N_1638);
and U2050 (N_2050,N_684,N_179);
xor U2051 (N_2051,N_191,N_453);
and U2052 (N_2052,N_1359,N_499);
nor U2053 (N_2053,N_1577,N_1098);
and U2054 (N_2054,N_122,N_1747);
and U2055 (N_2055,N_81,N_1450);
nor U2056 (N_2056,N_1845,N_1216);
nor U2057 (N_2057,N_1406,N_1916);
and U2058 (N_2058,N_1316,N_683);
or U2059 (N_2059,N_619,N_1160);
and U2060 (N_2060,N_319,N_271);
nor U2061 (N_2061,N_864,N_1444);
or U2062 (N_2062,N_400,N_458);
xor U2063 (N_2063,N_889,N_228);
or U2064 (N_2064,N_1386,N_1205);
nand U2065 (N_2065,N_1093,N_1989);
nand U2066 (N_2066,N_1769,N_451);
nand U2067 (N_2067,N_92,N_640);
nand U2068 (N_2068,N_1773,N_798);
or U2069 (N_2069,N_1367,N_840);
nand U2070 (N_2070,N_329,N_1542);
or U2071 (N_2071,N_1016,N_423);
and U2072 (N_2072,N_1913,N_598);
nor U2073 (N_2073,N_1471,N_788);
and U2074 (N_2074,N_1472,N_1741);
nand U2075 (N_2075,N_674,N_1592);
and U2076 (N_2076,N_1602,N_1932);
nand U2077 (N_2077,N_1644,N_1529);
and U2078 (N_2078,N_1279,N_1310);
and U2079 (N_2079,N_1108,N_11);
and U2080 (N_2080,N_1284,N_645);
nor U2081 (N_2081,N_877,N_1547);
and U2082 (N_2082,N_1374,N_1693);
nor U2083 (N_2083,N_1850,N_251);
and U2084 (N_2084,N_1757,N_1738);
nand U2085 (N_2085,N_18,N_1242);
or U2086 (N_2086,N_1699,N_1849);
nor U2087 (N_2087,N_415,N_697);
or U2088 (N_2088,N_379,N_666);
or U2089 (N_2089,N_430,N_766);
nand U2090 (N_2090,N_1661,N_716);
xor U2091 (N_2091,N_673,N_1537);
nand U2092 (N_2092,N_309,N_240);
nor U2093 (N_2093,N_1062,N_82);
nor U2094 (N_2094,N_1212,N_1154);
nor U2095 (N_2095,N_1189,N_343);
xor U2096 (N_2096,N_586,N_1518);
or U2097 (N_2097,N_1939,N_1040);
or U2098 (N_2098,N_1830,N_1117);
or U2099 (N_2099,N_471,N_1097);
and U2100 (N_2100,N_472,N_647);
and U2101 (N_2101,N_924,N_1128);
and U2102 (N_2102,N_442,N_1963);
and U2103 (N_2103,N_690,N_1213);
and U2104 (N_2104,N_181,N_771);
and U2105 (N_2105,N_900,N_1767);
or U2106 (N_2106,N_1899,N_1530);
and U2107 (N_2107,N_161,N_560);
or U2108 (N_2108,N_217,N_1502);
or U2109 (N_2109,N_960,N_14);
nor U2110 (N_2110,N_977,N_1750);
and U2111 (N_2111,N_48,N_1138);
and U2112 (N_2112,N_660,N_1516);
nand U2113 (N_2113,N_1658,N_367);
xor U2114 (N_2114,N_1864,N_427);
nor U2115 (N_2115,N_1796,N_1352);
nor U2116 (N_2116,N_1494,N_1424);
nor U2117 (N_2117,N_371,N_1775);
or U2118 (N_2118,N_1209,N_406);
nor U2119 (N_2119,N_1968,N_1026);
and U2120 (N_2120,N_1944,N_267);
nand U2121 (N_2121,N_1176,N_1140);
xnor U2122 (N_2122,N_63,N_1166);
nor U2123 (N_2123,N_268,N_528);
and U2124 (N_2124,N_1858,N_419);
nor U2125 (N_2125,N_153,N_1930);
xor U2126 (N_2126,N_1645,N_88);
nand U2127 (N_2127,N_314,N_3);
or U2128 (N_2128,N_617,N_1824);
and U2129 (N_2129,N_1457,N_1332);
nor U2130 (N_2130,N_1490,N_159);
or U2131 (N_2131,N_348,N_1178);
and U2132 (N_2132,N_1198,N_1555);
and U2133 (N_2133,N_172,N_1965);
nand U2134 (N_2134,N_327,N_304);
and U2135 (N_2135,N_548,N_1448);
and U2136 (N_2136,N_881,N_287);
xnor U2137 (N_2137,N_1749,N_538);
or U2138 (N_2138,N_1050,N_346);
nand U2139 (N_2139,N_175,N_1036);
nand U2140 (N_2140,N_1659,N_1463);
nand U2141 (N_2141,N_1334,N_1823);
and U2142 (N_2142,N_1941,N_701);
nand U2143 (N_2143,N_650,N_1066);
nor U2144 (N_2144,N_1868,N_740);
xnor U2145 (N_2145,N_782,N_791);
xnor U2146 (N_2146,N_296,N_1425);
nor U2147 (N_2147,N_714,N_370);
nor U2148 (N_2148,N_1718,N_1254);
or U2149 (N_2149,N_438,N_1832);
nand U2150 (N_2150,N_1072,N_1030);
nor U2151 (N_2151,N_1937,N_531);
xnor U2152 (N_2152,N_845,N_613);
nor U2153 (N_2153,N_917,N_1104);
or U2154 (N_2154,N_1075,N_283);
nand U2155 (N_2155,N_60,N_955);
nor U2156 (N_2156,N_237,N_58);
or U2157 (N_2157,N_71,N_250);
xor U2158 (N_2158,N_1363,N_829);
nand U2159 (N_2159,N_760,N_1045);
and U2160 (N_2160,N_986,N_678);
xor U2161 (N_2161,N_1979,N_1583);
and U2162 (N_2162,N_1617,N_285);
xor U2163 (N_2163,N_868,N_106);
nor U2164 (N_2164,N_1019,N_1194);
and U2165 (N_2165,N_1841,N_1318);
and U2166 (N_2166,N_1083,N_1111);
nand U2167 (N_2167,N_1788,N_860);
and U2168 (N_2168,N_1720,N_1096);
xor U2169 (N_2169,N_102,N_204);
and U2170 (N_2170,N_457,N_1287);
or U2171 (N_2171,N_1231,N_785);
xor U2172 (N_2172,N_1536,N_350);
xnor U2173 (N_2173,N_757,N_1986);
xnor U2174 (N_2174,N_230,N_1412);
nor U2175 (N_2175,N_133,N_1498);
and U2176 (N_2176,N_83,N_1984);
nor U2177 (N_2177,N_1311,N_1253);
or U2178 (N_2178,N_1183,N_361);
nand U2179 (N_2179,N_1032,N_1002);
or U2180 (N_2180,N_165,N_330);
xnor U2181 (N_2181,N_295,N_381);
and U2182 (N_2182,N_246,N_1430);
or U2183 (N_2183,N_1501,N_1283);
and U2184 (N_2184,N_837,N_797);
nor U2185 (N_2185,N_1298,N_1884);
nor U2186 (N_2186,N_447,N_292);
xor U2187 (N_2187,N_1517,N_364);
or U2188 (N_2188,N_1250,N_119);
and U2189 (N_2189,N_1006,N_1679);
or U2190 (N_2190,N_728,N_68);
and U2191 (N_2191,N_1714,N_562);
and U2192 (N_2192,N_1486,N_1709);
or U2193 (N_2193,N_424,N_389);
xnor U2194 (N_2194,N_28,N_1504);
nor U2195 (N_2195,N_1996,N_543);
or U2196 (N_2196,N_1058,N_1249);
nand U2197 (N_2197,N_1867,N_1317);
and U2198 (N_2198,N_1791,N_1204);
nand U2199 (N_2199,N_1987,N_320);
nand U2200 (N_2200,N_1308,N_1015);
nand U2201 (N_2201,N_1416,N_1948);
or U2202 (N_2202,N_518,N_527);
xnor U2203 (N_2203,N_599,N_1629);
nor U2204 (N_2204,N_1831,N_131);
xor U2205 (N_2205,N_890,N_614);
or U2206 (N_2206,N_156,N_115);
and U2207 (N_2207,N_95,N_944);
nor U2208 (N_2208,N_1698,N_850);
xnor U2209 (N_2209,N_951,N_1958);
nor U2210 (N_2210,N_1835,N_1088);
nand U2211 (N_2211,N_504,N_1202);
xnor U2212 (N_2212,N_316,N_1593);
nor U2213 (N_2213,N_1551,N_905);
nor U2214 (N_2214,N_956,N_1632);
or U2215 (N_2215,N_1263,N_1631);
and U2216 (N_2216,N_1109,N_1506);
nand U2217 (N_2217,N_1677,N_1982);
nor U2218 (N_2218,N_1268,N_1947);
nor U2219 (N_2219,N_1710,N_1765);
or U2220 (N_2220,N_1783,N_260);
xnor U2221 (N_2221,N_1708,N_769);
or U2222 (N_2222,N_460,N_974);
nor U2223 (N_2223,N_987,N_27);
nand U2224 (N_2224,N_224,N_1619);
nand U2225 (N_2225,N_689,N_1715);
and U2226 (N_2226,N_1481,N_628);
nand U2227 (N_2227,N_1116,N_382);
nand U2228 (N_2228,N_1942,N_1507);
nand U2229 (N_2229,N_901,N_1586);
xor U2230 (N_2230,N_903,N_1873);
nand U2231 (N_2231,N_152,N_1851);
and U2232 (N_2232,N_989,N_1614);
nor U2233 (N_2233,N_421,N_305);
or U2234 (N_2234,N_1524,N_1923);
xnor U2235 (N_2235,N_62,N_1641);
and U2236 (N_2236,N_121,N_491);
nand U2237 (N_2237,N_915,N_1820);
nor U2238 (N_2238,N_1400,N_469);
xnor U2239 (N_2239,N_1269,N_1427);
nand U2240 (N_2240,N_595,N_1459);
nand U2241 (N_2241,N_236,N_759);
xnor U2242 (N_2242,N_1819,N_1396);
nand U2243 (N_2243,N_863,N_1785);
xnor U2244 (N_2244,N_1571,N_711);
nor U2245 (N_2245,N_885,N_1742);
nor U2246 (N_2246,N_1856,N_1456);
nor U2247 (N_2247,N_1548,N_146);
nor U2248 (N_2248,N_1473,N_585);
nor U2249 (N_2249,N_1782,N_686);
xor U2250 (N_2250,N_433,N_1000);
nand U2251 (N_2251,N_1964,N_1566);
and U2252 (N_2252,N_1008,N_1346);
or U2253 (N_2253,N_904,N_1779);
nor U2254 (N_2254,N_459,N_922);
nand U2255 (N_2255,N_1642,N_164);
nor U2256 (N_2256,N_1112,N_1795);
or U2257 (N_2257,N_448,N_1553);
nor U2258 (N_2258,N_827,N_216);
xor U2259 (N_2259,N_1280,N_1696);
or U2260 (N_2260,N_1199,N_263);
nand U2261 (N_2261,N_804,N_635);
and U2262 (N_2262,N_13,N_806);
nand U2263 (N_2263,N_679,N_331);
xnor U2264 (N_2264,N_1053,N_1309);
nor U2265 (N_2265,N_1220,N_1059);
nand U2266 (N_2266,N_1376,N_532);
and U2267 (N_2267,N_157,N_128);
nor U2268 (N_2268,N_1405,N_1465);
or U2269 (N_2269,N_644,N_1667);
nand U2270 (N_2270,N_247,N_652);
or U2271 (N_2271,N_50,N_90);
xnor U2272 (N_2272,N_1181,N_39);
nor U2273 (N_2273,N_938,N_975);
xor U2274 (N_2274,N_838,N_129);
nand U2275 (N_2275,N_241,N_1458);
or U2276 (N_2276,N_1482,N_789);
nand U2277 (N_2277,N_1760,N_231);
or U2278 (N_2278,N_778,N_1364);
nand U2279 (N_2279,N_1578,N_872);
nor U2280 (N_2280,N_219,N_76);
nor U2281 (N_2281,N_188,N_468);
nor U2282 (N_2282,N_390,N_1957);
or U2283 (N_2283,N_773,N_1521);
nor U2284 (N_2284,N_276,N_1028);
nor U2285 (N_2285,N_1843,N_530);
nor U2286 (N_2286,N_1025,N_1252);
and U2287 (N_2287,N_751,N_1303);
xor U2288 (N_2288,N_1129,N_1248);
nand U2289 (N_2289,N_1727,N_1024);
or U2290 (N_2290,N_1432,N_908);
xor U2291 (N_2291,N_1929,N_473);
or U2292 (N_2292,N_1037,N_1127);
nor U2293 (N_2293,N_1612,N_1387);
and U2294 (N_2294,N_764,N_859);
nand U2295 (N_2295,N_1861,N_49);
xnor U2296 (N_2296,N_811,N_1685);
xor U2297 (N_2297,N_482,N_197);
or U2298 (N_2298,N_1124,N_1651);
or U2299 (N_2299,N_694,N_358);
or U2300 (N_2300,N_0,N_1620);
nor U2301 (N_2301,N_1161,N_1020);
or U2302 (N_2302,N_1665,N_793);
nand U2303 (N_2303,N_1225,N_952);
and U2304 (N_2304,N_277,N_1206);
or U2305 (N_2305,N_886,N_344);
xnor U2306 (N_2306,N_368,N_1927);
xnor U2307 (N_2307,N_1240,N_713);
or U2308 (N_2308,N_947,N_1801);
and U2309 (N_2309,N_1569,N_1561);
or U2310 (N_2310,N_1800,N_308);
or U2311 (N_2311,N_323,N_772);
nor U2312 (N_2312,N_608,N_1385);
or U2313 (N_2313,N_1389,N_1525);
and U2314 (N_2314,N_1196,N_1348);
xnor U2315 (N_2315,N_437,N_1492);
nor U2316 (N_2316,N_547,N_1258);
and U2317 (N_2317,N_1474,N_1134);
nand U2318 (N_2318,N_1192,N_1485);
or U2319 (N_2319,N_1234,N_1879);
nand U2320 (N_2320,N_998,N_591);
nor U2321 (N_2321,N_656,N_383);
nand U2322 (N_2322,N_155,N_297);
and U2323 (N_2323,N_1704,N_784);
or U2324 (N_2324,N_1604,N_220);
and U2325 (N_2325,N_754,N_89);
nand U2326 (N_2326,N_1145,N_1829);
nand U2327 (N_2327,N_1155,N_1780);
nor U2328 (N_2328,N_592,N_1195);
nor U2329 (N_2329,N_865,N_681);
nor U2330 (N_2330,N_1863,N_1331);
and U2331 (N_2331,N_670,N_46);
nand U2332 (N_2332,N_512,N_120);
xor U2333 (N_2333,N_1764,N_1132);
nand U2334 (N_2334,N_1513,N_177);
nand U2335 (N_2335,N_1866,N_1908);
nor U2336 (N_2336,N_661,N_1018);
and U2337 (N_2337,N_1345,N_1886);
xnor U2338 (N_2338,N_1454,N_441);
nor U2339 (N_2339,N_1022,N_313);
xor U2340 (N_2340,N_1426,N_577);
and U2341 (N_2341,N_291,N_258);
and U2342 (N_2342,N_335,N_1713);
nand U2343 (N_2343,N_1343,N_1811);
nand U2344 (N_2344,N_19,N_1029);
or U2345 (N_2345,N_1907,N_481);
nand U2346 (N_2346,N_34,N_1241);
and U2347 (N_2347,N_1271,N_1390);
and U2348 (N_2348,N_1141,N_1918);
or U2349 (N_2349,N_1557,N_1478);
nand U2350 (N_2350,N_1625,N_51);
and U2351 (N_2351,N_208,N_1429);
or U2352 (N_2352,N_253,N_1293);
or U2353 (N_2353,N_405,N_16);
nor U2354 (N_2354,N_1081,N_1071);
or U2355 (N_2355,N_1894,N_824);
or U2356 (N_2356,N_787,N_633);
and U2357 (N_2357,N_629,N_1113);
nand U2358 (N_2358,N_288,N_777);
or U2359 (N_2359,N_734,N_1330);
nand U2360 (N_2360,N_573,N_521);
and U2361 (N_2361,N_410,N_1323);
nand U2362 (N_2362,N_636,N_583);
xnor U2363 (N_2363,N_1333,N_1914);
and U2364 (N_2364,N_1902,N_269);
or U2365 (N_2365,N_1251,N_104);
nor U2366 (N_2366,N_213,N_6);
nor U2367 (N_2367,N_1671,N_1462);
and U2368 (N_2368,N_1859,N_856);
xnor U2369 (N_2369,N_32,N_456);
xnor U2370 (N_2370,N_823,N_1852);
and U2371 (N_2371,N_602,N_941);
and U2372 (N_2372,N_1574,N_495);
nand U2373 (N_2373,N_202,N_1981);
nor U2374 (N_2374,N_394,N_1174);
nor U2375 (N_2375,N_178,N_620);
or U2376 (N_2376,N_1590,N_653);
nand U2377 (N_2377,N_609,N_420);
and U2378 (N_2378,N_893,N_507);
nand U2379 (N_2379,N_779,N_215);
and U2380 (N_2380,N_1131,N_1943);
and U2381 (N_2381,N_273,N_554);
or U2382 (N_2382,N_1226,N_1934);
nand U2383 (N_2383,N_384,N_1118);
and U2384 (N_2384,N_1148,N_1799);
and U2385 (N_2385,N_557,N_1666);
and U2386 (N_2386,N_218,N_1621);
xnor U2387 (N_2387,N_470,N_1273);
nand U2388 (N_2388,N_1158,N_1535);
nor U2389 (N_2389,N_388,N_1301);
or U2390 (N_2390,N_1599,N_1003);
xor U2391 (N_2391,N_1522,N_800);
nor U2392 (N_2392,N_259,N_933);
nand U2393 (N_2393,N_1222,N_1255);
nand U2394 (N_2394,N_526,N_1825);
xnor U2395 (N_2395,N_869,N_357);
nand U2396 (N_2396,N_1978,N_1208);
or U2397 (N_2397,N_1689,N_1437);
and U2398 (N_2398,N_1550,N_1730);
or U2399 (N_2399,N_302,N_963);
and U2400 (N_2400,N_1828,N_1881);
nor U2401 (N_2401,N_38,N_972);
nor U2402 (N_2402,N_780,N_712);
nand U2403 (N_2403,N_1692,N_663);
nor U2404 (N_2404,N_930,N_736);
nand U2405 (N_2405,N_107,N_1275);
nor U2406 (N_2406,N_946,N_1959);
or U2407 (N_2407,N_244,N_1077);
xor U2408 (N_2408,N_511,N_480);
or U2409 (N_2409,N_568,N_347);
nand U2410 (N_2410,N_1186,N_988);
and U2411 (N_2411,N_127,N_173);
nor U2412 (N_2412,N_1669,N_733);
and U2413 (N_2413,N_132,N_746);
xnor U2414 (N_2414,N_688,N_1057);
nor U2415 (N_2415,N_1493,N_1549);
nor U2416 (N_2416,N_981,N_1805);
nand U2417 (N_2417,N_1300,N_1193);
or U2418 (N_2418,N_1114,N_1598);
xnor U2419 (N_2419,N_414,N_1105);
nor U2420 (N_2420,N_293,N_1101);
and U2421 (N_2421,N_1999,N_659);
nand U2422 (N_2422,N_488,N_730);
or U2423 (N_2423,N_928,N_1230);
nand U2424 (N_2424,N_1778,N_916);
or U2425 (N_2425,N_918,N_1684);
and U2426 (N_2426,N_294,N_1657);
nand U2427 (N_2427,N_639,N_391);
or U2428 (N_2428,N_1813,N_676);
or U2429 (N_2429,N_738,N_1371);
and U2430 (N_2430,N_959,N_1452);
nor U2431 (N_2431,N_832,N_1379);
or U2432 (N_2432,N_186,N_238);
nand U2433 (N_2433,N_1515,N_1312);
nand U2434 (N_2434,N_1688,N_729);
or U2435 (N_2435,N_1170,N_1403);
and U2436 (N_2436,N_396,N_1664);
nand U2437 (N_2437,N_1554,N_611);
nor U2438 (N_2438,N_53,N_1086);
xnor U2439 (N_2439,N_1774,N_1409);
nor U2440 (N_2440,N_820,N_925);
nand U2441 (N_2441,N_1144,N_1172);
nand U2442 (N_2442,N_449,N_1512);
nor U2443 (N_2443,N_1428,N_1357);
xnor U2444 (N_2444,N_1997,N_770);
nand U2445 (N_2445,N_1453,N_1177);
or U2446 (N_2446,N_1672,N_372);
and U2447 (N_2447,N_1998,N_1257);
nand U2448 (N_2448,N_1010,N_1286);
nor U2449 (N_2449,N_1675,N_851);
and U2450 (N_2450,N_1653,N_1609);
or U2451 (N_2451,N_1434,N_1270);
xor U2452 (N_2452,N_1798,N_1243);
nand U2453 (N_2453,N_1702,N_803);
xor U2454 (N_2454,N_1421,N_440);
nand U2455 (N_2455,N_1697,N_1060);
nor U2456 (N_2456,N_1683,N_1377);
or U2457 (N_2457,N_1534,N_1680);
nor U2458 (N_2458,N_279,N_1256);
and U2459 (N_2459,N_1344,N_1051);
and U2460 (N_2460,N_802,N_1139);
nand U2461 (N_2461,N_1505,N_66);
nand U2462 (N_2462,N_1038,N_641);
or U2463 (N_2463,N_1510,N_1857);
nand U2464 (N_2464,N_108,N_1260);
xnor U2465 (N_2465,N_529,N_1787);
and U2466 (N_2466,N_921,N_1564);
xor U2467 (N_2467,N_227,N_514);
nor U2468 (N_2468,N_597,N_5);
nand U2469 (N_2469,N_64,N_25);
nor U2470 (N_2470,N_604,N_1871);
xnor U2471 (N_2471,N_544,N_362);
nor U2472 (N_2472,N_1721,N_849);
nand U2473 (N_2473,N_1356,N_1776);
nand U2474 (N_2474,N_1495,N_1074);
nor U2475 (N_2475,N_1235,N_882);
or U2476 (N_2476,N_707,N_731);
nand U2477 (N_2477,N_1499,N_1967);
and U2478 (N_2478,N_1210,N_858);
xnor U2479 (N_2479,N_1267,N_1608);
xnor U2480 (N_2480,N_1878,N_632);
or U2481 (N_2481,N_1993,N_1203);
and U2482 (N_2482,N_1735,N_750);
xor U2483 (N_2483,N_1781,N_338);
and U2484 (N_2484,N_1565,N_919);
and U2485 (N_2485,N_80,N_439);
xor U2486 (N_2486,N_1758,N_337);
and U2487 (N_2487,N_718,N_968);
xnor U2488 (N_2488,N_1855,N_626);
nand U2489 (N_2489,N_4,N_428);
nand U2490 (N_2490,N_958,N_638);
and U2491 (N_2491,N_1084,N_786);
nor U2492 (N_2492,N_664,N_307);
xnor U2493 (N_2493,N_256,N_1337);
xnor U2494 (N_2494,N_1366,N_559);
xor U2495 (N_2495,N_1360,N_1951);
xnor U2496 (N_2496,N_398,N_758);
and U2497 (N_2497,N_1136,N_1572);
xnor U2498 (N_2498,N_884,N_699);
and U2499 (N_2499,N_1872,N_1476);
nor U2500 (N_2500,N_1520,N_333);
or U2501 (N_2501,N_342,N_945);
or U2502 (N_2502,N_1706,N_854);
xnor U2503 (N_2503,N_813,N_446);
or U2504 (N_2504,N_1743,N_1324);
nand U2505 (N_2505,N_1162,N_1305);
nor U2506 (N_2506,N_79,N_1440);
or U2507 (N_2507,N_1443,N_1729);
nand U2508 (N_2508,N_281,N_596);
xor U2509 (N_2509,N_1860,N_214);
nor U2510 (N_2510,N_1532,N_1446);
nand U2511 (N_2511,N_489,N_1837);
xor U2512 (N_2512,N_1351,N_206);
nand U2513 (N_2513,N_593,N_322);
nor U2514 (N_2514,N_205,N_1107);
nand U2515 (N_2515,N_1137,N_1687);
nand U2516 (N_2516,N_1314,N_634);
nor U2517 (N_2517,N_1091,N_817);
and U2518 (N_2518,N_1413,N_221);
xor U2519 (N_2519,N_210,N_1992);
xor U2520 (N_2520,N_1526,N_290);
nor U2521 (N_2521,N_136,N_1021);
nor U2522 (N_2522,N_739,N_1616);
nor U2523 (N_2523,N_1588,N_1771);
or U2524 (N_2524,N_1920,N_1630);
nand U2525 (N_2525,N_1748,N_1069);
xnor U2526 (N_2526,N_341,N_101);
or U2527 (N_2527,N_1282,N_1399);
xor U2528 (N_2528,N_1808,N_935);
xnor U2529 (N_2529,N_801,N_429);
xnor U2530 (N_2530,N_970,N_1078);
nand U2531 (N_2531,N_1422,N_143);
xor U2532 (N_2532,N_971,N_300);
and U2533 (N_2533,N_1793,N_1042);
nand U2534 (N_2534,N_812,N_56);
nand U2535 (N_2535,N_1328,N_35);
nor U2536 (N_2536,N_1394,N_1650);
or U2537 (N_2537,N_962,N_936);
and U2538 (N_2538,N_1342,N_748);
xnor U2539 (N_2539,N_141,N_318);
nor U2540 (N_2540,N_436,N_1533);
nand U2541 (N_2541,N_485,N_1772);
and U2542 (N_2542,N_1633,N_658);
and U2543 (N_2543,N_995,N_1906);
and U2544 (N_2544,N_225,N_193);
and U2545 (N_2545,N_1544,N_710);
or U2546 (N_2546,N_510,N_1438);
nor U2547 (N_2547,N_1110,N_1954);
xnor U2548 (N_2548,N_1,N_1905);
and U2549 (N_2549,N_1976,N_1232);
nand U2550 (N_2550,N_1646,N_1807);
xnor U2551 (N_2551,N_1049,N_1163);
nand U2552 (N_2552,N_1023,N_1289);
nand U2553 (N_2553,N_1180,N_1971);
nand U2554 (N_2554,N_1043,N_397);
nand U2555 (N_2555,N_280,N_47);
xnor U2556 (N_2556,N_148,N_715);
xnor U2557 (N_2557,N_1120,N_590);
nor U2558 (N_2558,N_444,N_558);
nor U2559 (N_2559,N_891,N_983);
nand U2560 (N_2560,N_375,N_498);
nand U2561 (N_2561,N_815,N_36);
nand U2562 (N_2562,N_118,N_1191);
and U2563 (N_2563,N_1378,N_1883);
and U2564 (N_2564,N_753,N_1960);
nand U2565 (N_2565,N_825,N_953);
xor U2566 (N_2566,N_1740,N_2);
and U2567 (N_2567,N_1563,N_1392);
nor U2568 (N_2568,N_1087,N_870);
xor U2569 (N_2569,N_732,N_1681);
xnor U2570 (N_2570,N_483,N_1261);
or U2571 (N_2571,N_1817,N_1909);
nand U2572 (N_2572,N_1703,N_1523);
xnor U2573 (N_2573,N_929,N_435);
and U2574 (N_2574,N_487,N_1962);
and U2575 (N_2575,N_363,N_387);
xor U2576 (N_2576,N_902,N_717);
nand U2577 (N_2577,N_654,N_112);
and U2578 (N_2578,N_403,N_187);
nand U2579 (N_2579,N_31,N_1734);
nor U2580 (N_2580,N_1833,N_10);
xor U2581 (N_2581,N_1338,N_1414);
nor U2582 (N_2582,N_571,N_1445);
nor U2583 (N_2583,N_747,N_1297);
or U2584 (N_2584,N_1167,N_326);
and U2585 (N_2585,N_892,N_1731);
nor U2586 (N_2586,N_899,N_1576);
nor U2587 (N_2587,N_1794,N_254);
nand U2588 (N_2588,N_1862,N_1827);
nor U2589 (N_2589,N_9,N_655);
nand U2590 (N_2590,N_1919,N_484);
nand U2591 (N_2591,N_174,N_1613);
and U2592 (N_2592,N_1953,N_1594);
xor U2593 (N_2593,N_1441,N_1244);
nor U2594 (N_2594,N_450,N_576);
and U2595 (N_2595,N_519,N_1726);
xor U2596 (N_2596,N_567,N_418);
or U2597 (N_2597,N_744,N_7);
or U2598 (N_2598,N_328,N_631);
and U2599 (N_2599,N_1068,N_1844);
and U2600 (N_2600,N_1295,N_623);
or U2601 (N_2601,N_98,N_73);
nand U2602 (N_2602,N_1307,N_392);
nand U2603 (N_2603,N_1239,N_1722);
and U2604 (N_2604,N_474,N_783);
xnor U2605 (N_2605,N_142,N_1277);
nor U2606 (N_2606,N_1717,N_1079);
nor U2607 (N_2607,N_1690,N_607);
and U2608 (N_2608,N_625,N_1603);
and U2609 (N_2609,N_1218,N_1756);
xnor U2610 (N_2610,N_1201,N_1393);
or U2611 (N_2611,N_1509,N_1488);
nor U2612 (N_2612,N_1925,N_702);
and U2613 (N_2613,N_467,N_1211);
nor U2614 (N_2614,N_8,N_266);
nand U2615 (N_2615,N_426,N_934);
or U2616 (N_2616,N_1395,N_564);
xor U2617 (N_2617,N_286,N_1173);
or U2618 (N_2618,N_502,N_1190);
or U2619 (N_2619,N_229,N_1373);
and U2620 (N_2620,N_84,N_1977);
nand U2621 (N_2621,N_1678,N_1700);
and U2622 (N_2622,N_1660,N_359);
xor U2623 (N_2623,N_1073,N_33);
or U2624 (N_2624,N_1875,N_1065);
nor U2625 (N_2625,N_665,N_234);
or U2626 (N_2626,N_1924,N_967);
nor U2627 (N_2627,N_792,N_570);
xor U2628 (N_2628,N_703,N_349);
nand U2629 (N_2629,N_883,N_853);
nor U2630 (N_2630,N_727,N_726);
nor U2631 (N_2631,N_494,N_1475);
and U2632 (N_2632,N_855,N_1739);
nand U2633 (N_2633,N_1970,N_1156);
nand U2634 (N_2634,N_1877,N_584);
nor U2635 (N_2635,N_1600,N_794);
and U2636 (N_2636,N_1326,N_605);
nor U2637 (N_2637,N_432,N_799);
nand U2638 (N_2638,N_722,N_755);
nor U2639 (N_2639,N_1623,N_1662);
nand U2640 (N_2640,N_1407,N_980);
nor U2641 (N_2641,N_1179,N_1272);
xor U2642 (N_2642,N_669,N_416);
and U2643 (N_2643,N_301,N_1611);
xor U2644 (N_2644,N_601,N_737);
nor U2645 (N_2645,N_1165,N_503);
xor U2646 (N_2646,N_1933,N_41);
xor U2647 (N_2647,N_662,N_325);
and U2648 (N_2648,N_52,N_1723);
and U2649 (N_2649,N_190,N_1415);
or U2650 (N_2650,N_1418,N_1848);
nor U2651 (N_2651,N_1126,N_1238);
nor U2652 (N_2652,N_1792,N_1763);
and U2653 (N_2653,N_1840,N_704);
xnor U2654 (N_2654,N_1966,N_1264);
or U2655 (N_2655,N_861,N_1339);
xor U2656 (N_2656,N_1246,N_1797);
nand U2657 (N_2657,N_1319,N_114);
nor U2658 (N_2658,N_1912,N_741);
and U2659 (N_2659,N_54,N_1988);
and U2660 (N_2660,N_1686,N_1768);
or U2661 (N_2661,N_695,N_111);
or U2662 (N_2662,N_589,N_158);
nand U2663 (N_2663,N_709,N_1184);
and U2664 (N_2664,N_1115,N_1067);
nand U2665 (N_2665,N_1541,N_492);
or U2666 (N_2666,N_790,N_1668);
nor U2667 (N_2667,N_1274,N_1080);
nor U2668 (N_2668,N_1663,N_805);
xor U2669 (N_2669,N_1995,N_866);
and U2670 (N_2670,N_1119,N_1595);
or U2671 (N_2671,N_756,N_270);
and U2672 (N_2672,N_1766,N_1839);
and U2673 (N_2673,N_875,N_183);
xor U2674 (N_2674,N_1527,N_1655);
xnor U2675 (N_2675,N_643,N_366);
or U2676 (N_2676,N_948,N_1188);
or U2677 (N_2677,N_169,N_1233);
and U2678 (N_2678,N_1955,N_982);
xnor U2679 (N_2679,N_1439,N_1508);
and U2680 (N_2680,N_1391,N_950);
xnor U2681 (N_2681,N_1935,N_1804);
nor U2682 (N_2682,N_407,N_1175);
nand U2683 (N_2683,N_1581,N_541);
nand U2684 (N_2684,N_465,N_749);
nor U2685 (N_2685,N_380,N_176);
xor U2686 (N_2686,N_1152,N_781);
nand U2687 (N_2687,N_1511,N_1648);
nor U2688 (N_2688,N_1123,N_1398);
or U2689 (N_2689,N_1011,N_1085);
or U2690 (N_2690,N_937,N_816);
and U2691 (N_2691,N_1514,N_1622);
nor U2692 (N_2692,N_1168,N_154);
or U2693 (N_2693,N_226,N_1146);
or U2694 (N_2694,N_1538,N_1401);
nor U2695 (N_2695,N_233,N_841);
xor U2696 (N_2696,N_1063,N_513);
and U2697 (N_2697,N_914,N_235);
nand U2698 (N_2698,N_262,N_535);
or U2699 (N_2699,N_606,N_464);
and U2700 (N_2700,N_1054,N_839);
and U2701 (N_2701,N_957,N_1903);
and U2702 (N_2702,N_1436,N_1358);
nor U2703 (N_2703,N_500,N_160);
xnor U2704 (N_2704,N_693,N_393);
or U2705 (N_2705,N_91,N_525);
or U2706 (N_2706,N_618,N_1150);
and U2707 (N_2707,N_1382,N_795);
xnor U2708 (N_2708,N_835,N_167);
nand U2709 (N_2709,N_834,N_1296);
or U2710 (N_2710,N_126,N_1014);
nor U2711 (N_2711,N_1607,N_1229);
xnor U2712 (N_2712,N_1122,N_1460);
and U2713 (N_2713,N_1135,N_516);
and U2714 (N_2714,N_552,N_1975);
and U2715 (N_2715,N_1946,N_1094);
nand U2716 (N_2716,N_1431,N_1215);
nand U2717 (N_2717,N_1634,N_1573);
or U2718 (N_2718,N_1876,N_1483);
xnor U2719 (N_2719,N_1313,N_1217);
and U2720 (N_2720,N_299,N_1707);
and U2721 (N_2721,N_1355,N_551);
or U2722 (N_2722,N_1911,N_1895);
and U2723 (N_2723,N_1896,N_961);
nand U2724 (N_2724,N_1469,N_125);
and U2725 (N_2725,N_321,N_198);
nand U2726 (N_2726,N_211,N_26);
xnor U2727 (N_2727,N_1724,N_743);
xor U2728 (N_2728,N_1285,N_1102);
nand U2729 (N_2729,N_1901,N_1562);
or U2730 (N_2730,N_408,N_1372);
nor U2731 (N_2731,N_1100,N_1853);
nor U2732 (N_2732,N_355,N_1882);
xor U2733 (N_2733,N_1846,N_1103);
nor U2734 (N_2734,N_976,N_232);
and U2735 (N_2735,N_1725,N_1606);
and U2736 (N_2736,N_1005,N_1556);
nand U2737 (N_2737,N_894,N_1004);
and U2738 (N_2738,N_249,N_1013);
nand U2739 (N_2739,N_404,N_1812);
nor U2740 (N_2740,N_195,N_651);
nand U2741 (N_2741,N_984,N_1985);
and U2742 (N_2742,N_1567,N_100);
xnor U2743 (N_2743,N_1803,N_828);
nand U2744 (N_2744,N_1802,N_1874);
or U2745 (N_2745,N_691,N_462);
and U2746 (N_2746,N_569,N_151);
xnor U2747 (N_2747,N_1245,N_831);
nor U2748 (N_2748,N_1869,N_1751);
nor U2749 (N_2749,N_565,N_365);
or U2750 (N_2750,N_1375,N_1336);
or U2751 (N_2751,N_455,N_1670);
or U2752 (N_2752,N_1676,N_72);
or U2753 (N_2753,N_1898,N_1639);
and U2754 (N_2754,N_1048,N_324);
nand U2755 (N_2755,N_385,N_994);
nor U2756 (N_2756,N_264,N_1716);
xnor U2757 (N_2757,N_200,N_675);
or U2758 (N_2758,N_610,N_1682);
and U2759 (N_2759,N_411,N_1784);
nand U2760 (N_2760,N_1640,N_1361);
and U2761 (N_2761,N_843,N_409);
xor U2762 (N_2762,N_1627,N_1834);
and U2763 (N_2763,N_1007,N_616);
or U2764 (N_2764,N_445,N_110);
xnor U2765 (N_2765,N_1052,N_1027);
or U2766 (N_2766,N_1945,N_1182);
nor U2767 (N_2767,N_1321,N_574);
nor U2768 (N_2768,N_1322,N_21);
or U2769 (N_2769,N_1605,N_637);
and U2770 (N_2770,N_1610,N_87);
nor U2771 (N_2771,N_24,N_1247);
nand U2772 (N_2772,N_1214,N_555);
and U2773 (N_2773,N_245,N_1790);
nand U2774 (N_2774,N_40,N_1732);
and U2775 (N_2775,N_871,N_399);
xnor U2776 (N_2776,N_1451,N_542);
nand U2777 (N_2777,N_561,N_1917);
nor U2778 (N_2778,N_1961,N_723);
and U2779 (N_2779,N_1596,N_209);
or U2780 (N_2780,N_763,N_20);
and U2781 (N_2781,N_1464,N_1539);
and U2782 (N_2782,N_1315,N_1200);
nor U2783 (N_2783,N_927,N_170);
nand U2784 (N_2784,N_579,N_15);
or U2785 (N_2785,N_808,N_1411);
xnor U2786 (N_2786,N_822,N_434);
nor U2787 (N_2787,N_1219,N_1880);
or U2788 (N_2788,N_943,N_725);
xnor U2789 (N_2789,N_212,N_846);
nor U2790 (N_2790,N_1656,N_199);
and U2791 (N_2791,N_768,N_1497);
or U2792 (N_2792,N_180,N_109);
nor U2793 (N_2793,N_1618,N_1035);
nor U2794 (N_2794,N_1106,N_1761);
nand U2795 (N_2795,N_77,N_171);
and U2796 (N_2796,N_1974,N_1888);
xor U2797 (N_2797,N_1503,N_1055);
and U2798 (N_2798,N_826,N_378);
or U2799 (N_2799,N_1368,N_1350);
and U2800 (N_2800,N_745,N_762);
xnor U2801 (N_2801,N_1197,N_137);
nor U2802 (N_2802,N_1149,N_1762);
nand U2803 (N_2803,N_96,N_1224);
nand U2804 (N_2804,N_1076,N_1649);
xor U2805 (N_2805,N_582,N_879);
nand U2806 (N_2806,N_135,N_533);
nand U2807 (N_2807,N_1582,N_242);
nand U2808 (N_2808,N_969,N_1302);
or U2809 (N_2809,N_1276,N_196);
nor U2810 (N_2810,N_821,N_896);
nand U2811 (N_2811,N_1931,N_243);
and U2812 (N_2812,N_336,N_509);
xor U2813 (N_2813,N_537,N_1531);
and U2814 (N_2814,N_622,N_752);
nand U2815 (N_2815,N_138,N_1151);
xnor U2816 (N_2816,N_1408,N_162);
nor U2817 (N_2817,N_1384,N_1500);
nor U2818 (N_2818,N_888,N_1636);
nor U2819 (N_2819,N_401,N_1365);
and U2820 (N_2820,N_1455,N_1223);
xor U2821 (N_2821,N_909,N_97);
or U2822 (N_2822,N_1477,N_184);
or U2823 (N_2823,N_985,N_452);
xnor U2824 (N_2824,N_534,N_1654);
nand U2825 (N_2825,N_1468,N_61);
xnor U2826 (N_2826,N_615,N_30);
xnor U2827 (N_2827,N_992,N_1842);
xnor U2828 (N_2828,N_848,N_425);
nand U2829 (N_2829,N_1064,N_373);
or U2830 (N_2830,N_966,N_873);
nand U2831 (N_2831,N_1733,N_621);
nor U2832 (N_2832,N_1809,N_1340);
nor U2833 (N_2833,N_284,N_145);
nor U2834 (N_2834,N_1673,N_1362);
or U2835 (N_2835,N_1227,N_563);
nand U2836 (N_2836,N_443,N_897);
nor U2837 (N_2837,N_150,N_69);
nor U2838 (N_2838,N_1628,N_1826);
xor U2839 (N_2839,N_1816,N_913);
nor U2840 (N_2840,N_1039,N_1125);
nand U2841 (N_2841,N_1291,N_493);
nor U2842 (N_2842,N_1589,N_1292);
xnor U2843 (N_2843,N_1591,N_1601);
xor U2844 (N_2844,N_942,N_70);
and U2845 (N_2845,N_876,N_466);
nor U2846 (N_2846,N_117,N_303);
nor U2847 (N_2847,N_1921,N_306);
nor U2848 (N_2848,N_721,N_1755);
xor U2849 (N_2849,N_692,N_282);
and U2850 (N_2850,N_255,N_1017);
nand U2851 (N_2851,N_386,N_1033);
nor U2852 (N_2852,N_964,N_1815);
nand U2853 (N_2853,N_1972,N_275);
and U2854 (N_2854,N_774,N_57);
nor U2855 (N_2855,N_149,N_1496);
nand U2856 (N_2856,N_1381,N_1491);
nor U2857 (N_2857,N_1335,N_515);
nor U2858 (N_2858,N_354,N_1810);
nand U2859 (N_2859,N_1637,N_1467);
nor U2860 (N_2860,N_1980,N_724);
or U2861 (N_2861,N_1447,N_1070);
nand U2862 (N_2862,N_1466,N_1587);
or U2863 (N_2863,N_1417,N_1266);
or U2864 (N_2864,N_996,N_1854);
and U2865 (N_2865,N_166,N_339);
nor U2866 (N_2866,N_1635,N_1712);
or U2867 (N_2867,N_852,N_612);
xor U2868 (N_2868,N_1410,N_1674);
nand U2869 (N_2869,N_312,N_1952);
xor U2870 (N_2870,N_627,N_1887);
or U2871 (N_2871,N_668,N_682);
nor U2872 (N_2872,N_671,N_649);
xnor U2873 (N_2873,N_311,N_105);
nor U2874 (N_2874,N_86,N_317);
nor U2875 (N_2875,N_1034,N_272);
nor U2876 (N_2876,N_463,N_1169);
xnor U2877 (N_2877,N_1744,N_508);
and U2878 (N_2878,N_1353,N_486);
and U2879 (N_2879,N_1306,N_973);
xnor U2880 (N_2880,N_1480,N_523);
xor U2881 (N_2881,N_1836,N_201);
and U2882 (N_2882,N_139,N_1990);
xor U2883 (N_2883,N_765,N_1736);
nand U2884 (N_2884,N_17,N_192);
nand U2885 (N_2885,N_1090,N_874);
and U2886 (N_2886,N_59,N_12);
and U2887 (N_2887,N_1380,N_906);
and U2888 (N_2888,N_1349,N_819);
nor U2889 (N_2889,N_1061,N_997);
xnor U2890 (N_2890,N_1299,N_1847);
and U2891 (N_2891,N_810,N_1559);
and U2892 (N_2892,N_708,N_910);
nand U2893 (N_2893,N_1545,N_814);
or U2894 (N_2894,N_431,N_377);
and U2895 (N_2895,N_1442,N_74);
and U2896 (N_2896,N_1265,N_1928);
xnor U2897 (N_2897,N_520,N_1892);
and U2898 (N_2898,N_999,N_761);
and U2899 (N_2899,N_1221,N_887);
or U2900 (N_2900,N_1479,N_991);
and U2901 (N_2901,N_422,N_274);
nand U2902 (N_2902,N_522,N_1420);
and U2903 (N_2903,N_657,N_587);
and U2904 (N_2904,N_954,N_261);
nor U2905 (N_2905,N_345,N_93);
nor U2906 (N_2906,N_1433,N_490);
or U2907 (N_2907,N_844,N_22);
nand U2908 (N_2908,N_1991,N_356);
and U2909 (N_2909,N_203,N_497);
and U2910 (N_2910,N_1865,N_842);
and U2911 (N_2911,N_1789,N_454);
or U2912 (N_2912,N_42,N_1143);
nor U2913 (N_2913,N_65,N_1423);
nand U2914 (N_2914,N_374,N_556);
nand U2915 (N_2915,N_168,N_147);
and U2916 (N_2916,N_144,N_1329);
or U2917 (N_2917,N_517,N_767);
xor U2918 (N_2918,N_553,N_833);
and U2919 (N_2919,N_1915,N_1099);
and U2920 (N_2920,N_505,N_476);
nand U2921 (N_2921,N_550,N_978);
and U2922 (N_2922,N_880,N_75);
or U2923 (N_2923,N_140,N_1694);
nand U2924 (N_2924,N_685,N_566);
and U2925 (N_2925,N_94,N_1568);
xnor U2926 (N_2926,N_461,N_1489);
and U2927 (N_2927,N_1870,N_1449);
or U2928 (N_2928,N_1237,N_1770);
nand U2929 (N_2929,N_182,N_857);
or U2930 (N_2930,N_239,N_706);
nand U2931 (N_2931,N_646,N_412);
xor U2932 (N_2932,N_1597,N_1528);
xor U2933 (N_2933,N_667,N_836);
nor U2934 (N_2934,N_1624,N_1327);
xnor U2935 (N_2935,N_1777,N_1753);
xor U2936 (N_2936,N_700,N_1890);
nand U2937 (N_2937,N_1938,N_578);
nor U2938 (N_2938,N_222,N_1402);
or U2939 (N_2939,N_1540,N_496);
nand U2940 (N_2940,N_1575,N_352);
nand U2941 (N_2941,N_1133,N_572);
nor U2942 (N_2942,N_1822,N_696);
and U2943 (N_2943,N_1585,N_278);
xor U2944 (N_2944,N_1818,N_1228);
nor U2945 (N_2945,N_1320,N_332);
xor U2946 (N_2946,N_1347,N_99);
or U2947 (N_2947,N_1821,N_130);
xor U2948 (N_2948,N_1354,N_1012);
or U2949 (N_2949,N_895,N_698);
and U2950 (N_2950,N_1041,N_478);
or U2951 (N_2951,N_310,N_1419);
and U2952 (N_2952,N_43,N_1157);
nor U2953 (N_2953,N_1705,N_417);
and U2954 (N_2954,N_1519,N_1786);
and U2955 (N_2955,N_1719,N_705);
and U2956 (N_2956,N_1001,N_1806);
nand U2957 (N_2957,N_932,N_624);
and U2958 (N_2958,N_23,N_940);
xor U2959 (N_2959,N_376,N_1983);
or U2960 (N_2960,N_1904,N_1164);
xnor U2961 (N_2961,N_1897,N_1397);
or U2962 (N_2962,N_719,N_116);
nand U2963 (N_2963,N_993,N_1259);
nand U2964 (N_2964,N_898,N_911);
xor U2965 (N_2965,N_1922,N_44);
xor U2966 (N_2966,N_1754,N_878);
nor U2967 (N_2967,N_298,N_549);
nor U2968 (N_2968,N_1910,N_1341);
nand U2969 (N_2969,N_926,N_402);
or U2970 (N_2970,N_1153,N_1031);
and U2971 (N_2971,N_124,N_1885);
nand U2972 (N_2972,N_223,N_185);
nand U2973 (N_2973,N_1615,N_1056);
nor U2974 (N_2974,N_67,N_1044);
xnor U2975 (N_2975,N_1558,N_37);
nor U2976 (N_2976,N_1560,N_540);
xor U2977 (N_2977,N_1370,N_1949);
nor U2978 (N_2978,N_862,N_189);
xor U2979 (N_2979,N_1584,N_1994);
nor U2980 (N_2980,N_1046,N_642);
and U2981 (N_2981,N_979,N_1089);
nor U2982 (N_2982,N_1759,N_163);
and U2983 (N_2983,N_1304,N_395);
and U2984 (N_2984,N_1891,N_847);
or U2985 (N_2985,N_1383,N_477);
or U2986 (N_2986,N_1652,N_55);
xor U2987 (N_2987,N_113,N_776);
xor U2988 (N_2988,N_257,N_78);
nand U2989 (N_2989,N_1543,N_1092);
nor U2990 (N_2990,N_134,N_912);
nand U2991 (N_2991,N_931,N_315);
or U2992 (N_2992,N_867,N_680);
xnor U2993 (N_2993,N_1695,N_1752);
xnor U2994 (N_2994,N_1294,N_475);
xnor U2995 (N_2995,N_1580,N_1969);
nor U2996 (N_2996,N_1435,N_818);
nor U2997 (N_2997,N_1838,N_1009);
nand U2998 (N_2998,N_1130,N_369);
nand U2999 (N_2999,N_1570,N_479);
or U3000 (N_3000,N_973,N_1127);
nor U3001 (N_3001,N_381,N_1418);
nor U3002 (N_3002,N_1473,N_1924);
xor U3003 (N_3003,N_687,N_58);
xor U3004 (N_3004,N_739,N_1664);
nand U3005 (N_3005,N_588,N_861);
or U3006 (N_3006,N_7,N_1551);
and U3007 (N_3007,N_198,N_376);
nand U3008 (N_3008,N_1104,N_1892);
or U3009 (N_3009,N_1322,N_1653);
and U3010 (N_3010,N_516,N_1072);
nand U3011 (N_3011,N_1215,N_1504);
or U3012 (N_3012,N_1218,N_357);
or U3013 (N_3013,N_1141,N_501);
or U3014 (N_3014,N_1476,N_1869);
xor U3015 (N_3015,N_1054,N_1749);
and U3016 (N_3016,N_1357,N_1113);
xor U3017 (N_3017,N_958,N_1772);
nor U3018 (N_3018,N_1051,N_1457);
or U3019 (N_3019,N_1219,N_1570);
or U3020 (N_3020,N_871,N_1461);
nor U3021 (N_3021,N_699,N_721);
xor U3022 (N_3022,N_1380,N_815);
or U3023 (N_3023,N_13,N_1341);
and U3024 (N_3024,N_563,N_1992);
nor U3025 (N_3025,N_1773,N_1104);
nand U3026 (N_3026,N_317,N_1690);
xor U3027 (N_3027,N_1693,N_299);
nand U3028 (N_3028,N_654,N_1840);
and U3029 (N_3029,N_1149,N_1274);
nor U3030 (N_3030,N_205,N_1045);
xnor U3031 (N_3031,N_1958,N_172);
and U3032 (N_3032,N_336,N_1028);
nor U3033 (N_3033,N_1709,N_897);
nand U3034 (N_3034,N_627,N_880);
and U3035 (N_3035,N_1119,N_1270);
nand U3036 (N_3036,N_1875,N_778);
and U3037 (N_3037,N_121,N_205);
and U3038 (N_3038,N_1361,N_1124);
nor U3039 (N_3039,N_639,N_1616);
xor U3040 (N_3040,N_684,N_1643);
nand U3041 (N_3041,N_1275,N_660);
or U3042 (N_3042,N_982,N_1860);
nand U3043 (N_3043,N_936,N_92);
or U3044 (N_3044,N_1789,N_1861);
or U3045 (N_3045,N_827,N_1032);
xnor U3046 (N_3046,N_395,N_1237);
xnor U3047 (N_3047,N_1294,N_1916);
xor U3048 (N_3048,N_261,N_1425);
nor U3049 (N_3049,N_488,N_1852);
nand U3050 (N_3050,N_1103,N_4);
and U3051 (N_3051,N_1150,N_933);
and U3052 (N_3052,N_639,N_1243);
and U3053 (N_3053,N_1498,N_1336);
or U3054 (N_3054,N_498,N_1599);
nand U3055 (N_3055,N_1297,N_1192);
or U3056 (N_3056,N_1996,N_982);
and U3057 (N_3057,N_606,N_1288);
nand U3058 (N_3058,N_1050,N_1108);
or U3059 (N_3059,N_704,N_99);
and U3060 (N_3060,N_1202,N_764);
nor U3061 (N_3061,N_1912,N_400);
xnor U3062 (N_3062,N_1667,N_1900);
xnor U3063 (N_3063,N_1343,N_386);
and U3064 (N_3064,N_1648,N_1459);
nand U3065 (N_3065,N_1335,N_314);
nor U3066 (N_3066,N_1874,N_1353);
nor U3067 (N_3067,N_1548,N_486);
xor U3068 (N_3068,N_796,N_902);
nand U3069 (N_3069,N_552,N_1743);
xor U3070 (N_3070,N_724,N_474);
nor U3071 (N_3071,N_482,N_1468);
xnor U3072 (N_3072,N_1091,N_1369);
and U3073 (N_3073,N_559,N_298);
xor U3074 (N_3074,N_1928,N_37);
or U3075 (N_3075,N_25,N_480);
nor U3076 (N_3076,N_1343,N_450);
nand U3077 (N_3077,N_821,N_1362);
nor U3078 (N_3078,N_1617,N_1672);
nand U3079 (N_3079,N_1175,N_174);
xnor U3080 (N_3080,N_1773,N_1942);
nand U3081 (N_3081,N_572,N_1534);
nor U3082 (N_3082,N_481,N_1344);
nor U3083 (N_3083,N_683,N_1856);
nor U3084 (N_3084,N_443,N_257);
nor U3085 (N_3085,N_72,N_1954);
xor U3086 (N_3086,N_10,N_1578);
xnor U3087 (N_3087,N_1086,N_309);
nor U3088 (N_3088,N_1638,N_1039);
or U3089 (N_3089,N_1732,N_199);
and U3090 (N_3090,N_808,N_1785);
or U3091 (N_3091,N_1125,N_1947);
xnor U3092 (N_3092,N_1737,N_1182);
nand U3093 (N_3093,N_1544,N_339);
or U3094 (N_3094,N_414,N_1200);
nor U3095 (N_3095,N_1010,N_1960);
and U3096 (N_3096,N_984,N_689);
or U3097 (N_3097,N_1841,N_1426);
and U3098 (N_3098,N_951,N_1105);
nand U3099 (N_3099,N_1816,N_1454);
nand U3100 (N_3100,N_1856,N_1221);
nor U3101 (N_3101,N_1220,N_95);
and U3102 (N_3102,N_1235,N_910);
or U3103 (N_3103,N_1353,N_1270);
or U3104 (N_3104,N_876,N_1685);
nand U3105 (N_3105,N_1606,N_1438);
nand U3106 (N_3106,N_1703,N_1626);
or U3107 (N_3107,N_1465,N_1107);
or U3108 (N_3108,N_1737,N_1922);
nand U3109 (N_3109,N_1009,N_575);
nor U3110 (N_3110,N_557,N_1101);
or U3111 (N_3111,N_237,N_543);
nor U3112 (N_3112,N_1830,N_457);
and U3113 (N_3113,N_656,N_1309);
or U3114 (N_3114,N_1835,N_1510);
xor U3115 (N_3115,N_1963,N_1681);
and U3116 (N_3116,N_1634,N_1605);
nand U3117 (N_3117,N_1835,N_1958);
and U3118 (N_3118,N_1077,N_1052);
and U3119 (N_3119,N_846,N_1167);
and U3120 (N_3120,N_1120,N_1683);
xor U3121 (N_3121,N_1564,N_995);
nor U3122 (N_3122,N_833,N_857);
and U3123 (N_3123,N_1632,N_179);
xor U3124 (N_3124,N_767,N_1203);
nand U3125 (N_3125,N_1613,N_51);
or U3126 (N_3126,N_1555,N_1995);
and U3127 (N_3127,N_1009,N_1549);
nor U3128 (N_3128,N_1575,N_1685);
or U3129 (N_3129,N_1853,N_1082);
or U3130 (N_3130,N_152,N_617);
nor U3131 (N_3131,N_1128,N_1922);
or U3132 (N_3132,N_790,N_343);
or U3133 (N_3133,N_18,N_638);
xor U3134 (N_3134,N_1870,N_556);
xor U3135 (N_3135,N_1671,N_26);
nor U3136 (N_3136,N_1392,N_1298);
nand U3137 (N_3137,N_1198,N_123);
xor U3138 (N_3138,N_1444,N_69);
and U3139 (N_3139,N_584,N_1444);
nand U3140 (N_3140,N_1383,N_1070);
nand U3141 (N_3141,N_1732,N_1686);
xnor U3142 (N_3142,N_1873,N_1665);
nor U3143 (N_3143,N_873,N_1851);
and U3144 (N_3144,N_1662,N_634);
xor U3145 (N_3145,N_513,N_182);
nor U3146 (N_3146,N_847,N_1);
nand U3147 (N_3147,N_1431,N_1959);
or U3148 (N_3148,N_52,N_872);
and U3149 (N_3149,N_444,N_1469);
or U3150 (N_3150,N_1751,N_745);
xnor U3151 (N_3151,N_1550,N_904);
nor U3152 (N_3152,N_1616,N_1093);
nor U3153 (N_3153,N_1981,N_604);
or U3154 (N_3154,N_1802,N_917);
and U3155 (N_3155,N_1885,N_444);
and U3156 (N_3156,N_951,N_1024);
xor U3157 (N_3157,N_1082,N_489);
nor U3158 (N_3158,N_1476,N_84);
or U3159 (N_3159,N_75,N_139);
or U3160 (N_3160,N_1155,N_1754);
and U3161 (N_3161,N_268,N_249);
xor U3162 (N_3162,N_1325,N_1192);
or U3163 (N_3163,N_1126,N_1266);
or U3164 (N_3164,N_989,N_496);
or U3165 (N_3165,N_302,N_958);
xnor U3166 (N_3166,N_1265,N_226);
or U3167 (N_3167,N_261,N_696);
xor U3168 (N_3168,N_118,N_1241);
nor U3169 (N_3169,N_142,N_1203);
xor U3170 (N_3170,N_1920,N_54);
nor U3171 (N_3171,N_811,N_136);
or U3172 (N_3172,N_290,N_907);
and U3173 (N_3173,N_219,N_1055);
nand U3174 (N_3174,N_727,N_1886);
and U3175 (N_3175,N_1685,N_1275);
xor U3176 (N_3176,N_485,N_336);
or U3177 (N_3177,N_1804,N_991);
nor U3178 (N_3178,N_719,N_1899);
and U3179 (N_3179,N_1568,N_312);
nand U3180 (N_3180,N_1852,N_1600);
nor U3181 (N_3181,N_1088,N_1343);
or U3182 (N_3182,N_723,N_331);
or U3183 (N_3183,N_1274,N_499);
xnor U3184 (N_3184,N_917,N_421);
xnor U3185 (N_3185,N_1139,N_753);
and U3186 (N_3186,N_1634,N_387);
nor U3187 (N_3187,N_403,N_145);
xnor U3188 (N_3188,N_615,N_1274);
nand U3189 (N_3189,N_1007,N_1817);
xor U3190 (N_3190,N_1203,N_1931);
xor U3191 (N_3191,N_353,N_1985);
nand U3192 (N_3192,N_563,N_476);
nor U3193 (N_3193,N_152,N_562);
nand U3194 (N_3194,N_1641,N_1862);
nand U3195 (N_3195,N_174,N_94);
or U3196 (N_3196,N_185,N_443);
and U3197 (N_3197,N_1474,N_175);
or U3198 (N_3198,N_694,N_1899);
nand U3199 (N_3199,N_375,N_416);
and U3200 (N_3200,N_1572,N_1165);
nor U3201 (N_3201,N_1342,N_1108);
and U3202 (N_3202,N_1851,N_164);
xnor U3203 (N_3203,N_1705,N_188);
and U3204 (N_3204,N_472,N_1426);
nand U3205 (N_3205,N_142,N_738);
nand U3206 (N_3206,N_1958,N_231);
or U3207 (N_3207,N_242,N_1850);
nand U3208 (N_3208,N_1233,N_1170);
nand U3209 (N_3209,N_1115,N_632);
and U3210 (N_3210,N_1996,N_1782);
nor U3211 (N_3211,N_95,N_400);
nor U3212 (N_3212,N_1526,N_1899);
and U3213 (N_3213,N_1083,N_1692);
and U3214 (N_3214,N_1879,N_923);
or U3215 (N_3215,N_251,N_692);
and U3216 (N_3216,N_1040,N_8);
nand U3217 (N_3217,N_193,N_616);
xor U3218 (N_3218,N_945,N_228);
nand U3219 (N_3219,N_175,N_416);
or U3220 (N_3220,N_627,N_689);
nand U3221 (N_3221,N_581,N_1423);
or U3222 (N_3222,N_1597,N_704);
xnor U3223 (N_3223,N_1121,N_260);
nand U3224 (N_3224,N_1467,N_1286);
and U3225 (N_3225,N_61,N_827);
or U3226 (N_3226,N_1261,N_977);
or U3227 (N_3227,N_152,N_711);
nand U3228 (N_3228,N_1583,N_281);
xor U3229 (N_3229,N_1686,N_1210);
or U3230 (N_3230,N_1246,N_683);
and U3231 (N_3231,N_1106,N_1927);
xor U3232 (N_3232,N_1930,N_1603);
and U3233 (N_3233,N_1682,N_1192);
nand U3234 (N_3234,N_197,N_1514);
or U3235 (N_3235,N_785,N_464);
or U3236 (N_3236,N_1339,N_643);
nor U3237 (N_3237,N_341,N_1102);
or U3238 (N_3238,N_1719,N_1341);
or U3239 (N_3239,N_1571,N_25);
and U3240 (N_3240,N_1917,N_1292);
nand U3241 (N_3241,N_118,N_289);
nand U3242 (N_3242,N_242,N_267);
nor U3243 (N_3243,N_1036,N_1809);
xnor U3244 (N_3244,N_743,N_1507);
or U3245 (N_3245,N_112,N_401);
or U3246 (N_3246,N_1597,N_1278);
nor U3247 (N_3247,N_1072,N_1617);
and U3248 (N_3248,N_578,N_504);
or U3249 (N_3249,N_869,N_254);
and U3250 (N_3250,N_1919,N_598);
nand U3251 (N_3251,N_1616,N_1390);
nor U3252 (N_3252,N_1185,N_1347);
or U3253 (N_3253,N_498,N_1539);
nand U3254 (N_3254,N_1532,N_1753);
and U3255 (N_3255,N_1925,N_1517);
xnor U3256 (N_3256,N_1406,N_1955);
nor U3257 (N_3257,N_1438,N_1526);
nand U3258 (N_3258,N_168,N_1213);
nor U3259 (N_3259,N_504,N_1676);
xnor U3260 (N_3260,N_1391,N_1190);
and U3261 (N_3261,N_197,N_1153);
or U3262 (N_3262,N_980,N_1723);
nand U3263 (N_3263,N_1043,N_1302);
nand U3264 (N_3264,N_524,N_1333);
or U3265 (N_3265,N_553,N_628);
nand U3266 (N_3266,N_714,N_1502);
nor U3267 (N_3267,N_1540,N_534);
or U3268 (N_3268,N_1337,N_393);
or U3269 (N_3269,N_1955,N_808);
nor U3270 (N_3270,N_1525,N_1218);
and U3271 (N_3271,N_1958,N_44);
and U3272 (N_3272,N_1558,N_1479);
and U3273 (N_3273,N_1987,N_1634);
xnor U3274 (N_3274,N_75,N_1926);
nor U3275 (N_3275,N_1464,N_1181);
or U3276 (N_3276,N_1195,N_539);
nand U3277 (N_3277,N_1283,N_845);
xor U3278 (N_3278,N_1377,N_1162);
nand U3279 (N_3279,N_1004,N_200);
or U3280 (N_3280,N_469,N_1113);
xor U3281 (N_3281,N_813,N_294);
xnor U3282 (N_3282,N_1327,N_1778);
or U3283 (N_3283,N_559,N_1434);
nor U3284 (N_3284,N_569,N_1933);
xnor U3285 (N_3285,N_97,N_1105);
or U3286 (N_3286,N_893,N_1264);
nand U3287 (N_3287,N_1251,N_986);
xor U3288 (N_3288,N_1503,N_395);
xnor U3289 (N_3289,N_626,N_604);
and U3290 (N_3290,N_290,N_280);
nand U3291 (N_3291,N_460,N_1397);
nand U3292 (N_3292,N_818,N_225);
xnor U3293 (N_3293,N_891,N_1842);
and U3294 (N_3294,N_1585,N_1579);
nand U3295 (N_3295,N_831,N_1747);
and U3296 (N_3296,N_1608,N_134);
nand U3297 (N_3297,N_990,N_1948);
nor U3298 (N_3298,N_966,N_911);
and U3299 (N_3299,N_1927,N_1779);
nand U3300 (N_3300,N_1797,N_852);
or U3301 (N_3301,N_1352,N_1852);
and U3302 (N_3302,N_1713,N_867);
nor U3303 (N_3303,N_469,N_1151);
nand U3304 (N_3304,N_889,N_673);
nand U3305 (N_3305,N_1164,N_126);
xor U3306 (N_3306,N_885,N_64);
or U3307 (N_3307,N_1961,N_286);
nor U3308 (N_3308,N_1271,N_1144);
nand U3309 (N_3309,N_471,N_962);
or U3310 (N_3310,N_58,N_47);
and U3311 (N_3311,N_1303,N_787);
or U3312 (N_3312,N_736,N_470);
xnor U3313 (N_3313,N_1183,N_1957);
and U3314 (N_3314,N_1202,N_1789);
and U3315 (N_3315,N_1038,N_1946);
nand U3316 (N_3316,N_459,N_376);
nand U3317 (N_3317,N_910,N_768);
nor U3318 (N_3318,N_403,N_1377);
nor U3319 (N_3319,N_1128,N_317);
and U3320 (N_3320,N_281,N_965);
nand U3321 (N_3321,N_954,N_9);
xor U3322 (N_3322,N_1146,N_747);
xor U3323 (N_3323,N_1744,N_234);
nand U3324 (N_3324,N_1781,N_810);
and U3325 (N_3325,N_1453,N_563);
and U3326 (N_3326,N_1561,N_96);
nand U3327 (N_3327,N_283,N_651);
nor U3328 (N_3328,N_934,N_142);
or U3329 (N_3329,N_519,N_1045);
nand U3330 (N_3330,N_1561,N_1705);
xor U3331 (N_3331,N_493,N_1048);
or U3332 (N_3332,N_832,N_1562);
nand U3333 (N_3333,N_1408,N_501);
or U3334 (N_3334,N_746,N_1270);
nand U3335 (N_3335,N_1787,N_100);
nor U3336 (N_3336,N_490,N_1373);
and U3337 (N_3337,N_1555,N_741);
xnor U3338 (N_3338,N_511,N_1938);
and U3339 (N_3339,N_248,N_1373);
nand U3340 (N_3340,N_1383,N_210);
and U3341 (N_3341,N_349,N_1163);
or U3342 (N_3342,N_369,N_1010);
and U3343 (N_3343,N_1953,N_1724);
xnor U3344 (N_3344,N_1685,N_1417);
nor U3345 (N_3345,N_1291,N_875);
nor U3346 (N_3346,N_1082,N_348);
or U3347 (N_3347,N_314,N_1578);
xnor U3348 (N_3348,N_1292,N_501);
nand U3349 (N_3349,N_1198,N_494);
nand U3350 (N_3350,N_111,N_1337);
xor U3351 (N_3351,N_1322,N_1400);
xnor U3352 (N_3352,N_55,N_1189);
xor U3353 (N_3353,N_431,N_781);
or U3354 (N_3354,N_388,N_1696);
nor U3355 (N_3355,N_1707,N_5);
or U3356 (N_3356,N_775,N_1084);
nand U3357 (N_3357,N_1895,N_1236);
and U3358 (N_3358,N_1540,N_1294);
nor U3359 (N_3359,N_1424,N_277);
nand U3360 (N_3360,N_889,N_1347);
and U3361 (N_3361,N_420,N_1149);
and U3362 (N_3362,N_512,N_1211);
or U3363 (N_3363,N_729,N_1889);
nor U3364 (N_3364,N_1566,N_879);
or U3365 (N_3365,N_294,N_677);
xnor U3366 (N_3366,N_1909,N_232);
nand U3367 (N_3367,N_201,N_1644);
and U3368 (N_3368,N_1646,N_1184);
nand U3369 (N_3369,N_503,N_1595);
or U3370 (N_3370,N_1519,N_1335);
nor U3371 (N_3371,N_1995,N_262);
or U3372 (N_3372,N_1996,N_1163);
or U3373 (N_3373,N_1207,N_1209);
and U3374 (N_3374,N_353,N_857);
xor U3375 (N_3375,N_1902,N_369);
nand U3376 (N_3376,N_393,N_776);
xnor U3377 (N_3377,N_921,N_1912);
nor U3378 (N_3378,N_1400,N_689);
nand U3379 (N_3379,N_359,N_1304);
xnor U3380 (N_3380,N_25,N_956);
nand U3381 (N_3381,N_1592,N_695);
nor U3382 (N_3382,N_888,N_897);
nand U3383 (N_3383,N_1565,N_822);
and U3384 (N_3384,N_737,N_1230);
nor U3385 (N_3385,N_616,N_1595);
nand U3386 (N_3386,N_367,N_966);
xor U3387 (N_3387,N_941,N_381);
nand U3388 (N_3388,N_548,N_929);
nor U3389 (N_3389,N_1590,N_503);
or U3390 (N_3390,N_1227,N_533);
nand U3391 (N_3391,N_893,N_1437);
nor U3392 (N_3392,N_1918,N_585);
xnor U3393 (N_3393,N_1639,N_1130);
or U3394 (N_3394,N_1842,N_1938);
nand U3395 (N_3395,N_1143,N_911);
or U3396 (N_3396,N_1226,N_305);
nor U3397 (N_3397,N_1186,N_905);
nand U3398 (N_3398,N_434,N_189);
and U3399 (N_3399,N_480,N_1623);
or U3400 (N_3400,N_289,N_1381);
nand U3401 (N_3401,N_234,N_1339);
or U3402 (N_3402,N_1096,N_1352);
xor U3403 (N_3403,N_41,N_45);
or U3404 (N_3404,N_1184,N_1117);
and U3405 (N_3405,N_608,N_1200);
or U3406 (N_3406,N_1438,N_1261);
xor U3407 (N_3407,N_189,N_1899);
xnor U3408 (N_3408,N_1208,N_277);
xnor U3409 (N_3409,N_875,N_1912);
and U3410 (N_3410,N_1331,N_1696);
xnor U3411 (N_3411,N_1240,N_1612);
nand U3412 (N_3412,N_17,N_250);
nor U3413 (N_3413,N_1286,N_1983);
and U3414 (N_3414,N_380,N_1984);
xor U3415 (N_3415,N_1239,N_482);
nand U3416 (N_3416,N_1429,N_943);
xor U3417 (N_3417,N_1915,N_981);
and U3418 (N_3418,N_204,N_1486);
and U3419 (N_3419,N_918,N_644);
and U3420 (N_3420,N_878,N_1276);
and U3421 (N_3421,N_286,N_1363);
or U3422 (N_3422,N_1269,N_1529);
and U3423 (N_3423,N_552,N_790);
nor U3424 (N_3424,N_1757,N_506);
nor U3425 (N_3425,N_535,N_1980);
or U3426 (N_3426,N_585,N_1551);
or U3427 (N_3427,N_332,N_1288);
nand U3428 (N_3428,N_1588,N_1467);
nand U3429 (N_3429,N_971,N_1942);
or U3430 (N_3430,N_640,N_665);
or U3431 (N_3431,N_1132,N_393);
or U3432 (N_3432,N_488,N_1177);
or U3433 (N_3433,N_1309,N_1680);
nand U3434 (N_3434,N_620,N_37);
nor U3435 (N_3435,N_1862,N_1233);
nand U3436 (N_3436,N_262,N_1830);
nor U3437 (N_3437,N_526,N_861);
nor U3438 (N_3438,N_639,N_16);
nand U3439 (N_3439,N_1503,N_1112);
nor U3440 (N_3440,N_1258,N_1153);
and U3441 (N_3441,N_1444,N_826);
or U3442 (N_3442,N_1340,N_1741);
and U3443 (N_3443,N_1439,N_397);
or U3444 (N_3444,N_1142,N_1328);
or U3445 (N_3445,N_7,N_297);
and U3446 (N_3446,N_1528,N_289);
or U3447 (N_3447,N_112,N_1284);
and U3448 (N_3448,N_1782,N_868);
xor U3449 (N_3449,N_465,N_1562);
nor U3450 (N_3450,N_1972,N_858);
or U3451 (N_3451,N_211,N_1571);
or U3452 (N_3452,N_1641,N_488);
xor U3453 (N_3453,N_61,N_948);
xor U3454 (N_3454,N_1690,N_613);
nor U3455 (N_3455,N_1413,N_761);
and U3456 (N_3456,N_1264,N_830);
xnor U3457 (N_3457,N_1480,N_341);
nand U3458 (N_3458,N_669,N_1522);
nand U3459 (N_3459,N_220,N_547);
nand U3460 (N_3460,N_390,N_500);
and U3461 (N_3461,N_517,N_1937);
nand U3462 (N_3462,N_1750,N_1533);
or U3463 (N_3463,N_433,N_1281);
or U3464 (N_3464,N_1847,N_1448);
nand U3465 (N_3465,N_41,N_195);
nand U3466 (N_3466,N_1959,N_1551);
nand U3467 (N_3467,N_1906,N_796);
and U3468 (N_3468,N_155,N_1822);
nor U3469 (N_3469,N_227,N_691);
nand U3470 (N_3470,N_726,N_493);
xnor U3471 (N_3471,N_833,N_1287);
xnor U3472 (N_3472,N_825,N_876);
nand U3473 (N_3473,N_114,N_143);
nor U3474 (N_3474,N_1719,N_326);
or U3475 (N_3475,N_97,N_1890);
nor U3476 (N_3476,N_379,N_946);
or U3477 (N_3477,N_1997,N_852);
and U3478 (N_3478,N_936,N_1661);
or U3479 (N_3479,N_367,N_883);
and U3480 (N_3480,N_228,N_1017);
or U3481 (N_3481,N_569,N_56);
nand U3482 (N_3482,N_1002,N_1560);
nor U3483 (N_3483,N_1597,N_497);
or U3484 (N_3484,N_1389,N_239);
nand U3485 (N_3485,N_151,N_1329);
nand U3486 (N_3486,N_673,N_592);
and U3487 (N_3487,N_1129,N_324);
and U3488 (N_3488,N_836,N_630);
or U3489 (N_3489,N_905,N_34);
xnor U3490 (N_3490,N_486,N_615);
nor U3491 (N_3491,N_1671,N_73);
nand U3492 (N_3492,N_1574,N_1304);
nand U3493 (N_3493,N_203,N_775);
and U3494 (N_3494,N_863,N_633);
nand U3495 (N_3495,N_653,N_960);
or U3496 (N_3496,N_1007,N_1370);
or U3497 (N_3497,N_720,N_622);
nand U3498 (N_3498,N_126,N_591);
and U3499 (N_3499,N_91,N_370);
nor U3500 (N_3500,N_1622,N_195);
and U3501 (N_3501,N_1979,N_1742);
nor U3502 (N_3502,N_1165,N_89);
nor U3503 (N_3503,N_499,N_916);
nor U3504 (N_3504,N_43,N_270);
nand U3505 (N_3505,N_245,N_1644);
nand U3506 (N_3506,N_0,N_568);
or U3507 (N_3507,N_682,N_756);
nor U3508 (N_3508,N_773,N_1913);
xor U3509 (N_3509,N_1004,N_925);
xor U3510 (N_3510,N_686,N_280);
xor U3511 (N_3511,N_116,N_817);
or U3512 (N_3512,N_1942,N_1730);
nor U3513 (N_3513,N_1438,N_1710);
or U3514 (N_3514,N_1562,N_1875);
nor U3515 (N_3515,N_988,N_1444);
xnor U3516 (N_3516,N_1990,N_1558);
nand U3517 (N_3517,N_481,N_256);
or U3518 (N_3518,N_907,N_1531);
and U3519 (N_3519,N_1216,N_913);
nand U3520 (N_3520,N_926,N_321);
nand U3521 (N_3521,N_1995,N_1375);
xnor U3522 (N_3522,N_205,N_197);
and U3523 (N_3523,N_1683,N_1890);
nor U3524 (N_3524,N_1631,N_879);
nor U3525 (N_3525,N_719,N_127);
nor U3526 (N_3526,N_535,N_1851);
nor U3527 (N_3527,N_74,N_849);
or U3528 (N_3528,N_504,N_1327);
nor U3529 (N_3529,N_1786,N_1768);
and U3530 (N_3530,N_274,N_1116);
nor U3531 (N_3531,N_1250,N_985);
nand U3532 (N_3532,N_934,N_149);
xnor U3533 (N_3533,N_1286,N_811);
nor U3534 (N_3534,N_488,N_1772);
nand U3535 (N_3535,N_1870,N_705);
xnor U3536 (N_3536,N_1797,N_1032);
and U3537 (N_3537,N_945,N_1965);
and U3538 (N_3538,N_152,N_1671);
and U3539 (N_3539,N_574,N_1352);
xnor U3540 (N_3540,N_887,N_690);
or U3541 (N_3541,N_1015,N_1851);
nand U3542 (N_3542,N_1896,N_221);
xor U3543 (N_3543,N_909,N_845);
nor U3544 (N_3544,N_1510,N_1764);
nor U3545 (N_3545,N_929,N_882);
or U3546 (N_3546,N_140,N_1042);
or U3547 (N_3547,N_902,N_1945);
or U3548 (N_3548,N_668,N_522);
xor U3549 (N_3549,N_1222,N_181);
xor U3550 (N_3550,N_644,N_1150);
xnor U3551 (N_3551,N_967,N_905);
xnor U3552 (N_3552,N_613,N_261);
xnor U3553 (N_3553,N_1814,N_1307);
or U3554 (N_3554,N_1548,N_1004);
nand U3555 (N_3555,N_425,N_1413);
or U3556 (N_3556,N_63,N_1135);
or U3557 (N_3557,N_659,N_597);
and U3558 (N_3558,N_562,N_1079);
xor U3559 (N_3559,N_1037,N_1534);
or U3560 (N_3560,N_690,N_1858);
nand U3561 (N_3561,N_1871,N_1245);
or U3562 (N_3562,N_1117,N_446);
xor U3563 (N_3563,N_1282,N_670);
and U3564 (N_3564,N_1045,N_1042);
nor U3565 (N_3565,N_1650,N_1513);
xnor U3566 (N_3566,N_570,N_707);
and U3567 (N_3567,N_793,N_510);
nor U3568 (N_3568,N_82,N_1495);
or U3569 (N_3569,N_1516,N_817);
nor U3570 (N_3570,N_1628,N_1980);
and U3571 (N_3571,N_1759,N_1763);
nand U3572 (N_3572,N_155,N_509);
and U3573 (N_3573,N_1717,N_360);
and U3574 (N_3574,N_1621,N_780);
nor U3575 (N_3575,N_354,N_1905);
xor U3576 (N_3576,N_749,N_1330);
xor U3577 (N_3577,N_1545,N_1426);
or U3578 (N_3578,N_1778,N_1532);
nand U3579 (N_3579,N_990,N_1775);
nand U3580 (N_3580,N_1173,N_1457);
or U3581 (N_3581,N_1859,N_303);
nand U3582 (N_3582,N_59,N_1755);
or U3583 (N_3583,N_481,N_764);
and U3584 (N_3584,N_1708,N_541);
nand U3585 (N_3585,N_1456,N_222);
nand U3586 (N_3586,N_1286,N_7);
nand U3587 (N_3587,N_1628,N_1542);
xor U3588 (N_3588,N_726,N_1810);
nand U3589 (N_3589,N_1181,N_330);
nor U3590 (N_3590,N_18,N_973);
and U3591 (N_3591,N_254,N_306);
or U3592 (N_3592,N_448,N_1471);
xor U3593 (N_3593,N_1190,N_964);
xnor U3594 (N_3594,N_1735,N_908);
xnor U3595 (N_3595,N_378,N_254);
or U3596 (N_3596,N_180,N_54);
and U3597 (N_3597,N_1213,N_1071);
xnor U3598 (N_3598,N_237,N_226);
xnor U3599 (N_3599,N_65,N_741);
nor U3600 (N_3600,N_1874,N_265);
xor U3601 (N_3601,N_250,N_268);
nand U3602 (N_3602,N_633,N_1119);
or U3603 (N_3603,N_311,N_1992);
xor U3604 (N_3604,N_436,N_365);
nor U3605 (N_3605,N_1980,N_1962);
and U3606 (N_3606,N_410,N_261);
xnor U3607 (N_3607,N_132,N_1514);
nor U3608 (N_3608,N_1931,N_458);
or U3609 (N_3609,N_1093,N_1395);
nor U3610 (N_3610,N_386,N_588);
and U3611 (N_3611,N_1498,N_1701);
nor U3612 (N_3612,N_1557,N_1876);
or U3613 (N_3613,N_391,N_1251);
xor U3614 (N_3614,N_586,N_1572);
and U3615 (N_3615,N_375,N_96);
nor U3616 (N_3616,N_1430,N_282);
nand U3617 (N_3617,N_885,N_1287);
xor U3618 (N_3618,N_968,N_860);
or U3619 (N_3619,N_199,N_1410);
nor U3620 (N_3620,N_1061,N_613);
nand U3621 (N_3621,N_1331,N_1470);
xnor U3622 (N_3622,N_1428,N_547);
xnor U3623 (N_3623,N_661,N_1787);
nor U3624 (N_3624,N_1456,N_1055);
or U3625 (N_3625,N_733,N_151);
or U3626 (N_3626,N_621,N_989);
xor U3627 (N_3627,N_1220,N_1315);
and U3628 (N_3628,N_76,N_1588);
nand U3629 (N_3629,N_212,N_221);
xor U3630 (N_3630,N_578,N_682);
xnor U3631 (N_3631,N_707,N_1166);
nor U3632 (N_3632,N_1461,N_457);
and U3633 (N_3633,N_1245,N_1758);
and U3634 (N_3634,N_1211,N_1583);
nand U3635 (N_3635,N_705,N_301);
nand U3636 (N_3636,N_1275,N_822);
and U3637 (N_3637,N_318,N_499);
nand U3638 (N_3638,N_452,N_1705);
nand U3639 (N_3639,N_1869,N_666);
nor U3640 (N_3640,N_362,N_1159);
nor U3641 (N_3641,N_1023,N_390);
nand U3642 (N_3642,N_1046,N_503);
or U3643 (N_3643,N_1849,N_1786);
nand U3644 (N_3644,N_1530,N_1246);
xor U3645 (N_3645,N_361,N_1429);
or U3646 (N_3646,N_141,N_299);
and U3647 (N_3647,N_1738,N_655);
or U3648 (N_3648,N_1772,N_1752);
xor U3649 (N_3649,N_466,N_1155);
xnor U3650 (N_3650,N_314,N_863);
nand U3651 (N_3651,N_1555,N_1869);
nand U3652 (N_3652,N_1452,N_1207);
nand U3653 (N_3653,N_1682,N_1877);
xor U3654 (N_3654,N_633,N_333);
and U3655 (N_3655,N_1481,N_1469);
xor U3656 (N_3656,N_939,N_1295);
or U3657 (N_3657,N_383,N_832);
or U3658 (N_3658,N_298,N_635);
xnor U3659 (N_3659,N_1838,N_1149);
nand U3660 (N_3660,N_67,N_956);
xnor U3661 (N_3661,N_1742,N_1579);
xor U3662 (N_3662,N_1904,N_1970);
xor U3663 (N_3663,N_740,N_1221);
or U3664 (N_3664,N_1243,N_568);
nor U3665 (N_3665,N_369,N_1672);
or U3666 (N_3666,N_1989,N_1481);
nor U3667 (N_3667,N_1777,N_1491);
xor U3668 (N_3668,N_1611,N_1418);
and U3669 (N_3669,N_654,N_187);
nand U3670 (N_3670,N_1454,N_1227);
nand U3671 (N_3671,N_1250,N_559);
nor U3672 (N_3672,N_1181,N_1018);
and U3673 (N_3673,N_1345,N_1996);
xor U3674 (N_3674,N_147,N_370);
xnor U3675 (N_3675,N_129,N_993);
or U3676 (N_3676,N_1250,N_1768);
nand U3677 (N_3677,N_950,N_1753);
or U3678 (N_3678,N_1803,N_1717);
or U3679 (N_3679,N_522,N_464);
nor U3680 (N_3680,N_1184,N_724);
nor U3681 (N_3681,N_154,N_184);
nor U3682 (N_3682,N_11,N_1201);
nor U3683 (N_3683,N_813,N_283);
xor U3684 (N_3684,N_1599,N_1577);
nor U3685 (N_3685,N_82,N_419);
nand U3686 (N_3686,N_1456,N_1969);
nor U3687 (N_3687,N_1474,N_750);
xor U3688 (N_3688,N_572,N_404);
nand U3689 (N_3689,N_546,N_324);
xnor U3690 (N_3690,N_699,N_569);
nand U3691 (N_3691,N_251,N_860);
nand U3692 (N_3692,N_1668,N_993);
and U3693 (N_3693,N_113,N_458);
nand U3694 (N_3694,N_897,N_1173);
nand U3695 (N_3695,N_993,N_1673);
and U3696 (N_3696,N_1725,N_1922);
nand U3697 (N_3697,N_1420,N_111);
xor U3698 (N_3698,N_1727,N_621);
xor U3699 (N_3699,N_113,N_638);
and U3700 (N_3700,N_1021,N_653);
or U3701 (N_3701,N_425,N_798);
nor U3702 (N_3702,N_1647,N_1637);
and U3703 (N_3703,N_426,N_743);
nor U3704 (N_3704,N_1847,N_293);
xor U3705 (N_3705,N_1284,N_1386);
or U3706 (N_3706,N_1707,N_1046);
or U3707 (N_3707,N_956,N_1791);
xnor U3708 (N_3708,N_802,N_1157);
or U3709 (N_3709,N_80,N_1213);
or U3710 (N_3710,N_1575,N_1145);
or U3711 (N_3711,N_1887,N_589);
xnor U3712 (N_3712,N_1648,N_315);
nand U3713 (N_3713,N_1277,N_377);
and U3714 (N_3714,N_1200,N_76);
xor U3715 (N_3715,N_340,N_483);
and U3716 (N_3716,N_629,N_973);
nand U3717 (N_3717,N_1598,N_678);
and U3718 (N_3718,N_1580,N_909);
xnor U3719 (N_3719,N_85,N_1411);
and U3720 (N_3720,N_1788,N_1560);
nor U3721 (N_3721,N_1477,N_1036);
nand U3722 (N_3722,N_43,N_159);
and U3723 (N_3723,N_440,N_1021);
or U3724 (N_3724,N_1483,N_1779);
or U3725 (N_3725,N_1679,N_1874);
xnor U3726 (N_3726,N_1097,N_1591);
xnor U3727 (N_3727,N_1557,N_40);
xnor U3728 (N_3728,N_1117,N_1879);
nor U3729 (N_3729,N_1016,N_900);
or U3730 (N_3730,N_1295,N_438);
and U3731 (N_3731,N_1593,N_143);
or U3732 (N_3732,N_28,N_529);
nand U3733 (N_3733,N_1308,N_626);
nor U3734 (N_3734,N_1479,N_1214);
nand U3735 (N_3735,N_1673,N_1645);
and U3736 (N_3736,N_1517,N_1394);
or U3737 (N_3737,N_671,N_631);
and U3738 (N_3738,N_1279,N_1024);
or U3739 (N_3739,N_1302,N_215);
or U3740 (N_3740,N_1515,N_242);
and U3741 (N_3741,N_1750,N_1680);
and U3742 (N_3742,N_1444,N_341);
xnor U3743 (N_3743,N_1416,N_1183);
nor U3744 (N_3744,N_690,N_112);
nand U3745 (N_3745,N_1237,N_1033);
nor U3746 (N_3746,N_515,N_167);
and U3747 (N_3747,N_146,N_646);
or U3748 (N_3748,N_370,N_59);
and U3749 (N_3749,N_484,N_612);
xor U3750 (N_3750,N_849,N_147);
nand U3751 (N_3751,N_1651,N_1910);
nor U3752 (N_3752,N_1805,N_1117);
nand U3753 (N_3753,N_1086,N_1984);
and U3754 (N_3754,N_475,N_1091);
and U3755 (N_3755,N_1951,N_54);
nand U3756 (N_3756,N_1732,N_1000);
xor U3757 (N_3757,N_1729,N_1515);
nor U3758 (N_3758,N_341,N_1375);
xor U3759 (N_3759,N_1766,N_222);
nor U3760 (N_3760,N_959,N_581);
or U3761 (N_3761,N_895,N_1339);
or U3762 (N_3762,N_269,N_1);
or U3763 (N_3763,N_775,N_1225);
nand U3764 (N_3764,N_166,N_934);
and U3765 (N_3765,N_556,N_1516);
nor U3766 (N_3766,N_1839,N_1728);
and U3767 (N_3767,N_876,N_314);
xnor U3768 (N_3768,N_941,N_664);
and U3769 (N_3769,N_1950,N_1044);
nand U3770 (N_3770,N_638,N_1047);
and U3771 (N_3771,N_1686,N_325);
nand U3772 (N_3772,N_1487,N_732);
nor U3773 (N_3773,N_1839,N_385);
nand U3774 (N_3774,N_211,N_1046);
xor U3775 (N_3775,N_451,N_375);
xnor U3776 (N_3776,N_1409,N_442);
xnor U3777 (N_3777,N_182,N_1269);
nand U3778 (N_3778,N_1154,N_1853);
or U3779 (N_3779,N_658,N_822);
nand U3780 (N_3780,N_497,N_414);
or U3781 (N_3781,N_1304,N_1012);
xor U3782 (N_3782,N_1896,N_130);
or U3783 (N_3783,N_1994,N_1056);
or U3784 (N_3784,N_1412,N_637);
nand U3785 (N_3785,N_1678,N_170);
xnor U3786 (N_3786,N_1489,N_243);
nand U3787 (N_3787,N_1296,N_1841);
nor U3788 (N_3788,N_324,N_1965);
nand U3789 (N_3789,N_1013,N_1158);
nand U3790 (N_3790,N_578,N_3);
xor U3791 (N_3791,N_1441,N_818);
nand U3792 (N_3792,N_1928,N_1163);
and U3793 (N_3793,N_984,N_1385);
and U3794 (N_3794,N_1860,N_479);
nand U3795 (N_3795,N_1489,N_1479);
nor U3796 (N_3796,N_550,N_171);
or U3797 (N_3797,N_936,N_498);
xor U3798 (N_3798,N_1013,N_469);
nand U3799 (N_3799,N_1117,N_1186);
or U3800 (N_3800,N_900,N_925);
nor U3801 (N_3801,N_1627,N_97);
nor U3802 (N_3802,N_602,N_597);
or U3803 (N_3803,N_1070,N_499);
nor U3804 (N_3804,N_1236,N_854);
xnor U3805 (N_3805,N_210,N_1540);
nand U3806 (N_3806,N_1255,N_372);
nand U3807 (N_3807,N_1684,N_1757);
and U3808 (N_3808,N_1218,N_1805);
nor U3809 (N_3809,N_1106,N_576);
xnor U3810 (N_3810,N_937,N_953);
nor U3811 (N_3811,N_72,N_1878);
and U3812 (N_3812,N_66,N_372);
or U3813 (N_3813,N_259,N_580);
nand U3814 (N_3814,N_1088,N_1595);
xor U3815 (N_3815,N_9,N_279);
nor U3816 (N_3816,N_598,N_1467);
or U3817 (N_3817,N_1578,N_136);
xnor U3818 (N_3818,N_1425,N_302);
nor U3819 (N_3819,N_970,N_1908);
nand U3820 (N_3820,N_1462,N_105);
and U3821 (N_3821,N_1290,N_1183);
or U3822 (N_3822,N_1755,N_663);
nand U3823 (N_3823,N_770,N_756);
xor U3824 (N_3824,N_1440,N_1646);
or U3825 (N_3825,N_56,N_137);
xor U3826 (N_3826,N_909,N_79);
nor U3827 (N_3827,N_1328,N_406);
or U3828 (N_3828,N_1847,N_499);
xnor U3829 (N_3829,N_371,N_1281);
nand U3830 (N_3830,N_951,N_1902);
and U3831 (N_3831,N_472,N_699);
and U3832 (N_3832,N_708,N_269);
nand U3833 (N_3833,N_1605,N_1666);
and U3834 (N_3834,N_748,N_402);
and U3835 (N_3835,N_947,N_1780);
or U3836 (N_3836,N_525,N_1299);
nor U3837 (N_3837,N_1744,N_1937);
nor U3838 (N_3838,N_1265,N_1231);
and U3839 (N_3839,N_675,N_1921);
and U3840 (N_3840,N_132,N_139);
nand U3841 (N_3841,N_571,N_156);
or U3842 (N_3842,N_789,N_1307);
and U3843 (N_3843,N_650,N_1537);
nand U3844 (N_3844,N_85,N_1753);
nand U3845 (N_3845,N_1779,N_1756);
and U3846 (N_3846,N_1133,N_1197);
xor U3847 (N_3847,N_706,N_617);
nor U3848 (N_3848,N_1978,N_1612);
nand U3849 (N_3849,N_1118,N_1234);
nor U3850 (N_3850,N_893,N_490);
nand U3851 (N_3851,N_827,N_1281);
and U3852 (N_3852,N_483,N_1123);
nand U3853 (N_3853,N_1332,N_604);
or U3854 (N_3854,N_1620,N_291);
and U3855 (N_3855,N_1536,N_70);
nor U3856 (N_3856,N_1811,N_598);
nand U3857 (N_3857,N_777,N_1607);
or U3858 (N_3858,N_1963,N_1927);
nor U3859 (N_3859,N_1622,N_336);
nand U3860 (N_3860,N_1553,N_1066);
nand U3861 (N_3861,N_194,N_483);
nand U3862 (N_3862,N_1777,N_898);
xor U3863 (N_3863,N_1336,N_705);
and U3864 (N_3864,N_589,N_1505);
xnor U3865 (N_3865,N_1564,N_1820);
nor U3866 (N_3866,N_662,N_836);
and U3867 (N_3867,N_1159,N_1496);
or U3868 (N_3868,N_1966,N_747);
xnor U3869 (N_3869,N_351,N_645);
xor U3870 (N_3870,N_476,N_706);
and U3871 (N_3871,N_1205,N_1042);
or U3872 (N_3872,N_1076,N_1530);
nor U3873 (N_3873,N_1089,N_1179);
nor U3874 (N_3874,N_408,N_485);
nor U3875 (N_3875,N_160,N_520);
or U3876 (N_3876,N_502,N_1584);
nand U3877 (N_3877,N_1847,N_1258);
nand U3878 (N_3878,N_243,N_744);
xnor U3879 (N_3879,N_1314,N_1970);
xnor U3880 (N_3880,N_1753,N_1135);
xor U3881 (N_3881,N_1053,N_915);
xnor U3882 (N_3882,N_1864,N_1537);
and U3883 (N_3883,N_898,N_1984);
nand U3884 (N_3884,N_1728,N_1708);
or U3885 (N_3885,N_1586,N_1136);
or U3886 (N_3886,N_332,N_151);
and U3887 (N_3887,N_511,N_1572);
and U3888 (N_3888,N_1691,N_253);
nor U3889 (N_3889,N_1861,N_1481);
or U3890 (N_3890,N_1548,N_999);
and U3891 (N_3891,N_1783,N_498);
nor U3892 (N_3892,N_1304,N_481);
and U3893 (N_3893,N_874,N_1427);
xor U3894 (N_3894,N_964,N_1126);
and U3895 (N_3895,N_1661,N_1461);
nor U3896 (N_3896,N_1755,N_56);
or U3897 (N_3897,N_271,N_769);
xnor U3898 (N_3898,N_119,N_1558);
xor U3899 (N_3899,N_1414,N_1401);
and U3900 (N_3900,N_186,N_1352);
nor U3901 (N_3901,N_112,N_1556);
nor U3902 (N_3902,N_605,N_164);
and U3903 (N_3903,N_622,N_751);
xor U3904 (N_3904,N_1619,N_1454);
nor U3905 (N_3905,N_1144,N_655);
and U3906 (N_3906,N_1223,N_1032);
or U3907 (N_3907,N_134,N_1413);
or U3908 (N_3908,N_462,N_1065);
and U3909 (N_3909,N_266,N_43);
nand U3910 (N_3910,N_745,N_1273);
xor U3911 (N_3911,N_1995,N_316);
xnor U3912 (N_3912,N_1291,N_1490);
xor U3913 (N_3913,N_807,N_1668);
nand U3914 (N_3914,N_1263,N_1466);
and U3915 (N_3915,N_1873,N_1210);
nor U3916 (N_3916,N_518,N_526);
and U3917 (N_3917,N_868,N_248);
nor U3918 (N_3918,N_1681,N_931);
and U3919 (N_3919,N_1051,N_1234);
nand U3920 (N_3920,N_852,N_1840);
nand U3921 (N_3921,N_495,N_1755);
and U3922 (N_3922,N_1156,N_227);
nor U3923 (N_3923,N_71,N_1884);
xor U3924 (N_3924,N_1963,N_88);
nor U3925 (N_3925,N_1913,N_1204);
nor U3926 (N_3926,N_1433,N_1573);
and U3927 (N_3927,N_965,N_316);
and U3928 (N_3928,N_58,N_470);
or U3929 (N_3929,N_578,N_1589);
nand U3930 (N_3930,N_469,N_326);
or U3931 (N_3931,N_333,N_493);
xnor U3932 (N_3932,N_1789,N_298);
nand U3933 (N_3933,N_215,N_315);
nor U3934 (N_3934,N_1311,N_1125);
or U3935 (N_3935,N_73,N_1768);
and U3936 (N_3936,N_352,N_114);
xnor U3937 (N_3937,N_350,N_187);
nand U3938 (N_3938,N_1577,N_470);
nand U3939 (N_3939,N_1445,N_943);
or U3940 (N_3940,N_1627,N_239);
xor U3941 (N_3941,N_1053,N_43);
or U3942 (N_3942,N_82,N_35);
or U3943 (N_3943,N_620,N_409);
and U3944 (N_3944,N_1706,N_236);
or U3945 (N_3945,N_1733,N_308);
and U3946 (N_3946,N_415,N_414);
xnor U3947 (N_3947,N_824,N_1361);
nand U3948 (N_3948,N_1555,N_1540);
xnor U3949 (N_3949,N_1120,N_840);
or U3950 (N_3950,N_1105,N_279);
nand U3951 (N_3951,N_202,N_1814);
or U3952 (N_3952,N_665,N_1119);
nand U3953 (N_3953,N_1854,N_1168);
or U3954 (N_3954,N_50,N_116);
xnor U3955 (N_3955,N_1670,N_1277);
nand U3956 (N_3956,N_1591,N_9);
nor U3957 (N_3957,N_53,N_396);
or U3958 (N_3958,N_786,N_1824);
nor U3959 (N_3959,N_1590,N_579);
nand U3960 (N_3960,N_184,N_1554);
nand U3961 (N_3961,N_646,N_1388);
nand U3962 (N_3962,N_1397,N_192);
or U3963 (N_3963,N_1709,N_813);
and U3964 (N_3964,N_1070,N_99);
nand U3965 (N_3965,N_1304,N_104);
and U3966 (N_3966,N_200,N_1657);
or U3967 (N_3967,N_315,N_910);
xnor U3968 (N_3968,N_1422,N_646);
xor U3969 (N_3969,N_1837,N_1121);
and U3970 (N_3970,N_276,N_1193);
nor U3971 (N_3971,N_388,N_1925);
and U3972 (N_3972,N_1948,N_139);
and U3973 (N_3973,N_329,N_1267);
or U3974 (N_3974,N_1285,N_490);
and U3975 (N_3975,N_574,N_1715);
nor U3976 (N_3976,N_1040,N_1723);
xor U3977 (N_3977,N_1114,N_1686);
nand U3978 (N_3978,N_1145,N_1431);
or U3979 (N_3979,N_648,N_178);
and U3980 (N_3980,N_967,N_1409);
and U3981 (N_3981,N_1012,N_567);
nand U3982 (N_3982,N_49,N_523);
and U3983 (N_3983,N_690,N_53);
or U3984 (N_3984,N_816,N_600);
xor U3985 (N_3985,N_484,N_361);
and U3986 (N_3986,N_672,N_437);
xor U3987 (N_3987,N_1322,N_1269);
nor U3988 (N_3988,N_817,N_899);
and U3989 (N_3989,N_1033,N_909);
and U3990 (N_3990,N_1302,N_1636);
xnor U3991 (N_3991,N_943,N_1768);
xnor U3992 (N_3992,N_1329,N_1155);
or U3993 (N_3993,N_25,N_802);
nor U3994 (N_3994,N_508,N_1815);
nor U3995 (N_3995,N_1695,N_209);
nor U3996 (N_3996,N_1013,N_14);
xor U3997 (N_3997,N_1316,N_450);
xor U3998 (N_3998,N_224,N_871);
nand U3999 (N_3999,N_1363,N_399);
and U4000 (N_4000,N_2712,N_3451);
nor U4001 (N_4001,N_3060,N_2825);
and U4002 (N_4002,N_3048,N_2340);
and U4003 (N_4003,N_3178,N_2626);
xor U4004 (N_4004,N_3753,N_3649);
or U4005 (N_4005,N_2111,N_2505);
or U4006 (N_4006,N_2030,N_2023);
and U4007 (N_4007,N_2837,N_2617);
and U4008 (N_4008,N_3425,N_2128);
and U4009 (N_4009,N_3518,N_2155);
or U4010 (N_4010,N_2765,N_2553);
and U4011 (N_4011,N_3865,N_2539);
xor U4012 (N_4012,N_2809,N_3303);
nor U4013 (N_4013,N_3053,N_2802);
xnor U4014 (N_4014,N_3429,N_2109);
and U4015 (N_4015,N_3251,N_3783);
or U4016 (N_4016,N_3078,N_2642);
or U4017 (N_4017,N_2671,N_3692);
nor U4018 (N_4018,N_2136,N_3482);
xor U4019 (N_4019,N_2740,N_3505);
and U4020 (N_4020,N_2010,N_3152);
or U4021 (N_4021,N_2885,N_2278);
and U4022 (N_4022,N_3222,N_2908);
nor U4023 (N_4023,N_2338,N_2421);
or U4024 (N_4024,N_3224,N_3587);
or U4025 (N_4025,N_2824,N_3698);
nor U4026 (N_4026,N_2643,N_2205);
or U4027 (N_4027,N_3439,N_3018);
or U4028 (N_4028,N_2273,N_3690);
nor U4029 (N_4029,N_2488,N_2558);
nand U4030 (N_4030,N_2075,N_3030);
nor U4031 (N_4031,N_2619,N_2601);
xnor U4032 (N_4032,N_2866,N_3094);
xor U4033 (N_4033,N_2146,N_2131);
nor U4034 (N_4034,N_2050,N_2298);
nor U4035 (N_4035,N_2310,N_2202);
nor U4036 (N_4036,N_3000,N_2172);
and U4037 (N_4037,N_2480,N_3384);
xnor U4038 (N_4038,N_3879,N_2972);
or U4039 (N_4039,N_2046,N_2141);
nor U4040 (N_4040,N_2938,N_2479);
and U4041 (N_4041,N_2341,N_3401);
nand U4042 (N_4042,N_3794,N_3723);
or U4043 (N_4043,N_2410,N_3497);
nor U4044 (N_4044,N_3234,N_3092);
or U4045 (N_4045,N_3858,N_2495);
nand U4046 (N_4046,N_3028,N_2428);
nor U4047 (N_4047,N_3928,N_3211);
or U4048 (N_4048,N_2876,N_3077);
nor U4049 (N_4049,N_3380,N_2035);
or U4050 (N_4050,N_3485,N_3866);
nor U4051 (N_4051,N_3165,N_2316);
nor U4052 (N_4052,N_3325,N_3336);
nand U4053 (N_4053,N_3186,N_3243);
and U4054 (N_4054,N_2174,N_2842);
or U4055 (N_4055,N_2276,N_2054);
nor U4056 (N_4056,N_3750,N_3113);
and U4057 (N_4057,N_3841,N_3472);
nor U4058 (N_4058,N_3755,N_3571);
nand U4059 (N_4059,N_2964,N_2510);
and U4060 (N_4060,N_2651,N_2058);
nor U4061 (N_4061,N_2548,N_3019);
xnor U4062 (N_4062,N_3507,N_2110);
nor U4063 (N_4063,N_2628,N_3300);
and U4064 (N_4064,N_3566,N_3233);
nand U4065 (N_4065,N_2597,N_2369);
and U4066 (N_4066,N_2300,N_3716);
and U4067 (N_4067,N_2345,N_2992);
or U4068 (N_4068,N_2019,N_2086);
nor U4069 (N_4069,N_3607,N_3326);
nor U4070 (N_4070,N_2847,N_2411);
nand U4071 (N_4071,N_2855,N_3670);
or U4072 (N_4072,N_2691,N_2040);
nor U4073 (N_4073,N_2520,N_3765);
xnor U4074 (N_4074,N_3985,N_3771);
or U4075 (N_4075,N_3150,N_3015);
and U4076 (N_4076,N_2875,N_2534);
xnor U4077 (N_4077,N_3864,N_2948);
or U4078 (N_4078,N_2192,N_2733);
and U4079 (N_4079,N_2043,N_2906);
and U4080 (N_4080,N_2929,N_3982);
and U4081 (N_4081,N_3634,N_2120);
nor U4082 (N_4082,N_3669,N_2838);
xor U4083 (N_4083,N_3702,N_2841);
nor U4084 (N_4084,N_2394,N_3084);
and U4085 (N_4085,N_3969,N_3544);
and U4086 (N_4086,N_2660,N_2937);
nand U4087 (N_4087,N_2468,N_3006);
nand U4088 (N_4088,N_2731,N_2004);
xor U4089 (N_4089,N_3342,N_2044);
xnor U4090 (N_4090,N_3455,N_2777);
nor U4091 (N_4091,N_2445,N_2674);
or U4092 (N_4092,N_3085,N_3091);
and U4093 (N_4093,N_3321,N_3148);
nor U4094 (N_4094,N_3740,N_3923);
or U4095 (N_4095,N_3469,N_2508);
nor U4096 (N_4096,N_2684,N_2730);
nand U4097 (N_4097,N_3288,N_2081);
or U4098 (N_4098,N_3855,N_3947);
and U4099 (N_4099,N_2658,N_3960);
and U4100 (N_4100,N_2181,N_2311);
or U4101 (N_4101,N_2159,N_3805);
and U4102 (N_4102,N_3108,N_2869);
and U4103 (N_4103,N_2725,N_2271);
nor U4104 (N_4104,N_2203,N_3216);
nand U4105 (N_4105,N_3473,N_2602);
and U4106 (N_4106,N_3868,N_3263);
nand U4107 (N_4107,N_2683,N_2576);
xnor U4108 (N_4108,N_2130,N_2523);
nand U4109 (N_4109,N_3900,N_2754);
xnor U4110 (N_4110,N_3075,N_3559);
nor U4111 (N_4111,N_3843,N_3857);
xor U4112 (N_4112,N_3652,N_3972);
nand U4113 (N_4113,N_2017,N_3047);
or U4114 (N_4114,N_2859,N_3218);
or U4115 (N_4115,N_3813,N_2543);
and U4116 (N_4116,N_3415,N_3361);
or U4117 (N_4117,N_2836,N_3659);
xor U4118 (N_4118,N_2060,N_2581);
nor U4119 (N_4119,N_2283,N_2582);
or U4120 (N_4120,N_2727,N_3207);
and U4121 (N_4121,N_2527,N_2724);
or U4122 (N_4122,N_2749,N_3126);
and U4123 (N_4123,N_3149,N_2280);
or U4124 (N_4124,N_2610,N_2812);
and U4125 (N_4125,N_3433,N_3671);
nand U4126 (N_4126,N_3219,N_3271);
and U4127 (N_4127,N_3264,N_2465);
and U4128 (N_4128,N_2206,N_2710);
nand U4129 (N_4129,N_3119,N_2393);
and U4130 (N_4130,N_3307,N_2641);
nand U4131 (N_4131,N_2541,N_3774);
or U4132 (N_4132,N_3529,N_2528);
or U4133 (N_4133,N_3557,N_2844);
xor U4134 (N_4134,N_2041,N_2827);
or U4135 (N_4135,N_3190,N_3594);
and U4136 (N_4136,N_3476,N_3435);
nor U4137 (N_4137,N_2376,N_2536);
and U4138 (N_4138,N_2819,N_3072);
and U4139 (N_4139,N_3260,N_3761);
and U4140 (N_4140,N_3672,N_3605);
nor U4141 (N_4141,N_3088,N_2336);
nand U4142 (N_4142,N_3886,N_3945);
xnor U4143 (N_4143,N_2848,N_3310);
and U4144 (N_4144,N_3167,N_3426);
nor U4145 (N_4145,N_2484,N_3188);
or U4146 (N_4146,N_2669,N_3952);
nand U4147 (N_4147,N_2834,N_2974);
nor U4148 (N_4148,N_3964,N_3316);
nand U4149 (N_4149,N_3498,N_3158);
xnor U4150 (N_4150,N_2121,N_2138);
xnor U4151 (N_4151,N_2059,N_3565);
xnor U4152 (N_4152,N_2144,N_2384);
nor U4153 (N_4153,N_3226,N_3798);
or U4154 (N_4154,N_2419,N_3474);
and U4155 (N_4155,N_2542,N_3296);
or U4156 (N_4156,N_3593,N_2170);
xnor U4157 (N_4157,N_3372,N_2851);
and U4158 (N_4158,N_3250,N_3647);
and U4159 (N_4159,N_3416,N_3424);
or U4160 (N_4160,N_2365,N_3773);
or U4161 (N_4161,N_3630,N_2688);
xnor U4162 (N_4162,N_2134,N_3792);
and U4163 (N_4163,N_3542,N_3290);
nand U4164 (N_4164,N_3730,N_3737);
nor U4165 (N_4165,N_2220,N_2563);
or U4166 (N_4166,N_2188,N_2180);
or U4167 (N_4167,N_3751,N_2404);
or U4168 (N_4168,N_2042,N_2962);
nor U4169 (N_4169,N_2627,N_3946);
nand U4170 (N_4170,N_3441,N_3231);
xor U4171 (N_4171,N_2092,N_3448);
nand U4172 (N_4172,N_2274,N_2381);
nor U4173 (N_4173,N_2647,N_3430);
or U4174 (N_4174,N_2382,N_2450);
and U4175 (N_4175,N_2103,N_3540);
xor U4176 (N_4176,N_3941,N_2313);
nor U4177 (N_4177,N_3450,N_3725);
xor U4178 (N_4178,N_2537,N_3990);
or U4179 (N_4179,N_3963,N_2097);
xnor U4180 (N_4180,N_2478,N_3143);
xnor U4181 (N_4181,N_3552,N_3099);
nor U4182 (N_4182,N_3357,N_3714);
nor U4183 (N_4183,N_2966,N_3703);
and U4184 (N_4184,N_3916,N_3490);
or U4185 (N_4185,N_3574,N_3353);
nor U4186 (N_4186,N_3686,N_2232);
nand U4187 (N_4187,N_3554,N_3056);
or U4188 (N_4188,N_3598,N_3790);
and U4189 (N_4189,N_3758,N_3892);
nor U4190 (N_4190,N_2608,N_3169);
and U4191 (N_4191,N_2227,N_2614);
nand U4192 (N_4192,N_2811,N_3459);
xor U4193 (N_4193,N_2516,N_3975);
or U4194 (N_4194,N_3155,N_2907);
and U4195 (N_4195,N_2293,N_2073);
nand U4196 (N_4196,N_2057,N_2920);
nand U4197 (N_4197,N_2100,N_3784);
xnor U4198 (N_4198,N_2151,N_3355);
and U4199 (N_4199,N_3971,N_3317);
xnor U4200 (N_4200,N_3715,N_3801);
or U4201 (N_4201,N_2234,N_3768);
or U4202 (N_4202,N_2678,N_2941);
nand U4203 (N_4203,N_2822,N_3050);
or U4204 (N_4204,N_3144,N_2464);
nand U4205 (N_4205,N_3732,N_2064);
or U4206 (N_4206,N_2716,N_3145);
and U4207 (N_4207,N_2457,N_3778);
and U4208 (N_4208,N_2786,N_2157);
and U4209 (N_4209,N_3181,N_3663);
xnor U4210 (N_4210,N_3406,N_2106);
nor U4211 (N_4211,N_2424,N_2037);
xnor U4212 (N_4212,N_2489,N_2795);
or U4213 (N_4213,N_2870,N_3277);
or U4214 (N_4214,N_3724,N_3107);
and U4215 (N_4215,N_3125,N_3951);
or U4216 (N_4216,N_3539,N_2009);
and U4217 (N_4217,N_2263,N_2705);
nor U4218 (N_4218,N_3039,N_3654);
or U4219 (N_4219,N_3022,N_2270);
nor U4220 (N_4220,N_2633,N_2832);
xnor U4221 (N_4221,N_2208,N_3863);
nor U4222 (N_4222,N_3292,N_2703);
or U4223 (N_4223,N_2997,N_3676);
nor U4224 (N_4224,N_2024,N_3710);
xor U4225 (N_4225,N_3176,N_2856);
and U4226 (N_4226,N_2281,N_3709);
or U4227 (N_4227,N_3489,N_2115);
nand U4228 (N_4228,N_2509,N_2448);
nand U4229 (N_4229,N_3583,N_2784);
or U4230 (N_4230,N_2342,N_3867);
or U4231 (N_4231,N_3405,N_3197);
nand U4232 (N_4232,N_3334,N_2659);
or U4233 (N_4233,N_3352,N_2061);
nor U4234 (N_4234,N_3066,N_2447);
or U4235 (N_4235,N_2596,N_2461);
or U4236 (N_4236,N_2118,N_3480);
nand U4237 (N_4237,N_3744,N_2360);
nor U4238 (N_4238,N_3931,N_2872);
nand U4239 (N_4239,N_3453,N_2820);
xor U4240 (N_4240,N_2637,N_3255);
or U4241 (N_4241,N_2918,N_2069);
xnor U4242 (N_4242,N_3180,N_3393);
nor U4243 (N_4243,N_2511,N_2089);
or U4244 (N_4244,N_3719,N_3688);
or U4245 (N_4245,N_2052,N_2254);
or U4246 (N_4246,N_2355,N_2493);
nand U4247 (N_4247,N_2752,N_2736);
and U4248 (N_4248,N_3562,N_3599);
xnor U4249 (N_4249,N_2771,N_2126);
nand U4250 (N_4250,N_2165,N_3872);
xnor U4251 (N_4251,N_2331,N_3697);
and U4252 (N_4252,N_2681,N_2833);
xor U4253 (N_4253,N_3658,N_3403);
or U4254 (N_4254,N_2446,N_2353);
xnor U4255 (N_4255,N_3936,N_2147);
xnor U4256 (N_4256,N_3713,N_3304);
nand U4257 (N_4257,N_2922,N_3524);
xnor U4258 (N_4258,N_2741,N_3641);
xnor U4259 (N_4259,N_3076,N_2850);
and U4260 (N_4260,N_2008,N_2378);
or U4261 (N_4261,N_2569,N_2169);
xor U4262 (N_4262,N_2803,N_3760);
or U4263 (N_4263,N_2959,N_3547);
and U4264 (N_4264,N_2645,N_2574);
nor U4265 (N_4265,N_3901,N_3828);
xor U4266 (N_4266,N_2570,N_3035);
xnor U4267 (N_4267,N_2142,N_3285);
nor U4268 (N_4268,N_2638,N_2483);
or U4269 (N_4269,N_3166,N_2277);
nor U4270 (N_4270,N_2506,N_3914);
xnor U4271 (N_4271,N_3021,N_2685);
xnor U4272 (N_4272,N_3071,N_2319);
and U4273 (N_4273,N_3185,N_3812);
xnor U4274 (N_4274,N_3272,N_2199);
and U4275 (N_4275,N_2031,N_3651);
nor U4276 (N_4276,N_2512,N_3718);
and U4277 (N_4277,N_2456,N_2807);
and U4278 (N_4278,N_3464,N_3973);
and U4279 (N_4279,N_3633,N_2482);
and U4280 (N_4280,N_3756,N_3907);
nor U4281 (N_4281,N_3515,N_2492);
xor U4282 (N_4282,N_3509,N_2474);
nand U4283 (N_4283,N_3266,N_2246);
or U4284 (N_4284,N_3838,N_3370);
and U4285 (N_4285,N_2919,N_2013);
nor U4286 (N_4286,N_3953,N_3995);
or U4287 (N_4287,N_2033,N_3189);
and U4288 (N_4288,N_2949,N_2207);
and U4289 (N_4289,N_3581,N_2719);
xor U4290 (N_4290,N_2379,N_2530);
xor U4291 (N_4291,N_2071,N_3532);
nand U4292 (N_4292,N_2646,N_3943);
nor U4293 (N_4293,N_3242,N_2987);
xnor U4294 (N_4294,N_2713,N_3994);
and U4295 (N_4295,N_3808,N_3880);
xnor U4296 (N_4296,N_2104,N_3116);
nor U4297 (N_4297,N_3111,N_3549);
nand U4298 (N_4298,N_3667,N_2268);
nand U4299 (N_4299,N_3417,N_3460);
or U4300 (N_4300,N_2229,N_2420);
xnor U4301 (N_4301,N_2176,N_2498);
and U4302 (N_4302,N_2472,N_3553);
or U4303 (N_4303,N_2590,N_3735);
nor U4304 (N_4304,N_2744,N_3885);
nand U4305 (N_4305,N_2965,N_3604);
nor U4306 (N_4306,N_3200,N_3741);
nor U4307 (N_4307,N_3032,N_3115);
xnor U4308 (N_4308,N_2201,N_2673);
and U4309 (N_4309,N_2654,N_2264);
nor U4310 (N_4310,N_2122,N_3580);
xor U4311 (N_4311,N_2587,N_3492);
nand U4312 (N_4312,N_2757,N_3785);
or U4313 (N_4313,N_2148,N_2153);
xnor U4314 (N_4314,N_3767,N_3289);
nand U4315 (N_4315,N_3625,N_2502);
xor U4316 (N_4316,N_2072,N_3984);
and U4317 (N_4317,N_3248,N_2934);
nor U4318 (N_4318,N_2611,N_2905);
xor U4319 (N_4319,N_3775,N_2171);
xor U4320 (N_4320,N_3269,N_2879);
nor U4321 (N_4321,N_3615,N_3376);
xor U4322 (N_4322,N_2209,N_3850);
and U4323 (N_4323,N_3062,N_3882);
nand U4324 (N_4324,N_2339,N_3466);
or U4325 (N_4325,N_3184,N_2032);
or U4326 (N_4326,N_3721,N_3086);
nor U4327 (N_4327,N_3146,N_2635);
xnor U4328 (N_4328,N_3930,N_3344);
and U4329 (N_4329,N_3367,N_3016);
and U4330 (N_4330,N_3873,N_3461);
nand U4331 (N_4331,N_3247,N_2257);
nor U4332 (N_4332,N_3738,N_2971);
xnor U4333 (N_4333,N_2723,N_3501);
xor U4334 (N_4334,N_2415,N_2515);
and U4335 (N_4335,N_2294,N_3766);
and U4336 (N_4336,N_3513,N_2720);
xnor U4337 (N_4337,N_3295,N_3987);
and U4338 (N_4338,N_2228,N_3249);
nand U4339 (N_4339,N_2640,N_2612);
xnor U4340 (N_4340,N_3495,N_3106);
nor U4341 (N_4341,N_3420,N_2904);
and U4342 (N_4342,N_3944,N_2951);
and U4343 (N_4343,N_3281,N_3592);
or U4344 (N_4344,N_2682,N_2615);
and U4345 (N_4345,N_3436,N_2299);
and U4346 (N_4346,N_3363,N_3918);
xor U4347 (N_4347,N_2163,N_3386);
or U4348 (N_4348,N_3989,N_2003);
and U4349 (N_4349,N_2901,N_2459);
xnor U4350 (N_4350,N_2963,N_3689);
xor U4351 (N_4351,N_2034,N_2302);
xor U4352 (N_4352,N_3128,N_3793);
xnor U4353 (N_4353,N_2857,N_2695);
nor U4354 (N_4354,N_2149,N_3954);
nand U4355 (N_4355,N_3471,N_3666);
and U4356 (N_4356,N_3967,N_3089);
and U4357 (N_4357,N_2195,N_2734);
xor U4358 (N_4358,N_2680,N_3707);
xnor U4359 (N_4359,N_2552,N_2475);
or U4360 (N_4360,N_2346,N_3095);
and U4361 (N_4361,N_3387,N_3313);
or U4362 (N_4362,N_2585,N_3042);
and U4363 (N_4363,N_3576,N_3530);
nor U4364 (N_4364,N_3220,N_2745);
nor U4365 (N_4365,N_3443,N_2430);
nor U4366 (N_4366,N_3815,N_3704);
xnor U4367 (N_4367,N_3419,N_2884);
and U4368 (N_4368,N_3159,N_2183);
nand U4369 (N_4369,N_2670,N_3842);
or U4370 (N_4370,N_2898,N_2012);
xnor U4371 (N_4371,N_3164,N_3992);
nor U4372 (N_4372,N_3170,N_3679);
or U4373 (N_4373,N_2864,N_3802);
xnor U4374 (N_4374,N_2375,N_2049);
nand U4375 (N_4375,N_3618,N_2463);
and U4376 (N_4376,N_3925,N_3871);
nor U4377 (N_4377,N_2036,N_2337);
nand U4378 (N_4378,N_3818,N_2551);
xor U4379 (N_4379,N_2737,N_3854);
or U4380 (N_4380,N_2418,N_3142);
and U4381 (N_4381,N_3375,N_3305);
nand U4382 (N_4382,N_2070,N_2413);
nand U4383 (N_4383,N_2307,N_3763);
or U4384 (N_4384,N_2191,N_2296);
nand U4385 (N_4385,N_3010,N_3770);
xnor U4386 (N_4386,N_2325,N_3267);
or U4387 (N_4387,N_2067,N_2406);
xor U4388 (N_4388,N_3942,N_3398);
xnor U4389 (N_4389,N_2503,N_2162);
nand U4390 (N_4390,N_2305,N_2091);
nor U4391 (N_4391,N_3575,N_2714);
nor U4392 (N_4392,N_3757,N_2599);
nor U4393 (N_4393,N_2279,N_3270);
xnor U4394 (N_4394,N_2014,N_3105);
nor U4395 (N_4395,N_2982,N_2787);
or U4396 (N_4396,N_2112,N_2332);
and U4397 (N_4397,N_3025,N_3927);
nand U4398 (N_4398,N_3632,N_3970);
nor U4399 (N_4399,N_3601,N_3463);
nor U4400 (N_4400,N_3020,N_2579);
xnor U4401 (N_4401,N_2429,N_2397);
nand U4402 (N_4402,N_2243,N_3005);
nor U4403 (N_4403,N_2835,N_2290);
nor U4404 (N_4404,N_3516,N_3311);
nor U4405 (N_4405,N_2976,N_2443);
or U4406 (N_4406,N_3488,N_3175);
or U4407 (N_4407,N_3577,N_2204);
or U4408 (N_4408,N_2666,N_3286);
or U4409 (N_4409,N_2873,N_2361);
nand U4410 (N_4410,N_2993,N_3265);
xnor U4411 (N_4411,N_2991,N_2212);
and U4412 (N_4412,N_3196,N_3215);
nand U4413 (N_4413,N_3561,N_3701);
nor U4414 (N_4414,N_3777,N_3043);
or U4415 (N_4415,N_3957,N_2862);
or U4416 (N_4416,N_3727,N_3225);
nand U4417 (N_4417,N_3685,N_2399);
nor U4418 (N_4418,N_3012,N_3291);
or U4419 (N_4419,N_3993,N_3645);
nand U4420 (N_4420,N_3301,N_2620);
nand U4421 (N_4421,N_3600,N_3769);
or U4422 (N_4422,N_3259,N_3780);
and U4423 (N_4423,N_2840,N_2808);
nand U4424 (N_4424,N_3083,N_2056);
and U4425 (N_4425,N_2224,N_2546);
nor U4426 (N_4426,N_3404,N_2335);
or U4427 (N_4427,N_2878,N_3747);
or U4428 (N_4428,N_3110,N_2675);
or U4429 (N_4429,N_3399,N_3227);
and U4430 (N_4430,N_2329,N_2481);
nand U4431 (N_4431,N_2794,N_3643);
or U4432 (N_4432,N_2370,N_3817);
xnor U4433 (N_4433,N_3183,N_2945);
xnor U4434 (N_4434,N_3383,N_2124);
and U4435 (N_4435,N_2926,N_3748);
nand U4436 (N_4436,N_3090,N_3899);
nand U4437 (N_4437,N_3391,N_2568);
or U4438 (N_4438,N_2175,N_2101);
nor U4439 (N_4439,N_2921,N_3396);
or U4440 (N_4440,N_2900,N_3423);
or U4441 (N_4441,N_2016,N_2916);
and U4442 (N_4442,N_3437,N_3734);
nor U4443 (N_4443,N_2460,N_3004);
nor U4444 (N_4444,N_2240,N_2051);
and U4445 (N_4445,N_3486,N_2769);
or U4446 (N_4446,N_2690,N_2883);
xnor U4447 (N_4447,N_2065,N_3595);
nor U4448 (N_4448,N_2373,N_2323);
and U4449 (N_4449,N_2077,N_3567);
and U4450 (N_4450,N_3308,N_3675);
nor U4451 (N_4451,N_2721,N_3776);
xor U4452 (N_4452,N_2961,N_2117);
or U4453 (N_4453,N_3320,N_3795);
nand U4454 (N_4454,N_2943,N_3681);
or U4455 (N_4455,N_3258,N_2935);
and U4456 (N_4456,N_2297,N_2657);
or U4457 (N_4457,N_2914,N_3079);
and U4458 (N_4458,N_2774,N_3397);
nor U4459 (N_4459,N_3810,N_2094);
or U4460 (N_4460,N_2200,N_3329);
and U4461 (N_4461,N_2778,N_2603);
or U4462 (N_4462,N_2285,N_2487);
nor U4463 (N_4463,N_3027,N_2132);
xor U4464 (N_4464,N_2001,N_2291);
nor U4465 (N_4465,N_3093,N_3161);
or U4466 (N_4466,N_2068,N_2606);
xor U4467 (N_4467,N_2613,N_2119);
and U4468 (N_4468,N_2631,N_3055);
and U4469 (N_4469,N_3058,N_2868);
nor U4470 (N_4470,N_2321,N_3191);
xor U4471 (N_4471,N_2435,N_3977);
nand U4472 (N_4472,N_2701,N_2589);
nor U4473 (N_4473,N_3849,N_3733);
nand U4474 (N_4474,N_3034,N_2417);
xor U4475 (N_4475,N_3306,N_2694);
xor U4476 (N_4476,N_2454,N_3739);
or U4477 (N_4477,N_2168,N_2954);
or U4478 (N_4478,N_3368,N_3351);
nor U4479 (N_4479,N_2473,N_3237);
xor U4480 (N_4480,N_2095,N_3366);
xor U4481 (N_4481,N_2387,N_3531);
and U4482 (N_4482,N_3331,N_3543);
nand U4483 (N_4483,N_2565,N_2252);
nor U4484 (N_4484,N_3822,N_3364);
nand U4485 (N_4485,N_3640,N_2785);
or U4486 (N_4486,N_2662,N_2630);
xor U4487 (N_4487,N_3546,N_3400);
or U4488 (N_4488,N_2910,N_2000);
or U4489 (N_4489,N_2352,N_2877);
nand U4490 (N_4490,N_2439,N_2977);
xor U4491 (N_4491,N_3328,N_3314);
nand U4492 (N_4492,N_2591,N_3359);
or U4493 (N_4493,N_2385,N_2082);
or U4494 (N_4494,N_3883,N_2249);
xnor U4495 (N_4495,N_3834,N_2780);
nor U4496 (N_4496,N_2793,N_3477);
nor U4497 (N_4497,N_3491,N_3627);
xor U4498 (N_4498,N_3104,N_2762);
and U4499 (N_4499,N_3354,N_2401);
nor U4500 (N_4500,N_3121,N_2927);
nand U4501 (N_4501,N_2556,N_2477);
xor U4502 (N_4502,N_3192,N_2891);
xor U4503 (N_4503,N_3402,N_2047);
nor U4504 (N_4504,N_2392,N_3392);
or U4505 (N_4505,N_2407,N_3348);
and U4506 (N_4506,N_3063,N_3337);
or U4507 (N_4507,N_2709,N_3535);
nor U4508 (N_4508,N_2773,N_3597);
xor U4509 (N_4509,N_2127,N_3049);
nand U4510 (N_4510,N_3029,N_3156);
nor U4511 (N_4511,N_3202,N_3746);
xnor U4512 (N_4512,N_2295,N_2099);
xor U4513 (N_4513,N_3065,N_3628);
and U4514 (N_4514,N_3141,N_2950);
and U4515 (N_4515,N_3230,N_2371);
or U4516 (N_4516,N_2960,N_2968);
nand U4517 (N_4517,N_3536,N_3635);
nor U4518 (N_4518,N_2235,N_3619);
xor U4519 (N_4519,N_3759,N_3123);
or U4520 (N_4520,N_3534,N_3414);
xnor U4521 (N_4521,N_2595,N_2677);
or U4522 (N_4522,N_3832,N_3136);
and U4523 (N_4523,N_2545,N_3614);
and U4524 (N_4524,N_3642,N_2799);
xor U4525 (N_4525,N_2214,N_2880);
nand U4526 (N_4526,N_2241,N_2315);
nand U4527 (N_4527,N_2665,N_2262);
nand U4528 (N_4528,N_2416,N_2458);
or U4529 (N_4529,N_2700,N_2917);
and U4530 (N_4530,N_3341,N_2303);
nand U4531 (N_4531,N_3194,N_3665);
xor U4532 (N_4532,N_2018,N_2308);
and U4533 (N_4533,N_2327,N_3609);
and U4534 (N_4534,N_2093,N_2453);
xnor U4535 (N_4535,N_2717,N_3988);
nor U4536 (N_4536,N_2222,N_2739);
nand U4537 (N_4537,N_2758,N_3287);
or U4538 (N_4538,N_3590,N_3319);
nand U4539 (N_4539,N_3087,N_3074);
and U4540 (N_4540,N_2261,N_3454);
xor U4541 (N_4541,N_3467,N_3422);
and U4542 (N_4542,N_2889,N_3040);
xnor U4543 (N_4543,N_2957,N_3890);
nor U4544 (N_4544,N_3965,N_3444);
nor U4545 (N_4545,N_3213,N_2783);
or U4546 (N_4546,N_3362,N_2363);
xnor U4547 (N_4547,N_2983,N_3373);
nor U4548 (N_4548,N_3935,N_3919);
and U4549 (N_4549,N_3442,N_3700);
nand U4550 (N_4550,N_3845,N_2496);
nor U4551 (N_4551,N_2726,N_3937);
and U4552 (N_4552,N_2686,N_2211);
and U4553 (N_4553,N_3059,N_2433);
and U4554 (N_4554,N_3282,N_3564);
and U4555 (N_4555,N_2782,N_2140);
nand U4556 (N_4556,N_3275,N_2679);
nand U4557 (N_4557,N_3036,N_3978);
or U4558 (N_4558,N_3228,N_2287);
nand U4559 (N_4559,N_2698,N_3745);
xnor U4560 (N_4560,N_2989,N_2839);
and U4561 (N_4561,N_2522,N_3496);
xor U4562 (N_4562,N_2554,N_3570);
nor U4563 (N_4563,N_3254,N_2015);
xor U4564 (N_4564,N_3133,N_3073);
nand U4565 (N_4565,N_3788,N_3550);
nor U4566 (N_4566,N_3377,N_3151);
xnor U4567 (N_4567,N_3449,N_3221);
and U4568 (N_4568,N_3897,N_3826);
nand U4569 (N_4569,N_2028,N_3621);
and U4570 (N_4570,N_3968,N_3860);
nand U4571 (N_4571,N_3938,N_3506);
xnor U4572 (N_4572,N_2011,N_3198);
nand U4573 (N_4573,N_2027,N_3418);
or U4574 (N_4574,N_3246,N_2063);
nor U4575 (N_4575,N_3139,N_3335);
nand U4576 (N_4576,N_2656,N_2928);
nor U4577 (N_4577,N_2796,N_3933);
nand U4578 (N_4578,N_2668,N_2791);
nor U4579 (N_4579,N_3712,N_3395);
and U4580 (N_4580,N_3668,N_2223);
nand U4581 (N_4581,N_3369,N_3327);
nor U4582 (N_4582,N_2766,N_3545);
xnor U4583 (N_4583,N_2449,N_3514);
xnor U4584 (N_4584,N_2078,N_2759);
and U4585 (N_4585,N_2810,N_2622);
and U4586 (N_4586,N_3130,N_3051);
xnor U4587 (N_4587,N_3742,N_2692);
or U4588 (N_4588,N_2217,N_3187);
nor U4589 (N_4589,N_2431,N_2828);
nor U4590 (N_4590,N_2105,N_3256);
nand U4591 (N_4591,N_2083,N_3637);
nor U4592 (N_4592,N_2999,N_3551);
nor U4593 (N_4593,N_2272,N_3568);
nor U4594 (N_4594,N_2025,N_3905);
xor U4595 (N_4595,N_3283,N_3479);
or U4596 (N_4596,N_2374,N_2107);
xor U4597 (N_4597,N_3132,N_3061);
nand U4598 (N_4598,N_2098,N_3431);
xor U4599 (N_4599,N_3582,N_2150);
or U4600 (N_4600,N_2894,N_3623);
and U4601 (N_4601,N_3884,N_3629);
nand U4602 (N_4602,N_3468,N_2529);
nor U4603 (N_4603,N_2756,N_2347);
or U4604 (N_4604,N_2532,N_3217);
xor U4605 (N_4605,N_3333,N_3657);
and U4606 (N_4606,N_2269,N_2776);
and U4607 (N_4607,N_3177,N_2746);
or U4608 (N_4608,N_3109,N_2230);
nor U4609 (N_4609,N_2892,N_2995);
xor U4610 (N_4610,N_3389,N_2088);
nand U4611 (N_4611,N_3533,N_3124);
or U4612 (N_4612,N_3527,N_2882);
and U4613 (N_4613,N_3360,N_2814);
or U4614 (N_4614,N_3394,N_3999);
nor U4615 (N_4615,N_2152,N_2586);
xnor U4616 (N_4616,N_2871,N_3475);
nand U4617 (N_4617,N_2116,N_3749);
nor U4618 (N_4618,N_2372,N_2253);
xor U4619 (N_4619,N_2286,N_3160);
nand U4620 (N_4620,N_2718,N_2096);
and U4621 (N_4621,N_3782,N_2967);
nor U4622 (N_4622,N_2572,N_3014);
and U4623 (N_4623,N_2789,N_2649);
or U4624 (N_4624,N_3955,N_3101);
xor U4625 (N_4625,N_2899,N_3098);
or U4626 (N_4626,N_3162,N_2958);
nor U4627 (N_4627,N_3346,N_2501);
xor U4628 (N_4628,N_2039,N_3209);
nor U4629 (N_4629,N_3888,N_3129);
xor U4630 (N_4630,N_2761,N_3438);
or U4631 (N_4631,N_3031,N_3961);
or U4632 (N_4632,N_3726,N_3606);
nor U4633 (N_4633,N_2550,N_2738);
nor U4634 (N_4634,N_3906,N_2362);
and U4635 (N_4635,N_2333,N_2854);
and U4636 (N_4636,N_2444,N_3869);
and U4637 (N_4637,N_3297,N_3626);
xnor U4638 (N_4638,N_2306,N_3508);
nor U4639 (N_4639,N_3253,N_2931);
and U4640 (N_4640,N_3608,N_2994);
and U4641 (N_4641,N_3315,N_3276);
xor U4642 (N_4642,N_3800,N_2575);
nand U4643 (N_4643,N_3309,N_3257);
nand U4644 (N_4644,N_2540,N_2102);
and U4645 (N_4645,N_2021,N_3007);
and U4646 (N_4646,N_3138,N_2952);
or U4647 (N_4647,N_2289,N_3980);
nor U4648 (N_4648,N_2400,N_3781);
nor U4649 (N_4649,N_2193,N_2237);
xnor U4650 (N_4650,N_3837,N_2388);
and U4651 (N_4651,N_2258,N_3610);
nor U4652 (N_4652,N_3193,N_2074);
or U4653 (N_4653,N_3974,N_3067);
nand U4654 (N_4654,N_2389,N_2781);
nand U4655 (N_4655,N_3786,N_3338);
xnor U4656 (N_4656,N_3274,N_3046);
xor U4657 (N_4657,N_2398,N_2790);
and U4658 (N_4658,N_3909,N_3240);
nor U4659 (N_4659,N_2422,N_3470);
nor U4660 (N_4660,N_3245,N_2427);
nand U4661 (N_4661,N_2114,N_3154);
xor U4662 (N_4662,N_3140,N_2621);
nor U4663 (N_4663,N_3052,N_3410);
nor U4664 (N_4664,N_3273,N_3135);
nand U4665 (N_4665,N_2377,N_2349);
nand U4666 (N_4666,N_3696,N_3493);
or U4667 (N_4667,N_3695,N_2275);
xnor U4668 (N_4668,N_2395,N_2600);
and U4669 (N_4669,N_2161,N_2242);
nand U4670 (N_4670,N_2970,N_3502);
or U4671 (N_4671,N_2005,N_2831);
xor U4672 (N_4672,N_2535,N_2650);
nand U4673 (N_4673,N_2707,N_3772);
nand U4674 (N_4674,N_2485,N_2218);
and U4675 (N_4675,N_3385,N_3407);
nand U4676 (N_4676,N_2753,N_2915);
nor U4677 (N_4677,N_3846,N_2231);
nand U4678 (N_4678,N_3829,N_3484);
or U4679 (N_4679,N_2804,N_2020);
xor U4680 (N_4680,N_2245,N_2770);
nand U4681 (N_4681,N_3411,N_3388);
xor U4682 (N_4682,N_2182,N_3011);
or U4683 (N_4683,N_3299,N_2085);
or U4684 (N_4684,N_3057,N_2732);
nand U4685 (N_4685,N_2158,N_3683);
or U4686 (N_4686,N_2816,N_2897);
nand U4687 (N_4687,N_2386,N_2383);
nand U4688 (N_4688,N_2661,N_3229);
nand U4689 (N_4689,N_3694,N_2942);
xor U4690 (N_4690,N_3081,N_3378);
nand U4691 (N_4691,N_3920,N_2247);
or U4692 (N_4692,N_2437,N_3412);
nor U4693 (N_4693,N_3537,N_2432);
or U4694 (N_4694,N_3462,N_2623);
or U4695 (N_4695,N_2507,N_2499);
xnor U4696 (N_4696,N_3660,N_3851);
or U4697 (N_4697,N_2062,N_3205);
nand U4698 (N_4698,N_2471,N_3238);
xor U4699 (N_4699,N_2317,N_2577);
nor U4700 (N_4700,N_3929,N_2890);
xnor U4701 (N_4701,N_3616,N_2652);
or U4702 (N_4702,N_3891,N_3820);
nor U4703 (N_4703,N_3045,N_3445);
nand U4704 (N_4704,N_2988,N_3428);
nand U4705 (N_4705,N_3456,N_3122);
xor U4706 (N_4706,N_3874,N_2521);
nand U4707 (N_4707,N_2173,N_3134);
or U4708 (N_4708,N_2933,N_3881);
nor U4709 (N_4709,N_2913,N_3082);
nor U4710 (N_4710,N_3706,N_3612);
or U4711 (N_4711,N_2390,N_3494);
xnor U4712 (N_4712,N_3520,N_2578);
or U4713 (N_4713,N_3806,N_3538);
nand U4714 (N_4714,N_3409,N_3578);
or U4715 (N_4715,N_3722,N_3163);
nand U4716 (N_4716,N_2768,N_3003);
nor U4717 (N_4717,N_3799,N_3887);
nor U4718 (N_4718,N_3998,N_3244);
nor U4719 (N_4719,N_2797,N_2625);
xnor U4720 (N_4720,N_2256,N_2438);
nor U4721 (N_4721,N_2978,N_3687);
and U4722 (N_4722,N_2980,N_3624);
nand U4723 (N_4723,N_3324,N_3949);
nand U4724 (N_4724,N_2874,N_3569);
and U4725 (N_4725,N_3434,N_2210);
and U4726 (N_4726,N_3894,N_2909);
nor U4727 (N_4727,N_3510,N_3563);
nand U4728 (N_4728,N_2775,N_2843);
xor U4729 (N_4729,N_2135,N_2531);
and U4730 (N_4730,N_2451,N_2902);
or U4731 (N_4731,N_2815,N_2066);
or U4732 (N_4732,N_2616,N_2947);
and U4733 (N_4733,N_3650,N_2996);
nor U4734 (N_4734,N_2852,N_3779);
nand U4735 (N_4735,N_3379,N_2979);
or U4736 (N_4736,N_3457,N_3382);
and U4737 (N_4737,N_3653,N_3103);
xor U4738 (N_4738,N_2185,N_2547);
nand U4739 (N_4739,N_3825,N_3268);
nand U4740 (N_4740,N_2594,N_2583);
nor U4741 (N_4741,N_3878,N_3525);
nor U4742 (N_4742,N_3620,N_3821);
nand U4743 (N_4743,N_3068,N_2549);
and U4744 (N_4744,N_3120,N_2517);
and U4745 (N_4745,N_2667,N_3208);
and U4746 (N_4746,N_2312,N_3877);
nor U4747 (N_4747,N_3284,N_3711);
and U4748 (N_4748,N_2186,N_2861);
and U4749 (N_4749,N_3648,N_2524);
and U4750 (N_4750,N_2233,N_2538);
and U4751 (N_4751,N_2139,N_2184);
xnor U4752 (N_4752,N_3204,N_3677);
xor U4753 (N_4753,N_3261,N_2137);
nor U4754 (N_4754,N_3895,N_3839);
nand U4755 (N_4755,N_2742,N_2805);
xor U4756 (N_4756,N_3114,N_3517);
xnor U4757 (N_4757,N_2216,N_3203);
or U4758 (N_4758,N_3452,N_2320);
and U4759 (N_4759,N_3356,N_2801);
and U4760 (N_4760,N_3588,N_3478);
xnor U4761 (N_4761,N_3127,N_2664);
or U4762 (N_4762,N_2125,N_2330);
or U4763 (N_4763,N_3241,N_3948);
and U4764 (N_4764,N_3720,N_3950);
and U4765 (N_4765,N_3662,N_2911);
xor U4766 (N_4766,N_3102,N_3236);
xnor U4767 (N_4767,N_2806,N_3298);
nand U4768 (N_4768,N_3558,N_2618);
nor U4769 (N_4769,N_2356,N_3330);
xnor U4770 (N_4770,N_3339,N_2813);
or U4771 (N_4771,N_3023,N_3898);
and U4772 (N_4772,N_3173,N_3374);
nor U4773 (N_4773,N_2648,N_3522);
nor U4774 (N_4774,N_2735,N_2514);
or U4775 (N_4775,N_2143,N_3819);
xnor U4776 (N_4776,N_2225,N_3343);
xnor U4777 (N_4777,N_3613,N_3638);
and U4778 (N_4778,N_3037,N_2426);
and U4779 (N_4779,N_2881,N_3831);
or U4780 (N_4780,N_2573,N_2519);
nand U4781 (N_4781,N_2309,N_3611);
and U4782 (N_4782,N_2895,N_3511);
and U4783 (N_4783,N_2055,N_3097);
xor U4784 (N_4784,N_3519,N_2722);
nor U4785 (N_4785,N_2634,N_2755);
or U4786 (N_4786,N_3617,N_3827);
xnor U4787 (N_4787,N_2955,N_2925);
nand U4788 (N_4788,N_2624,N_2946);
nand U4789 (N_4789,N_2053,N_3446);
or U4790 (N_4790,N_2343,N_2113);
nand U4791 (N_4791,N_3174,N_3499);
nand U4792 (N_4792,N_3958,N_3743);
nor U4793 (N_4793,N_2494,N_3981);
xor U4794 (N_4794,N_2689,N_3814);
and U4795 (N_4795,N_3483,N_2076);
xor U4796 (N_4796,N_2334,N_2663);
nand U4797 (N_4797,N_3796,N_2821);
nor U4798 (N_4798,N_3674,N_2324);
xor U4799 (N_4799,N_2936,N_2580);
xor U4800 (N_4800,N_3318,N_3131);
nor U4801 (N_4801,N_3503,N_2189);
nor U4802 (N_4802,N_2467,N_3168);
nand U4803 (N_4803,N_2351,N_2636);
xnor U4804 (N_4804,N_2026,N_3589);
or U4805 (N_4805,N_3816,N_3682);
and U4806 (N_4806,N_3809,N_3991);
and U4807 (N_4807,N_3691,N_3390);
nor U4808 (N_4808,N_2486,N_2038);
and U4809 (N_4809,N_3279,N_2470);
and U4810 (N_4810,N_2080,N_3179);
nor U4811 (N_4811,N_2358,N_3824);
nand U4812 (N_4812,N_2672,N_2409);
xor U4813 (N_4813,N_2178,N_2301);
nand U4814 (N_4814,N_3421,N_2609);
or U4815 (N_4815,N_2893,N_2366);
nand U4816 (N_4816,N_3201,N_3789);
nor U4817 (N_4817,N_3199,N_2975);
nand U4818 (N_4818,N_2219,N_2748);
nand U4819 (N_4819,N_2903,N_3622);
nor U4820 (N_4820,N_2166,N_2571);
and U4821 (N_4821,N_2326,N_3001);
nor U4822 (N_4822,N_2953,N_3172);
nand U4823 (N_4823,N_2533,N_3223);
xnor U4824 (N_4824,N_2239,N_2344);
nand U4825 (N_4825,N_3252,N_3997);
nand U4826 (N_4826,N_2408,N_2497);
or U4827 (N_4827,N_3100,N_2029);
and U4828 (N_4828,N_3902,N_2002);
nor U4829 (N_4829,N_3840,N_3017);
nor U4830 (N_4830,N_3408,N_3541);
and U4831 (N_4831,N_3171,N_2865);
and U4832 (N_4832,N_3876,N_3294);
xor U4833 (N_4833,N_3041,N_3699);
or U4834 (N_4834,N_2405,N_3731);
xor U4835 (N_4835,N_2973,N_2990);
nor U4836 (N_4836,N_2711,N_2860);
or U4837 (N_4837,N_2350,N_2544);
and U4838 (N_4838,N_2788,N_2328);
nand U4839 (N_4839,N_3893,N_3889);
nand U4840 (N_4840,N_2555,N_2830);
nor U4841 (N_4841,N_3602,N_3661);
xor U4842 (N_4842,N_2154,N_3487);
or U4843 (N_4843,N_2912,N_2145);
nor U4844 (N_4844,N_2354,N_3754);
and U4845 (N_4845,N_3848,N_3996);
nand U4846 (N_4846,N_3853,N_2322);
and U4847 (N_4847,N_2238,N_3262);
xor U4848 (N_4848,N_2985,N_3729);
nor U4849 (N_4849,N_2359,N_3934);
and U4850 (N_4850,N_3728,N_3044);
or U4851 (N_4851,N_2221,N_3959);
or U4852 (N_4852,N_3835,N_3926);
and U4853 (N_4853,N_2108,N_3064);
nand U4854 (N_4854,N_2491,N_2986);
or U4855 (N_4855,N_3278,N_2743);
and U4856 (N_4856,N_3054,N_3910);
nand U4857 (N_4857,N_3596,N_3708);
xor U4858 (N_4858,N_2526,N_2079);
and U4859 (N_4859,N_3585,N_3500);
and U4860 (N_4860,N_2440,N_3705);
xor U4861 (N_4861,N_2607,N_2760);
nand U4862 (N_4862,N_2706,N_2006);
xor U4863 (N_4863,N_2598,N_3349);
nand U4864 (N_4864,N_2226,N_2266);
or U4865 (N_4865,N_2605,N_2896);
xor U4866 (N_4866,N_2751,N_3591);
nand U4867 (N_4867,N_2823,N_3481);
nand U4868 (N_4868,N_2944,N_2696);
nor U4869 (N_4869,N_2022,N_2500);
nand U4870 (N_4870,N_3521,N_3639);
xnor U4871 (N_4871,N_2425,N_2194);
or U4872 (N_4872,N_2284,N_3870);
nand U4873 (N_4873,N_3118,N_3859);
nor U4874 (N_4874,N_2314,N_3033);
xnor U4875 (N_4875,N_3070,N_3908);
nand U4876 (N_4876,N_3214,N_3807);
nor U4877 (N_4877,N_2923,N_3603);
and U4878 (N_4878,N_3983,N_2566);
and U4879 (N_4879,N_2747,N_3340);
and U4880 (N_4880,N_3924,N_2213);
xor U4881 (N_4881,N_2123,N_3345);
nand U4882 (N_4882,N_3847,N_3080);
nand U4883 (N_4883,N_2704,N_2466);
nand U4884 (N_4884,N_3764,N_2932);
xnor U4885 (N_4885,N_3504,N_2007);
nor U4886 (N_4886,N_3664,N_2215);
and U4887 (N_4887,N_3680,N_2887);
and U4888 (N_4888,N_2886,N_3962);
or U4889 (N_4889,N_2593,N_2800);
nand U4890 (N_4890,N_3913,N_3212);
or U4891 (N_4891,N_3182,N_3350);
or U4892 (N_4892,N_2792,N_2629);
and U4893 (N_4893,N_2525,N_3804);
nand U4894 (N_4894,N_3655,N_3915);
xnor U4895 (N_4895,N_2653,N_2715);
or U4896 (N_4896,N_3465,N_3117);
and U4897 (N_4897,N_2423,N_2708);
nand U4898 (N_4898,N_2402,N_3069);
and U4899 (N_4899,N_2403,N_3903);
nand U4900 (N_4900,N_2729,N_3523);
and U4901 (N_4901,N_2867,N_2969);
or U4902 (N_4902,N_2045,N_2763);
and U4903 (N_4903,N_2452,N_3526);
xnor U4904 (N_4904,N_3556,N_3024);
xor U4905 (N_4905,N_2436,N_2087);
and U4906 (N_4906,N_3932,N_2849);
nor U4907 (N_4907,N_2164,N_3147);
or U4908 (N_4908,N_3966,N_2504);
and U4909 (N_4909,N_2826,N_2588);
nor U4910 (N_4910,N_2767,N_3586);
or U4911 (N_4911,N_3206,N_3644);
xnor U4912 (N_4912,N_2367,N_2469);
and U4913 (N_4913,N_3512,N_3572);
or U4914 (N_4914,N_2244,N_3008);
xnor U4915 (N_4915,N_3293,N_3573);
nor U4916 (N_4916,N_2697,N_2655);
xor U4917 (N_4917,N_3235,N_2084);
nor U4918 (N_4918,N_3322,N_2380);
nor U4919 (N_4919,N_2177,N_2853);
and U4920 (N_4920,N_3921,N_3458);
xor U4921 (N_4921,N_3861,N_3836);
xor U4922 (N_4922,N_2265,N_3862);
nand U4923 (N_4923,N_2817,N_3979);
or U4924 (N_4924,N_3875,N_2998);
nand U4925 (N_4925,N_2829,N_3656);
and U4926 (N_4926,N_2198,N_3232);
nor U4927 (N_4927,N_2160,N_3013);
nand U4928 (N_4928,N_3365,N_3752);
nor U4929 (N_4929,N_2236,N_3239);
nor U4930 (N_4930,N_3736,N_3762);
or U4931 (N_4931,N_2863,N_3646);
nand U4932 (N_4932,N_2939,N_2846);
xor U4933 (N_4933,N_3939,N_3153);
xor U4934 (N_4934,N_2592,N_2048);
nand U4935 (N_4935,N_2699,N_2728);
nor U4936 (N_4936,N_2129,N_2858);
xnor U4937 (N_4937,N_3940,N_2434);
nand U4938 (N_4938,N_2090,N_3157);
and U4939 (N_4939,N_3917,N_2639);
xor U4940 (N_4940,N_3579,N_3555);
xnor U4941 (N_4941,N_3432,N_2260);
and U4942 (N_4942,N_2518,N_3856);
or U4943 (N_4943,N_3636,N_2687);
or U4944 (N_4944,N_2348,N_2259);
nand U4945 (N_4945,N_3852,N_3922);
or U4946 (N_4946,N_2250,N_2772);
and U4947 (N_4947,N_2559,N_3823);
nand U4948 (N_4948,N_2267,N_3323);
or U4949 (N_4949,N_2304,N_2197);
or U4950 (N_4950,N_2818,N_2930);
xor U4951 (N_4951,N_3717,N_3210);
xor U4952 (N_4952,N_3584,N_3112);
nand U4953 (N_4953,N_2190,N_3195);
nor U4954 (N_4954,N_3797,N_2562);
nand U4955 (N_4955,N_2368,N_3912);
nor U4956 (N_4956,N_2798,N_2956);
xor U4957 (N_4957,N_3986,N_2462);
xor U4958 (N_4958,N_3911,N_3833);
xnor U4959 (N_4959,N_3678,N_2604);
nor U4960 (N_4960,N_2561,N_2490);
nor U4961 (N_4961,N_2187,N_3844);
nor U4962 (N_4962,N_3381,N_2357);
or U4963 (N_4963,N_2981,N_2282);
xor U4964 (N_4964,N_2414,N_2764);
or U4965 (N_4965,N_3803,N_2292);
nor U4966 (N_4966,N_2455,N_2248);
nand U4967 (N_4967,N_3096,N_3830);
nand U4968 (N_4968,N_2924,N_2441);
nand U4969 (N_4969,N_3002,N_3312);
nor U4970 (N_4970,N_2364,N_3347);
xnor U4971 (N_4971,N_2255,N_2412);
xor U4972 (N_4972,N_3976,N_3896);
and U4973 (N_4973,N_3811,N_3371);
nand U4974 (N_4974,N_2133,N_3904);
nand U4975 (N_4975,N_3447,N_3631);
xnor U4976 (N_4976,N_2644,N_2750);
and U4977 (N_4977,N_2396,N_3009);
nand U4978 (N_4978,N_2156,N_2702);
or U4979 (N_4979,N_3440,N_3548);
or U4980 (N_4980,N_3528,N_3280);
and U4981 (N_4981,N_2632,N_3427);
xor U4982 (N_4982,N_2288,N_3332);
nor U4983 (N_4983,N_2560,N_2779);
or U4984 (N_4984,N_2179,N_3791);
or U4985 (N_4985,N_2584,N_3137);
nor U4986 (N_4986,N_2196,N_2564);
nand U4987 (N_4987,N_3413,N_3358);
xnor U4988 (N_4988,N_3038,N_2984);
nand U4989 (N_4989,N_2251,N_3684);
and U4990 (N_4990,N_3787,N_2567);
nor U4991 (N_4991,N_2318,N_2442);
nand U4992 (N_4992,N_3302,N_3673);
nor U4993 (N_4993,N_2557,N_2888);
nor U4994 (N_4994,N_2513,N_3560);
nor U4995 (N_4995,N_2391,N_2676);
xnor U4996 (N_4996,N_2940,N_2167);
nor U4997 (N_4997,N_2693,N_3026);
nand U4998 (N_4998,N_3693,N_2476);
xnor U4999 (N_4999,N_3956,N_2845);
nand U5000 (N_5000,N_2637,N_3174);
nor U5001 (N_5001,N_3854,N_2839);
xnor U5002 (N_5002,N_3571,N_3765);
and U5003 (N_5003,N_2423,N_3716);
xor U5004 (N_5004,N_3929,N_3379);
xnor U5005 (N_5005,N_2481,N_3945);
or U5006 (N_5006,N_3024,N_3494);
xor U5007 (N_5007,N_3494,N_2389);
xnor U5008 (N_5008,N_2251,N_2712);
and U5009 (N_5009,N_3399,N_2843);
xor U5010 (N_5010,N_3755,N_3320);
or U5011 (N_5011,N_2615,N_3770);
nand U5012 (N_5012,N_3014,N_3012);
and U5013 (N_5013,N_3950,N_3761);
nor U5014 (N_5014,N_2116,N_3797);
nand U5015 (N_5015,N_2673,N_3575);
nand U5016 (N_5016,N_3922,N_3251);
nor U5017 (N_5017,N_2418,N_2397);
and U5018 (N_5018,N_3462,N_2723);
or U5019 (N_5019,N_3494,N_3625);
xnor U5020 (N_5020,N_2282,N_2547);
or U5021 (N_5021,N_3096,N_3941);
and U5022 (N_5022,N_3301,N_3396);
and U5023 (N_5023,N_3458,N_2051);
xor U5024 (N_5024,N_2718,N_2519);
or U5025 (N_5025,N_2032,N_3759);
xnor U5026 (N_5026,N_3576,N_3626);
nand U5027 (N_5027,N_2697,N_3896);
nor U5028 (N_5028,N_3567,N_2869);
nand U5029 (N_5029,N_3735,N_3552);
and U5030 (N_5030,N_2169,N_3548);
and U5031 (N_5031,N_3607,N_3907);
xnor U5032 (N_5032,N_3432,N_2366);
nor U5033 (N_5033,N_2152,N_2659);
or U5034 (N_5034,N_2876,N_3580);
xor U5035 (N_5035,N_2583,N_3079);
or U5036 (N_5036,N_3657,N_3699);
nor U5037 (N_5037,N_3384,N_2897);
or U5038 (N_5038,N_3527,N_2793);
and U5039 (N_5039,N_2063,N_2930);
and U5040 (N_5040,N_3817,N_3796);
nand U5041 (N_5041,N_2518,N_3173);
nor U5042 (N_5042,N_2721,N_3910);
nor U5043 (N_5043,N_3414,N_2076);
nand U5044 (N_5044,N_3145,N_3020);
and U5045 (N_5045,N_2841,N_3532);
nor U5046 (N_5046,N_2036,N_3944);
nor U5047 (N_5047,N_3065,N_2817);
and U5048 (N_5048,N_2221,N_3542);
and U5049 (N_5049,N_3251,N_3712);
xnor U5050 (N_5050,N_2304,N_3452);
or U5051 (N_5051,N_2691,N_3675);
nand U5052 (N_5052,N_2599,N_3033);
nand U5053 (N_5053,N_2158,N_3739);
or U5054 (N_5054,N_3477,N_3791);
or U5055 (N_5055,N_3893,N_3477);
nand U5056 (N_5056,N_3288,N_2437);
nand U5057 (N_5057,N_3642,N_3137);
xnor U5058 (N_5058,N_2266,N_3878);
nand U5059 (N_5059,N_2690,N_2509);
or U5060 (N_5060,N_3520,N_3405);
or U5061 (N_5061,N_3318,N_3301);
nor U5062 (N_5062,N_3693,N_3227);
nor U5063 (N_5063,N_2352,N_3748);
xor U5064 (N_5064,N_2324,N_2644);
xnor U5065 (N_5065,N_3410,N_3119);
and U5066 (N_5066,N_2569,N_3896);
xnor U5067 (N_5067,N_2487,N_3809);
nand U5068 (N_5068,N_3094,N_3417);
xnor U5069 (N_5069,N_2044,N_2147);
xnor U5070 (N_5070,N_3195,N_3691);
nand U5071 (N_5071,N_2433,N_3826);
nor U5072 (N_5072,N_3477,N_2229);
nand U5073 (N_5073,N_3884,N_2515);
and U5074 (N_5074,N_3964,N_3050);
and U5075 (N_5075,N_3642,N_2001);
or U5076 (N_5076,N_2138,N_3059);
nor U5077 (N_5077,N_3033,N_2711);
or U5078 (N_5078,N_3644,N_2942);
xnor U5079 (N_5079,N_3167,N_3398);
nor U5080 (N_5080,N_3172,N_3604);
xor U5081 (N_5081,N_2347,N_2642);
nand U5082 (N_5082,N_3235,N_2344);
nor U5083 (N_5083,N_3323,N_2185);
nor U5084 (N_5084,N_3729,N_2553);
or U5085 (N_5085,N_2409,N_2701);
or U5086 (N_5086,N_2439,N_2120);
xor U5087 (N_5087,N_2712,N_2304);
nor U5088 (N_5088,N_3827,N_2035);
and U5089 (N_5089,N_2859,N_3413);
nor U5090 (N_5090,N_2747,N_3429);
nand U5091 (N_5091,N_2202,N_2613);
nor U5092 (N_5092,N_2041,N_3705);
or U5093 (N_5093,N_2966,N_2833);
xnor U5094 (N_5094,N_3627,N_2759);
nor U5095 (N_5095,N_3815,N_2118);
or U5096 (N_5096,N_3325,N_2315);
xnor U5097 (N_5097,N_3354,N_2333);
nor U5098 (N_5098,N_3156,N_3040);
nor U5099 (N_5099,N_2104,N_2325);
xnor U5100 (N_5100,N_2892,N_3897);
or U5101 (N_5101,N_2970,N_3483);
nand U5102 (N_5102,N_3502,N_2672);
nor U5103 (N_5103,N_2854,N_2143);
nand U5104 (N_5104,N_2150,N_3290);
nor U5105 (N_5105,N_2440,N_2931);
xor U5106 (N_5106,N_3559,N_3724);
and U5107 (N_5107,N_2019,N_3428);
xor U5108 (N_5108,N_3030,N_2072);
or U5109 (N_5109,N_2846,N_2014);
nor U5110 (N_5110,N_3231,N_3234);
xnor U5111 (N_5111,N_2437,N_2524);
nand U5112 (N_5112,N_3955,N_2882);
xnor U5113 (N_5113,N_3856,N_3946);
or U5114 (N_5114,N_3033,N_3941);
and U5115 (N_5115,N_3888,N_2078);
or U5116 (N_5116,N_2978,N_2625);
nor U5117 (N_5117,N_2876,N_2403);
and U5118 (N_5118,N_3609,N_3297);
xor U5119 (N_5119,N_2255,N_2622);
nor U5120 (N_5120,N_2175,N_3705);
xnor U5121 (N_5121,N_3492,N_2083);
nor U5122 (N_5122,N_2364,N_3397);
and U5123 (N_5123,N_2255,N_2749);
and U5124 (N_5124,N_3170,N_2383);
and U5125 (N_5125,N_3748,N_3384);
xnor U5126 (N_5126,N_3756,N_2498);
nor U5127 (N_5127,N_2953,N_3645);
or U5128 (N_5128,N_2299,N_3638);
xnor U5129 (N_5129,N_2229,N_3434);
xor U5130 (N_5130,N_2848,N_2348);
nand U5131 (N_5131,N_3183,N_2751);
xor U5132 (N_5132,N_2810,N_3289);
and U5133 (N_5133,N_3691,N_2822);
xor U5134 (N_5134,N_2932,N_2927);
or U5135 (N_5135,N_3195,N_3026);
nand U5136 (N_5136,N_3323,N_3951);
nand U5137 (N_5137,N_3130,N_3348);
and U5138 (N_5138,N_3996,N_3486);
and U5139 (N_5139,N_2296,N_2785);
nor U5140 (N_5140,N_2777,N_2210);
and U5141 (N_5141,N_3071,N_3142);
nor U5142 (N_5142,N_3606,N_2644);
xor U5143 (N_5143,N_3499,N_2438);
and U5144 (N_5144,N_3026,N_2850);
or U5145 (N_5145,N_3858,N_2680);
and U5146 (N_5146,N_3561,N_2615);
nand U5147 (N_5147,N_2593,N_3232);
nand U5148 (N_5148,N_2645,N_3270);
and U5149 (N_5149,N_2747,N_3077);
xor U5150 (N_5150,N_3550,N_2642);
or U5151 (N_5151,N_3358,N_3340);
nor U5152 (N_5152,N_2830,N_2580);
xnor U5153 (N_5153,N_3567,N_2421);
nor U5154 (N_5154,N_2494,N_3020);
and U5155 (N_5155,N_2821,N_3396);
nand U5156 (N_5156,N_2758,N_2871);
nor U5157 (N_5157,N_2286,N_2265);
nand U5158 (N_5158,N_3458,N_2106);
nor U5159 (N_5159,N_3377,N_3340);
and U5160 (N_5160,N_2361,N_2813);
nand U5161 (N_5161,N_2682,N_3409);
nand U5162 (N_5162,N_2639,N_3531);
or U5163 (N_5163,N_3136,N_2418);
nand U5164 (N_5164,N_2397,N_3056);
xnor U5165 (N_5165,N_2017,N_3483);
and U5166 (N_5166,N_3242,N_2902);
nand U5167 (N_5167,N_2697,N_3420);
xnor U5168 (N_5168,N_2600,N_2873);
or U5169 (N_5169,N_2775,N_3845);
or U5170 (N_5170,N_3766,N_3512);
or U5171 (N_5171,N_3844,N_3818);
and U5172 (N_5172,N_2703,N_2960);
or U5173 (N_5173,N_2415,N_3954);
nor U5174 (N_5174,N_3973,N_3172);
xor U5175 (N_5175,N_2367,N_3880);
xnor U5176 (N_5176,N_3664,N_3689);
nand U5177 (N_5177,N_3125,N_3713);
nand U5178 (N_5178,N_3870,N_3974);
nand U5179 (N_5179,N_3856,N_2093);
and U5180 (N_5180,N_2440,N_2456);
xnor U5181 (N_5181,N_3477,N_2693);
and U5182 (N_5182,N_3861,N_2292);
nor U5183 (N_5183,N_3408,N_2435);
nor U5184 (N_5184,N_2588,N_2618);
and U5185 (N_5185,N_2580,N_2828);
or U5186 (N_5186,N_2222,N_2791);
and U5187 (N_5187,N_3752,N_2040);
and U5188 (N_5188,N_3652,N_3856);
nor U5189 (N_5189,N_3546,N_2029);
and U5190 (N_5190,N_3764,N_2308);
xnor U5191 (N_5191,N_2893,N_2061);
xor U5192 (N_5192,N_2911,N_2976);
and U5193 (N_5193,N_3395,N_2793);
xor U5194 (N_5194,N_3242,N_3987);
nor U5195 (N_5195,N_2213,N_2707);
and U5196 (N_5196,N_3001,N_2354);
nor U5197 (N_5197,N_2380,N_3862);
and U5198 (N_5198,N_3193,N_3949);
xnor U5199 (N_5199,N_2983,N_3584);
nand U5200 (N_5200,N_2789,N_3868);
xor U5201 (N_5201,N_2385,N_3214);
nand U5202 (N_5202,N_2347,N_2485);
or U5203 (N_5203,N_2112,N_2902);
nand U5204 (N_5204,N_2744,N_3105);
nor U5205 (N_5205,N_2964,N_3095);
nand U5206 (N_5206,N_3524,N_3044);
xor U5207 (N_5207,N_2636,N_2716);
xnor U5208 (N_5208,N_2541,N_3756);
and U5209 (N_5209,N_2397,N_2140);
and U5210 (N_5210,N_2141,N_2498);
nor U5211 (N_5211,N_2045,N_3466);
nor U5212 (N_5212,N_3213,N_3285);
xor U5213 (N_5213,N_2035,N_3031);
and U5214 (N_5214,N_2750,N_3779);
and U5215 (N_5215,N_3419,N_3262);
nand U5216 (N_5216,N_3601,N_3395);
or U5217 (N_5217,N_3099,N_3367);
and U5218 (N_5218,N_3943,N_3799);
xor U5219 (N_5219,N_2517,N_2022);
nand U5220 (N_5220,N_2844,N_2747);
nor U5221 (N_5221,N_3151,N_2292);
xor U5222 (N_5222,N_3702,N_3580);
nor U5223 (N_5223,N_3152,N_2064);
and U5224 (N_5224,N_3656,N_3348);
or U5225 (N_5225,N_2607,N_3308);
or U5226 (N_5226,N_3991,N_2576);
and U5227 (N_5227,N_2018,N_3103);
nor U5228 (N_5228,N_2107,N_2134);
nor U5229 (N_5229,N_3668,N_3029);
or U5230 (N_5230,N_3687,N_3710);
and U5231 (N_5231,N_3628,N_2450);
xnor U5232 (N_5232,N_3610,N_3977);
and U5233 (N_5233,N_2605,N_2311);
nor U5234 (N_5234,N_3701,N_3236);
or U5235 (N_5235,N_3325,N_2644);
and U5236 (N_5236,N_3300,N_2480);
or U5237 (N_5237,N_2123,N_3211);
xnor U5238 (N_5238,N_2729,N_2831);
nand U5239 (N_5239,N_3597,N_3878);
nand U5240 (N_5240,N_3484,N_2777);
or U5241 (N_5241,N_2740,N_2041);
xnor U5242 (N_5242,N_3641,N_2888);
and U5243 (N_5243,N_3100,N_3637);
nand U5244 (N_5244,N_2810,N_2572);
nand U5245 (N_5245,N_3312,N_3416);
or U5246 (N_5246,N_2186,N_2656);
nor U5247 (N_5247,N_3431,N_3902);
nand U5248 (N_5248,N_3890,N_3307);
or U5249 (N_5249,N_2356,N_3124);
and U5250 (N_5250,N_3495,N_3398);
or U5251 (N_5251,N_3574,N_3523);
xnor U5252 (N_5252,N_2178,N_3077);
nand U5253 (N_5253,N_3169,N_2667);
xnor U5254 (N_5254,N_2656,N_3152);
xnor U5255 (N_5255,N_3859,N_2945);
and U5256 (N_5256,N_3251,N_3234);
nand U5257 (N_5257,N_3556,N_2445);
nor U5258 (N_5258,N_3801,N_2206);
and U5259 (N_5259,N_2283,N_3225);
xnor U5260 (N_5260,N_2047,N_3150);
xor U5261 (N_5261,N_3763,N_2393);
or U5262 (N_5262,N_2854,N_2318);
xnor U5263 (N_5263,N_3510,N_3190);
nor U5264 (N_5264,N_2350,N_3872);
nand U5265 (N_5265,N_3156,N_2749);
nand U5266 (N_5266,N_2552,N_2562);
nand U5267 (N_5267,N_2311,N_2992);
nor U5268 (N_5268,N_3999,N_3143);
xor U5269 (N_5269,N_2112,N_3721);
and U5270 (N_5270,N_3878,N_3963);
xor U5271 (N_5271,N_3203,N_2415);
or U5272 (N_5272,N_2681,N_3475);
nand U5273 (N_5273,N_2846,N_2889);
or U5274 (N_5274,N_3973,N_2411);
nor U5275 (N_5275,N_3619,N_3272);
xor U5276 (N_5276,N_3196,N_2213);
nand U5277 (N_5277,N_3486,N_3418);
nand U5278 (N_5278,N_2708,N_2208);
nor U5279 (N_5279,N_3316,N_3907);
nand U5280 (N_5280,N_3778,N_2904);
and U5281 (N_5281,N_3197,N_3754);
nand U5282 (N_5282,N_3720,N_3782);
xnor U5283 (N_5283,N_3058,N_2149);
and U5284 (N_5284,N_3310,N_3495);
xnor U5285 (N_5285,N_2310,N_2825);
nor U5286 (N_5286,N_3981,N_2799);
nor U5287 (N_5287,N_2106,N_3434);
nor U5288 (N_5288,N_2816,N_3729);
nand U5289 (N_5289,N_3861,N_2964);
nand U5290 (N_5290,N_2379,N_2815);
or U5291 (N_5291,N_2049,N_2686);
nor U5292 (N_5292,N_3863,N_3067);
xor U5293 (N_5293,N_2607,N_3297);
xnor U5294 (N_5294,N_2155,N_2392);
and U5295 (N_5295,N_3617,N_2154);
or U5296 (N_5296,N_3300,N_3233);
or U5297 (N_5297,N_2798,N_2298);
nand U5298 (N_5298,N_2981,N_2074);
and U5299 (N_5299,N_3986,N_3943);
xnor U5300 (N_5300,N_2004,N_2384);
nand U5301 (N_5301,N_3428,N_2463);
nor U5302 (N_5302,N_2279,N_2272);
xnor U5303 (N_5303,N_2016,N_3498);
or U5304 (N_5304,N_2365,N_3220);
or U5305 (N_5305,N_3468,N_3142);
and U5306 (N_5306,N_3940,N_3865);
and U5307 (N_5307,N_3656,N_3045);
xor U5308 (N_5308,N_2711,N_2513);
or U5309 (N_5309,N_2418,N_2068);
nor U5310 (N_5310,N_2674,N_3689);
nor U5311 (N_5311,N_2401,N_2601);
xnor U5312 (N_5312,N_3088,N_2455);
or U5313 (N_5313,N_2645,N_3538);
or U5314 (N_5314,N_3778,N_2921);
xor U5315 (N_5315,N_3980,N_2528);
nand U5316 (N_5316,N_2144,N_2758);
or U5317 (N_5317,N_2042,N_3470);
or U5318 (N_5318,N_3680,N_2330);
nor U5319 (N_5319,N_2088,N_2780);
and U5320 (N_5320,N_3753,N_3882);
or U5321 (N_5321,N_2350,N_3153);
nand U5322 (N_5322,N_2331,N_2499);
or U5323 (N_5323,N_2098,N_2253);
nand U5324 (N_5324,N_3138,N_2587);
nand U5325 (N_5325,N_3852,N_3568);
nand U5326 (N_5326,N_3836,N_3443);
nand U5327 (N_5327,N_2355,N_3573);
or U5328 (N_5328,N_2400,N_2076);
nor U5329 (N_5329,N_2609,N_2960);
or U5330 (N_5330,N_3409,N_2612);
xnor U5331 (N_5331,N_3507,N_3677);
nand U5332 (N_5332,N_2957,N_2977);
nand U5333 (N_5333,N_3815,N_3805);
xnor U5334 (N_5334,N_3171,N_2699);
or U5335 (N_5335,N_3319,N_2630);
and U5336 (N_5336,N_3548,N_2898);
nand U5337 (N_5337,N_3072,N_2874);
nand U5338 (N_5338,N_3201,N_3814);
nor U5339 (N_5339,N_2596,N_2696);
or U5340 (N_5340,N_3805,N_2935);
nand U5341 (N_5341,N_3990,N_2277);
nor U5342 (N_5342,N_3671,N_3988);
xnor U5343 (N_5343,N_2277,N_3083);
and U5344 (N_5344,N_2673,N_2629);
xor U5345 (N_5345,N_3026,N_3557);
or U5346 (N_5346,N_3488,N_2971);
and U5347 (N_5347,N_3712,N_2022);
xnor U5348 (N_5348,N_2204,N_3579);
and U5349 (N_5349,N_3313,N_2065);
nand U5350 (N_5350,N_3408,N_2574);
xor U5351 (N_5351,N_2278,N_3223);
nor U5352 (N_5352,N_2972,N_3393);
nand U5353 (N_5353,N_2014,N_3903);
xor U5354 (N_5354,N_3166,N_3946);
nand U5355 (N_5355,N_2853,N_2532);
nand U5356 (N_5356,N_2111,N_3964);
nand U5357 (N_5357,N_2092,N_3451);
nor U5358 (N_5358,N_2529,N_2364);
nand U5359 (N_5359,N_3119,N_2124);
and U5360 (N_5360,N_3710,N_2133);
xor U5361 (N_5361,N_2764,N_2878);
or U5362 (N_5362,N_2363,N_2827);
or U5363 (N_5363,N_3348,N_3524);
xnor U5364 (N_5364,N_3845,N_3814);
nand U5365 (N_5365,N_2655,N_3931);
nand U5366 (N_5366,N_3813,N_2651);
nand U5367 (N_5367,N_2676,N_3514);
nor U5368 (N_5368,N_2637,N_3211);
or U5369 (N_5369,N_2478,N_3423);
nand U5370 (N_5370,N_3967,N_2399);
and U5371 (N_5371,N_3433,N_3633);
or U5372 (N_5372,N_3407,N_3896);
xor U5373 (N_5373,N_2875,N_3077);
or U5374 (N_5374,N_2520,N_2928);
nand U5375 (N_5375,N_2814,N_3771);
xnor U5376 (N_5376,N_3610,N_3620);
nor U5377 (N_5377,N_3514,N_2765);
and U5378 (N_5378,N_3833,N_2738);
or U5379 (N_5379,N_3075,N_2292);
nand U5380 (N_5380,N_3400,N_3071);
or U5381 (N_5381,N_2020,N_2439);
and U5382 (N_5382,N_3931,N_3716);
nor U5383 (N_5383,N_3112,N_3027);
nand U5384 (N_5384,N_3453,N_3691);
nand U5385 (N_5385,N_2730,N_2505);
nor U5386 (N_5386,N_3227,N_3318);
xor U5387 (N_5387,N_3347,N_3694);
or U5388 (N_5388,N_3703,N_3590);
nand U5389 (N_5389,N_2457,N_2004);
or U5390 (N_5390,N_3038,N_2170);
and U5391 (N_5391,N_3851,N_3057);
and U5392 (N_5392,N_2762,N_3380);
xnor U5393 (N_5393,N_3596,N_3484);
nor U5394 (N_5394,N_3477,N_2494);
xnor U5395 (N_5395,N_2879,N_2403);
and U5396 (N_5396,N_2901,N_2617);
nand U5397 (N_5397,N_2081,N_3920);
nor U5398 (N_5398,N_2811,N_2977);
and U5399 (N_5399,N_3262,N_3345);
nor U5400 (N_5400,N_3344,N_2259);
nor U5401 (N_5401,N_2327,N_2757);
xnor U5402 (N_5402,N_3548,N_3570);
nor U5403 (N_5403,N_2613,N_3145);
nand U5404 (N_5404,N_2075,N_3034);
nand U5405 (N_5405,N_3084,N_2091);
nor U5406 (N_5406,N_3231,N_3040);
or U5407 (N_5407,N_3141,N_2780);
xnor U5408 (N_5408,N_3326,N_2444);
nor U5409 (N_5409,N_2497,N_2928);
xor U5410 (N_5410,N_3079,N_2956);
xor U5411 (N_5411,N_2350,N_2133);
and U5412 (N_5412,N_2926,N_2111);
xor U5413 (N_5413,N_3105,N_3204);
xor U5414 (N_5414,N_2690,N_3413);
nor U5415 (N_5415,N_3961,N_2013);
or U5416 (N_5416,N_2088,N_3710);
xor U5417 (N_5417,N_3580,N_2474);
or U5418 (N_5418,N_2240,N_2511);
xnor U5419 (N_5419,N_2426,N_3306);
or U5420 (N_5420,N_2205,N_3347);
and U5421 (N_5421,N_2023,N_2958);
nor U5422 (N_5422,N_2656,N_3330);
nand U5423 (N_5423,N_2336,N_3045);
xnor U5424 (N_5424,N_2786,N_2289);
nand U5425 (N_5425,N_2784,N_2803);
nand U5426 (N_5426,N_2577,N_2063);
xor U5427 (N_5427,N_2203,N_3696);
nand U5428 (N_5428,N_3380,N_2121);
and U5429 (N_5429,N_3389,N_3529);
nor U5430 (N_5430,N_2141,N_2555);
nand U5431 (N_5431,N_2572,N_2014);
or U5432 (N_5432,N_2397,N_2336);
or U5433 (N_5433,N_3333,N_3744);
nand U5434 (N_5434,N_3880,N_2373);
nand U5435 (N_5435,N_3875,N_2779);
nor U5436 (N_5436,N_3878,N_2720);
nor U5437 (N_5437,N_2376,N_2441);
nand U5438 (N_5438,N_3361,N_3340);
xnor U5439 (N_5439,N_3591,N_2836);
nand U5440 (N_5440,N_3080,N_2915);
nor U5441 (N_5441,N_3438,N_3731);
nand U5442 (N_5442,N_2651,N_3824);
nand U5443 (N_5443,N_3227,N_2559);
xor U5444 (N_5444,N_2519,N_3231);
and U5445 (N_5445,N_2761,N_3704);
or U5446 (N_5446,N_3209,N_2005);
nand U5447 (N_5447,N_3084,N_3227);
or U5448 (N_5448,N_2002,N_2008);
and U5449 (N_5449,N_3332,N_3716);
nor U5450 (N_5450,N_3666,N_3098);
xor U5451 (N_5451,N_3210,N_3373);
nor U5452 (N_5452,N_2294,N_3485);
and U5453 (N_5453,N_2826,N_3100);
and U5454 (N_5454,N_2918,N_3585);
nand U5455 (N_5455,N_3425,N_3151);
and U5456 (N_5456,N_3091,N_3748);
xnor U5457 (N_5457,N_2268,N_3368);
and U5458 (N_5458,N_2547,N_2098);
xnor U5459 (N_5459,N_3481,N_2723);
nor U5460 (N_5460,N_3520,N_2600);
nand U5461 (N_5461,N_2186,N_3741);
nor U5462 (N_5462,N_3058,N_2026);
and U5463 (N_5463,N_3503,N_3657);
or U5464 (N_5464,N_2238,N_2297);
or U5465 (N_5465,N_2968,N_3370);
xor U5466 (N_5466,N_2085,N_2782);
and U5467 (N_5467,N_3178,N_2169);
and U5468 (N_5468,N_3284,N_3310);
or U5469 (N_5469,N_3060,N_2362);
xor U5470 (N_5470,N_2906,N_2214);
xnor U5471 (N_5471,N_2877,N_2462);
and U5472 (N_5472,N_3731,N_2191);
or U5473 (N_5473,N_2806,N_2305);
nand U5474 (N_5474,N_2206,N_3153);
or U5475 (N_5475,N_2619,N_3449);
nand U5476 (N_5476,N_2990,N_3582);
or U5477 (N_5477,N_3996,N_2797);
nand U5478 (N_5478,N_3100,N_2465);
and U5479 (N_5479,N_2236,N_3362);
nor U5480 (N_5480,N_2745,N_3447);
nand U5481 (N_5481,N_2316,N_3963);
or U5482 (N_5482,N_2302,N_3152);
xnor U5483 (N_5483,N_2990,N_3550);
and U5484 (N_5484,N_3281,N_2298);
or U5485 (N_5485,N_3421,N_3940);
xnor U5486 (N_5486,N_2988,N_3633);
nor U5487 (N_5487,N_2430,N_3313);
nand U5488 (N_5488,N_3803,N_2796);
nor U5489 (N_5489,N_3052,N_3163);
or U5490 (N_5490,N_2541,N_3181);
nor U5491 (N_5491,N_3997,N_2088);
xnor U5492 (N_5492,N_2276,N_2443);
and U5493 (N_5493,N_3283,N_3077);
nor U5494 (N_5494,N_3935,N_2456);
xor U5495 (N_5495,N_2627,N_3479);
nand U5496 (N_5496,N_3407,N_2066);
nor U5497 (N_5497,N_2340,N_2548);
or U5498 (N_5498,N_2740,N_2531);
or U5499 (N_5499,N_2679,N_2120);
nand U5500 (N_5500,N_3371,N_3634);
and U5501 (N_5501,N_3388,N_3636);
or U5502 (N_5502,N_2216,N_2572);
xnor U5503 (N_5503,N_2117,N_3048);
and U5504 (N_5504,N_3479,N_3974);
xor U5505 (N_5505,N_2967,N_3520);
nand U5506 (N_5506,N_3267,N_3506);
or U5507 (N_5507,N_3506,N_2485);
nand U5508 (N_5508,N_2599,N_3125);
nand U5509 (N_5509,N_2001,N_3673);
or U5510 (N_5510,N_2652,N_3413);
or U5511 (N_5511,N_2726,N_2078);
xor U5512 (N_5512,N_3302,N_2011);
or U5513 (N_5513,N_3318,N_2220);
nand U5514 (N_5514,N_2471,N_2659);
and U5515 (N_5515,N_3810,N_2935);
xor U5516 (N_5516,N_2417,N_2499);
xnor U5517 (N_5517,N_2573,N_3116);
and U5518 (N_5518,N_3620,N_2556);
nor U5519 (N_5519,N_2076,N_2729);
and U5520 (N_5520,N_2478,N_3705);
nand U5521 (N_5521,N_3861,N_3782);
xnor U5522 (N_5522,N_3440,N_3565);
nor U5523 (N_5523,N_2633,N_2199);
nor U5524 (N_5524,N_2633,N_3965);
nand U5525 (N_5525,N_2034,N_2095);
xor U5526 (N_5526,N_2421,N_3123);
or U5527 (N_5527,N_2456,N_2827);
or U5528 (N_5528,N_3521,N_3141);
nor U5529 (N_5529,N_2159,N_3628);
or U5530 (N_5530,N_2154,N_2347);
nand U5531 (N_5531,N_3758,N_2243);
nor U5532 (N_5532,N_2604,N_2357);
and U5533 (N_5533,N_2373,N_2759);
xnor U5534 (N_5534,N_3559,N_3215);
nand U5535 (N_5535,N_2596,N_3960);
or U5536 (N_5536,N_2799,N_2001);
or U5537 (N_5537,N_2914,N_2432);
xnor U5538 (N_5538,N_3793,N_2615);
nor U5539 (N_5539,N_3339,N_2926);
or U5540 (N_5540,N_2553,N_2877);
and U5541 (N_5541,N_3993,N_2386);
nand U5542 (N_5542,N_3606,N_3616);
or U5543 (N_5543,N_2034,N_2656);
and U5544 (N_5544,N_2988,N_2320);
nand U5545 (N_5545,N_2766,N_2183);
nand U5546 (N_5546,N_3815,N_3211);
and U5547 (N_5547,N_3843,N_3075);
nor U5548 (N_5548,N_2993,N_3206);
or U5549 (N_5549,N_3386,N_2899);
xor U5550 (N_5550,N_2382,N_2390);
or U5551 (N_5551,N_3721,N_2694);
nor U5552 (N_5552,N_2635,N_2295);
and U5553 (N_5553,N_2089,N_2934);
xor U5554 (N_5554,N_2827,N_3791);
nand U5555 (N_5555,N_2261,N_3209);
nand U5556 (N_5556,N_3457,N_2678);
or U5557 (N_5557,N_3935,N_3655);
or U5558 (N_5558,N_2562,N_3012);
xnor U5559 (N_5559,N_2391,N_2158);
nor U5560 (N_5560,N_2985,N_3553);
nand U5561 (N_5561,N_2831,N_2321);
nand U5562 (N_5562,N_3269,N_3915);
nand U5563 (N_5563,N_3678,N_2065);
nor U5564 (N_5564,N_2420,N_3061);
nand U5565 (N_5565,N_3343,N_3582);
or U5566 (N_5566,N_3739,N_3160);
and U5567 (N_5567,N_3008,N_2785);
and U5568 (N_5568,N_3402,N_3905);
and U5569 (N_5569,N_2984,N_2021);
nand U5570 (N_5570,N_3688,N_2166);
or U5571 (N_5571,N_3952,N_2936);
or U5572 (N_5572,N_3525,N_2880);
xnor U5573 (N_5573,N_3759,N_2602);
nand U5574 (N_5574,N_2827,N_3241);
and U5575 (N_5575,N_2751,N_2951);
nor U5576 (N_5576,N_2043,N_3500);
nand U5577 (N_5577,N_2690,N_2002);
nor U5578 (N_5578,N_2892,N_3787);
xor U5579 (N_5579,N_3616,N_3850);
nand U5580 (N_5580,N_3889,N_2368);
and U5581 (N_5581,N_2007,N_3568);
or U5582 (N_5582,N_3239,N_2797);
and U5583 (N_5583,N_3722,N_3247);
and U5584 (N_5584,N_3146,N_3556);
and U5585 (N_5585,N_3654,N_3988);
nor U5586 (N_5586,N_2791,N_2225);
nor U5587 (N_5587,N_3609,N_3384);
nand U5588 (N_5588,N_3289,N_3380);
and U5589 (N_5589,N_3467,N_2459);
or U5590 (N_5590,N_3289,N_3293);
or U5591 (N_5591,N_2626,N_2983);
xnor U5592 (N_5592,N_3305,N_3880);
xor U5593 (N_5593,N_2325,N_2227);
xor U5594 (N_5594,N_2939,N_3528);
nor U5595 (N_5595,N_2156,N_3770);
nand U5596 (N_5596,N_3002,N_2630);
nand U5597 (N_5597,N_2399,N_2110);
or U5598 (N_5598,N_3816,N_3717);
or U5599 (N_5599,N_2344,N_2120);
nand U5600 (N_5600,N_3074,N_2979);
and U5601 (N_5601,N_3553,N_3891);
xnor U5602 (N_5602,N_3286,N_2857);
and U5603 (N_5603,N_2674,N_3215);
and U5604 (N_5604,N_2446,N_2334);
xor U5605 (N_5605,N_2961,N_3497);
nand U5606 (N_5606,N_3587,N_2933);
xnor U5607 (N_5607,N_2692,N_2849);
and U5608 (N_5608,N_3448,N_2450);
and U5609 (N_5609,N_2812,N_3398);
xor U5610 (N_5610,N_3262,N_3465);
xnor U5611 (N_5611,N_3035,N_3871);
or U5612 (N_5612,N_3156,N_2331);
xnor U5613 (N_5613,N_3770,N_3674);
or U5614 (N_5614,N_2349,N_3656);
nor U5615 (N_5615,N_2874,N_2018);
nand U5616 (N_5616,N_3017,N_2617);
nand U5617 (N_5617,N_3737,N_2877);
nand U5618 (N_5618,N_2189,N_3182);
xnor U5619 (N_5619,N_2942,N_2517);
or U5620 (N_5620,N_3461,N_3562);
nand U5621 (N_5621,N_3741,N_3026);
nand U5622 (N_5622,N_2286,N_2503);
nor U5623 (N_5623,N_3314,N_2013);
and U5624 (N_5624,N_3822,N_2551);
xor U5625 (N_5625,N_2312,N_2424);
xor U5626 (N_5626,N_2933,N_3212);
and U5627 (N_5627,N_3397,N_3514);
or U5628 (N_5628,N_3672,N_2464);
nand U5629 (N_5629,N_3207,N_3836);
or U5630 (N_5630,N_3473,N_2106);
and U5631 (N_5631,N_2802,N_2805);
nor U5632 (N_5632,N_2363,N_3755);
xnor U5633 (N_5633,N_2801,N_3439);
and U5634 (N_5634,N_2130,N_2438);
xnor U5635 (N_5635,N_2684,N_3534);
and U5636 (N_5636,N_3738,N_3998);
or U5637 (N_5637,N_2714,N_2246);
xnor U5638 (N_5638,N_3468,N_2039);
and U5639 (N_5639,N_3938,N_2486);
or U5640 (N_5640,N_3265,N_2803);
or U5641 (N_5641,N_3063,N_3286);
and U5642 (N_5642,N_3556,N_2135);
xnor U5643 (N_5643,N_3151,N_2426);
nor U5644 (N_5644,N_3124,N_2165);
nand U5645 (N_5645,N_2081,N_2205);
nand U5646 (N_5646,N_2135,N_3017);
or U5647 (N_5647,N_2204,N_2962);
and U5648 (N_5648,N_2424,N_3879);
or U5649 (N_5649,N_3863,N_2858);
and U5650 (N_5650,N_2315,N_2471);
and U5651 (N_5651,N_3678,N_3361);
and U5652 (N_5652,N_2209,N_3251);
and U5653 (N_5653,N_3846,N_3658);
xnor U5654 (N_5654,N_3250,N_3982);
or U5655 (N_5655,N_3272,N_3029);
nand U5656 (N_5656,N_2625,N_3884);
xor U5657 (N_5657,N_2570,N_2306);
nand U5658 (N_5658,N_2048,N_3209);
nand U5659 (N_5659,N_2283,N_2340);
or U5660 (N_5660,N_3749,N_2882);
and U5661 (N_5661,N_2505,N_3356);
nand U5662 (N_5662,N_2950,N_2146);
and U5663 (N_5663,N_3669,N_2367);
nand U5664 (N_5664,N_2062,N_3938);
and U5665 (N_5665,N_3083,N_2645);
nor U5666 (N_5666,N_3471,N_2916);
nor U5667 (N_5667,N_2548,N_2332);
xor U5668 (N_5668,N_3067,N_3181);
xor U5669 (N_5669,N_3637,N_3796);
and U5670 (N_5670,N_3016,N_3160);
or U5671 (N_5671,N_3097,N_2617);
nor U5672 (N_5672,N_2684,N_3408);
or U5673 (N_5673,N_3566,N_2983);
xor U5674 (N_5674,N_2424,N_2766);
or U5675 (N_5675,N_2039,N_2947);
nand U5676 (N_5676,N_3655,N_2378);
and U5677 (N_5677,N_2413,N_3653);
or U5678 (N_5678,N_3055,N_2458);
and U5679 (N_5679,N_3989,N_3877);
and U5680 (N_5680,N_2966,N_3280);
nor U5681 (N_5681,N_3224,N_3167);
and U5682 (N_5682,N_2287,N_2326);
nand U5683 (N_5683,N_3096,N_2898);
nor U5684 (N_5684,N_2406,N_2961);
nand U5685 (N_5685,N_2888,N_2822);
or U5686 (N_5686,N_3402,N_2844);
and U5687 (N_5687,N_3187,N_3468);
nand U5688 (N_5688,N_3561,N_3721);
nor U5689 (N_5689,N_2761,N_2533);
and U5690 (N_5690,N_2630,N_3070);
or U5691 (N_5691,N_3215,N_2368);
or U5692 (N_5692,N_3113,N_3867);
xor U5693 (N_5693,N_3081,N_3517);
nor U5694 (N_5694,N_2922,N_2109);
and U5695 (N_5695,N_3988,N_3535);
and U5696 (N_5696,N_2920,N_2167);
or U5697 (N_5697,N_2034,N_2742);
nor U5698 (N_5698,N_2309,N_2403);
or U5699 (N_5699,N_2812,N_3864);
nor U5700 (N_5700,N_2105,N_2880);
nand U5701 (N_5701,N_2323,N_3054);
and U5702 (N_5702,N_3397,N_3138);
or U5703 (N_5703,N_3614,N_2590);
nand U5704 (N_5704,N_3776,N_2411);
nand U5705 (N_5705,N_3288,N_2023);
nor U5706 (N_5706,N_3747,N_2736);
xor U5707 (N_5707,N_3966,N_2995);
or U5708 (N_5708,N_2256,N_2328);
and U5709 (N_5709,N_3095,N_2921);
or U5710 (N_5710,N_3908,N_3618);
xor U5711 (N_5711,N_2354,N_3772);
and U5712 (N_5712,N_3883,N_2577);
or U5713 (N_5713,N_2249,N_2600);
and U5714 (N_5714,N_2389,N_2439);
or U5715 (N_5715,N_2843,N_2719);
and U5716 (N_5716,N_2686,N_2527);
xnor U5717 (N_5717,N_2261,N_3840);
nor U5718 (N_5718,N_2535,N_3400);
nor U5719 (N_5719,N_2563,N_2511);
xnor U5720 (N_5720,N_3540,N_3820);
nor U5721 (N_5721,N_2517,N_2063);
nor U5722 (N_5722,N_2049,N_2947);
or U5723 (N_5723,N_3123,N_2643);
and U5724 (N_5724,N_2631,N_2898);
nor U5725 (N_5725,N_2667,N_3552);
nor U5726 (N_5726,N_3394,N_2573);
nand U5727 (N_5727,N_2256,N_3987);
nand U5728 (N_5728,N_2933,N_3948);
and U5729 (N_5729,N_3704,N_2062);
nor U5730 (N_5730,N_3977,N_2132);
or U5731 (N_5731,N_2498,N_2726);
and U5732 (N_5732,N_3452,N_3136);
nand U5733 (N_5733,N_2035,N_2103);
nor U5734 (N_5734,N_2025,N_2752);
nor U5735 (N_5735,N_3827,N_2466);
nand U5736 (N_5736,N_2395,N_2152);
and U5737 (N_5737,N_3870,N_2155);
nand U5738 (N_5738,N_3579,N_2521);
or U5739 (N_5739,N_2336,N_3881);
and U5740 (N_5740,N_2154,N_3189);
xor U5741 (N_5741,N_2562,N_3385);
and U5742 (N_5742,N_3093,N_2281);
xor U5743 (N_5743,N_2207,N_2812);
xor U5744 (N_5744,N_2787,N_3783);
nand U5745 (N_5745,N_2725,N_2121);
or U5746 (N_5746,N_3760,N_3316);
or U5747 (N_5747,N_3546,N_3745);
nor U5748 (N_5748,N_2500,N_3706);
and U5749 (N_5749,N_3010,N_2004);
and U5750 (N_5750,N_2097,N_3118);
or U5751 (N_5751,N_2381,N_2116);
nor U5752 (N_5752,N_3478,N_2427);
xnor U5753 (N_5753,N_3683,N_3205);
or U5754 (N_5754,N_3327,N_3890);
and U5755 (N_5755,N_3132,N_3044);
nor U5756 (N_5756,N_2220,N_2492);
and U5757 (N_5757,N_3451,N_2105);
nand U5758 (N_5758,N_3903,N_3787);
or U5759 (N_5759,N_3922,N_3014);
and U5760 (N_5760,N_3112,N_3430);
xor U5761 (N_5761,N_3462,N_2504);
nand U5762 (N_5762,N_3688,N_3227);
xnor U5763 (N_5763,N_3506,N_2746);
nor U5764 (N_5764,N_2569,N_3528);
or U5765 (N_5765,N_2746,N_2963);
nand U5766 (N_5766,N_3305,N_2738);
and U5767 (N_5767,N_3498,N_3711);
nor U5768 (N_5768,N_2989,N_2080);
and U5769 (N_5769,N_3990,N_3027);
and U5770 (N_5770,N_2178,N_2451);
nand U5771 (N_5771,N_3101,N_3940);
and U5772 (N_5772,N_2149,N_3947);
nand U5773 (N_5773,N_3193,N_2861);
xor U5774 (N_5774,N_3003,N_3608);
nand U5775 (N_5775,N_3642,N_2931);
nand U5776 (N_5776,N_3279,N_2931);
xor U5777 (N_5777,N_2156,N_3496);
or U5778 (N_5778,N_3156,N_3716);
and U5779 (N_5779,N_3852,N_3103);
and U5780 (N_5780,N_3760,N_3614);
nand U5781 (N_5781,N_3903,N_2274);
nand U5782 (N_5782,N_3165,N_2822);
nand U5783 (N_5783,N_3118,N_2940);
or U5784 (N_5784,N_3527,N_3096);
or U5785 (N_5785,N_3785,N_2872);
and U5786 (N_5786,N_2595,N_3696);
or U5787 (N_5787,N_3120,N_2769);
nor U5788 (N_5788,N_3861,N_2939);
nand U5789 (N_5789,N_2624,N_2832);
nand U5790 (N_5790,N_2178,N_3702);
xor U5791 (N_5791,N_2293,N_3547);
nor U5792 (N_5792,N_3719,N_2559);
nor U5793 (N_5793,N_2498,N_2942);
or U5794 (N_5794,N_2420,N_2842);
nand U5795 (N_5795,N_3907,N_2301);
or U5796 (N_5796,N_2532,N_3963);
xor U5797 (N_5797,N_2255,N_3121);
xnor U5798 (N_5798,N_2481,N_3257);
nand U5799 (N_5799,N_2098,N_2042);
nand U5800 (N_5800,N_2306,N_3600);
xor U5801 (N_5801,N_2399,N_2982);
nor U5802 (N_5802,N_3975,N_2746);
xor U5803 (N_5803,N_3350,N_2822);
or U5804 (N_5804,N_2755,N_2169);
nor U5805 (N_5805,N_3287,N_3639);
nor U5806 (N_5806,N_2335,N_3768);
nand U5807 (N_5807,N_3553,N_3162);
nor U5808 (N_5808,N_2991,N_3148);
nand U5809 (N_5809,N_3220,N_3530);
and U5810 (N_5810,N_2106,N_3940);
or U5811 (N_5811,N_3993,N_2666);
nand U5812 (N_5812,N_3581,N_2874);
or U5813 (N_5813,N_2034,N_2511);
and U5814 (N_5814,N_2708,N_2783);
or U5815 (N_5815,N_3560,N_2904);
xor U5816 (N_5816,N_2302,N_3057);
xor U5817 (N_5817,N_2146,N_2756);
nor U5818 (N_5818,N_2111,N_3795);
and U5819 (N_5819,N_3040,N_2107);
or U5820 (N_5820,N_2173,N_3466);
and U5821 (N_5821,N_3335,N_2740);
nand U5822 (N_5822,N_2398,N_3498);
or U5823 (N_5823,N_2508,N_2777);
nand U5824 (N_5824,N_3004,N_3123);
xnor U5825 (N_5825,N_2263,N_3341);
and U5826 (N_5826,N_3249,N_3377);
xnor U5827 (N_5827,N_3459,N_2285);
xor U5828 (N_5828,N_3677,N_3271);
xnor U5829 (N_5829,N_3824,N_3679);
or U5830 (N_5830,N_2758,N_3477);
xor U5831 (N_5831,N_2232,N_3306);
xor U5832 (N_5832,N_3319,N_3600);
nor U5833 (N_5833,N_2068,N_3878);
and U5834 (N_5834,N_3489,N_2252);
and U5835 (N_5835,N_2742,N_2253);
xor U5836 (N_5836,N_2042,N_3783);
nand U5837 (N_5837,N_2012,N_3575);
or U5838 (N_5838,N_3155,N_3950);
and U5839 (N_5839,N_3858,N_3314);
nor U5840 (N_5840,N_3772,N_2941);
xnor U5841 (N_5841,N_2655,N_3818);
xor U5842 (N_5842,N_3375,N_2385);
nor U5843 (N_5843,N_2655,N_2385);
nand U5844 (N_5844,N_3793,N_2255);
nor U5845 (N_5845,N_3789,N_2073);
nand U5846 (N_5846,N_2215,N_3800);
xnor U5847 (N_5847,N_2924,N_2364);
or U5848 (N_5848,N_3376,N_3382);
and U5849 (N_5849,N_2651,N_3044);
or U5850 (N_5850,N_3404,N_2638);
and U5851 (N_5851,N_2019,N_3131);
and U5852 (N_5852,N_2101,N_3359);
nand U5853 (N_5853,N_2022,N_2230);
nor U5854 (N_5854,N_3920,N_3246);
xor U5855 (N_5855,N_2556,N_2974);
nand U5856 (N_5856,N_2651,N_2945);
xor U5857 (N_5857,N_2280,N_2288);
and U5858 (N_5858,N_2337,N_3550);
nor U5859 (N_5859,N_3824,N_2143);
and U5860 (N_5860,N_2563,N_3359);
nor U5861 (N_5861,N_2949,N_2356);
or U5862 (N_5862,N_2365,N_2626);
and U5863 (N_5863,N_3122,N_2740);
nand U5864 (N_5864,N_2175,N_2171);
or U5865 (N_5865,N_3532,N_2331);
or U5866 (N_5866,N_3348,N_2355);
xnor U5867 (N_5867,N_3712,N_3554);
or U5868 (N_5868,N_2758,N_3850);
nor U5869 (N_5869,N_3592,N_2082);
nor U5870 (N_5870,N_2615,N_2133);
and U5871 (N_5871,N_3737,N_3419);
or U5872 (N_5872,N_2312,N_3869);
and U5873 (N_5873,N_2658,N_2725);
and U5874 (N_5874,N_2207,N_2505);
nor U5875 (N_5875,N_2224,N_3279);
nor U5876 (N_5876,N_2355,N_3120);
and U5877 (N_5877,N_3179,N_2486);
nand U5878 (N_5878,N_2098,N_3330);
and U5879 (N_5879,N_2775,N_3725);
and U5880 (N_5880,N_2367,N_2527);
xor U5881 (N_5881,N_3066,N_3240);
or U5882 (N_5882,N_3342,N_2427);
xor U5883 (N_5883,N_2414,N_2972);
nand U5884 (N_5884,N_3704,N_2441);
nor U5885 (N_5885,N_3072,N_3378);
xor U5886 (N_5886,N_3151,N_3478);
xnor U5887 (N_5887,N_3055,N_3373);
and U5888 (N_5888,N_2219,N_3741);
nand U5889 (N_5889,N_2687,N_2765);
nand U5890 (N_5890,N_3019,N_2544);
nand U5891 (N_5891,N_3562,N_3366);
nor U5892 (N_5892,N_3676,N_3497);
nand U5893 (N_5893,N_2380,N_2144);
nand U5894 (N_5894,N_3858,N_2846);
or U5895 (N_5895,N_3827,N_2107);
xnor U5896 (N_5896,N_2793,N_2458);
nor U5897 (N_5897,N_3312,N_3684);
or U5898 (N_5898,N_3064,N_3040);
nor U5899 (N_5899,N_2946,N_2407);
nand U5900 (N_5900,N_2207,N_2799);
and U5901 (N_5901,N_3355,N_2709);
xnor U5902 (N_5902,N_2125,N_3441);
or U5903 (N_5903,N_3898,N_2215);
xor U5904 (N_5904,N_2186,N_3723);
nand U5905 (N_5905,N_2897,N_2158);
xor U5906 (N_5906,N_3120,N_3106);
nor U5907 (N_5907,N_3106,N_3139);
and U5908 (N_5908,N_3613,N_2927);
and U5909 (N_5909,N_2374,N_2698);
and U5910 (N_5910,N_2312,N_3455);
and U5911 (N_5911,N_2250,N_2519);
nand U5912 (N_5912,N_3426,N_3755);
xnor U5913 (N_5913,N_3796,N_2576);
and U5914 (N_5914,N_2758,N_3089);
and U5915 (N_5915,N_2987,N_3782);
nor U5916 (N_5916,N_3665,N_2190);
or U5917 (N_5917,N_3241,N_2464);
and U5918 (N_5918,N_3859,N_2727);
or U5919 (N_5919,N_2083,N_2474);
or U5920 (N_5920,N_3362,N_2063);
and U5921 (N_5921,N_3305,N_2302);
nand U5922 (N_5922,N_3537,N_3547);
nor U5923 (N_5923,N_2968,N_2678);
nand U5924 (N_5924,N_2665,N_3134);
xnor U5925 (N_5925,N_2801,N_2309);
nor U5926 (N_5926,N_2743,N_2199);
or U5927 (N_5927,N_3535,N_3787);
nor U5928 (N_5928,N_2725,N_3318);
nand U5929 (N_5929,N_2848,N_2277);
xnor U5930 (N_5930,N_2821,N_2027);
and U5931 (N_5931,N_3322,N_2768);
or U5932 (N_5932,N_2940,N_2032);
nor U5933 (N_5933,N_3804,N_3779);
xnor U5934 (N_5934,N_3828,N_3262);
nor U5935 (N_5935,N_2798,N_2904);
nor U5936 (N_5936,N_2656,N_3431);
nor U5937 (N_5937,N_3372,N_2351);
nor U5938 (N_5938,N_3689,N_3818);
and U5939 (N_5939,N_2826,N_2632);
nand U5940 (N_5940,N_3759,N_3798);
and U5941 (N_5941,N_3258,N_2866);
xnor U5942 (N_5942,N_2073,N_3956);
or U5943 (N_5943,N_3895,N_3367);
xor U5944 (N_5944,N_2469,N_2125);
xor U5945 (N_5945,N_2889,N_2775);
nor U5946 (N_5946,N_3112,N_3440);
and U5947 (N_5947,N_3982,N_3125);
nand U5948 (N_5948,N_3808,N_3261);
or U5949 (N_5949,N_3507,N_2748);
or U5950 (N_5950,N_2426,N_2379);
nand U5951 (N_5951,N_3362,N_2106);
or U5952 (N_5952,N_3184,N_3517);
nor U5953 (N_5953,N_2373,N_3202);
or U5954 (N_5954,N_2325,N_3498);
nor U5955 (N_5955,N_2648,N_2328);
and U5956 (N_5956,N_2451,N_2029);
xnor U5957 (N_5957,N_2852,N_2409);
or U5958 (N_5958,N_3600,N_3440);
or U5959 (N_5959,N_3814,N_2896);
and U5960 (N_5960,N_3121,N_2472);
nor U5961 (N_5961,N_3025,N_3592);
nand U5962 (N_5962,N_2138,N_2453);
xor U5963 (N_5963,N_2888,N_3761);
or U5964 (N_5964,N_2561,N_3256);
or U5965 (N_5965,N_3173,N_3540);
and U5966 (N_5966,N_2590,N_2723);
nand U5967 (N_5967,N_2415,N_3118);
nand U5968 (N_5968,N_2869,N_2893);
nor U5969 (N_5969,N_2817,N_2978);
or U5970 (N_5970,N_3060,N_3164);
or U5971 (N_5971,N_3155,N_2525);
nor U5972 (N_5972,N_2532,N_3284);
or U5973 (N_5973,N_2183,N_2479);
nand U5974 (N_5974,N_3816,N_3350);
and U5975 (N_5975,N_3237,N_3155);
or U5976 (N_5976,N_3095,N_2513);
nand U5977 (N_5977,N_3973,N_3769);
nor U5978 (N_5978,N_2744,N_2412);
and U5979 (N_5979,N_3265,N_2463);
nand U5980 (N_5980,N_3567,N_2593);
and U5981 (N_5981,N_2689,N_3069);
xnor U5982 (N_5982,N_2490,N_2990);
and U5983 (N_5983,N_2867,N_3612);
nor U5984 (N_5984,N_2355,N_3649);
nor U5985 (N_5985,N_2087,N_2567);
xnor U5986 (N_5986,N_2488,N_3313);
or U5987 (N_5987,N_2483,N_3201);
or U5988 (N_5988,N_3803,N_3150);
and U5989 (N_5989,N_2509,N_3784);
and U5990 (N_5990,N_2464,N_2813);
and U5991 (N_5991,N_2869,N_2659);
nor U5992 (N_5992,N_2467,N_2799);
and U5993 (N_5993,N_3567,N_2087);
nor U5994 (N_5994,N_2295,N_2864);
or U5995 (N_5995,N_2746,N_3189);
or U5996 (N_5996,N_2872,N_3747);
nand U5997 (N_5997,N_2498,N_2353);
nor U5998 (N_5998,N_3391,N_3817);
nand U5999 (N_5999,N_3089,N_2971);
or U6000 (N_6000,N_4364,N_5373);
and U6001 (N_6001,N_5809,N_5938);
or U6002 (N_6002,N_5076,N_5648);
nor U6003 (N_6003,N_4637,N_5299);
and U6004 (N_6004,N_4764,N_4942);
or U6005 (N_6005,N_5978,N_5724);
nand U6006 (N_6006,N_5031,N_5107);
nand U6007 (N_6007,N_4297,N_4019);
or U6008 (N_6008,N_4218,N_5420);
or U6009 (N_6009,N_4562,N_4514);
nand U6010 (N_6010,N_5423,N_4228);
and U6011 (N_6011,N_4099,N_5923);
or U6012 (N_6012,N_5541,N_5224);
or U6013 (N_6013,N_4648,N_5689);
nor U6014 (N_6014,N_4940,N_4187);
nor U6015 (N_6015,N_5879,N_4699);
xnor U6016 (N_6016,N_5343,N_5170);
nand U6017 (N_6017,N_5590,N_4947);
nor U6018 (N_6018,N_4663,N_4917);
and U6019 (N_6019,N_4118,N_4496);
xnor U6020 (N_6020,N_4376,N_4189);
nor U6021 (N_6021,N_5804,N_5968);
nand U6022 (N_6022,N_4055,N_4200);
and U6023 (N_6023,N_5433,N_5402);
nor U6024 (N_6024,N_5655,N_5412);
and U6025 (N_6025,N_5647,N_4698);
or U6026 (N_6026,N_5187,N_5759);
and U6027 (N_6027,N_5302,N_5554);
and U6028 (N_6028,N_4175,N_4421);
xnor U6029 (N_6029,N_4874,N_4669);
xnor U6030 (N_6030,N_4614,N_4989);
xnor U6031 (N_6031,N_4929,N_5900);
or U6032 (N_6032,N_4095,N_5816);
or U6033 (N_6033,N_4073,N_4380);
nand U6034 (N_6034,N_4239,N_5979);
nand U6035 (N_6035,N_5404,N_4120);
or U6036 (N_6036,N_5853,N_4913);
xor U6037 (N_6037,N_4456,N_4918);
or U6038 (N_6038,N_5636,N_4110);
or U6039 (N_6039,N_4369,N_4167);
nand U6040 (N_6040,N_4078,N_5767);
nand U6041 (N_6041,N_4279,N_5045);
or U6042 (N_6042,N_5068,N_5265);
xor U6043 (N_6043,N_5521,N_5523);
nor U6044 (N_6044,N_5162,N_5635);
or U6045 (N_6045,N_4311,N_4492);
and U6046 (N_6046,N_5277,N_5966);
nand U6047 (N_6047,N_5101,N_5425);
and U6048 (N_6048,N_4158,N_5323);
nand U6049 (N_6049,N_5610,N_4748);
or U6050 (N_6050,N_4464,N_4604);
nand U6051 (N_6051,N_5563,N_5390);
nor U6052 (N_6052,N_4815,N_5247);
nor U6053 (N_6053,N_4611,N_4309);
or U6054 (N_6054,N_5972,N_4303);
nor U6055 (N_6055,N_5232,N_5918);
xor U6056 (N_6056,N_5217,N_5686);
nand U6057 (N_6057,N_5559,N_4636);
or U6058 (N_6058,N_4792,N_5942);
or U6059 (N_6059,N_5450,N_5629);
or U6060 (N_6060,N_5890,N_5119);
or U6061 (N_6061,N_4139,N_5836);
nor U6062 (N_6062,N_5266,N_4635);
xor U6063 (N_6063,N_4084,N_4671);
xnor U6064 (N_6064,N_5441,N_5077);
nor U6065 (N_6065,N_4028,N_5043);
or U6066 (N_6066,N_4922,N_4825);
or U6067 (N_6067,N_4439,N_5086);
nand U6068 (N_6068,N_4463,N_4164);
nor U6069 (N_6069,N_4147,N_4951);
xor U6070 (N_6070,N_5271,N_5270);
nor U6071 (N_6071,N_4616,N_4857);
xor U6072 (N_6072,N_5062,N_4363);
nor U6073 (N_6073,N_5719,N_5651);
nor U6074 (N_6074,N_4871,N_5274);
or U6075 (N_6075,N_4282,N_5106);
nor U6076 (N_6076,N_5051,N_4255);
xor U6077 (N_6077,N_5079,N_5811);
nand U6078 (N_6078,N_4000,N_5206);
and U6079 (N_6079,N_4948,N_5919);
and U6080 (N_6080,N_5887,N_5478);
or U6081 (N_6081,N_5933,N_5452);
nor U6082 (N_6082,N_4711,N_4739);
or U6083 (N_6083,N_5906,N_4331);
nor U6084 (N_6084,N_4783,N_4687);
xnor U6085 (N_6085,N_5824,N_5133);
xor U6086 (N_6086,N_5418,N_4100);
nor U6087 (N_6087,N_4306,N_5771);
nor U6088 (N_6088,N_4640,N_5307);
nand U6089 (N_6089,N_4036,N_4564);
or U6090 (N_6090,N_4932,N_4257);
and U6091 (N_6091,N_5155,N_4325);
nand U6092 (N_6092,N_4862,N_5931);
nand U6093 (N_6093,N_4707,N_5607);
and U6094 (N_6094,N_5673,N_4323);
nor U6095 (N_6095,N_4312,N_4447);
nand U6096 (N_6096,N_4029,N_4859);
or U6097 (N_6097,N_5982,N_5503);
xor U6098 (N_6098,N_5118,N_5838);
xnor U6099 (N_6099,N_5616,N_4438);
xor U6100 (N_6100,N_4559,N_5877);
nor U6101 (N_6101,N_4620,N_4004);
nand U6102 (N_6102,N_5710,N_4659);
and U6103 (N_6103,N_5524,N_4983);
nor U6104 (N_6104,N_5235,N_4751);
or U6105 (N_6105,N_5231,N_4881);
nand U6106 (N_6106,N_5281,N_5336);
and U6107 (N_6107,N_5320,N_4109);
nor U6108 (N_6108,N_4544,N_4465);
xnor U6109 (N_6109,N_4225,N_5504);
nand U6110 (N_6110,N_5508,N_4488);
xnor U6111 (N_6111,N_5160,N_5226);
nor U6112 (N_6112,N_5246,N_4893);
nand U6113 (N_6113,N_4161,N_4368);
nor U6114 (N_6114,N_5069,N_5659);
or U6115 (N_6115,N_5352,N_4144);
xor U6116 (N_6116,N_4710,N_5749);
xnor U6117 (N_6117,N_4808,N_5248);
nor U6118 (N_6118,N_5748,N_5184);
and U6119 (N_6119,N_4322,N_5908);
and U6120 (N_6120,N_5324,N_4966);
or U6121 (N_6121,N_4641,N_5755);
and U6122 (N_6122,N_5500,N_4487);
nand U6123 (N_6123,N_4915,N_4720);
or U6124 (N_6124,N_4525,N_5483);
or U6125 (N_6125,N_5194,N_5993);
nand U6126 (N_6126,N_5568,N_5708);
nand U6127 (N_6127,N_5196,N_5734);
nand U6128 (N_6128,N_4081,N_4508);
and U6129 (N_6129,N_4778,N_4280);
and U6130 (N_6130,N_5571,N_4191);
nor U6131 (N_6131,N_4018,N_5063);
xnor U6132 (N_6132,N_4264,N_4682);
or U6133 (N_6133,N_4931,N_5499);
and U6134 (N_6134,N_5581,N_5419);
nor U6135 (N_6135,N_4262,N_5191);
or U6136 (N_6136,N_4160,N_5589);
xor U6137 (N_6137,N_5863,N_5641);
nor U6138 (N_6138,N_4259,N_5289);
xor U6139 (N_6139,N_4872,N_5388);
nor U6140 (N_6140,N_5800,N_4540);
nor U6141 (N_6141,N_5596,N_4198);
nand U6142 (N_6142,N_4043,N_4895);
and U6143 (N_6143,N_4665,N_4088);
and U6144 (N_6144,N_4761,N_5300);
xnor U6145 (N_6145,N_5652,N_4460);
or U6146 (N_6146,N_5986,N_4093);
and U6147 (N_6147,N_5383,N_4241);
xor U6148 (N_6148,N_4765,N_5866);
and U6149 (N_6149,N_4361,N_5539);
nor U6150 (N_6150,N_4847,N_5858);
and U6151 (N_6151,N_5766,N_4396);
and U6152 (N_6152,N_4375,N_4926);
nand U6153 (N_6153,N_4405,N_5021);
xor U6154 (N_6154,N_4401,N_5886);
xnor U6155 (N_6155,N_5762,N_4258);
xor U6156 (N_6156,N_5737,N_4071);
or U6157 (N_6157,N_5867,N_5746);
or U6158 (N_6158,N_4089,N_5127);
nor U6159 (N_6159,N_5882,N_4981);
xor U6160 (N_6160,N_4169,N_4359);
or U6161 (N_6161,N_4417,N_4468);
and U6162 (N_6162,N_5462,N_5860);
and U6163 (N_6163,N_4811,N_5244);
nand U6164 (N_6164,N_5309,N_5612);
nor U6165 (N_6165,N_4290,N_4656);
nand U6166 (N_6166,N_4680,N_4888);
nand U6167 (N_6167,N_5535,N_5620);
xnor U6168 (N_6168,N_4386,N_4840);
xnor U6169 (N_6169,N_5445,N_4197);
nor U6170 (N_6170,N_5959,N_5262);
xnor U6171 (N_6171,N_5774,N_4585);
nand U6172 (N_6172,N_4092,N_5338);
or U6173 (N_6173,N_5472,N_4580);
xor U6174 (N_6174,N_5609,N_4069);
nand U6175 (N_6175,N_5492,N_4556);
nand U6176 (N_6176,N_4494,N_4768);
nor U6177 (N_6177,N_5213,N_4830);
nand U6178 (N_6178,N_4434,N_5028);
nor U6179 (N_6179,N_4343,N_4987);
nand U6180 (N_6180,N_4121,N_4633);
or U6181 (N_6181,N_5456,N_4042);
or U6182 (N_6182,N_4621,N_5185);
nand U6183 (N_6183,N_4291,N_4355);
xnor U6184 (N_6184,N_4171,N_4701);
or U6185 (N_6185,N_5964,N_5792);
xnor U6186 (N_6186,N_5741,N_5256);
nand U6187 (N_6187,N_5066,N_5484);
nand U6188 (N_6188,N_5789,N_4988);
or U6189 (N_6189,N_5476,N_5742);
or U6190 (N_6190,N_4319,N_5178);
nor U6191 (N_6191,N_5208,N_5556);
nor U6192 (N_6192,N_4860,N_4523);
and U6193 (N_6193,N_4342,N_4798);
nor U6194 (N_6194,N_4208,N_5778);
and U6195 (N_6195,N_4841,N_4923);
and U6196 (N_6196,N_4021,N_4406);
or U6197 (N_6197,N_5382,N_4246);
nor U6198 (N_6198,N_5772,N_4469);
nand U6199 (N_6199,N_4300,N_4676);
xnor U6200 (N_6200,N_4195,N_5053);
or U6201 (N_6201,N_4662,N_4125);
nand U6202 (N_6202,N_5874,N_4425);
nand U6203 (N_6203,N_5228,N_5555);
nor U6204 (N_6204,N_4688,N_5627);
xnor U6205 (N_6205,N_5082,N_4743);
nor U6206 (N_6206,N_4480,N_5050);
or U6207 (N_6207,N_5192,N_4443);
nor U6208 (N_6208,N_4479,N_4172);
nand U6209 (N_6209,N_5552,N_5828);
nand U6210 (N_6210,N_5429,N_5222);
and U6211 (N_6211,N_5997,N_4301);
nor U6212 (N_6212,N_5143,N_5236);
xor U6213 (N_6213,N_5061,N_4672);
nand U6214 (N_6214,N_4563,N_4009);
nand U6215 (N_6215,N_5952,N_4617);
nor U6216 (N_6216,N_4423,N_4943);
and U6217 (N_6217,N_5670,N_5723);
xor U6218 (N_6218,N_5894,N_5657);
and U6219 (N_6219,N_4327,N_4212);
nand U6220 (N_6220,N_4738,N_4070);
nand U6221 (N_6221,N_5976,N_4236);
nand U6222 (N_6222,N_4788,N_4470);
nor U6223 (N_6223,N_5333,N_5448);
or U6224 (N_6224,N_4113,N_4952);
and U6225 (N_6225,N_4415,N_4557);
nand U6226 (N_6226,N_5891,N_5850);
xor U6227 (N_6227,N_5012,N_4111);
nand U6228 (N_6228,N_5873,N_5884);
and U6229 (N_6229,N_4571,N_5533);
xnor U6230 (N_6230,N_4861,N_5202);
xnor U6231 (N_6231,N_5920,N_5344);
nand U6232 (N_6232,N_4769,N_4047);
nand U6233 (N_6233,N_5696,N_5594);
nand U6234 (N_6234,N_5732,N_5743);
nor U6235 (N_6235,N_4873,N_4285);
nor U6236 (N_6236,N_4186,N_5714);
or U6237 (N_6237,N_5036,N_4734);
and U6238 (N_6238,N_5415,N_5384);
nand U6239 (N_6239,N_4424,N_4305);
or U6240 (N_6240,N_4579,N_5989);
nand U6241 (N_6241,N_4404,N_4346);
or U6242 (N_6242,N_5437,N_5457);
nand U6243 (N_6243,N_4308,N_4249);
nand U6244 (N_6244,N_5080,N_5955);
nand U6245 (N_6245,N_5164,N_5219);
and U6246 (N_6246,N_4281,N_4837);
nand U6247 (N_6247,N_5507,N_4289);
or U6248 (N_6248,N_4276,N_4130);
xor U6249 (N_6249,N_4834,N_4646);
nor U6250 (N_6250,N_5869,N_5180);
xnor U6251 (N_6251,N_5532,N_4786);
nor U6252 (N_6252,N_5864,N_4997);
xnor U6253 (N_6253,N_4967,N_5843);
or U6254 (N_6254,N_5435,N_4668);
and U6255 (N_6255,N_5371,N_4541);
nand U6256 (N_6256,N_5994,N_4753);
xnor U6257 (N_6257,N_4328,N_5971);
nor U6258 (N_6258,N_4863,N_4483);
and U6259 (N_6259,N_4724,N_4950);
nor U6260 (N_6260,N_4025,N_4221);
or U6261 (N_6261,N_4524,N_4341);
or U6262 (N_6262,N_5146,N_5859);
nor U6263 (N_6263,N_4429,N_5254);
xor U6264 (N_6264,N_5988,N_5760);
and U6265 (N_6265,N_4793,N_4574);
and U6266 (N_6266,N_5209,N_5842);
and U6267 (N_6267,N_5125,N_4677);
or U6268 (N_6268,N_5845,N_5930);
nor U6269 (N_6269,N_5372,N_4351);
nand U6270 (N_6270,N_4876,N_5453);
and U6271 (N_6271,N_5168,N_4419);
xor U6272 (N_6272,N_5094,N_5349);
xnor U6273 (N_6273,N_5706,N_5642);
and U6274 (N_6274,N_5121,N_4972);
nor U6275 (N_6275,N_5932,N_4575);
nand U6276 (N_6276,N_5661,N_5288);
and U6277 (N_6277,N_4002,N_4750);
nand U6278 (N_6278,N_4498,N_4461);
nor U6279 (N_6279,N_4824,N_4740);
nand U6280 (N_6280,N_4708,N_5833);
and U6281 (N_6281,N_4884,N_4486);
nand U6282 (N_6282,N_5872,N_4762);
nand U6283 (N_6283,N_4268,N_4274);
nand U6284 (N_6284,N_5334,N_5560);
xor U6285 (N_6285,N_5378,N_4296);
and U6286 (N_6286,N_4827,N_5922);
or U6287 (N_6287,N_5468,N_5455);
xnor U6288 (N_6288,N_4210,N_4394);
xnor U6289 (N_6289,N_5314,N_5322);
or U6290 (N_6290,N_5399,N_5510);
or U6291 (N_6291,N_5350,N_4887);
or U6292 (N_6292,N_5097,N_4866);
and U6293 (N_6293,N_4691,N_5411);
nand U6294 (N_6294,N_4155,N_4800);
and U6295 (N_6295,N_4377,N_5493);
or U6296 (N_6296,N_5572,N_5176);
and U6297 (N_6297,N_4224,N_5301);
or U6298 (N_6298,N_4057,N_4048);
and U6299 (N_6299,N_4014,N_5034);
nand U6300 (N_6300,N_4543,N_4576);
or U6301 (N_6301,N_5898,N_4956);
nand U6302 (N_6302,N_4911,N_5924);
nand U6303 (N_6303,N_4485,N_4512);
or U6304 (N_6304,N_4222,N_5148);
and U6305 (N_6305,N_5611,N_5934);
nand U6306 (N_6306,N_4610,N_4232);
xnor U6307 (N_6307,N_5156,N_4817);
nand U6308 (N_6308,N_5190,N_4506);
xnor U6309 (N_6309,N_4759,N_5907);
and U6310 (N_6310,N_5495,N_4696);
xnor U6311 (N_6311,N_5605,N_4642);
xnor U6312 (N_6312,N_4085,N_5841);
nor U6313 (N_6313,N_4234,N_5057);
xor U6314 (N_6314,N_4420,N_4944);
nand U6315 (N_6315,N_5750,N_5764);
xor U6316 (N_6316,N_4153,N_4385);
xor U6317 (N_6317,N_4962,N_4619);
nor U6318 (N_6318,N_5779,N_4476);
nand U6319 (N_6319,N_5812,N_5599);
xor U6320 (N_6320,N_4307,N_5946);
nand U6321 (N_6321,N_5392,N_5451);
or U6322 (N_6322,N_5279,N_5704);
xnor U6323 (N_6323,N_5022,N_4735);
or U6324 (N_6324,N_5188,N_5114);
nor U6325 (N_6325,N_4204,N_4038);
or U6326 (N_6326,N_4630,N_4584);
and U6327 (N_6327,N_4702,N_5081);
and U6328 (N_6328,N_5065,N_4521);
and U6329 (N_6329,N_4201,N_4194);
nand U6330 (N_6330,N_4607,N_4174);
nand U6331 (N_6331,N_4627,N_4921);
xnor U6332 (N_6332,N_5072,N_5780);
nand U6333 (N_6333,N_4026,N_4910);
and U6334 (N_6334,N_5332,N_5166);
and U6335 (N_6335,N_4062,N_4503);
nor U6336 (N_6336,N_5027,N_5130);
nor U6337 (N_6337,N_5911,N_5409);
or U6338 (N_6338,N_5707,N_5578);
or U6339 (N_6339,N_4454,N_4779);
xor U6340 (N_6340,N_4013,N_5600);
xor U6341 (N_6341,N_4728,N_4213);
xor U6342 (N_6342,N_5870,N_5788);
xnor U6343 (N_6343,N_4304,N_5104);
nor U6344 (N_6344,N_5857,N_5664);
xnor U6345 (N_6345,N_4250,N_5295);
xnor U6346 (N_6346,N_4226,N_5698);
xnor U6347 (N_6347,N_5085,N_5515);
xor U6348 (N_6348,N_5676,N_5024);
xnor U6349 (N_6349,N_4517,N_4713);
and U6350 (N_6350,N_4820,N_5912);
nand U6351 (N_6351,N_4409,N_4853);
nand U6352 (N_6352,N_4678,N_5049);
and U6353 (N_6353,N_5834,N_5396);
xnor U6354 (N_6354,N_5312,N_4252);
nand U6355 (N_6355,N_4546,N_4106);
xnor U6356 (N_6356,N_4313,N_5167);
or U6357 (N_6357,N_5327,N_4039);
nand U6358 (N_6358,N_4017,N_4030);
nor U6359 (N_6359,N_5849,N_4810);
or U6360 (N_6360,N_4934,N_4237);
xnor U6361 (N_6361,N_4657,N_5626);
or U6362 (N_6362,N_4833,N_4027);
nand U6363 (N_6363,N_4963,N_5356);
or U6364 (N_6364,N_5856,N_5880);
nand U6365 (N_6365,N_4372,N_5365);
xnor U6366 (N_6366,N_4985,N_4076);
and U6367 (N_6367,N_5726,N_4651);
xor U6368 (N_6368,N_4003,N_5267);
or U6369 (N_6369,N_4206,N_5210);
nor U6370 (N_6370,N_5929,N_5407);
xor U6371 (N_6371,N_4216,N_4565);
xnor U6372 (N_6372,N_5443,N_5868);
nand U6373 (N_6373,N_5678,N_4970);
nor U6374 (N_6374,N_4535,N_5374);
and U6375 (N_6375,N_5585,N_5434);
nor U6376 (N_6376,N_5969,N_5264);
nor U6377 (N_6377,N_4653,N_5163);
nor U6378 (N_6378,N_5477,N_5212);
nand U6379 (N_6379,N_4882,N_5351);
and U6380 (N_6380,N_5292,N_5649);
and U6381 (N_6381,N_4267,N_5528);
nand U6382 (N_6382,N_4270,N_4717);
nor U6383 (N_6383,N_5394,N_5199);
nand U6384 (N_6384,N_5278,N_4462);
nand U6385 (N_6385,N_5353,N_4570);
or U6386 (N_6386,N_5697,N_5040);
nor U6387 (N_6387,N_4080,N_5318);
or U6388 (N_6388,N_4482,N_5020);
nor U6389 (N_6389,N_4054,N_5367);
and U6390 (N_6390,N_4612,N_4745);
xnor U6391 (N_6391,N_4284,N_4338);
nor U6392 (N_6392,N_5709,N_5335);
and U6393 (N_6393,N_5927,N_5840);
xnor U6394 (N_6394,N_4340,N_5389);
or U6395 (N_6395,N_4097,N_5397);
nor U6396 (N_6396,N_4407,N_4266);
nor U6397 (N_6397,N_5469,N_5144);
or U6398 (N_6398,N_5103,N_5848);
xnor U6399 (N_6399,N_4230,N_5825);
xnor U6400 (N_6400,N_5925,N_4597);
nand U6401 (N_6401,N_4758,N_5177);
nand U6402 (N_6402,N_5340,N_5223);
or U6403 (N_6403,N_5449,N_4141);
and U6404 (N_6404,N_4977,N_5757);
or U6405 (N_6405,N_4528,N_5249);
and U6406 (N_6406,N_4392,N_5506);
nor U6407 (N_6407,N_5093,N_4945);
or U6408 (N_6408,N_5181,N_4165);
or U6409 (N_6409,N_4594,N_5883);
or U6410 (N_6410,N_5048,N_5835);
xor U6411 (N_6411,N_4927,N_4791);
nand U6412 (N_6412,N_5403,N_5214);
nand U6413 (N_6413,N_4723,N_4511);
or U6414 (N_6414,N_5878,N_4686);
nand U6415 (N_6415,N_4431,N_5613);
or U6416 (N_6416,N_4821,N_5820);
nand U6417 (N_6417,N_5534,N_5663);
nor U6418 (N_6418,N_5035,N_4532);
nor U6419 (N_6419,N_5525,N_5428);
and U6420 (N_6420,N_5775,N_4032);
nand U6421 (N_6421,N_5380,N_5470);
or U6422 (N_6422,N_4858,N_4384);
or U6423 (N_6423,N_5574,N_5783);
and U6424 (N_6424,N_4615,N_4879);
nand U6425 (N_6425,N_4205,N_4321);
xor U6426 (N_6426,N_4553,N_5639);
and U6427 (N_6427,N_5442,N_4244);
and U6428 (N_6428,N_5827,N_4441);
nand U6429 (N_6429,N_4561,N_5297);
nor U6430 (N_6430,N_4435,N_5579);
nand U6431 (N_6431,N_5044,N_4819);
xor U6432 (N_6432,N_5561,N_5668);
nor U6433 (N_6433,N_4041,N_4590);
and U6434 (N_6434,N_4248,N_5808);
nor U6435 (N_6435,N_5728,N_5718);
and U6436 (N_6436,N_5691,N_4173);
and U6437 (N_6437,N_4133,N_5893);
nor U6438 (N_6438,N_4243,N_5667);
nor U6439 (N_6439,N_5796,N_5003);
or U6440 (N_6440,N_4555,N_5137);
or U6441 (N_6441,N_5830,N_4362);
and U6442 (N_6442,N_5716,N_4196);
nor U6443 (N_6443,N_4192,N_5926);
nor U6444 (N_6444,N_4776,N_4516);
and U6445 (N_6445,N_4864,N_5122);
xor U6446 (N_6446,N_4684,N_5799);
xnor U6447 (N_6447,N_4716,N_4889);
or U6448 (N_6448,N_4763,N_4644);
nor U6449 (N_6449,N_4567,N_4854);
and U6450 (N_6450,N_5817,N_5273);
xor U6451 (N_6451,N_4430,N_5823);
nand U6452 (N_6452,N_4885,N_5060);
or U6453 (N_6453,N_5564,N_5348);
xnor U6454 (N_6454,N_5471,N_4269);
or U6455 (N_6455,N_5009,N_4356);
and U6456 (N_6456,N_5406,N_4693);
or U6457 (N_6457,N_4256,N_4709);
and U6458 (N_6458,N_4867,N_4497);
nand U6459 (N_6459,N_5680,N_4625);
or U6460 (N_6460,N_4601,N_5095);
nand U6461 (N_6461,N_5987,N_4427);
and U6462 (N_6462,N_5730,N_4245);
or U6463 (N_6463,N_4605,N_5328);
and U6464 (N_6464,N_5364,N_5790);
nand U6465 (N_6465,N_4531,N_4181);
and U6466 (N_6466,N_5509,N_5105);
nor U6467 (N_6467,N_4022,N_5801);
nor U6468 (N_6468,N_4755,N_4822);
nor U6469 (N_6469,N_5479,N_5111);
nor U6470 (N_6470,N_5522,N_5132);
nor U6471 (N_6471,N_5837,N_4298);
nand U6472 (N_6472,N_5090,N_5628);
nand U6473 (N_6473,N_5832,N_4148);
nor U6474 (N_6474,N_4957,N_4001);
xnor U6475 (N_6475,N_5366,N_4202);
nor U6476 (N_6476,N_5444,N_4850);
nor U6477 (N_6477,N_4675,N_5475);
and U6478 (N_6478,N_4623,N_5359);
nand U6479 (N_6479,N_4220,N_5237);
nand U6480 (N_6480,N_4715,N_4823);
and U6481 (N_6481,N_5276,N_5179);
xor U6482 (N_6482,N_4108,N_4844);
nor U6483 (N_6483,N_5290,N_4383);
nand U6484 (N_6484,N_4112,N_4935);
xnor U6485 (N_6485,N_4332,N_4378);
nor U6486 (N_6486,N_4122,N_5058);
nor U6487 (N_6487,N_4414,N_4527);
or U6488 (N_6488,N_5553,N_4333);
nor U6489 (N_6489,N_5227,N_4102);
or U6490 (N_6490,N_5075,N_4064);
nand U6491 (N_6491,N_5733,N_5683);
nand U6492 (N_6492,N_5438,N_5174);
nand U6493 (N_6493,N_5029,N_4442);
or U6494 (N_6494,N_4869,N_5195);
nor U6495 (N_6495,N_4647,N_5255);
nand U6496 (N_6496,N_4566,N_4596);
or U6497 (N_6497,N_4919,N_4519);
and U6498 (N_6498,N_4832,N_5129);
nor U6499 (N_6499,N_4638,N_5542);
nand U6500 (N_6500,N_4606,N_5238);
or U6501 (N_6501,N_5124,N_5722);
nand U6502 (N_6502,N_5645,N_5234);
nor U6503 (N_6503,N_4548,N_4458);
and U6504 (N_6504,N_5099,N_4134);
nor U6505 (N_6505,N_4538,N_4731);
or U6506 (N_6506,N_4166,N_5291);
or U6507 (N_6507,N_4838,N_4316);
nor U6508 (N_6508,N_4537,N_5720);
nand U6509 (N_6509,N_4398,N_5995);
or U6510 (N_6510,N_4880,N_4354);
or U6511 (N_6511,N_5606,N_5851);
xor U6512 (N_6512,N_4986,N_4939);
or U6513 (N_6513,N_4500,N_5703);
or U6514 (N_6514,N_4809,N_4598);
or U6515 (N_6515,N_5614,N_4547);
nand U6516 (N_6516,N_5424,N_5745);
nand U6517 (N_6517,N_4550,N_5253);
nand U6518 (N_6518,N_5401,N_5753);
or U6519 (N_6519,N_5393,N_5892);
nor U6520 (N_6520,N_4373,N_5282);
or U6521 (N_6521,N_5379,N_4586);
xor U6522 (N_6522,N_5604,N_4790);
nand U6523 (N_6523,N_5154,N_4079);
or U6524 (N_6524,N_4413,N_5865);
xor U6525 (N_6525,N_4335,N_5803);
nand U6526 (N_6526,N_5109,N_4773);
nand U6527 (N_6527,N_5646,N_4756);
and U6528 (N_6528,N_5829,N_4802);
or U6529 (N_6529,N_5064,N_5313);
or U6530 (N_6530,N_5183,N_4906);
nor U6531 (N_6531,N_5777,N_4536);
nand U6532 (N_6532,N_4909,N_4374);
and U6533 (N_6533,N_5608,N_4916);
and U6534 (N_6534,N_4992,N_4271);
or U6535 (N_6535,N_4408,N_4742);
xnor U6536 (N_6536,N_5315,N_4445);
nand U6537 (N_6537,N_4034,N_5377);
xor U6538 (N_6538,N_4053,N_5007);
and U6539 (N_6539,N_5557,N_5677);
or U6540 (N_6540,N_4904,N_4329);
nand U6541 (N_6541,N_5985,N_5632);
nor U6542 (N_6542,N_4704,N_5347);
nand U6543 (N_6543,N_5763,N_4679);
and U6544 (N_6544,N_4140,N_4273);
nand U6545 (N_6545,N_4897,N_5501);
and U6546 (N_6546,N_4722,N_4784);
and U6547 (N_6547,N_4358,N_4685);
nor U6548 (N_6548,N_5233,N_4733);
or U6549 (N_6549,N_4578,N_4499);
xor U6550 (N_6550,N_4422,N_5640);
nand U6551 (N_6551,N_5173,N_4689);
and U6552 (N_6552,N_4539,N_5120);
nor U6553 (N_6553,N_4628,N_4357);
nand U6554 (N_6554,N_4754,N_5427);
xor U6555 (N_6555,N_4242,N_5701);
and U6556 (N_6556,N_5795,N_5376);
xor U6557 (N_6557,N_4104,N_5660);
and U6558 (N_6558,N_4645,N_5145);
nand U6559 (N_6559,N_5055,N_5538);
and U6560 (N_6560,N_4851,N_4135);
or U6561 (N_6561,N_4466,N_5193);
and U6562 (N_6562,N_5806,N_4101);
xnor U6563 (N_6563,N_4278,N_5149);
and U6564 (N_6564,N_4275,N_4344);
and U6565 (N_6565,N_4115,N_5171);
nand U6566 (N_6566,N_4094,N_4182);
or U6567 (N_6567,N_5512,N_5046);
nand U6568 (N_6568,N_5592,N_4573);
nand U6569 (N_6569,N_4211,N_4955);
xnor U6570 (N_6570,N_4261,N_4116);
nor U6571 (N_6571,N_4016,N_5491);
xnor U6572 (N_6572,N_5684,N_4382);
nor U6573 (N_6573,N_4626,N_4162);
or U6574 (N_6574,N_5306,N_5134);
nand U6575 (N_6575,N_4011,N_4272);
xor U6576 (N_6576,N_4020,N_5567);
or U6577 (N_6577,N_5669,N_4787);
and U6578 (N_6578,N_4247,N_5439);
nand U6579 (N_6579,N_4912,N_4347);
nand U6580 (N_6580,N_5169,N_5071);
nor U6581 (N_6581,N_4785,N_5899);
xor U6582 (N_6582,N_5139,N_5293);
and U6583 (N_6583,N_5601,N_5126);
xor U6584 (N_6584,N_4444,N_4299);
nand U6585 (N_6585,N_5944,N_4719);
xor U6586 (N_6586,N_4156,N_4806);
or U6587 (N_6587,N_5474,N_4812);
nand U6588 (N_6588,N_4436,N_4450);
xnor U6589 (N_6589,N_4490,N_4217);
nor U6590 (N_6590,N_4365,N_5876);
or U6591 (N_6591,N_5844,N_4752);
nand U6592 (N_6592,N_5023,N_4288);
and U6593 (N_6593,N_5514,N_5765);
nand U6594 (N_6594,N_4856,N_4890);
nand U6595 (N_6595,N_5586,N_4969);
nand U6596 (N_6596,N_4868,N_4654);
nand U6597 (N_6597,N_5490,N_4658);
and U6598 (N_6598,N_4426,N_5935);
or U6599 (N_6599,N_4900,N_4072);
xor U6600 (N_6600,N_5440,N_4481);
xnor U6601 (N_6601,N_5702,N_5794);
nand U6602 (N_6602,N_4231,N_4082);
or U6603 (N_6603,N_4732,N_5569);
and U6604 (N_6604,N_5310,N_4599);
or U6605 (N_6605,N_4803,N_4741);
xor U6606 (N_6606,N_4367,N_4352);
nand U6607 (N_6607,N_4433,N_4501);
nor U6608 (N_6608,N_4159,N_4513);
and U6609 (N_6609,N_4805,N_5381);
xor U6610 (N_6610,N_4128,N_5426);
or U6611 (N_6611,N_4814,N_5643);
and U6612 (N_6612,N_4664,N_4891);
xor U6613 (N_6613,N_4185,N_5537);
xor U6614 (N_6614,N_5740,N_5410);
or U6615 (N_6615,N_5681,N_4877);
and U6616 (N_6616,N_5624,N_5502);
or U6617 (N_6617,N_4801,N_5017);
and U6618 (N_6618,N_4994,N_5562);
xor U6619 (N_6619,N_5672,N_4350);
and U6620 (N_6620,N_5284,N_4475);
nor U6621 (N_6621,N_5625,N_4031);
nand U6622 (N_6622,N_5889,N_4520);
and U6623 (N_6623,N_4736,N_4366);
nor U6624 (N_6624,N_5298,N_5937);
and U6625 (N_6625,N_5446,N_4103);
and U6626 (N_6626,N_4697,N_5054);
nor U6627 (N_6627,N_5136,N_4632);
xnor U6628 (N_6628,N_4980,N_5621);
nor U6629 (N_6629,N_5067,N_5311);
and U6630 (N_6630,N_5413,N_5725);
nand U6631 (N_6631,N_4397,N_4170);
nor U6632 (N_6632,N_4924,N_5161);
nor U6633 (N_6633,N_5421,N_5862);
or U6634 (N_6634,N_5000,N_4471);
xor U6635 (N_6635,N_4154,N_5319);
nor U6636 (N_6636,N_4705,N_5947);
and U6637 (N_6637,N_5638,N_5516);
xor U6638 (N_6638,N_4953,N_5172);
nand U6639 (N_6639,N_5422,N_4600);
nor U6640 (N_6640,N_4770,N_5436);
nand U6641 (N_6641,N_4489,N_4473);
and U6642 (N_6642,N_5666,N_5631);
nand U6643 (N_6643,N_5797,N_4818);
and U6644 (N_6644,N_4725,N_5131);
or U6645 (N_6645,N_5305,N_5117);
nand U6646 (N_6646,N_4979,N_4149);
xor U6647 (N_6647,N_4995,N_5566);
or U6648 (N_6648,N_5387,N_4515);
or U6649 (N_6649,N_4075,N_5700);
or U6650 (N_6650,N_4855,N_4813);
and U6651 (N_6651,N_5432,N_4582);
or U6652 (N_6652,N_5822,N_4775);
nand U6653 (N_6653,N_4502,N_5744);
nand U6654 (N_6654,N_4894,N_5128);
and U6655 (N_6655,N_5654,N_4941);
and U6656 (N_6656,N_5417,N_4505);
xnor U6657 (N_6657,N_4703,N_5786);
nor U6658 (N_6658,N_4302,N_5715);
nor U6659 (N_6659,N_5074,N_4152);
xnor U6660 (N_6660,N_5368,N_4381);
and U6661 (N_6661,N_4846,N_4314);
nand U6662 (N_6662,N_5218,N_5595);
or U6663 (N_6663,N_4826,N_5326);
xor U6664 (N_6664,N_4591,N_5038);
nand U6665 (N_6665,N_4318,N_5904);
nand U6666 (N_6666,N_4176,N_4902);
nand U6667 (N_6667,N_4428,N_4843);
nand U6668 (N_6668,N_4015,N_5198);
and U6669 (N_6669,N_5826,N_5004);
and U6670 (N_6670,N_5650,N_4634);
nand U6671 (N_6671,N_5839,N_5220);
nand U6672 (N_6672,N_4360,N_4683);
and U6673 (N_6673,N_5461,N_4892);
or U6674 (N_6674,N_5182,N_5953);
nor U6675 (N_6675,N_5201,N_4936);
xnor U6676 (N_6676,N_5294,N_4549);
or U6677 (N_6677,N_4044,N_5819);
xor U6678 (N_6678,N_5263,N_5230);
and U6679 (N_6679,N_5550,N_4074);
and U6680 (N_6680,N_5984,N_4726);
nor U6681 (N_6681,N_5693,N_5496);
nand U6682 (N_6682,N_4008,N_5756);
xnor U6683 (N_6683,N_4993,N_5902);
nor U6684 (N_6684,N_4649,N_5945);
xnor U6685 (N_6685,N_4114,N_5013);
nor U6686 (N_6686,N_4068,N_5773);
or U6687 (N_6687,N_5921,N_5330);
nand U6688 (N_6688,N_5940,N_4694);
nor U6689 (N_6689,N_5304,N_4453);
and U6690 (N_6690,N_5480,N_5818);
nand U6691 (N_6691,N_5776,N_5486);
xnor U6692 (N_6692,N_5385,N_4005);
xnor U6693 (N_6693,N_5949,N_5967);
or U6694 (N_6694,N_4455,N_4807);
and U6695 (N_6695,N_4146,N_4251);
xor U6696 (N_6696,N_5317,N_5215);
nand U6697 (N_6697,N_4618,N_4035);
or U6698 (N_6698,N_5141,N_5497);
or U6699 (N_6699,N_4294,N_5588);
xnor U6700 (N_6700,N_5257,N_4865);
xor U6701 (N_6701,N_5735,N_5617);
or U6702 (N_6702,N_4348,N_5855);
nand U6703 (N_6703,N_4209,N_4457);
xor U6704 (N_6704,N_5980,N_4903);
or U6705 (N_6705,N_4105,N_4448);
or U6706 (N_6706,N_4930,N_5002);
and U6707 (N_6707,N_5369,N_5791);
nor U6708 (N_6708,N_5430,N_4849);
nor U6709 (N_6709,N_5768,N_5229);
or U6710 (N_6710,N_4012,N_4781);
xnor U6711 (N_6711,N_4353,N_5885);
or U6712 (N_6712,N_5159,N_5685);
nor U6713 (N_6713,N_5098,N_4292);
xor U6714 (N_6714,N_4418,N_5658);
or U6715 (N_6715,N_4179,N_5634);
or U6716 (N_6716,N_4828,N_5464);
or U6717 (N_6717,N_4077,N_4132);
xnor U6718 (N_6718,N_5758,N_4509);
or U6719 (N_6719,N_4551,N_5943);
nand U6720 (N_6720,N_5536,N_4238);
xnor U6721 (N_6721,N_5260,N_5807);
xnor U6722 (N_6722,N_4495,N_4899);
nor U6723 (N_6723,N_5951,N_4760);
xor U6724 (N_6724,N_4655,N_4388);
xor U6725 (N_6725,N_4737,N_5974);
and U6726 (N_6726,N_4193,N_4142);
nand U6727 (N_6727,N_5110,N_4706);
nor U6728 (N_6728,N_4049,N_4946);
nand U6729 (N_6729,N_4098,N_4451);
xor U6730 (N_6730,N_5991,N_5975);
nand U6731 (N_6731,N_5543,N_4789);
xnor U6732 (N_6732,N_5901,N_4661);
nor U6733 (N_6733,N_5821,N_5798);
and U6734 (N_6734,N_4660,N_5280);
and U6735 (N_6735,N_5705,N_4393);
xor U6736 (N_6736,N_5400,N_4937);
nor U6737 (N_6737,N_4650,N_4287);
xor U6738 (N_6738,N_5083,N_4123);
and U6739 (N_6739,N_5084,N_4718);
nand U6740 (N_6740,N_5674,N_4960);
nand U6741 (N_6741,N_4265,N_4233);
and U6742 (N_6742,N_4554,N_4229);
and U6743 (N_6743,N_5970,N_4336);
nor U6744 (N_6744,N_5513,N_4190);
nor U6745 (N_6745,N_4954,N_5042);
nor U6746 (N_6746,N_5583,N_5917);
nand U6747 (N_6747,N_4184,N_5998);
and U6748 (N_6748,N_4795,N_4767);
or U6749 (N_6749,N_4349,N_5001);
or U6750 (N_6750,N_5408,N_4587);
nor U6751 (N_6751,N_5150,N_4320);
xnor U6752 (N_6752,N_5360,N_4609);
nand U6753 (N_6753,N_4138,N_4157);
or U6754 (N_6754,N_5467,N_5679);
xor U6755 (N_6755,N_5895,N_4978);
and U6756 (N_6756,N_4207,N_4602);
nand U6757 (N_6757,N_5618,N_4700);
and U6758 (N_6758,N_5965,N_4324);
or U6759 (N_6759,N_5570,N_4050);
nand U6760 (N_6760,N_5630,N_4522);
or U6761 (N_6761,N_5016,N_5785);
xnor U6762 (N_6762,N_5241,N_5547);
nor U6763 (N_6763,N_5548,N_5573);
nand U6764 (N_6764,N_5329,N_4371);
xor U6765 (N_6765,N_5962,N_4033);
xnor U6766 (N_6766,N_4124,N_5688);
or U6767 (N_6767,N_5852,N_5342);
nor U6768 (N_6768,N_5540,N_5252);
nand U6769 (N_6769,N_5308,N_5591);
or U6770 (N_6770,N_5981,N_4389);
nand U6771 (N_6771,N_5622,N_5112);
nor U6772 (N_6772,N_4835,N_5903);
or U6773 (N_6773,N_5152,N_5914);
and U6774 (N_6774,N_4045,N_5088);
nor U6775 (N_6775,N_5100,N_4914);
xor U6776 (N_6776,N_5948,N_5473);
nand U6777 (N_6777,N_5511,N_4477);
and U6778 (N_6778,N_4452,N_4052);
nor U6779 (N_6779,N_4065,N_5018);
nand U6780 (N_6780,N_5361,N_4771);
or U6781 (N_6781,N_4958,N_4472);
nor U6782 (N_6782,N_5239,N_4572);
xor U6783 (N_6783,N_5203,N_4845);
nand U6784 (N_6784,N_4747,N_5089);
and U6785 (N_6785,N_4690,N_4478);
xor U6786 (N_6786,N_4474,N_4905);
or U6787 (N_6787,N_4777,N_5269);
nor U6788 (N_6788,N_4568,N_4560);
and U6789 (N_6789,N_5992,N_5251);
nor U6790 (N_6790,N_5370,N_5897);
nor U6791 (N_6791,N_4938,N_5793);
xnor U6792 (N_6792,N_5587,N_5983);
nand U6793 (N_6793,N_4326,N_5519);
nand U6794 (N_6794,N_4875,N_4558);
xor U6795 (N_6795,N_4334,N_4117);
nand U6796 (N_6796,N_4137,N_5070);
xnor U6797 (N_6797,N_5915,N_4976);
and U6798 (N_6798,N_5037,N_4526);
and U6799 (N_6799,N_5357,N_4010);
xnor U6800 (N_6800,N_5671,N_4673);
nor U6801 (N_6801,N_4518,N_4542);
nor U6802 (N_6802,N_4780,N_5488);
xnor U6803 (N_6803,N_5362,N_5287);
nand U6804 (N_6804,N_5135,N_4996);
nand U6805 (N_6805,N_5151,N_5517);
nor U6806 (N_6806,N_5675,N_4842);
nor U6807 (N_6807,N_4293,N_5682);
nand U6808 (N_6808,N_4240,N_5831);
nor U6809 (N_6809,N_5200,N_4975);
nor U6810 (N_6810,N_4143,N_4150);
xnor U6811 (N_6811,N_5165,N_4552);
and U6812 (N_6812,N_4949,N_5073);
xor U6813 (N_6813,N_5854,N_5754);
xnor U6814 (N_6814,N_5025,N_5142);
xor U6815 (N_6815,N_5339,N_5153);
and U6816 (N_6816,N_4593,N_5459);
or U6817 (N_6817,N_4446,N_4058);
nor U6818 (N_6818,N_4729,N_4991);
nor U6819 (N_6819,N_5363,N_5096);
nand U6820 (N_6820,N_4974,N_4848);
and U6821 (N_6821,N_5355,N_5551);
xnor U6822 (N_6822,N_4254,N_5345);
xor U6823 (N_6823,N_4712,N_5416);
or U6824 (N_6824,N_4545,N_4484);
nor U6825 (N_6825,N_5582,N_4188);
nand U6826 (N_6826,N_4046,N_4295);
or U6827 (N_6827,N_4390,N_4907);
or U6828 (N_6828,N_5999,N_5087);
xnor U6829 (N_6829,N_4920,N_5498);
nand U6830 (N_6830,N_4583,N_4595);
and U6831 (N_6831,N_4090,N_4253);
and U6832 (N_6832,N_5465,N_5494);
and U6833 (N_6833,N_4395,N_4883);
xnor U6834 (N_6834,N_4163,N_4345);
xor U6835 (N_6835,N_5936,N_5531);
and U6836 (N_6836,N_5713,N_5189);
nor U6837 (N_6837,N_4529,N_4639);
xor U6838 (N_6838,N_5447,N_4643);
xor U6839 (N_6839,N_5712,N_5653);
nand U6840 (N_6840,N_4569,N_4666);
nor U6841 (N_6841,N_4432,N_4534);
nand U6842 (N_6842,N_4925,N_5115);
nand U6843 (N_6843,N_4402,N_4577);
xnor U6844 (N_6844,N_5546,N_5175);
nand U6845 (N_6845,N_4749,N_5814);
and U6846 (N_6846,N_4964,N_4219);
nand U6847 (N_6847,N_4315,N_5259);
and U6848 (N_6848,N_5694,N_5738);
xor U6849 (N_6849,N_5205,N_5727);
nor U6850 (N_6850,N_4908,N_4852);
nand U6851 (N_6851,N_5736,N_5623);
and U6852 (N_6852,N_4831,N_5871);
and U6853 (N_6853,N_5019,N_4886);
nor U6854 (N_6854,N_4235,N_4933);
nor U6855 (N_6855,N_5815,N_4387);
nor U6856 (N_6856,N_4260,N_5977);
xnor U6857 (N_6857,N_4652,N_5558);
xnor U6858 (N_6858,N_5665,N_4797);
nand U6859 (N_6859,N_5875,N_5078);
nand U6860 (N_6860,N_4670,N_4227);
nor U6861 (N_6861,N_5928,N_5597);
and U6862 (N_6862,N_4379,N_4714);
nand U6863 (N_6863,N_5395,N_5990);
and U6864 (N_6864,N_5813,N_5913);
and U6865 (N_6865,N_5108,N_5781);
xnor U6866 (N_6866,N_5784,N_5354);
xnor U6867 (N_6867,N_5769,N_5950);
nor U6868 (N_6868,N_5261,N_4056);
or U6869 (N_6869,N_4493,N_4183);
nand U6870 (N_6870,N_5603,N_5526);
nand U6871 (N_6871,N_4674,N_5272);
and U6872 (N_6872,N_5905,N_4067);
or U6873 (N_6873,N_5041,N_4370);
and U6874 (N_6874,N_4040,N_5138);
nand U6875 (N_6875,N_5711,N_4695);
or U6876 (N_6876,N_5751,N_5140);
nand U6877 (N_6877,N_4178,N_5242);
nand U6878 (N_6878,N_4007,N_5909);
nand U6879 (N_6879,N_5296,N_4510);
or U6880 (N_6880,N_5739,N_4391);
xor U6881 (N_6881,N_4136,N_5458);
xor U6882 (N_6882,N_4998,N_5881);
nand U6883 (N_6883,N_5752,N_5157);
or U6884 (N_6884,N_4129,N_5575);
or U6885 (N_6885,N_4203,N_5963);
nand U6886 (N_6886,N_4263,N_5544);
nand U6887 (N_6887,N_4744,N_5530);
nor U6888 (N_6888,N_5033,N_5303);
nand U6889 (N_6889,N_5032,N_4507);
nand U6890 (N_6890,N_5285,N_4467);
or U6891 (N_6891,N_5466,N_4965);
or U6892 (N_6892,N_4412,N_5059);
nor U6893 (N_6893,N_4131,N_5954);
and U6894 (N_6894,N_5358,N_5092);
or U6895 (N_6895,N_5197,N_4727);
and U6896 (N_6896,N_5695,N_5102);
or U6897 (N_6897,N_5910,N_4024);
nor U6898 (N_6898,N_4410,N_4961);
xor U6899 (N_6899,N_5485,N_5598);
xnor U6900 (N_6900,N_5225,N_5846);
or U6901 (N_6901,N_4059,N_5602);
or U6902 (N_6902,N_5956,N_5030);
and U6903 (N_6903,N_4437,N_5123);
or U6904 (N_6904,N_5633,N_5221);
and U6905 (N_6905,N_5460,N_4816);
and U6906 (N_6906,N_5847,N_4624);
xnor U6907 (N_6907,N_5545,N_5250);
and U6908 (N_6908,N_4829,N_5325);
and U6909 (N_6909,N_5529,N_5337);
and U6910 (N_6910,N_4107,N_4721);
nand U6911 (N_6911,N_5482,N_4746);
nor U6912 (N_6912,N_5580,N_5576);
or U6913 (N_6913,N_5386,N_4530);
and U6914 (N_6914,N_4083,N_4794);
xnor U6915 (N_6915,N_5615,N_4681);
nand U6916 (N_6916,N_5916,N_5010);
and U6917 (N_6917,N_5286,N_5245);
nand U6918 (N_6918,N_5113,N_5960);
xnor U6919 (N_6919,N_4339,N_5147);
nor U6920 (N_6920,N_5398,N_5584);
xor U6921 (N_6921,N_4400,N_5268);
nand U6922 (N_6922,N_4667,N_5431);
nand U6923 (N_6923,N_4973,N_4928);
and U6924 (N_6924,N_4145,N_5644);
xnor U6925 (N_6925,N_5961,N_4613);
nand U6926 (N_6926,N_5692,N_4898);
xnor U6927 (N_6927,N_5805,N_5527);
and U6928 (N_6928,N_4215,N_5463);
and U6929 (N_6929,N_5015,N_4504);
nand U6930 (N_6930,N_4214,N_4411);
or U6931 (N_6931,N_5518,N_4061);
or U6932 (N_6932,N_4692,N_4199);
and U6933 (N_6933,N_5091,N_4839);
and U6934 (N_6934,N_4440,N_4990);
xnor U6935 (N_6935,N_5996,N_4459);
nor U6936 (N_6936,N_5731,N_4772);
and U6937 (N_6937,N_4774,N_5346);
or U6938 (N_6938,N_5391,N_4337);
nand U6939 (N_6939,N_5240,N_5204);
xnor U6940 (N_6940,N_4177,N_4971);
nor U6941 (N_6941,N_4416,N_5721);
and U6942 (N_6942,N_5116,N_4403);
xnor U6943 (N_6943,N_5577,N_5414);
or U6944 (N_6944,N_4757,N_5487);
nor U6945 (N_6945,N_4310,N_5699);
and U6946 (N_6946,N_5321,N_4982);
nor U6947 (N_6947,N_5687,N_4984);
xor U6948 (N_6948,N_4283,N_5973);
nor U6949 (N_6949,N_4180,N_4999);
nor U6950 (N_6950,N_5283,N_5939);
xor U6951 (N_6951,N_5405,N_5243);
nand U6952 (N_6952,N_4796,N_4959);
and U6953 (N_6953,N_5520,N_5761);
and U6954 (N_6954,N_4023,N_4870);
nor U6955 (N_6955,N_4631,N_4091);
and U6956 (N_6956,N_5047,N_4399);
xnor U6957 (N_6957,N_5958,N_5770);
nand U6958 (N_6958,N_4622,N_5052);
or U6959 (N_6959,N_4533,N_4730);
or U6960 (N_6960,N_5619,N_5565);
and U6961 (N_6961,N_4603,N_5747);
nor U6962 (N_6962,N_5810,N_5593);
nand U6963 (N_6963,N_4096,N_4782);
nor U6964 (N_6964,N_4449,N_4896);
xnor U6965 (N_6965,N_5341,N_5489);
or U6966 (N_6966,N_5896,N_5802);
and U6967 (N_6967,N_4168,N_4063);
xnor U6968 (N_6968,N_4629,N_5957);
nand U6969 (N_6969,N_5787,N_4086);
nor U6970 (N_6970,N_4060,N_4799);
and U6971 (N_6971,N_5331,N_4151);
xor U6972 (N_6972,N_5211,N_5454);
xnor U6973 (N_6973,N_5275,N_5216);
nor U6974 (N_6974,N_5505,N_4223);
and U6975 (N_6975,N_5549,N_5782);
xnor U6976 (N_6976,N_5005,N_5011);
and U6977 (N_6977,N_4127,N_4968);
nor U6978 (N_6978,N_5008,N_4317);
or U6979 (N_6979,N_4581,N_4491);
nand U6980 (N_6980,N_4836,N_4037);
or U6981 (N_6981,N_4286,N_5186);
or U6982 (N_6982,N_5717,N_5006);
and U6983 (N_6983,N_4592,N_4608);
nand U6984 (N_6984,N_5014,N_5375);
nand U6985 (N_6985,N_5056,N_5258);
or U6986 (N_6986,N_5729,N_4766);
nand U6987 (N_6987,N_4878,N_5656);
nor U6988 (N_6988,N_4277,N_4006);
nand U6989 (N_6989,N_4126,N_5207);
or U6990 (N_6990,N_5039,N_5662);
or U6991 (N_6991,N_4066,N_4051);
nand U6992 (N_6992,N_5158,N_4087);
and U6993 (N_6993,N_4119,N_4589);
and U6994 (N_6994,N_4901,N_4330);
xor U6995 (N_6995,N_4588,N_5316);
xnor U6996 (N_6996,N_5888,N_5690);
xnor U6997 (N_6997,N_5026,N_5481);
xnor U6998 (N_6998,N_5941,N_5861);
or U6999 (N_6999,N_4804,N_5637);
or U7000 (N_7000,N_5698,N_4736);
nor U7001 (N_7001,N_5196,N_5862);
xnor U7002 (N_7002,N_4360,N_4788);
xor U7003 (N_7003,N_4915,N_5303);
or U7004 (N_7004,N_5671,N_5442);
and U7005 (N_7005,N_5913,N_5877);
nand U7006 (N_7006,N_5253,N_5762);
or U7007 (N_7007,N_5600,N_5578);
nand U7008 (N_7008,N_5704,N_5258);
or U7009 (N_7009,N_4793,N_5682);
xnor U7010 (N_7010,N_5510,N_5015);
xnor U7011 (N_7011,N_4594,N_5616);
or U7012 (N_7012,N_5328,N_5922);
and U7013 (N_7013,N_4561,N_4849);
or U7014 (N_7014,N_4899,N_5602);
nor U7015 (N_7015,N_5827,N_5701);
nand U7016 (N_7016,N_4407,N_4920);
or U7017 (N_7017,N_5520,N_5236);
or U7018 (N_7018,N_5665,N_4496);
or U7019 (N_7019,N_4246,N_5305);
nor U7020 (N_7020,N_4399,N_5970);
nor U7021 (N_7021,N_4738,N_4764);
and U7022 (N_7022,N_5202,N_4370);
and U7023 (N_7023,N_4357,N_4711);
nand U7024 (N_7024,N_5781,N_4274);
or U7025 (N_7025,N_5690,N_4504);
xor U7026 (N_7026,N_5749,N_5048);
nand U7027 (N_7027,N_5787,N_5328);
nor U7028 (N_7028,N_4869,N_4718);
or U7029 (N_7029,N_4981,N_5946);
or U7030 (N_7030,N_4191,N_4022);
nand U7031 (N_7031,N_5388,N_4900);
nand U7032 (N_7032,N_4775,N_4630);
xnor U7033 (N_7033,N_4385,N_5381);
and U7034 (N_7034,N_5304,N_4643);
or U7035 (N_7035,N_5257,N_5464);
and U7036 (N_7036,N_5905,N_4812);
xnor U7037 (N_7037,N_4774,N_4008);
and U7038 (N_7038,N_4421,N_4689);
nand U7039 (N_7039,N_5750,N_5299);
xor U7040 (N_7040,N_4270,N_5284);
nand U7041 (N_7041,N_5938,N_5437);
and U7042 (N_7042,N_4515,N_4891);
xor U7043 (N_7043,N_5185,N_4482);
xor U7044 (N_7044,N_5284,N_5679);
nand U7045 (N_7045,N_4004,N_4102);
nor U7046 (N_7046,N_4600,N_4034);
nand U7047 (N_7047,N_5292,N_5831);
nor U7048 (N_7048,N_4856,N_4359);
nand U7049 (N_7049,N_4984,N_4459);
or U7050 (N_7050,N_5527,N_4770);
nor U7051 (N_7051,N_4850,N_5348);
or U7052 (N_7052,N_5423,N_5876);
nand U7053 (N_7053,N_4344,N_5900);
nand U7054 (N_7054,N_4535,N_5760);
xor U7055 (N_7055,N_4999,N_5332);
or U7056 (N_7056,N_4623,N_4738);
nand U7057 (N_7057,N_5756,N_5094);
nor U7058 (N_7058,N_4898,N_4630);
nand U7059 (N_7059,N_5576,N_4990);
xor U7060 (N_7060,N_4439,N_5575);
or U7061 (N_7061,N_5736,N_5190);
or U7062 (N_7062,N_5178,N_4282);
or U7063 (N_7063,N_5942,N_4008);
nand U7064 (N_7064,N_5897,N_4548);
nand U7065 (N_7065,N_4483,N_4553);
or U7066 (N_7066,N_5533,N_5471);
nand U7067 (N_7067,N_4315,N_5262);
nor U7068 (N_7068,N_4303,N_4172);
xnor U7069 (N_7069,N_4217,N_4303);
or U7070 (N_7070,N_5905,N_5736);
nand U7071 (N_7071,N_4747,N_4042);
and U7072 (N_7072,N_4849,N_5880);
or U7073 (N_7073,N_4547,N_4555);
or U7074 (N_7074,N_4975,N_5487);
xnor U7075 (N_7075,N_4800,N_5631);
nand U7076 (N_7076,N_4417,N_4113);
or U7077 (N_7077,N_4229,N_5538);
and U7078 (N_7078,N_5979,N_5987);
xnor U7079 (N_7079,N_5526,N_5999);
xor U7080 (N_7080,N_5971,N_5888);
or U7081 (N_7081,N_5882,N_5162);
nor U7082 (N_7082,N_4515,N_5439);
nand U7083 (N_7083,N_4769,N_4129);
or U7084 (N_7084,N_5480,N_4635);
nor U7085 (N_7085,N_4634,N_5032);
and U7086 (N_7086,N_4807,N_5194);
or U7087 (N_7087,N_4864,N_5383);
and U7088 (N_7088,N_5204,N_5426);
or U7089 (N_7089,N_4702,N_4047);
xor U7090 (N_7090,N_4729,N_4440);
nand U7091 (N_7091,N_5014,N_5533);
or U7092 (N_7092,N_4754,N_4677);
or U7093 (N_7093,N_4653,N_5295);
and U7094 (N_7094,N_5162,N_4998);
and U7095 (N_7095,N_4377,N_4164);
nand U7096 (N_7096,N_4901,N_5455);
and U7097 (N_7097,N_4754,N_4319);
nand U7098 (N_7098,N_5284,N_4287);
nand U7099 (N_7099,N_4046,N_4527);
nor U7100 (N_7100,N_4556,N_4162);
nand U7101 (N_7101,N_4201,N_5823);
nor U7102 (N_7102,N_5215,N_4515);
or U7103 (N_7103,N_5157,N_5917);
or U7104 (N_7104,N_5795,N_5454);
nor U7105 (N_7105,N_4914,N_4081);
or U7106 (N_7106,N_4404,N_5918);
xor U7107 (N_7107,N_4247,N_4746);
and U7108 (N_7108,N_4564,N_4052);
nand U7109 (N_7109,N_4266,N_5670);
nor U7110 (N_7110,N_5717,N_5652);
nor U7111 (N_7111,N_5528,N_4017);
nor U7112 (N_7112,N_5782,N_4493);
xnor U7113 (N_7113,N_4446,N_5647);
and U7114 (N_7114,N_4110,N_4359);
xnor U7115 (N_7115,N_5665,N_4553);
xnor U7116 (N_7116,N_5852,N_4957);
or U7117 (N_7117,N_4012,N_4474);
or U7118 (N_7118,N_5278,N_4210);
nand U7119 (N_7119,N_5560,N_4780);
xor U7120 (N_7120,N_4736,N_5306);
nand U7121 (N_7121,N_4179,N_4409);
or U7122 (N_7122,N_5864,N_5807);
nor U7123 (N_7123,N_5438,N_5647);
xor U7124 (N_7124,N_4178,N_5337);
nand U7125 (N_7125,N_4947,N_5235);
and U7126 (N_7126,N_5543,N_5430);
or U7127 (N_7127,N_4327,N_5450);
nand U7128 (N_7128,N_5775,N_5976);
xnor U7129 (N_7129,N_4575,N_5027);
or U7130 (N_7130,N_5869,N_5563);
nand U7131 (N_7131,N_5153,N_4037);
nor U7132 (N_7132,N_4172,N_5869);
nand U7133 (N_7133,N_5208,N_5868);
nand U7134 (N_7134,N_4628,N_4072);
nand U7135 (N_7135,N_5445,N_5929);
and U7136 (N_7136,N_5792,N_5323);
xor U7137 (N_7137,N_4714,N_4450);
and U7138 (N_7138,N_4682,N_5127);
xor U7139 (N_7139,N_5413,N_5414);
and U7140 (N_7140,N_5089,N_4002);
and U7141 (N_7141,N_4935,N_4520);
and U7142 (N_7142,N_4610,N_4023);
nand U7143 (N_7143,N_5576,N_5684);
and U7144 (N_7144,N_4447,N_4617);
and U7145 (N_7145,N_5516,N_4646);
nor U7146 (N_7146,N_4014,N_5303);
or U7147 (N_7147,N_4972,N_4214);
xnor U7148 (N_7148,N_4947,N_4496);
nor U7149 (N_7149,N_4813,N_5395);
or U7150 (N_7150,N_4714,N_4693);
nor U7151 (N_7151,N_5690,N_5818);
xnor U7152 (N_7152,N_5242,N_4677);
nor U7153 (N_7153,N_4048,N_5958);
or U7154 (N_7154,N_4990,N_5712);
or U7155 (N_7155,N_5669,N_5788);
nor U7156 (N_7156,N_5352,N_5989);
nor U7157 (N_7157,N_5646,N_5917);
and U7158 (N_7158,N_5788,N_4254);
xnor U7159 (N_7159,N_5001,N_4531);
nor U7160 (N_7160,N_4180,N_5783);
xor U7161 (N_7161,N_5015,N_4406);
or U7162 (N_7162,N_4168,N_4530);
nand U7163 (N_7163,N_5767,N_4312);
or U7164 (N_7164,N_4570,N_4827);
and U7165 (N_7165,N_4214,N_5424);
xnor U7166 (N_7166,N_4416,N_5151);
nor U7167 (N_7167,N_5507,N_5840);
xor U7168 (N_7168,N_4036,N_4557);
or U7169 (N_7169,N_5315,N_4860);
xnor U7170 (N_7170,N_5540,N_4131);
or U7171 (N_7171,N_5514,N_5710);
nand U7172 (N_7172,N_4736,N_5416);
xnor U7173 (N_7173,N_5705,N_4103);
xnor U7174 (N_7174,N_4623,N_4108);
nand U7175 (N_7175,N_5360,N_4073);
xor U7176 (N_7176,N_4296,N_4985);
xor U7177 (N_7177,N_4201,N_5841);
and U7178 (N_7178,N_5567,N_4290);
nor U7179 (N_7179,N_4797,N_5488);
or U7180 (N_7180,N_4513,N_5649);
nor U7181 (N_7181,N_5821,N_4446);
nand U7182 (N_7182,N_5472,N_5359);
and U7183 (N_7183,N_5911,N_4553);
nand U7184 (N_7184,N_5052,N_5905);
xor U7185 (N_7185,N_5326,N_5074);
xnor U7186 (N_7186,N_4214,N_5018);
xor U7187 (N_7187,N_4478,N_4279);
and U7188 (N_7188,N_4439,N_4851);
nand U7189 (N_7189,N_4317,N_5348);
or U7190 (N_7190,N_4146,N_5840);
xnor U7191 (N_7191,N_4553,N_4058);
and U7192 (N_7192,N_4379,N_5394);
nand U7193 (N_7193,N_4971,N_4638);
nand U7194 (N_7194,N_5937,N_4509);
nand U7195 (N_7195,N_5578,N_4423);
nand U7196 (N_7196,N_4224,N_5034);
xnor U7197 (N_7197,N_5302,N_4889);
nand U7198 (N_7198,N_4077,N_4528);
or U7199 (N_7199,N_4144,N_4380);
and U7200 (N_7200,N_5471,N_5247);
and U7201 (N_7201,N_4861,N_5530);
nor U7202 (N_7202,N_5175,N_5745);
and U7203 (N_7203,N_5314,N_5855);
xor U7204 (N_7204,N_5467,N_5024);
or U7205 (N_7205,N_4613,N_4055);
xnor U7206 (N_7206,N_4158,N_5612);
nor U7207 (N_7207,N_5882,N_4336);
and U7208 (N_7208,N_4248,N_4056);
or U7209 (N_7209,N_5152,N_4300);
nand U7210 (N_7210,N_5071,N_5369);
nand U7211 (N_7211,N_5561,N_4927);
nand U7212 (N_7212,N_4257,N_5247);
or U7213 (N_7213,N_5352,N_4244);
nor U7214 (N_7214,N_4395,N_5491);
xor U7215 (N_7215,N_5976,N_5351);
nor U7216 (N_7216,N_5790,N_5858);
or U7217 (N_7217,N_5963,N_4775);
xnor U7218 (N_7218,N_4765,N_5003);
nand U7219 (N_7219,N_4328,N_5516);
and U7220 (N_7220,N_5582,N_4851);
nor U7221 (N_7221,N_4411,N_4920);
and U7222 (N_7222,N_5703,N_4875);
and U7223 (N_7223,N_4249,N_5496);
and U7224 (N_7224,N_5233,N_5494);
and U7225 (N_7225,N_5789,N_4828);
nor U7226 (N_7226,N_4080,N_5094);
and U7227 (N_7227,N_4882,N_5392);
nand U7228 (N_7228,N_5620,N_5882);
nor U7229 (N_7229,N_4456,N_4514);
and U7230 (N_7230,N_4641,N_4503);
or U7231 (N_7231,N_5961,N_4447);
or U7232 (N_7232,N_5826,N_5039);
or U7233 (N_7233,N_5058,N_5812);
nand U7234 (N_7234,N_4612,N_5022);
xnor U7235 (N_7235,N_5297,N_5178);
nor U7236 (N_7236,N_4979,N_4724);
nand U7237 (N_7237,N_5843,N_4527);
nand U7238 (N_7238,N_4126,N_4524);
xnor U7239 (N_7239,N_4378,N_4362);
nand U7240 (N_7240,N_4333,N_4206);
xnor U7241 (N_7241,N_4215,N_5262);
nor U7242 (N_7242,N_4850,N_4518);
nor U7243 (N_7243,N_5490,N_5201);
and U7244 (N_7244,N_5327,N_5945);
or U7245 (N_7245,N_4871,N_4154);
nor U7246 (N_7246,N_5367,N_5418);
and U7247 (N_7247,N_4018,N_4125);
nand U7248 (N_7248,N_4756,N_4742);
nor U7249 (N_7249,N_4272,N_5498);
nand U7250 (N_7250,N_4060,N_4992);
nand U7251 (N_7251,N_5833,N_4292);
nor U7252 (N_7252,N_5775,N_5172);
xnor U7253 (N_7253,N_4467,N_4882);
nor U7254 (N_7254,N_4274,N_5633);
and U7255 (N_7255,N_5535,N_4462);
and U7256 (N_7256,N_4225,N_5590);
and U7257 (N_7257,N_4074,N_4192);
xnor U7258 (N_7258,N_4144,N_4775);
nand U7259 (N_7259,N_5622,N_4048);
and U7260 (N_7260,N_5537,N_4616);
or U7261 (N_7261,N_5518,N_4287);
nor U7262 (N_7262,N_4013,N_4195);
xnor U7263 (N_7263,N_4475,N_5424);
nor U7264 (N_7264,N_4277,N_4545);
xor U7265 (N_7265,N_5843,N_4307);
or U7266 (N_7266,N_4282,N_5016);
nor U7267 (N_7267,N_4249,N_5334);
nor U7268 (N_7268,N_5600,N_4931);
xnor U7269 (N_7269,N_5328,N_4390);
nand U7270 (N_7270,N_5510,N_4213);
and U7271 (N_7271,N_4458,N_5637);
nor U7272 (N_7272,N_4044,N_5471);
nor U7273 (N_7273,N_4185,N_5799);
or U7274 (N_7274,N_4841,N_5129);
xor U7275 (N_7275,N_5099,N_5073);
xor U7276 (N_7276,N_4165,N_5429);
xnor U7277 (N_7277,N_4596,N_4841);
or U7278 (N_7278,N_4297,N_5168);
or U7279 (N_7279,N_5628,N_5626);
and U7280 (N_7280,N_4622,N_4260);
or U7281 (N_7281,N_5512,N_5922);
or U7282 (N_7282,N_5695,N_4192);
xor U7283 (N_7283,N_4121,N_5052);
nand U7284 (N_7284,N_5423,N_4631);
nand U7285 (N_7285,N_4889,N_5617);
nand U7286 (N_7286,N_4536,N_5634);
or U7287 (N_7287,N_5127,N_5251);
or U7288 (N_7288,N_4795,N_4455);
and U7289 (N_7289,N_5668,N_4126);
xnor U7290 (N_7290,N_5938,N_5286);
nand U7291 (N_7291,N_4448,N_4465);
nor U7292 (N_7292,N_5698,N_5134);
and U7293 (N_7293,N_4026,N_5310);
nand U7294 (N_7294,N_4360,N_5832);
nor U7295 (N_7295,N_5978,N_4175);
and U7296 (N_7296,N_4823,N_4737);
nand U7297 (N_7297,N_5386,N_5589);
xnor U7298 (N_7298,N_4737,N_5125);
nand U7299 (N_7299,N_5384,N_5017);
nand U7300 (N_7300,N_4979,N_5978);
nor U7301 (N_7301,N_5912,N_4469);
xor U7302 (N_7302,N_4290,N_5495);
or U7303 (N_7303,N_4812,N_4714);
nand U7304 (N_7304,N_5777,N_4539);
xnor U7305 (N_7305,N_5314,N_5290);
and U7306 (N_7306,N_5964,N_5790);
nor U7307 (N_7307,N_4995,N_4180);
xnor U7308 (N_7308,N_5355,N_5994);
xnor U7309 (N_7309,N_5023,N_4833);
xnor U7310 (N_7310,N_4503,N_4695);
nor U7311 (N_7311,N_4215,N_5516);
nor U7312 (N_7312,N_5094,N_5113);
nand U7313 (N_7313,N_4132,N_5713);
or U7314 (N_7314,N_4026,N_5744);
nor U7315 (N_7315,N_4987,N_5344);
xor U7316 (N_7316,N_4961,N_4287);
or U7317 (N_7317,N_5823,N_5973);
nor U7318 (N_7318,N_5575,N_4878);
nand U7319 (N_7319,N_5971,N_5047);
or U7320 (N_7320,N_4154,N_4458);
or U7321 (N_7321,N_4296,N_5804);
or U7322 (N_7322,N_4368,N_5863);
or U7323 (N_7323,N_4001,N_4456);
xnor U7324 (N_7324,N_5731,N_4424);
and U7325 (N_7325,N_4522,N_4655);
nand U7326 (N_7326,N_4897,N_4834);
xnor U7327 (N_7327,N_5657,N_5822);
and U7328 (N_7328,N_5184,N_4706);
xor U7329 (N_7329,N_4239,N_4847);
or U7330 (N_7330,N_4079,N_4604);
and U7331 (N_7331,N_5412,N_5629);
xor U7332 (N_7332,N_5444,N_5490);
nor U7333 (N_7333,N_5859,N_4550);
and U7334 (N_7334,N_4479,N_4596);
or U7335 (N_7335,N_5838,N_4083);
and U7336 (N_7336,N_5659,N_5190);
and U7337 (N_7337,N_5672,N_4346);
nor U7338 (N_7338,N_5691,N_5833);
and U7339 (N_7339,N_4196,N_4703);
nand U7340 (N_7340,N_5218,N_5234);
xor U7341 (N_7341,N_4537,N_4591);
and U7342 (N_7342,N_5784,N_4544);
nand U7343 (N_7343,N_5577,N_4655);
nor U7344 (N_7344,N_4055,N_5048);
and U7345 (N_7345,N_5414,N_4859);
xor U7346 (N_7346,N_5991,N_4137);
nand U7347 (N_7347,N_5865,N_5851);
nand U7348 (N_7348,N_4787,N_5208);
nor U7349 (N_7349,N_4060,N_5452);
xnor U7350 (N_7350,N_5367,N_5223);
and U7351 (N_7351,N_5889,N_5227);
xor U7352 (N_7352,N_4499,N_4548);
and U7353 (N_7353,N_4952,N_4140);
or U7354 (N_7354,N_5896,N_4645);
nor U7355 (N_7355,N_5510,N_4126);
nor U7356 (N_7356,N_4288,N_5668);
nor U7357 (N_7357,N_4041,N_5221);
or U7358 (N_7358,N_4722,N_4884);
nor U7359 (N_7359,N_4452,N_5579);
xor U7360 (N_7360,N_4962,N_5597);
nor U7361 (N_7361,N_5990,N_5470);
xor U7362 (N_7362,N_4045,N_4260);
and U7363 (N_7363,N_5236,N_5961);
xnor U7364 (N_7364,N_4786,N_4966);
and U7365 (N_7365,N_5150,N_5155);
xor U7366 (N_7366,N_4228,N_4882);
nand U7367 (N_7367,N_4962,N_4661);
and U7368 (N_7368,N_5355,N_4276);
nand U7369 (N_7369,N_4080,N_4116);
and U7370 (N_7370,N_5739,N_5049);
xor U7371 (N_7371,N_4119,N_5040);
and U7372 (N_7372,N_4002,N_4338);
nor U7373 (N_7373,N_5494,N_4566);
nor U7374 (N_7374,N_5472,N_5166);
or U7375 (N_7375,N_5834,N_4922);
xnor U7376 (N_7376,N_5581,N_5213);
nand U7377 (N_7377,N_5686,N_5619);
nor U7378 (N_7378,N_4730,N_4253);
nand U7379 (N_7379,N_4498,N_4260);
nand U7380 (N_7380,N_4118,N_5726);
nand U7381 (N_7381,N_4073,N_4735);
nand U7382 (N_7382,N_4911,N_5407);
and U7383 (N_7383,N_4615,N_5961);
xor U7384 (N_7384,N_4421,N_5995);
nand U7385 (N_7385,N_4208,N_5124);
and U7386 (N_7386,N_4386,N_4981);
or U7387 (N_7387,N_5745,N_5474);
or U7388 (N_7388,N_4092,N_5916);
and U7389 (N_7389,N_5722,N_5663);
nand U7390 (N_7390,N_5754,N_5382);
or U7391 (N_7391,N_5302,N_4431);
or U7392 (N_7392,N_4119,N_5852);
or U7393 (N_7393,N_4656,N_5599);
nor U7394 (N_7394,N_4929,N_5168);
nand U7395 (N_7395,N_4080,N_4589);
or U7396 (N_7396,N_5205,N_4533);
xnor U7397 (N_7397,N_5440,N_5024);
xor U7398 (N_7398,N_5357,N_5615);
nor U7399 (N_7399,N_4137,N_4528);
or U7400 (N_7400,N_5585,N_4398);
or U7401 (N_7401,N_4262,N_5055);
and U7402 (N_7402,N_4011,N_5303);
and U7403 (N_7403,N_5064,N_5585);
xor U7404 (N_7404,N_4587,N_4337);
xor U7405 (N_7405,N_4543,N_5986);
and U7406 (N_7406,N_5962,N_5310);
and U7407 (N_7407,N_5732,N_5674);
or U7408 (N_7408,N_5218,N_5538);
xor U7409 (N_7409,N_5376,N_4469);
nor U7410 (N_7410,N_5052,N_5032);
or U7411 (N_7411,N_4390,N_5387);
nand U7412 (N_7412,N_4454,N_5829);
or U7413 (N_7413,N_5978,N_4136);
xnor U7414 (N_7414,N_4751,N_4931);
or U7415 (N_7415,N_4653,N_5780);
xor U7416 (N_7416,N_4613,N_4726);
nor U7417 (N_7417,N_4852,N_5068);
xor U7418 (N_7418,N_4966,N_5903);
xor U7419 (N_7419,N_5067,N_4731);
nor U7420 (N_7420,N_5882,N_5506);
nand U7421 (N_7421,N_5305,N_4883);
xnor U7422 (N_7422,N_5479,N_4026);
xor U7423 (N_7423,N_4830,N_4791);
or U7424 (N_7424,N_5550,N_5416);
and U7425 (N_7425,N_5858,N_4462);
and U7426 (N_7426,N_4176,N_4329);
xor U7427 (N_7427,N_5100,N_5124);
and U7428 (N_7428,N_4678,N_4656);
xnor U7429 (N_7429,N_5347,N_5132);
xor U7430 (N_7430,N_4292,N_4412);
or U7431 (N_7431,N_4826,N_5034);
and U7432 (N_7432,N_4233,N_5935);
or U7433 (N_7433,N_5432,N_5372);
and U7434 (N_7434,N_4067,N_4037);
nand U7435 (N_7435,N_5790,N_5078);
xor U7436 (N_7436,N_5621,N_5378);
or U7437 (N_7437,N_4308,N_4772);
or U7438 (N_7438,N_5730,N_5310);
nand U7439 (N_7439,N_5956,N_5660);
nand U7440 (N_7440,N_4683,N_4094);
xnor U7441 (N_7441,N_5996,N_4169);
xnor U7442 (N_7442,N_5807,N_4052);
nand U7443 (N_7443,N_4943,N_5225);
xor U7444 (N_7444,N_4482,N_4500);
xnor U7445 (N_7445,N_4209,N_5283);
nand U7446 (N_7446,N_5973,N_5613);
nand U7447 (N_7447,N_5051,N_4455);
and U7448 (N_7448,N_5150,N_5283);
and U7449 (N_7449,N_5403,N_5518);
xnor U7450 (N_7450,N_4218,N_5949);
nor U7451 (N_7451,N_5330,N_5147);
xor U7452 (N_7452,N_4156,N_4497);
and U7453 (N_7453,N_4958,N_5076);
nor U7454 (N_7454,N_4306,N_4050);
nand U7455 (N_7455,N_5685,N_4611);
or U7456 (N_7456,N_4941,N_4800);
nor U7457 (N_7457,N_4206,N_4996);
or U7458 (N_7458,N_4019,N_4487);
or U7459 (N_7459,N_5810,N_5178);
and U7460 (N_7460,N_4741,N_5387);
nor U7461 (N_7461,N_4867,N_4298);
nor U7462 (N_7462,N_4064,N_4063);
or U7463 (N_7463,N_5659,N_5569);
nor U7464 (N_7464,N_5204,N_4859);
and U7465 (N_7465,N_5245,N_5677);
xor U7466 (N_7466,N_4737,N_4552);
or U7467 (N_7467,N_4362,N_5046);
and U7468 (N_7468,N_5994,N_4266);
xor U7469 (N_7469,N_4903,N_4478);
xor U7470 (N_7470,N_5568,N_4281);
xor U7471 (N_7471,N_5978,N_5874);
nor U7472 (N_7472,N_4045,N_4315);
and U7473 (N_7473,N_5138,N_4302);
nand U7474 (N_7474,N_4893,N_5114);
nor U7475 (N_7475,N_4845,N_4720);
nand U7476 (N_7476,N_5093,N_4362);
nor U7477 (N_7477,N_5910,N_5033);
nor U7478 (N_7478,N_4927,N_4853);
and U7479 (N_7479,N_5890,N_4605);
nand U7480 (N_7480,N_4172,N_4216);
and U7481 (N_7481,N_5032,N_5854);
nand U7482 (N_7482,N_5159,N_5344);
or U7483 (N_7483,N_4843,N_4860);
or U7484 (N_7484,N_4513,N_4739);
nand U7485 (N_7485,N_5008,N_4450);
nor U7486 (N_7486,N_4726,N_5246);
or U7487 (N_7487,N_4035,N_4750);
xnor U7488 (N_7488,N_5546,N_4224);
or U7489 (N_7489,N_4697,N_4258);
xor U7490 (N_7490,N_5728,N_5675);
or U7491 (N_7491,N_5825,N_5604);
nand U7492 (N_7492,N_5212,N_4016);
xnor U7493 (N_7493,N_4978,N_5121);
and U7494 (N_7494,N_5802,N_5063);
or U7495 (N_7495,N_5539,N_4245);
xor U7496 (N_7496,N_5038,N_5049);
and U7497 (N_7497,N_4804,N_5027);
nand U7498 (N_7498,N_4331,N_5316);
nor U7499 (N_7499,N_5127,N_4344);
or U7500 (N_7500,N_5981,N_5727);
xor U7501 (N_7501,N_5937,N_5944);
xnor U7502 (N_7502,N_5390,N_5033);
nor U7503 (N_7503,N_4443,N_5402);
xor U7504 (N_7504,N_4916,N_5510);
or U7505 (N_7505,N_5164,N_4500);
nand U7506 (N_7506,N_4940,N_4023);
and U7507 (N_7507,N_5694,N_4278);
or U7508 (N_7508,N_5274,N_4174);
and U7509 (N_7509,N_5339,N_5421);
or U7510 (N_7510,N_4899,N_4273);
and U7511 (N_7511,N_4060,N_4191);
xor U7512 (N_7512,N_4968,N_4602);
and U7513 (N_7513,N_5047,N_4487);
nand U7514 (N_7514,N_5805,N_5250);
nor U7515 (N_7515,N_5868,N_5647);
nand U7516 (N_7516,N_5021,N_4966);
xor U7517 (N_7517,N_4344,N_5244);
and U7518 (N_7518,N_5682,N_5420);
nor U7519 (N_7519,N_4658,N_5161);
or U7520 (N_7520,N_4743,N_5935);
xnor U7521 (N_7521,N_5564,N_5799);
nor U7522 (N_7522,N_5201,N_5649);
nor U7523 (N_7523,N_5253,N_5398);
nor U7524 (N_7524,N_5970,N_5310);
nand U7525 (N_7525,N_5505,N_4236);
xor U7526 (N_7526,N_4819,N_5468);
or U7527 (N_7527,N_4970,N_5134);
and U7528 (N_7528,N_5165,N_5275);
nor U7529 (N_7529,N_4299,N_5984);
and U7530 (N_7530,N_4826,N_4012);
nand U7531 (N_7531,N_4542,N_4427);
xor U7532 (N_7532,N_5521,N_4431);
xnor U7533 (N_7533,N_4476,N_5675);
nor U7534 (N_7534,N_5111,N_4225);
nand U7535 (N_7535,N_4937,N_5036);
or U7536 (N_7536,N_5812,N_4991);
nand U7537 (N_7537,N_5167,N_5959);
or U7538 (N_7538,N_4564,N_5473);
or U7539 (N_7539,N_5734,N_4458);
nand U7540 (N_7540,N_4624,N_4769);
or U7541 (N_7541,N_5300,N_5586);
nand U7542 (N_7542,N_5498,N_5239);
nand U7543 (N_7543,N_4139,N_4006);
xor U7544 (N_7544,N_4858,N_4643);
nor U7545 (N_7545,N_4940,N_4802);
xnor U7546 (N_7546,N_5157,N_5230);
or U7547 (N_7547,N_5112,N_4241);
xnor U7548 (N_7548,N_4980,N_4839);
and U7549 (N_7549,N_5828,N_5568);
and U7550 (N_7550,N_5836,N_4786);
nand U7551 (N_7551,N_5713,N_4996);
or U7552 (N_7552,N_5931,N_5737);
xor U7553 (N_7553,N_5522,N_4688);
and U7554 (N_7554,N_4428,N_4030);
and U7555 (N_7555,N_4092,N_5550);
and U7556 (N_7556,N_4436,N_4112);
or U7557 (N_7557,N_4648,N_4105);
nor U7558 (N_7558,N_4968,N_4080);
and U7559 (N_7559,N_5529,N_4709);
nor U7560 (N_7560,N_4058,N_5182);
and U7561 (N_7561,N_4713,N_4148);
and U7562 (N_7562,N_5574,N_5922);
and U7563 (N_7563,N_5364,N_4324);
nor U7564 (N_7564,N_4206,N_4014);
xnor U7565 (N_7565,N_4892,N_5655);
nand U7566 (N_7566,N_4259,N_5726);
nand U7567 (N_7567,N_4035,N_5055);
nand U7568 (N_7568,N_5116,N_4136);
and U7569 (N_7569,N_4555,N_5416);
and U7570 (N_7570,N_4012,N_4975);
xor U7571 (N_7571,N_5908,N_4025);
and U7572 (N_7572,N_5585,N_4213);
and U7573 (N_7573,N_5870,N_5573);
nand U7574 (N_7574,N_5327,N_5512);
nor U7575 (N_7575,N_4751,N_4797);
nor U7576 (N_7576,N_4397,N_4627);
nand U7577 (N_7577,N_4028,N_4542);
nand U7578 (N_7578,N_4475,N_4668);
nor U7579 (N_7579,N_5554,N_4127);
or U7580 (N_7580,N_5349,N_5128);
nor U7581 (N_7581,N_5572,N_4070);
and U7582 (N_7582,N_4499,N_5454);
xnor U7583 (N_7583,N_4549,N_4009);
xnor U7584 (N_7584,N_4852,N_5808);
nand U7585 (N_7585,N_4330,N_5603);
and U7586 (N_7586,N_4017,N_4121);
or U7587 (N_7587,N_4966,N_4475);
and U7588 (N_7588,N_4069,N_5904);
and U7589 (N_7589,N_5884,N_5600);
nand U7590 (N_7590,N_4070,N_5568);
nor U7591 (N_7591,N_4171,N_4037);
xnor U7592 (N_7592,N_4080,N_4935);
or U7593 (N_7593,N_4060,N_4805);
xor U7594 (N_7594,N_4017,N_4097);
nor U7595 (N_7595,N_4899,N_5922);
nand U7596 (N_7596,N_5260,N_5918);
nor U7597 (N_7597,N_4977,N_4526);
nor U7598 (N_7598,N_4400,N_4252);
or U7599 (N_7599,N_5684,N_4408);
xnor U7600 (N_7600,N_5500,N_5715);
nor U7601 (N_7601,N_4026,N_5524);
nand U7602 (N_7602,N_4811,N_4705);
or U7603 (N_7603,N_5069,N_5447);
nor U7604 (N_7604,N_5639,N_5218);
nor U7605 (N_7605,N_5268,N_4467);
nand U7606 (N_7606,N_5414,N_4334);
and U7607 (N_7607,N_5768,N_4757);
nand U7608 (N_7608,N_5832,N_4472);
nand U7609 (N_7609,N_5299,N_4471);
nor U7610 (N_7610,N_4903,N_4267);
and U7611 (N_7611,N_4272,N_4893);
nor U7612 (N_7612,N_5090,N_5022);
nand U7613 (N_7613,N_4099,N_5186);
xnor U7614 (N_7614,N_4876,N_5101);
nor U7615 (N_7615,N_5292,N_5549);
and U7616 (N_7616,N_4872,N_5386);
xnor U7617 (N_7617,N_4811,N_5731);
or U7618 (N_7618,N_5538,N_4791);
nor U7619 (N_7619,N_4009,N_5444);
and U7620 (N_7620,N_4634,N_4673);
xnor U7621 (N_7621,N_5614,N_4912);
and U7622 (N_7622,N_5646,N_4127);
and U7623 (N_7623,N_4275,N_4941);
xnor U7624 (N_7624,N_5305,N_5626);
xnor U7625 (N_7625,N_5197,N_5341);
nor U7626 (N_7626,N_4514,N_4134);
nor U7627 (N_7627,N_5834,N_5886);
nor U7628 (N_7628,N_4581,N_5569);
xor U7629 (N_7629,N_5132,N_5147);
and U7630 (N_7630,N_5737,N_4411);
or U7631 (N_7631,N_5919,N_4016);
and U7632 (N_7632,N_5865,N_5910);
xor U7633 (N_7633,N_4277,N_4583);
xnor U7634 (N_7634,N_4195,N_4942);
nor U7635 (N_7635,N_5938,N_4576);
xor U7636 (N_7636,N_4649,N_4690);
nor U7637 (N_7637,N_5368,N_4243);
nand U7638 (N_7638,N_4105,N_5921);
nor U7639 (N_7639,N_5282,N_5960);
xnor U7640 (N_7640,N_5763,N_5216);
nand U7641 (N_7641,N_5067,N_4197);
and U7642 (N_7642,N_5531,N_4297);
or U7643 (N_7643,N_5138,N_5392);
nand U7644 (N_7644,N_4946,N_4573);
and U7645 (N_7645,N_4421,N_5600);
xnor U7646 (N_7646,N_5855,N_5836);
nor U7647 (N_7647,N_4943,N_5696);
xor U7648 (N_7648,N_5764,N_5623);
and U7649 (N_7649,N_5873,N_5356);
nand U7650 (N_7650,N_5630,N_5729);
or U7651 (N_7651,N_5853,N_4739);
nand U7652 (N_7652,N_4580,N_4620);
nor U7653 (N_7653,N_5877,N_4352);
xnor U7654 (N_7654,N_5247,N_4569);
xnor U7655 (N_7655,N_5057,N_5536);
and U7656 (N_7656,N_4180,N_4790);
nand U7657 (N_7657,N_4287,N_5741);
nor U7658 (N_7658,N_4627,N_5837);
or U7659 (N_7659,N_4454,N_4346);
or U7660 (N_7660,N_5924,N_4542);
nor U7661 (N_7661,N_5483,N_5984);
or U7662 (N_7662,N_5214,N_5656);
and U7663 (N_7663,N_4440,N_4875);
nand U7664 (N_7664,N_4815,N_5466);
nor U7665 (N_7665,N_4109,N_5040);
nand U7666 (N_7666,N_4199,N_4750);
or U7667 (N_7667,N_5224,N_5742);
xor U7668 (N_7668,N_5812,N_4422);
and U7669 (N_7669,N_5659,N_4524);
nand U7670 (N_7670,N_5763,N_5596);
and U7671 (N_7671,N_4120,N_5491);
nor U7672 (N_7672,N_4659,N_4652);
or U7673 (N_7673,N_5845,N_5448);
and U7674 (N_7674,N_4002,N_4390);
or U7675 (N_7675,N_4912,N_5630);
or U7676 (N_7676,N_5231,N_5032);
nor U7677 (N_7677,N_4445,N_4306);
nor U7678 (N_7678,N_5102,N_4708);
nand U7679 (N_7679,N_5160,N_4925);
and U7680 (N_7680,N_5046,N_5983);
xor U7681 (N_7681,N_5722,N_4475);
nand U7682 (N_7682,N_4101,N_4411);
and U7683 (N_7683,N_5285,N_4527);
nor U7684 (N_7684,N_5527,N_5099);
or U7685 (N_7685,N_5949,N_5068);
and U7686 (N_7686,N_5598,N_5486);
or U7687 (N_7687,N_4335,N_5473);
or U7688 (N_7688,N_4315,N_5350);
and U7689 (N_7689,N_5676,N_5271);
nor U7690 (N_7690,N_5006,N_4403);
nor U7691 (N_7691,N_5844,N_5026);
xor U7692 (N_7692,N_4627,N_4943);
nor U7693 (N_7693,N_5911,N_5126);
and U7694 (N_7694,N_4823,N_5538);
and U7695 (N_7695,N_4272,N_5076);
nand U7696 (N_7696,N_5748,N_5688);
xor U7697 (N_7697,N_5922,N_4366);
xor U7698 (N_7698,N_5990,N_4382);
and U7699 (N_7699,N_4054,N_5391);
and U7700 (N_7700,N_5060,N_5166);
and U7701 (N_7701,N_5285,N_5543);
nand U7702 (N_7702,N_5576,N_5629);
nand U7703 (N_7703,N_5005,N_5154);
xnor U7704 (N_7704,N_5761,N_5027);
nand U7705 (N_7705,N_5991,N_4449);
nor U7706 (N_7706,N_4863,N_5702);
or U7707 (N_7707,N_4151,N_4339);
nand U7708 (N_7708,N_5482,N_5770);
or U7709 (N_7709,N_5598,N_4540);
nor U7710 (N_7710,N_4538,N_4322);
nor U7711 (N_7711,N_4700,N_4390);
or U7712 (N_7712,N_4039,N_5613);
nand U7713 (N_7713,N_4190,N_5549);
and U7714 (N_7714,N_5543,N_4228);
xor U7715 (N_7715,N_5839,N_5447);
nand U7716 (N_7716,N_4840,N_4252);
and U7717 (N_7717,N_4616,N_4159);
and U7718 (N_7718,N_4166,N_4255);
and U7719 (N_7719,N_5849,N_5623);
and U7720 (N_7720,N_5289,N_5787);
or U7721 (N_7721,N_4240,N_4423);
nand U7722 (N_7722,N_5096,N_4755);
or U7723 (N_7723,N_4215,N_4771);
xor U7724 (N_7724,N_4723,N_4437);
nor U7725 (N_7725,N_5415,N_4700);
and U7726 (N_7726,N_4122,N_4568);
nor U7727 (N_7727,N_5981,N_5442);
nor U7728 (N_7728,N_5185,N_5035);
and U7729 (N_7729,N_5334,N_5183);
xnor U7730 (N_7730,N_4676,N_5138);
nand U7731 (N_7731,N_5608,N_5481);
nand U7732 (N_7732,N_5557,N_4432);
nor U7733 (N_7733,N_5874,N_5799);
and U7734 (N_7734,N_5190,N_4589);
or U7735 (N_7735,N_5061,N_5460);
and U7736 (N_7736,N_4806,N_5204);
or U7737 (N_7737,N_4480,N_5920);
nand U7738 (N_7738,N_4915,N_5735);
and U7739 (N_7739,N_4924,N_5524);
xnor U7740 (N_7740,N_5561,N_5118);
nor U7741 (N_7741,N_5034,N_4228);
or U7742 (N_7742,N_5535,N_5700);
or U7743 (N_7743,N_4822,N_5174);
and U7744 (N_7744,N_5627,N_5789);
nor U7745 (N_7745,N_5673,N_4486);
and U7746 (N_7746,N_4147,N_4390);
or U7747 (N_7747,N_4609,N_5283);
or U7748 (N_7748,N_4943,N_4264);
xor U7749 (N_7749,N_5185,N_5203);
and U7750 (N_7750,N_5987,N_4670);
nor U7751 (N_7751,N_4197,N_5303);
and U7752 (N_7752,N_4072,N_4980);
and U7753 (N_7753,N_4843,N_4158);
nor U7754 (N_7754,N_5059,N_4618);
or U7755 (N_7755,N_5449,N_4741);
xnor U7756 (N_7756,N_4072,N_5872);
nor U7757 (N_7757,N_4843,N_4255);
and U7758 (N_7758,N_4850,N_5130);
and U7759 (N_7759,N_4304,N_5899);
xor U7760 (N_7760,N_5430,N_4678);
nor U7761 (N_7761,N_5419,N_4010);
nand U7762 (N_7762,N_4464,N_5240);
nor U7763 (N_7763,N_5074,N_5561);
and U7764 (N_7764,N_5641,N_5313);
or U7765 (N_7765,N_5081,N_5692);
nor U7766 (N_7766,N_4996,N_5152);
and U7767 (N_7767,N_4983,N_4576);
or U7768 (N_7768,N_5824,N_5007);
xnor U7769 (N_7769,N_4642,N_4573);
nand U7770 (N_7770,N_4658,N_5313);
xnor U7771 (N_7771,N_4501,N_4134);
and U7772 (N_7772,N_5900,N_5305);
nand U7773 (N_7773,N_5386,N_4498);
or U7774 (N_7774,N_4817,N_4171);
nor U7775 (N_7775,N_4922,N_5220);
xor U7776 (N_7776,N_5882,N_5584);
nor U7777 (N_7777,N_4932,N_4549);
nand U7778 (N_7778,N_4699,N_5749);
and U7779 (N_7779,N_4649,N_5371);
or U7780 (N_7780,N_4498,N_5100);
nand U7781 (N_7781,N_5104,N_5123);
nand U7782 (N_7782,N_5216,N_4988);
and U7783 (N_7783,N_5101,N_4611);
nor U7784 (N_7784,N_5157,N_5286);
or U7785 (N_7785,N_4601,N_5992);
nor U7786 (N_7786,N_4662,N_4160);
nor U7787 (N_7787,N_4088,N_4790);
nor U7788 (N_7788,N_5222,N_4649);
and U7789 (N_7789,N_4526,N_4412);
nor U7790 (N_7790,N_5347,N_5554);
nor U7791 (N_7791,N_4086,N_5006);
and U7792 (N_7792,N_4715,N_5375);
and U7793 (N_7793,N_4516,N_5105);
and U7794 (N_7794,N_4089,N_4747);
xor U7795 (N_7795,N_5160,N_4024);
xnor U7796 (N_7796,N_5092,N_4320);
and U7797 (N_7797,N_5150,N_4645);
nand U7798 (N_7798,N_5535,N_4266);
and U7799 (N_7799,N_4682,N_4492);
nand U7800 (N_7800,N_5879,N_4415);
xor U7801 (N_7801,N_5283,N_5743);
and U7802 (N_7802,N_4076,N_5035);
and U7803 (N_7803,N_4168,N_5121);
and U7804 (N_7804,N_4315,N_5725);
and U7805 (N_7805,N_4387,N_5476);
nand U7806 (N_7806,N_4108,N_4138);
nor U7807 (N_7807,N_4894,N_5318);
xnor U7808 (N_7808,N_4809,N_4400);
and U7809 (N_7809,N_5443,N_5046);
xor U7810 (N_7810,N_4819,N_4547);
and U7811 (N_7811,N_5766,N_4586);
nor U7812 (N_7812,N_4600,N_5743);
nand U7813 (N_7813,N_4742,N_4094);
and U7814 (N_7814,N_5494,N_5509);
or U7815 (N_7815,N_5847,N_4811);
nand U7816 (N_7816,N_5924,N_4868);
and U7817 (N_7817,N_5814,N_4580);
or U7818 (N_7818,N_5386,N_4944);
nand U7819 (N_7819,N_4696,N_5567);
nand U7820 (N_7820,N_5954,N_5310);
nor U7821 (N_7821,N_5635,N_4319);
or U7822 (N_7822,N_5424,N_5230);
nand U7823 (N_7823,N_5658,N_5640);
xnor U7824 (N_7824,N_4372,N_4597);
nor U7825 (N_7825,N_5720,N_5467);
or U7826 (N_7826,N_4683,N_5244);
xnor U7827 (N_7827,N_5502,N_4985);
nor U7828 (N_7828,N_4776,N_4093);
and U7829 (N_7829,N_5229,N_5126);
xnor U7830 (N_7830,N_4289,N_4372);
nor U7831 (N_7831,N_5634,N_5450);
nand U7832 (N_7832,N_5623,N_4542);
nor U7833 (N_7833,N_5830,N_5342);
or U7834 (N_7834,N_4146,N_5596);
or U7835 (N_7835,N_4613,N_5056);
or U7836 (N_7836,N_4098,N_4867);
nand U7837 (N_7837,N_4178,N_4380);
or U7838 (N_7838,N_5716,N_4899);
nor U7839 (N_7839,N_5052,N_4060);
nor U7840 (N_7840,N_5870,N_4771);
nor U7841 (N_7841,N_5632,N_5790);
or U7842 (N_7842,N_5269,N_5703);
xnor U7843 (N_7843,N_5349,N_5674);
xnor U7844 (N_7844,N_4761,N_5614);
or U7845 (N_7845,N_5657,N_5578);
and U7846 (N_7846,N_5377,N_4665);
nor U7847 (N_7847,N_4998,N_5259);
or U7848 (N_7848,N_5872,N_5694);
nand U7849 (N_7849,N_4927,N_4229);
xor U7850 (N_7850,N_5082,N_4404);
or U7851 (N_7851,N_4727,N_5960);
xor U7852 (N_7852,N_5583,N_5805);
or U7853 (N_7853,N_4730,N_5441);
or U7854 (N_7854,N_5826,N_5770);
nor U7855 (N_7855,N_4177,N_5989);
and U7856 (N_7856,N_4110,N_4047);
and U7857 (N_7857,N_4838,N_4871);
xnor U7858 (N_7858,N_5227,N_5275);
and U7859 (N_7859,N_5181,N_5423);
nand U7860 (N_7860,N_4615,N_4489);
and U7861 (N_7861,N_4151,N_4300);
and U7862 (N_7862,N_5702,N_5755);
nand U7863 (N_7863,N_4916,N_4798);
or U7864 (N_7864,N_5145,N_5437);
nor U7865 (N_7865,N_4431,N_4441);
and U7866 (N_7866,N_5595,N_5026);
nand U7867 (N_7867,N_4136,N_5420);
and U7868 (N_7868,N_4540,N_5589);
nor U7869 (N_7869,N_5632,N_5021);
and U7870 (N_7870,N_5961,N_5747);
and U7871 (N_7871,N_4417,N_4768);
nor U7872 (N_7872,N_5058,N_4334);
or U7873 (N_7873,N_4010,N_5965);
xor U7874 (N_7874,N_5531,N_4523);
xor U7875 (N_7875,N_4211,N_4461);
and U7876 (N_7876,N_5737,N_4365);
nor U7877 (N_7877,N_4279,N_4560);
or U7878 (N_7878,N_5908,N_4560);
nand U7879 (N_7879,N_5160,N_5924);
xor U7880 (N_7880,N_4936,N_4715);
or U7881 (N_7881,N_5732,N_5535);
nand U7882 (N_7882,N_5007,N_5040);
or U7883 (N_7883,N_4263,N_4607);
or U7884 (N_7884,N_5008,N_4931);
nor U7885 (N_7885,N_5669,N_4168);
xnor U7886 (N_7886,N_4338,N_5872);
nand U7887 (N_7887,N_5130,N_4873);
nor U7888 (N_7888,N_4610,N_4953);
or U7889 (N_7889,N_5202,N_5469);
nor U7890 (N_7890,N_4449,N_5411);
nor U7891 (N_7891,N_5183,N_4846);
or U7892 (N_7892,N_5825,N_5971);
nand U7893 (N_7893,N_4591,N_4138);
nor U7894 (N_7894,N_4970,N_4881);
nand U7895 (N_7895,N_4591,N_4123);
nand U7896 (N_7896,N_5586,N_5988);
xnor U7897 (N_7897,N_4356,N_4857);
xor U7898 (N_7898,N_5338,N_5306);
xor U7899 (N_7899,N_4517,N_4397);
nor U7900 (N_7900,N_5598,N_4329);
nor U7901 (N_7901,N_5577,N_4678);
nand U7902 (N_7902,N_4723,N_5231);
and U7903 (N_7903,N_5278,N_5408);
xnor U7904 (N_7904,N_4049,N_4074);
or U7905 (N_7905,N_5343,N_5397);
and U7906 (N_7906,N_5434,N_4702);
xor U7907 (N_7907,N_4942,N_4739);
nor U7908 (N_7908,N_4471,N_5851);
or U7909 (N_7909,N_4244,N_5095);
xor U7910 (N_7910,N_4310,N_5178);
and U7911 (N_7911,N_4708,N_4225);
xor U7912 (N_7912,N_4670,N_5411);
or U7913 (N_7913,N_5597,N_5836);
or U7914 (N_7914,N_5391,N_4175);
or U7915 (N_7915,N_4228,N_5797);
xnor U7916 (N_7916,N_4880,N_4610);
nand U7917 (N_7917,N_5866,N_4785);
nor U7918 (N_7918,N_4456,N_5764);
or U7919 (N_7919,N_5401,N_4947);
nor U7920 (N_7920,N_4171,N_4534);
nor U7921 (N_7921,N_4594,N_4905);
nand U7922 (N_7922,N_5915,N_4618);
and U7923 (N_7923,N_5682,N_5612);
nand U7924 (N_7924,N_4904,N_5163);
or U7925 (N_7925,N_5451,N_4629);
or U7926 (N_7926,N_4326,N_5137);
xor U7927 (N_7927,N_4947,N_4656);
and U7928 (N_7928,N_5390,N_5241);
or U7929 (N_7929,N_5145,N_4361);
xnor U7930 (N_7930,N_5121,N_5334);
xor U7931 (N_7931,N_5280,N_5835);
nor U7932 (N_7932,N_4510,N_4052);
and U7933 (N_7933,N_4361,N_4289);
xnor U7934 (N_7934,N_4787,N_4562);
or U7935 (N_7935,N_4863,N_4026);
nand U7936 (N_7936,N_4947,N_4802);
nor U7937 (N_7937,N_4357,N_4374);
and U7938 (N_7938,N_4751,N_5192);
or U7939 (N_7939,N_4664,N_5084);
and U7940 (N_7940,N_4396,N_5217);
nor U7941 (N_7941,N_4408,N_4158);
and U7942 (N_7942,N_4023,N_5344);
nand U7943 (N_7943,N_5449,N_4655);
xor U7944 (N_7944,N_4680,N_4326);
and U7945 (N_7945,N_5374,N_5503);
xnor U7946 (N_7946,N_5540,N_4092);
or U7947 (N_7947,N_5501,N_4530);
xnor U7948 (N_7948,N_4897,N_5308);
or U7949 (N_7949,N_4531,N_4787);
and U7950 (N_7950,N_5608,N_5663);
and U7951 (N_7951,N_4277,N_5719);
or U7952 (N_7952,N_5143,N_5058);
nand U7953 (N_7953,N_5006,N_5826);
xnor U7954 (N_7954,N_5802,N_4789);
xor U7955 (N_7955,N_4603,N_5807);
nand U7956 (N_7956,N_5794,N_5862);
nand U7957 (N_7957,N_5594,N_5436);
or U7958 (N_7958,N_5552,N_4405);
or U7959 (N_7959,N_5813,N_5753);
nor U7960 (N_7960,N_4596,N_4453);
nand U7961 (N_7961,N_5344,N_4294);
xor U7962 (N_7962,N_4559,N_4302);
xor U7963 (N_7963,N_4441,N_5839);
nand U7964 (N_7964,N_5982,N_4962);
xnor U7965 (N_7965,N_4519,N_4923);
nand U7966 (N_7966,N_5844,N_4679);
or U7967 (N_7967,N_4840,N_4767);
xor U7968 (N_7968,N_5205,N_5549);
nand U7969 (N_7969,N_4838,N_4846);
nor U7970 (N_7970,N_4095,N_4002);
or U7971 (N_7971,N_5452,N_5469);
nor U7972 (N_7972,N_5930,N_5006);
xor U7973 (N_7973,N_5062,N_5958);
and U7974 (N_7974,N_4015,N_5709);
nand U7975 (N_7975,N_5445,N_5895);
nor U7976 (N_7976,N_5510,N_5536);
nand U7977 (N_7977,N_4419,N_4655);
nand U7978 (N_7978,N_5897,N_5542);
nand U7979 (N_7979,N_4494,N_4227);
and U7980 (N_7980,N_5149,N_5425);
xor U7981 (N_7981,N_4897,N_4927);
nor U7982 (N_7982,N_4679,N_5166);
nand U7983 (N_7983,N_4255,N_4646);
or U7984 (N_7984,N_5121,N_5532);
nand U7985 (N_7985,N_4438,N_4746);
and U7986 (N_7986,N_5831,N_4496);
and U7987 (N_7987,N_5633,N_5203);
or U7988 (N_7988,N_4479,N_4437);
xor U7989 (N_7989,N_5067,N_5976);
xnor U7990 (N_7990,N_5843,N_5531);
xor U7991 (N_7991,N_5616,N_4184);
xnor U7992 (N_7992,N_5812,N_5255);
nand U7993 (N_7993,N_5084,N_4372);
and U7994 (N_7994,N_4011,N_5862);
nand U7995 (N_7995,N_4007,N_4155);
nand U7996 (N_7996,N_5787,N_5464);
and U7997 (N_7997,N_4695,N_4368);
xor U7998 (N_7998,N_4095,N_4908);
xnor U7999 (N_7999,N_5904,N_4363);
nand U8000 (N_8000,N_7871,N_7091);
nor U8001 (N_8001,N_6848,N_7760);
xor U8002 (N_8002,N_7503,N_7911);
or U8003 (N_8003,N_7113,N_6118);
nand U8004 (N_8004,N_6203,N_7588);
nand U8005 (N_8005,N_7912,N_6673);
xnor U8006 (N_8006,N_7762,N_7852);
xnor U8007 (N_8007,N_6488,N_6693);
and U8008 (N_8008,N_6401,N_7907);
nand U8009 (N_8009,N_7573,N_6264);
nor U8010 (N_8010,N_6459,N_6325);
nand U8011 (N_8011,N_6338,N_7578);
nand U8012 (N_8012,N_7053,N_6267);
nor U8013 (N_8013,N_6553,N_6419);
nand U8014 (N_8014,N_7829,N_7060);
nand U8015 (N_8015,N_7270,N_6501);
nor U8016 (N_8016,N_7181,N_7672);
nor U8017 (N_8017,N_7118,N_6932);
xnor U8018 (N_8018,N_6098,N_6744);
xor U8019 (N_8019,N_6705,N_6953);
and U8020 (N_8020,N_6321,N_7146);
or U8021 (N_8021,N_7376,N_6492);
and U8022 (N_8022,N_6233,N_6346);
xor U8023 (N_8023,N_6213,N_7169);
or U8024 (N_8024,N_7265,N_6897);
or U8025 (N_8025,N_6371,N_7096);
and U8026 (N_8026,N_7788,N_7010);
or U8027 (N_8027,N_7650,N_6397);
nor U8028 (N_8028,N_6797,N_7136);
and U8029 (N_8029,N_6446,N_6412);
xor U8030 (N_8030,N_7453,N_7652);
nor U8031 (N_8031,N_6631,N_7632);
and U8032 (N_8032,N_7132,N_6664);
nand U8033 (N_8033,N_6902,N_7383);
nor U8034 (N_8034,N_7687,N_7421);
xnor U8035 (N_8035,N_7474,N_6119);
or U8036 (N_8036,N_6234,N_7472);
nand U8037 (N_8037,N_7969,N_7732);
xnor U8038 (N_8038,N_7348,N_7694);
or U8039 (N_8039,N_6124,N_6508);
or U8040 (N_8040,N_7833,N_7357);
or U8041 (N_8041,N_7867,N_7950);
nor U8042 (N_8042,N_6512,N_6976);
or U8043 (N_8043,N_7860,N_7440);
xor U8044 (N_8044,N_7700,N_7241);
xor U8045 (N_8045,N_7373,N_6737);
or U8046 (N_8046,N_7576,N_7488);
xor U8047 (N_8047,N_6350,N_7078);
or U8048 (N_8048,N_7550,N_7959);
nand U8049 (N_8049,N_6465,N_7818);
nand U8050 (N_8050,N_6936,N_7894);
xnor U8051 (N_8051,N_6210,N_7556);
and U8052 (N_8052,N_6909,N_7901);
or U8053 (N_8053,N_7929,N_7423);
nor U8054 (N_8054,N_7039,N_6357);
or U8055 (N_8055,N_6109,N_6067);
or U8056 (N_8056,N_6417,N_7174);
xnor U8057 (N_8057,N_6448,N_7415);
nand U8058 (N_8058,N_6453,N_6431);
and U8059 (N_8059,N_7675,N_7221);
and U8060 (N_8060,N_6180,N_7756);
or U8061 (N_8061,N_7710,N_6777);
or U8062 (N_8062,N_7344,N_6018);
nand U8063 (N_8063,N_7935,N_6577);
nand U8064 (N_8064,N_6759,N_7076);
xor U8065 (N_8065,N_6855,N_7191);
or U8066 (N_8066,N_6318,N_6939);
nand U8067 (N_8067,N_6490,N_6340);
nand U8068 (N_8068,N_7057,N_6351);
or U8069 (N_8069,N_7522,N_7718);
or U8070 (N_8070,N_6965,N_7046);
or U8071 (N_8071,N_6838,N_6913);
nor U8072 (N_8072,N_7093,N_7305);
xnor U8073 (N_8073,N_6937,N_7562);
or U8074 (N_8074,N_6060,N_7134);
nand U8075 (N_8075,N_6454,N_7275);
and U8076 (N_8076,N_6919,N_7387);
nor U8077 (N_8077,N_7831,N_7048);
nand U8078 (N_8078,N_6395,N_6516);
nor U8079 (N_8079,N_7875,N_6150);
xnor U8080 (N_8080,N_7439,N_6510);
nor U8081 (N_8081,N_7869,N_7375);
or U8082 (N_8082,N_6772,N_7792);
nand U8083 (N_8083,N_7333,N_6557);
xor U8084 (N_8084,N_6404,N_7315);
and U8085 (N_8085,N_6598,N_7186);
nand U8086 (N_8086,N_6178,N_6741);
or U8087 (N_8087,N_7248,N_7783);
xnor U8088 (N_8088,N_6611,N_6266);
nor U8089 (N_8089,N_7560,N_6201);
and U8090 (N_8090,N_6407,N_7279);
and U8091 (N_8091,N_6829,N_6522);
or U8092 (N_8092,N_6602,N_6284);
xor U8093 (N_8093,N_7495,N_6593);
nand U8094 (N_8094,N_7544,N_6260);
nor U8095 (N_8095,N_7530,N_7583);
nand U8096 (N_8096,N_7317,N_7176);
xor U8097 (N_8097,N_6154,N_7160);
nor U8098 (N_8098,N_6388,N_7189);
and U8099 (N_8099,N_6658,N_6071);
or U8100 (N_8100,N_7660,N_7702);
nor U8101 (N_8101,N_7204,N_6344);
nor U8102 (N_8102,N_6339,N_6507);
nand U8103 (N_8103,N_7779,N_7830);
nand U8104 (N_8104,N_7516,N_7570);
nor U8105 (N_8105,N_6545,N_6819);
and U8106 (N_8106,N_7484,N_7065);
nor U8107 (N_8107,N_6229,N_6808);
and U8108 (N_8108,N_6943,N_7165);
and U8109 (N_8109,N_6596,N_7519);
nand U8110 (N_8110,N_6002,N_6420);
xor U8111 (N_8111,N_6620,N_6164);
nand U8112 (N_8112,N_6176,N_6136);
nor U8113 (N_8113,N_7904,N_6704);
xor U8114 (N_8114,N_6333,N_7567);
nor U8115 (N_8115,N_6426,N_6918);
xnor U8116 (N_8116,N_6722,N_7565);
and U8117 (N_8117,N_6949,N_6991);
and U8118 (N_8118,N_6539,N_7074);
or U8119 (N_8119,N_6096,N_7748);
nand U8120 (N_8120,N_7608,N_6125);
or U8121 (N_8121,N_7625,N_6640);
xor U8122 (N_8122,N_7478,N_6627);
xnor U8123 (N_8123,N_7858,N_7752);
xor U8124 (N_8124,N_6005,N_6615);
and U8125 (N_8125,N_6372,N_6961);
nor U8126 (N_8126,N_7533,N_7553);
and U8127 (N_8127,N_7686,N_6526);
or U8128 (N_8128,N_7329,N_6051);
xnor U8129 (N_8129,N_6236,N_6258);
xor U8130 (N_8130,N_6482,N_7507);
or U8131 (N_8131,N_7714,N_7701);
nand U8132 (N_8132,N_6847,N_7262);
nor U8133 (N_8133,N_7501,N_7443);
nand U8134 (N_8134,N_7704,N_6728);
nand U8135 (N_8135,N_6100,N_7386);
and U8136 (N_8136,N_7001,N_6194);
or U8137 (N_8137,N_6521,N_6581);
and U8138 (N_8138,N_7663,N_7446);
xor U8139 (N_8139,N_7953,N_6600);
and U8140 (N_8140,N_6089,N_7427);
nand U8141 (N_8141,N_7525,N_6850);
nand U8142 (N_8142,N_6588,N_6992);
nor U8143 (N_8143,N_6138,N_6319);
nor U8144 (N_8144,N_7476,N_7177);
nor U8145 (N_8145,N_6240,N_6671);
and U8146 (N_8146,N_7041,N_7033);
xnor U8147 (N_8147,N_6108,N_6066);
and U8148 (N_8148,N_6774,N_7677);
and U8149 (N_8149,N_6572,N_7623);
and U8150 (N_8150,N_6152,N_7441);
or U8151 (N_8151,N_6757,N_7541);
nor U8152 (N_8152,N_6126,N_7081);
nor U8153 (N_8153,N_7887,N_6544);
and U8154 (N_8154,N_7925,N_7910);
nor U8155 (N_8155,N_7771,N_6785);
nand U8156 (N_8156,N_6037,N_6479);
xnor U8157 (N_8157,N_7325,N_7171);
nand U8158 (N_8158,N_6987,N_6969);
xnor U8159 (N_8159,N_6549,N_7346);
or U8160 (N_8160,N_7938,N_7644);
nor U8161 (N_8161,N_6297,N_6908);
or U8162 (N_8162,N_6279,N_6123);
xor U8163 (N_8163,N_6439,N_6625);
nor U8164 (N_8164,N_6997,N_6696);
and U8165 (N_8165,N_7497,N_6043);
xor U8166 (N_8166,N_6677,N_7998);
and U8167 (N_8167,N_6276,N_6065);
nand U8168 (N_8168,N_6767,N_7297);
or U8169 (N_8169,N_6374,N_7500);
nor U8170 (N_8170,N_7207,N_7648);
nor U8171 (N_8171,N_7738,N_6172);
nand U8172 (N_8172,N_6585,N_6167);
nor U8173 (N_8173,N_6509,N_7984);
and U8174 (N_8174,N_6416,N_7278);
nor U8175 (N_8175,N_6537,N_6707);
nor U8176 (N_8176,N_7037,N_6894);
nand U8177 (N_8177,N_7784,N_6608);
nor U8178 (N_8178,N_6562,N_6183);
and U8179 (N_8179,N_6460,N_6144);
and U8180 (N_8180,N_7157,N_7908);
nand U8181 (N_8181,N_7754,N_7006);
nor U8182 (N_8182,N_7142,N_7896);
xnor U8183 (N_8183,N_6329,N_6674);
and U8184 (N_8184,N_6534,N_7244);
nor U8185 (N_8185,N_6189,N_6868);
xnor U8186 (N_8186,N_7296,N_7647);
nor U8187 (N_8187,N_7347,N_6307);
and U8188 (N_8188,N_6193,N_7891);
nor U8189 (N_8189,N_6896,N_6323);
and U8190 (N_8190,N_6034,N_7158);
or U8191 (N_8191,N_6146,N_7085);
nand U8192 (N_8192,N_7480,N_7836);
or U8193 (N_8193,N_7504,N_7673);
xnor U8194 (N_8194,N_6940,N_7363);
nand U8195 (N_8195,N_6216,N_6026);
and U8196 (N_8196,N_6445,N_7035);
or U8197 (N_8197,N_6480,N_6175);
nand U8198 (N_8198,N_7367,N_7155);
nor U8199 (N_8199,N_7414,N_7314);
nor U8200 (N_8200,N_7083,N_6352);
or U8201 (N_8201,N_7222,N_6017);
nor U8202 (N_8202,N_6773,N_7088);
and U8203 (N_8203,N_7259,N_7341);
xnor U8204 (N_8204,N_6105,N_7599);
or U8205 (N_8205,N_6709,N_7536);
and U8206 (N_8206,N_7388,N_6822);
nand U8207 (N_8207,N_6659,N_7437);
xor U8208 (N_8208,N_6881,N_6244);
xor U8209 (N_8209,N_6998,N_6610);
nor U8210 (N_8210,N_6502,N_6008);
or U8211 (N_8211,N_6062,N_6679);
nand U8212 (N_8212,N_7005,N_7403);
xnor U8213 (N_8213,N_7012,N_7619);
and U8214 (N_8214,N_7238,N_6301);
nor U8215 (N_8215,N_7506,N_7260);
nand U8216 (N_8216,N_6783,N_7895);
and U8217 (N_8217,N_7641,N_7202);
nor U8218 (N_8218,N_6921,N_7267);
or U8219 (N_8219,N_6725,N_6758);
or U8220 (N_8220,N_7196,N_6665);
nor U8221 (N_8221,N_7313,N_7825);
nor U8222 (N_8222,N_7511,N_7458);
xor U8223 (N_8223,N_6622,N_7678);
or U8224 (N_8224,N_7526,N_7144);
or U8225 (N_8225,N_6252,N_7050);
nand U8226 (N_8226,N_6145,N_6143);
or U8227 (N_8227,N_7351,N_6160);
nand U8228 (N_8228,N_7261,N_6487);
nor U8229 (N_8229,N_6700,N_7900);
xor U8230 (N_8230,N_6901,N_6683);
and U8231 (N_8231,N_7154,N_6038);
xnor U8232 (N_8232,N_7288,N_7483);
nand U8233 (N_8233,N_7429,N_6649);
xnor U8234 (N_8234,N_6692,N_7508);
xor U8235 (N_8235,N_7482,N_7442);
or U8236 (N_8236,N_7849,N_7264);
and U8237 (N_8237,N_7949,N_6583);
nor U8238 (N_8238,N_6449,N_7470);
and U8239 (N_8239,N_7521,N_7127);
nor U8240 (N_8240,N_6923,N_7569);
nor U8241 (N_8241,N_7843,N_6643);
xnor U8242 (N_8242,N_6481,N_7123);
xor U8243 (N_8243,N_7587,N_7454);
nor U8244 (N_8244,N_6751,N_6054);
nand U8245 (N_8245,N_6157,N_7767);
xnor U8246 (N_8246,N_6720,N_7234);
nand U8247 (N_8247,N_7232,N_7308);
nor U8248 (N_8248,N_6982,N_6462);
and U8249 (N_8249,N_7834,N_7943);
and U8250 (N_8250,N_7990,N_6666);
nor U8251 (N_8251,N_6314,N_7739);
nand U8252 (N_8252,N_6361,N_7581);
nor U8253 (N_8253,N_7527,N_6364);
nand U8254 (N_8254,N_6869,N_7820);
or U8255 (N_8255,N_6354,N_6827);
nand U8256 (N_8256,N_6116,N_7603);
nor U8257 (N_8257,N_7302,N_7185);
and U8258 (N_8258,N_6450,N_7575);
or U8259 (N_8259,N_7110,N_6898);
nand U8260 (N_8260,N_7662,N_7780);
xor U8261 (N_8261,N_7361,N_7517);
or U8262 (N_8262,N_6163,N_7156);
and U8263 (N_8263,N_6133,N_7218);
or U8264 (N_8264,N_6478,N_7636);
nand U8265 (N_8265,N_7448,N_7757);
and U8266 (N_8266,N_7397,N_6265);
nand U8267 (N_8267,N_7957,N_6697);
and U8268 (N_8268,N_6675,N_7306);
and U8269 (N_8269,N_6515,N_7332);
and U8270 (N_8270,N_7826,N_7774);
nand U8271 (N_8271,N_6379,N_6073);
nand U8272 (N_8272,N_7179,N_7293);
or U8273 (N_8273,N_6560,N_6957);
and U8274 (N_8274,N_7477,N_6775);
and U8275 (N_8275,N_6246,N_7324);
nor U8276 (N_8276,N_7170,N_6910);
and U8277 (N_8277,N_7642,N_7939);
xor U8278 (N_8278,N_7840,N_6699);
xnor U8279 (N_8279,N_7140,N_7976);
xnor U8280 (N_8280,N_6289,N_7954);
nand U8281 (N_8281,N_6520,N_7645);
nand U8282 (N_8282,N_7385,N_7251);
nor U8283 (N_8283,N_7696,N_6428);
and U8284 (N_8284,N_6800,N_6187);
or U8285 (N_8285,N_6025,N_7372);
nand U8286 (N_8286,N_6399,N_6142);
or U8287 (N_8287,N_7596,N_7974);
nor U8288 (N_8288,N_6712,N_7220);
nand U8289 (N_8289,N_6447,N_6542);
or U8290 (N_8290,N_6928,N_6540);
or U8291 (N_8291,N_6027,N_6418);
nor U8292 (N_8292,N_7068,N_6941);
nor U8293 (N_8293,N_6781,N_7670);
nand U8294 (N_8294,N_6646,N_6378);
nor U8295 (N_8295,N_7119,N_6635);
and U8296 (N_8296,N_6834,N_6215);
or U8297 (N_8297,N_6736,N_7310);
xnor U8298 (N_8298,N_7810,N_7630);
nand U8299 (N_8299,N_7613,N_7208);
or U8300 (N_8300,N_6155,N_7892);
xnor U8301 (N_8301,N_6900,N_6042);
nor U8302 (N_8302,N_6255,N_6220);
nand U8303 (N_8303,N_6195,N_7666);
xnor U8304 (N_8304,N_6802,N_7552);
xnor U8305 (N_8305,N_6655,N_6792);
xnor U8306 (N_8306,N_7451,N_6647);
xor U8307 (N_8307,N_7917,N_6995);
nor U8308 (N_8308,N_7152,N_6729);
nand U8309 (N_8309,N_6129,N_7029);
nor U8310 (N_8310,N_7649,N_6398);
nand U8311 (N_8311,N_7226,N_7610);
xnor U8312 (N_8312,N_6552,N_7182);
xnor U8313 (N_8313,N_7921,N_7209);
xnor U8314 (N_8314,N_6093,N_6040);
nand U8315 (N_8315,N_6111,N_7913);
nor U8316 (N_8316,N_6874,N_7611);
or U8317 (N_8317,N_6927,N_6636);
nand U8318 (N_8318,N_6415,N_7903);
nand U8319 (N_8319,N_7124,N_6656);
xnor U8320 (N_8320,N_6019,N_6857);
nand U8321 (N_8321,N_7729,N_6331);
xor U8322 (N_8322,N_7231,N_6559);
nand U8323 (N_8323,N_7628,N_7043);
and U8324 (N_8324,N_7680,N_6861);
or U8325 (N_8325,N_7551,N_7724);
and U8326 (N_8326,N_7456,N_7750);
xor U8327 (N_8327,N_6293,N_6298);
xor U8328 (N_8328,N_7566,N_6947);
xnor U8329 (N_8329,N_6077,N_6715);
nor U8330 (N_8330,N_6474,N_6531);
nand U8331 (N_8331,N_7047,N_7120);
nand U8332 (N_8332,N_6742,N_6001);
and U8333 (N_8333,N_7635,N_7633);
and U8334 (N_8334,N_7405,N_6814);
and U8335 (N_8335,N_6082,N_6734);
xnor U8336 (N_8336,N_6633,N_6669);
nand U8337 (N_8337,N_7066,N_6746);
xnor U8338 (N_8338,N_6930,N_7392);
and U8339 (N_8339,N_7095,N_6366);
and U8340 (N_8340,N_6546,N_6999);
nor U8341 (N_8341,N_6645,N_6393);
nand U8342 (N_8342,N_6566,N_6769);
and U8343 (N_8343,N_7758,N_7621);
and U8344 (N_8344,N_6326,N_7245);
xnor U8345 (N_8345,N_7092,N_7749);
and U8346 (N_8346,N_6074,N_6489);
nor U8347 (N_8347,N_6435,N_6239);
xor U8348 (N_8348,N_6343,N_6022);
xor U8349 (N_8349,N_6607,N_6871);
nand U8350 (N_8350,N_6069,N_7977);
nand U8351 (N_8351,N_7365,N_6994);
nor U8352 (N_8352,N_7547,N_6370);
and U8353 (N_8353,N_6626,N_6771);
nor U8354 (N_8354,N_7319,N_6532);
nand U8355 (N_8355,N_7434,N_6905);
or U8356 (N_8356,N_6832,N_6963);
nor U8357 (N_8357,N_6873,N_7580);
xor U8358 (N_8358,N_6859,N_7706);
and U8359 (N_8359,N_7883,N_6461);
or U8360 (N_8360,N_6437,N_6570);
nor U8361 (N_8361,N_6533,N_6687);
or U8362 (N_8362,N_6477,N_7125);
nand U8363 (N_8363,N_6342,N_6837);
nor U8364 (N_8364,N_6525,N_6754);
and U8365 (N_8365,N_6843,N_6595);
nand U8366 (N_8366,N_7751,N_7183);
xnor U8367 (N_8367,N_7004,N_6591);
and U8368 (N_8368,N_7283,N_6499);
xnor U8369 (N_8369,N_6968,N_6456);
xor U8370 (N_8370,N_6799,N_6468);
xnor U8371 (N_8371,N_7730,N_7989);
nand U8372 (N_8372,N_6724,N_6347);
nor U8373 (N_8373,N_7487,N_7590);
nor U8374 (N_8374,N_6204,N_6341);
and U8375 (N_8375,N_7072,N_7745);
nand U8376 (N_8376,N_6305,N_7795);
and U8377 (N_8377,N_7377,N_7847);
and U8378 (N_8378,N_6335,N_7129);
nand U8379 (N_8379,N_6429,N_6558);
or U8380 (N_8380,N_6384,N_6270);
nand U8381 (N_8381,N_7369,N_7736);
xor U8382 (N_8382,N_6668,N_6353);
and U8383 (N_8383,N_7726,N_6786);
or U8384 (N_8384,N_7548,N_7071);
and U8385 (N_8385,N_6422,N_7090);
nand U8386 (N_8386,N_6875,N_7335);
nand U8387 (N_8387,N_6807,N_7664);
xor U8388 (N_8388,N_6044,N_6836);
nor U8389 (N_8389,N_6660,N_6613);
or U8390 (N_8390,N_6275,N_7698);
or U8391 (N_8391,N_7802,N_7358);
nor U8392 (N_8392,N_6891,N_6726);
or U8393 (N_8393,N_7824,N_7098);
nand U8394 (N_8394,N_6153,N_7153);
or U8395 (N_8395,N_7854,N_7584);
xnor U8396 (N_8396,N_7469,N_7431);
nand U8397 (N_8397,N_6761,N_6962);
or U8398 (N_8398,N_6609,N_6020);
nand U8399 (N_8399,N_6784,N_7592);
or U8400 (N_8400,N_6983,N_7284);
nor U8401 (N_8401,N_6253,N_6322);
nor U8402 (N_8402,N_6592,N_6003);
nand U8403 (N_8403,N_6045,N_6653);
and U8404 (N_8404,N_7378,N_6817);
nor U8405 (N_8405,N_6245,N_6348);
xnor U8406 (N_8406,N_7709,N_7486);
nand U8407 (N_8407,N_6464,N_7671);
nand U8408 (N_8408,N_6458,N_7491);
and U8409 (N_8409,N_6496,N_6409);
and U8410 (N_8410,N_6095,N_7393);
xnor U8411 (N_8411,N_6466,N_7117);
and U8412 (N_8412,N_7946,N_6550);
nor U8413 (N_8413,N_6390,N_7199);
xor U8414 (N_8414,N_6711,N_7395);
xnor U8415 (N_8415,N_7693,N_6355);
and U8416 (N_8416,N_7545,N_7013);
nand U8417 (N_8417,N_6053,N_6391);
or U8418 (N_8418,N_7857,N_7087);
nand U8419 (N_8419,N_7586,N_7778);
nand U8420 (N_8420,N_7539,N_6920);
or U8421 (N_8421,N_6484,N_6251);
nor U8422 (N_8422,N_6052,N_6336);
nand U8423 (N_8423,N_7669,N_7410);
and U8424 (N_8424,N_7281,N_7513);
nor U8425 (N_8425,N_7941,N_6914);
and U8426 (N_8426,N_6756,N_7011);
nand U8427 (N_8427,N_7349,N_7064);
nand U8428 (N_8428,N_6916,N_6945);
or U8429 (N_8429,N_7389,N_7534);
xnor U8430 (N_8430,N_7430,N_6302);
nor U8431 (N_8431,N_6506,N_6046);
and U8432 (N_8432,N_6954,N_7808);
xor U8433 (N_8433,N_6638,N_7744);
or U8434 (N_8434,N_6548,N_7032);
nor U8435 (N_8435,N_6662,N_7356);
and U8436 (N_8436,N_6956,N_6684);
nor U8437 (N_8437,N_7067,N_6056);
xnor U8438 (N_8438,N_7416,N_7239);
xnor U8439 (N_8439,N_6132,N_6667);
xnor U8440 (N_8440,N_7390,N_6396);
and U8441 (N_8441,N_6670,N_6594);
and U8442 (N_8442,N_6958,N_6796);
nand U8443 (N_8443,N_6605,N_7121);
and U8444 (N_8444,N_6892,N_6358);
nand U8445 (N_8445,N_7657,N_6887);
or U8446 (N_8446,N_7639,N_7017);
or U8447 (N_8447,N_6114,N_7789);
xnor U8448 (N_8448,N_7916,N_7838);
nand U8449 (N_8449,N_6029,N_6717);
xor U8450 (N_8450,N_7790,N_6360);
nor U8451 (N_8451,N_7229,N_7277);
nand U8452 (N_8452,N_6639,N_6714);
xnor U8453 (N_8453,N_6543,N_6809);
nand U8454 (N_8454,N_6934,N_7112);
nor U8455 (N_8455,N_6547,N_6990);
nand U8456 (N_8456,N_6495,N_7817);
and U8457 (N_8457,N_6895,N_6064);
nand U8458 (N_8458,N_6863,N_6893);
nand U8459 (N_8459,N_6768,N_7148);
and U8460 (N_8460,N_6122,N_6048);
nor U8461 (N_8461,N_7918,N_6529);
nor U8462 (N_8462,N_7964,N_7885);
xor U8463 (N_8463,N_7192,N_7743);
nand U8464 (N_8464,N_6006,N_7816);
nand U8465 (N_8465,N_6970,N_6681);
xor U8466 (N_8466,N_6092,N_6831);
nand U8467 (N_8467,N_7518,N_6899);
nor U8468 (N_8468,N_7409,N_6231);
and U8469 (N_8469,N_7252,N_7955);
xor U8470 (N_8470,N_6966,N_6036);
xnor U8471 (N_8471,N_7591,N_7131);
nand U8472 (N_8472,N_6373,N_7995);
nor U8473 (N_8473,N_7832,N_6228);
nor U8474 (N_8474,N_7031,N_6030);
xor U8475 (N_8475,N_7028,N_7973);
xnor U8476 (N_8476,N_7674,N_6890);
and U8477 (N_8477,N_6188,N_6385);
nor U8478 (N_8478,N_6903,N_7256);
nor U8479 (N_8479,N_7294,N_6806);
xnor U8480 (N_8480,N_6821,N_6889);
xnor U8481 (N_8481,N_7606,N_6514);
or U8482 (N_8482,N_6198,N_7602);
or U8483 (N_8483,N_7133,N_6191);
and U8484 (N_8484,N_6214,N_6691);
xor U8485 (N_8485,N_7948,N_7617);
nor U8486 (N_8486,N_7203,N_7886);
nor U8487 (N_8487,N_7051,N_6565);
nor U8488 (N_8488,N_7352,N_7637);
xnor U8489 (N_8489,N_6106,N_7609);
or U8490 (N_8490,N_7007,N_7167);
nand U8491 (N_8491,N_7055,N_7366);
and U8492 (N_8492,N_6623,N_6951);
nor U8493 (N_8493,N_6402,N_6579);
nand U8494 (N_8494,N_6225,N_7727);
and U8495 (N_8495,N_7612,N_7558);
or U8496 (N_8496,N_6985,N_6942);
nand U8497 (N_8497,N_7682,N_7339);
nand U8498 (N_8498,N_7747,N_6567);
nor U8499 (N_8499,N_7016,N_6277);
or U8500 (N_8500,N_7321,N_6530);
nor U8501 (N_8501,N_6763,N_6624);
or U8502 (N_8502,N_7166,N_7360);
and U8503 (N_8503,N_6441,N_7881);
nand U8504 (N_8504,N_7723,N_6292);
xor U8505 (N_8505,N_7298,N_7931);
xor U8506 (N_8506,N_7985,N_7003);
nor U8507 (N_8507,N_7399,N_7899);
nand U8508 (N_8508,N_7851,N_7338);
and U8509 (N_8509,N_6291,N_7018);
xnor U8510 (N_8510,N_7691,N_7952);
nand U8511 (N_8511,N_6158,N_6476);
nand U8512 (N_8512,N_7850,N_7184);
and U8513 (N_8513,N_7906,N_6280);
or U8514 (N_8514,N_7620,N_7111);
xnor U8515 (N_8515,N_6877,N_6904);
or U8516 (N_8516,N_7105,N_7024);
xnor U8517 (N_8517,N_6375,N_6926);
nor U8518 (N_8518,N_6269,N_7301);
xnor U8519 (N_8519,N_6285,N_6128);
nor U8520 (N_8520,N_6173,N_7097);
and U8521 (N_8521,N_6882,N_7785);
nor U8522 (N_8522,N_7863,N_6755);
and U8523 (N_8523,N_7496,N_7336);
nand U8524 (N_8524,N_6286,N_6685);
nor U8525 (N_8525,N_7890,N_7063);
or U8526 (N_8526,N_6103,N_7042);
or U8527 (N_8527,N_6770,N_6306);
nand U8528 (N_8528,N_6504,N_6241);
or U8529 (N_8529,N_6411,N_6021);
xor U8530 (N_8530,N_6917,N_7845);
and U8531 (N_8531,N_6367,N_6294);
nor U8532 (N_8532,N_6973,N_7116);
nand U8533 (N_8533,N_6369,N_7417);
xor U8534 (N_8534,N_6224,N_7934);
nor U8535 (N_8535,N_6091,N_6642);
or U8536 (N_8536,N_7109,N_6181);
or U8537 (N_8537,N_7848,N_6612);
nand U8538 (N_8538,N_6629,N_7972);
xor U8539 (N_8539,N_6839,N_7510);
nor U8540 (N_8540,N_7607,N_7194);
nand U8541 (N_8541,N_7654,N_7303);
nor U8542 (N_8542,N_7280,N_6400);
nand U8543 (N_8543,N_6719,N_6498);
and U8544 (N_8544,N_6423,N_7282);
and U8545 (N_8545,N_7107,N_7772);
xor U8546 (N_8546,N_7180,N_7515);
and U8547 (N_8547,N_7930,N_6818);
xnor U8548 (N_8548,N_6686,N_7103);
and U8549 (N_8549,N_6107,N_7956);
and U8550 (N_8550,N_7658,N_6924);
and U8551 (N_8551,N_7475,N_6368);
nor U8552 (N_8552,N_6184,N_6059);
nand U8553 (N_8553,N_6117,N_6584);
and U8554 (N_8554,N_6324,N_7273);
nand U8555 (N_8555,N_7000,N_7712);
and U8556 (N_8556,N_7312,N_6867);
xnor U8557 (N_8557,N_7342,N_6804);
or U8558 (N_8558,N_7986,N_6483);
nand U8559 (N_8559,N_6813,N_7128);
nor U8560 (N_8560,N_6413,N_6823);
or U8561 (N_8561,N_6242,N_6151);
xnor U8562 (N_8562,N_6967,N_6055);
nand U8563 (N_8563,N_7624,N_7407);
xnor U8564 (N_8564,N_6356,N_6197);
xor U8565 (N_8565,N_7467,N_7631);
xor U8566 (N_8566,N_7286,N_6312);
or U8567 (N_8567,N_7782,N_7733);
or U8568 (N_8568,N_6386,N_7626);
or U8569 (N_8569,N_7554,N_7145);
and U8570 (N_8570,N_6110,N_6888);
and U8571 (N_8571,N_6938,N_6207);
xor U8572 (N_8572,N_7008,N_7036);
or U8573 (N_8573,N_7276,N_6041);
xor U8574 (N_8574,N_7371,N_6009);
and U8575 (N_8575,N_7629,N_7077);
and U8576 (N_8576,N_7528,N_6731);
nand U8577 (N_8577,N_6256,N_6438);
or U8578 (N_8578,N_6517,N_7940);
nor U8579 (N_8579,N_6977,N_6851);
nand U8580 (N_8580,N_6115,N_7295);
or U8581 (N_8581,N_7141,N_6617);
nor U8582 (N_8582,N_7945,N_6406);
and U8583 (N_8583,N_7402,N_6171);
nor U8584 (N_8584,N_6915,N_7193);
xnor U8585 (N_8585,N_6752,N_6443);
nand U8586 (N_8586,N_7796,N_7999);
xnor U8587 (N_8587,N_7015,N_7418);
nand U8588 (N_8588,N_7520,N_7787);
nor U8589 (N_8589,N_6858,N_6328);
and U8590 (N_8590,N_6313,N_7919);
or U8591 (N_8591,N_6491,N_6986);
nor U8592 (N_8592,N_7540,N_6451);
and U8593 (N_8593,N_6296,N_6028);
and U8594 (N_8594,N_7876,N_7811);
xor U8595 (N_8595,N_6805,N_6782);
or U8596 (N_8596,N_6885,N_7841);
nand U8597 (N_8597,N_7898,N_7485);
nor U8598 (N_8598,N_6505,N_6237);
or U8599 (N_8599,N_6876,N_6090);
nand U8600 (N_8600,N_6238,N_7355);
nor U8601 (N_8601,N_6248,N_7728);
nor U8602 (N_8602,N_6906,N_7692);
nor U8603 (N_8603,N_7126,N_6790);
nand U8604 (N_8604,N_6864,N_7428);
nor U8605 (N_8605,N_7804,N_7837);
xor U8606 (N_8606,N_7217,N_7695);
nand U8607 (N_8607,N_7873,N_7178);
and U8608 (N_8608,N_7924,N_6295);
xnor U8609 (N_8609,N_6621,N_6268);
and U8610 (N_8610,N_7106,N_6290);
nand U8611 (N_8611,N_7761,N_7821);
nor U8612 (N_8612,N_7164,N_6382);
nor U8613 (N_8613,N_7272,N_6708);
nand U8614 (N_8614,N_7889,N_7406);
or U8615 (N_8615,N_6713,N_6582);
or U8616 (N_8616,N_7137,N_7162);
nor U8617 (N_8617,N_6227,N_7021);
xor U8618 (N_8618,N_7471,N_6247);
or U8619 (N_8619,N_6536,N_7579);
nor U8620 (N_8620,N_7061,N_6471);
nand U8621 (N_8621,N_6738,N_7759);
or U8622 (N_8622,N_7791,N_7075);
and U8623 (N_8623,N_6085,N_7400);
and U8624 (N_8624,N_7914,N_6376);
or U8625 (N_8625,N_7734,N_7069);
and U8626 (N_8626,N_7676,N_7699);
and U8627 (N_8627,N_7130,N_7763);
and U8628 (N_8628,N_7543,N_7893);
nor U8629 (N_8629,N_6652,N_6206);
xor U8630 (N_8630,N_7257,N_7404);
and U8631 (N_8631,N_7258,N_6249);
nor U8632 (N_8632,N_7653,N_7786);
nand U8633 (N_8633,N_7823,N_7382);
and U8634 (N_8634,N_6835,N_7215);
xor U8635 (N_8635,N_7535,N_6830);
xnor U8636 (N_8636,N_7689,N_7054);
nor U8637 (N_8637,N_6815,N_6212);
and U8638 (N_8638,N_6563,N_6551);
and U8639 (N_8639,N_7711,N_7195);
nor U8640 (N_8640,N_6812,N_6689);
nor U8641 (N_8641,N_7766,N_6981);
xor U8642 (N_8642,N_7741,N_7902);
or U8643 (N_8643,N_7114,N_6000);
or U8644 (N_8644,N_7084,N_7568);
nor U8645 (N_8645,N_6230,N_7290);
nand U8646 (N_8646,N_7122,N_6849);
or U8647 (N_8647,N_6010,N_6853);
nor U8648 (N_8648,N_7697,N_7794);
or U8649 (N_8649,N_6569,N_6597);
or U8650 (N_8650,N_6068,N_7493);
xnor U8651 (N_8651,N_7197,N_7835);
nand U8652 (N_8652,N_7923,N_6221);
xor U8653 (N_8653,N_6263,N_7979);
nand U8654 (N_8654,N_6886,N_6337);
nand U8655 (N_8655,N_6523,N_6304);
and U8656 (N_8656,N_6688,N_6541);
nand U8657 (N_8657,N_6076,N_6564);
xor U8658 (N_8658,N_6634,N_6993);
nand U8659 (N_8659,N_6856,N_6978);
nand U8660 (N_8660,N_6589,N_6147);
nand U8661 (N_8661,N_7524,N_7214);
nor U8662 (N_8662,N_7216,N_7419);
and U8663 (N_8663,N_7755,N_7715);
nand U8664 (N_8664,N_6650,N_7665);
xor U8665 (N_8665,N_6190,N_6139);
nand U8666 (N_8666,N_7420,N_7266);
or U8667 (N_8667,N_7449,N_7593);
nor U8668 (N_8668,N_7634,N_6186);
nand U8669 (N_8669,N_7572,N_7236);
xor U8670 (N_8670,N_6408,N_6603);
nand U8671 (N_8671,N_7384,N_6442);
nand U8672 (N_8672,N_6219,N_7034);
nand U8673 (N_8673,N_7464,N_6765);
and U8674 (N_8674,N_6698,N_6810);
nor U8675 (N_8675,N_7815,N_7716);
and U8676 (N_8676,N_6485,N_7198);
nor U8677 (N_8677,N_6753,N_7492);
and U8678 (N_8678,N_6980,N_7531);
nor U8679 (N_8679,N_7374,N_7546);
nand U8680 (N_8680,N_7115,N_6014);
nor U8681 (N_8681,N_7598,N_7651);
nor U8682 (N_8682,N_7460,N_7933);
nor U8683 (N_8683,N_7812,N_7842);
and U8684 (N_8684,N_7853,N_7457);
or U8685 (N_8685,N_7806,N_7960);
xnor U8686 (N_8686,N_7020,N_7646);
and U8687 (N_8687,N_7961,N_7882);
nand U8688 (N_8688,N_6473,N_7062);
or U8689 (N_8689,N_6223,N_7023);
or U8690 (N_8690,N_6779,N_7864);
xor U8691 (N_8691,N_6243,N_7438);
xor U8692 (N_8692,N_6578,N_6907);
and U8693 (N_8693,N_7433,N_6039);
nand U8694 (N_8694,N_7233,N_7793);
xnor U8695 (N_8695,N_6130,N_7987);
nor U8696 (N_8696,N_6254,N_7877);
xnor U8697 (N_8697,N_6880,N_6573);
and U8698 (N_8698,N_7862,N_7685);
and U8699 (N_8699,N_6984,N_7951);
and U8700 (N_8700,N_7391,N_7396);
or U8701 (N_8701,N_7499,N_6262);
nand U8702 (N_8702,N_6518,N_6735);
nand U8703 (N_8703,N_6950,N_7304);
and U8704 (N_8704,N_7574,N_7025);
and U8705 (N_8705,N_6272,N_6935);
or U8706 (N_8706,N_6690,N_6884);
or U8707 (N_8707,N_6568,N_7479);
xnor U8708 (N_8708,N_7147,N_6257);
or U8709 (N_8709,N_6094,N_7905);
or U8710 (N_8710,N_7809,N_7401);
nor U8711 (N_8711,N_7915,N_6989);
nand U8712 (N_8712,N_7223,N_7868);
and U8713 (N_8713,N_6556,N_7188);
or U8714 (N_8714,N_7537,N_6580);
xor U8715 (N_8715,N_6200,N_6854);
nor U8716 (N_8716,N_6701,N_6641);
or U8717 (N_8717,N_6179,N_7713);
or U8718 (N_8718,N_6619,N_6023);
nand U8719 (N_8719,N_7212,N_7082);
or U8720 (N_8720,N_7595,N_6467);
nor U8721 (N_8721,N_7542,N_7200);
nand U8722 (N_8722,N_6209,N_7615);
or U8723 (N_8723,N_6182,N_6486);
nor U8724 (N_8724,N_7667,N_7398);
xor U8725 (N_8725,N_7827,N_6031);
nand U8726 (N_8726,N_7523,N_6300);
nand U8727 (N_8727,N_7978,N_7455);
nor U8728 (N_8728,N_6159,N_7139);
nand U8729 (N_8729,N_6475,N_7300);
nand U8730 (N_8730,N_6405,N_7370);
nand U8731 (N_8731,N_7163,N_7775);
or U8732 (N_8732,N_7502,N_6299);
and U8733 (N_8733,N_7285,N_6599);
or U8734 (N_8734,N_6791,N_7104);
or U8735 (N_8735,N_7089,N_7268);
and U8736 (N_8736,N_6320,N_6140);
nor U8737 (N_8737,N_7059,N_6760);
nand U8738 (N_8738,N_6842,N_6648);
xnor U8739 (N_8739,N_7769,N_7094);
or U8740 (N_8740,N_6733,N_7627);
nor U8741 (N_8741,N_6727,N_6463);
xnor U8742 (N_8742,N_7509,N_6586);
nor U8743 (N_8743,N_7354,N_6912);
nor U8744 (N_8744,N_6271,N_6303);
nor U8745 (N_8745,N_6811,N_6047);
and U8746 (N_8746,N_7340,N_7045);
xnor U8747 (N_8747,N_6121,N_6099);
nor U8748 (N_8748,N_7345,N_6127);
nand U8749 (N_8749,N_6571,N_6387);
and U8750 (N_8750,N_7928,N_7450);
or U8751 (N_8751,N_7086,N_6576);
nor U8752 (N_8752,N_7425,N_6826);
nand U8753 (N_8753,N_6788,N_7965);
nand U8754 (N_8754,N_7394,N_7291);
nand U8755 (N_8755,N_7705,N_7498);
nand U8756 (N_8756,N_6084,N_6032);
nor U8757 (N_8757,N_6259,N_7235);
or U8758 (N_8758,N_6680,N_7210);
and U8759 (N_8759,N_6493,N_7942);
nand U8760 (N_8760,N_6527,N_7444);
or U8761 (N_8761,N_6497,N_6316);
or U8762 (N_8762,N_7962,N_6503);
nand U8763 (N_8763,N_7413,N_6972);
nor U8764 (N_8764,N_6651,N_7740);
or U8765 (N_8765,N_6218,N_6535);
or U8766 (N_8766,N_7219,N_7683);
and U8767 (N_8767,N_7505,N_7143);
or U8768 (N_8768,N_7980,N_7049);
nor U8769 (N_8769,N_7781,N_7320);
xor U8770 (N_8770,N_7604,N_7445);
and U8771 (N_8771,N_6310,N_6766);
and U8772 (N_8772,N_7982,N_6101);
nor U8773 (N_8773,N_7030,N_6955);
nand U8774 (N_8774,N_7101,N_7462);
xnor U8775 (N_8775,N_6776,N_7201);
nand U8776 (N_8776,N_7230,N_7009);
xor U8777 (N_8777,N_6013,N_7981);
xor U8778 (N_8778,N_7975,N_7263);
nor U8779 (N_8779,N_7582,N_6410);
or U8780 (N_8780,N_6840,N_7897);
nand U8781 (N_8781,N_6825,N_7800);
nand U8782 (N_8782,N_6403,N_6964);
nand U8783 (N_8783,N_6274,N_7255);
xnor U8784 (N_8784,N_6168,N_6911);
and U8785 (N_8785,N_6702,N_7019);
xor U8786 (N_8786,N_6365,N_6278);
nand U8787 (N_8787,N_7819,N_6971);
nor U8788 (N_8788,N_7655,N_7330);
or U8789 (N_8789,N_6606,N_6764);
nand U8790 (N_8790,N_6317,N_6747);
nor U8791 (N_8791,N_7411,N_6575);
nor U8792 (N_8792,N_6120,N_6433);
and U8793 (N_8793,N_6795,N_6745);
nor U8794 (N_8794,N_6470,N_7426);
nor U8795 (N_8795,N_7846,N_7968);
or U8796 (N_8796,N_6165,N_6087);
and U8797 (N_8797,N_7797,N_6762);
or U8798 (N_8798,N_7865,N_7490);
and U8799 (N_8799,N_7656,N_7870);
nand U8800 (N_8800,N_7274,N_6933);
nor U8801 (N_8801,N_7512,N_6794);
nor U8802 (N_8802,N_6327,N_6952);
nor U8803 (N_8803,N_7211,N_7991);
nor U8804 (N_8804,N_7079,N_6377);
or U8805 (N_8805,N_7271,N_7844);
xor U8806 (N_8806,N_7722,N_6308);
or U8807 (N_8807,N_6996,N_7359);
or U8808 (N_8808,N_7436,N_6925);
or U8809 (N_8809,N_6929,N_7659);
nor U8810 (N_8810,N_7432,N_7532);
or U8811 (N_8811,N_7878,N_6174);
and U8812 (N_8812,N_6614,N_6345);
nor U8813 (N_8813,N_7684,N_6706);
or U8814 (N_8814,N_7073,N_6959);
xnor U8815 (N_8815,N_6205,N_6618);
nand U8816 (N_8816,N_6113,N_7622);
nor U8817 (N_8817,N_6222,N_7643);
and U8818 (N_8818,N_7481,N_7316);
or U8819 (N_8819,N_6672,N_7161);
nor U8820 (N_8820,N_6102,N_6135);
nand U8821 (N_8821,N_6872,N_7737);
nor U8822 (N_8822,N_7461,N_7725);
nand U8823 (N_8823,N_7240,N_7594);
and U8824 (N_8824,N_6703,N_7318);
xnor U8825 (N_8825,N_6434,N_7719);
nand U8826 (N_8826,N_6948,N_6349);
xnor U8827 (N_8827,N_7328,N_7289);
nand U8828 (N_8828,N_7249,N_7473);
xor U8829 (N_8829,N_6519,N_7100);
nand U8830 (N_8830,N_6226,N_7828);
nand U8831 (N_8831,N_7424,N_6392);
nand U8832 (N_8832,N_6362,N_6538);
or U8833 (N_8833,N_6657,N_6162);
nand U8834 (N_8834,N_7102,N_6833);
xnor U8835 (N_8835,N_7243,N_7640);
nor U8836 (N_8836,N_6841,N_7465);
or U8837 (N_8837,N_7253,N_7764);
and U8838 (N_8838,N_6820,N_6787);
nand U8839 (N_8839,N_7466,N_6716);
and U8840 (N_8840,N_6682,N_6217);
nor U8841 (N_8841,N_7350,N_6554);
nor U8842 (N_8842,N_7966,N_7368);
and U8843 (N_8843,N_7364,N_6088);
and U8844 (N_8844,N_6381,N_7616);
xnor U8845 (N_8845,N_6922,N_6137);
or U8846 (N_8846,N_6616,N_7206);
and U8847 (N_8847,N_7307,N_7707);
xnor U8848 (N_8848,N_6780,N_7661);
nor U8849 (N_8849,N_7922,N_6080);
nor U8850 (N_8850,N_6211,N_6801);
and U8851 (N_8851,N_6261,N_6587);
xor U8852 (N_8852,N_7988,N_6199);
and U8853 (N_8853,N_6288,N_7920);
and U8854 (N_8854,N_6035,N_6513);
and U8855 (N_8855,N_7880,N_6011);
xor U8856 (N_8856,N_6332,N_6421);
nand U8857 (N_8857,N_7237,N_6974);
and U8858 (N_8858,N_6383,N_7463);
or U8859 (N_8859,N_6630,N_6196);
nor U8860 (N_8860,N_7571,N_7052);
xor U8861 (N_8861,N_6192,N_7703);
nor U8862 (N_8862,N_7983,N_6436);
or U8863 (N_8863,N_6749,N_6710);
or U8864 (N_8864,N_6081,N_6789);
nand U8865 (N_8865,N_7605,N_6828);
or U8866 (N_8866,N_6104,N_7997);
nand U8867 (N_8867,N_6208,N_6072);
nor U8868 (N_8868,N_7247,N_7334);
or U8869 (N_8869,N_7813,N_7269);
and U8870 (N_8870,N_7468,N_6457);
and U8871 (N_8871,N_6654,N_6148);
or U8872 (N_8872,N_7026,N_6852);
nor U8873 (N_8873,N_7770,N_7559);
or U8874 (N_8874,N_6430,N_7563);
nand U8875 (N_8875,N_6330,N_7600);
xor U8876 (N_8876,N_6232,N_7967);
xor U8877 (N_8877,N_6112,N_7173);
xnor U8878 (N_8878,N_7717,N_7963);
and U8879 (N_8879,N_6721,N_6427);
nor U8880 (N_8880,N_6033,N_7058);
nand U8881 (N_8881,N_6282,N_7175);
nand U8882 (N_8882,N_6281,N_7027);
and U8883 (N_8883,N_6024,N_7529);
or U8884 (N_8884,N_6078,N_7447);
nand U8885 (N_8885,N_6472,N_7926);
or U8886 (N_8886,N_7149,N_6944);
nor U8887 (N_8887,N_7322,N_7798);
nor U8888 (N_8888,N_6846,N_6131);
nor U8889 (N_8889,N_7993,N_7227);
or U8890 (N_8890,N_6058,N_6086);
nor U8891 (N_8891,N_6803,N_7353);
and U8892 (N_8892,N_7690,N_6424);
and U8893 (N_8893,N_7856,N_6561);
or U8894 (N_8894,N_6166,N_6860);
nand U8895 (N_8895,N_6177,N_6816);
and U8896 (N_8896,N_6414,N_7814);
or U8897 (N_8897,N_6311,N_7742);
nand U8898 (N_8898,N_7287,N_7014);
and U8899 (N_8899,N_6979,N_7638);
xnor U8900 (N_8900,N_7681,N_7803);
nand U8901 (N_8901,N_7768,N_6975);
or U8902 (N_8902,N_7292,N_6740);
and U8903 (N_8903,N_7555,N_7150);
and U8904 (N_8904,N_7970,N_6315);
and U8905 (N_8905,N_7937,N_7250);
nor U8906 (N_8906,N_6015,N_7879);
or U8907 (N_8907,N_6862,N_6469);
and U8908 (N_8908,N_7549,N_6632);
or U8909 (N_8909,N_6004,N_6007);
nand U8910 (N_8910,N_7668,N_7056);
xor U8911 (N_8911,N_7944,N_7224);
and U8912 (N_8912,N_7168,N_6050);
or U8913 (N_8913,N_7379,N_6425);
nor U8914 (N_8914,N_6663,N_7753);
xnor U8915 (N_8915,N_7585,N_7564);
and U8916 (N_8916,N_7746,N_7589);
or U8917 (N_8917,N_6075,N_7228);
xnor U8918 (N_8918,N_7708,N_6678);
nor U8919 (N_8919,N_7514,N_6309);
or U8920 (N_8920,N_6250,N_7412);
and U8921 (N_8921,N_7597,N_7309);
xor U8922 (N_8922,N_6283,N_6590);
nand U8923 (N_8923,N_6695,N_6432);
or U8924 (N_8924,N_6063,N_7489);
or U8925 (N_8925,N_7246,N_7731);
xnor U8926 (N_8926,N_7861,N_7044);
nand U8927 (N_8927,N_6637,N_6718);
and U8928 (N_8928,N_6287,N_7872);
and U8929 (N_8929,N_7362,N_6732);
nor U8930 (N_8930,N_6946,N_6070);
xor U8931 (N_8931,N_7187,N_7326);
and U8932 (N_8932,N_7765,N_7022);
or U8933 (N_8933,N_6845,N_7799);
and U8934 (N_8934,N_7538,N_6750);
and U8935 (N_8935,N_7936,N_6960);
xor U8936 (N_8936,N_7958,N_7038);
or U8937 (N_8937,N_7932,N_7614);
xor U8938 (N_8938,N_7225,N_7080);
and U8939 (N_8939,N_6440,N_6049);
nand U8940 (N_8940,N_7172,N_6865);
nand U8941 (N_8941,N_6793,N_6604);
and U8942 (N_8942,N_7822,N_7459);
and U8943 (N_8943,N_6644,N_6730);
xor U8944 (N_8944,N_6988,N_6083);
xnor U8945 (N_8945,N_6134,N_7884);
and U8946 (N_8946,N_6097,N_7909);
or U8947 (N_8947,N_7688,N_6185);
nand U8948 (N_8948,N_6748,N_6235);
nand U8949 (N_8949,N_7494,N_7190);
and U8950 (N_8950,N_6743,N_6061);
nor U8951 (N_8951,N_7205,N_6334);
or U8952 (N_8952,N_7380,N_7618);
and U8953 (N_8953,N_7773,N_7323);
and U8954 (N_8954,N_7138,N_6555);
xnor U8955 (N_8955,N_6149,N_7070);
and U8956 (N_8956,N_6156,N_6511);
nor U8957 (N_8957,N_6012,N_6363);
or U8958 (N_8958,N_7331,N_7577);
xor U8959 (N_8959,N_6739,N_7801);
nor U8960 (N_8960,N_6202,N_7327);
and U8961 (N_8961,N_6394,N_7839);
or U8962 (N_8962,N_7135,N_6380);
and U8963 (N_8963,N_7435,N_7735);
or U8964 (N_8964,N_6844,N_6661);
or U8965 (N_8965,N_7159,N_6878);
nand U8966 (N_8966,N_7561,N_7299);
or U8967 (N_8967,N_6694,N_7408);
xor U8968 (N_8968,N_6931,N_6389);
nor U8969 (N_8969,N_6016,N_6079);
nand U8970 (N_8970,N_6169,N_7422);
nand U8971 (N_8971,N_7242,N_7343);
nand U8972 (N_8972,N_6524,N_6866);
xor U8973 (N_8973,N_7720,N_7381);
nand U8974 (N_8974,N_7874,N_6798);
xnor U8975 (N_8975,N_7601,N_6574);
and U8976 (N_8976,N_6170,N_6883);
nand U8977 (N_8977,N_7337,N_6500);
and U8978 (N_8978,N_7254,N_7213);
nand U8979 (N_8979,N_7994,N_6676);
nand U8980 (N_8980,N_7971,N_7311);
or U8981 (N_8981,N_7947,N_6455);
nor U8982 (N_8982,N_6161,N_6444);
or U8983 (N_8983,N_6778,N_7927);
and U8984 (N_8984,N_7679,N_7866);
xor U8985 (N_8985,N_6452,N_6528);
nand U8986 (N_8986,N_7807,N_6879);
xor U8987 (N_8987,N_7002,N_6141);
and U8988 (N_8988,N_6824,N_7777);
and U8989 (N_8989,N_7888,N_7557);
nand U8990 (N_8990,N_7776,N_6494);
nor U8991 (N_8991,N_7099,N_7721);
nand U8992 (N_8992,N_7452,N_7992);
nor U8993 (N_8993,N_7040,N_7859);
nand U8994 (N_8994,N_6359,N_6870);
or U8995 (N_8995,N_7855,N_7805);
nand U8996 (N_8996,N_6601,N_7108);
xnor U8997 (N_8997,N_6723,N_6057);
nand U8998 (N_8998,N_7996,N_6628);
nor U8999 (N_8999,N_6273,N_7151);
nor U9000 (N_9000,N_6869,N_6749);
nor U9001 (N_9001,N_6896,N_7730);
and U9002 (N_9002,N_6947,N_7423);
nor U9003 (N_9003,N_7566,N_6296);
or U9004 (N_9004,N_6791,N_7449);
nor U9005 (N_9005,N_7843,N_6163);
and U9006 (N_9006,N_6076,N_7709);
nor U9007 (N_9007,N_7621,N_7529);
xnor U9008 (N_9008,N_7213,N_7577);
and U9009 (N_9009,N_7312,N_6035);
nand U9010 (N_9010,N_7181,N_6124);
xnor U9011 (N_9011,N_6431,N_7907);
nor U9012 (N_9012,N_7315,N_7689);
or U9013 (N_9013,N_7268,N_7373);
or U9014 (N_9014,N_6734,N_6215);
and U9015 (N_9015,N_6660,N_7203);
xor U9016 (N_9016,N_6254,N_7735);
and U9017 (N_9017,N_6841,N_6388);
and U9018 (N_9018,N_6602,N_6683);
or U9019 (N_9019,N_6766,N_7175);
or U9020 (N_9020,N_6197,N_7900);
and U9021 (N_9021,N_7299,N_7962);
or U9022 (N_9022,N_7754,N_7798);
xnor U9023 (N_9023,N_6216,N_6263);
xnor U9024 (N_9024,N_6021,N_7445);
nor U9025 (N_9025,N_7843,N_7215);
nor U9026 (N_9026,N_7316,N_6600);
xnor U9027 (N_9027,N_7327,N_7797);
xnor U9028 (N_9028,N_7537,N_7906);
nand U9029 (N_9029,N_7479,N_7398);
and U9030 (N_9030,N_6502,N_7478);
and U9031 (N_9031,N_7238,N_7748);
nand U9032 (N_9032,N_7231,N_7026);
nand U9033 (N_9033,N_7114,N_7781);
nor U9034 (N_9034,N_7732,N_6006);
or U9035 (N_9035,N_6162,N_7093);
nor U9036 (N_9036,N_7960,N_7647);
xnor U9037 (N_9037,N_6322,N_6672);
xnor U9038 (N_9038,N_7693,N_7083);
nor U9039 (N_9039,N_7122,N_7677);
and U9040 (N_9040,N_7902,N_6085);
xnor U9041 (N_9041,N_7167,N_7673);
and U9042 (N_9042,N_6790,N_7895);
and U9043 (N_9043,N_7656,N_6662);
xnor U9044 (N_9044,N_6703,N_7207);
xor U9045 (N_9045,N_6052,N_7168);
nor U9046 (N_9046,N_6878,N_7575);
and U9047 (N_9047,N_6145,N_7912);
or U9048 (N_9048,N_6511,N_7360);
nor U9049 (N_9049,N_7237,N_7470);
nand U9050 (N_9050,N_6529,N_6009);
xnor U9051 (N_9051,N_7736,N_6419);
nand U9052 (N_9052,N_6859,N_7658);
xor U9053 (N_9053,N_6898,N_7583);
or U9054 (N_9054,N_6490,N_7705);
xor U9055 (N_9055,N_7616,N_7489);
and U9056 (N_9056,N_7495,N_6604);
nand U9057 (N_9057,N_6485,N_6517);
or U9058 (N_9058,N_6132,N_6357);
nand U9059 (N_9059,N_7362,N_7620);
or U9060 (N_9060,N_6801,N_7295);
or U9061 (N_9061,N_6874,N_7497);
nor U9062 (N_9062,N_6060,N_7135);
xor U9063 (N_9063,N_7674,N_6067);
nor U9064 (N_9064,N_6050,N_7173);
or U9065 (N_9065,N_6505,N_7441);
xor U9066 (N_9066,N_7611,N_6292);
xor U9067 (N_9067,N_6010,N_6157);
and U9068 (N_9068,N_7825,N_6572);
and U9069 (N_9069,N_7472,N_7805);
xnor U9070 (N_9070,N_7177,N_7939);
or U9071 (N_9071,N_6084,N_6833);
xor U9072 (N_9072,N_7429,N_7607);
xor U9073 (N_9073,N_7246,N_6656);
and U9074 (N_9074,N_6234,N_7277);
and U9075 (N_9075,N_7998,N_7945);
or U9076 (N_9076,N_6288,N_6644);
or U9077 (N_9077,N_7065,N_6563);
or U9078 (N_9078,N_6667,N_7360);
xnor U9079 (N_9079,N_6894,N_6759);
and U9080 (N_9080,N_7759,N_6457);
nor U9081 (N_9081,N_6912,N_6817);
nor U9082 (N_9082,N_7462,N_6597);
xor U9083 (N_9083,N_6651,N_7045);
nor U9084 (N_9084,N_7837,N_7722);
nor U9085 (N_9085,N_7268,N_7672);
nor U9086 (N_9086,N_7113,N_6051);
or U9087 (N_9087,N_7714,N_7886);
nor U9088 (N_9088,N_7450,N_7881);
or U9089 (N_9089,N_6939,N_6025);
nand U9090 (N_9090,N_7293,N_7849);
and U9091 (N_9091,N_6497,N_6898);
nor U9092 (N_9092,N_6865,N_7944);
nand U9093 (N_9093,N_6219,N_7362);
nand U9094 (N_9094,N_7913,N_7569);
nor U9095 (N_9095,N_7741,N_7543);
xor U9096 (N_9096,N_7484,N_6030);
xnor U9097 (N_9097,N_7029,N_6349);
and U9098 (N_9098,N_7328,N_6869);
or U9099 (N_9099,N_7883,N_7780);
nor U9100 (N_9100,N_7443,N_6307);
and U9101 (N_9101,N_6062,N_6827);
xnor U9102 (N_9102,N_6461,N_7757);
and U9103 (N_9103,N_6407,N_6334);
nor U9104 (N_9104,N_7887,N_6034);
nor U9105 (N_9105,N_6241,N_6987);
and U9106 (N_9106,N_6501,N_7442);
or U9107 (N_9107,N_7851,N_7585);
nand U9108 (N_9108,N_6474,N_7529);
xor U9109 (N_9109,N_6520,N_7313);
nor U9110 (N_9110,N_6423,N_6029);
nand U9111 (N_9111,N_6370,N_6831);
nand U9112 (N_9112,N_7237,N_6306);
nand U9113 (N_9113,N_6799,N_6807);
or U9114 (N_9114,N_7362,N_7204);
nor U9115 (N_9115,N_6234,N_7658);
or U9116 (N_9116,N_7136,N_7655);
or U9117 (N_9117,N_6459,N_6730);
nor U9118 (N_9118,N_6698,N_7940);
and U9119 (N_9119,N_7562,N_7236);
or U9120 (N_9120,N_7436,N_6461);
nor U9121 (N_9121,N_7394,N_6576);
or U9122 (N_9122,N_6202,N_7368);
nand U9123 (N_9123,N_6275,N_7182);
nand U9124 (N_9124,N_7195,N_6690);
nand U9125 (N_9125,N_6632,N_7051);
xor U9126 (N_9126,N_7896,N_7893);
nand U9127 (N_9127,N_7232,N_6587);
nor U9128 (N_9128,N_7437,N_7972);
or U9129 (N_9129,N_7520,N_7921);
and U9130 (N_9130,N_6967,N_6939);
or U9131 (N_9131,N_7206,N_7927);
or U9132 (N_9132,N_6785,N_7995);
xor U9133 (N_9133,N_7953,N_6197);
nor U9134 (N_9134,N_6718,N_7299);
xor U9135 (N_9135,N_6021,N_7652);
and U9136 (N_9136,N_7198,N_6857);
nand U9137 (N_9137,N_6759,N_6052);
xnor U9138 (N_9138,N_6369,N_7284);
xnor U9139 (N_9139,N_7791,N_6553);
nand U9140 (N_9140,N_7691,N_6437);
and U9141 (N_9141,N_6539,N_7551);
xor U9142 (N_9142,N_7301,N_7331);
nor U9143 (N_9143,N_7342,N_7638);
nand U9144 (N_9144,N_6082,N_6257);
nor U9145 (N_9145,N_6026,N_6612);
nor U9146 (N_9146,N_6674,N_6442);
or U9147 (N_9147,N_7650,N_6599);
nand U9148 (N_9148,N_6440,N_7999);
and U9149 (N_9149,N_6585,N_7892);
nor U9150 (N_9150,N_6798,N_6108);
nor U9151 (N_9151,N_6079,N_6963);
nor U9152 (N_9152,N_6590,N_7891);
nand U9153 (N_9153,N_7605,N_6845);
nand U9154 (N_9154,N_7066,N_6172);
nor U9155 (N_9155,N_6185,N_6243);
or U9156 (N_9156,N_6759,N_7712);
nand U9157 (N_9157,N_7895,N_7236);
and U9158 (N_9158,N_7485,N_6079);
and U9159 (N_9159,N_7119,N_7863);
nor U9160 (N_9160,N_7846,N_7549);
nand U9161 (N_9161,N_7329,N_6241);
nor U9162 (N_9162,N_7326,N_6762);
nor U9163 (N_9163,N_7944,N_7867);
or U9164 (N_9164,N_7253,N_6905);
nor U9165 (N_9165,N_7652,N_7254);
xnor U9166 (N_9166,N_7550,N_7159);
or U9167 (N_9167,N_6174,N_6316);
and U9168 (N_9168,N_6867,N_7838);
xnor U9169 (N_9169,N_7876,N_7484);
or U9170 (N_9170,N_7951,N_7588);
and U9171 (N_9171,N_6020,N_7073);
nand U9172 (N_9172,N_6776,N_6515);
and U9173 (N_9173,N_7999,N_7041);
nor U9174 (N_9174,N_6182,N_7761);
nand U9175 (N_9175,N_7719,N_7992);
nand U9176 (N_9176,N_6538,N_6223);
and U9177 (N_9177,N_7644,N_6932);
nor U9178 (N_9178,N_6153,N_6245);
or U9179 (N_9179,N_6579,N_7989);
nor U9180 (N_9180,N_7536,N_6927);
or U9181 (N_9181,N_6168,N_6001);
nand U9182 (N_9182,N_6874,N_6272);
nor U9183 (N_9183,N_6181,N_7301);
nor U9184 (N_9184,N_6881,N_7959);
nand U9185 (N_9185,N_7018,N_6253);
or U9186 (N_9186,N_7467,N_7882);
or U9187 (N_9187,N_6074,N_7977);
nor U9188 (N_9188,N_7778,N_6590);
xor U9189 (N_9189,N_6683,N_7240);
xnor U9190 (N_9190,N_7145,N_7302);
or U9191 (N_9191,N_6665,N_7171);
or U9192 (N_9192,N_7977,N_7700);
xor U9193 (N_9193,N_7242,N_7718);
xor U9194 (N_9194,N_6950,N_7176);
and U9195 (N_9195,N_6073,N_6859);
and U9196 (N_9196,N_6202,N_6398);
and U9197 (N_9197,N_6052,N_6004);
nand U9198 (N_9198,N_7487,N_6830);
or U9199 (N_9199,N_6949,N_6318);
and U9200 (N_9200,N_6978,N_7133);
nor U9201 (N_9201,N_7783,N_7397);
nor U9202 (N_9202,N_6071,N_7046);
nor U9203 (N_9203,N_6721,N_7859);
nand U9204 (N_9204,N_7938,N_6723);
nand U9205 (N_9205,N_6682,N_7305);
nor U9206 (N_9206,N_6918,N_7228);
or U9207 (N_9207,N_6368,N_7588);
nor U9208 (N_9208,N_7673,N_7967);
xnor U9209 (N_9209,N_6796,N_6719);
and U9210 (N_9210,N_6856,N_6049);
xnor U9211 (N_9211,N_7751,N_7437);
nor U9212 (N_9212,N_7576,N_6759);
or U9213 (N_9213,N_7031,N_6846);
xnor U9214 (N_9214,N_7280,N_7608);
nand U9215 (N_9215,N_6081,N_6359);
and U9216 (N_9216,N_6224,N_6431);
nor U9217 (N_9217,N_7821,N_7816);
nand U9218 (N_9218,N_6299,N_6558);
and U9219 (N_9219,N_7691,N_7019);
nand U9220 (N_9220,N_6833,N_7758);
nand U9221 (N_9221,N_6566,N_7911);
or U9222 (N_9222,N_7808,N_6436);
and U9223 (N_9223,N_6912,N_7508);
nand U9224 (N_9224,N_7642,N_7609);
nor U9225 (N_9225,N_7375,N_6511);
xnor U9226 (N_9226,N_6627,N_6936);
xor U9227 (N_9227,N_7521,N_6576);
or U9228 (N_9228,N_6817,N_6600);
and U9229 (N_9229,N_7245,N_7517);
and U9230 (N_9230,N_6701,N_6415);
and U9231 (N_9231,N_7111,N_7875);
xnor U9232 (N_9232,N_7796,N_6943);
and U9233 (N_9233,N_6885,N_7746);
nor U9234 (N_9234,N_6771,N_7497);
and U9235 (N_9235,N_7926,N_6268);
or U9236 (N_9236,N_6398,N_6530);
xor U9237 (N_9237,N_7663,N_7490);
or U9238 (N_9238,N_7724,N_6382);
nand U9239 (N_9239,N_6071,N_7459);
xor U9240 (N_9240,N_6552,N_7846);
nor U9241 (N_9241,N_7414,N_7831);
and U9242 (N_9242,N_7519,N_7423);
or U9243 (N_9243,N_6381,N_6372);
and U9244 (N_9244,N_6911,N_7035);
and U9245 (N_9245,N_6552,N_7633);
or U9246 (N_9246,N_6386,N_6663);
or U9247 (N_9247,N_7797,N_6458);
nor U9248 (N_9248,N_7429,N_7069);
nand U9249 (N_9249,N_6142,N_6562);
or U9250 (N_9250,N_7321,N_6633);
or U9251 (N_9251,N_7277,N_7570);
nor U9252 (N_9252,N_7506,N_7185);
and U9253 (N_9253,N_6710,N_6102);
nand U9254 (N_9254,N_7166,N_7208);
nor U9255 (N_9255,N_7920,N_6911);
and U9256 (N_9256,N_7516,N_7587);
and U9257 (N_9257,N_6674,N_6291);
nor U9258 (N_9258,N_6476,N_6732);
or U9259 (N_9259,N_7190,N_6714);
xor U9260 (N_9260,N_7305,N_7160);
and U9261 (N_9261,N_6312,N_7508);
nand U9262 (N_9262,N_6635,N_6437);
xor U9263 (N_9263,N_6865,N_6107);
nand U9264 (N_9264,N_7292,N_7021);
nor U9265 (N_9265,N_6126,N_7458);
nor U9266 (N_9266,N_6147,N_6423);
nand U9267 (N_9267,N_6747,N_6297);
and U9268 (N_9268,N_7578,N_7157);
nor U9269 (N_9269,N_6704,N_6295);
xnor U9270 (N_9270,N_6550,N_7562);
or U9271 (N_9271,N_7631,N_6538);
and U9272 (N_9272,N_7218,N_7573);
xnor U9273 (N_9273,N_7529,N_7522);
or U9274 (N_9274,N_7952,N_6406);
nor U9275 (N_9275,N_7821,N_7086);
nand U9276 (N_9276,N_6683,N_7634);
and U9277 (N_9277,N_6392,N_6731);
xor U9278 (N_9278,N_7554,N_7072);
nor U9279 (N_9279,N_6310,N_7391);
or U9280 (N_9280,N_6185,N_6389);
or U9281 (N_9281,N_6467,N_7737);
or U9282 (N_9282,N_6584,N_7041);
or U9283 (N_9283,N_7042,N_6654);
nor U9284 (N_9284,N_6159,N_7450);
or U9285 (N_9285,N_6558,N_6815);
or U9286 (N_9286,N_7891,N_6955);
nand U9287 (N_9287,N_6026,N_6669);
and U9288 (N_9288,N_7810,N_6459);
nand U9289 (N_9289,N_6905,N_7561);
xor U9290 (N_9290,N_6610,N_7616);
nor U9291 (N_9291,N_6659,N_7070);
or U9292 (N_9292,N_6633,N_6891);
nor U9293 (N_9293,N_6214,N_7408);
and U9294 (N_9294,N_6004,N_6459);
xor U9295 (N_9295,N_6112,N_6716);
nand U9296 (N_9296,N_7501,N_6113);
nor U9297 (N_9297,N_6643,N_6504);
nand U9298 (N_9298,N_7151,N_7708);
xor U9299 (N_9299,N_6226,N_6482);
xor U9300 (N_9300,N_6644,N_7075);
and U9301 (N_9301,N_6270,N_7253);
or U9302 (N_9302,N_6830,N_7260);
and U9303 (N_9303,N_7701,N_6475);
or U9304 (N_9304,N_6036,N_6597);
and U9305 (N_9305,N_7350,N_6975);
nor U9306 (N_9306,N_6501,N_7757);
nand U9307 (N_9307,N_7114,N_6234);
nand U9308 (N_9308,N_6170,N_7483);
xor U9309 (N_9309,N_6386,N_6534);
nand U9310 (N_9310,N_7197,N_7471);
and U9311 (N_9311,N_7541,N_6317);
nor U9312 (N_9312,N_7090,N_7684);
and U9313 (N_9313,N_6261,N_7870);
nand U9314 (N_9314,N_6181,N_6701);
nand U9315 (N_9315,N_6628,N_6426);
xnor U9316 (N_9316,N_6512,N_6383);
nand U9317 (N_9317,N_7255,N_6982);
xnor U9318 (N_9318,N_6393,N_7071);
xor U9319 (N_9319,N_7118,N_6630);
xnor U9320 (N_9320,N_7828,N_6922);
and U9321 (N_9321,N_7855,N_7227);
nand U9322 (N_9322,N_6674,N_6508);
nor U9323 (N_9323,N_6296,N_7375);
and U9324 (N_9324,N_7129,N_6305);
or U9325 (N_9325,N_6575,N_7020);
and U9326 (N_9326,N_6454,N_7683);
xnor U9327 (N_9327,N_6066,N_7934);
nand U9328 (N_9328,N_7660,N_7771);
and U9329 (N_9329,N_7117,N_7698);
or U9330 (N_9330,N_7426,N_6188);
nor U9331 (N_9331,N_7126,N_7211);
or U9332 (N_9332,N_6807,N_7764);
xor U9333 (N_9333,N_6350,N_6343);
nand U9334 (N_9334,N_6982,N_7208);
xnor U9335 (N_9335,N_7910,N_7275);
xor U9336 (N_9336,N_7123,N_7253);
and U9337 (N_9337,N_7345,N_7519);
nand U9338 (N_9338,N_6304,N_7371);
nand U9339 (N_9339,N_6136,N_6470);
nand U9340 (N_9340,N_7564,N_6096);
nor U9341 (N_9341,N_6623,N_6548);
nor U9342 (N_9342,N_7205,N_7941);
nor U9343 (N_9343,N_6783,N_6569);
or U9344 (N_9344,N_7872,N_7151);
nor U9345 (N_9345,N_7502,N_6727);
nand U9346 (N_9346,N_6645,N_7928);
nor U9347 (N_9347,N_7401,N_6121);
and U9348 (N_9348,N_6721,N_6600);
or U9349 (N_9349,N_6311,N_6909);
nor U9350 (N_9350,N_7257,N_7168);
nor U9351 (N_9351,N_6988,N_7356);
xor U9352 (N_9352,N_7798,N_7426);
nor U9353 (N_9353,N_6982,N_7569);
and U9354 (N_9354,N_7658,N_6066);
nand U9355 (N_9355,N_7874,N_7755);
or U9356 (N_9356,N_7934,N_7377);
or U9357 (N_9357,N_6145,N_6343);
or U9358 (N_9358,N_6130,N_6213);
nand U9359 (N_9359,N_7922,N_6567);
nand U9360 (N_9360,N_7135,N_7226);
and U9361 (N_9361,N_6389,N_6911);
and U9362 (N_9362,N_6302,N_7530);
nand U9363 (N_9363,N_6792,N_6661);
or U9364 (N_9364,N_6924,N_7453);
or U9365 (N_9365,N_6443,N_6556);
and U9366 (N_9366,N_7266,N_6911);
or U9367 (N_9367,N_6910,N_7403);
xor U9368 (N_9368,N_6343,N_7656);
nand U9369 (N_9369,N_6398,N_7335);
nand U9370 (N_9370,N_7837,N_6856);
nor U9371 (N_9371,N_7689,N_6557);
or U9372 (N_9372,N_6936,N_6843);
or U9373 (N_9373,N_6014,N_7467);
and U9374 (N_9374,N_6530,N_6230);
xnor U9375 (N_9375,N_7928,N_7186);
nand U9376 (N_9376,N_7429,N_7373);
xnor U9377 (N_9377,N_7777,N_7925);
or U9378 (N_9378,N_6815,N_7254);
nand U9379 (N_9379,N_7454,N_6384);
or U9380 (N_9380,N_7580,N_6905);
or U9381 (N_9381,N_7467,N_6472);
or U9382 (N_9382,N_7705,N_6938);
nand U9383 (N_9383,N_7452,N_7365);
and U9384 (N_9384,N_6168,N_7909);
and U9385 (N_9385,N_6836,N_7512);
xnor U9386 (N_9386,N_6883,N_7787);
nor U9387 (N_9387,N_6857,N_6610);
nor U9388 (N_9388,N_6158,N_7257);
nor U9389 (N_9389,N_6201,N_7697);
xnor U9390 (N_9390,N_7225,N_6066);
xor U9391 (N_9391,N_7079,N_7873);
and U9392 (N_9392,N_7430,N_7823);
nor U9393 (N_9393,N_7251,N_7473);
and U9394 (N_9394,N_6520,N_6926);
and U9395 (N_9395,N_6202,N_7202);
xor U9396 (N_9396,N_6745,N_7389);
nor U9397 (N_9397,N_7027,N_7044);
and U9398 (N_9398,N_7976,N_6156);
or U9399 (N_9399,N_6465,N_6064);
and U9400 (N_9400,N_7030,N_6506);
xnor U9401 (N_9401,N_6286,N_7413);
xnor U9402 (N_9402,N_6906,N_7162);
xnor U9403 (N_9403,N_6187,N_7349);
nand U9404 (N_9404,N_6229,N_6981);
nand U9405 (N_9405,N_6682,N_6590);
nor U9406 (N_9406,N_7276,N_7502);
and U9407 (N_9407,N_7186,N_6712);
nor U9408 (N_9408,N_7131,N_7320);
and U9409 (N_9409,N_6011,N_7063);
nand U9410 (N_9410,N_6624,N_7924);
nor U9411 (N_9411,N_6344,N_7738);
xnor U9412 (N_9412,N_7179,N_6822);
and U9413 (N_9413,N_7807,N_6284);
and U9414 (N_9414,N_6002,N_7164);
or U9415 (N_9415,N_7833,N_7443);
and U9416 (N_9416,N_7274,N_7270);
nor U9417 (N_9417,N_6729,N_7707);
or U9418 (N_9418,N_6802,N_6024);
and U9419 (N_9419,N_6611,N_7111);
nand U9420 (N_9420,N_7205,N_6669);
and U9421 (N_9421,N_7098,N_7592);
or U9422 (N_9422,N_6032,N_6282);
nand U9423 (N_9423,N_6935,N_6492);
xnor U9424 (N_9424,N_7881,N_7082);
xor U9425 (N_9425,N_6174,N_6874);
or U9426 (N_9426,N_6449,N_7430);
or U9427 (N_9427,N_6662,N_7740);
xnor U9428 (N_9428,N_7404,N_7461);
nor U9429 (N_9429,N_6087,N_6422);
nor U9430 (N_9430,N_7223,N_7973);
and U9431 (N_9431,N_7174,N_7375);
or U9432 (N_9432,N_6130,N_6402);
and U9433 (N_9433,N_7139,N_7827);
and U9434 (N_9434,N_7262,N_7149);
xnor U9435 (N_9435,N_6959,N_6726);
nand U9436 (N_9436,N_7051,N_6293);
nor U9437 (N_9437,N_6783,N_7354);
and U9438 (N_9438,N_7637,N_7040);
nor U9439 (N_9439,N_6957,N_7879);
nand U9440 (N_9440,N_6895,N_7595);
and U9441 (N_9441,N_7518,N_7890);
and U9442 (N_9442,N_6715,N_6606);
xor U9443 (N_9443,N_6208,N_6631);
and U9444 (N_9444,N_7967,N_6567);
xnor U9445 (N_9445,N_6498,N_6265);
or U9446 (N_9446,N_6383,N_7813);
or U9447 (N_9447,N_7994,N_6481);
nand U9448 (N_9448,N_7724,N_7828);
xor U9449 (N_9449,N_7523,N_7146);
nand U9450 (N_9450,N_6573,N_6339);
xnor U9451 (N_9451,N_7486,N_6004);
nand U9452 (N_9452,N_6467,N_7258);
nor U9453 (N_9453,N_7200,N_6979);
nor U9454 (N_9454,N_7234,N_6823);
nor U9455 (N_9455,N_6576,N_6632);
nor U9456 (N_9456,N_6001,N_7366);
and U9457 (N_9457,N_6052,N_6244);
or U9458 (N_9458,N_6568,N_7192);
nand U9459 (N_9459,N_7021,N_6066);
or U9460 (N_9460,N_6876,N_7994);
and U9461 (N_9461,N_7693,N_6049);
xnor U9462 (N_9462,N_7915,N_6173);
and U9463 (N_9463,N_6876,N_7102);
xor U9464 (N_9464,N_6784,N_6409);
nor U9465 (N_9465,N_7569,N_7831);
or U9466 (N_9466,N_7154,N_7885);
xnor U9467 (N_9467,N_7720,N_7589);
nor U9468 (N_9468,N_6158,N_7844);
nor U9469 (N_9469,N_7817,N_6262);
and U9470 (N_9470,N_7411,N_7353);
and U9471 (N_9471,N_6263,N_6066);
and U9472 (N_9472,N_6986,N_6722);
xor U9473 (N_9473,N_7504,N_7008);
and U9474 (N_9474,N_6010,N_6005);
nor U9475 (N_9475,N_7414,N_7178);
xnor U9476 (N_9476,N_6154,N_6178);
nand U9477 (N_9477,N_7428,N_6684);
xnor U9478 (N_9478,N_7101,N_7937);
or U9479 (N_9479,N_7773,N_6856);
xor U9480 (N_9480,N_6198,N_6365);
nand U9481 (N_9481,N_6928,N_6431);
nor U9482 (N_9482,N_7127,N_7666);
nand U9483 (N_9483,N_6578,N_7703);
nand U9484 (N_9484,N_6976,N_7901);
nand U9485 (N_9485,N_7686,N_7234);
or U9486 (N_9486,N_6396,N_6342);
and U9487 (N_9487,N_7588,N_6852);
and U9488 (N_9488,N_7792,N_6008);
and U9489 (N_9489,N_7503,N_6065);
xor U9490 (N_9490,N_6687,N_6078);
xor U9491 (N_9491,N_7193,N_6922);
nor U9492 (N_9492,N_6652,N_6674);
and U9493 (N_9493,N_7583,N_7223);
or U9494 (N_9494,N_7410,N_7261);
nor U9495 (N_9495,N_7019,N_6617);
nand U9496 (N_9496,N_6906,N_7655);
xor U9497 (N_9497,N_7812,N_6402);
xor U9498 (N_9498,N_6196,N_7391);
nor U9499 (N_9499,N_7083,N_6245);
nor U9500 (N_9500,N_7429,N_7511);
and U9501 (N_9501,N_6651,N_7912);
or U9502 (N_9502,N_6139,N_7699);
nor U9503 (N_9503,N_7407,N_6589);
nor U9504 (N_9504,N_6292,N_7268);
and U9505 (N_9505,N_7352,N_7319);
nor U9506 (N_9506,N_7018,N_7948);
nor U9507 (N_9507,N_6410,N_7306);
or U9508 (N_9508,N_7861,N_7750);
nor U9509 (N_9509,N_7656,N_7330);
nor U9510 (N_9510,N_6205,N_7413);
or U9511 (N_9511,N_6859,N_6934);
xor U9512 (N_9512,N_6689,N_7739);
or U9513 (N_9513,N_7845,N_6210);
and U9514 (N_9514,N_7876,N_7312);
nand U9515 (N_9515,N_6996,N_6831);
or U9516 (N_9516,N_7320,N_7153);
nand U9517 (N_9517,N_6026,N_7579);
and U9518 (N_9518,N_6304,N_7640);
and U9519 (N_9519,N_6499,N_7905);
or U9520 (N_9520,N_7639,N_7613);
or U9521 (N_9521,N_6542,N_6210);
nor U9522 (N_9522,N_7488,N_7746);
nor U9523 (N_9523,N_6785,N_6555);
or U9524 (N_9524,N_7368,N_6701);
and U9525 (N_9525,N_7739,N_7949);
nor U9526 (N_9526,N_7730,N_6153);
nor U9527 (N_9527,N_7940,N_7625);
nor U9528 (N_9528,N_7960,N_7535);
nor U9529 (N_9529,N_7714,N_6506);
xor U9530 (N_9530,N_6002,N_6284);
xnor U9531 (N_9531,N_7914,N_6919);
xor U9532 (N_9532,N_6429,N_6613);
nor U9533 (N_9533,N_7732,N_6950);
and U9534 (N_9534,N_6675,N_7204);
or U9535 (N_9535,N_6354,N_7376);
or U9536 (N_9536,N_7044,N_7969);
and U9537 (N_9537,N_7171,N_6927);
xnor U9538 (N_9538,N_7508,N_7165);
or U9539 (N_9539,N_6293,N_7431);
nand U9540 (N_9540,N_6977,N_7579);
nor U9541 (N_9541,N_7256,N_6104);
nand U9542 (N_9542,N_7741,N_6497);
and U9543 (N_9543,N_7084,N_6737);
nand U9544 (N_9544,N_7712,N_6449);
and U9545 (N_9545,N_6463,N_7898);
or U9546 (N_9546,N_6159,N_6622);
and U9547 (N_9547,N_7671,N_6265);
xor U9548 (N_9548,N_6053,N_6111);
nand U9549 (N_9549,N_6406,N_6378);
xor U9550 (N_9550,N_6245,N_7856);
xnor U9551 (N_9551,N_6793,N_7177);
and U9552 (N_9552,N_6936,N_6341);
xnor U9553 (N_9553,N_6771,N_7193);
or U9554 (N_9554,N_6954,N_6716);
or U9555 (N_9555,N_7950,N_6664);
nor U9556 (N_9556,N_6033,N_6213);
or U9557 (N_9557,N_6389,N_7650);
or U9558 (N_9558,N_7121,N_6390);
nor U9559 (N_9559,N_6617,N_7200);
nand U9560 (N_9560,N_7532,N_6285);
nor U9561 (N_9561,N_6459,N_7150);
nor U9562 (N_9562,N_6371,N_7294);
or U9563 (N_9563,N_6165,N_7934);
xnor U9564 (N_9564,N_6536,N_7266);
or U9565 (N_9565,N_7461,N_6478);
xor U9566 (N_9566,N_6176,N_6411);
and U9567 (N_9567,N_6967,N_7727);
xor U9568 (N_9568,N_7582,N_7586);
or U9569 (N_9569,N_7363,N_7459);
nor U9570 (N_9570,N_7269,N_6218);
nand U9571 (N_9571,N_6865,N_7196);
nand U9572 (N_9572,N_6497,N_6852);
nand U9573 (N_9573,N_6031,N_6167);
nand U9574 (N_9574,N_7368,N_6656);
nand U9575 (N_9575,N_6834,N_6832);
nand U9576 (N_9576,N_6284,N_7454);
nand U9577 (N_9577,N_6632,N_7136);
xnor U9578 (N_9578,N_6619,N_7390);
nor U9579 (N_9579,N_6235,N_7461);
nor U9580 (N_9580,N_7175,N_7881);
nand U9581 (N_9581,N_6334,N_7340);
or U9582 (N_9582,N_7677,N_6995);
nand U9583 (N_9583,N_6811,N_7218);
and U9584 (N_9584,N_6919,N_6494);
or U9585 (N_9585,N_6377,N_6994);
xor U9586 (N_9586,N_6607,N_7561);
xor U9587 (N_9587,N_6750,N_6339);
nor U9588 (N_9588,N_7139,N_7982);
and U9589 (N_9589,N_6981,N_7717);
xnor U9590 (N_9590,N_6193,N_6921);
nand U9591 (N_9591,N_7167,N_6336);
and U9592 (N_9592,N_6844,N_6317);
and U9593 (N_9593,N_7423,N_7662);
nand U9594 (N_9594,N_7595,N_6843);
nand U9595 (N_9595,N_6884,N_6473);
and U9596 (N_9596,N_6777,N_6510);
xor U9597 (N_9597,N_6280,N_7381);
nor U9598 (N_9598,N_7401,N_6253);
or U9599 (N_9599,N_6319,N_7901);
xnor U9600 (N_9600,N_7739,N_7258);
nor U9601 (N_9601,N_7455,N_6920);
xor U9602 (N_9602,N_6684,N_7154);
nand U9603 (N_9603,N_6777,N_7076);
nor U9604 (N_9604,N_6388,N_6073);
or U9605 (N_9605,N_7328,N_7412);
nor U9606 (N_9606,N_6966,N_7039);
and U9607 (N_9607,N_7538,N_6035);
xnor U9608 (N_9608,N_6878,N_6232);
xnor U9609 (N_9609,N_7133,N_6332);
nor U9610 (N_9610,N_7289,N_7569);
nor U9611 (N_9611,N_7726,N_6966);
and U9612 (N_9612,N_7193,N_7248);
nand U9613 (N_9613,N_6469,N_7251);
xor U9614 (N_9614,N_7560,N_7241);
nor U9615 (N_9615,N_7467,N_6616);
and U9616 (N_9616,N_6253,N_7048);
nand U9617 (N_9617,N_6701,N_6649);
xnor U9618 (N_9618,N_7107,N_7584);
nand U9619 (N_9619,N_7652,N_7232);
and U9620 (N_9620,N_6418,N_7389);
nand U9621 (N_9621,N_6421,N_6486);
nor U9622 (N_9622,N_6388,N_7759);
and U9623 (N_9623,N_7010,N_6204);
nand U9624 (N_9624,N_7537,N_7626);
xor U9625 (N_9625,N_6711,N_6839);
and U9626 (N_9626,N_7317,N_6775);
and U9627 (N_9627,N_7508,N_7390);
and U9628 (N_9628,N_7384,N_6626);
nor U9629 (N_9629,N_7643,N_7383);
xnor U9630 (N_9630,N_6036,N_7834);
nand U9631 (N_9631,N_6450,N_7585);
nand U9632 (N_9632,N_7509,N_6561);
and U9633 (N_9633,N_6026,N_7230);
nand U9634 (N_9634,N_6111,N_7102);
or U9635 (N_9635,N_7114,N_6774);
and U9636 (N_9636,N_7055,N_7856);
nor U9637 (N_9637,N_7635,N_7339);
and U9638 (N_9638,N_6567,N_6436);
and U9639 (N_9639,N_7486,N_6577);
and U9640 (N_9640,N_7345,N_7386);
nand U9641 (N_9641,N_7498,N_6536);
xnor U9642 (N_9642,N_6186,N_6033);
nor U9643 (N_9643,N_7258,N_7611);
and U9644 (N_9644,N_6782,N_7656);
xnor U9645 (N_9645,N_6645,N_7135);
nor U9646 (N_9646,N_6798,N_7378);
or U9647 (N_9647,N_7679,N_6742);
nand U9648 (N_9648,N_7893,N_7355);
and U9649 (N_9649,N_7638,N_6552);
and U9650 (N_9650,N_7287,N_6523);
nand U9651 (N_9651,N_7128,N_6548);
xnor U9652 (N_9652,N_6156,N_7520);
and U9653 (N_9653,N_6281,N_7274);
nor U9654 (N_9654,N_6163,N_6107);
xnor U9655 (N_9655,N_7092,N_6999);
and U9656 (N_9656,N_7079,N_6081);
xor U9657 (N_9657,N_7290,N_7493);
xor U9658 (N_9658,N_7292,N_6329);
xnor U9659 (N_9659,N_7890,N_6813);
nand U9660 (N_9660,N_6166,N_6789);
nand U9661 (N_9661,N_7218,N_6707);
xnor U9662 (N_9662,N_6510,N_6233);
nand U9663 (N_9663,N_7007,N_7240);
nand U9664 (N_9664,N_7661,N_7070);
nor U9665 (N_9665,N_6850,N_7808);
nand U9666 (N_9666,N_6345,N_6249);
xor U9667 (N_9667,N_6121,N_7807);
and U9668 (N_9668,N_6361,N_6938);
or U9669 (N_9669,N_6971,N_6628);
xor U9670 (N_9670,N_7552,N_7961);
xnor U9671 (N_9671,N_7733,N_7209);
and U9672 (N_9672,N_6259,N_6095);
or U9673 (N_9673,N_7548,N_7317);
and U9674 (N_9674,N_6033,N_7166);
nor U9675 (N_9675,N_7389,N_6823);
nand U9676 (N_9676,N_6004,N_7439);
and U9677 (N_9677,N_7642,N_6860);
xor U9678 (N_9678,N_6797,N_6686);
or U9679 (N_9679,N_7243,N_7183);
nor U9680 (N_9680,N_6567,N_6447);
xor U9681 (N_9681,N_7976,N_7525);
and U9682 (N_9682,N_7828,N_7173);
nand U9683 (N_9683,N_6666,N_7603);
xnor U9684 (N_9684,N_7928,N_6506);
nor U9685 (N_9685,N_7257,N_6458);
nand U9686 (N_9686,N_7687,N_7083);
or U9687 (N_9687,N_6823,N_7964);
xnor U9688 (N_9688,N_7786,N_7598);
nor U9689 (N_9689,N_6610,N_6835);
and U9690 (N_9690,N_7817,N_7474);
or U9691 (N_9691,N_7013,N_7104);
nand U9692 (N_9692,N_6175,N_6354);
or U9693 (N_9693,N_6729,N_7940);
nand U9694 (N_9694,N_6360,N_6778);
nor U9695 (N_9695,N_6099,N_6517);
and U9696 (N_9696,N_7389,N_7346);
nand U9697 (N_9697,N_6129,N_7293);
and U9698 (N_9698,N_7769,N_6975);
nor U9699 (N_9699,N_7089,N_6713);
and U9700 (N_9700,N_6665,N_7245);
and U9701 (N_9701,N_7306,N_6638);
xnor U9702 (N_9702,N_7758,N_7267);
xor U9703 (N_9703,N_6590,N_7249);
and U9704 (N_9704,N_6296,N_6749);
nor U9705 (N_9705,N_6478,N_6172);
xnor U9706 (N_9706,N_7300,N_6776);
or U9707 (N_9707,N_6505,N_6104);
nand U9708 (N_9708,N_7755,N_7855);
and U9709 (N_9709,N_7713,N_7087);
or U9710 (N_9710,N_6807,N_7002);
xnor U9711 (N_9711,N_7961,N_7487);
xor U9712 (N_9712,N_6786,N_7118);
xor U9713 (N_9713,N_7972,N_7297);
nor U9714 (N_9714,N_6004,N_6380);
nand U9715 (N_9715,N_6885,N_7595);
and U9716 (N_9716,N_6955,N_7816);
or U9717 (N_9717,N_7557,N_6560);
nor U9718 (N_9718,N_6100,N_7994);
nor U9719 (N_9719,N_7071,N_6441);
or U9720 (N_9720,N_6331,N_7000);
nor U9721 (N_9721,N_6141,N_7369);
nand U9722 (N_9722,N_7779,N_6444);
xor U9723 (N_9723,N_7365,N_7380);
nor U9724 (N_9724,N_7533,N_6506);
xor U9725 (N_9725,N_7891,N_7552);
nor U9726 (N_9726,N_6710,N_6261);
nor U9727 (N_9727,N_7587,N_7450);
nand U9728 (N_9728,N_6098,N_6290);
and U9729 (N_9729,N_6077,N_7526);
nand U9730 (N_9730,N_7618,N_6557);
xnor U9731 (N_9731,N_7395,N_7620);
nor U9732 (N_9732,N_6902,N_7254);
xor U9733 (N_9733,N_6873,N_6774);
nand U9734 (N_9734,N_6494,N_6778);
and U9735 (N_9735,N_7869,N_7026);
or U9736 (N_9736,N_7123,N_7723);
nor U9737 (N_9737,N_6044,N_6773);
xor U9738 (N_9738,N_6378,N_7849);
and U9739 (N_9739,N_7331,N_6556);
nor U9740 (N_9740,N_6913,N_6628);
and U9741 (N_9741,N_6303,N_6711);
and U9742 (N_9742,N_6447,N_6689);
xnor U9743 (N_9743,N_6045,N_7447);
nand U9744 (N_9744,N_6616,N_7834);
nor U9745 (N_9745,N_7947,N_7366);
nor U9746 (N_9746,N_7518,N_6391);
nor U9747 (N_9747,N_6239,N_6125);
xnor U9748 (N_9748,N_6951,N_6020);
nand U9749 (N_9749,N_6786,N_7827);
nand U9750 (N_9750,N_7308,N_6899);
nor U9751 (N_9751,N_6047,N_7222);
xnor U9752 (N_9752,N_7708,N_6212);
nand U9753 (N_9753,N_6365,N_6017);
or U9754 (N_9754,N_7260,N_7104);
nand U9755 (N_9755,N_6976,N_7527);
nand U9756 (N_9756,N_7730,N_7413);
nand U9757 (N_9757,N_7358,N_7725);
and U9758 (N_9758,N_7580,N_7329);
nor U9759 (N_9759,N_7008,N_6669);
or U9760 (N_9760,N_7933,N_7224);
and U9761 (N_9761,N_7354,N_7662);
nor U9762 (N_9762,N_6620,N_6958);
nand U9763 (N_9763,N_7508,N_7870);
xnor U9764 (N_9764,N_6906,N_6289);
and U9765 (N_9765,N_6941,N_6236);
nand U9766 (N_9766,N_7357,N_7054);
and U9767 (N_9767,N_6706,N_6908);
xor U9768 (N_9768,N_7740,N_7669);
or U9769 (N_9769,N_6235,N_7866);
xor U9770 (N_9770,N_7525,N_6559);
and U9771 (N_9771,N_7038,N_7834);
nor U9772 (N_9772,N_6553,N_6358);
nand U9773 (N_9773,N_7559,N_7797);
nand U9774 (N_9774,N_6634,N_6566);
and U9775 (N_9775,N_6222,N_7145);
nor U9776 (N_9776,N_6077,N_6073);
and U9777 (N_9777,N_7091,N_7586);
xnor U9778 (N_9778,N_7217,N_6366);
and U9779 (N_9779,N_6712,N_6250);
xor U9780 (N_9780,N_7217,N_6094);
xnor U9781 (N_9781,N_6016,N_7587);
or U9782 (N_9782,N_6628,N_6093);
and U9783 (N_9783,N_7365,N_7510);
xor U9784 (N_9784,N_6147,N_7729);
xor U9785 (N_9785,N_6433,N_6177);
or U9786 (N_9786,N_6024,N_6392);
nand U9787 (N_9787,N_7718,N_7909);
nor U9788 (N_9788,N_6349,N_7640);
nand U9789 (N_9789,N_6652,N_6439);
and U9790 (N_9790,N_6339,N_7772);
and U9791 (N_9791,N_7512,N_7298);
nand U9792 (N_9792,N_7931,N_7794);
nand U9793 (N_9793,N_7532,N_7680);
xor U9794 (N_9794,N_7173,N_7660);
and U9795 (N_9795,N_6516,N_7232);
nor U9796 (N_9796,N_7372,N_7025);
xnor U9797 (N_9797,N_7800,N_7538);
or U9798 (N_9798,N_7714,N_6153);
nand U9799 (N_9799,N_7672,N_6141);
nor U9800 (N_9800,N_7561,N_7011);
xor U9801 (N_9801,N_6662,N_6919);
or U9802 (N_9802,N_7815,N_6182);
or U9803 (N_9803,N_7002,N_7866);
or U9804 (N_9804,N_6968,N_6301);
or U9805 (N_9805,N_7421,N_6756);
nand U9806 (N_9806,N_7933,N_6101);
or U9807 (N_9807,N_7664,N_7774);
or U9808 (N_9808,N_6245,N_6790);
or U9809 (N_9809,N_6666,N_7417);
or U9810 (N_9810,N_7717,N_6761);
and U9811 (N_9811,N_7706,N_7431);
nor U9812 (N_9812,N_6698,N_6788);
nor U9813 (N_9813,N_6965,N_6880);
and U9814 (N_9814,N_7786,N_7628);
nand U9815 (N_9815,N_7822,N_6715);
xor U9816 (N_9816,N_7564,N_6577);
or U9817 (N_9817,N_6938,N_7799);
and U9818 (N_9818,N_7311,N_7718);
xor U9819 (N_9819,N_7244,N_6554);
nand U9820 (N_9820,N_6677,N_7100);
and U9821 (N_9821,N_6108,N_7664);
nand U9822 (N_9822,N_7171,N_7607);
nor U9823 (N_9823,N_6575,N_7989);
xnor U9824 (N_9824,N_6314,N_6681);
nand U9825 (N_9825,N_6845,N_7658);
nand U9826 (N_9826,N_7179,N_6688);
and U9827 (N_9827,N_7694,N_6697);
nor U9828 (N_9828,N_6769,N_6320);
or U9829 (N_9829,N_7044,N_6493);
and U9830 (N_9830,N_6720,N_7143);
and U9831 (N_9831,N_6956,N_6965);
nand U9832 (N_9832,N_6343,N_7323);
nand U9833 (N_9833,N_6078,N_6510);
or U9834 (N_9834,N_7417,N_7193);
xor U9835 (N_9835,N_6881,N_6394);
nor U9836 (N_9836,N_6680,N_7468);
xnor U9837 (N_9837,N_6108,N_6697);
and U9838 (N_9838,N_7267,N_6910);
xnor U9839 (N_9839,N_7380,N_7457);
and U9840 (N_9840,N_6464,N_6882);
nand U9841 (N_9841,N_7043,N_6361);
and U9842 (N_9842,N_6174,N_7267);
nand U9843 (N_9843,N_6807,N_7323);
nor U9844 (N_9844,N_7066,N_6816);
xor U9845 (N_9845,N_6058,N_6254);
or U9846 (N_9846,N_6818,N_6900);
and U9847 (N_9847,N_6657,N_7358);
nand U9848 (N_9848,N_6360,N_7260);
nand U9849 (N_9849,N_6603,N_6190);
and U9850 (N_9850,N_6289,N_7007);
nor U9851 (N_9851,N_7201,N_7774);
and U9852 (N_9852,N_6112,N_6882);
xor U9853 (N_9853,N_6955,N_6918);
and U9854 (N_9854,N_7666,N_6285);
xnor U9855 (N_9855,N_7876,N_6436);
xnor U9856 (N_9856,N_6315,N_6346);
xor U9857 (N_9857,N_7111,N_7545);
nor U9858 (N_9858,N_7857,N_7568);
nand U9859 (N_9859,N_7025,N_7166);
nor U9860 (N_9860,N_6450,N_6006);
nor U9861 (N_9861,N_6470,N_7713);
or U9862 (N_9862,N_7754,N_7034);
nand U9863 (N_9863,N_6749,N_6243);
nor U9864 (N_9864,N_7699,N_6664);
nand U9865 (N_9865,N_7605,N_7666);
or U9866 (N_9866,N_6598,N_6190);
xnor U9867 (N_9867,N_7429,N_6926);
xnor U9868 (N_9868,N_6285,N_7184);
and U9869 (N_9869,N_7584,N_6025);
and U9870 (N_9870,N_6071,N_6881);
and U9871 (N_9871,N_7470,N_7835);
xnor U9872 (N_9872,N_7412,N_6940);
or U9873 (N_9873,N_7090,N_6688);
xor U9874 (N_9874,N_7776,N_7439);
nor U9875 (N_9875,N_7658,N_7015);
nand U9876 (N_9876,N_7027,N_7191);
and U9877 (N_9877,N_7840,N_6727);
xor U9878 (N_9878,N_7326,N_7584);
nor U9879 (N_9879,N_7680,N_6705);
and U9880 (N_9880,N_6169,N_7541);
xor U9881 (N_9881,N_7696,N_7456);
xor U9882 (N_9882,N_7789,N_7934);
nor U9883 (N_9883,N_6838,N_6694);
or U9884 (N_9884,N_7047,N_7629);
nor U9885 (N_9885,N_6905,N_6050);
and U9886 (N_9886,N_7253,N_6790);
nand U9887 (N_9887,N_6858,N_6802);
or U9888 (N_9888,N_7863,N_7156);
and U9889 (N_9889,N_7239,N_6067);
nor U9890 (N_9890,N_6298,N_7586);
xnor U9891 (N_9891,N_7691,N_6800);
nand U9892 (N_9892,N_6661,N_7802);
nor U9893 (N_9893,N_7553,N_6187);
nand U9894 (N_9894,N_6806,N_6635);
or U9895 (N_9895,N_7718,N_7218);
nand U9896 (N_9896,N_7893,N_6299);
nand U9897 (N_9897,N_6130,N_6304);
xnor U9898 (N_9898,N_7239,N_6251);
nor U9899 (N_9899,N_6593,N_6655);
nand U9900 (N_9900,N_7556,N_6824);
xor U9901 (N_9901,N_7334,N_7918);
nor U9902 (N_9902,N_6208,N_7678);
nor U9903 (N_9903,N_7256,N_7886);
xnor U9904 (N_9904,N_6866,N_6471);
and U9905 (N_9905,N_7623,N_6713);
nor U9906 (N_9906,N_7693,N_7928);
xnor U9907 (N_9907,N_7933,N_7714);
xnor U9908 (N_9908,N_7034,N_6972);
nor U9909 (N_9909,N_7710,N_7160);
or U9910 (N_9910,N_7426,N_6392);
xnor U9911 (N_9911,N_7023,N_7223);
nand U9912 (N_9912,N_6634,N_7414);
and U9913 (N_9913,N_7684,N_7999);
nand U9914 (N_9914,N_7397,N_6547);
nor U9915 (N_9915,N_6036,N_6429);
or U9916 (N_9916,N_6267,N_6567);
or U9917 (N_9917,N_6702,N_6564);
and U9918 (N_9918,N_7515,N_6585);
xnor U9919 (N_9919,N_7884,N_7495);
nand U9920 (N_9920,N_7811,N_6131);
xnor U9921 (N_9921,N_6600,N_6459);
nand U9922 (N_9922,N_7707,N_6340);
nor U9923 (N_9923,N_6880,N_7893);
nand U9924 (N_9924,N_7111,N_6159);
nor U9925 (N_9925,N_6585,N_7117);
and U9926 (N_9926,N_6368,N_7666);
xnor U9927 (N_9927,N_7961,N_6734);
and U9928 (N_9928,N_6807,N_7717);
xnor U9929 (N_9929,N_7978,N_7987);
or U9930 (N_9930,N_6091,N_6959);
and U9931 (N_9931,N_7292,N_7385);
or U9932 (N_9932,N_6388,N_7527);
nand U9933 (N_9933,N_7404,N_7144);
nor U9934 (N_9934,N_7761,N_7341);
nand U9935 (N_9935,N_6065,N_7379);
and U9936 (N_9936,N_6343,N_7840);
nor U9937 (N_9937,N_7500,N_6097);
xnor U9938 (N_9938,N_7144,N_7336);
xnor U9939 (N_9939,N_6114,N_7208);
nor U9940 (N_9940,N_7093,N_7462);
and U9941 (N_9941,N_7003,N_6955);
or U9942 (N_9942,N_7841,N_7246);
and U9943 (N_9943,N_7655,N_6826);
or U9944 (N_9944,N_7533,N_6578);
nand U9945 (N_9945,N_7004,N_7495);
and U9946 (N_9946,N_6255,N_6768);
or U9947 (N_9947,N_7264,N_7816);
xnor U9948 (N_9948,N_7964,N_7209);
xnor U9949 (N_9949,N_6386,N_6192);
nand U9950 (N_9950,N_7703,N_6605);
nand U9951 (N_9951,N_6438,N_6752);
nand U9952 (N_9952,N_6560,N_7586);
nand U9953 (N_9953,N_6694,N_6942);
and U9954 (N_9954,N_6929,N_6802);
or U9955 (N_9955,N_7819,N_7412);
nand U9956 (N_9956,N_7649,N_7594);
or U9957 (N_9957,N_7458,N_6571);
xor U9958 (N_9958,N_7798,N_7871);
xor U9959 (N_9959,N_7036,N_6001);
nand U9960 (N_9960,N_6338,N_6893);
xnor U9961 (N_9961,N_6840,N_7329);
nand U9962 (N_9962,N_7667,N_7479);
xnor U9963 (N_9963,N_7482,N_7058);
and U9964 (N_9964,N_6307,N_7253);
nand U9965 (N_9965,N_6570,N_6295);
or U9966 (N_9966,N_7186,N_7476);
xnor U9967 (N_9967,N_6092,N_6083);
nand U9968 (N_9968,N_6805,N_7092);
nor U9969 (N_9969,N_7578,N_7240);
and U9970 (N_9970,N_6677,N_7443);
nand U9971 (N_9971,N_6692,N_6140);
or U9972 (N_9972,N_6402,N_6246);
nor U9973 (N_9973,N_7659,N_7364);
nor U9974 (N_9974,N_7393,N_6595);
and U9975 (N_9975,N_6966,N_7879);
or U9976 (N_9976,N_7373,N_6665);
or U9977 (N_9977,N_7490,N_7528);
or U9978 (N_9978,N_6833,N_6634);
nor U9979 (N_9979,N_7493,N_7480);
and U9980 (N_9980,N_6221,N_6381);
nor U9981 (N_9981,N_6894,N_7435);
nand U9982 (N_9982,N_6797,N_7471);
or U9983 (N_9983,N_6339,N_6883);
nor U9984 (N_9984,N_6056,N_7196);
nor U9985 (N_9985,N_6024,N_7688);
or U9986 (N_9986,N_6932,N_7886);
and U9987 (N_9987,N_7639,N_7833);
nor U9988 (N_9988,N_7749,N_7634);
nand U9989 (N_9989,N_6280,N_7294);
or U9990 (N_9990,N_7482,N_7408);
or U9991 (N_9991,N_7303,N_7882);
or U9992 (N_9992,N_7367,N_6713);
nand U9993 (N_9993,N_6342,N_7686);
and U9994 (N_9994,N_6721,N_6374);
and U9995 (N_9995,N_7891,N_7875);
xnor U9996 (N_9996,N_6329,N_7369);
nor U9997 (N_9997,N_7548,N_6115);
nor U9998 (N_9998,N_6093,N_6442);
nand U9999 (N_9999,N_7902,N_7932);
nor U10000 (N_10000,N_8305,N_9712);
or U10001 (N_10001,N_8211,N_8647);
nand U10002 (N_10002,N_8417,N_9402);
nor U10003 (N_10003,N_9890,N_8412);
or U10004 (N_10004,N_9656,N_8878);
and U10005 (N_10005,N_9071,N_8166);
xor U10006 (N_10006,N_9796,N_8349);
nor U10007 (N_10007,N_9439,N_8142);
nor U10008 (N_10008,N_8099,N_9948);
or U10009 (N_10009,N_8549,N_9468);
nor U10010 (N_10010,N_8177,N_8885);
nand U10011 (N_10011,N_8192,N_8038);
xnor U10012 (N_10012,N_8152,N_8804);
xor U10013 (N_10013,N_8010,N_8794);
nor U10014 (N_10014,N_9204,N_9535);
and U10015 (N_10015,N_9283,N_8614);
and U10016 (N_10016,N_9777,N_8932);
or U10017 (N_10017,N_8429,N_9149);
xor U10018 (N_10018,N_9376,N_8447);
nor U10019 (N_10019,N_8572,N_9597);
xor U10020 (N_10020,N_8227,N_8013);
nor U10021 (N_10021,N_9703,N_8726);
or U10022 (N_10022,N_8992,N_8999);
nor U10023 (N_10023,N_8656,N_9737);
or U10024 (N_10024,N_9857,N_8964);
nor U10025 (N_10025,N_9619,N_8242);
nand U10026 (N_10026,N_9643,N_9031);
nor U10027 (N_10027,N_9942,N_8293);
nor U10028 (N_10028,N_9486,N_8256);
xor U10029 (N_10029,N_8959,N_9772);
xnor U10030 (N_10030,N_8302,N_8213);
and U10031 (N_10031,N_8460,N_9269);
nand U10032 (N_10032,N_9244,N_8048);
and U10033 (N_10033,N_8503,N_9934);
or U10034 (N_10034,N_8587,N_9202);
nand U10035 (N_10035,N_8043,N_9629);
nor U10036 (N_10036,N_9655,N_9590);
xnor U10037 (N_10037,N_8845,N_8011);
and U10038 (N_10038,N_9545,N_9697);
and U10039 (N_10039,N_8171,N_9055);
and U10040 (N_10040,N_8299,N_9841);
nor U10041 (N_10041,N_8626,N_9518);
or U10042 (N_10042,N_9346,N_8107);
or U10043 (N_10043,N_8100,N_9318);
nor U10044 (N_10044,N_9524,N_8632);
or U10045 (N_10045,N_8955,N_9785);
nor U10046 (N_10046,N_8122,N_9152);
xor U10047 (N_10047,N_9749,N_8078);
xor U10048 (N_10048,N_9199,N_8251);
and U10049 (N_10049,N_9039,N_8223);
xnor U10050 (N_10050,N_8623,N_9561);
nor U10051 (N_10051,N_9853,N_8901);
nand U10052 (N_10052,N_8390,N_9583);
nor U10053 (N_10053,N_9610,N_8609);
or U10054 (N_10054,N_8655,N_8432);
or U10055 (N_10055,N_9370,N_8454);
nor U10056 (N_10056,N_8336,N_9862);
xnor U10057 (N_10057,N_9715,N_8364);
xnor U10058 (N_10058,N_8457,N_8443);
and U10059 (N_10059,N_9121,N_8513);
and U10060 (N_10060,N_9194,N_9906);
and U10061 (N_10061,N_8442,N_9374);
xor U10062 (N_10062,N_9157,N_9787);
nand U10063 (N_10063,N_9773,N_9297);
nand U10064 (N_10064,N_9153,N_9998);
xor U10065 (N_10065,N_9236,N_8874);
xor U10066 (N_10066,N_9064,N_8176);
xnor U10067 (N_10067,N_8820,N_8556);
xor U10068 (N_10068,N_8406,N_9633);
or U10069 (N_10069,N_8009,N_8965);
or U10070 (N_10070,N_9483,N_8568);
nor U10071 (N_10071,N_9427,N_8659);
or U10072 (N_10072,N_9249,N_8024);
and U10073 (N_10073,N_8034,N_9366);
and U10074 (N_10074,N_8883,N_9081);
nor U10075 (N_10075,N_9650,N_8800);
and U10076 (N_10076,N_9696,N_8924);
or U10077 (N_10077,N_9133,N_8830);
nand U10078 (N_10078,N_8561,N_8813);
xor U10079 (N_10079,N_9181,N_8335);
or U10080 (N_10080,N_8271,N_9587);
nor U10081 (N_10081,N_8080,N_8927);
xor U10082 (N_10082,N_9635,N_9222);
nand U10083 (N_10083,N_9471,N_8421);
xor U10084 (N_10084,N_8347,N_9276);
nor U10085 (N_10085,N_9909,N_9437);
nand U10086 (N_10086,N_9451,N_9176);
nor U10087 (N_10087,N_8154,N_8770);
and U10088 (N_10088,N_8319,N_9676);
and U10089 (N_10089,N_9810,N_8797);
nand U10090 (N_10090,N_8052,N_9821);
nand U10091 (N_10091,N_9245,N_8359);
or U10092 (N_10092,N_8836,N_8323);
nand U10093 (N_10093,N_9294,N_9111);
and U10094 (N_10094,N_9602,N_8473);
nor U10095 (N_10095,N_8670,N_8534);
nand U10096 (N_10096,N_8189,N_9992);
or U10097 (N_10097,N_9018,N_8546);
or U10098 (N_10098,N_8768,N_8680);
nand U10099 (N_10099,N_8907,N_9229);
or U10100 (N_10100,N_8428,N_8725);
or U10101 (N_10101,N_8554,N_9735);
xnor U10102 (N_10102,N_8968,N_8764);
nand U10103 (N_10103,N_8182,N_8969);
or U10104 (N_10104,N_9322,N_9621);
nor U10105 (N_10105,N_9497,N_9617);
or U10106 (N_10106,N_9137,N_9690);
or U10107 (N_10107,N_8005,N_8237);
nand U10108 (N_10108,N_8779,N_9344);
and U10109 (N_10109,N_8222,N_8277);
nand U10110 (N_10110,N_8066,N_9500);
and U10111 (N_10111,N_8583,N_8749);
nand U10112 (N_10112,N_8346,N_8669);
nand U10113 (N_10113,N_8200,N_8648);
or U10114 (N_10114,N_9469,N_8115);
xor U10115 (N_10115,N_8516,N_9160);
xor U10116 (N_10116,N_9396,N_8449);
xor U10117 (N_10117,N_8098,N_9799);
xnor U10118 (N_10118,N_9037,N_8668);
xnor U10119 (N_10119,N_8003,N_9104);
or U10120 (N_10120,N_8709,N_9743);
and U10121 (N_10121,N_9642,N_9755);
and U10122 (N_10122,N_9571,N_8821);
and U10123 (N_10123,N_9110,N_9963);
nand U10124 (N_10124,N_8151,N_8582);
and U10125 (N_10125,N_8119,N_8146);
xor U10126 (N_10126,N_9254,N_8689);
nor U10127 (N_10127,N_8717,N_9896);
and U10128 (N_10128,N_9720,N_9534);
and U10129 (N_10129,N_8723,N_8475);
or U10130 (N_10130,N_9593,N_8812);
and U10131 (N_10131,N_9769,N_9701);
nand U10132 (N_10132,N_9581,N_8488);
nand U10133 (N_10133,N_9837,N_9774);
or U10134 (N_10134,N_9714,N_8399);
nor U10135 (N_10135,N_8016,N_8258);
and U10136 (N_10136,N_9393,N_8472);
and U10137 (N_10137,N_9813,N_9052);
xnor U10138 (N_10138,N_8594,N_9231);
nand U10139 (N_10139,N_8934,N_9739);
or U10140 (N_10140,N_8133,N_9567);
or U10141 (N_10141,N_8480,N_9733);
xor U10142 (N_10142,N_9060,N_8795);
xnor U10143 (N_10143,N_9513,N_8906);
or U10144 (N_10144,N_8398,N_9214);
and U10145 (N_10145,N_8361,N_9291);
xnor U10146 (N_10146,N_9702,N_9098);
nor U10147 (N_10147,N_9219,N_8089);
nand U10148 (N_10148,N_9442,N_8411);
or U10149 (N_10149,N_9713,N_9887);
xnor U10150 (N_10150,N_8756,N_9203);
xnor U10151 (N_10151,N_9107,N_8807);
or U10152 (N_10152,N_8339,N_8840);
and U10153 (N_10153,N_8490,N_8774);
and U10154 (N_10154,N_9109,N_8922);
nor U10155 (N_10155,N_8022,N_8719);
nor U10156 (N_10156,N_8953,N_8937);
nor U10157 (N_10157,N_8851,N_9260);
or U10158 (N_10158,N_9449,N_8837);
or U10159 (N_10159,N_9757,N_8909);
xnor U10160 (N_10160,N_8504,N_9191);
and U10161 (N_10161,N_8716,N_9049);
or U10162 (N_10162,N_8117,N_8198);
nand U10163 (N_10163,N_8091,N_8073);
xor U10164 (N_10164,N_8778,N_8983);
and U10165 (N_10165,N_8848,N_9316);
or U10166 (N_10166,N_8598,N_8752);
xor U10167 (N_10167,N_9788,N_9336);
xnor U10168 (N_10168,N_8703,N_8573);
nand U10169 (N_10169,N_8026,N_9870);
and U10170 (N_10170,N_9674,N_8645);
xnor U10171 (N_10171,N_8380,N_9280);
xor U10172 (N_10172,N_8287,N_8739);
xor U10173 (N_10173,N_9122,N_9016);
nor U10174 (N_10174,N_8585,N_9424);
nor U10175 (N_10175,N_8579,N_9683);
and U10176 (N_10176,N_9675,N_9649);
or U10177 (N_10177,N_9577,N_9613);
or U10178 (N_10178,N_9846,N_9335);
and U10179 (N_10179,N_8341,N_8039);
or U10180 (N_10180,N_8613,N_8118);
and U10181 (N_10181,N_9419,N_8537);
xor U10182 (N_10182,N_9200,N_9716);
xor U10183 (N_10183,N_9038,N_9072);
or U10184 (N_10184,N_8963,N_9169);
nor U10185 (N_10185,N_9786,N_9937);
and U10186 (N_10186,N_9802,N_9227);
and U10187 (N_10187,N_9759,N_9827);
nor U10188 (N_10188,N_9069,N_9804);
nor U10189 (N_10189,N_8315,N_9671);
xor U10190 (N_10190,N_8199,N_9453);
nand U10191 (N_10191,N_8831,N_9412);
xor U10192 (N_10192,N_9916,N_9271);
xor U10193 (N_10193,N_8126,N_8741);
xor U10194 (N_10194,N_9085,N_8371);
nand U10195 (N_10195,N_9845,N_8744);
or U10196 (N_10196,N_8178,N_9794);
or U10197 (N_10197,N_8025,N_8289);
and U10198 (N_10198,N_8044,N_8345);
or U10199 (N_10199,N_9398,N_8675);
or U10200 (N_10200,N_8788,N_9797);
xor U10201 (N_10201,N_9900,N_8765);
nand U10202 (N_10202,N_8030,N_8738);
or U10203 (N_10203,N_9170,N_9615);
nand U10204 (N_10204,N_8793,N_9340);
xor U10205 (N_10205,N_8275,N_8140);
and U10206 (N_10206,N_8174,N_9985);
xor U10207 (N_10207,N_9901,N_9997);
xor U10208 (N_10208,N_8300,N_9144);
nor U10209 (N_10209,N_9084,N_9263);
and U10210 (N_10210,N_8654,N_8902);
and U10211 (N_10211,N_8230,N_8958);
and U10212 (N_10212,N_9397,N_9850);
or U10213 (N_10213,N_9476,N_8858);
and U10214 (N_10214,N_9988,N_8402);
and U10215 (N_10215,N_8015,N_8479);
and U10216 (N_10216,N_9126,N_9407);
nand U10217 (N_10217,N_9261,N_9265);
xor U10218 (N_10218,N_8577,N_8520);
nand U10219 (N_10219,N_9529,N_9717);
and U10220 (N_10220,N_9413,N_9557);
xor U10221 (N_10221,N_8621,N_8850);
xor U10222 (N_10222,N_9552,N_8388);
xor U10223 (N_10223,N_8045,N_8826);
xnor U10224 (N_10224,N_9303,N_8041);
xor U10225 (N_10225,N_8747,N_9333);
and U10226 (N_10226,N_8083,N_9032);
and U10227 (N_10227,N_8849,N_8167);
nor U10228 (N_10228,N_8913,N_9512);
xnor U10229 (N_10229,N_9582,N_8129);
and U10230 (N_10230,N_8781,N_9048);
and U10231 (N_10231,N_9741,N_8046);
and U10232 (N_10232,N_8921,N_8735);
or U10233 (N_10233,N_8569,N_9530);
or U10234 (N_10234,N_8827,N_8674);
or U10235 (N_10235,N_8375,N_8097);
or U10236 (N_10236,N_8019,N_9080);
or U10237 (N_10237,N_9975,N_9403);
or U10238 (N_10238,N_9299,N_9030);
nand U10239 (N_10239,N_8630,N_9738);
xnor U10240 (N_10240,N_9317,N_9806);
and U10241 (N_10241,N_9921,N_8545);
xnor U10242 (N_10242,N_8303,N_8441);
and U10243 (N_10243,N_8558,N_9467);
and U10244 (N_10244,N_8617,N_8606);
xor U10245 (N_10245,N_8920,N_8929);
xor U10246 (N_10246,N_9851,N_8517);
nor U10247 (N_10247,N_9815,N_9764);
and U10248 (N_10248,N_8508,N_9885);
nand U10249 (N_10249,N_9286,N_8027);
or U10250 (N_10250,N_9595,N_8282);
xor U10251 (N_10251,N_9950,N_9563);
nor U10252 (N_10252,N_8387,N_9522);
or U10253 (N_10253,N_9953,N_9814);
nand U10254 (N_10254,N_9805,N_8642);
nand U10255 (N_10255,N_8350,N_8591);
nor U10256 (N_10256,N_9225,N_9996);
xnor U10257 (N_10257,N_9196,N_8497);
xor U10258 (N_10258,N_9478,N_9097);
nand U10259 (N_10259,N_8772,N_9586);
nand U10260 (N_10260,N_8981,N_9003);
or U10261 (N_10261,N_9417,N_9936);
and U10262 (N_10262,N_9112,N_8215);
xnor U10263 (N_10263,N_9051,N_8759);
nand U10264 (N_10264,N_8210,N_9094);
nor U10265 (N_10265,N_9010,N_9295);
nor U10266 (N_10266,N_8148,N_9803);
or U10267 (N_10267,N_8419,N_9977);
nand U10268 (N_10268,N_8001,N_8751);
and U10269 (N_10269,N_9433,N_9927);
nor U10270 (N_10270,N_9059,N_8529);
nor U10271 (N_10271,N_8757,N_8366);
or U10272 (N_10272,N_8578,N_8970);
nor U10273 (N_10273,N_9005,N_9627);
nand U10274 (N_10274,N_8020,N_8787);
nor U10275 (N_10275,N_8047,N_8708);
xnor U10276 (N_10276,N_8574,N_9751);
xnor U10277 (N_10277,N_9239,N_8718);
and U10278 (N_10278,N_8935,N_9960);
or U10279 (N_10279,N_8822,N_8195);
xnor U10280 (N_10280,N_8157,N_8159);
or U10281 (N_10281,N_9224,N_8553);
and U10282 (N_10282,N_9371,N_8530);
or U10283 (N_10283,N_8264,N_8903);
or U10284 (N_10284,N_9641,N_8590);
xor U10285 (N_10285,N_9025,N_8061);
and U10286 (N_10286,N_9677,N_8312);
and U10287 (N_10287,N_9892,N_9723);
or U10288 (N_10288,N_9142,N_8514);
and U10289 (N_10289,N_8183,N_9447);
or U10290 (N_10290,N_8743,N_8095);
and U10291 (N_10291,N_8301,N_8252);
nor U10292 (N_10292,N_9315,N_9982);
nor U10293 (N_10293,N_9466,N_8263);
nand U10294 (N_10294,N_9822,N_8522);
xnor U10295 (N_10295,N_9753,N_8990);
xnor U10296 (N_10296,N_8662,N_9425);
or U10297 (N_10297,N_9117,N_8538);
xnor U10298 (N_10298,N_8801,N_9767);
or U10299 (N_10299,N_9289,N_9812);
nand U10300 (N_10300,N_8945,N_9281);
nand U10301 (N_10301,N_9480,N_9611);
and U10302 (N_10302,N_9957,N_8123);
nor U10303 (N_10303,N_8681,N_8007);
and U10304 (N_10304,N_8491,N_9429);
or U10305 (N_10305,N_9275,N_8313);
nand U10306 (N_10306,N_8403,N_9377);
xnor U10307 (N_10307,N_9658,N_8678);
xnor U10308 (N_10308,N_9124,N_8511);
nor U10309 (N_10309,N_8435,N_9994);
or U10310 (N_10310,N_8108,N_9130);
nand U10311 (N_10311,N_8754,N_8898);
xor U10312 (N_10312,N_9448,N_9680);
nand U10313 (N_10313,N_9257,N_9848);
nand U10314 (N_10314,N_9247,N_8724);
or U10315 (N_10315,N_8438,N_9362);
and U10316 (N_10316,N_9365,N_9243);
nand U10317 (N_10317,N_8104,N_8110);
nor U10318 (N_10318,N_8567,N_8467);
xnor U10319 (N_10319,N_9493,N_9017);
xnor U10320 (N_10320,N_9798,N_8592);
nor U10321 (N_10321,N_9542,N_8374);
nor U10322 (N_10322,N_9015,N_9668);
and U10323 (N_10323,N_9589,N_8695);
or U10324 (N_10324,N_8424,N_9095);
or U10325 (N_10325,N_9919,N_8141);
nand U10326 (N_10326,N_8410,N_8641);
nand U10327 (N_10327,N_8649,N_8112);
or U10328 (N_10328,N_9186,N_8803);
or U10329 (N_10329,N_9849,N_8239);
and U10330 (N_10330,N_9073,N_8607);
and U10331 (N_10331,N_9758,N_9113);
and U10332 (N_10332,N_9746,N_9925);
or U10333 (N_10333,N_9301,N_8204);
nor U10334 (N_10334,N_8862,N_8377);
xor U10335 (N_10335,N_9657,N_8124);
or U10336 (N_10336,N_8487,N_8181);
or U10337 (N_10337,N_8518,N_9965);
or U10338 (N_10338,N_8939,N_9601);
xnor U10339 (N_10339,N_8062,N_8891);
xnor U10340 (N_10340,N_8519,N_9915);
xor U10341 (N_10341,N_9351,N_9521);
nor U10342 (N_10342,N_8633,N_9310);
xor U10343 (N_10343,N_9387,N_9938);
nor U10344 (N_10344,N_9820,N_8688);
xor U10345 (N_10345,N_8832,N_8805);
nor U10346 (N_10346,N_9431,N_9562);
and U10347 (N_10347,N_9604,N_8967);
or U10348 (N_10348,N_8249,N_9838);
xnor U10349 (N_10349,N_8042,N_9995);
xnor U10350 (N_10350,N_8385,N_8175);
nand U10351 (N_10351,N_8186,N_8557);
nor U10352 (N_10352,N_9359,N_9883);
and U10353 (N_10353,N_9300,N_8393);
nor U10354 (N_10354,N_9308,N_9272);
or U10355 (N_10355,N_9775,N_8564);
or U10356 (N_10356,N_8236,N_8815);
nor U10357 (N_10357,N_9125,N_8401);
and U10358 (N_10358,N_9893,N_8462);
or U10359 (N_10359,N_9205,N_8995);
xnor U10360 (N_10360,N_8373,N_9736);
nor U10361 (N_10361,N_9970,N_8610);
xor U10362 (N_10362,N_9600,N_9544);
and U10363 (N_10363,N_9436,N_8855);
and U10364 (N_10364,N_8431,N_9665);
xor U10365 (N_10365,N_8079,N_9311);
or U10366 (N_10366,N_9296,N_9592);
nand U10367 (N_10367,N_9539,N_8414);
nor U10368 (N_10368,N_8288,N_9666);
nor U10369 (N_10369,N_9819,N_9831);
xnor U10370 (N_10370,N_9498,N_8881);
nand U10371 (N_10371,N_8773,N_9750);
nor U10372 (N_10372,N_8279,N_8000);
xnor U10373 (N_10373,N_8331,N_8687);
nor U10374 (N_10374,N_8321,N_8396);
nand U10375 (N_10375,N_8919,N_8165);
nand U10376 (N_10376,N_8704,N_9083);
or U10377 (N_10377,N_8527,N_8444);
and U10378 (N_10378,N_8698,N_8814);
xor U10379 (N_10379,N_9201,N_9728);
and U10380 (N_10380,N_8470,N_9704);
xor U10381 (N_10381,N_9584,N_9783);
or U10382 (N_10382,N_8535,N_9711);
and U10383 (N_10383,N_9150,N_9268);
xnor U10384 (N_10384,N_9001,N_9390);
nand U10385 (N_10385,N_9895,N_9978);
nand U10386 (N_10386,N_8789,N_9019);
and U10387 (N_10387,N_8624,N_8074);
nand U10388 (N_10388,N_8326,N_8382);
xnor U10389 (N_10389,N_9686,N_9780);
or U10390 (N_10390,N_8317,N_9879);
xor U10391 (N_10391,N_9458,N_8143);
nor U10392 (N_10392,N_9914,N_8111);
nand U10393 (N_10393,N_8087,N_9006);
nand U10394 (N_10394,N_8232,N_8458);
or U10395 (N_10395,N_9155,N_9389);
or U10396 (N_10396,N_8600,N_9826);
nand U10397 (N_10397,N_9158,N_9246);
and U10398 (N_10398,N_8481,N_8705);
nor U10399 (N_10399,N_9935,N_8163);
or U10400 (N_10400,N_9099,N_9103);
and U10401 (N_10401,N_9989,N_8523);
nor U10402 (N_10402,N_8168,N_8076);
or U10403 (N_10403,N_8340,N_8267);
and U10404 (N_10404,N_9947,N_8077);
xnor U10405 (N_10405,N_9605,N_8265);
xor U10406 (N_10406,N_8653,N_8309);
nand U10407 (N_10407,N_8865,N_9218);
nand U10408 (N_10408,N_8559,N_8397);
xnor U10409 (N_10409,N_8116,N_9543);
and U10410 (N_10410,N_9752,N_8203);
nand U10411 (N_10411,N_9430,N_8188);
xnor U10412 (N_10412,N_8482,N_8890);
xor U10413 (N_10413,N_9718,N_9760);
xor U10414 (N_10414,N_8502,N_8816);
nor U10415 (N_10415,N_8464,N_8531);
or U10416 (N_10416,N_8551,N_8905);
xnor U10417 (N_10417,N_9208,N_8158);
and U10418 (N_10418,N_9279,N_9569);
nand U10419 (N_10419,N_8780,N_9050);
xnor U10420 (N_10420,N_9404,N_8147);
and U10421 (N_10421,N_9648,N_8325);
or U10422 (N_10422,N_8253,N_8418);
or U10423 (N_10423,N_8231,N_8950);
or U10424 (N_10424,N_8144,N_9022);
nor U10425 (N_10425,N_8835,N_8775);
xor U10426 (N_10426,N_9609,N_9386);
and U10427 (N_10427,N_9740,N_9782);
and U10428 (N_10428,N_9210,N_8248);
nor U10429 (N_10429,N_8547,N_8067);
nor U10430 (N_10430,N_8295,N_9159);
nand U10431 (N_10431,N_8852,N_9585);
xnor U10432 (N_10432,N_8539,N_9598);
or U10433 (N_10433,N_9646,N_9987);
or U10434 (N_10434,N_9999,N_8246);
or U10435 (N_10435,N_8785,N_8071);
and U10436 (N_10436,N_8220,N_8075);
or U10437 (N_10437,N_9504,N_8348);
nor U10438 (N_10438,N_8971,N_8873);
and U10439 (N_10439,N_8028,N_9452);
nand U10440 (N_10440,N_9105,N_8944);
xor U10441 (N_10441,N_8525,N_9614);
or U10442 (N_10442,N_9045,N_9742);
nor U10443 (N_10443,N_8229,N_9756);
nor U10444 (N_10444,N_9670,N_8450);
nor U10445 (N_10445,N_8996,N_9762);
xnor U10446 (N_10446,N_9363,N_9488);
nand U10447 (N_10447,N_8818,N_8928);
nand U10448 (N_10448,N_8580,N_9020);
and U10449 (N_10449,N_8702,N_9913);
and U10450 (N_10450,N_8576,N_9630);
xor U10451 (N_10451,N_9139,N_9911);
and U10452 (N_10452,N_9014,N_9177);
nand U10453 (N_10453,N_9548,N_8221);
and U10454 (N_10454,N_8180,N_8002);
or U10455 (N_10455,N_9042,N_9454);
nand U10456 (N_10456,N_9538,N_8892);
nor U10457 (N_10457,N_9008,N_8201);
xnor U10458 (N_10458,N_9259,N_9379);
xor U10459 (N_10459,N_9930,N_8652);
and U10460 (N_10460,N_9933,N_8243);
and U10461 (N_10461,N_9355,N_9328);
nor U10462 (N_10462,N_9537,N_9361);
and U10463 (N_10463,N_9178,N_9274);
and U10464 (N_10464,N_8439,N_9375);
nand U10465 (N_10465,N_8162,N_9596);
or U10466 (N_10466,N_9881,N_8871);
or U10467 (N_10467,N_9345,N_8542);
xor U10468 (N_10468,N_8059,N_9213);
xnor U10469 (N_10469,N_9145,N_9863);
nand U10470 (N_10470,N_8064,N_9108);
and U10471 (N_10471,N_9624,N_8226);
xor U10472 (N_10472,N_9556,N_9520);
xor U10473 (N_10473,N_8761,N_9817);
nor U10474 (N_10474,N_9106,N_8494);
nand U10475 (N_10475,N_9441,N_9146);
nand U10476 (N_10476,N_9705,N_8185);
xor U10477 (N_10477,N_9331,N_8120);
or U10478 (N_10478,N_9876,N_9868);
or U10479 (N_10479,N_9215,N_8218);
nor U10480 (N_10480,N_9367,N_8870);
nor U10481 (N_10481,N_9664,N_9415);
xor U10482 (N_10482,N_8381,N_8661);
nor U10483 (N_10483,N_9706,N_8395);
xor U10484 (N_10484,N_9087,N_9574);
nor U10485 (N_10485,N_9047,N_8135);
or U10486 (N_10486,N_9645,N_9551);
nor U10487 (N_10487,N_8828,N_8427);
and U10488 (N_10488,N_9843,N_9682);
or U10489 (N_10489,N_9727,N_8139);
xor U10490 (N_10490,N_9482,N_8506);
or U10491 (N_10491,N_9182,N_9477);
or U10492 (N_10492,N_9349,N_9284);
nand U10493 (N_10493,N_9304,N_9902);
or U10494 (N_10494,N_9491,N_8868);
nor U10495 (N_10495,N_9855,N_8543);
or U10496 (N_10496,N_8817,N_9102);
or U10497 (N_10497,N_9140,N_8261);
or U10498 (N_10498,N_8351,N_9654);
xnor U10499 (N_10499,N_9662,N_9894);
nor U10500 (N_10500,N_8172,N_9864);
and U10501 (N_10501,N_9632,N_8477);
nor U10502 (N_10502,N_8560,N_8466);
nand U10503 (N_10503,N_8550,N_9258);
and U10504 (N_10504,N_8671,N_8276);
nand U10505 (N_10505,N_8650,N_9348);
xor U10506 (N_10506,N_8006,N_9233);
xor U10507 (N_10507,N_9305,N_9460);
and U10508 (N_10508,N_9667,N_8362);
nand U10509 (N_10509,N_9079,N_8235);
nor U10510 (N_10510,N_9066,N_8008);
xor U10511 (N_10511,N_8233,N_8501);
xnor U10512 (N_10512,N_8899,N_9681);
nor U10513 (N_10513,N_8984,N_8665);
nand U10514 (N_10514,N_8054,N_8127);
nand U10515 (N_10515,N_8468,N_9165);
nand U10516 (N_10516,N_8285,N_9332);
or U10517 (N_10517,N_9253,N_9958);
nand U10518 (N_10518,N_9410,N_9496);
and U10519 (N_10519,N_9041,N_9114);
nand U10520 (N_10520,N_8191,N_9639);
or U10521 (N_10521,N_9119,N_9399);
xor U10522 (N_10522,N_9588,N_9264);
xnor U10523 (N_10523,N_9388,N_8733);
nor U10524 (N_10524,N_8948,N_9195);
and U10525 (N_10525,N_9226,N_8699);
nor U10526 (N_10526,N_9575,N_9086);
and U10527 (N_10527,N_8337,N_8031);
and U10528 (N_10528,N_8440,N_9063);
or U10529 (N_10529,N_9197,N_8416);
nand U10530 (N_10530,N_8365,N_8876);
nor U10531 (N_10531,N_8982,N_9494);
nor U10532 (N_10532,N_8692,N_9473);
and U10533 (N_10533,N_8618,N_8925);
nand U10534 (N_10534,N_9499,N_9235);
xnor U10535 (N_10535,N_9354,N_9678);
nor U10536 (N_10536,N_8274,N_8933);
nor U10537 (N_10537,N_8409,N_9972);
xor U10538 (N_10538,N_8776,N_8798);
and U10539 (N_10539,N_9212,N_8114);
nand U10540 (N_10540,N_8352,N_9628);
xor U10541 (N_10541,N_8400,N_9012);
nand U10542 (N_10542,N_8672,N_8334);
nand U10543 (N_10543,N_8021,N_8386);
and U10544 (N_10544,N_8853,N_9409);
or U10545 (N_10545,N_9240,N_8755);
nand U10546 (N_10546,N_8985,N_9731);
or U10547 (N_10547,N_9078,N_9465);
or U10548 (N_10548,N_8307,N_8096);
nand U10549 (N_10549,N_9091,N_9237);
and U10550 (N_10550,N_8161,N_9382);
or U10551 (N_10551,N_8035,N_9256);
xor U10552 (N_10552,N_9185,N_8247);
xnor U10553 (N_10553,N_9961,N_8993);
nor U10554 (N_10554,N_8225,N_8344);
xnor U10555 (N_10555,N_9070,N_8316);
xnor U10556 (N_10556,N_9011,N_8997);
and U10557 (N_10557,N_8732,N_9000);
nand U10558 (N_10558,N_9606,N_8555);
nor U10559 (N_10559,N_9183,N_9461);
nand U10560 (N_10560,N_9156,N_9341);
nand U10561 (N_10561,N_8420,N_9368);
nand U10562 (N_10562,N_8639,N_9871);
or U10563 (N_10563,N_9339,N_8053);
or U10564 (N_10564,N_9984,N_8838);
nor U10565 (N_10565,N_9120,N_8570);
or U10566 (N_10566,N_9710,N_9991);
nor U10567 (N_10567,N_9854,N_9959);
xnor U10568 (N_10568,N_9096,N_9401);
nand U10569 (N_10569,N_8994,N_9287);
xor U10570 (N_10570,N_8338,N_8908);
nor U10571 (N_10571,N_9492,N_9192);
nor U10572 (N_10572,N_8036,N_9298);
xnor U10573 (N_10573,N_8640,N_9004);
nor U10574 (N_10574,N_8452,N_9986);
or U10575 (N_10575,N_9456,N_8631);
or U10576 (N_10576,N_9035,N_8512);
and U10577 (N_10577,N_8392,N_9459);
nand U10578 (N_10578,N_9912,N_8268);
nor U10579 (N_10579,N_8912,N_9860);
nand U10580 (N_10580,N_8946,N_9818);
nand U10581 (N_10581,N_8763,N_8938);
nor U10582 (N_10582,N_8823,N_9053);
nand U10583 (N_10583,N_9330,N_9129);
or U10584 (N_10584,N_8012,N_8029);
xnor U10585 (N_10585,N_8563,N_9168);
xnor U10586 (N_10586,N_8691,N_8040);
xnor U10587 (N_10587,N_8426,N_9904);
or U10588 (N_10588,N_9056,N_9100);
nor U10589 (N_10589,N_9910,N_9941);
xnor U10590 (N_10590,N_8138,N_9745);
or U10591 (N_10591,N_8956,N_9891);
xnor U10592 (N_10592,N_9463,N_9013);
nor U10593 (N_10593,N_8360,N_9669);
nand U10594 (N_10594,N_8679,N_8446);
nor U10595 (N_10595,N_8685,N_8977);
or U10596 (N_10596,N_9148,N_8734);
xor U10597 (N_10597,N_8297,N_9694);
nor U10598 (N_10598,N_8354,N_8290);
xor U10599 (N_10599,N_8391,N_9517);
or U10600 (N_10600,N_9372,N_9940);
xor U10601 (N_10601,N_9768,N_9184);
xnor U10602 (N_10602,N_8923,N_9781);
or U10603 (N_10603,N_8343,N_8461);
nand U10604 (N_10604,N_9625,N_9880);
and U10605 (N_10605,N_8260,N_8566);
xor U10606 (N_10606,N_8496,N_8164);
nand U10607 (N_10607,N_8859,N_9443);
and U10608 (N_10608,N_8690,N_9440);
xor U10609 (N_10609,N_8526,N_9151);
nand U10610 (N_10610,N_8842,N_8824);
xnor U10611 (N_10611,N_9693,N_9293);
or U10612 (N_10612,N_9220,N_8790);
nand U10613 (N_10613,N_9692,N_8485);
nand U10614 (N_10614,N_9190,N_9928);
nand U10615 (N_10615,N_8667,N_9572);
nor U10616 (N_10616,N_9926,N_9479);
and U10617 (N_10617,N_9721,N_9554);
nand U10618 (N_10618,N_9278,N_9509);
xor U10619 (N_10619,N_8136,N_9623);
xor U10620 (N_10620,N_9503,N_9874);
xnor U10621 (N_10621,N_8004,N_8294);
and U10622 (N_10622,N_8658,N_8942);
or U10623 (N_10623,N_9290,N_8284);
nand U10624 (N_10624,N_9288,N_8978);
and U10625 (N_10625,N_9882,N_8379);
and U10626 (N_10626,N_9949,N_9180);
or U10627 (N_10627,N_8806,N_8729);
nand U10628 (N_10628,N_8941,N_8489);
and U10629 (N_10629,N_9067,N_8507);
nand U10630 (N_10630,N_8125,N_9068);
xnor U10631 (N_10631,N_9307,N_8562);
nand U10632 (N_10632,N_8094,N_9699);
xor U10633 (N_10633,N_8254,N_8930);
and U10634 (N_10634,N_8949,N_9426);
and U10635 (N_10635,N_8082,N_8808);
nand U10636 (N_10636,N_8711,N_9968);
nand U10637 (N_10637,N_9147,N_9266);
nand U10638 (N_10638,N_8771,N_8864);
nand U10639 (N_10639,N_9839,N_9406);
or U10640 (N_10640,N_9434,N_9899);
xor U10641 (N_10641,N_8792,N_9023);
nor U10642 (N_10642,N_8216,N_9411);
xnor U10643 (N_10643,N_8536,N_8961);
nor U10644 (N_10644,N_9285,N_8611);
nor U10645 (N_10645,N_9724,N_8088);
and U10646 (N_10646,N_8620,N_8532);
or U10647 (N_10647,N_8612,N_9432);
nand U10648 (N_10648,N_9836,N_9391);
or U10649 (N_10649,N_9709,N_9962);
xor U10650 (N_10650,N_8072,N_8666);
xnor U10651 (N_10651,N_9455,N_8451);
nand U10652 (N_10652,N_9270,N_8799);
nand U10653 (N_10653,N_9983,N_9776);
nor U10654 (N_10654,N_8697,N_8783);
nand U10655 (N_10655,N_8484,N_9135);
nor U10656 (N_10656,N_9966,N_9092);
xnor U10657 (N_10657,N_8483,N_8280);
nand U10658 (N_10658,N_9867,N_8311);
nor U10659 (N_10659,N_8184,N_9878);
and U10660 (N_10660,N_9062,N_9034);
nand U10661 (N_10661,N_9976,N_9093);
xnor U10662 (N_10662,N_9725,N_9075);
or U10663 (N_10663,N_8713,N_8193);
nand U10664 (N_10664,N_9421,N_8809);
and U10665 (N_10665,N_9043,N_9834);
nor U10666 (N_10666,N_8540,N_9967);
nand U10667 (N_10667,N_8701,N_9905);
or U10668 (N_10668,N_9793,N_9580);
and U10669 (N_10669,N_9599,N_8308);
xnor U10670 (N_10670,N_9685,N_8132);
xor U10671 (N_10671,N_8742,N_9400);
xnor U10672 (N_10672,N_8367,N_8767);
xor U10673 (N_10673,N_8476,N_8664);
nand U10674 (N_10674,N_8109,N_9134);
xnor U10675 (N_10675,N_8604,N_9550);
and U10676 (N_10676,N_8296,N_8453);
nor U10677 (N_10677,N_8037,N_9323);
nand U10678 (N_10678,N_9964,N_8106);
xnor U10679 (N_10679,N_8422,N_8465);
nand U10680 (N_10680,N_8057,N_8050);
nand U10681 (N_10681,N_8936,N_9188);
nor U10682 (N_10682,N_8829,N_9637);
or U10683 (N_10683,N_9326,N_8190);
xnor U10684 (N_10684,N_8292,N_9353);
xor U10685 (N_10685,N_9128,N_9033);
or U10686 (N_10686,N_8269,N_9536);
xor U10687 (N_10687,N_9687,N_9856);
nand U10688 (N_10688,N_9282,N_9262);
nor U10689 (N_10689,N_9695,N_8746);
nor U10690 (N_10690,N_8207,N_9620);
and U10691 (N_10691,N_8895,N_8715);
and U10692 (N_10692,N_9352,N_8926);
nand U10693 (N_10693,N_8459,N_9811);
and U10694 (N_10694,N_8628,N_9872);
or U10695 (N_10695,N_9040,N_8962);
or U10696 (N_10696,N_8205,N_8304);
or U10697 (N_10697,N_8291,N_9221);
xnor U10698 (N_10698,N_9519,N_9241);
nor U10699 (N_10699,N_9061,N_8081);
nor U10700 (N_10700,N_9700,N_9765);
nor U10701 (N_10701,N_9136,N_8219);
xnor U10702 (N_10702,N_8255,N_9252);
and U10703 (N_10703,N_9771,N_8068);
and U10704 (N_10704,N_8306,N_8405);
and U10705 (N_10705,N_8722,N_9462);
nor U10706 (N_10706,N_8844,N_9444);
xor U10707 (N_10707,N_9313,N_8437);
nor U10708 (N_10708,N_8358,N_8056);
xor U10709 (N_10709,N_8436,N_8974);
xor U10710 (N_10710,N_9044,N_8646);
and U10711 (N_10711,N_9384,N_9779);
nor U10712 (N_10712,N_8430,N_8445);
xnor U10713 (N_10713,N_8493,N_8515);
or U10714 (N_10714,N_8149,N_9578);
or U10715 (N_10715,N_8196,N_8627);
xor U10716 (N_10716,N_8879,N_9659);
xor U10717 (N_10717,N_9175,N_9510);
and U10718 (N_10718,N_9560,N_8637);
xnor U10719 (N_10719,N_9791,N_8694);
or U10720 (N_10720,N_8069,N_8603);
and U10721 (N_10721,N_9546,N_8372);
or U10722 (N_10722,N_8018,N_9242);
xnor U10723 (N_10723,N_9945,N_9334);
and U10724 (N_10724,N_9644,N_9358);
nor U10725 (N_10725,N_9719,N_9356);
or U10726 (N_10726,N_9943,N_8987);
xor U10727 (N_10727,N_9474,N_8330);
xnor U10728 (N_10728,N_8954,N_8943);
or U10729 (N_10729,N_8867,N_8212);
or U10730 (N_10730,N_8368,N_8931);
xnor U10731 (N_10731,N_9594,N_9501);
xor U10732 (N_10732,N_9689,N_8134);
or U10733 (N_10733,N_9918,N_9360);
nand U10734 (N_10734,N_9167,N_8677);
and U10735 (N_10735,N_8363,N_9487);
nor U10736 (N_10736,N_9445,N_9844);
and U10737 (N_10737,N_8745,N_8651);
and U10738 (N_10738,N_8615,N_8857);
or U10739 (N_10739,N_9127,N_9636);
or U10740 (N_10740,N_8769,N_9923);
nor U10741 (N_10741,N_8415,N_8032);
xnor U10742 (N_10742,N_9903,N_9971);
or U10743 (N_10743,N_8169,N_9932);
and U10744 (N_10744,N_8055,N_9405);
xnor U10745 (N_10745,N_9485,N_9591);
and U10746 (N_10746,N_8278,N_8998);
xor U10747 (N_10747,N_9907,N_9884);
and U10748 (N_10748,N_9508,N_8113);
xnor U10749 (N_10749,N_9869,N_9684);
or U10750 (N_10750,N_8262,N_9920);
nand U10751 (N_10751,N_9292,N_9211);
nor U10752 (N_10752,N_9579,N_8802);
or U10753 (N_10753,N_8533,N_9990);
nand U10754 (N_10754,N_9277,N_8173);
nor U10755 (N_10755,N_9707,N_9832);
nor U10756 (N_10756,N_9842,N_9321);
and U10757 (N_10757,N_9954,N_9823);
nor U10758 (N_10758,N_9533,N_9054);
nand U10759 (N_10759,N_8214,N_9074);
and U10760 (N_10760,N_9217,N_8407);
xnor U10761 (N_10761,N_8318,N_9663);
nand U10762 (N_10762,N_9250,N_8988);
nand U10763 (N_10763,N_9414,N_9490);
nor U10764 (N_10764,N_9526,N_9481);
and U10765 (N_10765,N_9570,N_9889);
xor U10766 (N_10766,N_9174,N_9255);
nand U10767 (N_10767,N_9897,N_8811);
and U10768 (N_10768,N_9638,N_8888);
nor U10769 (N_10769,N_9395,N_9754);
and U10770 (N_10770,N_8972,N_9438);
and U10771 (N_10771,N_8619,N_8332);
nand U10772 (N_10772,N_8721,N_9828);
nand U10773 (N_10773,N_8896,N_9408);
and U10774 (N_10774,N_8084,N_8866);
nor U10775 (N_10775,N_9024,N_8228);
xnor U10776 (N_10776,N_9830,N_8796);
or U10777 (N_10777,N_8413,N_9541);
nand U10778 (N_10778,N_9939,N_8825);
nand U10779 (N_10779,N_9981,N_9314);
xnor U10780 (N_10780,N_8153,N_9929);
and U10781 (N_10781,N_8856,N_8731);
nand U10782 (N_10782,N_9428,N_8408);
xnor U10783 (N_10783,N_9337,N_9329);
or U10784 (N_10784,N_9320,N_8707);
xor U10785 (N_10785,N_9232,N_8571);
nand U10786 (N_10786,N_8914,N_9946);
xor U10787 (N_10787,N_9306,N_8884);
and U10788 (N_10788,N_8875,N_9847);
or U10789 (N_10789,N_8486,N_8748);
or U10790 (N_10790,N_9640,N_8986);
nand U10791 (N_10791,N_8565,N_8102);
and U10792 (N_10792,N_8712,N_9908);
nand U10793 (N_10793,N_8777,N_8989);
nand U10794 (N_10794,N_9917,N_9730);
nor U10795 (N_10795,N_8601,N_9888);
nand U10796 (N_10796,N_9525,N_8544);
and U10797 (N_10797,N_9824,N_8455);
xor U10798 (N_10798,N_8588,N_9143);
xnor U10799 (N_10799,N_9324,N_9209);
nor U10800 (N_10800,N_9866,N_8105);
nor U10801 (N_10801,N_9422,N_8714);
nand U10802 (N_10802,N_9154,N_9618);
and U10803 (N_10803,N_9065,N_9082);
or U10804 (N_10804,N_9002,N_8049);
nand U10805 (N_10805,N_8595,N_8217);
and U10806 (N_10806,N_8495,N_8209);
or U10807 (N_10807,N_9172,N_9944);
or U10808 (N_10808,N_8663,N_9801);
or U10809 (N_10809,N_9951,N_9343);
or U10810 (N_10810,N_9364,N_8456);
nand U10811 (N_10811,N_8498,N_8854);
and U10812 (N_10812,N_9688,N_8657);
xor U10813 (N_10813,N_9325,N_8322);
or U10814 (N_10814,N_9875,N_8638);
or U10815 (N_10815,N_9672,N_8593);
nor U10816 (N_10816,N_9319,N_8684);
xor U10817 (N_10817,N_8194,N_8833);
or U10818 (N_10818,N_8910,N_8310);
or U10819 (N_10819,N_9446,N_8070);
nand U10820 (N_10820,N_8017,N_8499);
nor U10821 (N_10821,N_8737,N_8728);
nor U10822 (N_10822,N_9852,N_9612);
xnor U10823 (N_10823,N_9327,N_9956);
or U10824 (N_10824,N_8384,N_8179);
nor U10825 (N_10825,N_9974,N_8103);
xnor U10826 (N_10826,N_9123,N_9540);
nand U10827 (N_10827,N_8947,N_8644);
or U10828 (N_10828,N_9251,N_9568);
xnor U10829 (N_10829,N_9189,N_8602);
nand U10830 (N_10830,N_9835,N_9164);
nand U10831 (N_10831,N_8170,N_8492);
nor U10832 (N_10832,N_9565,N_8584);
xor U10833 (N_10833,N_9416,N_9784);
nor U10834 (N_10834,N_8145,N_8940);
or U10835 (N_10835,N_9865,N_9732);
and U10836 (N_10836,N_8766,N_8589);
or U10837 (N_10837,N_9077,N_8272);
and U10838 (N_10838,N_8758,N_9532);
and U10839 (N_10839,N_8206,N_8634);
and U10840 (N_10840,N_8469,N_9631);
or U10841 (N_10841,N_8324,N_9514);
or U10842 (N_10842,N_8991,N_8882);
nand U10843 (N_10843,N_8886,N_9969);
nor U10844 (N_10844,N_8887,N_9734);
and U10845 (N_10845,N_9116,N_8524);
or U10846 (N_10846,N_9026,N_8900);
and U10847 (N_10847,N_9979,N_9161);
or U10848 (N_10848,N_9385,N_8425);
or U10849 (N_10849,N_9502,N_9187);
and U10850 (N_10850,N_8880,N_8861);
nor U10851 (N_10851,N_8033,N_9859);
or U10852 (N_10852,N_8342,N_9131);
nand U10853 (N_10853,N_8383,N_9179);
xnor U10854 (N_10854,N_8463,N_9495);
or U10855 (N_10855,N_8753,N_8051);
nand U10856 (N_10856,N_9511,N_9223);
or U10857 (N_10857,N_9993,N_8841);
and U10858 (N_10858,N_8509,N_8389);
xor U10859 (N_10859,N_8682,N_8376);
and U10860 (N_10860,N_9861,N_9338);
nor U10861 (N_10861,N_8283,N_9369);
nor U10862 (N_10862,N_8625,N_8710);
or U10863 (N_10863,N_9886,N_9816);
and U10864 (N_10864,N_8581,N_9980);
nor U10865 (N_10865,N_9549,N_9506);
and U10866 (N_10866,N_8329,N_9559);
nand U10867 (N_10867,N_8023,N_8298);
or U10868 (N_10868,N_9634,N_8683);
nor U10869 (N_10869,N_8250,N_9877);
xnor U10870 (N_10870,N_9516,N_8086);
and U10871 (N_10871,N_8819,N_9373);
nand U10872 (N_10872,N_9778,N_9118);
and U10873 (N_10873,N_8060,N_8150);
nand U10874 (N_10874,N_8357,N_9248);
or U10875 (N_10875,N_9651,N_9952);
nand U10876 (N_10876,N_9475,N_9029);
or U10877 (N_10877,N_8314,N_9898);
xnor U10878 (N_10878,N_8863,N_8877);
and U10879 (N_10879,N_8394,N_9115);
nand U10880 (N_10880,N_9564,N_9829);
xor U10881 (N_10881,N_9342,N_8636);
or U10882 (N_10882,N_8635,N_8605);
or U10883 (N_10883,N_9840,N_9507);
nand U10884 (N_10884,N_9484,N_9955);
xnor U10885 (N_10885,N_9558,N_9566);
and U10886 (N_10886,N_9380,N_9141);
or U10887 (N_10887,N_8693,N_8090);
xnor U10888 (N_10888,N_8960,N_9347);
xnor U10889 (N_10889,N_9673,N_8197);
nor U10890 (N_10890,N_9171,N_8599);
xor U10891 (N_10891,N_8234,N_8706);
and U10892 (N_10892,N_9607,N_9708);
nor U10893 (N_10893,N_9470,N_8575);
and U10894 (N_10894,N_8320,N_8063);
nand U10895 (N_10895,N_9858,N_8951);
and U10896 (N_10896,N_9789,N_8782);
nand U10897 (N_10897,N_8736,N_9547);
xnor U10898 (N_10898,N_8762,N_9228);
xnor U10899 (N_10899,N_8894,N_8156);
xnor U10900 (N_10900,N_8730,N_9198);
or U10901 (N_10901,N_8676,N_9457);
or U10902 (N_10902,N_9726,N_8889);
and U10903 (N_10903,N_8966,N_8092);
xnor U10904 (N_10904,N_8975,N_8085);
or U10905 (N_10905,N_8916,N_9273);
or U10906 (N_10906,N_9729,N_8952);
nor U10907 (N_10907,N_9101,N_9698);
nand U10908 (N_10908,N_9435,N_8448);
nor U10909 (N_10909,N_9378,N_8869);
nor U10910 (N_10910,N_9661,N_8327);
and U10911 (N_10911,N_8750,N_8596);
or U10912 (N_10912,N_9057,N_8784);
or U10913 (N_10913,N_8471,N_9652);
or U10914 (N_10914,N_9088,N_9973);
and U10915 (N_10915,N_9653,N_8328);
nor U10916 (N_10916,N_9450,N_8058);
nand U10917 (N_10917,N_8155,N_8353);
or U10918 (N_10918,N_9691,N_8433);
nand U10919 (N_10919,N_8643,N_8286);
xor U10920 (N_10920,N_8541,N_9392);
or U10921 (N_10921,N_9931,N_9163);
or U10922 (N_10922,N_8130,N_8131);
nor U10923 (N_10923,N_8093,N_9350);
or U10924 (N_10924,N_9770,N_9312);
and U10925 (N_10925,N_8500,N_8521);
nand U10926 (N_10926,N_9036,N_9747);
and U10927 (N_10927,N_9238,N_8245);
nand U10928 (N_10928,N_9722,N_8872);
nand U10929 (N_10929,N_8834,N_8510);
or U10930 (N_10930,N_9555,N_8240);
and U10931 (N_10931,N_9027,N_9309);
or U10932 (N_10932,N_9523,N_8740);
xor U10933 (N_10933,N_8370,N_9922);
nand U10934 (N_10934,N_9576,N_9267);
xor U10935 (N_10935,N_9660,N_9162);
nor U10936 (N_10936,N_9464,N_9748);
nand U10937 (N_10937,N_8957,N_8897);
nor U10938 (N_10938,N_8720,N_8244);
xnor U10939 (N_10939,N_8700,N_9795);
or U10940 (N_10940,N_9528,N_9381);
and U10941 (N_10941,N_9383,N_9790);
nand U10942 (N_10942,N_8281,N_9230);
xor U10943 (N_10943,N_8238,N_8423);
nand U10944 (N_10944,N_8616,N_9766);
nand U10945 (N_10945,N_8356,N_8846);
or U10946 (N_10946,N_9166,N_8727);
or U10947 (N_10947,N_9009,N_8369);
and U10948 (N_10948,N_8786,N_9924);
or U10949 (N_10949,N_8202,N_8548);
nand U10950 (N_10950,N_9302,N_8187);
xnor U10951 (N_10951,N_9809,N_9206);
nand U10952 (N_10952,N_8976,N_9394);
or U10953 (N_10953,N_8597,N_8673);
and U10954 (N_10954,N_8860,N_9527);
nand U10955 (N_10955,N_8014,N_8622);
and U10956 (N_10956,N_8552,N_8528);
xor U10957 (N_10957,N_8760,N_9058);
and U10958 (N_10958,N_9089,N_9216);
or U10959 (N_10959,N_8660,N_8979);
or U10960 (N_10960,N_9021,N_9825);
xnor U10961 (N_10961,N_9472,N_9808);
xnor U10962 (N_10962,N_8843,N_9357);
nor U10963 (N_10963,N_9647,N_8608);
nor U10964 (N_10964,N_8810,N_9515);
and U10965 (N_10965,N_8241,N_8065);
xnor U10966 (N_10966,N_9800,N_8586);
nand U10967 (N_10967,N_8160,N_9792);
and U10968 (N_10968,N_8355,N_9873);
nand U10969 (N_10969,N_9761,N_9622);
xor U10970 (N_10970,N_9679,N_8101);
nand U10971 (N_10971,N_9626,N_8378);
and U10972 (N_10972,N_9420,N_8973);
nor U10973 (N_10973,N_8257,N_9616);
and U10974 (N_10974,N_9418,N_8911);
and U10975 (N_10975,N_9531,N_8259);
and U10976 (N_10976,N_8918,N_8333);
and U10977 (N_10977,N_8208,N_9608);
and U10978 (N_10978,N_9763,N_8478);
xnor U10979 (N_10979,N_9046,N_8696);
or U10980 (N_10980,N_9234,N_9833);
and U10981 (N_10981,N_9173,N_9193);
or U10982 (N_10982,N_8904,N_8270);
nor U10983 (N_10983,N_9132,N_9505);
or U10984 (N_10984,N_8266,N_8224);
or U10985 (N_10985,N_8137,N_9603);
and U10986 (N_10986,N_8980,N_9138);
and U10987 (N_10987,N_9090,N_9553);
nand U10988 (N_10988,N_8917,N_8839);
xor U10989 (N_10989,N_9007,N_9028);
nor U10990 (N_10990,N_9076,N_9207);
nand U10991 (N_10991,N_9573,N_9807);
and U10992 (N_10992,N_9744,N_8505);
and U10993 (N_10993,N_8128,N_8686);
nor U10994 (N_10994,N_8629,N_8434);
and U10995 (N_10995,N_8474,N_8847);
nand U10996 (N_10996,N_9489,N_8121);
or U10997 (N_10997,N_8915,N_8273);
nand U10998 (N_10998,N_8791,N_8404);
nand U10999 (N_10999,N_8893,N_9423);
nor U11000 (N_11000,N_9849,N_9024);
or U11001 (N_11001,N_9396,N_9381);
and U11002 (N_11002,N_8051,N_8714);
and U11003 (N_11003,N_9095,N_8835);
nor U11004 (N_11004,N_9626,N_9527);
xor U11005 (N_11005,N_9515,N_9056);
nand U11006 (N_11006,N_8873,N_9269);
and U11007 (N_11007,N_9716,N_9044);
nand U11008 (N_11008,N_9703,N_8981);
nand U11009 (N_11009,N_8973,N_8859);
and U11010 (N_11010,N_9667,N_9578);
xor U11011 (N_11011,N_8978,N_9909);
nand U11012 (N_11012,N_9947,N_9831);
nor U11013 (N_11013,N_9126,N_8156);
or U11014 (N_11014,N_9981,N_9273);
or U11015 (N_11015,N_8167,N_8484);
nand U11016 (N_11016,N_9592,N_8527);
and U11017 (N_11017,N_9877,N_9210);
and U11018 (N_11018,N_9325,N_9682);
xor U11019 (N_11019,N_8673,N_8359);
and U11020 (N_11020,N_8810,N_9900);
nor U11021 (N_11021,N_8085,N_8484);
nor U11022 (N_11022,N_8497,N_8116);
or U11023 (N_11023,N_9390,N_8036);
nand U11024 (N_11024,N_8332,N_9108);
xor U11025 (N_11025,N_8571,N_8812);
nand U11026 (N_11026,N_9643,N_9482);
and U11027 (N_11027,N_8904,N_8661);
or U11028 (N_11028,N_8288,N_8628);
or U11029 (N_11029,N_9005,N_9217);
nand U11030 (N_11030,N_8127,N_9345);
xor U11031 (N_11031,N_8653,N_9417);
xnor U11032 (N_11032,N_8739,N_8517);
or U11033 (N_11033,N_9118,N_8998);
nand U11034 (N_11034,N_8093,N_9322);
and U11035 (N_11035,N_9760,N_9924);
xor U11036 (N_11036,N_8211,N_8899);
or U11037 (N_11037,N_8023,N_9161);
nor U11038 (N_11038,N_9963,N_8118);
nand U11039 (N_11039,N_8700,N_9188);
nor U11040 (N_11040,N_9255,N_9126);
or U11041 (N_11041,N_8664,N_9965);
xor U11042 (N_11042,N_9627,N_8480);
or U11043 (N_11043,N_9213,N_9949);
or U11044 (N_11044,N_8386,N_8834);
xnor U11045 (N_11045,N_8852,N_9742);
nand U11046 (N_11046,N_9351,N_9219);
and U11047 (N_11047,N_8544,N_9025);
or U11048 (N_11048,N_8922,N_9981);
nor U11049 (N_11049,N_9517,N_8609);
nand U11050 (N_11050,N_8778,N_8023);
nor U11051 (N_11051,N_9310,N_9888);
nand U11052 (N_11052,N_9585,N_8426);
or U11053 (N_11053,N_9990,N_8145);
nand U11054 (N_11054,N_9192,N_9474);
nor U11055 (N_11055,N_9812,N_8810);
nand U11056 (N_11056,N_8180,N_9198);
and U11057 (N_11057,N_9530,N_8242);
or U11058 (N_11058,N_8865,N_9478);
xor U11059 (N_11059,N_8810,N_9623);
xor U11060 (N_11060,N_9831,N_8167);
xor U11061 (N_11061,N_8075,N_8032);
nand U11062 (N_11062,N_8718,N_9867);
nor U11063 (N_11063,N_9777,N_9804);
and U11064 (N_11064,N_9213,N_8975);
nor U11065 (N_11065,N_8832,N_9148);
and U11066 (N_11066,N_8317,N_8027);
xnor U11067 (N_11067,N_9240,N_8044);
or U11068 (N_11068,N_8717,N_9940);
nand U11069 (N_11069,N_9743,N_8694);
and U11070 (N_11070,N_9518,N_8957);
nor U11071 (N_11071,N_9216,N_9949);
and U11072 (N_11072,N_8136,N_9173);
nand U11073 (N_11073,N_8013,N_8957);
nand U11074 (N_11074,N_8558,N_9091);
xnor U11075 (N_11075,N_8616,N_8745);
nand U11076 (N_11076,N_9404,N_9130);
and U11077 (N_11077,N_8925,N_8824);
and U11078 (N_11078,N_9413,N_8041);
and U11079 (N_11079,N_9662,N_8947);
xor U11080 (N_11080,N_9923,N_9166);
and U11081 (N_11081,N_8365,N_8429);
nand U11082 (N_11082,N_8673,N_9591);
nand U11083 (N_11083,N_8709,N_8410);
nor U11084 (N_11084,N_9369,N_8066);
xor U11085 (N_11085,N_9819,N_8461);
or U11086 (N_11086,N_8354,N_9020);
nand U11087 (N_11087,N_9489,N_8039);
xor U11088 (N_11088,N_9776,N_9892);
and U11089 (N_11089,N_9317,N_9002);
nand U11090 (N_11090,N_8988,N_9928);
xnor U11091 (N_11091,N_8936,N_9313);
nor U11092 (N_11092,N_8271,N_9574);
nand U11093 (N_11093,N_8022,N_9795);
nor U11094 (N_11094,N_8204,N_8254);
and U11095 (N_11095,N_8901,N_8284);
and U11096 (N_11096,N_9214,N_9302);
nand U11097 (N_11097,N_8842,N_8366);
and U11098 (N_11098,N_9046,N_9464);
nor U11099 (N_11099,N_8229,N_8789);
nand U11100 (N_11100,N_9870,N_9649);
nand U11101 (N_11101,N_9578,N_8400);
and U11102 (N_11102,N_9693,N_8223);
nand U11103 (N_11103,N_8273,N_9165);
nand U11104 (N_11104,N_9445,N_9363);
xor U11105 (N_11105,N_9858,N_9845);
xor U11106 (N_11106,N_8189,N_8209);
or U11107 (N_11107,N_8331,N_9370);
and U11108 (N_11108,N_9436,N_9644);
xor U11109 (N_11109,N_9344,N_9025);
and U11110 (N_11110,N_8517,N_9051);
or U11111 (N_11111,N_8173,N_8849);
xnor U11112 (N_11112,N_8485,N_9435);
nor U11113 (N_11113,N_8986,N_9843);
nand U11114 (N_11114,N_9639,N_9869);
nor U11115 (N_11115,N_8305,N_8038);
xnor U11116 (N_11116,N_8407,N_9092);
or U11117 (N_11117,N_9658,N_8906);
nand U11118 (N_11118,N_9485,N_8333);
or U11119 (N_11119,N_9466,N_8514);
xnor U11120 (N_11120,N_9236,N_8733);
xnor U11121 (N_11121,N_9256,N_8797);
and U11122 (N_11122,N_8443,N_8045);
nor U11123 (N_11123,N_9888,N_8788);
and U11124 (N_11124,N_8564,N_9311);
or U11125 (N_11125,N_9028,N_8734);
nand U11126 (N_11126,N_9931,N_8751);
nand U11127 (N_11127,N_9303,N_9728);
or U11128 (N_11128,N_9361,N_8649);
and U11129 (N_11129,N_9098,N_8737);
nand U11130 (N_11130,N_8913,N_9475);
nand U11131 (N_11131,N_8642,N_9000);
or U11132 (N_11132,N_9129,N_8790);
nor U11133 (N_11133,N_9325,N_9156);
nand U11134 (N_11134,N_8068,N_8613);
nand U11135 (N_11135,N_8272,N_8057);
nand U11136 (N_11136,N_9820,N_9059);
or U11137 (N_11137,N_8850,N_8120);
nand U11138 (N_11138,N_9153,N_8366);
or U11139 (N_11139,N_8282,N_8987);
and U11140 (N_11140,N_9353,N_8935);
nand U11141 (N_11141,N_8362,N_9080);
nand U11142 (N_11142,N_8546,N_8895);
or U11143 (N_11143,N_8086,N_8466);
and U11144 (N_11144,N_9713,N_8123);
xor U11145 (N_11145,N_9270,N_9717);
nor U11146 (N_11146,N_8327,N_8886);
nor U11147 (N_11147,N_9839,N_8286);
nand U11148 (N_11148,N_8307,N_9423);
xor U11149 (N_11149,N_9962,N_8008);
nor U11150 (N_11150,N_9336,N_8757);
and U11151 (N_11151,N_9198,N_9938);
xor U11152 (N_11152,N_9909,N_9724);
or U11153 (N_11153,N_9332,N_9900);
nand U11154 (N_11154,N_8927,N_9028);
or U11155 (N_11155,N_8887,N_9490);
or U11156 (N_11156,N_9696,N_8339);
nand U11157 (N_11157,N_9019,N_9926);
nor U11158 (N_11158,N_8658,N_9488);
xnor U11159 (N_11159,N_9617,N_9949);
nand U11160 (N_11160,N_8044,N_9169);
or U11161 (N_11161,N_8044,N_9713);
and U11162 (N_11162,N_9189,N_9606);
xnor U11163 (N_11163,N_9151,N_9621);
nand U11164 (N_11164,N_8532,N_9879);
nand U11165 (N_11165,N_9670,N_8165);
xor U11166 (N_11166,N_9445,N_9939);
nor U11167 (N_11167,N_8129,N_9647);
xnor U11168 (N_11168,N_8138,N_8963);
and U11169 (N_11169,N_8190,N_9724);
nand U11170 (N_11170,N_8204,N_8896);
nand U11171 (N_11171,N_8731,N_8651);
or U11172 (N_11172,N_8001,N_8004);
and U11173 (N_11173,N_8417,N_9581);
nor U11174 (N_11174,N_8964,N_8816);
or U11175 (N_11175,N_8879,N_9360);
and U11176 (N_11176,N_8899,N_8309);
and U11177 (N_11177,N_8289,N_8452);
nor U11178 (N_11178,N_9981,N_9833);
and U11179 (N_11179,N_8880,N_8688);
xnor U11180 (N_11180,N_8137,N_8225);
nor U11181 (N_11181,N_9949,N_9053);
nand U11182 (N_11182,N_8948,N_9096);
nor U11183 (N_11183,N_8165,N_9300);
nand U11184 (N_11184,N_9184,N_8203);
and U11185 (N_11185,N_9054,N_8981);
and U11186 (N_11186,N_8583,N_8352);
nand U11187 (N_11187,N_8311,N_8051);
and U11188 (N_11188,N_8131,N_9062);
or U11189 (N_11189,N_8698,N_8529);
xor U11190 (N_11190,N_9492,N_8481);
and U11191 (N_11191,N_8761,N_9788);
nand U11192 (N_11192,N_8540,N_9337);
xnor U11193 (N_11193,N_9714,N_8123);
nand U11194 (N_11194,N_9813,N_9597);
and U11195 (N_11195,N_8759,N_9810);
and U11196 (N_11196,N_8884,N_9367);
and U11197 (N_11197,N_9334,N_8168);
and U11198 (N_11198,N_9498,N_8386);
nor U11199 (N_11199,N_9378,N_9404);
or U11200 (N_11200,N_8174,N_9642);
and U11201 (N_11201,N_9108,N_8329);
nand U11202 (N_11202,N_8940,N_8615);
or U11203 (N_11203,N_9674,N_8584);
nor U11204 (N_11204,N_9988,N_8929);
and U11205 (N_11205,N_8558,N_9101);
or U11206 (N_11206,N_9440,N_9975);
nor U11207 (N_11207,N_9181,N_8958);
xor U11208 (N_11208,N_8381,N_8713);
and U11209 (N_11209,N_9530,N_9301);
nand U11210 (N_11210,N_9579,N_8937);
nor U11211 (N_11211,N_9449,N_8593);
nor U11212 (N_11212,N_9509,N_8477);
and U11213 (N_11213,N_9756,N_9372);
nand U11214 (N_11214,N_8074,N_8572);
or U11215 (N_11215,N_8306,N_9132);
and U11216 (N_11216,N_8556,N_9957);
nand U11217 (N_11217,N_8390,N_9621);
nor U11218 (N_11218,N_9750,N_9322);
or U11219 (N_11219,N_9687,N_9909);
nand U11220 (N_11220,N_8091,N_8455);
and U11221 (N_11221,N_8291,N_8749);
xnor U11222 (N_11222,N_9112,N_8769);
and U11223 (N_11223,N_9314,N_9885);
nor U11224 (N_11224,N_9666,N_8263);
xor U11225 (N_11225,N_9799,N_9284);
nor U11226 (N_11226,N_8982,N_9283);
xnor U11227 (N_11227,N_8283,N_9363);
and U11228 (N_11228,N_9742,N_9105);
nor U11229 (N_11229,N_9926,N_9160);
nand U11230 (N_11230,N_8568,N_9668);
nor U11231 (N_11231,N_8871,N_9907);
or U11232 (N_11232,N_8073,N_8144);
and U11233 (N_11233,N_8491,N_8019);
or U11234 (N_11234,N_8099,N_8781);
and U11235 (N_11235,N_8249,N_9752);
and U11236 (N_11236,N_9535,N_8725);
nand U11237 (N_11237,N_9614,N_8021);
nand U11238 (N_11238,N_9944,N_8888);
or U11239 (N_11239,N_8535,N_9920);
xor U11240 (N_11240,N_9976,N_8499);
nand U11241 (N_11241,N_8086,N_8352);
or U11242 (N_11242,N_9949,N_8950);
xor U11243 (N_11243,N_9241,N_9678);
nor U11244 (N_11244,N_9925,N_9945);
nand U11245 (N_11245,N_9158,N_8489);
nand U11246 (N_11246,N_9387,N_9960);
nor U11247 (N_11247,N_9200,N_9491);
nand U11248 (N_11248,N_8024,N_8786);
nor U11249 (N_11249,N_9772,N_8523);
nand U11250 (N_11250,N_8767,N_8665);
nand U11251 (N_11251,N_9728,N_9501);
and U11252 (N_11252,N_9958,N_9154);
xor U11253 (N_11253,N_9246,N_9517);
nor U11254 (N_11254,N_8222,N_9271);
nor U11255 (N_11255,N_8901,N_8113);
nand U11256 (N_11256,N_8362,N_9071);
or U11257 (N_11257,N_9814,N_9272);
nor U11258 (N_11258,N_8683,N_9612);
or U11259 (N_11259,N_8158,N_8708);
and U11260 (N_11260,N_9850,N_9919);
and U11261 (N_11261,N_8681,N_9189);
xnor U11262 (N_11262,N_9631,N_8325);
nand U11263 (N_11263,N_8812,N_8012);
or U11264 (N_11264,N_8276,N_9205);
xor U11265 (N_11265,N_9733,N_9882);
and U11266 (N_11266,N_8390,N_9931);
and U11267 (N_11267,N_9671,N_8768);
xor U11268 (N_11268,N_9883,N_8908);
xor U11269 (N_11269,N_8477,N_8613);
nand U11270 (N_11270,N_8100,N_9337);
or U11271 (N_11271,N_9818,N_8876);
or U11272 (N_11272,N_8297,N_8969);
or U11273 (N_11273,N_9046,N_8756);
nand U11274 (N_11274,N_8454,N_9692);
and U11275 (N_11275,N_9106,N_8141);
nor U11276 (N_11276,N_8811,N_8496);
nand U11277 (N_11277,N_9144,N_8869);
nor U11278 (N_11278,N_9369,N_8935);
xnor U11279 (N_11279,N_8774,N_8053);
and U11280 (N_11280,N_9908,N_9283);
and U11281 (N_11281,N_8750,N_9327);
xor U11282 (N_11282,N_9902,N_9789);
nor U11283 (N_11283,N_8003,N_8018);
nor U11284 (N_11284,N_9671,N_8349);
nor U11285 (N_11285,N_8235,N_9941);
or U11286 (N_11286,N_9467,N_8605);
or U11287 (N_11287,N_8855,N_8448);
xnor U11288 (N_11288,N_8885,N_9401);
and U11289 (N_11289,N_9516,N_8095);
or U11290 (N_11290,N_8070,N_8159);
or U11291 (N_11291,N_9901,N_9415);
xnor U11292 (N_11292,N_9593,N_8735);
xnor U11293 (N_11293,N_8329,N_9610);
and U11294 (N_11294,N_9052,N_9620);
or U11295 (N_11295,N_8628,N_8040);
xnor U11296 (N_11296,N_8962,N_9606);
and U11297 (N_11297,N_8297,N_9477);
and U11298 (N_11298,N_9740,N_9868);
and U11299 (N_11299,N_9899,N_9626);
nand U11300 (N_11300,N_9876,N_9598);
or U11301 (N_11301,N_8684,N_9214);
nor U11302 (N_11302,N_9878,N_9253);
nand U11303 (N_11303,N_8552,N_9228);
nor U11304 (N_11304,N_9599,N_9636);
or U11305 (N_11305,N_8959,N_8811);
nand U11306 (N_11306,N_8668,N_8802);
and U11307 (N_11307,N_8896,N_9007);
xnor U11308 (N_11308,N_8749,N_8117);
or U11309 (N_11309,N_8810,N_9306);
xnor U11310 (N_11310,N_9848,N_9461);
xnor U11311 (N_11311,N_9252,N_9125);
and U11312 (N_11312,N_8138,N_8236);
and U11313 (N_11313,N_9443,N_9941);
nor U11314 (N_11314,N_8594,N_9196);
xnor U11315 (N_11315,N_9044,N_9067);
xnor U11316 (N_11316,N_9702,N_9203);
or U11317 (N_11317,N_9881,N_9591);
and U11318 (N_11318,N_9592,N_8293);
nor U11319 (N_11319,N_8677,N_9729);
or U11320 (N_11320,N_8132,N_9311);
nand U11321 (N_11321,N_8321,N_8206);
and U11322 (N_11322,N_9390,N_9724);
and U11323 (N_11323,N_8112,N_8524);
nor U11324 (N_11324,N_9794,N_9985);
or U11325 (N_11325,N_9957,N_9754);
and U11326 (N_11326,N_8440,N_9569);
and U11327 (N_11327,N_8419,N_9660);
or U11328 (N_11328,N_9976,N_8881);
or U11329 (N_11329,N_8082,N_9260);
and U11330 (N_11330,N_8911,N_9705);
nand U11331 (N_11331,N_9974,N_8801);
and U11332 (N_11332,N_8093,N_9096);
xnor U11333 (N_11333,N_9383,N_9009);
nor U11334 (N_11334,N_9934,N_8401);
nor U11335 (N_11335,N_8795,N_8789);
and U11336 (N_11336,N_9833,N_9605);
xnor U11337 (N_11337,N_9166,N_8306);
nor U11338 (N_11338,N_9988,N_9462);
and U11339 (N_11339,N_8013,N_9057);
nand U11340 (N_11340,N_8057,N_8503);
xor U11341 (N_11341,N_9828,N_9811);
xor U11342 (N_11342,N_8347,N_8558);
or U11343 (N_11343,N_9021,N_8799);
or U11344 (N_11344,N_9753,N_8437);
and U11345 (N_11345,N_9716,N_8610);
nand U11346 (N_11346,N_8510,N_9367);
xnor U11347 (N_11347,N_9179,N_8273);
nand U11348 (N_11348,N_8891,N_9006);
nand U11349 (N_11349,N_8228,N_8823);
xor U11350 (N_11350,N_8712,N_9766);
xor U11351 (N_11351,N_8411,N_8291);
and U11352 (N_11352,N_9064,N_9204);
and U11353 (N_11353,N_8592,N_8436);
xnor U11354 (N_11354,N_8055,N_8528);
nand U11355 (N_11355,N_8549,N_8792);
or U11356 (N_11356,N_9234,N_8446);
nand U11357 (N_11357,N_9481,N_9802);
or U11358 (N_11358,N_8745,N_9864);
nor U11359 (N_11359,N_8062,N_9119);
xnor U11360 (N_11360,N_9914,N_9828);
nand U11361 (N_11361,N_8013,N_8952);
or U11362 (N_11362,N_9358,N_9803);
nor U11363 (N_11363,N_8867,N_8454);
nand U11364 (N_11364,N_9528,N_9076);
xnor U11365 (N_11365,N_8363,N_8396);
nand U11366 (N_11366,N_9142,N_9082);
and U11367 (N_11367,N_9987,N_9847);
nand U11368 (N_11368,N_8411,N_9313);
or U11369 (N_11369,N_9616,N_9819);
nor U11370 (N_11370,N_8336,N_8614);
nor U11371 (N_11371,N_9974,N_8457);
nand U11372 (N_11372,N_8146,N_8333);
nor U11373 (N_11373,N_8010,N_9810);
and U11374 (N_11374,N_8332,N_8815);
and U11375 (N_11375,N_9433,N_8243);
or U11376 (N_11376,N_8634,N_9534);
nor U11377 (N_11377,N_8874,N_8306);
nand U11378 (N_11378,N_8326,N_8733);
xor U11379 (N_11379,N_9021,N_8218);
xnor U11380 (N_11380,N_9018,N_8423);
and U11381 (N_11381,N_9070,N_9742);
nor U11382 (N_11382,N_9736,N_8254);
and U11383 (N_11383,N_8861,N_8708);
nor U11384 (N_11384,N_9468,N_8422);
or U11385 (N_11385,N_9321,N_9989);
nor U11386 (N_11386,N_8422,N_8195);
nand U11387 (N_11387,N_9727,N_8634);
nor U11388 (N_11388,N_8508,N_9909);
and U11389 (N_11389,N_8145,N_8104);
and U11390 (N_11390,N_8218,N_8243);
and U11391 (N_11391,N_9734,N_9231);
or U11392 (N_11392,N_9473,N_8630);
nor U11393 (N_11393,N_9483,N_9538);
nor U11394 (N_11394,N_9225,N_8394);
nor U11395 (N_11395,N_9947,N_9280);
or U11396 (N_11396,N_9472,N_8340);
and U11397 (N_11397,N_8079,N_8693);
xnor U11398 (N_11398,N_9485,N_9729);
nor U11399 (N_11399,N_9255,N_8769);
nand U11400 (N_11400,N_8413,N_8392);
or U11401 (N_11401,N_8642,N_9694);
or U11402 (N_11402,N_9079,N_9730);
or U11403 (N_11403,N_9697,N_8133);
and U11404 (N_11404,N_9435,N_9242);
and U11405 (N_11405,N_9639,N_9173);
xnor U11406 (N_11406,N_9257,N_9965);
nand U11407 (N_11407,N_8900,N_9310);
or U11408 (N_11408,N_8479,N_8776);
xor U11409 (N_11409,N_8414,N_9246);
or U11410 (N_11410,N_8535,N_9851);
nand U11411 (N_11411,N_9961,N_9974);
or U11412 (N_11412,N_8742,N_8477);
nand U11413 (N_11413,N_9529,N_8781);
nor U11414 (N_11414,N_8091,N_9709);
or U11415 (N_11415,N_9121,N_8203);
nand U11416 (N_11416,N_9240,N_9473);
nand U11417 (N_11417,N_9741,N_8256);
xor U11418 (N_11418,N_8976,N_8256);
or U11419 (N_11419,N_8441,N_8976);
xor U11420 (N_11420,N_9484,N_9515);
and U11421 (N_11421,N_8186,N_9306);
nor U11422 (N_11422,N_9168,N_9833);
or U11423 (N_11423,N_8067,N_8015);
xnor U11424 (N_11424,N_9896,N_8769);
and U11425 (N_11425,N_8933,N_9951);
nand U11426 (N_11426,N_9917,N_9138);
or U11427 (N_11427,N_8118,N_8376);
nand U11428 (N_11428,N_9621,N_9224);
nor U11429 (N_11429,N_9222,N_8581);
or U11430 (N_11430,N_9396,N_9798);
and U11431 (N_11431,N_9052,N_8809);
or U11432 (N_11432,N_9656,N_9640);
and U11433 (N_11433,N_9154,N_9103);
nand U11434 (N_11434,N_9549,N_8379);
nand U11435 (N_11435,N_8391,N_9857);
nor U11436 (N_11436,N_8031,N_8647);
nor U11437 (N_11437,N_8782,N_8761);
or U11438 (N_11438,N_8760,N_9736);
and U11439 (N_11439,N_8609,N_8193);
nand U11440 (N_11440,N_9372,N_8229);
or U11441 (N_11441,N_8855,N_9086);
nor U11442 (N_11442,N_9010,N_8274);
nand U11443 (N_11443,N_8207,N_8402);
nand U11444 (N_11444,N_9748,N_8242);
nor U11445 (N_11445,N_9841,N_9281);
and U11446 (N_11446,N_9720,N_9772);
nand U11447 (N_11447,N_8210,N_8710);
or U11448 (N_11448,N_9477,N_8044);
and U11449 (N_11449,N_8306,N_8901);
or U11450 (N_11450,N_8824,N_9842);
xnor U11451 (N_11451,N_8357,N_8815);
nor U11452 (N_11452,N_9194,N_8737);
nand U11453 (N_11453,N_8205,N_8506);
nand U11454 (N_11454,N_9578,N_8928);
xnor U11455 (N_11455,N_9061,N_8159);
nand U11456 (N_11456,N_9230,N_8340);
nor U11457 (N_11457,N_8818,N_8197);
and U11458 (N_11458,N_8715,N_8684);
xnor U11459 (N_11459,N_9766,N_9095);
nand U11460 (N_11460,N_8315,N_9319);
or U11461 (N_11461,N_8259,N_8987);
or U11462 (N_11462,N_9754,N_9005);
or U11463 (N_11463,N_8565,N_8064);
and U11464 (N_11464,N_8635,N_9719);
xnor U11465 (N_11465,N_9684,N_9578);
or U11466 (N_11466,N_8424,N_9344);
xnor U11467 (N_11467,N_9494,N_9293);
nor U11468 (N_11468,N_8779,N_8470);
nor U11469 (N_11469,N_8195,N_9007);
nor U11470 (N_11470,N_8444,N_8665);
and U11471 (N_11471,N_8261,N_9831);
nor U11472 (N_11472,N_9885,N_8835);
nand U11473 (N_11473,N_8509,N_8222);
nor U11474 (N_11474,N_8648,N_9299);
nor U11475 (N_11475,N_8271,N_8540);
or U11476 (N_11476,N_9539,N_8566);
nor U11477 (N_11477,N_8397,N_8130);
nor U11478 (N_11478,N_8865,N_8555);
xnor U11479 (N_11479,N_8294,N_8487);
nor U11480 (N_11480,N_9530,N_9675);
or U11481 (N_11481,N_9658,N_8003);
nand U11482 (N_11482,N_9095,N_8649);
and U11483 (N_11483,N_9082,N_8890);
nand U11484 (N_11484,N_8142,N_9551);
nor U11485 (N_11485,N_8563,N_9096);
or U11486 (N_11486,N_9523,N_9919);
and U11487 (N_11487,N_8638,N_8683);
nand U11488 (N_11488,N_9318,N_8579);
or U11489 (N_11489,N_9697,N_9870);
and U11490 (N_11490,N_8377,N_9695);
xnor U11491 (N_11491,N_9955,N_8110);
and U11492 (N_11492,N_9054,N_8126);
xnor U11493 (N_11493,N_8570,N_8974);
nor U11494 (N_11494,N_9207,N_9459);
nand U11495 (N_11495,N_9787,N_8676);
nor U11496 (N_11496,N_9387,N_9710);
xor U11497 (N_11497,N_9157,N_8817);
xnor U11498 (N_11498,N_8009,N_8048);
or U11499 (N_11499,N_9123,N_8771);
or U11500 (N_11500,N_9868,N_8969);
nand U11501 (N_11501,N_8346,N_9896);
and U11502 (N_11502,N_8855,N_8192);
nor U11503 (N_11503,N_9790,N_8729);
and U11504 (N_11504,N_8664,N_9895);
nand U11505 (N_11505,N_9649,N_8480);
and U11506 (N_11506,N_8869,N_8332);
xnor U11507 (N_11507,N_8311,N_9741);
xor U11508 (N_11508,N_8833,N_8534);
nand U11509 (N_11509,N_9424,N_9682);
xnor U11510 (N_11510,N_9699,N_8613);
nor U11511 (N_11511,N_9879,N_9469);
or U11512 (N_11512,N_8242,N_8183);
nand U11513 (N_11513,N_9057,N_8089);
xor U11514 (N_11514,N_8297,N_9640);
nand U11515 (N_11515,N_9727,N_9498);
xor U11516 (N_11516,N_8555,N_9003);
nand U11517 (N_11517,N_9847,N_8543);
nand U11518 (N_11518,N_9003,N_8222);
xnor U11519 (N_11519,N_9743,N_9932);
nand U11520 (N_11520,N_9912,N_8799);
nor U11521 (N_11521,N_9790,N_8799);
nor U11522 (N_11522,N_8350,N_9095);
and U11523 (N_11523,N_8596,N_9948);
nand U11524 (N_11524,N_9186,N_9260);
xor U11525 (N_11525,N_9818,N_9247);
nor U11526 (N_11526,N_9779,N_8169);
nand U11527 (N_11527,N_9648,N_8757);
xnor U11528 (N_11528,N_9806,N_9802);
or U11529 (N_11529,N_9157,N_8844);
xor U11530 (N_11530,N_9920,N_9071);
xor U11531 (N_11531,N_8982,N_8711);
xor U11532 (N_11532,N_8362,N_8373);
and U11533 (N_11533,N_8975,N_9271);
and U11534 (N_11534,N_8556,N_9464);
xnor U11535 (N_11535,N_9005,N_9049);
xnor U11536 (N_11536,N_8680,N_8456);
nand U11537 (N_11537,N_9343,N_9915);
or U11538 (N_11538,N_9911,N_8290);
xor U11539 (N_11539,N_8333,N_9823);
nor U11540 (N_11540,N_8254,N_8760);
or U11541 (N_11541,N_9756,N_9426);
and U11542 (N_11542,N_9644,N_9579);
and U11543 (N_11543,N_8402,N_8007);
and U11544 (N_11544,N_8521,N_9807);
or U11545 (N_11545,N_8245,N_9569);
or U11546 (N_11546,N_8898,N_8293);
nor U11547 (N_11547,N_9343,N_8063);
nor U11548 (N_11548,N_9842,N_9631);
or U11549 (N_11549,N_9851,N_8760);
nor U11550 (N_11550,N_8615,N_8830);
nor U11551 (N_11551,N_8065,N_9186);
xor U11552 (N_11552,N_8639,N_9911);
nand U11553 (N_11553,N_9250,N_9326);
nor U11554 (N_11554,N_8126,N_9890);
xnor U11555 (N_11555,N_8091,N_9146);
xnor U11556 (N_11556,N_9002,N_9994);
xor U11557 (N_11557,N_8740,N_8625);
and U11558 (N_11558,N_9163,N_8050);
and U11559 (N_11559,N_9128,N_8186);
and U11560 (N_11560,N_9012,N_8167);
and U11561 (N_11561,N_8794,N_9385);
and U11562 (N_11562,N_8786,N_9514);
xor U11563 (N_11563,N_8872,N_8589);
or U11564 (N_11564,N_9511,N_9966);
and U11565 (N_11565,N_8640,N_8043);
xor U11566 (N_11566,N_8172,N_8017);
xnor U11567 (N_11567,N_8834,N_8784);
or U11568 (N_11568,N_9015,N_8910);
nand U11569 (N_11569,N_9962,N_9372);
or U11570 (N_11570,N_9344,N_9785);
or U11571 (N_11571,N_9994,N_9546);
or U11572 (N_11572,N_9574,N_9663);
and U11573 (N_11573,N_9124,N_8120);
nor U11574 (N_11574,N_9403,N_9840);
nor U11575 (N_11575,N_8240,N_8581);
nor U11576 (N_11576,N_8096,N_8289);
xnor U11577 (N_11577,N_9651,N_8509);
nor U11578 (N_11578,N_9090,N_9968);
xnor U11579 (N_11579,N_9030,N_9878);
and U11580 (N_11580,N_9477,N_9635);
or U11581 (N_11581,N_8571,N_8433);
xor U11582 (N_11582,N_9659,N_9549);
nor U11583 (N_11583,N_8649,N_9777);
or U11584 (N_11584,N_8291,N_9558);
or U11585 (N_11585,N_8073,N_9481);
and U11586 (N_11586,N_9646,N_8670);
nor U11587 (N_11587,N_8948,N_9720);
or U11588 (N_11588,N_8848,N_8851);
or U11589 (N_11589,N_9012,N_9102);
nor U11590 (N_11590,N_8028,N_8402);
or U11591 (N_11591,N_9968,N_8906);
or U11592 (N_11592,N_8702,N_8355);
nor U11593 (N_11593,N_8678,N_8969);
nor U11594 (N_11594,N_8616,N_8215);
nand U11595 (N_11595,N_9825,N_9827);
nor U11596 (N_11596,N_9461,N_8145);
and U11597 (N_11597,N_8622,N_8902);
nand U11598 (N_11598,N_8917,N_8670);
nor U11599 (N_11599,N_8574,N_8228);
or U11600 (N_11600,N_8134,N_8938);
nor U11601 (N_11601,N_8231,N_8215);
xnor U11602 (N_11602,N_8294,N_8189);
nand U11603 (N_11603,N_8789,N_8375);
or U11604 (N_11604,N_9302,N_9206);
or U11605 (N_11605,N_9828,N_8930);
xnor U11606 (N_11606,N_8956,N_9548);
nand U11607 (N_11607,N_8049,N_8760);
and U11608 (N_11608,N_9686,N_8420);
or U11609 (N_11609,N_8986,N_9397);
nand U11610 (N_11610,N_9311,N_8941);
nor U11611 (N_11611,N_8155,N_8612);
and U11612 (N_11612,N_8135,N_8456);
and U11613 (N_11613,N_8837,N_8338);
or U11614 (N_11614,N_9065,N_8034);
nand U11615 (N_11615,N_9755,N_8306);
xnor U11616 (N_11616,N_8508,N_8217);
xor U11617 (N_11617,N_9317,N_9702);
xor U11618 (N_11618,N_9691,N_8532);
and U11619 (N_11619,N_8706,N_8945);
xor U11620 (N_11620,N_8855,N_9517);
nor U11621 (N_11621,N_8791,N_9160);
nor U11622 (N_11622,N_9653,N_8761);
xnor U11623 (N_11623,N_9862,N_8951);
or U11624 (N_11624,N_8284,N_8875);
xor U11625 (N_11625,N_8048,N_9833);
nand U11626 (N_11626,N_8206,N_8834);
nor U11627 (N_11627,N_8567,N_8995);
xnor U11628 (N_11628,N_9257,N_9663);
and U11629 (N_11629,N_8451,N_9721);
or U11630 (N_11630,N_9768,N_8374);
and U11631 (N_11631,N_9713,N_8900);
nand U11632 (N_11632,N_8283,N_9580);
nand U11633 (N_11633,N_8811,N_8414);
and U11634 (N_11634,N_9655,N_8762);
nor U11635 (N_11635,N_8269,N_8029);
and U11636 (N_11636,N_8513,N_8476);
and U11637 (N_11637,N_9707,N_8823);
and U11638 (N_11638,N_8850,N_8652);
nand U11639 (N_11639,N_9803,N_8282);
nor U11640 (N_11640,N_9432,N_9698);
or U11641 (N_11641,N_9217,N_9410);
nand U11642 (N_11642,N_9092,N_9428);
or U11643 (N_11643,N_8625,N_9399);
and U11644 (N_11644,N_9515,N_8842);
or U11645 (N_11645,N_9343,N_8767);
nand U11646 (N_11646,N_9343,N_8695);
and U11647 (N_11647,N_8282,N_8105);
nand U11648 (N_11648,N_8338,N_9464);
xnor U11649 (N_11649,N_9351,N_9118);
nor U11650 (N_11650,N_8857,N_9901);
nand U11651 (N_11651,N_9799,N_9982);
nor U11652 (N_11652,N_9887,N_8885);
or U11653 (N_11653,N_8213,N_8845);
nor U11654 (N_11654,N_8193,N_9460);
xor U11655 (N_11655,N_9585,N_9258);
or U11656 (N_11656,N_9816,N_9479);
or U11657 (N_11657,N_8580,N_9200);
xnor U11658 (N_11658,N_9196,N_9669);
or U11659 (N_11659,N_9785,N_9388);
and U11660 (N_11660,N_9486,N_9719);
nor U11661 (N_11661,N_9353,N_8556);
nor U11662 (N_11662,N_9034,N_8988);
nand U11663 (N_11663,N_8197,N_8169);
nor U11664 (N_11664,N_8189,N_8483);
or U11665 (N_11665,N_8049,N_9993);
nor U11666 (N_11666,N_8294,N_9074);
xor U11667 (N_11667,N_9185,N_8660);
xor U11668 (N_11668,N_9440,N_8296);
or U11669 (N_11669,N_8147,N_9243);
nand U11670 (N_11670,N_8445,N_8434);
nor U11671 (N_11671,N_9983,N_8201);
or U11672 (N_11672,N_8356,N_9064);
or U11673 (N_11673,N_8723,N_8566);
and U11674 (N_11674,N_8561,N_8932);
and U11675 (N_11675,N_9144,N_8043);
nand U11676 (N_11676,N_8770,N_8391);
and U11677 (N_11677,N_9728,N_9834);
nor U11678 (N_11678,N_9271,N_8481);
nor U11679 (N_11679,N_9776,N_8285);
or U11680 (N_11680,N_9476,N_9773);
or U11681 (N_11681,N_9359,N_8947);
xor U11682 (N_11682,N_9266,N_8783);
or U11683 (N_11683,N_8799,N_8995);
and U11684 (N_11684,N_8423,N_9005);
and U11685 (N_11685,N_8082,N_9532);
nand U11686 (N_11686,N_9828,N_8596);
xnor U11687 (N_11687,N_8741,N_9272);
or U11688 (N_11688,N_9451,N_9970);
nor U11689 (N_11689,N_9179,N_8118);
xor U11690 (N_11690,N_9567,N_9628);
or U11691 (N_11691,N_8558,N_9237);
nand U11692 (N_11692,N_8625,N_8858);
or U11693 (N_11693,N_9065,N_8960);
xnor U11694 (N_11694,N_9919,N_9430);
nor U11695 (N_11695,N_9636,N_9833);
xor U11696 (N_11696,N_9293,N_8254);
nor U11697 (N_11697,N_9884,N_8181);
or U11698 (N_11698,N_8939,N_8420);
nor U11699 (N_11699,N_9115,N_8784);
nand U11700 (N_11700,N_8944,N_8510);
nand U11701 (N_11701,N_9475,N_9550);
nor U11702 (N_11702,N_9487,N_9016);
nand U11703 (N_11703,N_8934,N_9183);
or U11704 (N_11704,N_8745,N_8888);
and U11705 (N_11705,N_9334,N_9776);
or U11706 (N_11706,N_9315,N_9122);
or U11707 (N_11707,N_9887,N_9803);
or U11708 (N_11708,N_9830,N_8981);
nand U11709 (N_11709,N_9104,N_9411);
nand U11710 (N_11710,N_9525,N_8046);
nand U11711 (N_11711,N_8107,N_9965);
xor U11712 (N_11712,N_9463,N_8151);
or U11713 (N_11713,N_8806,N_8533);
nand U11714 (N_11714,N_8705,N_8860);
nor U11715 (N_11715,N_8824,N_8583);
xnor U11716 (N_11716,N_8133,N_8217);
xnor U11717 (N_11717,N_8840,N_9567);
and U11718 (N_11718,N_9500,N_8360);
or U11719 (N_11719,N_9066,N_8438);
xnor U11720 (N_11720,N_9387,N_9572);
and U11721 (N_11721,N_9142,N_9681);
or U11722 (N_11722,N_9954,N_9155);
or U11723 (N_11723,N_8824,N_9568);
and U11724 (N_11724,N_9001,N_8684);
nor U11725 (N_11725,N_8640,N_8200);
and U11726 (N_11726,N_9213,N_8610);
nor U11727 (N_11727,N_8395,N_9400);
nor U11728 (N_11728,N_9494,N_9831);
or U11729 (N_11729,N_9682,N_8143);
and U11730 (N_11730,N_9717,N_8403);
and U11731 (N_11731,N_8554,N_9996);
xnor U11732 (N_11732,N_9238,N_8604);
nand U11733 (N_11733,N_8447,N_8387);
xnor U11734 (N_11734,N_9111,N_8998);
nand U11735 (N_11735,N_9540,N_8204);
nor U11736 (N_11736,N_9831,N_9621);
and U11737 (N_11737,N_9675,N_8467);
and U11738 (N_11738,N_8137,N_8533);
nand U11739 (N_11739,N_9316,N_8056);
and U11740 (N_11740,N_9489,N_8219);
nor U11741 (N_11741,N_9226,N_9366);
nor U11742 (N_11742,N_8364,N_9045);
or U11743 (N_11743,N_9367,N_8258);
xnor U11744 (N_11744,N_9721,N_8587);
nand U11745 (N_11745,N_8233,N_8137);
or U11746 (N_11746,N_8244,N_9144);
or U11747 (N_11747,N_8346,N_9955);
nor U11748 (N_11748,N_8853,N_9551);
nand U11749 (N_11749,N_9811,N_9052);
nand U11750 (N_11750,N_9995,N_8189);
nand U11751 (N_11751,N_9593,N_9034);
xor U11752 (N_11752,N_8941,N_8682);
xnor U11753 (N_11753,N_9981,N_8343);
and U11754 (N_11754,N_9301,N_8334);
nor U11755 (N_11755,N_9178,N_8783);
nor U11756 (N_11756,N_8391,N_9359);
xor U11757 (N_11757,N_8865,N_9733);
or U11758 (N_11758,N_9870,N_8083);
and U11759 (N_11759,N_9297,N_8057);
xnor U11760 (N_11760,N_8337,N_9944);
or U11761 (N_11761,N_8787,N_8806);
and U11762 (N_11762,N_8033,N_8480);
nor U11763 (N_11763,N_9875,N_9780);
or U11764 (N_11764,N_8964,N_9920);
or U11765 (N_11765,N_8476,N_9614);
nor U11766 (N_11766,N_8737,N_9890);
nor U11767 (N_11767,N_8248,N_8217);
nor U11768 (N_11768,N_9057,N_8675);
nor U11769 (N_11769,N_8025,N_9052);
nor U11770 (N_11770,N_9600,N_8026);
nand U11771 (N_11771,N_9049,N_9260);
or U11772 (N_11772,N_8758,N_8845);
nor U11773 (N_11773,N_9454,N_9605);
xor U11774 (N_11774,N_8156,N_8834);
nand U11775 (N_11775,N_9856,N_9535);
nor U11776 (N_11776,N_8740,N_9220);
and U11777 (N_11777,N_9010,N_9469);
or U11778 (N_11778,N_8723,N_9844);
and U11779 (N_11779,N_9324,N_8204);
xnor U11780 (N_11780,N_9573,N_8404);
xnor U11781 (N_11781,N_8871,N_8832);
xnor U11782 (N_11782,N_8584,N_9219);
or U11783 (N_11783,N_8660,N_9049);
nor U11784 (N_11784,N_8667,N_9689);
nand U11785 (N_11785,N_8566,N_8199);
xor U11786 (N_11786,N_8882,N_8676);
or U11787 (N_11787,N_9854,N_9962);
nand U11788 (N_11788,N_8780,N_9339);
and U11789 (N_11789,N_9302,N_9522);
or U11790 (N_11790,N_9702,N_8439);
nand U11791 (N_11791,N_9123,N_9256);
xor U11792 (N_11792,N_9833,N_9506);
nor U11793 (N_11793,N_9655,N_9998);
nand U11794 (N_11794,N_9527,N_8004);
nand U11795 (N_11795,N_8901,N_9771);
xnor U11796 (N_11796,N_8826,N_8565);
xor U11797 (N_11797,N_9551,N_8581);
nand U11798 (N_11798,N_9844,N_8246);
nor U11799 (N_11799,N_8777,N_9082);
and U11800 (N_11800,N_8545,N_8475);
xnor U11801 (N_11801,N_9588,N_9150);
or U11802 (N_11802,N_9240,N_9955);
or U11803 (N_11803,N_8594,N_9264);
and U11804 (N_11804,N_8383,N_8281);
nor U11805 (N_11805,N_8848,N_8042);
nand U11806 (N_11806,N_8251,N_9390);
nor U11807 (N_11807,N_8075,N_9657);
nor U11808 (N_11808,N_9070,N_9428);
or U11809 (N_11809,N_9506,N_8817);
nor U11810 (N_11810,N_8386,N_8486);
nand U11811 (N_11811,N_9065,N_8590);
and U11812 (N_11812,N_9447,N_9008);
or U11813 (N_11813,N_8412,N_9152);
and U11814 (N_11814,N_8600,N_8259);
xnor U11815 (N_11815,N_9793,N_9502);
nand U11816 (N_11816,N_9304,N_9223);
or U11817 (N_11817,N_8493,N_8392);
and U11818 (N_11818,N_8046,N_9688);
or U11819 (N_11819,N_9119,N_9687);
xor U11820 (N_11820,N_9087,N_9814);
nand U11821 (N_11821,N_8289,N_8243);
nand U11822 (N_11822,N_8156,N_9841);
or U11823 (N_11823,N_8533,N_8588);
nor U11824 (N_11824,N_9302,N_8943);
xnor U11825 (N_11825,N_8390,N_9606);
nor U11826 (N_11826,N_8628,N_9599);
or U11827 (N_11827,N_8767,N_8379);
xor U11828 (N_11828,N_9296,N_9897);
nor U11829 (N_11829,N_9673,N_8819);
nand U11830 (N_11830,N_9729,N_8116);
xnor U11831 (N_11831,N_9875,N_9279);
nor U11832 (N_11832,N_8994,N_8630);
and U11833 (N_11833,N_8807,N_9257);
nor U11834 (N_11834,N_9227,N_8100);
nand U11835 (N_11835,N_9930,N_9826);
or U11836 (N_11836,N_8892,N_9065);
xor U11837 (N_11837,N_9638,N_8867);
nand U11838 (N_11838,N_9560,N_9372);
xnor U11839 (N_11839,N_8518,N_9918);
nor U11840 (N_11840,N_9791,N_8759);
or U11841 (N_11841,N_9565,N_8831);
nor U11842 (N_11842,N_9845,N_9536);
xor U11843 (N_11843,N_9790,N_8690);
or U11844 (N_11844,N_9118,N_9258);
xor U11845 (N_11845,N_9615,N_9234);
xor U11846 (N_11846,N_9032,N_9356);
and U11847 (N_11847,N_9211,N_9785);
xnor U11848 (N_11848,N_9979,N_8162);
nand U11849 (N_11849,N_9300,N_8847);
and U11850 (N_11850,N_9641,N_8040);
nand U11851 (N_11851,N_8575,N_8855);
nor U11852 (N_11852,N_9813,N_8277);
xnor U11853 (N_11853,N_8492,N_9544);
or U11854 (N_11854,N_9655,N_9194);
nor U11855 (N_11855,N_9980,N_8030);
xnor U11856 (N_11856,N_9883,N_8432);
and U11857 (N_11857,N_9774,N_9449);
nand U11858 (N_11858,N_8257,N_9165);
nor U11859 (N_11859,N_9667,N_8570);
xor U11860 (N_11860,N_8218,N_9014);
or U11861 (N_11861,N_9257,N_9524);
or U11862 (N_11862,N_9023,N_8247);
nand U11863 (N_11863,N_9804,N_9240);
nor U11864 (N_11864,N_9940,N_9917);
xnor U11865 (N_11865,N_8387,N_8911);
and U11866 (N_11866,N_8614,N_9102);
xor U11867 (N_11867,N_8628,N_9212);
and U11868 (N_11868,N_8056,N_9228);
or U11869 (N_11869,N_8189,N_8269);
and U11870 (N_11870,N_9301,N_8723);
nor U11871 (N_11871,N_9725,N_9628);
and U11872 (N_11872,N_8862,N_9316);
xnor U11873 (N_11873,N_8068,N_9491);
nor U11874 (N_11874,N_8913,N_9439);
nor U11875 (N_11875,N_8847,N_9904);
nand U11876 (N_11876,N_8014,N_9480);
nor U11877 (N_11877,N_8466,N_9196);
or U11878 (N_11878,N_8759,N_9968);
nand U11879 (N_11879,N_8933,N_8922);
and U11880 (N_11880,N_8401,N_8311);
or U11881 (N_11881,N_8933,N_9944);
nor U11882 (N_11882,N_9152,N_8242);
xnor U11883 (N_11883,N_8874,N_8726);
nor U11884 (N_11884,N_8591,N_9438);
and U11885 (N_11885,N_9172,N_9060);
or U11886 (N_11886,N_8761,N_8250);
nor U11887 (N_11887,N_8438,N_9925);
xnor U11888 (N_11888,N_8055,N_9019);
nor U11889 (N_11889,N_9498,N_8809);
nand U11890 (N_11890,N_9025,N_8213);
nand U11891 (N_11891,N_8349,N_9876);
nand U11892 (N_11892,N_8882,N_9561);
or U11893 (N_11893,N_8864,N_8514);
or U11894 (N_11894,N_9505,N_8930);
xnor U11895 (N_11895,N_8335,N_9413);
and U11896 (N_11896,N_8969,N_9725);
nor U11897 (N_11897,N_9323,N_9468);
nand U11898 (N_11898,N_8158,N_8401);
or U11899 (N_11899,N_9335,N_9194);
nor U11900 (N_11900,N_9050,N_9518);
xor U11901 (N_11901,N_9316,N_9273);
and U11902 (N_11902,N_8717,N_8586);
and U11903 (N_11903,N_8156,N_9414);
and U11904 (N_11904,N_9538,N_9637);
xnor U11905 (N_11905,N_9265,N_8978);
or U11906 (N_11906,N_9002,N_9057);
xor U11907 (N_11907,N_9527,N_9242);
and U11908 (N_11908,N_8758,N_9589);
and U11909 (N_11909,N_9619,N_9169);
xnor U11910 (N_11910,N_8976,N_9065);
xnor U11911 (N_11911,N_8118,N_9786);
xor U11912 (N_11912,N_9664,N_8325);
nand U11913 (N_11913,N_8452,N_8887);
and U11914 (N_11914,N_8593,N_9709);
and U11915 (N_11915,N_9829,N_8656);
and U11916 (N_11916,N_9016,N_9064);
and U11917 (N_11917,N_9655,N_8943);
and U11918 (N_11918,N_9683,N_9867);
or U11919 (N_11919,N_9768,N_8762);
nand U11920 (N_11920,N_9858,N_8898);
or U11921 (N_11921,N_9989,N_8250);
nand U11922 (N_11922,N_8303,N_9928);
nand U11923 (N_11923,N_8447,N_8510);
and U11924 (N_11924,N_8982,N_9655);
or U11925 (N_11925,N_8943,N_8373);
xnor U11926 (N_11926,N_9892,N_9261);
nand U11927 (N_11927,N_9218,N_9664);
xnor U11928 (N_11928,N_9970,N_9233);
and U11929 (N_11929,N_8863,N_8754);
xnor U11930 (N_11930,N_8630,N_8726);
or U11931 (N_11931,N_9208,N_8354);
or U11932 (N_11932,N_8660,N_8377);
nor U11933 (N_11933,N_9838,N_9641);
or U11934 (N_11934,N_9157,N_9635);
or U11935 (N_11935,N_9300,N_8559);
xnor U11936 (N_11936,N_8610,N_9986);
xor U11937 (N_11937,N_9542,N_8801);
and U11938 (N_11938,N_9826,N_9235);
nand U11939 (N_11939,N_9360,N_9556);
nand U11940 (N_11940,N_8911,N_9886);
nand U11941 (N_11941,N_8342,N_9493);
xnor U11942 (N_11942,N_8591,N_8173);
or U11943 (N_11943,N_9343,N_8633);
nor U11944 (N_11944,N_9952,N_9936);
and U11945 (N_11945,N_8472,N_9778);
and U11946 (N_11946,N_8697,N_8364);
nor U11947 (N_11947,N_8183,N_8560);
nand U11948 (N_11948,N_8176,N_8333);
or U11949 (N_11949,N_9300,N_8157);
nand U11950 (N_11950,N_8439,N_8506);
nand U11951 (N_11951,N_8882,N_8745);
nand U11952 (N_11952,N_8294,N_9972);
nand U11953 (N_11953,N_8191,N_9538);
nor U11954 (N_11954,N_9643,N_9722);
nand U11955 (N_11955,N_8259,N_8000);
nand U11956 (N_11956,N_9094,N_8502);
nor U11957 (N_11957,N_9096,N_8986);
xor U11958 (N_11958,N_8967,N_9565);
or U11959 (N_11959,N_8951,N_9028);
xnor U11960 (N_11960,N_9054,N_8299);
nor U11961 (N_11961,N_8072,N_8956);
nor U11962 (N_11962,N_9078,N_8593);
and U11963 (N_11963,N_9059,N_9389);
or U11964 (N_11964,N_8057,N_9538);
and U11965 (N_11965,N_8759,N_9282);
nor U11966 (N_11966,N_9884,N_9901);
or U11967 (N_11967,N_9452,N_9077);
and U11968 (N_11968,N_9851,N_9732);
nand U11969 (N_11969,N_8142,N_8338);
nand U11970 (N_11970,N_8151,N_9641);
xnor U11971 (N_11971,N_8700,N_8127);
and U11972 (N_11972,N_9503,N_8395);
nand U11973 (N_11973,N_9872,N_9321);
nor U11974 (N_11974,N_8352,N_8187);
xnor U11975 (N_11975,N_9671,N_8132);
nand U11976 (N_11976,N_8252,N_8382);
nor U11977 (N_11977,N_9290,N_9298);
nor U11978 (N_11978,N_9316,N_9221);
or U11979 (N_11979,N_8832,N_9694);
nand U11980 (N_11980,N_9229,N_8181);
or U11981 (N_11981,N_9680,N_8240);
and U11982 (N_11982,N_9572,N_8456);
or U11983 (N_11983,N_9702,N_9060);
nand U11984 (N_11984,N_8141,N_9744);
and U11985 (N_11985,N_8691,N_9867);
or U11986 (N_11986,N_8279,N_8946);
nor U11987 (N_11987,N_8509,N_9645);
nand U11988 (N_11988,N_8794,N_9539);
and U11989 (N_11989,N_9088,N_8052);
nand U11990 (N_11990,N_8727,N_8505);
or U11991 (N_11991,N_8783,N_9941);
or U11992 (N_11992,N_8696,N_9894);
and U11993 (N_11993,N_9343,N_8754);
nand U11994 (N_11994,N_9203,N_8400);
nand U11995 (N_11995,N_9029,N_8935);
nor U11996 (N_11996,N_9660,N_9971);
or U11997 (N_11997,N_9866,N_9167);
and U11998 (N_11998,N_8501,N_9655);
and U11999 (N_11999,N_9019,N_8549);
nand U12000 (N_12000,N_10301,N_10261);
or U12001 (N_12001,N_10453,N_11449);
nand U12002 (N_12002,N_10111,N_11855);
and U12003 (N_12003,N_11119,N_10653);
nor U12004 (N_12004,N_10449,N_10953);
xor U12005 (N_12005,N_11423,N_10973);
nand U12006 (N_12006,N_11814,N_10756);
xnor U12007 (N_12007,N_10047,N_11463);
or U12008 (N_12008,N_10750,N_10969);
and U12009 (N_12009,N_10888,N_10843);
nand U12010 (N_12010,N_11764,N_10733);
nand U12011 (N_12011,N_10074,N_11918);
xnor U12012 (N_12012,N_10338,N_11835);
nor U12013 (N_12013,N_11400,N_11544);
nand U12014 (N_12014,N_10977,N_10860);
and U12015 (N_12015,N_11832,N_11729);
xnor U12016 (N_12016,N_10207,N_11316);
xnor U12017 (N_12017,N_11638,N_10367);
xnor U12018 (N_12018,N_10251,N_11741);
or U12019 (N_12019,N_10451,N_11494);
xnor U12020 (N_12020,N_10492,N_11102);
and U12021 (N_12021,N_10085,N_11677);
xnor U12022 (N_12022,N_11435,N_10407);
and U12023 (N_12023,N_10294,N_10565);
nor U12024 (N_12024,N_10838,N_10830);
xnor U12025 (N_12025,N_10109,N_10813);
xor U12026 (N_12026,N_10757,N_10610);
xor U12027 (N_12027,N_11086,N_11155);
and U12028 (N_12028,N_10581,N_11490);
or U12029 (N_12029,N_10429,N_10753);
nand U12030 (N_12030,N_10516,N_10069);
nor U12031 (N_12031,N_10238,N_10172);
xor U12032 (N_12032,N_11129,N_11412);
xnor U12033 (N_12033,N_10186,N_11325);
or U12034 (N_12034,N_11334,N_10649);
xor U12035 (N_12035,N_10450,N_10715);
nand U12036 (N_12036,N_11089,N_10404);
and U12037 (N_12037,N_10331,N_10349);
xnor U12038 (N_12038,N_11194,N_10842);
xnor U12039 (N_12039,N_11784,N_10320);
nand U12040 (N_12040,N_10816,N_11320);
nor U12041 (N_12041,N_10457,N_11515);
and U12042 (N_12042,N_10542,N_11639);
xnor U12043 (N_12043,N_10789,N_10030);
and U12044 (N_12044,N_11927,N_10477);
and U12045 (N_12045,N_11620,N_11486);
and U12046 (N_12046,N_10209,N_11592);
or U12047 (N_12047,N_10532,N_10835);
or U12048 (N_12048,N_10593,N_11771);
and U12049 (N_12049,N_10932,N_10180);
nand U12050 (N_12050,N_11507,N_10052);
or U12051 (N_12051,N_11475,N_11642);
nand U12052 (N_12052,N_10206,N_11734);
and U12053 (N_12053,N_10306,N_10271);
or U12054 (N_12054,N_10812,N_11285);
or U12055 (N_12055,N_10675,N_11436);
nor U12056 (N_12056,N_10595,N_10668);
xor U12057 (N_12057,N_10926,N_11870);
and U12058 (N_12058,N_10295,N_10431);
and U12059 (N_12059,N_11452,N_10131);
and U12060 (N_12060,N_11021,N_10316);
nand U12061 (N_12061,N_11221,N_11836);
xnor U12062 (N_12062,N_10585,N_11117);
or U12063 (N_12063,N_10469,N_10865);
or U12064 (N_12064,N_10168,N_11665);
or U12065 (N_12065,N_11231,N_10150);
or U12066 (N_12066,N_10483,N_11902);
and U12067 (N_12067,N_11685,N_11422);
and U12068 (N_12068,N_10101,N_11492);
nor U12069 (N_12069,N_11479,N_10397);
xnor U12070 (N_12070,N_11396,N_10994);
nor U12071 (N_12071,N_11482,N_11889);
xnor U12072 (N_12072,N_10541,N_10575);
and U12073 (N_12073,N_11055,N_10600);
nand U12074 (N_12074,N_11225,N_11719);
or U12075 (N_12075,N_10126,N_11458);
and U12076 (N_12076,N_11159,N_10672);
xor U12077 (N_12077,N_11499,N_11502);
or U12078 (N_12078,N_11590,N_10577);
and U12079 (N_12079,N_10006,N_10696);
nor U12080 (N_12080,N_10856,N_11358);
xor U12081 (N_12081,N_10745,N_10480);
or U12082 (N_12082,N_11271,N_11846);
and U12083 (N_12083,N_10989,N_11333);
and U12084 (N_12084,N_11104,N_10032);
and U12085 (N_12085,N_11017,N_11774);
xor U12086 (N_12086,N_11331,N_10370);
nor U12087 (N_12087,N_11024,N_11687);
xor U12088 (N_12088,N_10341,N_11173);
nand U12089 (N_12089,N_10748,N_11063);
nand U12090 (N_12090,N_11748,N_10354);
and U12091 (N_12091,N_10970,N_10523);
nor U12092 (N_12092,N_11361,N_10257);
or U12093 (N_12093,N_11876,N_10592);
nand U12094 (N_12094,N_10702,N_11552);
nor U12095 (N_12095,N_10667,N_10379);
and U12096 (N_12096,N_11978,N_10440);
xor U12097 (N_12097,N_11064,N_11296);
nor U12098 (N_12098,N_10158,N_11007);
xnor U12099 (N_12099,N_11852,N_11935);
xnor U12100 (N_12100,N_10405,N_10080);
or U12101 (N_12101,N_10014,N_11817);
and U12102 (N_12102,N_11197,N_10227);
xnor U12103 (N_12103,N_11939,N_10285);
xor U12104 (N_12104,N_11897,N_10466);
or U12105 (N_12105,N_11663,N_11560);
or U12106 (N_12106,N_10139,N_11212);
nor U12107 (N_12107,N_10004,N_11951);
nor U12108 (N_12108,N_11455,N_10627);
or U12109 (N_12109,N_11954,N_10554);
nand U12110 (N_12110,N_10693,N_10375);
and U12111 (N_12111,N_11080,N_11156);
nor U12112 (N_12112,N_10252,N_10095);
xnor U12113 (N_12113,N_10652,N_11795);
or U12114 (N_12114,N_10707,N_11359);
nor U12115 (N_12115,N_11084,N_11972);
xnor U12116 (N_12116,N_10722,N_11550);
nand U12117 (N_12117,N_11009,N_11912);
or U12118 (N_12118,N_11374,N_11780);
nand U12119 (N_12119,N_11433,N_10659);
or U12120 (N_12120,N_11875,N_11793);
nand U12121 (N_12121,N_10670,N_11506);
and U12122 (N_12122,N_10894,N_10275);
or U12123 (N_12123,N_11208,N_11997);
nand U12124 (N_12124,N_11066,N_10372);
nor U12125 (N_12125,N_10007,N_11969);
nor U12126 (N_12126,N_10233,N_10679);
nor U12127 (N_12127,N_10226,N_11987);
nor U12128 (N_12128,N_10084,N_10521);
nor U12129 (N_12129,N_11848,N_11467);
or U12130 (N_12130,N_11085,N_11022);
xnor U12131 (N_12131,N_10414,N_11146);
and U12132 (N_12132,N_11603,N_11018);
xor U12133 (N_12133,N_11892,N_11053);
or U12134 (N_12134,N_10852,N_10986);
or U12135 (N_12135,N_11770,N_10772);
and U12136 (N_12136,N_10921,N_11858);
nand U12137 (N_12137,N_11723,N_10942);
nand U12138 (N_12138,N_10923,N_10828);
nor U12139 (N_12139,N_11120,N_11382);
xor U12140 (N_12140,N_10694,N_11006);
nand U12141 (N_12141,N_10445,N_10773);
nor U12142 (N_12142,N_11167,N_10132);
nand U12143 (N_12143,N_11440,N_11177);
nand U12144 (N_12144,N_11641,N_11478);
nand U12145 (N_12145,N_10955,N_11329);
and U12146 (N_12146,N_11139,N_10931);
nand U12147 (N_12147,N_10505,N_10943);
or U12148 (N_12148,N_11984,N_10690);
or U12149 (N_12149,N_10784,N_11392);
xnor U12150 (N_12150,N_10189,N_11035);
nand U12151 (N_12151,N_11791,N_10870);
and U12152 (N_12152,N_11658,N_11121);
or U12153 (N_12153,N_10990,N_10157);
nor U12154 (N_12154,N_11568,N_11404);
and U12155 (N_12155,N_11803,N_11008);
nand U12156 (N_12156,N_11116,N_10272);
nand U12157 (N_12157,N_11686,N_11558);
or U12158 (N_12158,N_11352,N_11726);
and U12159 (N_12159,N_10120,N_10549);
and U12160 (N_12160,N_10012,N_10650);
and U12161 (N_12161,N_10358,N_10642);
xnor U12162 (N_12162,N_11232,N_11027);
or U12163 (N_12163,N_10918,N_10009);
and U12164 (N_12164,N_11067,N_11344);
xnor U12165 (N_12165,N_11189,N_11087);
or U12166 (N_12166,N_10082,N_10321);
xnor U12167 (N_12167,N_10826,N_10971);
nor U12168 (N_12168,N_10562,N_10395);
and U12169 (N_12169,N_11673,N_11269);
and U12170 (N_12170,N_11806,N_11815);
nor U12171 (N_12171,N_11058,N_10844);
and U12172 (N_12172,N_10897,N_10558);
nor U12173 (N_12173,N_11300,N_10712);
and U12174 (N_12174,N_11763,N_10570);
and U12175 (N_12175,N_10956,N_10783);
xor U12176 (N_12176,N_11580,N_10478);
nand U12177 (N_12177,N_11323,N_11233);
and U12178 (N_12178,N_11666,N_11701);
and U12179 (N_12179,N_11275,N_10669);
xor U12180 (N_12180,N_10017,N_10485);
nand U12181 (N_12181,N_10335,N_11670);
xor U12182 (N_12182,N_10311,N_11536);
and U12183 (N_12183,N_11766,N_10064);
xor U12184 (N_12184,N_11759,N_11346);
and U12185 (N_12185,N_11448,N_10645);
and U12186 (N_12186,N_11838,N_10471);
xor U12187 (N_12187,N_11483,N_11512);
xnor U12188 (N_12188,N_10269,N_10966);
and U12189 (N_12189,N_10329,N_11210);
nor U12190 (N_12190,N_11469,N_11775);
xnor U12191 (N_12191,N_11958,N_10183);
nand U12192 (N_12192,N_11270,N_11751);
nand U12193 (N_12193,N_11122,N_11924);
and U12194 (N_12194,N_10768,N_10054);
or U12195 (N_12195,N_10576,N_11188);
nor U12196 (N_12196,N_10435,N_10152);
nor U12197 (N_12197,N_11247,N_10347);
and U12198 (N_12198,N_11281,N_11330);
xnor U12199 (N_12199,N_10447,N_10851);
nor U12200 (N_12200,N_11576,N_10845);
or U12201 (N_12201,N_11733,N_11611);
nand U12202 (N_12202,N_10617,N_10580);
or U12203 (N_12203,N_11246,N_10114);
or U12204 (N_12204,N_10859,N_11446);
nand U12205 (N_12205,N_11174,N_10099);
nor U12206 (N_12206,N_11394,N_11150);
nor U12207 (N_12207,N_11800,N_10946);
or U12208 (N_12208,N_10657,N_10190);
or U12209 (N_12209,N_11740,N_11822);
nand U12210 (N_12210,N_10706,N_11204);
and U12211 (N_12211,N_10680,N_11168);
and U12212 (N_12212,N_10950,N_10105);
nand U12213 (N_12213,N_11322,N_11657);
nor U12214 (N_12214,N_11427,N_11886);
and U12215 (N_12215,N_11471,N_10598);
and U12216 (N_12216,N_10513,N_10040);
and U12217 (N_12217,N_11501,N_10046);
nor U12218 (N_12218,N_10217,N_11513);
or U12219 (N_12219,N_11096,N_10028);
and U12220 (N_12220,N_11082,N_11138);
or U12221 (N_12221,N_11586,N_11634);
nand U12222 (N_12222,N_11708,N_10276);
and U12223 (N_12223,N_10980,N_11454);
or U12224 (N_12224,N_10059,N_11481);
or U12225 (N_12225,N_11625,N_10042);
nor U12226 (N_12226,N_11294,N_11306);
or U12227 (N_12227,N_11430,N_11011);
and U12228 (N_12228,N_11600,N_10005);
or U12229 (N_12229,N_10391,N_10023);
or U12230 (N_12230,N_10530,N_11079);
xnor U12231 (N_12231,N_11010,N_11083);
nand U12232 (N_12232,N_10548,N_11851);
and U12233 (N_12233,N_10566,N_11599);
nor U12234 (N_12234,N_10991,N_11738);
nand U12235 (N_12235,N_10602,N_10146);
xnor U12236 (N_12236,N_10929,N_10547);
and U12237 (N_12237,N_11746,N_11187);
nand U12238 (N_12238,N_10415,N_11960);
and U12239 (N_12239,N_10070,N_10409);
or U12240 (N_12240,N_10277,N_11991);
nor U12241 (N_12241,N_11183,N_11700);
nand U12242 (N_12242,N_11389,N_11111);
nand U12243 (N_12243,N_11750,N_11514);
nor U12244 (N_12244,N_10605,N_10197);
nand U12245 (N_12245,N_11714,N_11324);
xnor U12246 (N_12246,N_10102,N_11240);
nor U12247 (N_12247,N_10458,N_11098);
nor U12248 (N_12248,N_11789,N_11092);
and U12249 (N_12249,N_11107,N_11805);
or U12250 (N_12250,N_11689,N_11033);
and U12251 (N_12251,N_10219,N_10319);
xnor U12252 (N_12252,N_11443,N_11439);
nand U12253 (N_12253,N_11676,N_10303);
nor U12254 (N_12254,N_10965,N_10116);
nand U12255 (N_12255,N_10947,N_10903);
xnor U12256 (N_12256,N_10976,N_11180);
nand U12257 (N_12257,N_11543,N_11635);
xnor U12258 (N_12258,N_10821,N_10591);
or U12259 (N_12259,N_10951,N_11172);
xnor U12260 (N_12260,N_11081,N_10635);
xnor U12261 (N_12261,N_10801,N_11266);
xnor U12262 (N_12262,N_11200,N_11056);
or U12263 (N_12263,N_10434,N_10160);
xnor U12264 (N_12264,N_10736,N_11794);
nand U12265 (N_12265,N_11853,N_11061);
or U12266 (N_12266,N_10872,N_11651);
xor U12267 (N_12267,N_11702,N_11533);
and U12268 (N_12268,N_11088,N_11664);
xor U12269 (N_12269,N_11253,N_11953);
and U12270 (N_12270,N_10960,N_11153);
or U12271 (N_12271,N_11798,N_11627);
and U12272 (N_12272,N_11785,N_11591);
nand U12273 (N_12273,N_10709,N_11048);
or U12274 (N_12274,N_10608,N_10130);
nor U12275 (N_12275,N_10545,N_10169);
and U12276 (N_12276,N_11967,N_11808);
xnor U12277 (N_12277,N_10170,N_11069);
and U12278 (N_12278,N_10215,N_11585);
nor U12279 (N_12279,N_10840,N_10460);
and U12280 (N_12280,N_10156,N_10728);
and U12281 (N_12281,N_10462,N_11337);
xnor U12282 (N_12282,N_11224,N_10097);
xor U12283 (N_12283,N_10839,N_11047);
nand U12284 (N_12284,N_11818,N_11961);
or U12285 (N_12285,N_11531,N_11721);
and U12286 (N_12286,N_11937,N_11660);
nand U12287 (N_12287,N_11100,N_10421);
nor U12288 (N_12288,N_10297,N_11621);
nand U12289 (N_12289,N_11850,N_10355);
and U12290 (N_12290,N_10448,N_10310);
or U12291 (N_12291,N_10270,N_10501);
and U12292 (N_12292,N_11199,N_10472);
nand U12293 (N_12293,N_10230,N_10735);
nand U12294 (N_12294,N_11613,N_11073);
and U12295 (N_12295,N_11674,N_10115);
xnor U12296 (N_12296,N_10802,N_11354);
xor U12297 (N_12297,N_11162,N_11557);
nor U12298 (N_12298,N_10142,N_10616);
or U12299 (N_12299,N_10621,N_10896);
or U12300 (N_12300,N_10198,N_11273);
or U12301 (N_12301,N_10825,N_11608);
nor U12302 (N_12302,N_10351,N_11095);
nor U12303 (N_12303,N_11518,N_11843);
or U12304 (N_12304,N_10237,N_10881);
or U12305 (N_12305,N_11690,N_10491);
xor U12306 (N_12306,N_11348,N_11259);
xor U12307 (N_12307,N_11052,N_11920);
xnor U12308 (N_12308,N_11353,N_10535);
or U12309 (N_12309,N_11014,N_11787);
or U12310 (N_12310,N_10326,N_11547);
nand U12311 (N_12311,N_10242,N_10473);
nor U12312 (N_12312,N_11417,N_10537);
nand U12313 (N_12313,N_11143,N_11712);
and U12314 (N_12314,N_11632,N_10727);
nor U12315 (N_12315,N_11828,N_11526);
or U12316 (N_12316,N_10543,N_11881);
or U12317 (N_12317,N_10436,N_10412);
and U12318 (N_12318,N_10454,N_10569);
or U12319 (N_12319,N_10673,N_11649);
nand U12320 (N_12320,N_11235,N_11288);
nor U12321 (N_12321,N_11768,N_10777);
nand U12322 (N_12322,N_10360,N_10018);
or U12323 (N_12323,N_11470,N_11196);
nand U12324 (N_12324,N_11145,N_10873);
nand U12325 (N_12325,N_10463,N_10117);
xor U12326 (N_12326,N_11908,N_11391);
xnor U12327 (N_12327,N_10193,N_10599);
xor U12328 (N_12328,N_10705,N_10999);
nor U12329 (N_12329,N_11308,N_10945);
xnor U12330 (N_12330,N_11801,N_11041);
nand U12331 (N_12331,N_11704,N_11519);
xor U12332 (N_12332,N_10258,N_10920);
nand U12333 (N_12333,N_10879,N_11681);
or U12334 (N_12334,N_10380,N_10824);
nand U12335 (N_12335,N_10368,N_10939);
nand U12336 (N_12336,N_11819,N_10557);
nand U12337 (N_12337,N_11957,N_11248);
or U12338 (N_12338,N_10254,N_10717);
nand U12339 (N_12339,N_11466,N_10244);
nand U12340 (N_12340,N_10029,N_10222);
xnor U12341 (N_12341,N_11134,N_10744);
nand U12342 (N_12342,N_11037,N_11877);
and U12343 (N_12343,N_11860,N_11866);
or U12344 (N_12344,N_11534,N_10459);
or U12345 (N_12345,N_10519,N_10282);
nand U12346 (N_12346,N_11979,N_11397);
or U12347 (N_12347,N_11165,N_11461);
xnor U12348 (N_12348,N_10893,N_10857);
nor U12349 (N_12349,N_10922,N_10787);
and U12350 (N_12350,N_10676,N_11522);
or U12351 (N_12351,N_11103,N_10377);
nand U12352 (N_12352,N_11065,N_10967);
and U12353 (N_12353,N_11113,N_10406);
or U12354 (N_12354,N_11636,N_10781);
or U12355 (N_12355,N_10629,N_11698);
xnor U12356 (N_12356,N_11899,N_10867);
nor U12357 (N_12357,N_10214,N_11661);
and U12358 (N_12358,N_11562,N_11890);
nand U12359 (N_12359,N_11807,N_10475);
nand U12360 (N_12360,N_11206,N_10666);
xnor U12361 (N_12361,N_11549,N_11442);
nand U12362 (N_12362,N_10411,N_10098);
nor U12363 (N_12363,N_10831,N_11377);
nand U12364 (N_12364,N_10509,N_10941);
xor U12365 (N_12365,N_11587,N_11809);
or U12366 (N_12366,N_10201,N_10034);
or U12367 (N_12367,N_11276,N_11693);
or U12368 (N_12368,N_11026,N_11133);
xor U12369 (N_12369,N_11216,N_10268);
nand U12370 (N_12370,N_10322,N_11643);
nor U12371 (N_12371,N_10742,N_10441);
xnor U12372 (N_12372,N_10100,N_11307);
nor U12373 (N_12373,N_11730,N_10484);
nand U12374 (N_12374,N_10353,N_11871);
and U12375 (N_12375,N_11123,N_11078);
nand U12376 (N_12376,N_10935,N_11313);
xor U12377 (N_12377,N_10620,N_11994);
nor U12378 (N_12378,N_11101,N_11000);
and U12379 (N_12379,N_10318,N_10253);
xor U12380 (N_12380,N_10751,N_11472);
or U12381 (N_12381,N_11706,N_11769);
and U12382 (N_12382,N_11570,N_11343);
nor U12383 (N_12383,N_11754,N_10737);
xnor U12384 (N_12384,N_10281,N_10755);
and U12385 (N_12385,N_10399,N_10661);
xor U12386 (N_12386,N_10804,N_10770);
xor U12387 (N_12387,N_11952,N_11198);
xor U12388 (N_12388,N_10936,N_10136);
and U12389 (N_12389,N_10555,N_11465);
and U12390 (N_12390,N_11955,N_10361);
nand U12391 (N_12391,N_10489,N_10015);
nor U12392 (N_12392,N_11287,N_11906);
nor U12393 (N_12393,N_10741,N_10641);
or U12394 (N_12394,N_10563,N_10604);
or U12395 (N_12395,N_10263,N_10300);
or U12396 (N_12396,N_11255,N_11388);
and U12397 (N_12397,N_11596,N_10432);
xnor U12398 (N_12398,N_10766,N_10815);
xnor U12399 (N_12399,N_11130,N_11094);
nor U12400 (N_12400,N_10344,N_11762);
xor U12401 (N_12401,N_11564,N_10568);
nand U12402 (N_12402,N_10143,N_11756);
nor U12403 (N_12403,N_11630,N_11301);
nor U12404 (N_12404,N_10293,N_10056);
xnor U12405 (N_12405,N_10880,N_11873);
nand U12406 (N_12406,N_10767,N_11421);
nor U12407 (N_12407,N_10041,N_11988);
or U12408 (N_12408,N_10243,N_10240);
and U12409 (N_12409,N_10248,N_10882);
nand U12410 (N_12410,N_10154,N_10914);
xor U12411 (N_12411,N_10196,N_11995);
and U12412 (N_12412,N_10901,N_11757);
or U12413 (N_12413,N_11171,N_10119);
xnor U12414 (N_12414,N_10045,N_11857);
xor U12415 (N_12415,N_11732,N_11508);
nor U12416 (N_12416,N_11106,N_10841);
and U12417 (N_12417,N_11409,N_11679);
nand U12418 (N_12418,N_10993,N_10356);
and U12419 (N_12419,N_10020,N_10692);
nand U12420 (N_12420,N_11824,N_10691);
nor U12421 (N_12421,N_10072,N_10155);
and U12422 (N_12422,N_11050,N_10374);
nand U12423 (N_12423,N_11245,N_11473);
nor U12424 (N_12424,N_11616,N_10503);
nand U12425 (N_12425,N_11584,N_11124);
or U12426 (N_12426,N_10615,N_10493);
nand U12427 (N_12427,N_11090,N_11390);
nand U12428 (N_12428,N_10626,N_10224);
xnor U12429 (N_12429,N_11191,N_11727);
or U12430 (N_12430,N_11413,N_11802);
or U12431 (N_12431,N_11662,N_10556);
xor U12432 (N_12432,N_10027,N_10531);
xor U12433 (N_12433,N_10400,N_10799);
and U12434 (N_12434,N_10518,N_11609);
or U12435 (N_12435,N_10315,N_11274);
xnor U12436 (N_12436,N_10797,N_10091);
or U12437 (N_12437,N_10868,N_10245);
and U12438 (N_12438,N_11251,N_11796);
nand U12439 (N_12439,N_11511,N_11811);
and U12440 (N_12440,N_11215,N_11707);
or U12441 (N_12441,N_11856,N_10975);
nor U12442 (N_12442,N_10529,N_11783);
nor U12443 (N_12443,N_10247,N_10948);
nor U12444 (N_12444,N_10752,N_11864);
nor U12445 (N_12445,N_10810,N_11882);
and U12446 (N_12446,N_11309,N_11367);
and U12447 (N_12447,N_10633,N_10063);
or U12448 (N_12448,N_11234,N_11581);
nand U12449 (N_12449,N_10749,N_10776);
or U12450 (N_12450,N_10145,N_10731);
nor U12451 (N_12451,N_10520,N_11767);
and U12452 (N_12452,N_10836,N_10452);
xor U12453 (N_12453,N_10166,N_10930);
nor U12454 (N_12454,N_11051,N_10678);
xnor U12455 (N_12455,N_11114,N_10758);
nor U12456 (N_12456,N_10236,N_11914);
nor U12457 (N_12457,N_11545,N_10759);
nand U12458 (N_12458,N_11804,N_11347);
nor U12459 (N_12459,N_10979,N_11487);
nor U12460 (N_12460,N_11001,N_11559);
or U12461 (N_12461,N_10579,N_10181);
xnor U12462 (N_12462,N_10113,N_11386);
nand U12463 (N_12463,N_11148,N_10078);
and U12464 (N_12464,N_10439,N_11016);
or U12465 (N_12465,N_11823,N_10832);
nor U12466 (N_12466,N_10764,N_11077);
xnor U12467 (N_12467,N_11284,N_10444);
nor U12468 (N_12468,N_11297,N_10195);
and U12469 (N_12469,N_11376,N_10220);
nor U12470 (N_12470,N_10647,N_11108);
or U12471 (N_12471,N_11779,N_11341);
xnor U12472 (N_12472,N_10202,N_10433);
nor U12473 (N_12473,N_10507,N_11151);
xor U12474 (N_12474,N_10008,N_10044);
nand U12475 (N_12475,N_10818,N_10286);
xnor U12476 (N_12476,N_10022,N_10417);
or U12477 (N_12477,N_11761,N_11626);
or U12478 (N_12478,N_11911,N_11099);
or U12479 (N_12479,N_11737,N_10192);
and U12480 (N_12480,N_11202,N_11656);
or U12481 (N_12481,N_11773,N_10010);
nand U12482 (N_12482,N_11910,N_10339);
or U12483 (N_12483,N_10144,N_10333);
and U12484 (N_12484,N_11476,N_11311);
and U12485 (N_12485,N_11985,N_10389);
nor U12486 (N_12486,N_10283,N_11975);
xnor U12487 (N_12487,N_10438,N_10304);
xor U12488 (N_12488,N_10289,N_10849);
nand U12489 (N_12489,N_10944,N_10016);
nand U12490 (N_12490,N_10365,N_10687);
nand U12491 (N_12491,N_10985,N_11989);
nor U12492 (N_12492,N_10298,N_11993);
xor U12493 (N_12493,N_11220,N_11068);
nor U12494 (N_12494,N_11414,N_11060);
and U12495 (N_12495,N_10163,N_10246);
or U12496 (N_12496,N_10915,N_10790);
xnor U12497 (N_12497,N_10949,N_11368);
nor U12498 (N_12498,N_11419,N_10239);
or U12499 (N_12499,N_10278,N_10508);
and U12500 (N_12500,N_11525,N_11878);
nand U12501 (N_12501,N_11540,N_11527);
nor U12502 (N_12502,N_11810,N_11227);
and U12503 (N_12503,N_10628,N_11426);
or U12504 (N_12504,N_11236,N_11922);
xor U12505 (N_12505,N_11678,N_10601);
or U12506 (N_12506,N_10031,N_10437);
xnor U12507 (N_12507,N_10234,N_11289);
and U12508 (N_12508,N_10798,N_10771);
and U12509 (N_12509,N_11556,N_10681);
nand U12510 (N_12510,N_11593,N_11614);
nor U12511 (N_12511,N_10874,N_10885);
nor U12512 (N_12512,N_11012,N_10788);
nor U12513 (N_12513,N_11725,N_10995);
nor U12514 (N_12514,N_11328,N_10952);
nor U12515 (N_12515,N_11578,N_10890);
xnor U12516 (N_12516,N_11900,N_10066);
nand U12517 (N_12517,N_11713,N_11896);
or U12518 (N_12518,N_10312,N_11555);
nand U12519 (N_12519,N_10465,N_10820);
and U12520 (N_12520,N_11976,N_10786);
xnor U12521 (N_12521,N_10829,N_10288);
and U12522 (N_12522,N_10905,N_10408);
nand U12523 (N_12523,N_10211,N_10637);
and U12524 (N_12524,N_11589,N_11990);
and U12525 (N_12525,N_10262,N_11260);
or U12526 (N_12526,N_10050,N_11447);
xnor U12527 (N_12527,N_10654,N_10382);
or U12528 (N_12528,N_10422,N_11229);
nand U12529 (N_12529,N_11749,N_11974);
or U12530 (N_12530,N_10928,N_11901);
nand U12531 (N_12531,N_11597,N_10803);
nor U12532 (N_12532,N_11885,N_10345);
xnor U12533 (N_12533,N_11028,N_10589);
nor U12534 (N_12534,N_11040,N_10959);
or U12535 (N_12535,N_10596,N_11338);
and U12536 (N_12536,N_10369,N_10517);
nand U12537 (N_12537,N_10396,N_11977);
nor U12538 (N_12538,N_10001,N_11314);
or U12539 (N_12539,N_11049,N_10583);
nand U12540 (N_12540,N_11854,N_11075);
xnor U12541 (N_12541,N_11500,N_10175);
and U12542 (N_12542,N_11760,N_11339);
nor U12543 (N_12543,N_10231,N_10121);
xor U12544 (N_12544,N_10747,N_10571);
nor U12545 (N_12545,N_10188,N_11318);
nand U12546 (N_12546,N_10340,N_10809);
and U12547 (N_12547,N_10038,N_10096);
or U12548 (N_12548,N_10313,N_11302);
nor U12549 (N_12549,N_11485,N_10076);
nand U12550 (N_12550,N_11640,N_11812);
or U12551 (N_12551,N_11601,N_10714);
and U12552 (N_12552,N_10847,N_10765);
or U12553 (N_12553,N_10291,N_10364);
or U12554 (N_12554,N_10148,N_11573);
nor U12555 (N_12555,N_11753,N_11820);
xnor U12556 (N_12556,N_10336,N_11934);
or U12557 (N_12557,N_10643,N_11916);
and U12558 (N_12558,N_10587,N_11859);
or U12559 (N_12559,N_10264,N_11747);
xnor U12560 (N_12560,N_10323,N_11940);
and U12561 (N_12561,N_11249,N_10983);
nor U12562 (N_12562,N_11862,N_11965);
nor U12563 (N_12563,N_10249,N_10997);
nand U12564 (N_12564,N_10792,N_11699);
or U12565 (N_12565,N_10837,N_10470);
and U12566 (N_12566,N_11628,N_10387);
xor U12567 (N_12567,N_11264,N_10394);
or U12568 (N_12568,N_11416,N_10039);
nor U12569 (N_12569,N_11046,N_11034);
nand U12570 (N_12570,N_10625,N_11157);
and U12571 (N_12571,N_11244,N_11542);
nor U12572 (N_12572,N_11709,N_11497);
nand U12573 (N_12573,N_11036,N_10062);
xnor U12574 (N_12574,N_11336,N_10512);
nand U12575 (N_12575,N_11136,N_10924);
nand U12576 (N_12576,N_10068,N_10332);
xnor U12577 (N_12577,N_10123,N_11583);
and U12578 (N_12578,N_10863,N_10684);
nor U12579 (N_12579,N_11291,N_10938);
xnor U12580 (N_12580,N_11831,N_10055);
xor U12581 (N_12581,N_11379,N_11647);
or U12582 (N_12582,N_10464,N_10425);
or U12583 (N_12583,N_10586,N_10682);
or U12584 (N_12584,N_11618,N_10528);
and U12585 (N_12585,N_10685,N_10497);
nand U12586 (N_12586,N_11013,N_11813);
nand U12587 (N_12587,N_10533,N_10194);
nor U12588 (N_12588,N_11261,N_10711);
nand U12589 (N_12589,N_10800,N_11450);
nand U12590 (N_12590,N_11335,N_10594);
and U12591 (N_12591,N_11844,N_11312);
and U12592 (N_12592,N_11943,N_11303);
xnor U12593 (N_12593,N_10919,N_11538);
or U12594 (N_12594,N_11509,N_10255);
nor U12595 (N_12595,N_10287,N_10567);
nor U12596 (N_12596,N_11403,N_10392);
nand U12597 (N_12597,N_11680,N_10504);
xor U12598 (N_12598,N_10461,N_10739);
xor U12599 (N_12599,N_11968,N_11837);
nor U12600 (N_12600,N_11149,N_11267);
and U12601 (N_12601,N_11137,N_10796);
or U12602 (N_12602,N_10762,N_11605);
nand U12603 (N_12603,N_11371,N_10573);
xnor U12604 (N_12604,N_10913,N_10216);
and U12605 (N_12605,N_10546,N_11459);
and U12606 (N_12606,N_10002,N_11032);
nand U12607 (N_12607,N_11863,N_10662);
nor U12608 (N_12608,N_10071,N_10700);
nand U12609 (N_12609,N_10147,N_11893);
nor U12610 (N_12610,N_11743,N_10420);
or U12611 (N_12611,N_11326,N_10636);
nor U12612 (N_12612,N_10309,N_10371);
nand U12613 (N_12613,N_11973,N_11283);
and U12614 (N_12614,N_10141,N_10611);
nand U12615 (N_12615,N_11201,N_11282);
or U12616 (N_12616,N_11938,N_10877);
and U12617 (N_12617,N_10419,N_11539);
xor U12618 (N_12618,N_10205,N_11395);
or U12619 (N_12619,N_10984,N_11744);
nor U12620 (N_12620,N_10384,N_11002);
or U12621 (N_12621,N_11265,N_10560);
nand U12622 (N_12622,N_11728,N_11140);
and U12623 (N_12623,N_11410,N_10021);
and U12624 (N_12624,N_11521,N_10607);
nand U12625 (N_12625,N_10992,N_11998);
or U12626 (N_12626,N_10934,N_10362);
nand U12627 (N_12627,N_10525,N_11147);
or U12628 (N_12628,N_10719,N_11909);
xnor U12629 (N_12629,N_11385,N_11498);
nand U12630 (N_12630,N_10357,N_10515);
xor U12631 (N_12631,N_10699,N_10378);
or U12632 (N_12632,N_10634,N_11716);
nor U12633 (N_12633,N_11765,N_10574);
and U12634 (N_12634,N_10035,N_11703);
nand U12635 (N_12635,N_11420,N_10916);
and U12636 (N_12636,N_10721,N_11424);
and U12637 (N_12637,N_10416,N_11905);
xnor U12638 (N_12638,N_11895,N_10184);
xor U12639 (N_12639,N_10743,N_10875);
nand U12640 (N_12640,N_11445,N_11160);
nor U12641 (N_12641,N_10663,N_10496);
xnor U12642 (N_12642,N_11141,N_10486);
nand U12643 (N_12643,N_10363,N_10089);
and U12644 (N_12644,N_10499,N_11127);
nor U12645 (N_12645,N_10446,N_10551);
nand U12646 (N_12646,N_11971,N_10088);
xor U12647 (N_12647,N_11484,N_11963);
and U12648 (N_12648,N_10094,N_10871);
and U12649 (N_12649,N_10129,N_11238);
and U12650 (N_12650,N_10987,N_10887);
nand U12651 (N_12651,N_11691,N_11154);
or U12652 (N_12652,N_11203,N_10514);
nand U12653 (N_12653,N_11186,N_10500);
nand U12654 (N_12654,N_10876,N_10122);
nand U12655 (N_12655,N_10037,N_11115);
nor U12656 (N_12656,N_11671,N_11668);
and U12657 (N_12657,N_11169,N_11563);
or U12658 (N_12658,N_11982,N_11411);
and U12659 (N_12659,N_10302,N_10228);
nand U12660 (N_12660,N_11782,N_11223);
nor U12661 (N_12661,N_10390,N_11582);
nor U12662 (N_12662,N_11948,N_10899);
or U12663 (N_12663,N_11894,N_11933);
nor U12664 (N_12664,N_10061,N_11964);
xnor U12665 (N_12665,N_10232,N_11370);
or U12666 (N_12666,N_10495,N_10386);
xor U12667 (N_12667,N_11565,N_11305);
xnor U12668 (N_12668,N_11250,N_11356);
or U12669 (N_12669,N_11504,N_11262);
and U12670 (N_12670,N_10171,N_11529);
nor U12671 (N_12671,N_10638,N_11554);
xor U12672 (N_12672,N_11402,N_11380);
nor U12673 (N_12673,N_11752,N_11623);
xor U12674 (N_12674,N_11710,N_11474);
and U12675 (N_12675,N_10077,N_10424);
xor U12676 (N_12676,N_11816,N_10266);
nand U12677 (N_12677,N_11441,N_11840);
or U12678 (N_12678,N_10648,N_10352);
or U12679 (N_12679,N_10290,N_11755);
nor U12680 (N_12680,N_10698,N_10808);
nor U12681 (N_12681,N_11694,N_11675);
xor U12682 (N_12682,N_10393,N_11891);
or U12683 (N_12683,N_10218,N_10883);
xor U12684 (N_12684,N_10443,N_10468);
xor U12685 (N_12685,N_10153,N_10730);
or U12686 (N_12686,N_10664,N_11986);
and U12687 (N_12687,N_10426,N_10348);
nand U12688 (N_12688,N_10972,N_10740);
nand U12689 (N_12689,N_11936,N_10273);
and U12690 (N_12690,N_11193,N_10774);
nand U12691 (N_12691,N_11546,N_11867);
or U12692 (N_12692,N_11105,N_10746);
nor U12693 (N_12693,N_11595,N_11383);
nor U12694 (N_12694,N_10689,N_11688);
and U12695 (N_12695,N_11252,N_10927);
xnor U12696 (N_12696,N_11239,N_11925);
nor U12697 (N_12697,N_10794,N_10279);
nand U12698 (N_12698,N_10902,N_11503);
and U12699 (N_12699,N_11125,N_10734);
or U12700 (N_12700,N_10553,N_11829);
and U12701 (N_12701,N_11959,N_11054);
or U12702 (N_12702,N_11790,N_10049);
nand U12703 (N_12703,N_10241,N_11434);
nor U12704 (N_12704,N_11869,N_11489);
nor U12705 (N_12705,N_10137,N_10853);
nor U12706 (N_12706,N_11219,N_11834);
xor U12707 (N_12707,N_11031,N_11057);
xnor U12708 (N_12708,N_11650,N_10892);
or U12709 (N_12709,N_11321,N_10149);
xor U12710 (N_12710,N_10866,N_10342);
and U12711 (N_12711,N_11042,N_11144);
nor U12712 (N_12712,N_11181,N_10869);
nor U12713 (N_12713,N_11841,N_11606);
xor U12714 (N_12714,N_10125,N_10961);
or U12715 (N_12715,N_10498,N_11038);
nor U12716 (N_12716,N_11904,N_11158);
xnor U12717 (N_12717,N_11254,N_10597);
or U12718 (N_12718,N_11879,N_10671);
or U12719 (N_12719,N_11921,N_11428);
nor U12720 (N_12720,N_11293,N_11928);
nor U12721 (N_12721,N_11023,N_10474);
nor U12722 (N_12722,N_10284,N_10974);
nor U12723 (N_12723,N_11365,N_10819);
nand U12724 (N_12724,N_10187,N_10785);
nand U12725 (N_12725,N_11659,N_10564);
xor U12726 (N_12726,N_11517,N_11742);
and U12727 (N_12727,N_10858,N_11408);
xnor U12728 (N_12728,N_10805,N_11849);
nor U12729 (N_12729,N_11243,N_10527);
and U12730 (N_12730,N_10978,N_11541);
xnor U12731 (N_12731,N_10907,N_10539);
nor U12732 (N_12732,N_10060,N_10609);
or U12733 (N_12733,N_10724,N_10011);
or U12734 (N_12734,N_10274,N_11496);
and U12735 (N_12735,N_11437,N_10381);
nand U12736 (N_12736,N_10162,N_10526);
and U12737 (N_12737,N_10630,N_10817);
nor U12738 (N_12738,N_10401,N_10086);
and U12739 (N_12739,N_11228,N_11351);
and U12740 (N_12740,N_11072,N_10613);
or U12741 (N_12741,N_11175,N_10308);
nor U12742 (N_12742,N_10823,N_10780);
and U12743 (N_12743,N_11778,N_11566);
nand U12744 (N_12744,N_10834,N_11372);
and U12745 (N_12745,N_10754,N_11561);
or U12746 (N_12746,N_10128,N_11135);
nor U12747 (N_12747,N_11735,N_11532);
and U12748 (N_12748,N_11950,N_11292);
or U12749 (N_12749,N_11418,N_10683);
xor U12750 (N_12750,N_11505,N_10710);
nor U12751 (N_12751,N_10442,N_11381);
xnor U12752 (N_12752,N_11363,N_10723);
or U12753 (N_12753,N_11258,N_11142);
xnor U12754 (N_12754,N_11369,N_11654);
and U12755 (N_12755,N_10036,N_10779);
or U12756 (N_12756,N_10127,N_11722);
or U12757 (N_12757,N_11683,N_10656);
nor U12758 (N_12758,N_11777,N_11184);
nand U12759 (N_12759,N_10134,N_11833);
nand U12760 (N_12760,N_11364,N_11949);
or U12761 (N_12761,N_11029,N_10940);
nor U12762 (N_12762,N_10572,N_10769);
xor U12763 (N_12763,N_11272,N_10481);
xnor U12764 (N_12764,N_11401,N_11295);
nand U12765 (N_12765,N_11366,N_10259);
and U12766 (N_12766,N_10688,N_11880);
or U12767 (N_12767,N_11847,N_11280);
xnor U12768 (N_12768,N_10488,N_10182);
xnor U12769 (N_12769,N_11132,N_10346);
and U12770 (N_12770,N_10701,N_11530);
or U12771 (N_12771,N_11929,N_10807);
and U12772 (N_12772,N_11926,N_10456);
nor U12773 (N_12773,N_10891,N_10048);
xor U12774 (N_12774,N_10328,N_10075);
nor U12775 (N_12775,N_11572,N_11340);
nand U12776 (N_12776,N_10674,N_11631);
and U12777 (N_12777,N_10658,N_11030);
nor U12778 (N_12778,N_10033,N_11724);
nand U12779 (N_12779,N_11692,N_10112);
nor U12780 (N_12780,N_11211,N_10314);
nor U12781 (N_12781,N_10092,N_10763);
nand U12782 (N_12782,N_11332,N_10811);
nor U12783 (N_12783,N_10161,N_10855);
xor U12784 (N_12784,N_11015,N_11405);
nand U12785 (N_12785,N_11398,N_10343);
or U12786 (N_12786,N_11888,N_11577);
xnor U12787 (N_12787,N_11617,N_10511);
or U12788 (N_12788,N_11646,N_10614);
xor U12789 (N_12789,N_11362,N_10013);
and U12790 (N_12790,N_11788,N_11097);
xnor U12791 (N_12791,N_11131,N_10848);
xnor U12792 (N_12792,N_11695,N_10908);
and U12793 (N_12793,N_11602,N_10212);
nor U12794 (N_12794,N_10200,N_10760);
xor U12795 (N_12795,N_11164,N_10864);
nand U12796 (N_12796,N_11913,N_11575);
nor U12797 (N_12797,N_10655,N_10898);
or U12798 (N_12798,N_10878,N_11179);
nand U12799 (N_12799,N_10026,N_10057);
and U12800 (N_12800,N_11842,N_10660);
nor U12801 (N_12801,N_10164,N_11970);
xnor U12802 (N_12802,N_10646,N_11887);
or U12803 (N_12803,N_11579,N_10140);
nand U12804 (N_12804,N_10703,N_11652);
and U12805 (N_12805,N_11178,N_11610);
and U12806 (N_12806,N_10093,N_10720);
or U12807 (N_12807,N_11516,N_11930);
nor U12808 (N_12808,N_11242,N_11185);
nand U12809 (N_12809,N_11387,N_10476);
and U12810 (N_12810,N_11237,N_10925);
xor U12811 (N_12811,N_11192,N_10761);
nor U12812 (N_12812,N_10410,N_11845);
xor U12813 (N_12813,N_11112,N_10305);
nand U12814 (N_12814,N_11003,N_11745);
nor U12815 (N_12815,N_11821,N_10640);
xnor U12816 (N_12816,N_11872,N_11415);
nor U12817 (N_12817,N_11407,N_11432);
xnor U12818 (N_12818,N_10697,N_10376);
nand U12819 (N_12819,N_11128,N_10296);
xnor U12820 (N_12820,N_10850,N_10191);
or U12821 (N_12821,N_10884,N_10330);
xor U12822 (N_12822,N_11629,N_10912);
nor U12823 (N_12823,N_10827,N_10584);
and U12824 (N_12824,N_10632,N_11510);
xor U12825 (N_12825,N_11786,N_11304);
nand U12826 (N_12826,N_10911,N_11996);
xnor U12827 (N_12827,N_10260,N_11524);
nor U12828 (N_12828,N_11062,N_11567);
or U12829 (N_12829,N_11256,N_10619);
or U12830 (N_12830,N_11992,N_10403);
or U12831 (N_12831,N_11020,N_10307);
xnor U12832 (N_12832,N_10677,N_11826);
or U12833 (N_12833,N_10174,N_11645);
nand U12834 (N_12834,N_10494,N_10110);
and U12835 (N_12835,N_10964,N_11357);
or U12836 (N_12836,N_10388,N_11653);
and U12837 (N_12837,N_11429,N_11980);
nand U12838 (N_12838,N_10482,N_11451);
nor U12839 (N_12839,N_10204,N_10073);
xnor U12840 (N_12840,N_11839,N_10561);
nor U12841 (N_12841,N_10177,N_10350);
xnor U12842 (N_12842,N_11217,N_11043);
or U12843 (N_12843,N_11999,N_11731);
nand U12844 (N_12844,N_10053,N_11528);
nor U12845 (N_12845,N_10550,N_10003);
and U12846 (N_12846,N_10552,N_11176);
or U12847 (N_12847,N_11983,N_10176);
nor U12848 (N_12848,N_11378,N_11622);
or U12849 (N_12849,N_11696,N_11739);
xor U12850 (N_12850,N_10065,N_10524);
xnor U12851 (N_12851,N_11286,N_10299);
nand U12852 (N_12852,N_10933,N_11349);
or U12853 (N_12853,N_11919,N_10108);
nor U12854 (N_12854,N_10588,N_10578);
or U12855 (N_12855,N_10067,N_10982);
or U12856 (N_12856,N_10280,N_11797);
or U12857 (N_12857,N_11981,N_11607);
nand U12858 (N_12858,N_11355,N_11624);
nor U12859 (N_12859,N_11931,N_10886);
or U12860 (N_12860,N_11644,N_11907);
nor U12861 (N_12861,N_10631,N_11711);
or U12862 (N_12862,N_10334,N_11004);
and U12863 (N_12863,N_11457,N_11861);
nor U12864 (N_12864,N_11491,N_11612);
nor U12865 (N_12865,N_10225,N_11781);
and U12866 (N_12866,N_11720,N_11604);
and U12867 (N_12867,N_10958,N_11045);
and U12868 (N_12868,N_11207,N_11548);
nand U12869 (N_12869,N_10256,N_10814);
and U12870 (N_12870,N_11883,N_10043);
xor U12871 (N_12871,N_10178,N_11438);
or U12872 (N_12872,N_11682,N_11350);
or U12873 (N_12873,N_11226,N_11736);
or U12874 (N_12874,N_11947,N_10917);
or U12875 (N_12875,N_10833,N_11594);
and U12876 (N_12876,N_11152,N_11697);
xnor U12877 (N_12877,N_10385,N_10910);
or U12878 (N_12878,N_11551,N_11345);
nor U12879 (N_12879,N_10665,N_11044);
xnor U12880 (N_12880,N_11667,N_11195);
nand U12881 (N_12881,N_10430,N_11319);
nand U12882 (N_12882,N_11537,N_10791);
xnor U12883 (N_12883,N_10981,N_10079);
and U12884 (N_12884,N_10538,N_11480);
and U12885 (N_12885,N_11946,N_10133);
xnor U12886 (N_12886,N_10582,N_10778);
xor U12887 (N_12887,N_10559,N_10713);
and U12888 (N_12888,N_11342,N_10467);
xnor U12889 (N_12889,N_11941,N_10418);
nor U12890 (N_12890,N_10383,N_11182);
and U12891 (N_12891,N_11071,N_10138);
or U12892 (N_12892,N_10900,N_10623);
and U12893 (N_12893,N_11257,N_11317);
xnor U12894 (N_12894,N_10413,N_10019);
xor U12895 (N_12895,N_11375,N_10024);
or U12896 (N_12896,N_11648,N_11222);
nor U12897 (N_12897,N_11110,N_10267);
and U12898 (N_12898,N_11799,N_10118);
nor U12899 (N_12899,N_11456,N_10612);
and U12900 (N_12900,N_11758,N_10265);
or U12901 (N_12901,N_10159,N_10846);
and U12902 (N_12902,N_11059,N_10686);
nand U12903 (N_12903,N_10904,N_11091);
xor U12904 (N_12904,N_10324,N_10544);
nor U12905 (N_12905,N_10862,N_10795);
xor U12906 (N_12906,N_10510,N_10861);
nor U12907 (N_12907,N_11493,N_10622);
xnor U12908 (N_12908,N_10782,N_10996);
and U12909 (N_12909,N_11705,N_10502);
and U12910 (N_12910,N_10729,N_11327);
or U12911 (N_12911,N_11425,N_10822);
and U12912 (N_12912,N_10793,N_10402);
nor U12913 (N_12913,N_11495,N_11205);
nor U12914 (N_12914,N_10250,N_11074);
xnor U12915 (N_12915,N_11717,N_10428);
nand U12916 (N_12916,N_10337,N_10025);
nor U12917 (N_12917,N_10213,N_11477);
xor U12918 (N_12918,N_11874,N_10534);
nor U12919 (N_12919,N_10606,N_11520);
nor U12920 (N_12920,N_10081,N_11241);
nor U12921 (N_12921,N_11718,N_10968);
nor U12922 (N_12922,N_11039,N_10644);
nand U12923 (N_12923,N_10618,N_11230);
and U12924 (N_12924,N_11213,N_11290);
or U12925 (N_12925,N_11827,N_10522);
or U12926 (N_12926,N_11170,N_10725);
nor U12927 (N_12927,N_10366,N_11966);
nor U12928 (N_12928,N_10235,N_11865);
xor U12929 (N_12929,N_10179,N_10058);
nor U12930 (N_12930,N_10988,N_10726);
nor U12931 (N_12931,N_11588,N_10325);
and U12932 (N_12932,N_10104,N_11672);
and U12933 (N_12933,N_10221,N_11792);
xor U12934 (N_12934,N_11310,N_11715);
or U12935 (N_12935,N_11190,N_10373);
xnor U12936 (N_12936,N_11884,N_11637);
nand U12937 (N_12937,N_10208,N_10229);
and U12938 (N_12938,N_11898,N_11942);
and U12939 (N_12939,N_11535,N_10962);
nor U12940 (N_12940,N_10590,N_11462);
nor U12941 (N_12941,N_11868,N_11093);
nand U12942 (N_12942,N_10199,N_11431);
nor U12943 (N_12943,N_10479,N_11574);
nand U12944 (N_12944,N_11277,N_10540);
xnor U12945 (N_12945,N_11669,N_10708);
nor U12946 (N_12946,N_10455,N_10490);
xor U12947 (N_12947,N_10124,N_11268);
xnor U12948 (N_12948,N_11298,N_10317);
nand U12949 (N_12949,N_11109,N_11830);
or U12950 (N_12950,N_10223,N_10090);
nand U12951 (N_12951,N_11488,N_11460);
xnor U12952 (N_12952,N_11917,N_11932);
or U12953 (N_12953,N_11005,N_10909);
or U12954 (N_12954,N_10998,N_11464);
xnor U12955 (N_12955,N_11956,N_11278);
nor U12956 (N_12956,N_11915,N_10732);
nand U12957 (N_12957,N_11163,N_10000);
nand U12958 (N_12958,N_10603,N_10738);
nand U12959 (N_12959,N_10203,N_11444);
nand U12960 (N_12960,N_11945,N_11468);
or U12961 (N_12961,N_11373,N_10716);
and U12962 (N_12962,N_11553,N_10427);
xor U12963 (N_12963,N_10103,N_11126);
xnor U12964 (N_12964,N_10107,N_10704);
or U12965 (N_12965,N_11633,N_11903);
or U12966 (N_12966,N_10359,N_11214);
nor U12967 (N_12967,N_10957,N_10624);
or U12968 (N_12968,N_11406,N_10651);
or U12969 (N_12969,N_11076,N_11598);
or U12970 (N_12970,N_10087,N_11118);
nand U12971 (N_12971,N_10806,N_11523);
nor U12972 (N_12972,N_10775,N_10536);
and U12973 (N_12973,N_10889,N_10854);
or U12974 (N_12974,N_10963,N_10167);
nor U12975 (N_12975,N_10327,N_10083);
nor U12976 (N_12976,N_11776,N_10135);
nand U12977 (N_12977,N_10639,N_10185);
and U12978 (N_12978,N_11399,N_11944);
nand U12979 (N_12979,N_10398,N_10051);
or U12980 (N_12980,N_10487,N_11315);
xor U12981 (N_12981,N_10423,N_11384);
or U12982 (N_12982,N_11684,N_11655);
xnor U12983 (N_12983,N_11962,N_11772);
or U12984 (N_12984,N_10937,N_11453);
nor U12985 (N_12985,N_11360,N_10106);
nor U12986 (N_12986,N_10506,N_10165);
xor U12987 (N_12987,N_11209,N_11615);
nand U12988 (N_12988,N_11019,N_11923);
nor U12989 (N_12989,N_10210,N_11025);
or U12990 (N_12990,N_11070,N_11279);
or U12991 (N_12991,N_10954,N_10906);
and U12992 (N_12992,N_11571,N_11263);
nand U12993 (N_12993,N_11218,N_10718);
nand U12994 (N_12994,N_11393,N_10895);
and U12995 (N_12995,N_11161,N_11569);
xor U12996 (N_12996,N_10292,N_11299);
xor U12997 (N_12997,N_11825,N_10695);
and U12998 (N_12998,N_11166,N_11619);
nand U12999 (N_12999,N_10151,N_10173);
xnor U13000 (N_13000,N_10429,N_11599);
or U13001 (N_13001,N_11911,N_11416);
xor U13002 (N_13002,N_11377,N_10548);
nand U13003 (N_13003,N_11889,N_11513);
nor U13004 (N_13004,N_10117,N_11627);
xnor U13005 (N_13005,N_11727,N_10079);
nand U13006 (N_13006,N_10726,N_11161);
or U13007 (N_13007,N_11955,N_10124);
or U13008 (N_13008,N_11681,N_10316);
xor U13009 (N_13009,N_10818,N_10829);
nand U13010 (N_13010,N_11450,N_11808);
xnor U13011 (N_13011,N_11895,N_11273);
nand U13012 (N_13012,N_11163,N_10276);
nor U13013 (N_13013,N_11766,N_11193);
xor U13014 (N_13014,N_11898,N_10245);
and U13015 (N_13015,N_10393,N_11553);
and U13016 (N_13016,N_11899,N_10955);
nor U13017 (N_13017,N_10293,N_11288);
or U13018 (N_13018,N_11663,N_10179);
nor U13019 (N_13019,N_10063,N_11143);
nand U13020 (N_13020,N_11931,N_11524);
and U13021 (N_13021,N_10850,N_11068);
nand U13022 (N_13022,N_10520,N_11349);
nor U13023 (N_13023,N_10780,N_10179);
xnor U13024 (N_13024,N_10731,N_11663);
nand U13025 (N_13025,N_10190,N_11611);
xor U13026 (N_13026,N_10632,N_10670);
xor U13027 (N_13027,N_10584,N_10836);
xnor U13028 (N_13028,N_10905,N_10761);
or U13029 (N_13029,N_10516,N_10594);
nor U13030 (N_13030,N_11742,N_10480);
xor U13031 (N_13031,N_10998,N_10402);
and U13032 (N_13032,N_10870,N_10799);
or U13033 (N_13033,N_11311,N_10862);
or U13034 (N_13034,N_10129,N_10561);
and U13035 (N_13035,N_10097,N_10057);
and U13036 (N_13036,N_11948,N_11045);
nand U13037 (N_13037,N_11459,N_10377);
xnor U13038 (N_13038,N_11319,N_11329);
nand U13039 (N_13039,N_11021,N_10731);
nor U13040 (N_13040,N_10233,N_11160);
nand U13041 (N_13041,N_11076,N_10540);
and U13042 (N_13042,N_11351,N_10024);
nor U13043 (N_13043,N_11055,N_10940);
nor U13044 (N_13044,N_10778,N_11568);
xnor U13045 (N_13045,N_11986,N_10936);
nor U13046 (N_13046,N_10478,N_10933);
xor U13047 (N_13047,N_11444,N_10967);
nand U13048 (N_13048,N_10864,N_11708);
nor U13049 (N_13049,N_11268,N_11412);
nand U13050 (N_13050,N_11964,N_10984);
xnor U13051 (N_13051,N_11968,N_11119);
or U13052 (N_13052,N_10201,N_10307);
nor U13053 (N_13053,N_10936,N_11538);
nand U13054 (N_13054,N_11112,N_11297);
and U13055 (N_13055,N_10720,N_10319);
xnor U13056 (N_13056,N_10946,N_10578);
xor U13057 (N_13057,N_11413,N_11668);
xnor U13058 (N_13058,N_11698,N_11520);
nand U13059 (N_13059,N_11419,N_10486);
xnor U13060 (N_13060,N_10030,N_11261);
nand U13061 (N_13061,N_10700,N_11638);
nor U13062 (N_13062,N_11359,N_11058);
nor U13063 (N_13063,N_10456,N_11296);
nand U13064 (N_13064,N_11101,N_11546);
or U13065 (N_13065,N_11443,N_10088);
xor U13066 (N_13066,N_10141,N_10876);
nor U13067 (N_13067,N_10921,N_11277);
and U13068 (N_13068,N_11987,N_10075);
or U13069 (N_13069,N_10123,N_10551);
and U13070 (N_13070,N_10486,N_10218);
and U13071 (N_13071,N_10198,N_11399);
nand U13072 (N_13072,N_11380,N_11561);
xor U13073 (N_13073,N_11610,N_10029);
nand U13074 (N_13074,N_10007,N_10776);
nand U13075 (N_13075,N_10848,N_11016);
nand U13076 (N_13076,N_10909,N_11691);
or U13077 (N_13077,N_10652,N_10925);
xnor U13078 (N_13078,N_10039,N_10013);
and U13079 (N_13079,N_11491,N_11020);
xor U13080 (N_13080,N_11295,N_10249);
nor U13081 (N_13081,N_11021,N_11623);
xnor U13082 (N_13082,N_10294,N_11855);
or U13083 (N_13083,N_11882,N_10792);
nor U13084 (N_13084,N_11965,N_10638);
nor U13085 (N_13085,N_10091,N_11837);
xor U13086 (N_13086,N_10703,N_10083);
and U13087 (N_13087,N_11528,N_10853);
nand U13088 (N_13088,N_11913,N_10202);
nand U13089 (N_13089,N_11539,N_11860);
nor U13090 (N_13090,N_10377,N_11924);
or U13091 (N_13091,N_10050,N_11313);
xnor U13092 (N_13092,N_10284,N_11638);
nor U13093 (N_13093,N_10932,N_11133);
or U13094 (N_13094,N_10792,N_11714);
or U13095 (N_13095,N_10364,N_10871);
xnor U13096 (N_13096,N_11826,N_11004);
xor U13097 (N_13097,N_11554,N_10814);
nor U13098 (N_13098,N_10765,N_10511);
nor U13099 (N_13099,N_10072,N_10418);
nor U13100 (N_13100,N_10484,N_10068);
nand U13101 (N_13101,N_10052,N_10997);
nand U13102 (N_13102,N_11511,N_10138);
nand U13103 (N_13103,N_10246,N_10035);
nand U13104 (N_13104,N_11569,N_11687);
and U13105 (N_13105,N_11166,N_11713);
xor U13106 (N_13106,N_11127,N_10818);
xnor U13107 (N_13107,N_11174,N_10991);
nor U13108 (N_13108,N_10569,N_11780);
nand U13109 (N_13109,N_11090,N_11288);
or U13110 (N_13110,N_10059,N_11446);
xor U13111 (N_13111,N_10130,N_11761);
nand U13112 (N_13112,N_11582,N_10174);
nand U13113 (N_13113,N_11052,N_11094);
and U13114 (N_13114,N_10745,N_11534);
nor U13115 (N_13115,N_11922,N_10127);
and U13116 (N_13116,N_10904,N_10918);
xor U13117 (N_13117,N_10511,N_11550);
xnor U13118 (N_13118,N_11189,N_11688);
or U13119 (N_13119,N_11676,N_10531);
xor U13120 (N_13120,N_10099,N_11267);
xnor U13121 (N_13121,N_11940,N_10467);
xnor U13122 (N_13122,N_11539,N_11068);
xor U13123 (N_13123,N_10086,N_10250);
and U13124 (N_13124,N_10671,N_11180);
and U13125 (N_13125,N_11575,N_10342);
xnor U13126 (N_13126,N_10496,N_11182);
and U13127 (N_13127,N_11003,N_11418);
or U13128 (N_13128,N_10455,N_10259);
nand U13129 (N_13129,N_11537,N_11160);
nor U13130 (N_13130,N_11552,N_10885);
xor U13131 (N_13131,N_11483,N_10306);
or U13132 (N_13132,N_11640,N_10703);
nor U13133 (N_13133,N_11647,N_10914);
nand U13134 (N_13134,N_11305,N_10871);
xor U13135 (N_13135,N_11383,N_11875);
xor U13136 (N_13136,N_11102,N_11785);
or U13137 (N_13137,N_11678,N_10373);
nor U13138 (N_13138,N_11308,N_11208);
nor U13139 (N_13139,N_10280,N_10680);
nor U13140 (N_13140,N_11381,N_10592);
and U13141 (N_13141,N_10222,N_11327);
and U13142 (N_13142,N_10940,N_10857);
xor U13143 (N_13143,N_10192,N_10264);
xor U13144 (N_13144,N_11790,N_10441);
xor U13145 (N_13145,N_10734,N_11108);
and U13146 (N_13146,N_11423,N_11792);
and U13147 (N_13147,N_10486,N_11037);
and U13148 (N_13148,N_11952,N_11094);
nand U13149 (N_13149,N_11766,N_10007);
xnor U13150 (N_13150,N_10125,N_10902);
nand U13151 (N_13151,N_10773,N_10500);
nand U13152 (N_13152,N_10667,N_11600);
xor U13153 (N_13153,N_11611,N_11787);
and U13154 (N_13154,N_10921,N_10864);
nor U13155 (N_13155,N_11105,N_11804);
xnor U13156 (N_13156,N_10173,N_11662);
xor U13157 (N_13157,N_10861,N_10476);
nor U13158 (N_13158,N_10948,N_11550);
nand U13159 (N_13159,N_10073,N_10833);
or U13160 (N_13160,N_10789,N_11140);
nand U13161 (N_13161,N_10959,N_10527);
or U13162 (N_13162,N_10640,N_10429);
or U13163 (N_13163,N_11059,N_10114);
xnor U13164 (N_13164,N_10191,N_10671);
and U13165 (N_13165,N_11691,N_11436);
xor U13166 (N_13166,N_10336,N_10912);
nand U13167 (N_13167,N_10190,N_11849);
nor U13168 (N_13168,N_11126,N_11995);
xnor U13169 (N_13169,N_11975,N_10431);
or U13170 (N_13170,N_11672,N_11192);
or U13171 (N_13171,N_11902,N_10245);
xor U13172 (N_13172,N_11424,N_11800);
and U13173 (N_13173,N_11122,N_11322);
and U13174 (N_13174,N_10402,N_11268);
and U13175 (N_13175,N_10119,N_11165);
or U13176 (N_13176,N_11477,N_11780);
or U13177 (N_13177,N_10923,N_11337);
nand U13178 (N_13178,N_11227,N_10941);
or U13179 (N_13179,N_11793,N_10202);
nor U13180 (N_13180,N_11816,N_11311);
nor U13181 (N_13181,N_11324,N_10317);
and U13182 (N_13182,N_11409,N_10959);
or U13183 (N_13183,N_10919,N_10519);
nand U13184 (N_13184,N_10535,N_10285);
xor U13185 (N_13185,N_10406,N_11134);
nor U13186 (N_13186,N_10596,N_11940);
or U13187 (N_13187,N_11628,N_11135);
xnor U13188 (N_13188,N_11360,N_11664);
nand U13189 (N_13189,N_11813,N_11307);
nand U13190 (N_13190,N_11666,N_11574);
or U13191 (N_13191,N_10499,N_11696);
or U13192 (N_13192,N_10525,N_10195);
nor U13193 (N_13193,N_10400,N_11334);
nand U13194 (N_13194,N_11390,N_11035);
nor U13195 (N_13195,N_10220,N_11508);
xnor U13196 (N_13196,N_10222,N_11050);
xor U13197 (N_13197,N_10975,N_11801);
and U13198 (N_13198,N_11016,N_10504);
and U13199 (N_13199,N_11931,N_11681);
and U13200 (N_13200,N_11887,N_10280);
xor U13201 (N_13201,N_11909,N_11168);
and U13202 (N_13202,N_10065,N_10069);
nand U13203 (N_13203,N_10933,N_10905);
xnor U13204 (N_13204,N_10506,N_11712);
nor U13205 (N_13205,N_10523,N_10922);
and U13206 (N_13206,N_11811,N_11152);
or U13207 (N_13207,N_11448,N_10815);
nor U13208 (N_13208,N_10126,N_11756);
xor U13209 (N_13209,N_10914,N_11113);
and U13210 (N_13210,N_11704,N_10357);
nor U13211 (N_13211,N_10087,N_11023);
and U13212 (N_13212,N_10614,N_10064);
xor U13213 (N_13213,N_10382,N_10919);
nand U13214 (N_13214,N_11206,N_11138);
nor U13215 (N_13215,N_11531,N_11348);
nor U13216 (N_13216,N_11322,N_11965);
and U13217 (N_13217,N_10364,N_10105);
and U13218 (N_13218,N_11498,N_11135);
nor U13219 (N_13219,N_10409,N_10148);
or U13220 (N_13220,N_11528,N_11899);
and U13221 (N_13221,N_10734,N_10540);
or U13222 (N_13222,N_11809,N_11461);
xor U13223 (N_13223,N_10085,N_10992);
nor U13224 (N_13224,N_11950,N_11530);
nand U13225 (N_13225,N_11242,N_10023);
or U13226 (N_13226,N_10858,N_11985);
or U13227 (N_13227,N_10457,N_11333);
nand U13228 (N_13228,N_10056,N_11339);
or U13229 (N_13229,N_10745,N_11314);
nand U13230 (N_13230,N_11798,N_10491);
nor U13231 (N_13231,N_10433,N_10188);
nor U13232 (N_13232,N_10587,N_10661);
and U13233 (N_13233,N_10105,N_10218);
xnor U13234 (N_13234,N_11961,N_11602);
nor U13235 (N_13235,N_10955,N_11541);
nand U13236 (N_13236,N_10137,N_11639);
xnor U13237 (N_13237,N_11305,N_11223);
nand U13238 (N_13238,N_10979,N_11734);
nand U13239 (N_13239,N_11433,N_11387);
nor U13240 (N_13240,N_11547,N_11970);
xnor U13241 (N_13241,N_11021,N_10360);
nor U13242 (N_13242,N_11524,N_10020);
and U13243 (N_13243,N_10424,N_10023);
xor U13244 (N_13244,N_11291,N_11321);
or U13245 (N_13245,N_11749,N_10457);
and U13246 (N_13246,N_10474,N_10773);
nor U13247 (N_13247,N_10255,N_10384);
or U13248 (N_13248,N_11065,N_10813);
or U13249 (N_13249,N_11402,N_10024);
or U13250 (N_13250,N_11293,N_11186);
nand U13251 (N_13251,N_10139,N_10359);
or U13252 (N_13252,N_11331,N_10986);
or U13253 (N_13253,N_11826,N_11162);
nand U13254 (N_13254,N_10971,N_10736);
or U13255 (N_13255,N_10945,N_11146);
or U13256 (N_13256,N_11885,N_11907);
and U13257 (N_13257,N_10548,N_10003);
nand U13258 (N_13258,N_11270,N_10794);
xnor U13259 (N_13259,N_10772,N_11588);
nand U13260 (N_13260,N_10929,N_10817);
nand U13261 (N_13261,N_11794,N_11682);
or U13262 (N_13262,N_10520,N_10484);
nor U13263 (N_13263,N_10186,N_11593);
xnor U13264 (N_13264,N_11252,N_10758);
and U13265 (N_13265,N_11172,N_11364);
nor U13266 (N_13266,N_10586,N_10274);
and U13267 (N_13267,N_10859,N_10436);
nand U13268 (N_13268,N_10258,N_10025);
and U13269 (N_13269,N_10542,N_11460);
xnor U13270 (N_13270,N_10076,N_11335);
or U13271 (N_13271,N_11782,N_11070);
or U13272 (N_13272,N_11558,N_11597);
and U13273 (N_13273,N_10109,N_10838);
and U13274 (N_13274,N_11554,N_11975);
nand U13275 (N_13275,N_10273,N_11926);
xor U13276 (N_13276,N_11913,N_10752);
or U13277 (N_13277,N_10088,N_11362);
or U13278 (N_13278,N_10020,N_10078);
and U13279 (N_13279,N_11439,N_10279);
nand U13280 (N_13280,N_10714,N_10290);
nor U13281 (N_13281,N_10170,N_10002);
xor U13282 (N_13282,N_11231,N_10408);
and U13283 (N_13283,N_11722,N_11109);
and U13284 (N_13284,N_11155,N_11663);
or U13285 (N_13285,N_11625,N_10185);
nand U13286 (N_13286,N_11122,N_10593);
xor U13287 (N_13287,N_10653,N_11070);
nor U13288 (N_13288,N_11254,N_10040);
nand U13289 (N_13289,N_10066,N_10040);
and U13290 (N_13290,N_11954,N_10153);
xnor U13291 (N_13291,N_10714,N_10835);
xor U13292 (N_13292,N_11869,N_11768);
nand U13293 (N_13293,N_11215,N_10810);
nor U13294 (N_13294,N_11384,N_11122);
and U13295 (N_13295,N_10441,N_11310);
nor U13296 (N_13296,N_11812,N_10528);
nor U13297 (N_13297,N_11975,N_10676);
or U13298 (N_13298,N_11275,N_10526);
or U13299 (N_13299,N_10516,N_10938);
and U13300 (N_13300,N_11257,N_10934);
xor U13301 (N_13301,N_11326,N_11146);
nor U13302 (N_13302,N_10345,N_10792);
and U13303 (N_13303,N_10750,N_10757);
or U13304 (N_13304,N_11366,N_11122);
xor U13305 (N_13305,N_10032,N_11414);
nand U13306 (N_13306,N_10592,N_11288);
xor U13307 (N_13307,N_11938,N_11688);
nor U13308 (N_13308,N_11483,N_11395);
and U13309 (N_13309,N_11144,N_10752);
nor U13310 (N_13310,N_10581,N_11243);
nor U13311 (N_13311,N_11016,N_11705);
xnor U13312 (N_13312,N_10682,N_10457);
or U13313 (N_13313,N_10370,N_10407);
or U13314 (N_13314,N_10777,N_11628);
nor U13315 (N_13315,N_10732,N_10470);
nor U13316 (N_13316,N_11962,N_11851);
and U13317 (N_13317,N_10546,N_10265);
xor U13318 (N_13318,N_10456,N_11675);
nor U13319 (N_13319,N_11765,N_10738);
nand U13320 (N_13320,N_11212,N_11829);
xor U13321 (N_13321,N_11889,N_11405);
xor U13322 (N_13322,N_10805,N_10225);
and U13323 (N_13323,N_10592,N_10715);
nor U13324 (N_13324,N_11209,N_11796);
nand U13325 (N_13325,N_10061,N_10027);
nand U13326 (N_13326,N_10961,N_10453);
and U13327 (N_13327,N_11290,N_11454);
xor U13328 (N_13328,N_11483,N_10197);
or U13329 (N_13329,N_10660,N_10525);
nor U13330 (N_13330,N_11057,N_11323);
nand U13331 (N_13331,N_10378,N_11433);
or U13332 (N_13332,N_10459,N_11527);
and U13333 (N_13333,N_10197,N_11125);
nand U13334 (N_13334,N_10392,N_10615);
or U13335 (N_13335,N_11250,N_11264);
or U13336 (N_13336,N_11908,N_11694);
nor U13337 (N_13337,N_10127,N_11147);
and U13338 (N_13338,N_11409,N_10119);
xnor U13339 (N_13339,N_10150,N_11490);
nor U13340 (N_13340,N_11679,N_11715);
and U13341 (N_13341,N_10523,N_10292);
and U13342 (N_13342,N_11068,N_10660);
xor U13343 (N_13343,N_11387,N_11853);
nor U13344 (N_13344,N_11090,N_11467);
or U13345 (N_13345,N_11306,N_10428);
and U13346 (N_13346,N_10200,N_10587);
nand U13347 (N_13347,N_11268,N_11494);
nor U13348 (N_13348,N_11686,N_11447);
xor U13349 (N_13349,N_11407,N_11295);
nor U13350 (N_13350,N_11582,N_10627);
nand U13351 (N_13351,N_11662,N_11400);
nor U13352 (N_13352,N_10774,N_10288);
and U13353 (N_13353,N_11948,N_11866);
or U13354 (N_13354,N_11305,N_11005);
or U13355 (N_13355,N_10068,N_11862);
nand U13356 (N_13356,N_10340,N_10102);
xor U13357 (N_13357,N_10282,N_10908);
nand U13358 (N_13358,N_11046,N_10368);
nand U13359 (N_13359,N_11037,N_10589);
nor U13360 (N_13360,N_10070,N_10301);
or U13361 (N_13361,N_10576,N_11733);
xnor U13362 (N_13362,N_11411,N_11264);
or U13363 (N_13363,N_10065,N_11532);
nor U13364 (N_13364,N_11950,N_11239);
nand U13365 (N_13365,N_10595,N_11833);
or U13366 (N_13366,N_11971,N_11848);
nor U13367 (N_13367,N_11197,N_11256);
xor U13368 (N_13368,N_10326,N_10664);
nor U13369 (N_13369,N_10548,N_10315);
or U13370 (N_13370,N_10290,N_10148);
and U13371 (N_13371,N_10672,N_10413);
nor U13372 (N_13372,N_10542,N_10167);
nor U13373 (N_13373,N_11154,N_11653);
xor U13374 (N_13374,N_11466,N_11033);
nand U13375 (N_13375,N_11311,N_11354);
or U13376 (N_13376,N_10791,N_11344);
and U13377 (N_13377,N_10478,N_11470);
and U13378 (N_13378,N_11399,N_11159);
xnor U13379 (N_13379,N_11017,N_11056);
nand U13380 (N_13380,N_11202,N_10798);
and U13381 (N_13381,N_10810,N_11771);
or U13382 (N_13382,N_11464,N_10726);
xor U13383 (N_13383,N_10884,N_11738);
or U13384 (N_13384,N_10828,N_10647);
and U13385 (N_13385,N_11167,N_10751);
nand U13386 (N_13386,N_10246,N_10552);
or U13387 (N_13387,N_11521,N_10226);
nand U13388 (N_13388,N_10047,N_10550);
or U13389 (N_13389,N_11719,N_11319);
nand U13390 (N_13390,N_11830,N_11313);
xor U13391 (N_13391,N_10735,N_11001);
xnor U13392 (N_13392,N_10148,N_11746);
and U13393 (N_13393,N_11047,N_11122);
nor U13394 (N_13394,N_11603,N_11079);
xor U13395 (N_13395,N_10159,N_11033);
nand U13396 (N_13396,N_11767,N_10802);
and U13397 (N_13397,N_11324,N_11415);
nor U13398 (N_13398,N_10211,N_10870);
and U13399 (N_13399,N_11607,N_10176);
nand U13400 (N_13400,N_11545,N_11828);
nand U13401 (N_13401,N_10778,N_10298);
nor U13402 (N_13402,N_11783,N_10394);
xor U13403 (N_13403,N_10933,N_10415);
nor U13404 (N_13404,N_10623,N_11876);
and U13405 (N_13405,N_10321,N_10799);
and U13406 (N_13406,N_11630,N_11437);
or U13407 (N_13407,N_11748,N_10030);
or U13408 (N_13408,N_11634,N_11959);
nor U13409 (N_13409,N_10392,N_11253);
or U13410 (N_13410,N_10387,N_10862);
and U13411 (N_13411,N_11003,N_11347);
nor U13412 (N_13412,N_11265,N_11967);
xor U13413 (N_13413,N_11644,N_10442);
or U13414 (N_13414,N_10083,N_10596);
nor U13415 (N_13415,N_11138,N_10067);
nor U13416 (N_13416,N_10324,N_11801);
and U13417 (N_13417,N_11671,N_11820);
nor U13418 (N_13418,N_11170,N_10314);
or U13419 (N_13419,N_11898,N_11116);
xnor U13420 (N_13420,N_11931,N_11866);
xnor U13421 (N_13421,N_11181,N_10015);
nand U13422 (N_13422,N_10762,N_10731);
or U13423 (N_13423,N_11759,N_11638);
and U13424 (N_13424,N_11521,N_11057);
or U13425 (N_13425,N_11482,N_10844);
nor U13426 (N_13426,N_10073,N_10197);
nand U13427 (N_13427,N_11336,N_10260);
and U13428 (N_13428,N_10370,N_11060);
or U13429 (N_13429,N_11098,N_10925);
or U13430 (N_13430,N_11902,N_11797);
nor U13431 (N_13431,N_11405,N_10959);
or U13432 (N_13432,N_10779,N_10718);
and U13433 (N_13433,N_11350,N_11253);
and U13434 (N_13434,N_11199,N_11273);
and U13435 (N_13435,N_11775,N_10069);
nor U13436 (N_13436,N_11670,N_10649);
and U13437 (N_13437,N_11304,N_11053);
nand U13438 (N_13438,N_11393,N_10272);
and U13439 (N_13439,N_10379,N_10153);
xor U13440 (N_13440,N_10022,N_10673);
nand U13441 (N_13441,N_10093,N_11382);
xnor U13442 (N_13442,N_10363,N_10444);
or U13443 (N_13443,N_10583,N_10697);
nand U13444 (N_13444,N_10638,N_10463);
xnor U13445 (N_13445,N_11935,N_10839);
xnor U13446 (N_13446,N_11456,N_10802);
xnor U13447 (N_13447,N_11859,N_11636);
nand U13448 (N_13448,N_11887,N_11681);
nand U13449 (N_13449,N_10553,N_10166);
xnor U13450 (N_13450,N_10165,N_10891);
nand U13451 (N_13451,N_11914,N_11584);
nor U13452 (N_13452,N_10498,N_11493);
nor U13453 (N_13453,N_11718,N_10880);
or U13454 (N_13454,N_11906,N_11627);
nand U13455 (N_13455,N_10105,N_10775);
and U13456 (N_13456,N_10525,N_11293);
and U13457 (N_13457,N_10561,N_10788);
nand U13458 (N_13458,N_10702,N_10159);
or U13459 (N_13459,N_10678,N_10816);
and U13460 (N_13460,N_11605,N_11127);
or U13461 (N_13461,N_10139,N_10179);
xnor U13462 (N_13462,N_10560,N_11014);
or U13463 (N_13463,N_10996,N_11116);
xor U13464 (N_13464,N_10783,N_10412);
xnor U13465 (N_13465,N_11800,N_10512);
and U13466 (N_13466,N_10373,N_11458);
nand U13467 (N_13467,N_10327,N_10639);
or U13468 (N_13468,N_10446,N_11867);
or U13469 (N_13469,N_11349,N_10826);
and U13470 (N_13470,N_10259,N_11735);
xnor U13471 (N_13471,N_10025,N_11936);
nand U13472 (N_13472,N_11829,N_10168);
nor U13473 (N_13473,N_11040,N_11786);
or U13474 (N_13474,N_10269,N_11593);
nor U13475 (N_13475,N_10930,N_11188);
nand U13476 (N_13476,N_10815,N_11948);
nand U13477 (N_13477,N_11948,N_10787);
nor U13478 (N_13478,N_10092,N_11841);
xor U13479 (N_13479,N_10641,N_10827);
nand U13480 (N_13480,N_10587,N_10808);
or U13481 (N_13481,N_11496,N_11988);
and U13482 (N_13482,N_11371,N_11458);
or U13483 (N_13483,N_11976,N_10520);
nor U13484 (N_13484,N_10590,N_10532);
nor U13485 (N_13485,N_10615,N_11813);
nor U13486 (N_13486,N_11735,N_10569);
xor U13487 (N_13487,N_11899,N_10264);
or U13488 (N_13488,N_10121,N_11885);
nor U13489 (N_13489,N_10179,N_11542);
or U13490 (N_13490,N_10028,N_11932);
xor U13491 (N_13491,N_10330,N_10301);
xor U13492 (N_13492,N_11614,N_10827);
nor U13493 (N_13493,N_10869,N_10182);
nand U13494 (N_13494,N_10623,N_11260);
nand U13495 (N_13495,N_11369,N_11823);
and U13496 (N_13496,N_10421,N_10459);
xnor U13497 (N_13497,N_10926,N_10630);
and U13498 (N_13498,N_11388,N_11520);
nand U13499 (N_13499,N_10690,N_10543);
or U13500 (N_13500,N_11552,N_11780);
nor U13501 (N_13501,N_11229,N_10595);
nand U13502 (N_13502,N_10431,N_10726);
xor U13503 (N_13503,N_11141,N_10493);
or U13504 (N_13504,N_10791,N_11171);
and U13505 (N_13505,N_10877,N_11859);
or U13506 (N_13506,N_10722,N_11306);
or U13507 (N_13507,N_11639,N_10061);
xor U13508 (N_13508,N_11363,N_11022);
nand U13509 (N_13509,N_11378,N_11432);
or U13510 (N_13510,N_11619,N_10833);
xnor U13511 (N_13511,N_11086,N_10260);
nor U13512 (N_13512,N_11215,N_10260);
or U13513 (N_13513,N_10763,N_11720);
nand U13514 (N_13514,N_10752,N_10411);
nor U13515 (N_13515,N_10944,N_11979);
and U13516 (N_13516,N_10171,N_11877);
and U13517 (N_13517,N_10912,N_11110);
or U13518 (N_13518,N_10683,N_11343);
and U13519 (N_13519,N_10364,N_10546);
xnor U13520 (N_13520,N_10634,N_10147);
nand U13521 (N_13521,N_11235,N_10341);
and U13522 (N_13522,N_11243,N_11892);
and U13523 (N_13523,N_11842,N_10149);
nor U13524 (N_13524,N_10106,N_10531);
or U13525 (N_13525,N_11021,N_11015);
xor U13526 (N_13526,N_10296,N_10623);
nor U13527 (N_13527,N_10244,N_11915);
xnor U13528 (N_13528,N_11363,N_10915);
or U13529 (N_13529,N_11384,N_10940);
nand U13530 (N_13530,N_10814,N_11056);
or U13531 (N_13531,N_11829,N_11013);
xor U13532 (N_13532,N_11105,N_11866);
nand U13533 (N_13533,N_10307,N_11151);
or U13534 (N_13534,N_11163,N_11421);
nand U13535 (N_13535,N_11897,N_11325);
and U13536 (N_13536,N_10567,N_10176);
and U13537 (N_13537,N_10880,N_10952);
and U13538 (N_13538,N_10136,N_10472);
and U13539 (N_13539,N_11754,N_10265);
or U13540 (N_13540,N_10468,N_10234);
xnor U13541 (N_13541,N_11262,N_10399);
and U13542 (N_13542,N_10283,N_11221);
nand U13543 (N_13543,N_11766,N_10372);
nor U13544 (N_13544,N_10587,N_11957);
and U13545 (N_13545,N_10134,N_11741);
or U13546 (N_13546,N_11930,N_11652);
nor U13547 (N_13547,N_11966,N_10722);
and U13548 (N_13548,N_10053,N_10184);
nor U13549 (N_13549,N_11022,N_10578);
and U13550 (N_13550,N_11190,N_11746);
nand U13551 (N_13551,N_11650,N_10894);
nand U13552 (N_13552,N_11697,N_11472);
xnor U13553 (N_13553,N_10687,N_11588);
and U13554 (N_13554,N_10535,N_10203);
nand U13555 (N_13555,N_10139,N_11201);
and U13556 (N_13556,N_10937,N_10670);
nand U13557 (N_13557,N_10095,N_11601);
or U13558 (N_13558,N_10148,N_11071);
nand U13559 (N_13559,N_11933,N_11762);
and U13560 (N_13560,N_11802,N_10771);
nand U13561 (N_13561,N_11965,N_11873);
nor U13562 (N_13562,N_10802,N_11165);
or U13563 (N_13563,N_11060,N_11291);
nand U13564 (N_13564,N_11269,N_11737);
and U13565 (N_13565,N_10677,N_11819);
xnor U13566 (N_13566,N_10306,N_10412);
or U13567 (N_13567,N_11602,N_10184);
nor U13568 (N_13568,N_11147,N_10272);
nor U13569 (N_13569,N_11515,N_10671);
xor U13570 (N_13570,N_11297,N_11158);
or U13571 (N_13571,N_10646,N_11961);
xnor U13572 (N_13572,N_11515,N_11187);
xnor U13573 (N_13573,N_10102,N_10890);
xor U13574 (N_13574,N_11647,N_11887);
nand U13575 (N_13575,N_10354,N_10374);
and U13576 (N_13576,N_10228,N_11594);
or U13577 (N_13577,N_11284,N_11653);
nor U13578 (N_13578,N_10072,N_10053);
and U13579 (N_13579,N_11089,N_10439);
and U13580 (N_13580,N_10305,N_11267);
and U13581 (N_13581,N_11386,N_10223);
or U13582 (N_13582,N_11724,N_10446);
nor U13583 (N_13583,N_11162,N_11373);
nand U13584 (N_13584,N_11081,N_10753);
nand U13585 (N_13585,N_11582,N_11870);
or U13586 (N_13586,N_10890,N_10399);
nor U13587 (N_13587,N_10759,N_11395);
nor U13588 (N_13588,N_11092,N_11074);
xnor U13589 (N_13589,N_10667,N_11868);
and U13590 (N_13590,N_10535,N_11183);
or U13591 (N_13591,N_10043,N_10687);
nand U13592 (N_13592,N_10822,N_10092);
and U13593 (N_13593,N_10249,N_11139);
and U13594 (N_13594,N_10529,N_11822);
or U13595 (N_13595,N_11495,N_10966);
or U13596 (N_13596,N_11420,N_11044);
xor U13597 (N_13597,N_11153,N_11652);
nand U13598 (N_13598,N_10417,N_10052);
nor U13599 (N_13599,N_11050,N_11233);
nand U13600 (N_13600,N_10375,N_10958);
nor U13601 (N_13601,N_11056,N_11810);
nor U13602 (N_13602,N_11751,N_10228);
nor U13603 (N_13603,N_11334,N_11701);
nand U13604 (N_13604,N_11217,N_10023);
nand U13605 (N_13605,N_11491,N_11475);
nand U13606 (N_13606,N_11859,N_10965);
xor U13607 (N_13607,N_11651,N_10153);
or U13608 (N_13608,N_11045,N_11539);
nand U13609 (N_13609,N_10127,N_10981);
xor U13610 (N_13610,N_11043,N_11440);
nand U13611 (N_13611,N_10944,N_11888);
nand U13612 (N_13612,N_10342,N_10478);
xor U13613 (N_13613,N_11773,N_11296);
and U13614 (N_13614,N_11902,N_11187);
or U13615 (N_13615,N_10845,N_11812);
xor U13616 (N_13616,N_10445,N_11914);
nor U13617 (N_13617,N_10688,N_10338);
or U13618 (N_13618,N_10347,N_10987);
or U13619 (N_13619,N_10654,N_11948);
nor U13620 (N_13620,N_11968,N_11317);
nand U13621 (N_13621,N_10313,N_10707);
and U13622 (N_13622,N_10019,N_11212);
xnor U13623 (N_13623,N_10019,N_10317);
nor U13624 (N_13624,N_11269,N_10872);
xor U13625 (N_13625,N_11691,N_10279);
nor U13626 (N_13626,N_11869,N_11895);
nand U13627 (N_13627,N_11855,N_10785);
nor U13628 (N_13628,N_10289,N_10865);
nand U13629 (N_13629,N_10422,N_11131);
xor U13630 (N_13630,N_10127,N_10722);
nand U13631 (N_13631,N_11845,N_10727);
xor U13632 (N_13632,N_10370,N_11077);
nor U13633 (N_13633,N_10724,N_11731);
nand U13634 (N_13634,N_10274,N_11752);
nor U13635 (N_13635,N_11541,N_11716);
nor U13636 (N_13636,N_11793,N_11941);
nor U13637 (N_13637,N_11098,N_11936);
nand U13638 (N_13638,N_11903,N_10000);
or U13639 (N_13639,N_11456,N_11727);
nor U13640 (N_13640,N_11413,N_10614);
or U13641 (N_13641,N_11590,N_11593);
nor U13642 (N_13642,N_11614,N_11291);
and U13643 (N_13643,N_10917,N_11194);
nor U13644 (N_13644,N_11073,N_10370);
and U13645 (N_13645,N_11396,N_11011);
nor U13646 (N_13646,N_10163,N_10324);
and U13647 (N_13647,N_10543,N_11243);
nor U13648 (N_13648,N_10380,N_10093);
nand U13649 (N_13649,N_10928,N_11557);
nand U13650 (N_13650,N_10503,N_10927);
and U13651 (N_13651,N_10389,N_11447);
and U13652 (N_13652,N_11338,N_11102);
nor U13653 (N_13653,N_11109,N_11917);
nand U13654 (N_13654,N_10144,N_11022);
and U13655 (N_13655,N_11731,N_10107);
xor U13656 (N_13656,N_10934,N_10454);
or U13657 (N_13657,N_11816,N_10070);
nand U13658 (N_13658,N_10294,N_11447);
nor U13659 (N_13659,N_11886,N_11080);
xor U13660 (N_13660,N_11665,N_10801);
nor U13661 (N_13661,N_11365,N_11063);
xnor U13662 (N_13662,N_10986,N_11787);
or U13663 (N_13663,N_11232,N_11377);
nor U13664 (N_13664,N_10798,N_11086);
nand U13665 (N_13665,N_11126,N_10577);
xnor U13666 (N_13666,N_11581,N_11303);
or U13667 (N_13667,N_11032,N_11166);
nand U13668 (N_13668,N_11932,N_10829);
xnor U13669 (N_13669,N_10281,N_11810);
xnor U13670 (N_13670,N_11838,N_10456);
and U13671 (N_13671,N_11820,N_10673);
nor U13672 (N_13672,N_11747,N_11331);
nor U13673 (N_13673,N_10657,N_10384);
nor U13674 (N_13674,N_11091,N_11706);
or U13675 (N_13675,N_11437,N_11490);
or U13676 (N_13676,N_11867,N_10517);
nor U13677 (N_13677,N_11879,N_10079);
and U13678 (N_13678,N_11211,N_11915);
nor U13679 (N_13679,N_10576,N_11318);
nand U13680 (N_13680,N_10202,N_10926);
nand U13681 (N_13681,N_11028,N_10518);
xnor U13682 (N_13682,N_10194,N_10953);
xnor U13683 (N_13683,N_11998,N_11430);
nor U13684 (N_13684,N_11944,N_10017);
or U13685 (N_13685,N_11465,N_10337);
nand U13686 (N_13686,N_10576,N_11551);
and U13687 (N_13687,N_11229,N_10738);
or U13688 (N_13688,N_10756,N_11139);
xnor U13689 (N_13689,N_10808,N_10192);
nor U13690 (N_13690,N_10420,N_10961);
nand U13691 (N_13691,N_11724,N_10274);
xor U13692 (N_13692,N_10886,N_10361);
nand U13693 (N_13693,N_10168,N_10842);
nand U13694 (N_13694,N_10872,N_11883);
nor U13695 (N_13695,N_11649,N_10851);
xor U13696 (N_13696,N_11256,N_11015);
xnor U13697 (N_13697,N_11051,N_10950);
nor U13698 (N_13698,N_10537,N_11164);
nor U13699 (N_13699,N_10751,N_11632);
nand U13700 (N_13700,N_10328,N_11858);
xnor U13701 (N_13701,N_10927,N_11343);
and U13702 (N_13702,N_11180,N_10039);
and U13703 (N_13703,N_11127,N_10847);
nand U13704 (N_13704,N_10514,N_10721);
nand U13705 (N_13705,N_10563,N_11591);
xnor U13706 (N_13706,N_10944,N_10319);
or U13707 (N_13707,N_10404,N_10255);
nand U13708 (N_13708,N_10609,N_11931);
or U13709 (N_13709,N_11037,N_11576);
nor U13710 (N_13710,N_10501,N_10705);
or U13711 (N_13711,N_10146,N_11545);
and U13712 (N_13712,N_10407,N_11838);
xor U13713 (N_13713,N_11750,N_11931);
nand U13714 (N_13714,N_10909,N_11009);
nor U13715 (N_13715,N_11696,N_10880);
or U13716 (N_13716,N_10057,N_11378);
xor U13717 (N_13717,N_10406,N_10577);
and U13718 (N_13718,N_10960,N_11309);
nand U13719 (N_13719,N_10979,N_10081);
or U13720 (N_13720,N_11030,N_10550);
and U13721 (N_13721,N_11335,N_11478);
xnor U13722 (N_13722,N_10392,N_10756);
and U13723 (N_13723,N_10797,N_11630);
nor U13724 (N_13724,N_11639,N_10568);
xor U13725 (N_13725,N_11767,N_11247);
xor U13726 (N_13726,N_10735,N_11201);
nand U13727 (N_13727,N_10632,N_11392);
or U13728 (N_13728,N_11108,N_10658);
xnor U13729 (N_13729,N_10734,N_11750);
or U13730 (N_13730,N_10975,N_10862);
nor U13731 (N_13731,N_11723,N_10722);
xor U13732 (N_13732,N_11624,N_11647);
nor U13733 (N_13733,N_11558,N_10145);
xor U13734 (N_13734,N_11748,N_10029);
xnor U13735 (N_13735,N_11105,N_10757);
nor U13736 (N_13736,N_11319,N_11542);
nand U13737 (N_13737,N_11485,N_11412);
or U13738 (N_13738,N_10346,N_10715);
nor U13739 (N_13739,N_10393,N_11203);
and U13740 (N_13740,N_11218,N_10269);
nand U13741 (N_13741,N_10798,N_10506);
and U13742 (N_13742,N_10246,N_11302);
nand U13743 (N_13743,N_11419,N_10621);
nand U13744 (N_13744,N_10204,N_10916);
xor U13745 (N_13745,N_11049,N_11383);
nand U13746 (N_13746,N_11325,N_10594);
nor U13747 (N_13747,N_10665,N_11473);
and U13748 (N_13748,N_10842,N_11854);
xor U13749 (N_13749,N_10983,N_11642);
or U13750 (N_13750,N_10021,N_11664);
nor U13751 (N_13751,N_11171,N_11714);
nand U13752 (N_13752,N_10120,N_11305);
nor U13753 (N_13753,N_11513,N_11858);
xor U13754 (N_13754,N_11025,N_10587);
nand U13755 (N_13755,N_11656,N_10731);
or U13756 (N_13756,N_11587,N_10045);
xnor U13757 (N_13757,N_11449,N_10472);
xnor U13758 (N_13758,N_10996,N_10806);
nor U13759 (N_13759,N_11783,N_11156);
nand U13760 (N_13760,N_10120,N_11580);
xor U13761 (N_13761,N_11891,N_10309);
or U13762 (N_13762,N_10289,N_10137);
or U13763 (N_13763,N_11423,N_11450);
and U13764 (N_13764,N_10599,N_10078);
or U13765 (N_13765,N_11088,N_11251);
nand U13766 (N_13766,N_11475,N_10934);
xnor U13767 (N_13767,N_10048,N_11512);
xor U13768 (N_13768,N_10733,N_10262);
nand U13769 (N_13769,N_11651,N_10966);
nor U13770 (N_13770,N_10063,N_11210);
nand U13771 (N_13771,N_10046,N_10705);
nand U13772 (N_13772,N_10142,N_11176);
or U13773 (N_13773,N_11313,N_10289);
nor U13774 (N_13774,N_10046,N_10515);
xnor U13775 (N_13775,N_10014,N_10255);
or U13776 (N_13776,N_11142,N_11290);
xnor U13777 (N_13777,N_11821,N_11548);
xor U13778 (N_13778,N_10589,N_10449);
nand U13779 (N_13779,N_11582,N_10778);
or U13780 (N_13780,N_11213,N_10241);
and U13781 (N_13781,N_11891,N_10839);
or U13782 (N_13782,N_10959,N_11968);
or U13783 (N_13783,N_11744,N_10902);
and U13784 (N_13784,N_10732,N_10158);
nand U13785 (N_13785,N_11422,N_11332);
nor U13786 (N_13786,N_10451,N_10076);
and U13787 (N_13787,N_10029,N_11903);
xnor U13788 (N_13788,N_11745,N_10275);
or U13789 (N_13789,N_11915,N_10965);
and U13790 (N_13790,N_10826,N_10818);
or U13791 (N_13791,N_11210,N_10457);
nor U13792 (N_13792,N_10834,N_11652);
or U13793 (N_13793,N_11714,N_10713);
nor U13794 (N_13794,N_10014,N_10052);
nor U13795 (N_13795,N_10301,N_11985);
and U13796 (N_13796,N_10973,N_10000);
or U13797 (N_13797,N_11796,N_10869);
nand U13798 (N_13798,N_11553,N_11080);
nand U13799 (N_13799,N_10520,N_11229);
or U13800 (N_13800,N_11943,N_11649);
nor U13801 (N_13801,N_11225,N_10481);
xor U13802 (N_13802,N_11162,N_11030);
xor U13803 (N_13803,N_11732,N_10590);
nand U13804 (N_13804,N_11780,N_11351);
and U13805 (N_13805,N_11417,N_11075);
and U13806 (N_13806,N_11144,N_10144);
and U13807 (N_13807,N_10288,N_10942);
and U13808 (N_13808,N_10577,N_11705);
nand U13809 (N_13809,N_11441,N_10099);
nand U13810 (N_13810,N_10847,N_10420);
nand U13811 (N_13811,N_10775,N_11945);
and U13812 (N_13812,N_11339,N_10367);
and U13813 (N_13813,N_11702,N_10657);
nor U13814 (N_13814,N_10265,N_10821);
nand U13815 (N_13815,N_10381,N_11894);
nor U13816 (N_13816,N_11825,N_11917);
nor U13817 (N_13817,N_11304,N_11232);
nand U13818 (N_13818,N_10644,N_11379);
nand U13819 (N_13819,N_10574,N_10173);
or U13820 (N_13820,N_10356,N_11872);
xor U13821 (N_13821,N_11213,N_10278);
xnor U13822 (N_13822,N_10726,N_11486);
nor U13823 (N_13823,N_10576,N_10397);
or U13824 (N_13824,N_10317,N_11624);
or U13825 (N_13825,N_11868,N_11548);
nor U13826 (N_13826,N_10083,N_10915);
and U13827 (N_13827,N_10007,N_11945);
and U13828 (N_13828,N_11461,N_11345);
and U13829 (N_13829,N_11524,N_10078);
and U13830 (N_13830,N_10848,N_11652);
nor U13831 (N_13831,N_11723,N_10673);
or U13832 (N_13832,N_10221,N_10744);
nand U13833 (N_13833,N_10364,N_10477);
nor U13834 (N_13834,N_10909,N_10525);
xnor U13835 (N_13835,N_10200,N_10253);
and U13836 (N_13836,N_10074,N_11100);
or U13837 (N_13837,N_11806,N_11426);
nor U13838 (N_13838,N_10307,N_10356);
or U13839 (N_13839,N_10475,N_11852);
and U13840 (N_13840,N_10696,N_10932);
nor U13841 (N_13841,N_11064,N_11737);
nor U13842 (N_13842,N_11554,N_11555);
and U13843 (N_13843,N_11080,N_10218);
and U13844 (N_13844,N_10152,N_10085);
xnor U13845 (N_13845,N_10133,N_11123);
xor U13846 (N_13846,N_11235,N_10679);
nor U13847 (N_13847,N_10481,N_10266);
xnor U13848 (N_13848,N_11438,N_11058);
nand U13849 (N_13849,N_11871,N_10454);
or U13850 (N_13850,N_10888,N_10987);
xor U13851 (N_13851,N_10126,N_11768);
nand U13852 (N_13852,N_10781,N_10047);
nor U13853 (N_13853,N_11579,N_10095);
nor U13854 (N_13854,N_11256,N_11342);
and U13855 (N_13855,N_11949,N_10969);
and U13856 (N_13856,N_11916,N_10447);
nor U13857 (N_13857,N_11773,N_11585);
nand U13858 (N_13858,N_10906,N_11840);
or U13859 (N_13859,N_10617,N_10380);
and U13860 (N_13860,N_11568,N_10232);
nand U13861 (N_13861,N_10553,N_10629);
xor U13862 (N_13862,N_11221,N_11047);
nor U13863 (N_13863,N_10930,N_10530);
nor U13864 (N_13864,N_10618,N_10200);
or U13865 (N_13865,N_11847,N_11419);
and U13866 (N_13866,N_10860,N_11684);
or U13867 (N_13867,N_10771,N_10449);
or U13868 (N_13868,N_11596,N_10573);
nand U13869 (N_13869,N_10750,N_11237);
nand U13870 (N_13870,N_10786,N_11051);
and U13871 (N_13871,N_10821,N_11797);
or U13872 (N_13872,N_10659,N_11568);
and U13873 (N_13873,N_11262,N_10908);
xnor U13874 (N_13874,N_10928,N_11062);
nand U13875 (N_13875,N_11240,N_11039);
and U13876 (N_13876,N_10209,N_11674);
or U13877 (N_13877,N_10770,N_11055);
xnor U13878 (N_13878,N_10678,N_10569);
nor U13879 (N_13879,N_11328,N_10386);
or U13880 (N_13880,N_11631,N_11815);
xnor U13881 (N_13881,N_10089,N_11945);
nor U13882 (N_13882,N_11416,N_10164);
nor U13883 (N_13883,N_10123,N_11664);
or U13884 (N_13884,N_11154,N_10735);
or U13885 (N_13885,N_11334,N_11234);
nand U13886 (N_13886,N_11570,N_11937);
nand U13887 (N_13887,N_11653,N_10045);
nand U13888 (N_13888,N_11107,N_10554);
nor U13889 (N_13889,N_11820,N_10991);
and U13890 (N_13890,N_11416,N_10085);
nand U13891 (N_13891,N_10336,N_11166);
and U13892 (N_13892,N_10220,N_11756);
xnor U13893 (N_13893,N_11793,N_10201);
nor U13894 (N_13894,N_11430,N_10609);
nor U13895 (N_13895,N_11616,N_11732);
and U13896 (N_13896,N_11514,N_11348);
nor U13897 (N_13897,N_10756,N_10508);
nand U13898 (N_13898,N_11903,N_11139);
or U13899 (N_13899,N_10018,N_11040);
or U13900 (N_13900,N_11433,N_10629);
xor U13901 (N_13901,N_10817,N_11442);
and U13902 (N_13902,N_11036,N_10134);
and U13903 (N_13903,N_10207,N_10987);
xnor U13904 (N_13904,N_10178,N_10843);
xnor U13905 (N_13905,N_10227,N_10010);
and U13906 (N_13906,N_10187,N_11024);
nor U13907 (N_13907,N_10089,N_10336);
or U13908 (N_13908,N_10599,N_10362);
xor U13909 (N_13909,N_10320,N_10686);
nor U13910 (N_13910,N_11169,N_11153);
or U13911 (N_13911,N_11797,N_11539);
nor U13912 (N_13912,N_10007,N_11299);
or U13913 (N_13913,N_11655,N_11633);
and U13914 (N_13914,N_11216,N_11846);
and U13915 (N_13915,N_10939,N_10478);
nor U13916 (N_13916,N_11835,N_10118);
xor U13917 (N_13917,N_11328,N_11102);
nand U13918 (N_13918,N_11282,N_11529);
xnor U13919 (N_13919,N_10959,N_10098);
or U13920 (N_13920,N_10393,N_11689);
xor U13921 (N_13921,N_11808,N_10785);
or U13922 (N_13922,N_10653,N_10847);
xnor U13923 (N_13923,N_10084,N_11901);
and U13924 (N_13924,N_10912,N_10483);
and U13925 (N_13925,N_10070,N_10650);
and U13926 (N_13926,N_11133,N_10899);
nand U13927 (N_13927,N_11889,N_10809);
nor U13928 (N_13928,N_10924,N_10614);
and U13929 (N_13929,N_10013,N_10653);
xor U13930 (N_13930,N_11832,N_10477);
and U13931 (N_13931,N_11329,N_11246);
xnor U13932 (N_13932,N_11380,N_11412);
xor U13933 (N_13933,N_10723,N_10904);
or U13934 (N_13934,N_11211,N_11649);
nand U13935 (N_13935,N_11772,N_11614);
nor U13936 (N_13936,N_11810,N_10733);
nor U13937 (N_13937,N_11580,N_10414);
and U13938 (N_13938,N_10979,N_11474);
or U13939 (N_13939,N_11992,N_10483);
nor U13940 (N_13940,N_11745,N_11506);
and U13941 (N_13941,N_11857,N_11552);
xor U13942 (N_13942,N_11919,N_10268);
nor U13943 (N_13943,N_11797,N_11213);
xnor U13944 (N_13944,N_11306,N_10140);
nand U13945 (N_13945,N_10303,N_11348);
nand U13946 (N_13946,N_11670,N_11800);
nor U13947 (N_13947,N_10963,N_11555);
nor U13948 (N_13948,N_11435,N_10331);
nand U13949 (N_13949,N_10933,N_11071);
nor U13950 (N_13950,N_10719,N_11863);
or U13951 (N_13951,N_11353,N_11000);
or U13952 (N_13952,N_11148,N_10174);
or U13953 (N_13953,N_10793,N_11920);
and U13954 (N_13954,N_10046,N_10909);
nand U13955 (N_13955,N_11689,N_11342);
nor U13956 (N_13956,N_11441,N_10676);
or U13957 (N_13957,N_10359,N_11243);
nand U13958 (N_13958,N_11461,N_11377);
and U13959 (N_13959,N_11212,N_10977);
nand U13960 (N_13960,N_10945,N_10642);
or U13961 (N_13961,N_11278,N_11503);
xor U13962 (N_13962,N_11648,N_11328);
nand U13963 (N_13963,N_10844,N_11047);
nand U13964 (N_13964,N_10168,N_10490);
nand U13965 (N_13965,N_10370,N_11491);
nand U13966 (N_13966,N_10301,N_10635);
or U13967 (N_13967,N_10872,N_10146);
xor U13968 (N_13968,N_11425,N_11614);
nand U13969 (N_13969,N_10499,N_10803);
and U13970 (N_13970,N_11928,N_11963);
nor U13971 (N_13971,N_11749,N_11292);
and U13972 (N_13972,N_11887,N_10010);
nor U13973 (N_13973,N_10176,N_10139);
and U13974 (N_13974,N_11014,N_11321);
nor U13975 (N_13975,N_10231,N_11733);
xor U13976 (N_13976,N_11192,N_10069);
nand U13977 (N_13977,N_11136,N_11545);
and U13978 (N_13978,N_11014,N_11392);
and U13979 (N_13979,N_11022,N_10753);
and U13980 (N_13980,N_11585,N_10990);
or U13981 (N_13981,N_11763,N_11355);
nand U13982 (N_13982,N_11358,N_10833);
and U13983 (N_13983,N_11846,N_11406);
nor U13984 (N_13984,N_11335,N_10762);
or U13985 (N_13985,N_11225,N_10007);
nor U13986 (N_13986,N_10931,N_11515);
or U13987 (N_13987,N_10192,N_11270);
or U13988 (N_13988,N_11400,N_10308);
and U13989 (N_13989,N_10852,N_10972);
and U13990 (N_13990,N_11711,N_10404);
xnor U13991 (N_13991,N_11400,N_11831);
nor U13992 (N_13992,N_11681,N_11384);
and U13993 (N_13993,N_10943,N_11005);
and U13994 (N_13994,N_10616,N_11578);
and U13995 (N_13995,N_11381,N_10892);
or U13996 (N_13996,N_10822,N_11773);
nor U13997 (N_13997,N_11439,N_10246);
or U13998 (N_13998,N_11864,N_10383);
and U13999 (N_13999,N_10978,N_10141);
nand U14000 (N_14000,N_13677,N_12095);
nor U14001 (N_14001,N_13541,N_13657);
nand U14002 (N_14002,N_13321,N_12917);
and U14003 (N_14003,N_12425,N_12962);
or U14004 (N_14004,N_13522,N_13899);
and U14005 (N_14005,N_13653,N_12499);
xnor U14006 (N_14006,N_13027,N_12163);
or U14007 (N_14007,N_12831,N_13111);
nor U14008 (N_14008,N_12070,N_12302);
or U14009 (N_14009,N_13010,N_12398);
nor U14010 (N_14010,N_12493,N_12053);
and U14011 (N_14011,N_13096,N_13146);
nor U14012 (N_14012,N_13727,N_12538);
and U14013 (N_14013,N_12675,N_13021);
and U14014 (N_14014,N_13118,N_12607);
xor U14015 (N_14015,N_12769,N_12122);
nor U14016 (N_14016,N_13125,N_12423);
and U14017 (N_14017,N_13767,N_12435);
xor U14018 (N_14018,N_12983,N_12746);
nor U14019 (N_14019,N_13614,N_12691);
nor U14020 (N_14020,N_12217,N_13768);
nand U14021 (N_14021,N_13559,N_13849);
nor U14022 (N_14022,N_13317,N_13120);
or U14023 (N_14023,N_12145,N_13031);
nor U14024 (N_14024,N_13943,N_13372);
nand U14025 (N_14025,N_13500,N_12484);
xor U14026 (N_14026,N_12738,N_12574);
xnor U14027 (N_14027,N_13515,N_13831);
xor U14028 (N_14028,N_13718,N_12380);
xnor U14029 (N_14029,N_12043,N_12376);
nand U14030 (N_14030,N_13877,N_12830);
and U14031 (N_14031,N_13085,N_13762);
xor U14032 (N_14032,N_13544,N_12035);
and U14033 (N_14033,N_13624,N_13475);
nor U14034 (N_14034,N_12033,N_13458);
nor U14035 (N_14035,N_12149,N_12552);
nor U14036 (N_14036,N_12878,N_13946);
nor U14037 (N_14037,N_12566,N_12848);
nand U14038 (N_14038,N_13088,N_13092);
xor U14039 (N_14039,N_12890,N_12846);
nand U14040 (N_14040,N_12599,N_12268);
xor U14041 (N_14041,N_12120,N_12176);
nor U14042 (N_14042,N_12925,N_13628);
nor U14043 (N_14043,N_13290,N_12190);
and U14044 (N_14044,N_12926,N_13870);
and U14045 (N_14045,N_13952,N_12107);
nand U14046 (N_14046,N_12580,N_12375);
or U14047 (N_14047,N_12845,N_13533);
or U14048 (N_14048,N_12100,N_13399);
nor U14049 (N_14049,N_13776,N_12565);
or U14050 (N_14050,N_12515,N_13525);
nor U14051 (N_14051,N_13929,N_13385);
xnor U14052 (N_14052,N_13045,N_12781);
nor U14053 (N_14053,N_13959,N_12361);
or U14054 (N_14054,N_13467,N_13143);
or U14055 (N_14055,N_12803,N_12736);
nor U14056 (N_14056,N_12147,N_13422);
and U14057 (N_14057,N_12224,N_12821);
or U14058 (N_14058,N_13220,N_13038);
xnor U14059 (N_14059,N_12312,N_13410);
nor U14060 (N_14060,N_12577,N_13023);
nor U14061 (N_14061,N_12218,N_13856);
or U14062 (N_14062,N_12490,N_12478);
or U14063 (N_14063,N_12052,N_12152);
and U14064 (N_14064,N_12175,N_13574);
nand U14065 (N_14065,N_12753,N_12004);
nor U14066 (N_14066,N_13961,N_12920);
and U14067 (N_14067,N_12382,N_12928);
and U14068 (N_14068,N_13479,N_13578);
and U14069 (N_14069,N_12256,N_13030);
or U14070 (N_14070,N_12245,N_12048);
nor U14071 (N_14071,N_13466,N_12936);
nand U14072 (N_14072,N_13642,N_13145);
nand U14073 (N_14073,N_13015,N_13556);
nor U14074 (N_14074,N_12481,N_13606);
or U14075 (N_14075,N_13006,N_13409);
or U14076 (N_14076,N_13491,N_13552);
or U14077 (N_14077,N_13345,N_12286);
and U14078 (N_14078,N_12270,N_12628);
or U14079 (N_14079,N_13095,N_12165);
nor U14080 (N_14080,N_13549,N_12167);
and U14081 (N_14081,N_13867,N_13369);
nand U14082 (N_14082,N_13602,N_13885);
nor U14083 (N_14083,N_13881,N_12192);
or U14084 (N_14084,N_12404,N_12251);
or U14085 (N_14085,N_12014,N_13262);
nand U14086 (N_14086,N_12174,N_12386);
or U14087 (N_14087,N_12600,N_12989);
xnor U14088 (N_14088,N_12862,N_13570);
nand U14089 (N_14089,N_13197,N_12057);
and U14090 (N_14090,N_13836,N_12324);
nor U14091 (N_14091,N_12916,N_12437);
xnor U14092 (N_14092,N_12111,N_12209);
xor U14093 (N_14093,N_13189,N_13065);
and U14094 (N_14094,N_13802,N_12416);
and U14095 (N_14095,N_12329,N_12693);
nor U14096 (N_14096,N_12258,N_12353);
or U14097 (N_14097,N_13381,N_12702);
xnor U14098 (N_14098,N_12887,N_12685);
nor U14099 (N_14099,N_12207,N_12308);
or U14100 (N_14100,N_12318,N_13748);
nand U14101 (N_14101,N_12912,N_12009);
and U14102 (N_14102,N_12899,N_12266);
or U14103 (N_14103,N_12334,N_12332);
and U14104 (N_14104,N_12443,N_12118);
nor U14105 (N_14105,N_13608,N_12602);
and U14106 (N_14106,N_13577,N_12992);
xnor U14107 (N_14107,N_13966,N_12520);
or U14108 (N_14108,N_13744,N_13244);
xnor U14109 (N_14109,N_12452,N_13872);
xnor U14110 (N_14110,N_12188,N_12724);
nand U14111 (N_14111,N_13136,N_13584);
or U14112 (N_14112,N_13984,N_13322);
xor U14113 (N_14113,N_13432,N_13108);
nand U14114 (N_14114,N_13873,N_12798);
xor U14115 (N_14115,N_12045,N_12841);
or U14116 (N_14116,N_12428,N_13518);
or U14117 (N_14117,N_13237,N_12123);
xnor U14118 (N_14118,N_12875,N_13086);
nor U14119 (N_14119,N_12979,N_12264);
or U14120 (N_14120,N_12792,N_12480);
nor U14121 (N_14121,N_12117,N_12840);
or U14122 (N_14122,N_12473,N_13889);
nor U14123 (N_14123,N_13816,N_13383);
xor U14124 (N_14124,N_12470,N_12720);
or U14125 (N_14125,N_12299,N_13560);
or U14126 (N_14126,N_13427,N_12756);
nor U14127 (N_14127,N_13115,N_13182);
nand U14128 (N_14128,N_12072,N_12856);
and U14129 (N_14129,N_12189,N_12692);
nor U14130 (N_14130,N_13306,N_12106);
nor U14131 (N_14131,N_12179,N_13282);
or U14132 (N_14132,N_13405,N_13772);
or U14133 (N_14133,N_12390,N_13723);
nand U14134 (N_14134,N_13168,N_12153);
nand U14135 (N_14135,N_12988,N_12140);
nand U14136 (N_14136,N_12460,N_12968);
or U14137 (N_14137,N_12146,N_13913);
nor U14138 (N_14138,N_13489,N_13105);
or U14139 (N_14139,N_13785,N_13914);
or U14140 (N_14140,N_13598,N_13530);
or U14141 (N_14141,N_12465,N_13271);
nand U14142 (N_14142,N_13411,N_13490);
nor U14143 (N_14143,N_13535,N_12468);
nor U14144 (N_14144,N_13621,N_12960);
and U14145 (N_14145,N_12085,N_12378);
or U14146 (N_14146,N_13415,N_13974);
nand U14147 (N_14147,N_12414,N_13364);
nor U14148 (N_14148,N_13078,N_13194);
nor U14149 (N_14149,N_12557,N_12415);
nand U14150 (N_14150,N_13887,N_13007);
and U14151 (N_14151,N_12825,N_12389);
xnor U14152 (N_14152,N_12688,N_13298);
and U14153 (N_14153,N_12281,N_12248);
nand U14154 (N_14154,N_12737,N_12502);
nor U14155 (N_14155,N_12952,N_12313);
nand U14156 (N_14156,N_12171,N_13452);
nand U14157 (N_14157,N_12168,N_13353);
nand U14158 (N_14158,N_12942,N_13547);
nand U14159 (N_14159,N_12016,N_13763);
or U14160 (N_14160,N_13663,N_12818);
nand U14161 (N_14161,N_13033,N_12496);
and U14162 (N_14162,N_13536,N_12008);
xor U14163 (N_14163,N_12653,N_12665);
nand U14164 (N_14164,N_13198,N_13729);
nand U14165 (N_14165,N_13299,N_12026);
nor U14166 (N_14166,N_13694,N_12674);
and U14167 (N_14167,N_12901,N_13215);
nor U14168 (N_14168,N_12497,N_13580);
nor U14169 (N_14169,N_13854,N_13796);
xnor U14170 (N_14170,N_13991,N_13810);
or U14171 (N_14171,N_12214,N_12835);
or U14172 (N_14172,N_12352,N_12886);
or U14173 (N_14173,N_12158,N_13679);
nor U14174 (N_14174,N_12037,N_13423);
nor U14175 (N_14175,N_13397,N_12402);
nand U14176 (N_14176,N_13609,N_12625);
and U14177 (N_14177,N_13706,N_13403);
nand U14178 (N_14178,N_13797,N_12569);
nand U14179 (N_14179,N_12613,N_12283);
xnor U14180 (N_14180,N_12729,N_13281);
and U14181 (N_14181,N_13869,N_13823);
nor U14182 (N_14182,N_13435,N_12802);
xor U14183 (N_14183,N_12529,N_12780);
nor U14184 (N_14184,N_12159,N_13993);
xnor U14185 (N_14185,N_13235,N_13428);
nor U14186 (N_14186,N_12477,N_12278);
and U14187 (N_14187,N_13840,N_13922);
xor U14188 (N_14188,N_12131,N_12227);
xor U14189 (N_14189,N_13018,N_13070);
nor U14190 (N_14190,N_12485,N_12896);
or U14191 (N_14191,N_12592,N_13496);
nand U14192 (N_14192,N_13184,N_12754);
nand U14193 (N_14193,N_12424,N_13738);
nand U14194 (N_14194,N_13789,N_12967);
or U14195 (N_14195,N_12943,N_13592);
nor U14196 (N_14196,N_13732,N_13890);
and U14197 (N_14197,N_12377,N_12865);
or U14198 (N_14198,N_12110,N_12526);
and U14199 (N_14199,N_13293,N_12432);
and U14200 (N_14200,N_13342,N_12407);
xnor U14201 (N_14201,N_13319,N_13268);
or U14202 (N_14202,N_12647,N_13457);
nand U14203 (N_14203,N_13291,N_12621);
nand U14204 (N_14204,N_12451,N_13004);
and U14205 (N_14205,N_13002,N_12020);
xnor U14206 (N_14206,N_13465,N_13450);
nor U14207 (N_14207,N_13080,N_13682);
nor U14208 (N_14208,N_13819,N_13223);
nor U14209 (N_14209,N_12205,N_13186);
nor U14210 (N_14210,N_13148,N_12860);
xor U14211 (N_14211,N_13178,N_12002);
nand U14212 (N_14212,N_13527,N_13071);
or U14213 (N_14213,N_12805,N_12196);
xor U14214 (N_14214,N_12273,N_12114);
nand U14215 (N_14215,N_13431,N_12635);
nor U14216 (N_14216,N_12986,N_13062);
nor U14217 (N_14217,N_12543,N_12459);
nand U14218 (N_14218,N_13040,N_12046);
nor U14219 (N_14219,N_13066,N_12819);
xnor U14220 (N_14220,N_13177,N_13000);
nor U14221 (N_14221,N_13107,N_13554);
nor U14222 (N_14222,N_12454,N_13703);
nor U14223 (N_14223,N_12202,N_13637);
xnor U14224 (N_14224,N_13528,N_13339);
xor U14225 (N_14225,N_12689,N_13671);
xnor U14226 (N_14226,N_13907,N_13855);
nor U14227 (N_14227,N_13736,N_13356);
or U14228 (N_14228,N_12981,N_12065);
xor U14229 (N_14229,N_12271,N_12610);
xnor U14230 (N_14230,N_13859,N_13257);
nor U14231 (N_14231,N_13905,N_12582);
or U14232 (N_14232,N_12588,N_12813);
or U14233 (N_14233,N_12984,N_12243);
nand U14234 (N_14234,N_13393,N_12034);
nor U14235 (N_14235,N_13585,N_13822);
nand U14236 (N_14236,N_12839,N_13206);
nand U14237 (N_14237,N_13927,N_13246);
and U14238 (N_14238,N_13801,N_13950);
or U14239 (N_14239,N_13507,N_13099);
xor U14240 (N_14240,N_13942,N_12127);
or U14241 (N_14241,N_13800,N_12093);
xor U14242 (N_14242,N_13935,N_13516);
and U14243 (N_14243,N_13582,N_12327);
nand U14244 (N_14244,N_12551,N_13692);
nor U14245 (N_14245,N_12121,N_12115);
nor U14246 (N_14246,N_13534,N_12698);
xnor U14247 (N_14247,N_12346,N_13627);
nor U14248 (N_14248,N_13140,N_13478);
and U14249 (N_14249,N_13986,N_12556);
xor U14250 (N_14250,N_12779,N_13894);
nor U14251 (N_14251,N_12368,N_13448);
nor U14252 (N_14252,N_12649,N_12479);
nor U14253 (N_14253,N_12973,N_13312);
or U14254 (N_14254,N_13531,N_12799);
xnor U14255 (N_14255,N_12269,N_13999);
xnor U14256 (N_14256,N_13586,N_13688);
xor U14257 (N_14257,N_12006,N_12410);
and U14258 (N_14258,N_12527,N_12314);
xor U14259 (N_14259,N_13416,N_13611);
or U14260 (N_14260,N_12969,N_12274);
or U14261 (N_14261,N_13445,N_12124);
xnor U14262 (N_14262,N_12631,N_13809);
nor U14263 (N_14263,N_13827,N_12130);
nand U14264 (N_14264,N_12669,N_13851);
xor U14265 (N_14265,N_12793,N_13765);
nor U14266 (N_14266,N_12932,N_13508);
nand U14267 (N_14267,N_12365,N_13886);
or U14268 (N_14268,N_12408,N_12101);
or U14269 (N_14269,N_12730,N_12164);
nor U14270 (N_14270,N_13649,N_12047);
nor U14271 (N_14271,N_13799,N_13437);
or U14272 (N_14272,N_13540,N_13109);
nand U14273 (N_14273,N_12907,N_12705);
and U14274 (N_14274,N_12879,N_13263);
or U14275 (N_14275,N_12098,N_12622);
and U14276 (N_14276,N_13449,N_12934);
xnor U14277 (N_14277,N_12340,N_12683);
nand U14278 (N_14278,N_12089,N_12672);
and U14279 (N_14279,N_12507,N_13617);
nand U14280 (N_14280,N_12636,N_12842);
nand U14281 (N_14281,N_13407,N_13362);
or U14282 (N_14282,N_13937,N_12306);
or U14283 (N_14283,N_12918,N_12677);
nand U14284 (N_14284,N_12541,N_13893);
or U14285 (N_14285,N_13605,N_13731);
or U14286 (N_14286,N_13970,N_13975);
nor U14287 (N_14287,N_12446,N_12676);
and U14288 (N_14288,N_12280,N_12108);
and U14289 (N_14289,N_12138,N_12609);
and U14290 (N_14290,N_13013,N_12086);
or U14291 (N_14291,N_13089,N_12961);
and U14292 (N_14292,N_13848,N_13563);
nand U14293 (N_14293,N_13259,N_12049);
nor U14294 (N_14294,N_13805,N_12029);
or U14295 (N_14295,N_13075,N_13163);
nor U14296 (N_14296,N_13813,N_12595);
nand U14297 (N_14297,N_13239,N_12186);
xnor U14298 (N_14298,N_13674,N_13245);
and U14299 (N_14299,N_12594,N_12247);
or U14300 (N_14300,N_12391,N_12032);
xor U14301 (N_14301,N_12113,N_13687);
nor U14302 (N_14302,N_12215,N_13127);
and U14303 (N_14303,N_12701,N_12417);
nand U14304 (N_14304,N_13456,N_12082);
nor U14305 (N_14305,N_13581,N_12656);
and U14306 (N_14306,N_12195,N_13757);
and U14307 (N_14307,N_12547,N_13055);
and U14308 (N_14308,N_13998,N_12231);
and U14309 (N_14309,N_13623,N_13591);
nor U14310 (N_14310,N_13100,N_13324);
or U14311 (N_14311,N_12212,N_12954);
and U14312 (N_14312,N_13532,N_12142);
xor U14313 (N_14313,N_13149,N_13691);
or U14314 (N_14314,N_13648,N_13685);
or U14315 (N_14315,N_12620,N_12272);
or U14316 (N_14316,N_13520,N_13121);
and U14317 (N_14317,N_13229,N_12658);
and U14318 (N_14318,N_13218,N_13046);
nor U14319 (N_14319,N_13561,N_13832);
or U14320 (N_14320,N_13355,N_13326);
or U14321 (N_14321,N_13020,N_12230);
nor U14322 (N_14322,N_12360,N_13473);
xnor U14323 (N_14323,N_13328,N_13707);
or U14324 (N_14324,N_13863,N_12814);
nor U14325 (N_14325,N_13794,N_12909);
nor U14326 (N_14326,N_13963,N_13242);
or U14327 (N_14327,N_13357,N_13944);
nand U14328 (N_14328,N_12458,N_12870);
nand U14329 (N_14329,N_12170,N_13542);
xor U14330 (N_14330,N_13625,N_12544);
or U14331 (N_14331,N_13468,N_12940);
nor U14332 (N_14332,N_13665,N_12974);
and U14333 (N_14333,N_12471,N_13626);
nor U14334 (N_14334,N_13702,N_12596);
nand U14335 (N_14335,N_12099,N_13862);
nand U14336 (N_14336,N_12648,N_13255);
nor U14337 (N_14337,N_13204,N_12567);
and U14338 (N_14338,N_13583,N_13752);
nand U14339 (N_14339,N_13057,N_13190);
nand U14340 (N_14340,N_13633,N_13464);
or U14341 (N_14341,N_13933,N_12593);
nor U14342 (N_14342,N_13784,N_12449);
or U14343 (N_14343,N_12789,N_13017);
nand U14344 (N_14344,N_13394,N_13699);
and U14345 (N_14345,N_13953,N_12549);
nor U14346 (N_14346,N_13745,N_13673);
and U14347 (N_14347,N_12203,N_13664);
nand U14348 (N_14348,N_13750,N_13351);
xnor U14349 (N_14349,N_13643,N_12645);
xor U14350 (N_14350,N_12184,N_12125);
nor U14351 (N_14351,N_13517,N_12833);
nand U14352 (N_14352,N_12201,N_13129);
or U14353 (N_14353,N_13879,N_12448);
xnor U14354 (N_14354,N_13955,N_13787);
nor U14355 (N_14355,N_12143,N_13142);
xnor U14356 (N_14356,N_12900,N_12554);
and U14357 (N_14357,N_12359,N_12128);
or U14358 (N_14358,N_12169,N_13067);
and U14359 (N_14359,N_12347,N_13334);
or U14360 (N_14360,N_12650,N_13301);
or U14361 (N_14361,N_12197,N_12811);
xor U14362 (N_14362,N_12298,N_13826);
and U14363 (N_14363,N_12476,N_12405);
nand U14364 (N_14364,N_13636,N_12718);
xor U14365 (N_14365,N_13945,N_13158);
and U14366 (N_14366,N_12482,N_13343);
and U14367 (N_14367,N_13746,N_13521);
or U14368 (N_14368,N_13928,N_12654);
nand U14369 (N_14369,N_13181,N_13714);
nor U14370 (N_14370,N_12996,N_13737);
and U14371 (N_14371,N_13670,N_13811);
or U14372 (N_14372,N_13981,N_12985);
and U14373 (N_14373,N_12442,N_13666);
nand U14374 (N_14374,N_12396,N_13104);
and U14375 (N_14375,N_13072,N_12714);
xor U14376 (N_14376,N_13137,N_13270);
and U14377 (N_14377,N_13575,N_13191);
or U14378 (N_14378,N_12558,N_13579);
xnor U14379 (N_14379,N_12068,N_13376);
and U14380 (N_14380,N_13365,N_13771);
or U14381 (N_14381,N_13052,N_13675);
xor U14382 (N_14382,N_12290,N_12267);
xor U14383 (N_14383,N_13083,N_12548);
and U14384 (N_14384,N_12559,N_13056);
nand U14385 (N_14385,N_12311,N_13414);
and U14386 (N_14386,N_13792,N_13434);
or U14387 (N_14387,N_13014,N_12221);
and U14388 (N_14388,N_13164,N_13283);
xnor U14389 (N_14389,N_12987,N_13461);
nor U14390 (N_14390,N_13847,N_13076);
nor U14391 (N_14391,N_13883,N_12467);
xnor U14392 (N_14392,N_13476,N_12898);
nand U14393 (N_14393,N_12679,N_12075);
xnor U14394 (N_14394,N_13429,N_13153);
and U14395 (N_14395,N_12137,N_13420);
and U14396 (N_14396,N_13025,N_12810);
and U14397 (N_14397,N_13860,N_13916);
and U14398 (N_14398,N_13367,N_13593);
nand U14399 (N_14399,N_12555,N_13700);
nor U14400 (N_14400,N_12296,N_13501);
nand U14401 (N_14401,N_12518,N_12585);
nand U14402 (N_14402,N_12466,N_12709);
nand U14403 (N_14403,N_12090,N_12277);
and U14404 (N_14404,N_12604,N_12322);
and U14405 (N_14405,N_13236,N_13202);
xor U14406 (N_14406,N_12104,N_13936);
xnor U14407 (N_14407,N_13932,N_12657);
or U14408 (N_14408,N_13980,N_12028);
and U14409 (N_14409,N_12259,N_12542);
and U14410 (N_14410,N_13634,N_13297);
xor U14411 (N_14411,N_12775,N_13059);
nor U14412 (N_14412,N_13804,N_12024);
or U14413 (N_14413,N_12826,N_12643);
nor U14414 (N_14414,N_12584,N_13509);
and U14415 (N_14415,N_12000,N_12463);
xor U14416 (N_14416,N_12788,N_13599);
nand U14417 (N_14417,N_12511,N_13068);
or U14418 (N_14418,N_13043,N_13327);
xnor U14419 (N_14419,N_12409,N_12545);
and U14420 (N_14420,N_13469,N_12447);
nor U14421 (N_14421,N_13151,N_13338);
nor U14422 (N_14422,N_13413,N_13240);
nand U14423 (N_14423,N_13035,N_13562);
xnor U14424 (N_14424,N_12880,N_12083);
or U14425 (N_14425,N_13843,N_12357);
and U14426 (N_14426,N_12105,N_12297);
nor U14427 (N_14427,N_12512,N_12637);
xor U14428 (N_14428,N_13011,N_12684);
or U14429 (N_14429,N_12895,N_12400);
nand U14430 (N_14430,N_13812,N_13224);
xnor U14431 (N_14431,N_12439,N_13173);
and U14432 (N_14432,N_13041,N_12249);
nor U14433 (N_14433,N_13837,N_12902);
or U14434 (N_14434,N_12486,N_13098);
xor U14435 (N_14435,N_12686,N_13747);
nand U14436 (N_14436,N_12939,N_13635);
xnor U14437 (N_14437,N_12305,N_12444);
and U14438 (N_14438,N_13391,N_12180);
or U14439 (N_14439,N_13987,N_12946);
xor U14440 (N_14440,N_12503,N_12434);
nand U14441 (N_14441,N_12399,N_13217);
nand U14442 (N_14442,N_13588,N_12838);
and U14443 (N_14443,N_12751,N_13940);
xor U14444 (N_14444,N_12027,N_12616);
and U14445 (N_14445,N_13493,N_12626);
or U14446 (N_14446,N_12007,N_12535);
nor U14447 (N_14447,N_13252,N_13788);
and U14448 (N_14448,N_13770,N_13690);
nand U14449 (N_14449,N_12022,N_12238);
nand U14450 (N_14450,N_12505,N_13352);
nand U14451 (N_14451,N_12933,N_12904);
nand U14452 (N_14452,N_12732,N_13972);
nor U14453 (N_14453,N_13506,N_13705);
nand U14454 (N_14454,N_13101,N_12829);
and U14455 (N_14455,N_13400,N_13354);
nor U14456 (N_14456,N_13103,N_12678);
nand U14457 (N_14457,N_12550,N_12608);
nand U14458 (N_14458,N_13730,N_12563);
nand U14459 (N_14459,N_13278,N_13795);
or U14460 (N_14460,N_13495,N_13511);
nor U14461 (N_14461,N_13113,N_12500);
and U14462 (N_14462,N_13680,N_12787);
nand U14463 (N_14463,N_13920,N_12854);
or U14464 (N_14464,N_13047,N_13419);
xor U14465 (N_14465,N_13444,N_12713);
nand U14466 (N_14466,N_12156,N_12173);
xor U14467 (N_14467,N_13954,N_13751);
or U14468 (N_14468,N_12013,N_12641);
nand U14469 (N_14469,N_12742,N_12074);
and U14470 (N_14470,N_13721,N_12785);
nor U14471 (N_14471,N_13514,N_13008);
nor U14472 (N_14472,N_13123,N_13210);
or U14473 (N_14473,N_13630,N_13632);
or U14474 (N_14474,N_13077,N_12039);
and U14475 (N_14475,N_12652,N_13571);
and U14476 (N_14476,N_12717,N_13696);
or U14477 (N_14477,N_12615,N_13659);
xor U14478 (N_14478,N_13526,N_12017);
nand U14479 (N_14479,N_12977,N_13265);
nor U14480 (N_14480,N_12379,N_12949);
nand U14481 (N_14481,N_12284,N_13743);
and U14482 (N_14482,N_13948,N_13346);
or U14483 (N_14483,N_12629,N_13285);
nor U14484 (N_14484,N_12148,N_13230);
nand U14485 (N_14485,N_13631,N_13924);
nor U14486 (N_14486,N_13212,N_12419);
or U14487 (N_14487,N_13835,N_13587);
nor U14488 (N_14488,N_12315,N_13782);
nand U14489 (N_14489,N_12784,N_12706);
nand U14490 (N_14490,N_13320,N_12572);
nand U14491 (N_14491,N_13742,N_13717);
and U14492 (N_14492,N_13766,N_13335);
nand U14493 (N_14493,N_12807,N_12970);
and U14494 (N_14494,N_12537,N_13036);
and U14495 (N_14495,N_12351,N_12663);
xnor U14496 (N_14496,N_12136,N_13174);
or U14497 (N_14497,N_12116,N_12495);
and U14498 (N_14498,N_13167,N_13994);
nand U14499 (N_14499,N_12316,N_13878);
and U14500 (N_14500,N_12040,N_12162);
and U14501 (N_14501,N_13214,N_13375);
nand U14502 (N_14502,N_12743,N_13486);
xnor U14503 (N_14503,N_13331,N_13310);
and U14504 (N_14504,N_12287,N_12081);
nor U14505 (N_14505,N_12133,N_12078);
xor U14506 (N_14506,N_12474,N_12690);
nand U14507 (N_14507,N_12630,N_13388);
and U14508 (N_14508,N_13725,N_12328);
and U14509 (N_14509,N_13156,N_12877);
nor U14510 (N_14510,N_12355,N_12226);
xor U14511 (N_14511,N_12883,N_12019);
nand U14512 (N_14512,N_12061,N_13477);
or U14513 (N_14513,N_12291,N_12707);
or U14514 (N_14514,N_13443,N_13807);
or U14515 (N_14515,N_12166,N_12155);
and U14516 (N_14516,N_12060,N_12944);
xor U14517 (N_14517,N_13132,N_12680);
nor U14518 (N_14518,N_12583,N_13144);
nand U14519 (N_14519,N_12185,N_13272);
and U14520 (N_14520,N_13576,N_13607);
nor U14521 (N_14521,N_13838,N_12073);
xor U14522 (N_14522,N_12096,N_12990);
xor U14523 (N_14523,N_12430,N_13081);
nor U14524 (N_14524,N_12889,N_12003);
or U14525 (N_14525,N_13087,N_12517);
xnor U14526 (N_14526,N_13462,N_12362);
or U14527 (N_14527,N_12741,N_13295);
nand U14528 (N_14528,N_13311,N_13019);
and U14529 (N_14529,N_12950,N_12882);
nor U14530 (N_14530,N_12058,N_13865);
xor U14531 (N_14531,N_13844,N_13160);
nand U14532 (N_14532,N_13256,N_12749);
and U14533 (N_14533,N_12513,N_12363);
nor U14534 (N_14534,N_13117,N_12721);
nand U14535 (N_14535,N_12345,N_12229);
nor U14536 (N_14536,N_12697,N_13740);
nand U14537 (N_14537,N_13336,N_13808);
or U14538 (N_14538,N_12823,N_13106);
nor U14539 (N_14539,N_13309,N_12568);
or U14540 (N_14540,N_13901,N_13009);
and U14541 (N_14541,N_12966,N_12619);
xor U14542 (N_14542,N_13551,N_13203);
nand U14543 (N_14543,N_13639,N_12254);
xnor U14544 (N_14544,N_12366,N_12605);
nor U14545 (N_14545,N_13681,N_12786);
nand U14546 (N_14546,N_12758,N_13231);
and U14547 (N_14547,N_13192,N_12208);
and U14548 (N_14548,N_12491,N_13726);
or U14549 (N_14549,N_12897,N_13857);
xnor U14550 (N_14550,N_13201,N_13460);
and U14551 (N_14551,N_12546,N_13300);
or U14552 (N_14552,N_13939,N_13371);
and U14553 (N_14553,N_12102,N_13775);
nor U14554 (N_14554,N_13654,N_13992);
or U14555 (N_14555,N_13550,N_12903);
or U14556 (N_14556,N_12836,N_12772);
and U14557 (N_14557,N_13573,N_13222);
nor U14558 (N_14558,N_13193,N_13951);
xor U14559 (N_14559,N_12614,N_13292);
xor U14560 (N_14560,N_12172,N_12531);
and U14561 (N_14561,N_13363,N_12655);
and U14562 (N_14562,N_13647,N_13296);
nand U14563 (N_14563,N_12455,N_13803);
nor U14564 (N_14564,N_13110,N_12927);
or U14565 (N_14565,N_13917,N_12618);
xor U14566 (N_14566,N_12181,N_13756);
and U14567 (N_14567,N_13537,N_12553);
and U14568 (N_14568,N_12905,N_12282);
or U14569 (N_14569,N_12010,N_13135);
xor U14570 (N_14570,N_13128,N_12711);
nor U14571 (N_14571,N_12937,N_13668);
and U14572 (N_14572,N_12914,N_13658);
xnor U14573 (N_14573,N_13048,N_13512);
xnor U14574 (N_14574,N_12257,N_13861);
or U14575 (N_14575,N_12590,N_12206);
or U14576 (N_14576,N_13739,N_13842);
or U14577 (N_14577,N_13119,N_13909);
or U14578 (N_14578,N_13660,N_13781);
or U14579 (N_14579,N_13629,N_12031);
and U14580 (N_14580,N_12844,N_12712);
xor U14581 (N_14581,N_13157,N_12087);
or U14582 (N_14582,N_13387,N_13425);
and U14583 (N_14583,N_13958,N_12253);
and U14584 (N_14584,N_13404,N_13806);
xnor U14585 (N_14585,N_12919,N_12338);
nand U14586 (N_14586,N_12733,N_12971);
or U14587 (N_14587,N_13438,N_12367);
nand U14588 (N_14588,N_12276,N_12727);
and U14589 (N_14589,N_13442,N_13200);
nor U14590 (N_14590,N_12863,N_12199);
and U14591 (N_14591,N_12646,N_13484);
nand U14592 (N_14592,N_12699,N_13502);
xor U14593 (N_14593,N_12748,N_13930);
nor U14594 (N_14594,N_13016,N_12234);
xnor U14595 (N_14595,N_13715,N_13188);
and U14596 (N_14596,N_12667,N_13172);
and U14597 (N_14597,N_12827,N_13641);
and U14598 (N_14598,N_12540,N_12335);
xnor U14599 (N_14599,N_12498,N_12300);
nor U14600 (N_14600,N_13761,N_13358);
xor U14601 (N_14601,N_13780,N_12516);
nand U14602 (N_14602,N_13402,N_12331);
or U14603 (N_14603,N_13060,N_13711);
xnor U14604 (N_14604,N_13139,N_12528);
and U14605 (N_14605,N_13377,N_13091);
nor U14606 (N_14606,N_13303,N_12640);
nor U14607 (N_14607,N_12030,N_13251);
nand U14608 (N_14608,N_12617,N_12119);
xor U14609 (N_14609,N_13124,N_13276);
nor U14610 (N_14610,N_13005,N_12976);
xnor U14611 (N_14611,N_13398,N_12888);
and U14612 (N_14612,N_13919,N_12852);
nand U14613 (N_14613,N_12941,N_13938);
nand U14614 (N_14614,N_12959,N_12980);
and U14615 (N_14615,N_12571,N_12427);
nor U14616 (N_14616,N_13504,N_12354);
xnor U14617 (N_14617,N_12673,N_13166);
nand U14618 (N_14618,N_13170,N_13451);
or U14619 (N_14619,N_13258,N_12232);
nand U14620 (N_14620,N_13455,N_13112);
nor U14621 (N_14621,N_12524,N_12791);
and U14622 (N_14622,N_12606,N_12938);
nand U14623 (N_14623,N_13693,N_13433);
nand U14624 (N_14624,N_12795,N_13412);
xor U14625 (N_14625,N_12369,N_12144);
or U14626 (N_14626,N_12109,N_13906);
nand U14627 (N_14627,N_12762,N_13382);
or U14628 (N_14628,N_13672,N_13488);
nand U14629 (N_14629,N_12358,N_13989);
xor U14630 (N_14630,N_13701,N_13454);
nand U14631 (N_14631,N_13225,N_12598);
or U14632 (N_14632,N_12440,N_13314);
and U14633 (N_14633,N_13279,N_13260);
and U14634 (N_14634,N_13875,N_13463);
or U14635 (N_14635,N_13102,N_12644);
and U14636 (N_14636,N_12388,N_13510);
nand U14637 (N_14637,N_13439,N_13595);
nor U14638 (N_14638,N_12892,N_12385);
and U14639 (N_14639,N_13709,N_12945);
and U14640 (N_14640,N_13483,N_13024);
and U14641 (N_14641,N_13042,N_13208);
nor U14642 (N_14642,N_13361,N_12948);
or U14643 (N_14643,N_13858,N_12722);
nor U14644 (N_14644,N_12715,N_13053);
and U14645 (N_14645,N_13976,N_13874);
nor U14646 (N_14646,N_13565,N_12999);
and U14647 (N_14647,N_12700,N_12429);
and U14648 (N_14648,N_12850,N_13392);
nor U14649 (N_14649,N_13289,N_13162);
xnor U14650 (N_14650,N_13620,N_13074);
and U14651 (N_14651,N_13028,N_13094);
nand U14652 (N_14652,N_12824,N_13818);
nor U14653 (N_14653,N_13436,N_12632);
or U14654 (N_14654,N_12364,N_13154);
and U14655 (N_14655,N_13097,N_12383);
xor U14656 (N_14656,N_12233,N_12228);
nor U14657 (N_14657,N_13254,N_12381);
nand U14658 (N_14658,N_13446,N_12963);
and U14659 (N_14659,N_13418,N_13308);
nand U14660 (N_14660,N_13965,N_12456);
or U14661 (N_14661,N_12964,N_12800);
and U14662 (N_14662,N_13141,N_13305);
and U14663 (N_14663,N_13175,N_13934);
and U14664 (N_14664,N_13114,N_12740);
nor U14665 (N_14665,N_12832,N_13661);
or U14666 (N_14666,N_12659,N_12913);
nor U14667 (N_14667,N_12223,N_12077);
nand U14668 (N_14668,N_12350,N_12851);
and U14669 (N_14669,N_12472,N_12450);
nor U14670 (N_14670,N_13619,N_13390);
nand U14671 (N_14671,N_12132,N_12576);
xor U14672 (N_14672,N_13337,N_13273);
or U14673 (N_14673,N_12747,N_13814);
xor U14674 (N_14674,N_13183,N_12822);
and U14675 (N_14675,N_12216,N_13902);
or U14676 (N_14676,N_13374,N_12508);
and U14677 (N_14677,N_12804,N_13567);
nor U14678 (N_14678,N_12323,N_13615);
nor U14679 (N_14679,N_13001,N_13054);
nand U14680 (N_14680,N_13871,N_13651);
and U14681 (N_14681,N_12387,N_13719);
xnor U14682 (N_14682,N_12219,N_12225);
xnor U14683 (N_14683,N_13205,N_13676);
or U14684 (N_14684,N_12084,N_12993);
xor U14685 (N_14685,N_13498,N_12891);
nor U14686 (N_14686,N_12349,N_13925);
nand U14687 (N_14687,N_12975,N_13825);
nand U14688 (N_14688,N_13180,N_12337);
or U14689 (N_14689,N_13199,N_13380);
and U14690 (N_14690,N_13820,N_13485);
or U14691 (N_14691,N_13389,N_13910);
and U14692 (N_14692,N_13926,N_12773);
xor U14693 (N_14693,N_13791,N_12317);
nor U14694 (N_14694,N_12682,N_12341);
nand U14695 (N_14695,N_12651,N_13474);
and U14696 (N_14696,N_13969,N_13187);
xor U14697 (N_14697,N_13610,N_13241);
and U14698 (N_14698,N_12194,N_12642);
and U14699 (N_14699,N_12930,N_12694);
nand U14700 (N_14700,N_12664,N_13126);
nor U14701 (N_14701,N_12348,N_13880);
xnor U14702 (N_14702,N_12151,N_12242);
or U14703 (N_14703,N_13266,N_12489);
nand U14704 (N_14704,N_12872,N_13708);
nor U14705 (N_14705,N_12668,N_13908);
nand U14706 (N_14706,N_12812,N_12514);
nand U14707 (N_14707,N_12200,N_13850);
nor U14708 (N_14708,N_13082,N_13247);
xor U14709 (N_14709,N_12573,N_13459);
or U14710 (N_14710,N_12704,N_12309);
xor U14711 (N_14711,N_12532,N_12343);
and U14712 (N_14712,N_12246,N_13386);
or U14713 (N_14713,N_13882,N_13755);
and U14714 (N_14714,N_12288,N_12601);
nor U14715 (N_14715,N_13779,N_13716);
or U14716 (N_14716,N_12808,N_13304);
and U14717 (N_14717,N_12177,N_12055);
nor U14718 (N_14718,N_13505,N_13487);
or U14719 (N_14719,N_13373,N_13773);
nor U14720 (N_14720,N_13284,N_12394);
and U14721 (N_14721,N_12041,N_12750);
nand U14722 (N_14722,N_12797,N_13558);
nand U14723 (N_14723,N_13482,N_12160);
and U14724 (N_14724,N_12182,N_12235);
nor U14725 (N_14725,N_13735,N_12884);
nand U14726 (N_14726,N_12790,N_12858);
xnor U14727 (N_14727,N_13572,N_13962);
or U14728 (N_14728,N_12336,N_13323);
xor U14729 (N_14729,N_12054,N_12603);
or U14730 (N_14730,N_13618,N_12326);
or U14731 (N_14731,N_12431,N_13884);
or U14732 (N_14732,N_12260,N_13895);
nand U14733 (N_14733,N_12506,N_13161);
nor U14734 (N_14734,N_13704,N_13783);
and U14735 (N_14735,N_12076,N_12771);
nor U14736 (N_14736,N_13652,N_12384);
xor U14737 (N_14737,N_12768,N_13417);
and U14738 (N_14738,N_13898,N_13684);
or U14739 (N_14739,N_13749,N_12562);
and U14740 (N_14740,N_13470,N_13169);
and U14741 (N_14741,N_13274,N_12412);
xor U14742 (N_14742,N_12044,N_13472);
xor U14743 (N_14743,N_12777,N_13497);
nor U14744 (N_14744,N_12411,N_12866);
nand U14745 (N_14745,N_12294,N_12765);
and U14746 (N_14746,N_12063,N_13545);
xnor U14747 (N_14747,N_12509,N_13689);
nand U14748 (N_14748,N_12307,N_12911);
xnor U14749 (N_14749,N_12796,N_12403);
nand U14750 (N_14750,N_13264,N_12855);
or U14751 (N_14751,N_13248,N_12998);
nand U14752 (N_14752,N_12639,N_12213);
nor U14753 (N_14753,N_12372,N_12716);
nor U14754 (N_14754,N_12112,N_12204);
and U14755 (N_14755,N_12401,N_13275);
or U14756 (N_14756,N_12764,N_12708);
nor U14757 (N_14757,N_13494,N_13287);
nand U14758 (N_14758,N_12774,N_13982);
xnor U14759 (N_14759,N_13824,N_13378);
or U14760 (N_14760,N_12469,N_12079);
and U14761 (N_14761,N_12995,N_12303);
nor U14762 (N_14762,N_13543,N_12339);
or U14763 (N_14763,N_12965,N_12735);
and U14764 (N_14764,N_13063,N_12018);
xnor U14765 (N_14765,N_13754,N_12623);
or U14766 (N_14766,N_13032,N_13758);
nand U14767 (N_14767,N_12488,N_12239);
xor U14768 (N_14768,N_12957,N_13853);
or U14769 (N_14769,N_12533,N_12521);
nand U14770 (N_14770,N_12275,N_12139);
nor U14771 (N_14771,N_13138,N_13179);
nand U14772 (N_14772,N_12457,N_13333);
nand U14773 (N_14773,N_13697,N_13211);
and U14774 (N_14774,N_13720,N_12126);
nor U14775 (N_14775,N_12534,N_12038);
xnor U14776 (N_14776,N_12023,N_12634);
or U14777 (N_14777,N_13548,N_13209);
xnor U14778 (N_14778,N_13395,N_13159);
nor U14779 (N_14779,N_13228,N_12241);
nor U14780 (N_14780,N_13774,N_13616);
or U14781 (N_14781,N_12579,N_13710);
or U14782 (N_14782,N_12728,N_12670);
nand U14783 (N_14783,N_12587,N_13234);
or U14784 (N_14784,N_13165,N_13957);
xnor U14785 (N_14785,N_13261,N_13539);
nand U14786 (N_14786,N_12183,N_13213);
and U14787 (N_14787,N_12857,N_12530);
xnor U14788 (N_14788,N_13622,N_13195);
and U14789 (N_14789,N_13786,N_12187);
xnor U14790 (N_14790,N_13995,N_12262);
and U14791 (N_14791,N_12853,N_12525);
nor U14792 (N_14792,N_13600,N_12837);
nand U14793 (N_14793,N_12236,N_12397);
nand U14794 (N_14794,N_13249,N_13546);
xnor U14795 (N_14795,N_12295,N_13238);
xnor U14796 (N_14796,N_13288,N_13695);
nand U14797 (N_14797,N_12660,N_13555);
nor U14798 (N_14798,N_12958,N_12103);
nor U14799 (N_14799,N_12069,N_13613);
nand U14800 (N_14800,N_12627,N_12624);
or U14801 (N_14801,N_13596,N_13964);
nor U14802 (N_14802,N_12861,N_12150);
xnor U14803 (N_14803,N_13828,N_12012);
nor U14804 (N_14804,N_13829,N_12420);
nor U14805 (N_14805,N_12539,N_12178);
nand U14806 (N_14806,N_13973,N_13370);
nor U14807 (N_14807,N_12666,N_13232);
or U14808 (N_14808,N_13594,N_12695);
nor U14809 (N_14809,N_12894,N_12575);
nor U14810 (N_14810,N_12056,N_13640);
xnor U14811 (N_14811,N_12325,N_12910);
nor U14812 (N_14812,N_12923,N_12929);
xnor U14813 (N_14813,N_12092,N_12947);
nor U14814 (N_14814,N_12874,N_13852);
nand U14815 (N_14815,N_13359,N_12211);
xnor U14816 (N_14816,N_12873,N_13644);
or U14817 (N_14817,N_13131,N_12237);
nor U14818 (N_14818,N_12597,N_13253);
or U14819 (N_14819,N_13152,N_12342);
xnor U14820 (N_14820,N_13084,N_12817);
and U14821 (N_14821,N_12492,N_12744);
nand U14822 (N_14822,N_13344,N_13568);
xnor U14823 (N_14823,N_12560,N_12906);
nor U14824 (N_14824,N_12611,N_13891);
or U14825 (N_14825,N_13646,N_12869);
and U14826 (N_14826,N_12752,N_12671);
and U14827 (N_14827,N_13921,N_13778);
and U14828 (N_14828,N_12261,N_12719);
nor U14829 (N_14829,N_13834,N_13150);
and U14830 (N_14830,N_13441,N_13892);
xnor U14831 (N_14831,N_13227,N_12445);
xnor U14832 (N_14832,N_13090,N_13904);
xor U14833 (N_14833,N_12161,N_13026);
and U14834 (N_14834,N_12922,N_13221);
nand U14835 (N_14835,N_12522,N_13286);
and U14836 (N_14836,N_13039,N_13650);
and U14837 (N_14837,N_12464,N_13603);
xor U14838 (N_14838,N_12696,N_13233);
and U14839 (N_14839,N_13207,N_12051);
and U14840 (N_14840,N_12504,N_12794);
and U14841 (N_14841,N_12483,N_12461);
nor U14842 (N_14842,N_12222,N_13686);
nand U14843 (N_14843,N_12725,N_12763);
and U14844 (N_14844,N_12908,N_12828);
nor U14845 (N_14845,N_12523,N_13777);
nand U14846 (N_14846,N_12997,N_13219);
xor U14847 (N_14847,N_12413,N_13977);
or U14848 (N_14848,N_13741,N_13316);
or U14849 (N_14849,N_13347,N_12395);
xor U14850 (N_14850,N_12776,N_12876);
or U14851 (N_14851,N_13471,N_12710);
and U14852 (N_14852,N_13330,N_12755);
nor U14853 (N_14853,N_12956,N_13513);
nand U14854 (N_14854,N_12820,N_13590);
xnor U14855 (N_14855,N_12373,N_12433);
or U14856 (N_14856,N_13798,N_12661);
nand U14857 (N_14857,N_12292,N_13728);
nor U14858 (N_14858,N_13421,N_12953);
nor U14859 (N_14859,N_13044,N_12220);
nand U14860 (N_14860,N_13947,N_13956);
nand U14861 (N_14861,N_13918,N_13453);
and U14862 (N_14862,N_12638,N_12578);
nor U14863 (N_14863,N_13985,N_13817);
nor U14864 (N_14864,N_12703,N_12252);
xnor U14865 (N_14865,N_13503,N_12767);
nand U14866 (N_14866,N_13313,N_13396);
nand U14867 (N_14867,N_12494,N_13034);
or U14868 (N_14868,N_13983,N_13793);
and U14869 (N_14869,N_12982,N_13569);
xnor U14870 (N_14870,N_13226,N_12994);
or U14871 (N_14871,N_12071,N_12064);
and U14872 (N_14872,N_13722,N_12263);
xnor U14873 (N_14873,N_13996,N_13990);
or U14874 (N_14874,N_13868,N_13564);
or U14875 (N_14875,N_13911,N_12250);
and U14876 (N_14876,N_13379,N_12893);
or U14877 (N_14877,N_13022,N_13678);
xnor U14878 (N_14878,N_13073,N_12760);
and U14879 (N_14879,N_12586,N_13216);
nor U14880 (N_14880,N_12393,N_12847);
and U14881 (N_14881,N_12868,N_13971);
and U14882 (N_14882,N_12436,N_12770);
nand U14883 (N_14883,N_13147,N_13277);
and U14884 (N_14884,N_13424,N_13764);
xor U14885 (N_14885,N_12761,N_13079);
xor U14886 (N_14886,N_12809,N_13557);
and U14887 (N_14887,N_12193,N_12091);
or U14888 (N_14888,N_12871,N_13130);
and U14889 (N_14889,N_13923,N_12344);
or U14890 (N_14890,N_12731,N_12681);
and U14891 (N_14891,N_13949,N_13360);
nor U14892 (N_14892,N_13667,N_13662);
and U14893 (N_14893,N_12406,N_13401);
or U14894 (N_14894,N_13669,N_13406);
and U14895 (N_14895,N_12371,N_12279);
and U14896 (N_14896,N_13134,N_12834);
nand U14897 (N_14897,N_12591,N_13366);
and U14898 (N_14898,N_12885,N_12134);
xnor U14899 (N_14899,N_13341,N_12723);
or U14900 (N_14900,N_12867,N_12453);
nand U14901 (N_14901,N_13176,N_12021);
and U14902 (N_14902,N_12766,N_12129);
xnor U14903 (N_14903,N_12088,N_12441);
xor U14904 (N_14904,N_12392,N_13589);
and U14905 (N_14905,N_12633,N_12589);
nor U14906 (N_14906,N_13012,N_12759);
nand U14907 (N_14907,N_13845,N_13896);
and U14908 (N_14908,N_13903,N_12310);
nor U14909 (N_14909,N_12330,N_13171);
and U14910 (N_14910,N_13760,N_13384);
or U14911 (N_14911,N_13440,N_13524);
and U14912 (N_14912,N_13888,N_12801);
nand U14913 (N_14913,N_12816,N_12198);
nand U14914 (N_14914,N_13093,N_13051);
xor U14915 (N_14915,N_13307,N_13915);
nand U14916 (N_14916,N_12475,N_13724);
xnor U14917 (N_14917,N_13061,N_12011);
nand U14918 (N_14918,N_12881,N_13350);
xnor U14919 (N_14919,N_13243,N_12739);
or U14920 (N_14920,N_13049,N_13329);
or U14921 (N_14921,N_13050,N_12062);
xor U14922 (N_14922,N_12244,N_12191);
nand U14923 (N_14923,N_13523,N_12519);
and U14924 (N_14924,N_12734,N_12066);
nor U14925 (N_14925,N_13846,N_12080);
or U14926 (N_14926,N_13492,N_13645);
or U14927 (N_14927,N_12240,N_12293);
nand U14928 (N_14928,N_13481,N_12001);
nand U14929 (N_14929,N_13897,N_13294);
nor U14930 (N_14930,N_12438,N_12157);
and U14931 (N_14931,N_13196,N_13250);
xor U14932 (N_14932,N_13349,N_12564);
nand U14933 (N_14933,N_12921,N_13769);
or U14934 (N_14934,N_12285,N_13967);
nand U14935 (N_14935,N_12067,N_13003);
nand U14936 (N_14936,N_13759,N_13597);
and U14937 (N_14937,N_13978,N_13815);
and U14938 (N_14938,N_13656,N_12972);
or U14939 (N_14939,N_12510,N_12141);
nand U14940 (N_14940,N_12501,N_13900);
and U14941 (N_14941,N_12210,N_13876);
and U14942 (N_14942,N_12320,N_12726);
nand U14943 (N_14943,N_13753,N_13790);
xor U14944 (N_14944,N_13655,N_12783);
xnor U14945 (N_14945,N_13734,N_12931);
xor U14946 (N_14946,N_12059,N_13604);
xor U14947 (N_14947,N_13960,N_12991);
or U14948 (N_14948,N_12843,N_13116);
or U14949 (N_14949,N_12757,N_12422);
and U14950 (N_14950,N_13519,N_12304);
nand U14951 (N_14951,N_13499,N_13058);
xnor U14952 (N_14952,N_13426,N_12094);
nor U14953 (N_14953,N_12935,N_12487);
xor U14954 (N_14954,N_12025,N_12319);
nor U14955 (N_14955,N_12374,N_13821);
and U14956 (N_14956,N_13447,N_13866);
xnor U14957 (N_14957,N_12462,N_12859);
and U14958 (N_14958,N_12289,N_12782);
nand U14959 (N_14959,N_12536,N_13185);
nand U14960 (N_14960,N_13122,N_12356);
nor U14961 (N_14961,N_13332,N_13430);
xor U14962 (N_14962,N_13408,N_13133);
nand U14963 (N_14963,N_12687,N_12581);
nor U14964 (N_14964,N_12951,N_12154);
or U14965 (N_14965,N_12255,N_13269);
or U14966 (N_14966,N_12745,N_13480);
and U14967 (N_14967,N_12321,N_12426);
nand U14968 (N_14968,N_12418,N_12778);
and U14969 (N_14969,N_12333,N_12864);
nor U14970 (N_14970,N_13553,N_13733);
nand U14971 (N_14971,N_13997,N_12015);
nor U14972 (N_14972,N_13638,N_13864);
xnor U14973 (N_14973,N_13529,N_12561);
nor U14974 (N_14974,N_13698,N_13315);
and U14975 (N_14975,N_12915,N_13340);
or U14976 (N_14976,N_12570,N_13302);
or U14977 (N_14977,N_13069,N_12806);
nand U14978 (N_14978,N_13267,N_12955);
or U14979 (N_14979,N_13029,N_13713);
nand U14980 (N_14980,N_13064,N_12815);
nor U14981 (N_14981,N_12042,N_13348);
or U14982 (N_14982,N_12301,N_13538);
and U14983 (N_14983,N_12849,N_12135);
nor U14984 (N_14984,N_13941,N_13931);
xnor U14985 (N_14985,N_13712,N_13612);
nand U14986 (N_14986,N_13833,N_13912);
or U14987 (N_14987,N_13155,N_13979);
nand U14988 (N_14988,N_13683,N_12050);
nand U14989 (N_14989,N_13318,N_12265);
or U14990 (N_14990,N_12005,N_13566);
xor U14991 (N_14991,N_12662,N_13601);
nor U14992 (N_14992,N_13325,N_12421);
nor U14993 (N_14993,N_12612,N_12097);
and U14994 (N_14994,N_12370,N_13988);
nand U14995 (N_14995,N_13280,N_12036);
or U14996 (N_14996,N_13830,N_13037);
and U14997 (N_14997,N_13968,N_12924);
or U14998 (N_14998,N_13841,N_13839);
nand U14999 (N_14999,N_13368,N_12978);
xor U15000 (N_15000,N_13758,N_13419);
and U15001 (N_15001,N_12243,N_13134);
nor U15002 (N_15002,N_13265,N_13019);
nand U15003 (N_15003,N_12276,N_13042);
nand U15004 (N_15004,N_13565,N_12128);
nand U15005 (N_15005,N_13070,N_13466);
and U15006 (N_15006,N_13533,N_13505);
nand U15007 (N_15007,N_12779,N_12787);
nor U15008 (N_15008,N_13233,N_12279);
and U15009 (N_15009,N_12080,N_12966);
nand U15010 (N_15010,N_12863,N_12188);
nand U15011 (N_15011,N_13562,N_12188);
and U15012 (N_15012,N_12982,N_12903);
xor U15013 (N_15013,N_12574,N_13795);
or U15014 (N_15014,N_12681,N_13820);
or U15015 (N_15015,N_12947,N_13920);
nor U15016 (N_15016,N_12220,N_12234);
xor U15017 (N_15017,N_13268,N_12727);
xor U15018 (N_15018,N_12351,N_13968);
xor U15019 (N_15019,N_13040,N_12800);
nor U15020 (N_15020,N_13578,N_13071);
or U15021 (N_15021,N_13805,N_13983);
nand U15022 (N_15022,N_12876,N_13135);
or U15023 (N_15023,N_12099,N_12904);
or U15024 (N_15024,N_13177,N_12166);
nand U15025 (N_15025,N_13153,N_13406);
xnor U15026 (N_15026,N_13130,N_13887);
xor U15027 (N_15027,N_13677,N_12035);
nand U15028 (N_15028,N_13079,N_12134);
nand U15029 (N_15029,N_13247,N_12857);
nor U15030 (N_15030,N_12172,N_13694);
or U15031 (N_15031,N_12650,N_12850);
and U15032 (N_15032,N_12083,N_12839);
or U15033 (N_15033,N_12701,N_13789);
nand U15034 (N_15034,N_13577,N_13056);
nor U15035 (N_15035,N_12469,N_13216);
or U15036 (N_15036,N_12727,N_13215);
or U15037 (N_15037,N_13441,N_13351);
nor U15038 (N_15038,N_12988,N_12841);
nor U15039 (N_15039,N_13288,N_13839);
xnor U15040 (N_15040,N_13209,N_12040);
nand U15041 (N_15041,N_12322,N_13501);
or U15042 (N_15042,N_12876,N_13731);
nand U15043 (N_15043,N_13233,N_12689);
nand U15044 (N_15044,N_12941,N_13274);
nand U15045 (N_15045,N_13171,N_13834);
xor U15046 (N_15046,N_12003,N_12707);
nand U15047 (N_15047,N_13610,N_12292);
nor U15048 (N_15048,N_13454,N_13657);
or U15049 (N_15049,N_13310,N_12405);
nand U15050 (N_15050,N_12408,N_12536);
nor U15051 (N_15051,N_12037,N_13330);
nor U15052 (N_15052,N_12958,N_13315);
or U15053 (N_15053,N_13939,N_13655);
nand U15054 (N_15054,N_12741,N_13635);
xor U15055 (N_15055,N_12285,N_13816);
and U15056 (N_15056,N_13513,N_13249);
or U15057 (N_15057,N_13246,N_13118);
or U15058 (N_15058,N_12866,N_12481);
nand U15059 (N_15059,N_12791,N_13861);
nand U15060 (N_15060,N_13280,N_12484);
nor U15061 (N_15061,N_13037,N_12944);
nand U15062 (N_15062,N_13501,N_13035);
xnor U15063 (N_15063,N_12314,N_13412);
and U15064 (N_15064,N_13623,N_12635);
and U15065 (N_15065,N_13867,N_13539);
or U15066 (N_15066,N_13916,N_12149);
nor U15067 (N_15067,N_13830,N_13433);
nor U15068 (N_15068,N_13894,N_13273);
and U15069 (N_15069,N_13122,N_12580);
nor U15070 (N_15070,N_12710,N_13680);
and U15071 (N_15071,N_13081,N_12096);
xor U15072 (N_15072,N_13586,N_13591);
and U15073 (N_15073,N_13395,N_13219);
xnor U15074 (N_15074,N_12210,N_12865);
and U15075 (N_15075,N_13366,N_12839);
nand U15076 (N_15076,N_13624,N_12814);
nor U15077 (N_15077,N_12346,N_13501);
nor U15078 (N_15078,N_12195,N_13429);
nand U15079 (N_15079,N_13924,N_13925);
nand U15080 (N_15080,N_12447,N_12265);
nand U15081 (N_15081,N_12065,N_13188);
and U15082 (N_15082,N_13659,N_12540);
nand U15083 (N_15083,N_13993,N_13608);
nand U15084 (N_15084,N_12338,N_12868);
and U15085 (N_15085,N_12737,N_12336);
or U15086 (N_15086,N_12432,N_13037);
and U15087 (N_15087,N_13801,N_13628);
or U15088 (N_15088,N_13185,N_13103);
or U15089 (N_15089,N_12371,N_12132);
or U15090 (N_15090,N_13331,N_13983);
and U15091 (N_15091,N_12009,N_12901);
or U15092 (N_15092,N_13216,N_12380);
nor U15093 (N_15093,N_12091,N_13486);
nor U15094 (N_15094,N_13213,N_12018);
nand U15095 (N_15095,N_13087,N_12687);
nor U15096 (N_15096,N_13204,N_13775);
or U15097 (N_15097,N_12014,N_12575);
nor U15098 (N_15098,N_12474,N_13100);
or U15099 (N_15099,N_12081,N_12048);
nor U15100 (N_15100,N_12084,N_12935);
and U15101 (N_15101,N_13690,N_12713);
xor U15102 (N_15102,N_12757,N_13982);
nor U15103 (N_15103,N_13761,N_13062);
or U15104 (N_15104,N_12255,N_13565);
or U15105 (N_15105,N_13450,N_13110);
and U15106 (N_15106,N_13405,N_12266);
xor U15107 (N_15107,N_13087,N_12470);
xor U15108 (N_15108,N_13553,N_13483);
nand U15109 (N_15109,N_12183,N_13848);
and U15110 (N_15110,N_12697,N_13421);
nor U15111 (N_15111,N_13139,N_12669);
and U15112 (N_15112,N_13160,N_13636);
or U15113 (N_15113,N_12005,N_12469);
or U15114 (N_15114,N_13677,N_12805);
xnor U15115 (N_15115,N_12971,N_13134);
or U15116 (N_15116,N_12612,N_12749);
and U15117 (N_15117,N_13050,N_12313);
nor U15118 (N_15118,N_13818,N_12719);
nand U15119 (N_15119,N_12292,N_12374);
or U15120 (N_15120,N_12146,N_13719);
nor U15121 (N_15121,N_12418,N_12553);
xor U15122 (N_15122,N_12578,N_12986);
nand U15123 (N_15123,N_12881,N_13586);
nand U15124 (N_15124,N_13468,N_13006);
nand U15125 (N_15125,N_12851,N_12309);
nor U15126 (N_15126,N_12733,N_12773);
nand U15127 (N_15127,N_13508,N_12778);
nand U15128 (N_15128,N_13385,N_12312);
and U15129 (N_15129,N_13991,N_13435);
nor U15130 (N_15130,N_12223,N_13402);
nand U15131 (N_15131,N_12318,N_13648);
or U15132 (N_15132,N_13881,N_13596);
and U15133 (N_15133,N_13509,N_13224);
and U15134 (N_15134,N_13506,N_13620);
and U15135 (N_15135,N_12753,N_13102);
nand U15136 (N_15136,N_13928,N_13415);
or U15137 (N_15137,N_12970,N_12601);
nand U15138 (N_15138,N_12681,N_12600);
or U15139 (N_15139,N_13604,N_12192);
nand U15140 (N_15140,N_12831,N_12256);
xnor U15141 (N_15141,N_12106,N_12702);
nand U15142 (N_15142,N_12626,N_13998);
or U15143 (N_15143,N_12366,N_13127);
or U15144 (N_15144,N_12158,N_13358);
nand U15145 (N_15145,N_12920,N_12941);
nand U15146 (N_15146,N_13964,N_13510);
or U15147 (N_15147,N_13489,N_12796);
nor U15148 (N_15148,N_13051,N_13274);
nor U15149 (N_15149,N_12578,N_12921);
or U15150 (N_15150,N_13986,N_13389);
nand U15151 (N_15151,N_13899,N_13661);
xnor U15152 (N_15152,N_13711,N_12842);
xor U15153 (N_15153,N_12971,N_13891);
or U15154 (N_15154,N_13136,N_12686);
and U15155 (N_15155,N_12062,N_13112);
and U15156 (N_15156,N_13217,N_12620);
and U15157 (N_15157,N_13578,N_12859);
and U15158 (N_15158,N_12431,N_13837);
and U15159 (N_15159,N_12944,N_12134);
xor U15160 (N_15160,N_13567,N_12913);
xor U15161 (N_15161,N_13694,N_12468);
or U15162 (N_15162,N_12010,N_12455);
xnor U15163 (N_15163,N_13055,N_13457);
nand U15164 (N_15164,N_13993,N_12088);
nor U15165 (N_15165,N_12955,N_13206);
xnor U15166 (N_15166,N_12690,N_13642);
and U15167 (N_15167,N_12834,N_12728);
or U15168 (N_15168,N_12744,N_13027);
nand U15169 (N_15169,N_13261,N_12751);
nor U15170 (N_15170,N_12457,N_12292);
nor U15171 (N_15171,N_12423,N_13172);
nand U15172 (N_15172,N_13433,N_13602);
and U15173 (N_15173,N_13767,N_13851);
xor U15174 (N_15174,N_13940,N_13271);
and U15175 (N_15175,N_12655,N_13163);
nand U15176 (N_15176,N_13935,N_12030);
nand U15177 (N_15177,N_12280,N_12381);
or U15178 (N_15178,N_12702,N_12777);
nand U15179 (N_15179,N_13702,N_12611);
nand U15180 (N_15180,N_13205,N_13409);
or U15181 (N_15181,N_13301,N_13782);
or U15182 (N_15182,N_12357,N_12447);
nor U15183 (N_15183,N_12257,N_13272);
and U15184 (N_15184,N_12979,N_13316);
and U15185 (N_15185,N_12746,N_13093);
nand U15186 (N_15186,N_12398,N_12863);
and U15187 (N_15187,N_13597,N_13494);
and U15188 (N_15188,N_13629,N_13553);
nor U15189 (N_15189,N_12947,N_13014);
and U15190 (N_15190,N_12462,N_12135);
and U15191 (N_15191,N_13736,N_13500);
xor U15192 (N_15192,N_12773,N_13564);
nor U15193 (N_15193,N_12106,N_13409);
nand U15194 (N_15194,N_12261,N_13879);
nor U15195 (N_15195,N_12081,N_13425);
and U15196 (N_15196,N_12040,N_12639);
or U15197 (N_15197,N_12898,N_12324);
or U15198 (N_15198,N_13279,N_12375);
xnor U15199 (N_15199,N_12798,N_12807);
or U15200 (N_15200,N_13623,N_12819);
or U15201 (N_15201,N_12298,N_13557);
xnor U15202 (N_15202,N_12713,N_13413);
nand U15203 (N_15203,N_13461,N_12128);
nor U15204 (N_15204,N_13469,N_12815);
nor U15205 (N_15205,N_13950,N_12227);
or U15206 (N_15206,N_12449,N_13534);
and U15207 (N_15207,N_13388,N_13262);
and U15208 (N_15208,N_12837,N_12533);
nor U15209 (N_15209,N_13596,N_13784);
and U15210 (N_15210,N_12034,N_13251);
xor U15211 (N_15211,N_13164,N_12347);
xnor U15212 (N_15212,N_12083,N_12558);
nor U15213 (N_15213,N_12829,N_12949);
nor U15214 (N_15214,N_13776,N_13724);
nand U15215 (N_15215,N_13388,N_12940);
xnor U15216 (N_15216,N_13365,N_13246);
xor U15217 (N_15217,N_13619,N_13676);
nand U15218 (N_15218,N_13441,N_13008);
nand U15219 (N_15219,N_12785,N_12446);
and U15220 (N_15220,N_12046,N_13505);
and U15221 (N_15221,N_12984,N_13995);
nand U15222 (N_15222,N_12917,N_13964);
xor U15223 (N_15223,N_12176,N_12486);
xnor U15224 (N_15224,N_13964,N_13440);
nor U15225 (N_15225,N_12045,N_13223);
or U15226 (N_15226,N_12474,N_13432);
or U15227 (N_15227,N_13340,N_12583);
nor U15228 (N_15228,N_12542,N_12641);
nor U15229 (N_15229,N_12711,N_12200);
and U15230 (N_15230,N_12173,N_13147);
nor U15231 (N_15231,N_13047,N_12396);
nor U15232 (N_15232,N_12140,N_13601);
nor U15233 (N_15233,N_13088,N_13503);
and U15234 (N_15234,N_12281,N_13591);
xnor U15235 (N_15235,N_13512,N_13067);
and U15236 (N_15236,N_12167,N_12359);
nor U15237 (N_15237,N_12346,N_13387);
xnor U15238 (N_15238,N_12635,N_12787);
and U15239 (N_15239,N_12598,N_12032);
nand U15240 (N_15240,N_12304,N_12866);
nand U15241 (N_15241,N_12497,N_12330);
xnor U15242 (N_15242,N_12304,N_12639);
and U15243 (N_15243,N_13773,N_13510);
nand U15244 (N_15244,N_12021,N_13963);
or U15245 (N_15245,N_12438,N_13872);
nand U15246 (N_15246,N_12674,N_13465);
or U15247 (N_15247,N_12114,N_13521);
and U15248 (N_15248,N_13841,N_12235);
or U15249 (N_15249,N_12865,N_13296);
xnor U15250 (N_15250,N_13791,N_12774);
or U15251 (N_15251,N_13066,N_13726);
nor U15252 (N_15252,N_13716,N_12350);
nor U15253 (N_15253,N_12510,N_13161);
nor U15254 (N_15254,N_13192,N_13854);
nor U15255 (N_15255,N_13878,N_12078);
nand U15256 (N_15256,N_12653,N_12651);
nand U15257 (N_15257,N_12749,N_12147);
and U15258 (N_15258,N_12599,N_12767);
xnor U15259 (N_15259,N_12639,N_12955);
and U15260 (N_15260,N_13421,N_12939);
and U15261 (N_15261,N_13131,N_13395);
or U15262 (N_15262,N_12232,N_13167);
or U15263 (N_15263,N_12087,N_13512);
and U15264 (N_15264,N_13072,N_12434);
nor U15265 (N_15265,N_12493,N_13111);
and U15266 (N_15266,N_13311,N_12427);
and U15267 (N_15267,N_12755,N_12377);
or U15268 (N_15268,N_12087,N_13929);
xor U15269 (N_15269,N_13187,N_12898);
nand U15270 (N_15270,N_12719,N_13013);
and U15271 (N_15271,N_13922,N_12242);
and U15272 (N_15272,N_12588,N_12864);
and U15273 (N_15273,N_12707,N_12180);
nor U15274 (N_15274,N_13309,N_13912);
and U15275 (N_15275,N_13083,N_12105);
or U15276 (N_15276,N_12456,N_12090);
nor U15277 (N_15277,N_13600,N_13837);
nand U15278 (N_15278,N_13719,N_12715);
nand U15279 (N_15279,N_12753,N_12665);
nor U15280 (N_15280,N_13875,N_12884);
or U15281 (N_15281,N_12169,N_13881);
and U15282 (N_15282,N_12026,N_13392);
xor U15283 (N_15283,N_12771,N_12711);
and U15284 (N_15284,N_12386,N_12894);
or U15285 (N_15285,N_12203,N_13673);
xor U15286 (N_15286,N_13029,N_13745);
xnor U15287 (N_15287,N_12278,N_13109);
and U15288 (N_15288,N_13868,N_12370);
nor U15289 (N_15289,N_13374,N_13195);
and U15290 (N_15290,N_13116,N_13854);
or U15291 (N_15291,N_13304,N_13032);
nor U15292 (N_15292,N_12416,N_12807);
and U15293 (N_15293,N_13159,N_12948);
nand U15294 (N_15294,N_12778,N_13485);
and U15295 (N_15295,N_13997,N_12120);
and U15296 (N_15296,N_12092,N_13704);
xnor U15297 (N_15297,N_13622,N_12453);
xnor U15298 (N_15298,N_13453,N_13631);
nor U15299 (N_15299,N_12335,N_12836);
nor U15300 (N_15300,N_12251,N_12081);
nand U15301 (N_15301,N_13674,N_12497);
and U15302 (N_15302,N_12877,N_13758);
nand U15303 (N_15303,N_13290,N_13684);
nand U15304 (N_15304,N_12456,N_12184);
nor U15305 (N_15305,N_13665,N_13772);
and U15306 (N_15306,N_13659,N_12082);
and U15307 (N_15307,N_13793,N_12070);
and U15308 (N_15308,N_12295,N_13481);
xor U15309 (N_15309,N_13831,N_12647);
xnor U15310 (N_15310,N_12051,N_13356);
or U15311 (N_15311,N_13044,N_13837);
nor U15312 (N_15312,N_13187,N_13181);
and U15313 (N_15313,N_13466,N_12072);
and U15314 (N_15314,N_12926,N_13615);
and U15315 (N_15315,N_13173,N_12994);
or U15316 (N_15316,N_12257,N_12813);
nand U15317 (N_15317,N_12006,N_12611);
nor U15318 (N_15318,N_12724,N_12223);
xor U15319 (N_15319,N_13933,N_13492);
or U15320 (N_15320,N_13095,N_12465);
and U15321 (N_15321,N_13888,N_12455);
xnor U15322 (N_15322,N_12230,N_13237);
and U15323 (N_15323,N_12230,N_12585);
nand U15324 (N_15324,N_13848,N_12555);
nor U15325 (N_15325,N_12581,N_12736);
and U15326 (N_15326,N_13347,N_12251);
and U15327 (N_15327,N_13957,N_12180);
nor U15328 (N_15328,N_12664,N_13195);
xnor U15329 (N_15329,N_13245,N_12710);
and U15330 (N_15330,N_13152,N_12880);
and U15331 (N_15331,N_13473,N_12111);
and U15332 (N_15332,N_13329,N_13728);
or U15333 (N_15333,N_12418,N_12601);
nor U15334 (N_15334,N_13036,N_12885);
nor U15335 (N_15335,N_13188,N_13639);
or U15336 (N_15336,N_12326,N_13142);
nor U15337 (N_15337,N_12844,N_12355);
xnor U15338 (N_15338,N_13054,N_12418);
xnor U15339 (N_15339,N_13815,N_12021);
nor U15340 (N_15340,N_13245,N_13873);
nor U15341 (N_15341,N_13438,N_12008);
nand U15342 (N_15342,N_12569,N_12199);
xnor U15343 (N_15343,N_13061,N_12760);
nand U15344 (N_15344,N_13728,N_12953);
nand U15345 (N_15345,N_12719,N_13420);
nand U15346 (N_15346,N_12864,N_12038);
xnor U15347 (N_15347,N_13632,N_12505);
or U15348 (N_15348,N_13015,N_13030);
or U15349 (N_15349,N_12713,N_13835);
nor U15350 (N_15350,N_13971,N_12254);
or U15351 (N_15351,N_13183,N_12530);
and U15352 (N_15352,N_13134,N_12522);
and U15353 (N_15353,N_13876,N_13383);
nand U15354 (N_15354,N_13637,N_12073);
xor U15355 (N_15355,N_13605,N_12521);
and U15356 (N_15356,N_13649,N_12192);
nor U15357 (N_15357,N_13325,N_13697);
nand U15358 (N_15358,N_13588,N_12490);
xnor U15359 (N_15359,N_12745,N_13068);
or U15360 (N_15360,N_12789,N_12221);
and U15361 (N_15361,N_13261,N_13560);
nor U15362 (N_15362,N_13519,N_13745);
nor U15363 (N_15363,N_12047,N_13969);
or U15364 (N_15364,N_12852,N_13908);
or U15365 (N_15365,N_12210,N_13687);
nor U15366 (N_15366,N_13458,N_12522);
nand U15367 (N_15367,N_13569,N_12198);
and U15368 (N_15368,N_13161,N_13519);
or U15369 (N_15369,N_12091,N_12271);
or U15370 (N_15370,N_12608,N_13380);
nor U15371 (N_15371,N_12039,N_12820);
nand U15372 (N_15372,N_13984,N_13666);
nand U15373 (N_15373,N_13779,N_13576);
nand U15374 (N_15374,N_13070,N_12414);
and U15375 (N_15375,N_12693,N_13385);
and U15376 (N_15376,N_13188,N_12387);
nand U15377 (N_15377,N_13842,N_13015);
xor U15378 (N_15378,N_12904,N_13969);
or U15379 (N_15379,N_12963,N_13186);
nand U15380 (N_15380,N_12163,N_12453);
or U15381 (N_15381,N_13906,N_12045);
nand U15382 (N_15382,N_13841,N_13101);
or U15383 (N_15383,N_13608,N_12383);
nand U15384 (N_15384,N_13262,N_13816);
xor U15385 (N_15385,N_13717,N_13562);
and U15386 (N_15386,N_13592,N_12252);
xor U15387 (N_15387,N_12224,N_13505);
or U15388 (N_15388,N_13852,N_13181);
and U15389 (N_15389,N_13569,N_12862);
or U15390 (N_15390,N_13876,N_13943);
and U15391 (N_15391,N_12272,N_12868);
nand U15392 (N_15392,N_13597,N_13960);
or U15393 (N_15393,N_13660,N_12432);
xor U15394 (N_15394,N_12061,N_13413);
nand U15395 (N_15395,N_13029,N_12779);
xor U15396 (N_15396,N_13838,N_13631);
nand U15397 (N_15397,N_13035,N_12410);
and U15398 (N_15398,N_12625,N_13483);
and U15399 (N_15399,N_13958,N_12364);
or U15400 (N_15400,N_12960,N_13653);
or U15401 (N_15401,N_12121,N_12756);
and U15402 (N_15402,N_13787,N_12990);
and U15403 (N_15403,N_12427,N_12838);
xor U15404 (N_15404,N_12308,N_12268);
and U15405 (N_15405,N_12764,N_13999);
and U15406 (N_15406,N_13780,N_13513);
or U15407 (N_15407,N_13325,N_13715);
and U15408 (N_15408,N_12458,N_13468);
xor U15409 (N_15409,N_12165,N_13756);
or U15410 (N_15410,N_12463,N_13811);
and U15411 (N_15411,N_12562,N_13673);
and U15412 (N_15412,N_13040,N_13067);
nor U15413 (N_15413,N_12325,N_13587);
and U15414 (N_15414,N_12051,N_13900);
and U15415 (N_15415,N_13822,N_12819);
and U15416 (N_15416,N_12592,N_12290);
and U15417 (N_15417,N_12816,N_13335);
nor U15418 (N_15418,N_12127,N_13828);
or U15419 (N_15419,N_13160,N_13132);
or U15420 (N_15420,N_12958,N_13793);
nor U15421 (N_15421,N_13361,N_12819);
xor U15422 (N_15422,N_13374,N_13556);
xnor U15423 (N_15423,N_13534,N_12354);
nor U15424 (N_15424,N_13723,N_12034);
or U15425 (N_15425,N_12753,N_13603);
or U15426 (N_15426,N_13444,N_12746);
xnor U15427 (N_15427,N_12688,N_13655);
nor U15428 (N_15428,N_12877,N_13410);
nor U15429 (N_15429,N_13434,N_13188);
or U15430 (N_15430,N_12594,N_13324);
or U15431 (N_15431,N_13753,N_12182);
or U15432 (N_15432,N_12867,N_13961);
nor U15433 (N_15433,N_13451,N_12594);
xnor U15434 (N_15434,N_12606,N_13547);
xnor U15435 (N_15435,N_13309,N_12505);
nand U15436 (N_15436,N_13637,N_12367);
and U15437 (N_15437,N_13415,N_12564);
and U15438 (N_15438,N_13883,N_13763);
xor U15439 (N_15439,N_13521,N_12228);
and U15440 (N_15440,N_13740,N_13805);
and U15441 (N_15441,N_12292,N_12858);
and U15442 (N_15442,N_13760,N_12312);
nor U15443 (N_15443,N_12723,N_13048);
and U15444 (N_15444,N_12484,N_12158);
and U15445 (N_15445,N_13507,N_13000);
xor U15446 (N_15446,N_13914,N_13122);
nand U15447 (N_15447,N_12269,N_12418);
and U15448 (N_15448,N_13235,N_13058);
and U15449 (N_15449,N_12994,N_12884);
xnor U15450 (N_15450,N_13633,N_12620);
nand U15451 (N_15451,N_13805,N_12026);
or U15452 (N_15452,N_12382,N_12874);
and U15453 (N_15453,N_13774,N_12004);
nand U15454 (N_15454,N_12884,N_13775);
xnor U15455 (N_15455,N_12129,N_12052);
nand U15456 (N_15456,N_12505,N_12135);
xnor U15457 (N_15457,N_13167,N_12968);
and U15458 (N_15458,N_13171,N_13808);
xnor U15459 (N_15459,N_12003,N_13541);
or U15460 (N_15460,N_12557,N_13016);
nand U15461 (N_15461,N_12440,N_13154);
and U15462 (N_15462,N_13707,N_13380);
nor U15463 (N_15463,N_12582,N_12418);
or U15464 (N_15464,N_13932,N_12969);
and U15465 (N_15465,N_13904,N_12734);
nand U15466 (N_15466,N_12473,N_12600);
nand U15467 (N_15467,N_13439,N_13659);
and U15468 (N_15468,N_13934,N_13897);
xor U15469 (N_15469,N_12738,N_13500);
or U15470 (N_15470,N_12364,N_12110);
xnor U15471 (N_15471,N_13134,N_13785);
nand U15472 (N_15472,N_13896,N_13883);
or U15473 (N_15473,N_13094,N_12615);
or U15474 (N_15474,N_13000,N_12486);
nand U15475 (N_15475,N_12530,N_12431);
or U15476 (N_15476,N_13063,N_13569);
xnor U15477 (N_15477,N_12791,N_12608);
or U15478 (N_15478,N_12801,N_12970);
nor U15479 (N_15479,N_13513,N_13494);
xnor U15480 (N_15480,N_12949,N_13378);
nor U15481 (N_15481,N_13190,N_13106);
and U15482 (N_15482,N_12776,N_12491);
nand U15483 (N_15483,N_12987,N_13289);
and U15484 (N_15484,N_13278,N_12618);
xor U15485 (N_15485,N_13257,N_12045);
or U15486 (N_15486,N_12995,N_12319);
and U15487 (N_15487,N_13775,N_12792);
nand U15488 (N_15488,N_12815,N_12471);
nand U15489 (N_15489,N_12883,N_12024);
or U15490 (N_15490,N_13658,N_13790);
xnor U15491 (N_15491,N_13098,N_12028);
nor U15492 (N_15492,N_12502,N_12361);
or U15493 (N_15493,N_12161,N_13331);
or U15494 (N_15494,N_12523,N_13839);
or U15495 (N_15495,N_12859,N_13320);
nand U15496 (N_15496,N_13552,N_12636);
and U15497 (N_15497,N_13706,N_12862);
nand U15498 (N_15498,N_13390,N_13184);
and U15499 (N_15499,N_13307,N_12853);
nor U15500 (N_15500,N_12507,N_12838);
or U15501 (N_15501,N_13423,N_12991);
nor U15502 (N_15502,N_13777,N_13926);
nand U15503 (N_15503,N_13513,N_12194);
and U15504 (N_15504,N_13901,N_13097);
and U15505 (N_15505,N_13083,N_12576);
xor U15506 (N_15506,N_12094,N_12350);
or U15507 (N_15507,N_12726,N_13050);
nand U15508 (N_15508,N_12308,N_13095);
xnor U15509 (N_15509,N_13359,N_12215);
and U15510 (N_15510,N_12868,N_12973);
and U15511 (N_15511,N_12863,N_13652);
nand U15512 (N_15512,N_12104,N_13546);
xnor U15513 (N_15513,N_12203,N_13478);
and U15514 (N_15514,N_13790,N_12797);
or U15515 (N_15515,N_13174,N_12286);
or U15516 (N_15516,N_12839,N_13409);
nand U15517 (N_15517,N_13526,N_12294);
nand U15518 (N_15518,N_12295,N_13410);
nor U15519 (N_15519,N_12349,N_13271);
or U15520 (N_15520,N_13490,N_12384);
nor U15521 (N_15521,N_13881,N_13530);
nand U15522 (N_15522,N_13890,N_12170);
or U15523 (N_15523,N_13106,N_13012);
xor U15524 (N_15524,N_12185,N_13285);
nor U15525 (N_15525,N_13605,N_12286);
or U15526 (N_15526,N_12878,N_12103);
nand U15527 (N_15527,N_13492,N_12750);
nand U15528 (N_15528,N_13082,N_12147);
nand U15529 (N_15529,N_12415,N_12335);
xnor U15530 (N_15530,N_13887,N_12904);
xor U15531 (N_15531,N_13436,N_13891);
nand U15532 (N_15532,N_13282,N_13196);
nand U15533 (N_15533,N_12056,N_13180);
or U15534 (N_15534,N_12528,N_12621);
nand U15535 (N_15535,N_13876,N_12932);
and U15536 (N_15536,N_13893,N_13475);
nor U15537 (N_15537,N_13344,N_13564);
nor U15538 (N_15538,N_12595,N_12206);
or U15539 (N_15539,N_13979,N_12095);
nand U15540 (N_15540,N_12323,N_13777);
xnor U15541 (N_15541,N_12373,N_12183);
nor U15542 (N_15542,N_13547,N_13024);
nand U15543 (N_15543,N_13139,N_12386);
xor U15544 (N_15544,N_13280,N_13113);
or U15545 (N_15545,N_12241,N_12680);
nand U15546 (N_15546,N_13489,N_12793);
or U15547 (N_15547,N_12040,N_12715);
xor U15548 (N_15548,N_12313,N_12746);
and U15549 (N_15549,N_12568,N_13316);
and U15550 (N_15550,N_12547,N_12662);
or U15551 (N_15551,N_13377,N_12836);
xnor U15552 (N_15552,N_13050,N_13061);
nor U15553 (N_15553,N_12655,N_13077);
xnor U15554 (N_15554,N_13089,N_12752);
nand U15555 (N_15555,N_13882,N_13598);
or U15556 (N_15556,N_12334,N_12878);
nor U15557 (N_15557,N_12057,N_13665);
and U15558 (N_15558,N_13749,N_13018);
nand U15559 (N_15559,N_13398,N_12848);
or U15560 (N_15560,N_12294,N_13480);
and U15561 (N_15561,N_12722,N_13992);
and U15562 (N_15562,N_13774,N_13739);
or U15563 (N_15563,N_13152,N_12243);
xor U15564 (N_15564,N_13378,N_12414);
xnor U15565 (N_15565,N_12801,N_12900);
or U15566 (N_15566,N_12537,N_12816);
nor U15567 (N_15567,N_13454,N_12355);
or U15568 (N_15568,N_13307,N_13437);
nor U15569 (N_15569,N_13351,N_13872);
nor U15570 (N_15570,N_12268,N_13264);
and U15571 (N_15571,N_12920,N_12708);
nor U15572 (N_15572,N_12259,N_12764);
xnor U15573 (N_15573,N_13785,N_12954);
and U15574 (N_15574,N_12604,N_13066);
nor U15575 (N_15575,N_13735,N_13361);
or U15576 (N_15576,N_12435,N_13519);
xor U15577 (N_15577,N_13536,N_13411);
nor U15578 (N_15578,N_12610,N_12794);
nand U15579 (N_15579,N_12790,N_13805);
xnor U15580 (N_15580,N_12755,N_12870);
or U15581 (N_15581,N_13237,N_13393);
or U15582 (N_15582,N_12005,N_13511);
or U15583 (N_15583,N_12802,N_13863);
and U15584 (N_15584,N_12462,N_13397);
xor U15585 (N_15585,N_12000,N_12834);
and U15586 (N_15586,N_13917,N_13881);
or U15587 (N_15587,N_13219,N_13905);
xnor U15588 (N_15588,N_12582,N_12719);
or U15589 (N_15589,N_13566,N_13010);
and U15590 (N_15590,N_13101,N_13934);
and U15591 (N_15591,N_13578,N_13155);
nand U15592 (N_15592,N_12395,N_12259);
nor U15593 (N_15593,N_13890,N_13749);
nand U15594 (N_15594,N_12980,N_12784);
nand U15595 (N_15595,N_13732,N_13591);
nand U15596 (N_15596,N_13417,N_12244);
xor U15597 (N_15597,N_12607,N_13137);
and U15598 (N_15598,N_13816,N_13349);
and U15599 (N_15599,N_12708,N_13459);
nor U15600 (N_15600,N_12695,N_12197);
or U15601 (N_15601,N_13779,N_13507);
nand U15602 (N_15602,N_12259,N_13629);
or U15603 (N_15603,N_13426,N_12048);
xor U15604 (N_15604,N_13437,N_13732);
nand U15605 (N_15605,N_12718,N_13218);
and U15606 (N_15606,N_13359,N_13746);
and U15607 (N_15607,N_12694,N_12447);
nand U15608 (N_15608,N_12764,N_12839);
xnor U15609 (N_15609,N_12612,N_12831);
and U15610 (N_15610,N_13247,N_12318);
xnor U15611 (N_15611,N_13850,N_12613);
nor U15612 (N_15612,N_12295,N_12792);
nand U15613 (N_15613,N_13223,N_13135);
and U15614 (N_15614,N_12172,N_12555);
nand U15615 (N_15615,N_12972,N_13126);
nand U15616 (N_15616,N_13178,N_13270);
or U15617 (N_15617,N_13340,N_12363);
nor U15618 (N_15618,N_13593,N_13774);
xnor U15619 (N_15619,N_12170,N_12951);
nand U15620 (N_15620,N_12485,N_12854);
and U15621 (N_15621,N_13798,N_13144);
or U15622 (N_15622,N_13440,N_12327);
and U15623 (N_15623,N_12463,N_12484);
xnor U15624 (N_15624,N_13554,N_12038);
and U15625 (N_15625,N_13570,N_12263);
and U15626 (N_15626,N_13554,N_13391);
or U15627 (N_15627,N_13533,N_13758);
or U15628 (N_15628,N_13172,N_12685);
or U15629 (N_15629,N_13311,N_12342);
or U15630 (N_15630,N_13307,N_13585);
nor U15631 (N_15631,N_13855,N_12309);
nand U15632 (N_15632,N_12032,N_12534);
and U15633 (N_15633,N_12755,N_13317);
xnor U15634 (N_15634,N_13643,N_12287);
xnor U15635 (N_15635,N_12242,N_13595);
nor U15636 (N_15636,N_13132,N_12869);
xnor U15637 (N_15637,N_12700,N_12655);
xnor U15638 (N_15638,N_12876,N_12839);
or U15639 (N_15639,N_13002,N_12794);
xnor U15640 (N_15640,N_12423,N_12493);
nand U15641 (N_15641,N_12071,N_12139);
nand U15642 (N_15642,N_13131,N_13559);
or U15643 (N_15643,N_12786,N_12850);
xnor U15644 (N_15644,N_12442,N_12925);
nor U15645 (N_15645,N_13449,N_13679);
nor U15646 (N_15646,N_12483,N_13281);
nand U15647 (N_15647,N_13328,N_13464);
and U15648 (N_15648,N_12922,N_13559);
and U15649 (N_15649,N_12815,N_13406);
or U15650 (N_15650,N_13391,N_13164);
and U15651 (N_15651,N_13541,N_13110);
nor U15652 (N_15652,N_12242,N_12256);
and U15653 (N_15653,N_12646,N_13820);
nand U15654 (N_15654,N_13850,N_13858);
or U15655 (N_15655,N_13296,N_12190);
or U15656 (N_15656,N_13314,N_12838);
nor U15657 (N_15657,N_13100,N_13720);
nor U15658 (N_15658,N_12944,N_12923);
or U15659 (N_15659,N_13653,N_12514);
xnor U15660 (N_15660,N_13013,N_13328);
xnor U15661 (N_15661,N_13871,N_13335);
nor U15662 (N_15662,N_13294,N_12097);
or U15663 (N_15663,N_13287,N_12054);
and U15664 (N_15664,N_12972,N_12196);
nand U15665 (N_15665,N_13725,N_13503);
nand U15666 (N_15666,N_13660,N_12706);
nand U15667 (N_15667,N_12724,N_12980);
nand U15668 (N_15668,N_13043,N_13525);
nand U15669 (N_15669,N_13616,N_12104);
nor U15670 (N_15670,N_12601,N_13220);
xor U15671 (N_15671,N_13336,N_12822);
and U15672 (N_15672,N_12044,N_12455);
nor U15673 (N_15673,N_12584,N_12655);
or U15674 (N_15674,N_13276,N_12393);
nor U15675 (N_15675,N_13062,N_13663);
nand U15676 (N_15676,N_12959,N_13784);
or U15677 (N_15677,N_13917,N_12280);
nand U15678 (N_15678,N_13869,N_13297);
nand U15679 (N_15679,N_12029,N_13111);
and U15680 (N_15680,N_12003,N_12258);
nand U15681 (N_15681,N_13398,N_12430);
nor U15682 (N_15682,N_13753,N_13337);
or U15683 (N_15683,N_12122,N_12140);
xor U15684 (N_15684,N_12260,N_13953);
and U15685 (N_15685,N_12436,N_12764);
or U15686 (N_15686,N_12891,N_13062);
nor U15687 (N_15687,N_12287,N_13368);
nor U15688 (N_15688,N_12985,N_12911);
and U15689 (N_15689,N_13763,N_13992);
and U15690 (N_15690,N_12232,N_12482);
or U15691 (N_15691,N_12553,N_13992);
nand U15692 (N_15692,N_12800,N_12069);
nand U15693 (N_15693,N_13606,N_12534);
nor U15694 (N_15694,N_12001,N_13868);
nand U15695 (N_15695,N_13480,N_13344);
nand U15696 (N_15696,N_12951,N_13985);
xnor U15697 (N_15697,N_13019,N_12507);
and U15698 (N_15698,N_12926,N_13786);
xor U15699 (N_15699,N_13440,N_13442);
nor U15700 (N_15700,N_12310,N_13422);
and U15701 (N_15701,N_13583,N_13645);
or U15702 (N_15702,N_12330,N_13264);
and U15703 (N_15703,N_13303,N_13672);
and U15704 (N_15704,N_12960,N_12445);
or U15705 (N_15705,N_13407,N_12949);
or U15706 (N_15706,N_12690,N_13936);
nand U15707 (N_15707,N_13913,N_13478);
or U15708 (N_15708,N_13545,N_13519);
and U15709 (N_15709,N_13667,N_12778);
nor U15710 (N_15710,N_12842,N_13846);
nand U15711 (N_15711,N_13147,N_13934);
nand U15712 (N_15712,N_13520,N_12226);
or U15713 (N_15713,N_12694,N_13360);
and U15714 (N_15714,N_12574,N_12515);
nand U15715 (N_15715,N_13042,N_12039);
xor U15716 (N_15716,N_12140,N_12653);
or U15717 (N_15717,N_13276,N_13261);
or U15718 (N_15718,N_12789,N_12204);
or U15719 (N_15719,N_12043,N_12598);
xor U15720 (N_15720,N_13840,N_13517);
or U15721 (N_15721,N_13611,N_12852);
nand U15722 (N_15722,N_13454,N_13123);
nor U15723 (N_15723,N_13685,N_12799);
xor U15724 (N_15724,N_12016,N_12600);
nand U15725 (N_15725,N_13141,N_13990);
and U15726 (N_15726,N_12002,N_12278);
or U15727 (N_15727,N_12213,N_12108);
xor U15728 (N_15728,N_12877,N_12274);
nand U15729 (N_15729,N_12134,N_12940);
nor U15730 (N_15730,N_13947,N_13653);
or U15731 (N_15731,N_13475,N_13391);
nand U15732 (N_15732,N_13575,N_13877);
xor U15733 (N_15733,N_12765,N_12897);
xnor U15734 (N_15734,N_12207,N_13997);
and U15735 (N_15735,N_13274,N_13680);
xnor U15736 (N_15736,N_12869,N_12770);
and U15737 (N_15737,N_12463,N_12776);
xnor U15738 (N_15738,N_12866,N_13854);
or U15739 (N_15739,N_13933,N_13943);
xor U15740 (N_15740,N_12786,N_13109);
nand U15741 (N_15741,N_13065,N_12575);
and U15742 (N_15742,N_13682,N_13176);
and U15743 (N_15743,N_12086,N_13150);
xnor U15744 (N_15744,N_13936,N_13392);
or U15745 (N_15745,N_13570,N_13825);
nand U15746 (N_15746,N_12767,N_12429);
and U15747 (N_15747,N_13537,N_12600);
nor U15748 (N_15748,N_12984,N_13914);
nor U15749 (N_15749,N_13200,N_12324);
and U15750 (N_15750,N_13700,N_12185);
and U15751 (N_15751,N_13470,N_13939);
nor U15752 (N_15752,N_13674,N_13770);
xor U15753 (N_15753,N_13031,N_12834);
and U15754 (N_15754,N_12357,N_13323);
nand U15755 (N_15755,N_12215,N_13351);
nor U15756 (N_15756,N_12377,N_13872);
nand U15757 (N_15757,N_13498,N_12608);
nand U15758 (N_15758,N_13283,N_12204);
and U15759 (N_15759,N_13833,N_12852);
or U15760 (N_15760,N_13996,N_12968);
nor U15761 (N_15761,N_12972,N_12355);
and U15762 (N_15762,N_12898,N_13488);
nor U15763 (N_15763,N_12016,N_12250);
nand U15764 (N_15764,N_12945,N_13570);
and U15765 (N_15765,N_12491,N_13947);
nand U15766 (N_15766,N_13657,N_12953);
xnor U15767 (N_15767,N_12283,N_12954);
xnor U15768 (N_15768,N_12070,N_12288);
nand U15769 (N_15769,N_13803,N_13425);
xnor U15770 (N_15770,N_12046,N_12396);
and U15771 (N_15771,N_12739,N_12956);
or U15772 (N_15772,N_12290,N_12873);
and U15773 (N_15773,N_12772,N_13844);
nor U15774 (N_15774,N_12176,N_12423);
xor U15775 (N_15775,N_13081,N_12819);
xor U15776 (N_15776,N_12453,N_12925);
or U15777 (N_15777,N_12690,N_13950);
and U15778 (N_15778,N_12939,N_12716);
or U15779 (N_15779,N_12101,N_12288);
and U15780 (N_15780,N_12226,N_12153);
or U15781 (N_15781,N_13358,N_13985);
nor U15782 (N_15782,N_12521,N_13188);
nand U15783 (N_15783,N_12760,N_12834);
and U15784 (N_15784,N_12885,N_13331);
and U15785 (N_15785,N_12601,N_12584);
xor U15786 (N_15786,N_13680,N_12871);
nor U15787 (N_15787,N_13335,N_13853);
nor U15788 (N_15788,N_12569,N_13089);
and U15789 (N_15789,N_13567,N_13799);
xor U15790 (N_15790,N_13764,N_12936);
nor U15791 (N_15791,N_12757,N_13141);
xnor U15792 (N_15792,N_12646,N_12697);
xor U15793 (N_15793,N_12350,N_12739);
or U15794 (N_15794,N_13117,N_12951);
nand U15795 (N_15795,N_12639,N_13144);
or U15796 (N_15796,N_12233,N_13844);
xor U15797 (N_15797,N_12841,N_13748);
or U15798 (N_15798,N_13356,N_12993);
xnor U15799 (N_15799,N_12765,N_13228);
xor U15800 (N_15800,N_12610,N_13533);
or U15801 (N_15801,N_12765,N_13490);
nand U15802 (N_15802,N_13249,N_13684);
and U15803 (N_15803,N_13509,N_12388);
nor U15804 (N_15804,N_12408,N_13387);
or U15805 (N_15805,N_13491,N_12290);
nand U15806 (N_15806,N_12906,N_13111);
nor U15807 (N_15807,N_13643,N_13806);
or U15808 (N_15808,N_12502,N_12342);
nand U15809 (N_15809,N_12522,N_13706);
and U15810 (N_15810,N_12545,N_13810);
or U15811 (N_15811,N_12472,N_12917);
or U15812 (N_15812,N_12803,N_13131);
xor U15813 (N_15813,N_12630,N_12120);
nand U15814 (N_15814,N_13706,N_13195);
nand U15815 (N_15815,N_12827,N_13164);
xnor U15816 (N_15816,N_12475,N_12902);
xor U15817 (N_15817,N_13617,N_12827);
and U15818 (N_15818,N_12036,N_12504);
or U15819 (N_15819,N_13084,N_12796);
nor U15820 (N_15820,N_13249,N_13487);
nor U15821 (N_15821,N_13048,N_12722);
nand U15822 (N_15822,N_12952,N_13839);
and U15823 (N_15823,N_13067,N_12353);
and U15824 (N_15824,N_13515,N_12077);
nor U15825 (N_15825,N_12822,N_13672);
nor U15826 (N_15826,N_13869,N_13130);
and U15827 (N_15827,N_13909,N_12790);
xor U15828 (N_15828,N_13909,N_13059);
nor U15829 (N_15829,N_12495,N_13632);
xnor U15830 (N_15830,N_12332,N_12666);
xor U15831 (N_15831,N_13735,N_13298);
or U15832 (N_15832,N_13942,N_13780);
xnor U15833 (N_15833,N_13855,N_12368);
or U15834 (N_15834,N_12977,N_13962);
or U15835 (N_15835,N_13098,N_12341);
nor U15836 (N_15836,N_12275,N_13288);
nand U15837 (N_15837,N_13854,N_13531);
xor U15838 (N_15838,N_12943,N_13690);
and U15839 (N_15839,N_13005,N_12006);
xnor U15840 (N_15840,N_13553,N_13602);
or U15841 (N_15841,N_12379,N_12217);
nand U15842 (N_15842,N_12574,N_13585);
or U15843 (N_15843,N_12656,N_13239);
or U15844 (N_15844,N_12888,N_12103);
nor U15845 (N_15845,N_12579,N_12493);
nor U15846 (N_15846,N_13398,N_13584);
or U15847 (N_15847,N_12392,N_13531);
or U15848 (N_15848,N_13577,N_12718);
nor U15849 (N_15849,N_13850,N_13574);
nand U15850 (N_15850,N_13944,N_12677);
or U15851 (N_15851,N_13976,N_12690);
nand U15852 (N_15852,N_13099,N_13422);
and U15853 (N_15853,N_12684,N_12589);
nand U15854 (N_15854,N_12542,N_12051);
xnor U15855 (N_15855,N_13682,N_12327);
and U15856 (N_15856,N_13862,N_13153);
or U15857 (N_15857,N_13735,N_13760);
and U15858 (N_15858,N_12431,N_13352);
nor U15859 (N_15859,N_13592,N_12577);
nand U15860 (N_15860,N_12275,N_13839);
nor U15861 (N_15861,N_12016,N_13883);
nor U15862 (N_15862,N_12346,N_13726);
nand U15863 (N_15863,N_13572,N_13079);
and U15864 (N_15864,N_13750,N_12963);
and U15865 (N_15865,N_13872,N_13506);
nand U15866 (N_15866,N_12739,N_12477);
nor U15867 (N_15867,N_13769,N_13542);
nand U15868 (N_15868,N_12517,N_13514);
xnor U15869 (N_15869,N_12653,N_13485);
xor U15870 (N_15870,N_12570,N_12080);
nand U15871 (N_15871,N_12800,N_12738);
or U15872 (N_15872,N_12844,N_12280);
and U15873 (N_15873,N_12853,N_13505);
or U15874 (N_15874,N_12376,N_12214);
nand U15875 (N_15875,N_13595,N_13187);
nor U15876 (N_15876,N_12213,N_13835);
xor U15877 (N_15877,N_13488,N_13385);
nor U15878 (N_15878,N_13108,N_12981);
or U15879 (N_15879,N_13478,N_12638);
and U15880 (N_15880,N_12242,N_13736);
and U15881 (N_15881,N_12818,N_12757);
xor U15882 (N_15882,N_13780,N_12588);
and U15883 (N_15883,N_13439,N_12302);
nor U15884 (N_15884,N_13197,N_12869);
xor U15885 (N_15885,N_13047,N_12259);
nor U15886 (N_15886,N_12293,N_12217);
and U15887 (N_15887,N_12518,N_12762);
xnor U15888 (N_15888,N_12939,N_12456);
nand U15889 (N_15889,N_13712,N_13266);
xor U15890 (N_15890,N_12851,N_13729);
xnor U15891 (N_15891,N_12156,N_13693);
or U15892 (N_15892,N_12869,N_13736);
and U15893 (N_15893,N_13700,N_12371);
and U15894 (N_15894,N_13447,N_13259);
nor U15895 (N_15895,N_13801,N_13013);
xnor U15896 (N_15896,N_12959,N_12742);
nand U15897 (N_15897,N_13032,N_13336);
and U15898 (N_15898,N_13696,N_13439);
xor U15899 (N_15899,N_13835,N_12917);
and U15900 (N_15900,N_13034,N_13265);
and U15901 (N_15901,N_12856,N_12548);
or U15902 (N_15902,N_13849,N_12889);
nand U15903 (N_15903,N_12022,N_12392);
or U15904 (N_15904,N_13687,N_12017);
xnor U15905 (N_15905,N_13340,N_13430);
or U15906 (N_15906,N_13638,N_13049);
nor U15907 (N_15907,N_13338,N_13307);
or U15908 (N_15908,N_12729,N_12442);
nor U15909 (N_15909,N_13173,N_13960);
nor U15910 (N_15910,N_12127,N_12542);
nor U15911 (N_15911,N_13690,N_13890);
nor U15912 (N_15912,N_13126,N_13838);
nand U15913 (N_15913,N_12747,N_12346);
xor U15914 (N_15914,N_12471,N_12449);
nand U15915 (N_15915,N_13390,N_13845);
xnor U15916 (N_15916,N_12110,N_13464);
nand U15917 (N_15917,N_12639,N_12431);
and U15918 (N_15918,N_12853,N_13503);
nor U15919 (N_15919,N_12804,N_13414);
or U15920 (N_15920,N_12635,N_13131);
xnor U15921 (N_15921,N_12511,N_12543);
or U15922 (N_15922,N_13951,N_12018);
xor U15923 (N_15923,N_13938,N_13404);
nand U15924 (N_15924,N_13070,N_12466);
xnor U15925 (N_15925,N_13555,N_13850);
nor U15926 (N_15926,N_12653,N_13336);
xnor U15927 (N_15927,N_12498,N_12082);
or U15928 (N_15928,N_13479,N_12395);
xor U15929 (N_15929,N_12610,N_12719);
or U15930 (N_15930,N_12820,N_13986);
or U15931 (N_15931,N_12607,N_12692);
or U15932 (N_15932,N_12672,N_12791);
xor U15933 (N_15933,N_12105,N_12242);
nand U15934 (N_15934,N_12939,N_12331);
xor U15935 (N_15935,N_13401,N_12728);
nand U15936 (N_15936,N_12376,N_13403);
and U15937 (N_15937,N_12372,N_12567);
nor U15938 (N_15938,N_13130,N_12892);
xnor U15939 (N_15939,N_13361,N_13979);
nand U15940 (N_15940,N_12236,N_13497);
xnor U15941 (N_15941,N_13362,N_13314);
nor U15942 (N_15942,N_12665,N_12619);
or U15943 (N_15943,N_12529,N_12116);
nor U15944 (N_15944,N_12870,N_13329);
nand U15945 (N_15945,N_12785,N_12689);
and U15946 (N_15946,N_12151,N_12107);
xor U15947 (N_15947,N_12459,N_12833);
or U15948 (N_15948,N_13580,N_12946);
and U15949 (N_15949,N_13516,N_13448);
xnor U15950 (N_15950,N_12646,N_13305);
nor U15951 (N_15951,N_13313,N_13971);
nor U15952 (N_15952,N_12120,N_13246);
nand U15953 (N_15953,N_13679,N_13234);
nand U15954 (N_15954,N_13018,N_13244);
and U15955 (N_15955,N_12930,N_12887);
xnor U15956 (N_15956,N_12938,N_13233);
nand U15957 (N_15957,N_12619,N_13020);
and U15958 (N_15958,N_12869,N_13420);
xnor U15959 (N_15959,N_13471,N_13978);
nor U15960 (N_15960,N_13711,N_12174);
nor U15961 (N_15961,N_13112,N_13337);
or U15962 (N_15962,N_12237,N_12348);
nor U15963 (N_15963,N_13521,N_13091);
nor U15964 (N_15964,N_13413,N_13989);
nor U15965 (N_15965,N_13405,N_12819);
xor U15966 (N_15966,N_13697,N_13590);
nor U15967 (N_15967,N_12571,N_12903);
xnor U15968 (N_15968,N_13303,N_13707);
or U15969 (N_15969,N_12055,N_13789);
nor U15970 (N_15970,N_12368,N_13369);
and U15971 (N_15971,N_12484,N_12721);
or U15972 (N_15972,N_13487,N_13355);
or U15973 (N_15973,N_13809,N_12541);
or U15974 (N_15974,N_12204,N_12092);
or U15975 (N_15975,N_13930,N_12664);
nand U15976 (N_15976,N_13456,N_12544);
or U15977 (N_15977,N_13629,N_13937);
xnor U15978 (N_15978,N_12021,N_13091);
or U15979 (N_15979,N_13324,N_13961);
or U15980 (N_15980,N_13473,N_13725);
nor U15981 (N_15981,N_13477,N_12584);
xor U15982 (N_15982,N_12500,N_13292);
or U15983 (N_15983,N_13867,N_12440);
and U15984 (N_15984,N_13937,N_12003);
and U15985 (N_15985,N_13052,N_13280);
or U15986 (N_15986,N_13022,N_13345);
xor U15987 (N_15987,N_12419,N_12301);
xnor U15988 (N_15988,N_12170,N_12835);
nor U15989 (N_15989,N_12509,N_12629);
nor U15990 (N_15990,N_12810,N_13889);
nor U15991 (N_15991,N_13375,N_12253);
nand U15992 (N_15992,N_12983,N_13380);
nand U15993 (N_15993,N_12214,N_12494);
nand U15994 (N_15994,N_12946,N_13560);
nand U15995 (N_15995,N_13315,N_12389);
xor U15996 (N_15996,N_13986,N_13247);
xor U15997 (N_15997,N_12463,N_12103);
nor U15998 (N_15998,N_13178,N_12587);
or U15999 (N_15999,N_12120,N_12108);
or U16000 (N_16000,N_14375,N_15822);
nor U16001 (N_16001,N_14574,N_14676);
nor U16002 (N_16002,N_14209,N_14718);
or U16003 (N_16003,N_15940,N_15254);
xnor U16004 (N_16004,N_15406,N_14990);
nor U16005 (N_16005,N_14808,N_14492);
nor U16006 (N_16006,N_14138,N_15531);
nor U16007 (N_16007,N_15325,N_15123);
xnor U16008 (N_16008,N_15943,N_15681);
or U16009 (N_16009,N_14053,N_14128);
xor U16010 (N_16010,N_15608,N_14343);
or U16011 (N_16011,N_14979,N_15557);
nand U16012 (N_16012,N_15138,N_15604);
nor U16013 (N_16013,N_14806,N_15274);
nor U16014 (N_16014,N_14988,N_15830);
and U16015 (N_16015,N_15964,N_14126);
nor U16016 (N_16016,N_14899,N_14028);
xnor U16017 (N_16017,N_15602,N_15414);
xor U16018 (N_16018,N_14940,N_14578);
or U16019 (N_16019,N_15308,N_15927);
nor U16020 (N_16020,N_14432,N_14660);
nand U16021 (N_16021,N_15579,N_15051);
xnor U16022 (N_16022,N_15412,N_15311);
and U16023 (N_16023,N_14233,N_15529);
nor U16024 (N_16024,N_15615,N_15566);
nor U16025 (N_16025,N_14112,N_15097);
nand U16026 (N_16026,N_14405,N_15721);
nor U16027 (N_16027,N_15072,N_15585);
xor U16028 (N_16028,N_14282,N_14687);
nand U16029 (N_16029,N_15955,N_15399);
xnor U16030 (N_16030,N_14524,N_15278);
nand U16031 (N_16031,N_15786,N_14843);
nor U16032 (N_16032,N_14333,N_15185);
and U16033 (N_16033,N_14096,N_14707);
and U16034 (N_16034,N_14228,N_15977);
nand U16035 (N_16035,N_15680,N_14819);
nand U16036 (N_16036,N_15963,N_15860);
and U16037 (N_16037,N_14728,N_14294);
or U16038 (N_16038,N_14370,N_14244);
nor U16039 (N_16039,N_15332,N_14188);
xnor U16040 (N_16040,N_15926,N_14602);
nor U16041 (N_16041,N_14266,N_15990);
and U16042 (N_16042,N_15347,N_14727);
nor U16043 (N_16043,N_14224,N_15104);
and U16044 (N_16044,N_15280,N_14065);
nand U16045 (N_16045,N_15191,N_14450);
xnor U16046 (N_16046,N_15416,N_15288);
nand U16047 (N_16047,N_15142,N_14299);
nand U16048 (N_16048,N_15059,N_15112);
or U16049 (N_16049,N_15451,N_14541);
and U16050 (N_16050,N_15887,N_15912);
nand U16051 (N_16051,N_15540,N_14336);
nand U16052 (N_16052,N_14166,N_14378);
or U16053 (N_16053,N_15544,N_14879);
or U16054 (N_16054,N_14841,N_15891);
nand U16055 (N_16055,N_15477,N_15530);
nor U16056 (N_16056,N_15390,N_15918);
and U16057 (N_16057,N_14621,N_14555);
or U16058 (N_16058,N_14009,N_15302);
xnor U16059 (N_16059,N_15473,N_14110);
nand U16060 (N_16060,N_14323,N_15485);
nor U16061 (N_16061,N_14793,N_14455);
nand U16062 (N_16062,N_14335,N_14840);
and U16063 (N_16063,N_15453,N_14208);
nand U16064 (N_16064,N_15182,N_15813);
or U16065 (N_16065,N_14436,N_15016);
xnor U16066 (N_16066,N_15994,N_14195);
nor U16067 (N_16067,N_15386,N_15703);
nand U16068 (N_16068,N_15210,N_15186);
or U16069 (N_16069,N_15641,N_14585);
or U16070 (N_16070,N_14024,N_14225);
xnor U16071 (N_16071,N_14365,N_15944);
nor U16072 (N_16072,N_15082,N_14174);
and U16073 (N_16073,N_14035,N_14157);
xor U16074 (N_16074,N_15591,N_15146);
and U16075 (N_16075,N_14963,N_14387);
and U16076 (N_16076,N_14094,N_14172);
xnor U16077 (N_16077,N_14736,N_15486);
nor U16078 (N_16078,N_15304,N_14263);
and U16079 (N_16079,N_15455,N_14501);
nand U16080 (N_16080,N_15610,N_15915);
and U16081 (N_16081,N_14640,N_15581);
and U16082 (N_16082,N_15647,N_14362);
nor U16083 (N_16083,N_15179,N_15770);
and U16084 (N_16084,N_15193,N_15756);
or U16085 (N_16085,N_15420,N_15046);
and U16086 (N_16086,N_15835,N_14962);
or U16087 (N_16087,N_15925,N_15656);
or U16088 (N_16088,N_14137,N_15003);
nand U16089 (N_16089,N_15374,N_15783);
xnor U16090 (N_16090,N_14748,N_14120);
nand U16091 (N_16091,N_15518,N_15643);
xor U16092 (N_16092,N_14192,N_14489);
xor U16093 (N_16093,N_14904,N_15144);
and U16094 (N_16094,N_14567,N_14632);
xor U16095 (N_16095,N_15836,N_14477);
and U16096 (N_16096,N_14042,N_14264);
xor U16097 (N_16097,N_15899,N_15755);
and U16098 (N_16098,N_15221,N_14101);
or U16099 (N_16099,N_15165,N_15659);
nand U16100 (N_16100,N_14245,N_15991);
xor U16101 (N_16101,N_15778,N_14831);
nor U16102 (N_16102,N_14587,N_14597);
nor U16103 (N_16103,N_15364,N_15825);
nand U16104 (N_16104,N_14794,N_15381);
xnor U16105 (N_16105,N_15238,N_15969);
or U16106 (N_16106,N_15653,N_15949);
and U16107 (N_16107,N_15058,N_15597);
nor U16108 (N_16108,N_14629,N_14685);
nor U16109 (N_16109,N_15978,N_14625);
xor U16110 (N_16110,N_14402,N_14221);
nor U16111 (N_16111,N_15404,N_15303);
nor U16112 (N_16112,N_15872,N_14022);
nand U16113 (N_16113,N_15468,N_14865);
or U16114 (N_16114,N_15295,N_14826);
nand U16115 (N_16115,N_15137,N_14784);
nand U16116 (N_16116,N_14770,N_15898);
nand U16117 (N_16117,N_14662,N_15605);
nand U16118 (N_16118,N_14124,N_15296);
xnor U16119 (N_16119,N_14652,N_15574);
nor U16120 (N_16120,N_15411,N_15121);
xnor U16121 (N_16121,N_14945,N_14534);
or U16122 (N_16122,N_15299,N_15110);
xor U16123 (N_16123,N_15713,N_14134);
and U16124 (N_16124,N_14683,N_15122);
nand U16125 (N_16125,N_15514,N_14372);
xor U16126 (N_16126,N_15795,N_14003);
or U16127 (N_16127,N_15229,N_14763);
nor U16128 (N_16128,N_14733,N_15619);
and U16129 (N_16129,N_14371,N_14391);
nand U16130 (N_16130,N_14158,N_14705);
or U16131 (N_16131,N_15556,N_14497);
nand U16132 (N_16132,N_14358,N_14435);
and U16133 (N_16133,N_15388,N_15446);
and U16134 (N_16134,N_15230,N_14251);
nor U16135 (N_16135,N_15108,N_15312);
and U16136 (N_16136,N_15538,N_15373);
and U16137 (N_16137,N_15508,N_15471);
xor U16138 (N_16138,N_15673,N_15816);
and U16139 (N_16139,N_14440,N_14952);
nand U16140 (N_16140,N_15131,N_14661);
nor U16141 (N_16141,N_15054,N_14599);
nor U16142 (N_16142,N_15031,N_15043);
or U16143 (N_16143,N_15157,N_14173);
nand U16144 (N_16144,N_15310,N_14059);
and U16145 (N_16145,N_14725,N_15655);
or U16146 (N_16146,N_15202,N_15617);
nand U16147 (N_16147,N_15164,N_14563);
nand U16148 (N_16148,N_15194,N_14605);
xnor U16149 (N_16149,N_14400,N_14752);
or U16150 (N_16150,N_14768,N_15358);
or U16151 (N_16151,N_15021,N_14889);
nand U16152 (N_16152,N_14229,N_15959);
nand U16153 (N_16153,N_14293,N_15090);
or U16154 (N_16154,N_14697,N_14778);
nand U16155 (N_16155,N_14056,N_15953);
xor U16156 (N_16156,N_14617,N_14993);
and U16157 (N_16157,N_15539,N_15187);
nand U16158 (N_16158,N_14050,N_14906);
or U16159 (N_16159,N_15433,N_14189);
nor U16160 (N_16160,N_15751,N_15675);
and U16161 (N_16161,N_14301,N_15847);
nand U16162 (N_16162,N_15981,N_14551);
xnor U16163 (N_16163,N_14797,N_15839);
and U16164 (N_16164,N_15845,N_14956);
nor U16165 (N_16165,N_15988,N_14711);
nand U16166 (N_16166,N_15309,N_14849);
nand U16167 (N_16167,N_15070,N_15056);
or U16168 (N_16168,N_14407,N_15710);
or U16169 (N_16169,N_14423,N_15008);
xnor U16170 (N_16170,N_14890,N_14769);
nor U16171 (N_16171,N_14891,N_14483);
and U16172 (N_16172,N_15793,N_14898);
nor U16173 (N_16173,N_15287,N_15026);
nand U16174 (N_16174,N_14029,N_15078);
nand U16175 (N_16175,N_15668,N_14925);
and U16176 (N_16176,N_15985,N_15984);
and U16177 (N_16177,N_14399,N_15696);
nand U16178 (N_16178,N_15626,N_15178);
nor U16179 (N_16179,N_14242,N_14720);
nor U16180 (N_16180,N_14281,N_14951);
nand U16181 (N_16181,N_15419,N_15598);
xor U16182 (N_16182,N_14329,N_14084);
or U16183 (N_16183,N_14033,N_15161);
or U16184 (N_16184,N_15725,N_15007);
or U16185 (N_16185,N_14047,N_15478);
nand U16186 (N_16186,N_14664,N_15039);
and U16187 (N_16187,N_14085,N_15498);
and U16188 (N_16188,N_14976,N_15063);
or U16189 (N_16189,N_15867,N_15688);
and U16190 (N_16190,N_14820,N_14066);
and U16191 (N_16191,N_15812,N_15649);
nand U16192 (N_16192,N_15614,N_14967);
xor U16193 (N_16193,N_14352,N_15520);
xor U16194 (N_16194,N_15245,N_14917);
nand U16195 (N_16195,N_14448,N_14417);
and U16196 (N_16196,N_14751,N_14971);
or U16197 (N_16197,N_15428,N_15938);
nand U16198 (N_16198,N_15004,N_14508);
or U16199 (N_16199,N_15041,N_15997);
and U16200 (N_16200,N_15716,N_14918);
nor U16201 (N_16201,N_15865,N_14321);
or U16202 (N_16202,N_14255,N_15513);
xor U16203 (N_16203,N_15177,N_14610);
nor U16204 (N_16204,N_15960,N_15686);
nand U16205 (N_16205,N_14929,N_15425);
nor U16206 (N_16206,N_15341,N_15805);
or U16207 (N_16207,N_14213,N_14064);
xnor U16208 (N_16208,N_15521,N_14558);
and U16209 (N_16209,N_14862,N_14493);
nand U16210 (N_16210,N_14550,N_15741);
and U16211 (N_16211,N_14291,N_15447);
and U16212 (N_16212,N_15038,N_15583);
xor U16213 (N_16213,N_14108,N_15732);
nand U16214 (N_16214,N_15140,N_14284);
xor U16215 (N_16215,N_15558,N_15316);
xnor U16216 (N_16216,N_14430,N_15369);
nand U16217 (N_16217,N_15424,N_15678);
or U16218 (N_16218,N_15523,N_14637);
nor U16219 (N_16219,N_15223,N_15698);
xor U16220 (N_16220,N_15661,N_14735);
or U16221 (N_16221,N_14876,N_15754);
nor U16222 (N_16222,N_14783,N_14915);
nand U16223 (N_16223,N_14606,N_15742);
or U16224 (N_16224,N_15166,N_14256);
xor U16225 (N_16225,N_14133,N_15875);
xor U16226 (N_16226,N_14207,N_14027);
and U16227 (N_16227,N_15774,N_15149);
nor U16228 (N_16228,N_14782,N_14471);
nor U16229 (N_16229,N_15706,N_15017);
and U16230 (N_16230,N_15378,N_14531);
nand U16231 (N_16231,N_15219,N_15737);
or U16232 (N_16232,N_15368,N_15248);
xor U16233 (N_16233,N_14373,N_15705);
and U16234 (N_16234,N_15509,N_14756);
or U16235 (N_16235,N_15993,N_15375);
nand U16236 (N_16236,N_15240,N_15376);
xor U16237 (N_16237,N_14626,N_15359);
xnor U16238 (N_16238,N_14877,N_15027);
nor U16239 (N_16239,N_15427,N_14540);
xnor U16240 (N_16240,N_14590,N_14422);
xnor U16241 (N_16241,N_14892,N_15200);
and U16242 (N_16242,N_15232,N_15336);
and U16243 (N_16243,N_14360,N_14986);
and U16244 (N_16244,N_14746,N_15644);
nand U16245 (N_16245,N_14475,N_15268);
and U16246 (N_16246,N_14351,N_14203);
or U16247 (N_16247,N_15844,N_15738);
nor U16248 (N_16248,N_15061,N_14647);
and U16249 (N_16249,N_15169,N_14342);
nor U16250 (N_16250,N_15565,N_14595);
nand U16251 (N_16251,N_14528,N_14267);
nor U16252 (N_16252,N_14071,N_14686);
xor U16253 (N_16253,N_15115,N_15136);
nand U16254 (N_16254,N_14655,N_15854);
nand U16255 (N_16255,N_15151,N_14468);
and U16256 (N_16256,N_14445,N_15707);
nor U16257 (N_16257,N_15951,N_14943);
and U16258 (N_16258,N_15467,N_15664);
nor U16259 (N_16259,N_15630,N_14488);
and U16260 (N_16260,N_14757,N_14178);
and U16261 (N_16261,N_15018,N_15189);
nand U16262 (N_16262,N_14562,N_14609);
nand U16263 (N_16263,N_14845,N_14583);
xor U16264 (N_16264,N_14818,N_14216);
nor U16265 (N_16265,N_14078,N_14368);
and U16266 (N_16266,N_15904,N_14013);
nand U16267 (N_16267,N_14506,N_15559);
and U16268 (N_16268,N_14165,N_14579);
and U16269 (N_16269,N_15492,N_15073);
or U16270 (N_16270,N_15005,N_15129);
nor U16271 (N_16271,N_14830,N_14914);
or U16272 (N_16272,N_14616,N_15040);
or U16273 (N_16273,N_15444,N_15265);
and U16274 (N_16274,N_14187,N_15249);
xnor U16275 (N_16275,N_15636,N_14045);
xnor U16276 (N_16276,N_15134,N_14996);
nor U16277 (N_16277,N_14260,N_14775);
nor U16278 (N_16278,N_14498,N_14090);
nor U16279 (N_16279,N_14667,N_15118);
or U16280 (N_16280,N_14153,N_15128);
and U16281 (N_16281,N_14582,N_15360);
xnor U16282 (N_16282,N_15011,N_15517);
and U16283 (N_16283,N_14999,N_14997);
xnor U16284 (N_16284,N_15768,N_14779);
xor U16285 (N_16285,N_14302,N_14023);
nor U16286 (N_16286,N_14103,N_15549);
or U16287 (N_16287,N_14600,N_14331);
nor U16288 (N_16288,N_14960,N_15057);
or U16289 (N_16289,N_14622,N_15727);
or U16290 (N_16290,N_14349,N_14886);
xor U16291 (N_16291,N_15799,N_14011);
and U16292 (N_16292,N_15633,N_14995);
xnor U16293 (N_16293,N_14088,N_15717);
or U16294 (N_16294,N_14312,N_15398);
nand U16295 (N_16295,N_14116,N_15474);
or U16296 (N_16296,N_14314,N_14543);
nor U16297 (N_16297,N_14481,N_14984);
or U16298 (N_16298,N_15297,N_15000);
xor U16299 (N_16299,N_14320,N_14571);
nor U16300 (N_16300,N_15315,N_15580);
xnor U16301 (N_16301,N_14656,N_15113);
xor U16302 (N_16302,N_14082,N_14535);
nand U16303 (N_16303,N_14955,N_15323);
and U16304 (N_16304,N_15366,N_14604);
nand U16305 (N_16305,N_14888,N_14451);
nor U16306 (N_16306,N_15116,N_15470);
nand U16307 (N_16307,N_14798,N_14791);
xnor U16308 (N_16308,N_14805,N_15820);
nand U16309 (N_16309,N_14220,N_14449);
or U16310 (N_16310,N_14698,N_14796);
and U16311 (N_16311,N_14992,N_14125);
nand U16312 (N_16312,N_15015,N_15338);
xor U16313 (N_16313,N_14815,N_14893);
nor U16314 (N_16314,N_14810,N_14322);
or U16315 (N_16315,N_14525,N_14223);
nor U16316 (N_16316,N_15667,N_14714);
or U16317 (N_16317,N_14395,N_14139);
nand U16318 (N_16318,N_15127,N_14415);
and U16319 (N_16319,N_15334,N_14470);
and U16320 (N_16320,N_14480,N_14318);
or U16321 (N_16321,N_14016,N_14901);
or U16322 (N_16322,N_14953,N_14202);
nand U16323 (N_16323,N_14874,N_15462);
xor U16324 (N_16324,N_15241,N_15395);
and U16325 (N_16325,N_15772,N_15036);
and U16326 (N_16326,N_15109,N_14719);
nand U16327 (N_16327,N_15159,N_15083);
xor U16328 (N_16328,N_14485,N_15807);
nor U16329 (N_16329,N_14106,N_14265);
xnor U16330 (N_16330,N_14944,N_15196);
or U16331 (N_16331,N_15851,N_15266);
or U16332 (N_16332,N_15009,N_15394);
nand U16333 (N_16333,N_14743,N_15937);
or U16334 (N_16334,N_14392,N_14019);
and U16335 (N_16335,N_15611,N_15607);
nand U16336 (N_16336,N_14717,N_15947);
nand U16337 (N_16337,N_14026,N_14155);
nor U16338 (N_16338,N_14337,N_14315);
xnor U16339 (N_16339,N_14749,N_15354);
xor U16340 (N_16340,N_15685,N_15212);
and U16341 (N_16341,N_15117,N_14650);
and U16342 (N_16342,N_15924,N_15679);
and U16343 (N_16343,N_14482,N_15405);
or U16344 (N_16344,N_14277,N_14691);
and U16345 (N_16345,N_14427,N_15261);
or U16346 (N_16346,N_14347,N_15989);
xnor U16347 (N_16347,N_15651,N_14846);
xor U16348 (N_16348,N_15576,N_15689);
nor U16349 (N_16349,N_14121,N_15568);
or U16350 (N_16350,N_14708,N_14665);
nor U16351 (N_16351,N_14644,N_14657);
xnor U16352 (N_16352,N_15400,N_15488);
and U16353 (N_16353,N_15349,N_14693);
nand U16354 (N_16354,N_15283,N_14651);
or U16355 (N_16355,N_15760,N_15735);
nor U16356 (N_16356,N_14290,N_14142);
or U16357 (N_16357,N_14565,N_15570);
xor U16358 (N_16358,N_15044,N_15501);
nand U16359 (N_16359,N_15533,N_15372);
xnor U16360 (N_16360,N_14150,N_15234);
xor U16361 (N_16361,N_14416,N_14222);
nor U16362 (N_16362,N_15101,N_15790);
nand U16363 (N_16363,N_15069,N_15880);
xnor U16364 (N_16364,N_14308,N_14702);
and U16365 (N_16365,N_14473,N_14215);
xnor U16366 (N_16366,N_14152,N_15060);
xnor U16367 (N_16367,N_15857,N_14135);
nor U16368 (N_16368,N_15817,N_15763);
xor U16369 (N_16369,N_14273,N_14713);
nor U16370 (N_16370,N_14658,N_15806);
and U16371 (N_16371,N_14589,N_15652);
xor U16372 (N_16372,N_14038,N_14077);
nor U16373 (N_16373,N_14390,N_15328);
xnor U16374 (N_16374,N_14759,N_15019);
nor U16375 (N_16375,N_15171,N_15983);
nor U16376 (N_16376,N_15764,N_15147);
xnor U16377 (N_16377,N_14409,N_15236);
nor U16378 (N_16378,N_15827,N_14678);
and U16379 (N_16379,N_15257,N_15148);
xor U16380 (N_16380,N_15337,N_15911);
nand U16381 (N_16381,N_15356,N_14792);
or U16382 (N_16382,N_14032,N_15638);
nor U16383 (N_16383,N_15826,N_14734);
and U16384 (N_16384,N_15033,N_15259);
and U16385 (N_16385,N_14092,N_15423);
nand U16386 (N_16386,N_15824,N_14210);
xor U16387 (N_16387,N_15049,N_15849);
nand U16388 (N_16388,N_15114,N_15294);
nand U16389 (N_16389,N_14146,N_15535);
xor U16390 (N_16390,N_15671,N_14460);
and U16391 (N_16391,N_15702,N_14109);
and U16392 (N_16392,N_14654,N_14307);
nand U16393 (N_16393,N_14408,N_15340);
or U16394 (N_16394,N_14700,N_15396);
nor U16395 (N_16395,N_15749,N_14389);
xnor U16396 (N_16396,N_14067,N_15237);
xor U16397 (N_16397,N_14183,N_15465);
or U16398 (N_16398,N_14348,N_14633);
nor U16399 (N_16399,N_15645,N_15861);
or U16400 (N_16400,N_15906,N_15639);
nand U16401 (N_16401,N_15589,N_15204);
nor U16402 (N_16402,N_15298,N_14978);
and U16403 (N_16403,N_14051,N_14628);
nand U16404 (N_16404,N_14154,N_14823);
or U16405 (N_16405,N_15184,N_14227);
and U16406 (N_16406,N_15603,N_15869);
or U16407 (N_16407,N_14296,N_14547);
nand U16408 (N_16408,N_15582,N_15174);
nand U16409 (N_16409,N_15543,N_15883);
nor U16410 (N_16410,N_15350,N_14570);
xnor U16411 (N_16411,N_15222,N_15318);
nor U16412 (N_16412,N_15495,N_14802);
or U16413 (N_16413,N_14167,N_15107);
and U16414 (N_16414,N_15279,N_14706);
nor U16415 (N_16415,N_14428,N_15690);
and U16416 (N_16416,N_15901,N_14184);
and U16417 (N_16417,N_15413,N_14036);
nand U16418 (N_16418,N_14684,N_14297);
nor U16419 (N_16419,N_14552,N_15491);
and U16420 (N_16420,N_15479,N_15874);
or U16421 (N_16421,N_14958,N_15469);
nand U16422 (N_16422,N_15804,N_15214);
and U16423 (N_16423,N_14837,N_15065);
or U16424 (N_16424,N_14504,N_14847);
nand U16425 (N_16425,N_14515,N_15519);
nor U16426 (N_16426,N_15648,N_14758);
nor U16427 (N_16427,N_15028,N_14766);
or U16428 (N_16428,N_14382,N_14959);
or U16429 (N_16429,N_14828,N_15348);
nand U16430 (N_16430,N_15272,N_15343);
nand U16431 (N_16431,N_14271,N_15052);
xor U16432 (N_16432,N_15313,N_14780);
nand U16433 (N_16433,N_14316,N_14008);
nor U16434 (N_16434,N_14283,N_15974);
nand U16435 (N_16435,N_14093,N_14194);
nand U16436 (N_16436,N_14377,N_14231);
nor U16437 (N_16437,N_14040,N_15393);
or U16438 (N_16438,N_15440,N_15956);
or U16439 (N_16439,N_15666,N_15970);
or U16440 (N_16440,N_15885,N_14932);
or U16441 (N_16441,N_14669,N_14095);
or U16442 (N_16442,N_14860,N_15216);
nor U16443 (N_16443,N_15429,N_14080);
nand U16444 (N_16444,N_14285,N_14479);
nand U16445 (N_16445,N_14429,N_15119);
nand U16446 (N_16446,N_15600,N_15946);
and U16447 (N_16447,N_15683,N_15892);
nand U16448 (N_16448,N_15934,N_15578);
xor U16449 (N_16449,N_14068,N_15198);
nand U16450 (N_16450,N_14197,N_15014);
nor U16451 (N_16451,N_15551,N_15766);
xor U16452 (N_16452,N_14406,N_14058);
nor U16453 (N_16453,N_14253,N_15842);
or U16454 (N_16454,N_14868,N_14801);
or U16455 (N_16455,N_15852,N_15153);
or U16456 (N_16456,N_15840,N_15418);
or U16457 (N_16457,N_14396,N_14279);
or U16458 (N_16458,N_15629,N_15720);
nor U16459 (N_16459,N_14760,N_15595);
xnor U16460 (N_16460,N_15935,N_15919);
nand U16461 (N_16461,N_14044,N_14894);
and U16462 (N_16462,N_15162,N_15777);
nor U16463 (N_16463,N_15506,N_14907);
xor U16464 (N_16464,N_15802,N_14981);
or U16465 (N_16465,N_14190,N_14920);
nor U16466 (N_16466,N_15239,N_15493);
nor U16467 (N_16467,N_14006,N_15357);
nor U16468 (N_16468,N_14612,N_15922);
or U16469 (N_16469,N_14864,N_14141);
and U16470 (N_16470,N_15695,N_15961);
and U16471 (N_16471,N_14624,N_15663);
or U16472 (N_16472,N_14062,N_14467);
or U16473 (N_16473,N_14593,N_14105);
nand U16474 (N_16474,N_15168,N_14715);
or U16475 (N_16475,N_15289,N_15837);
xnor U16476 (N_16476,N_15782,N_15436);
and U16477 (N_16477,N_14274,N_15227);
and U16478 (N_16478,N_15628,N_15654);
or U16479 (N_16479,N_14014,N_14364);
nand U16480 (N_16480,N_15715,N_15814);
or U16481 (N_16481,N_14672,N_14747);
nor U16482 (N_16482,N_14186,N_14179);
and U16483 (N_16483,N_14458,N_15389);
nor U16484 (N_16484,N_14356,N_15800);
xnor U16485 (N_16485,N_15561,N_15750);
nand U16486 (N_16486,N_14511,N_15285);
and U16487 (N_16487,N_15281,N_14638);
or U16488 (N_16488,N_14086,N_15532);
or U16489 (N_16489,N_14544,N_14731);
or U16490 (N_16490,N_15577,N_15862);
xnor U16491 (N_16491,N_14131,N_15733);
xnor U16492 (N_16492,N_14611,N_14645);
or U16493 (N_16493,N_15554,N_15346);
xor U16494 (N_16494,N_14034,N_14677);
xnor U16495 (N_16495,N_14942,N_14114);
and U16496 (N_16496,N_15599,N_14198);
and U16497 (N_16497,N_15331,N_15693);
nor U16498 (N_16498,N_14581,N_15461);
nand U16499 (N_16499,N_14568,N_15012);
and U16500 (N_16500,N_14304,N_14286);
or U16501 (N_16501,N_14910,N_14829);
nor U16502 (N_16502,N_14924,N_14520);
and U16503 (N_16503,N_15753,N_15260);
and U16504 (N_16504,N_14816,N_15900);
nand U16505 (N_16505,N_14326,N_15913);
nand U16506 (N_16506,N_14873,N_14682);
nor U16507 (N_16507,N_15062,N_14834);
or U16508 (N_16508,N_14002,N_15256);
and U16509 (N_16509,N_15030,N_14262);
or U16510 (N_16510,N_15291,N_14259);
xnor U16511 (N_16511,N_14973,N_14140);
and U16512 (N_16512,N_15077,N_15392);
and U16513 (N_16513,N_15454,N_15660);
nand U16514 (N_16514,N_15430,N_14836);
nor U16515 (N_16515,N_14113,N_15320);
xnor U16516 (N_16516,N_14319,N_14446);
and U16517 (N_16517,N_15377,N_14902);
or U16518 (N_16518,N_15371,N_15625);
nor U16519 (N_16519,N_14909,N_14908);
and U16520 (N_16520,N_14694,N_14037);
xnor U16521 (N_16521,N_15843,N_15743);
nand U16522 (N_16522,N_14098,N_14170);
xnor U16523 (N_16523,N_14217,N_15697);
xnor U16524 (N_16524,N_14355,N_15088);
or U16525 (N_16525,N_15801,N_15475);
nand U16526 (N_16526,N_15546,N_14591);
and U16527 (N_16527,N_15096,N_15572);
xor U16528 (N_16528,N_15275,N_14171);
and U16529 (N_16529,N_14017,N_15013);
nor U16530 (N_16530,N_14418,N_14376);
or U16531 (N_16531,N_14755,N_15457);
nor U16532 (N_16532,N_14619,N_14168);
nor U16533 (N_16533,N_14539,N_15409);
or U16534 (N_16534,N_15868,N_15158);
nand U16535 (N_16535,N_15718,N_14148);
nor U16536 (N_16536,N_14021,N_14887);
nor U16537 (N_16537,N_14311,N_14772);
nor U16538 (N_16538,N_14239,N_15794);
or U16539 (N_16539,N_15143,N_14921);
nand U16540 (N_16540,N_15658,N_14313);
xnor U16541 (N_16541,N_14767,N_14070);
or U16542 (N_16542,N_14374,N_14247);
or U16543 (N_16543,N_14659,N_15086);
nand U16544 (N_16544,N_14452,N_15258);
and U16545 (N_16545,N_15367,N_14526);
xor U16546 (N_16546,N_15779,N_14413);
nor U16547 (N_16547,N_14839,N_14099);
nor U16548 (N_16548,N_15687,N_15821);
xnor U16549 (N_16549,N_14922,N_14969);
xor U16550 (N_16550,N_15352,N_15780);
xor U16551 (N_16551,N_14310,N_14761);
and U16552 (N_16552,N_14903,N_14900);
or U16553 (N_16553,N_15719,N_14627);
nor U16554 (N_16554,N_14275,N_15456);
xor U16555 (N_16555,N_15255,N_14254);
and U16556 (N_16556,N_15226,N_14030);
nor U16557 (N_16557,N_15512,N_14704);
and U16558 (N_16558,N_14936,N_14000);
and U16559 (N_16559,N_15575,N_15646);
nand U16560 (N_16560,N_15798,N_15293);
nand U16561 (N_16561,N_14938,N_14433);
nor U16562 (N_16562,N_15307,N_14964);
and U16563 (N_16563,N_15075,N_14776);
nor U16564 (N_16564,N_15933,N_15677);
xnor U16565 (N_16565,N_15384,N_14856);
nor U16566 (N_16566,N_14001,N_15966);
or U16567 (N_16567,N_14895,N_15522);
and U16568 (N_16568,N_15130,N_14821);
nor U16569 (N_16569,N_14218,N_14057);
xor U16570 (N_16570,N_15879,N_14673);
or U16571 (N_16571,N_14557,N_14989);
and U16572 (N_16572,N_14235,N_14773);
nand U16573 (N_16573,N_15081,N_14982);
nor U16574 (N_16574,N_14248,N_15435);
or U16575 (N_16575,N_14164,N_14340);
and U16576 (N_16576,N_15220,N_15276);
and U16577 (N_16577,N_15776,N_15103);
xnor U16578 (N_16578,N_14151,N_15884);
and U16579 (N_16579,N_14814,N_14354);
or U16580 (N_16580,N_14205,N_15618);
xor U16581 (N_16581,N_14569,N_14510);
nand U16582 (N_16582,N_15206,N_14043);
and U16583 (N_16583,N_15550,N_14100);
and U16584 (N_16584,N_14598,N_14919);
nor U16585 (N_16585,N_15034,N_15606);
or U16586 (N_16586,N_14330,N_14507);
and U16587 (N_16587,N_15167,N_14073);
and U16588 (N_16588,N_15306,N_14201);
and U16589 (N_16589,N_14812,N_14670);
nor U16590 (N_16590,N_14401,N_14974);
nor U16591 (N_16591,N_15642,N_15023);
nor U16592 (N_16592,N_15132,N_15785);
nand U16593 (N_16593,N_15620,N_14144);
or U16594 (N_16594,N_15330,N_15890);
and U16595 (N_16595,N_14411,N_14542);
or U16596 (N_16596,N_15897,N_15333);
and U16597 (N_16597,N_14811,N_14160);
and U16598 (N_16598,N_14803,N_15180);
xnor U16599 (N_16599,N_14465,N_14442);
xnor U16600 (N_16600,N_14346,N_15269);
and U16601 (N_16601,N_14663,N_15909);
and U16602 (N_16602,N_14463,N_15560);
xnor U16603 (N_16603,N_14980,N_15277);
and U16604 (N_16604,N_15124,N_15841);
and U16605 (N_16605,N_15907,N_15211);
nor U16606 (N_16606,N_14384,N_15421);
nor U16607 (N_16607,N_15945,N_14353);
nand U16608 (N_16608,N_14857,N_15908);
nor U16609 (N_16609,N_14175,N_15921);
nor U16610 (N_16610,N_14118,N_15536);
and U16611 (N_16611,N_14785,N_15045);
nand U16612 (N_16612,N_14339,N_14513);
nor U16613 (N_16613,N_15100,N_15431);
and U16614 (N_16614,N_14545,N_14226);
and U16615 (N_16615,N_15920,N_14709);
nand U16616 (N_16616,N_15452,N_15744);
or U16617 (N_16617,N_15590,N_15809);
nor U16618 (N_16618,N_15002,N_14270);
or U16619 (N_16619,N_14863,N_14977);
nor U16620 (N_16620,N_14437,N_15476);
xnor U16621 (N_16621,N_15627,N_14466);
xor U16622 (N_16622,N_14443,N_15672);
nor U16623 (N_16623,N_15218,N_14858);
nand U16624 (N_16624,N_14985,N_15724);
or U16625 (N_16625,N_14494,N_15192);
nand U16626 (N_16626,N_14212,N_15301);
or U16627 (N_16627,N_14844,N_15877);
nand U16628 (N_16628,N_14722,N_14012);
and U16629 (N_16629,N_15541,N_14854);
xor U16630 (N_16630,N_15609,N_15442);
and U16631 (N_16631,N_15999,N_14199);
nand U16632 (N_16632,N_14147,N_15723);
nor U16633 (N_16633,N_15329,N_15850);
and U16634 (N_16634,N_14338,N_15207);
nand U16635 (N_16635,N_15502,N_14393);
or U16636 (N_16636,N_15950,N_15071);
xor U16637 (N_16637,N_14268,N_15217);
nor U16638 (N_16638,N_15889,N_14586);
nor U16639 (N_16639,N_14699,N_14607);
xnor U16640 (N_16640,N_15437,N_15537);
nor U16641 (N_16641,N_14935,N_15699);
xor U16642 (N_16642,N_15593,N_14232);
nand U16643 (N_16643,N_15781,N_14580);
xnor U16644 (N_16644,N_15387,N_15982);
nor U16645 (N_16645,N_15484,N_14824);
nor U16646 (N_16646,N_14076,N_15525);
xnor U16647 (N_16647,N_15767,N_14957);
xor U16648 (N_16648,N_14983,N_15853);
nor U16649 (N_16649,N_14278,N_15032);
nor U16650 (N_16650,N_14419,N_15832);
nand U16651 (N_16651,N_14642,N_14643);
nor U16652 (N_16652,N_14257,N_15111);
and U16653 (N_16653,N_15976,N_14514);
and U16654 (N_16654,N_14991,N_15251);
xor U16655 (N_16655,N_14527,N_15209);
and U16656 (N_16656,N_15942,N_15569);
nand U16657 (N_16657,N_14689,N_15024);
xnor U16658 (N_16658,N_14025,N_14789);
and U16659 (N_16659,N_15657,N_15747);
xnor U16660 (N_16660,N_14970,N_15682);
nor U16661 (N_16661,N_14937,N_15722);
nor U16662 (N_16662,N_14237,N_14548);
nand U16663 (N_16663,N_15006,N_14115);
and U16664 (N_16664,N_15391,N_15466);
xnor U16665 (N_16665,N_15480,N_14870);
nor U16666 (N_16666,N_15001,N_15510);
and U16667 (N_16667,N_15962,N_14518);
xor U16668 (N_16668,N_14556,N_15759);
or U16669 (N_16669,N_14911,N_14532);
and U16670 (N_16670,N_14363,N_14750);
nor U16671 (N_16671,N_15588,N_15856);
nand U16672 (N_16672,N_14441,N_14156);
nor U16673 (N_16673,N_15321,N_14679);
or U16674 (N_16674,N_14359,N_14288);
or U16675 (N_16675,N_14309,N_14939);
or U16676 (N_16676,N_15385,N_15818);
and U16677 (N_16677,N_15235,N_15085);
nand U16678 (N_16678,N_14594,N_14947);
nand U16679 (N_16679,N_15120,N_14478);
nand U16680 (N_16680,N_14464,N_14741);
xor U16681 (N_16681,N_15995,N_15992);
xor U16682 (N_16682,N_14072,N_15730);
and U16683 (N_16683,N_14883,N_15203);
nand U16684 (N_16684,N_14905,N_14739);
xnor U16685 (N_16685,N_14149,N_15106);
xor U16686 (N_16686,N_14380,N_15224);
nand U16687 (N_16687,N_15172,N_15215);
nor U16688 (N_16688,N_15758,N_15035);
nor U16689 (N_16689,N_15098,N_14852);
nor U16690 (N_16690,N_15160,N_14204);
xnor U16691 (N_16691,N_15383,N_14869);
nand U16692 (N_16692,N_14069,N_15838);
or U16693 (N_16693,N_14280,N_15201);
or U16694 (N_16694,N_14630,N_15434);
nand U16695 (N_16695,N_15213,N_15662);
nor U16696 (N_16696,N_15464,N_15634);
xnor U16697 (N_16697,N_14738,N_15930);
xnor U16698 (N_16698,N_14397,N_15928);
and U16699 (N_16699,N_15397,N_14934);
or U16700 (N_16700,N_14822,N_14817);
xnor U16701 (N_16701,N_15552,N_15326);
xor U16702 (N_16702,N_14063,N_15534);
nor U16703 (N_16703,N_14180,N_15048);
xor U16704 (N_16704,N_15286,N_15050);
xor U16705 (N_16705,N_14079,N_14649);
nand U16706 (N_16706,N_14007,N_15916);
nor U16707 (N_16707,N_15902,N_15370);
xnor U16708 (N_16708,N_14447,N_14102);
or U16709 (N_16709,N_14258,N_15426);
nand U16710 (N_16710,N_15833,N_14505);
nand U16711 (N_16711,N_15365,N_14087);
nor U16712 (N_16712,N_14136,N_14795);
nor U16713 (N_16713,N_15882,N_14601);
or U16714 (N_16714,N_14383,N_15761);
and U16715 (N_16715,N_15823,N_14117);
and U16716 (N_16716,N_14648,N_15528);
nor U16717 (N_16717,N_14701,N_15270);
nand U16718 (N_16718,N_14787,N_14615);
xor U16719 (N_16719,N_14564,N_14074);
nor U16720 (N_16720,N_14219,N_15936);
nor U16721 (N_16721,N_15505,N_15594);
and U16722 (N_16722,N_14425,N_14182);
nand U16723 (N_16723,N_15954,N_14762);
xnor U16724 (N_16724,N_14523,N_15573);
or U16725 (N_16725,N_15152,N_15562);
nand U16726 (N_16726,N_15066,N_14623);
and U16727 (N_16727,N_14196,N_14703);
or U16728 (N_16728,N_15622,N_14306);
or U16729 (N_16729,N_14931,N_14412);
or U16730 (N_16730,N_15866,N_14809);
xnor U16731 (N_16731,N_14366,N_14529);
xor U16732 (N_16732,N_15345,N_14521);
nand U16733 (N_16733,N_15621,N_15472);
and U16734 (N_16734,N_15975,N_15601);
or U16735 (N_16735,N_15410,N_14692);
and U16736 (N_16736,N_15709,N_14386);
xnor U16737 (N_16737,N_14054,N_14462);
xnor U16738 (N_16738,N_14049,N_15815);
xor U16739 (N_16739,N_15190,N_14031);
xnor U16740 (N_16740,N_15403,N_15834);
xnor U16741 (N_16741,N_15731,N_14777);
or U16742 (N_16742,N_14075,N_14575);
nor U16743 (N_16743,N_14716,N_15163);
nand U16744 (N_16744,N_15704,N_15787);
and U16745 (N_16745,N_15154,N_14424);
and U16746 (N_16746,N_15351,N_14538);
nor U16747 (N_16747,N_15155,N_14896);
xnor U16748 (N_16748,N_14833,N_14410);
xnor U16749 (N_16749,N_15613,N_15415);
xor U16750 (N_16750,N_15917,N_15941);
nand U16751 (N_16751,N_14674,N_15339);
xor U16752 (N_16752,N_14261,N_14123);
or U16753 (N_16753,N_14861,N_14191);
nor U16754 (N_16754,N_14832,N_14853);
or U16755 (N_16755,N_15923,N_15871);
nand U16756 (N_16756,N_14132,N_14954);
nor U16757 (N_16757,N_15811,N_14882);
nand U16758 (N_16758,N_15752,N_15091);
nor U16759 (N_16759,N_15150,N_15527);
xor U16760 (N_16760,N_15361,N_14827);
nor U16761 (N_16761,N_15612,N_15745);
or U16762 (N_16762,N_14554,N_15076);
and U16763 (N_16763,N_15099,N_14866);
nand U16764 (N_16764,N_14799,N_15188);
nand U16765 (N_16765,N_15439,N_15487);
xnor U16766 (N_16766,N_14576,N_14723);
nand U16767 (N_16767,N_15762,N_15511);
or U16768 (N_16768,N_14252,N_15504);
and U16769 (N_16769,N_15126,N_15483);
nor U16770 (N_16770,N_15555,N_15445);
and U16771 (N_16771,N_15692,N_14913);
or U16772 (N_16772,N_15973,N_14324);
xor U16773 (N_16773,N_14091,N_14737);
nand U16774 (N_16774,N_14681,N_15135);
or U16775 (N_16775,N_14603,N_15788);
xnor U16776 (N_16776,N_15789,N_14675);
and U16777 (N_16777,N_14438,N_14842);
xor U16778 (N_16778,N_15499,N_14414);
nand U16779 (N_16779,N_14696,N_15181);
and U16780 (N_16780,N_15886,N_14459);
nand U16781 (N_16781,N_15064,N_14193);
nand U16782 (N_16782,N_15791,N_15979);
nand U16783 (N_16783,N_14546,N_15775);
nand U16784 (N_16784,N_15500,N_14474);
xor U16785 (N_16785,N_14439,N_15967);
nor U16786 (N_16786,N_15183,N_14020);
or U16787 (N_16787,N_14653,N_14420);
and U16788 (N_16788,N_15490,N_15986);
nand U16789 (N_16789,N_15449,N_14941);
nand U16790 (N_16790,N_14048,N_15773);
nor U16791 (N_16791,N_14145,N_14461);
xnor U16792 (N_16792,N_14491,N_15362);
nor U16793 (N_16793,N_15247,N_15864);
and U16794 (N_16794,N_14350,N_14859);
and U16795 (N_16795,N_14965,N_14503);
nand U16796 (N_16796,N_14041,N_14200);
nand U16797 (N_16797,N_14159,N_15665);
and U16798 (N_16798,N_15708,N_14848);
or U16799 (N_16799,N_15564,N_14710);
and U16800 (N_16800,N_15547,N_14129);
xor U16801 (N_16801,N_15829,N_15881);
xnor U16802 (N_16802,N_14246,N_15765);
xor U16803 (N_16803,N_14881,N_14754);
xor U16804 (N_16804,N_14453,N_14305);
xor U16805 (N_16805,N_14484,N_15380);
and U16806 (N_16806,N_15587,N_15463);
and U16807 (N_16807,N_15342,N_14851);
nor U16808 (N_16808,N_15105,N_15586);
xor U16809 (N_16809,N_14553,N_15896);
nor U16810 (N_16810,N_15089,N_14249);
nand U16811 (N_16811,N_14712,N_14972);
xor U16812 (N_16812,N_14403,N_15087);
and U16813 (N_16813,N_15176,N_14998);
and U16814 (N_16814,N_15173,N_14083);
and U16815 (N_16815,N_15243,N_15624);
xnor U16816 (N_16816,N_15074,N_15740);
nor U16817 (N_16817,N_14061,N_14897);
nor U16818 (N_16818,N_15448,N_15417);
or U16819 (N_16819,N_14269,N_15910);
and U16820 (N_16820,N_15092,N_15141);
nor U16821 (N_16821,N_15402,N_15769);
and U16822 (N_16822,N_14052,N_15355);
and U16823 (N_16823,N_14444,N_15873);
nor U16824 (N_16824,N_14588,N_14549);
and U16825 (N_16825,N_15808,N_14688);
and U16826 (N_16826,N_15273,N_15503);
nand U16827 (N_16827,N_15596,N_15526);
nor U16828 (N_16828,N_15810,N_15637);
nor U16829 (N_16829,N_14388,N_14015);
and U16830 (N_16830,N_14169,N_15831);
nor U16831 (N_16831,N_14163,N_14512);
nand U16832 (N_16832,N_15327,N_15407);
nand U16833 (N_16833,N_14671,N_15025);
nor U16834 (N_16834,N_14838,N_15819);
nand U16835 (N_16835,N_15441,N_15987);
and U16836 (N_16836,N_14634,N_14618);
nand U16837 (N_16837,N_15670,N_14162);
nand U16838 (N_16838,N_15694,N_15623);
nand U16839 (N_16839,N_14317,N_14695);
or U16840 (N_16840,N_15079,N_15497);
xor U16841 (N_16841,N_15952,N_14039);
or U16842 (N_16842,N_14369,N_15481);
and U16843 (N_16843,N_14537,N_15567);
or U16844 (N_16844,N_15729,N_14010);
or U16845 (N_16845,N_14005,N_14740);
xnor U16846 (N_16846,N_15282,N_15010);
nor U16847 (N_16847,N_15746,N_14379);
or U16848 (N_16848,N_15996,N_14499);
xor U16849 (N_16849,N_14875,N_14680);
nand U16850 (N_16850,N_14298,N_15632);
nand U16851 (N_16851,N_14303,N_14788);
and U16852 (N_16852,N_15635,N_15968);
nor U16853 (N_16853,N_14790,N_14122);
nand U16854 (N_16854,N_15205,N_14398);
xnor U16855 (N_16855,N_15542,N_15691);
nand U16856 (N_16856,N_15084,N_14111);
nor U16857 (N_16857,N_14885,N_15631);
and U16858 (N_16858,N_14107,N_14835);
nand U16859 (N_16859,N_15322,N_15401);
nand U16860 (N_16860,N_14850,N_15545);
or U16861 (N_16861,N_15460,N_15208);
or U16862 (N_16862,N_15971,N_15080);
xnor U16863 (N_16863,N_15870,N_14855);
xnor U16864 (N_16864,N_15888,N_15711);
and U16865 (N_16865,N_14272,N_15878);
or U16866 (N_16866,N_14771,N_15939);
nand U16867 (N_16867,N_14608,N_14060);
nor U16868 (N_16868,N_15739,N_14566);
nor U16869 (N_16869,N_14536,N_14341);
or U16870 (N_16870,N_14631,N_14635);
nor U16871 (N_16871,N_15093,N_15022);
nor U16872 (N_16872,N_14968,N_14381);
or U16873 (N_16873,N_14807,N_14495);
nand U16874 (N_16874,N_14295,N_15863);
nand U16875 (N_16875,N_14636,N_15053);
nor U16876 (N_16876,N_15714,N_15094);
and U16877 (N_16877,N_15650,N_15125);
xor U16878 (N_16878,N_14732,N_14097);
and U16879 (N_16879,N_15482,N_14729);
nor U16880 (N_16880,N_14161,N_15319);
and U16881 (N_16881,N_15233,N_15029);
nor U16882 (N_16882,N_15244,N_14933);
or U16883 (N_16883,N_15515,N_15020);
nand U16884 (N_16884,N_14872,N_15139);
nand U16885 (N_16885,N_15443,N_14994);
nor U16886 (N_16886,N_14325,N_15267);
or U16887 (N_16887,N_14975,N_14177);
nand U16888 (N_16888,N_14250,N_15284);
nand U16889 (N_16889,N_14641,N_15728);
or U16890 (N_16890,N_14289,N_14573);
nor U16891 (N_16891,N_15584,N_15855);
nor U16892 (N_16892,N_14081,N_14961);
and U16893 (N_16893,N_15263,N_14230);
and U16894 (N_16894,N_15195,N_15524);
xor U16895 (N_16895,N_15507,N_14345);
xnor U16896 (N_16896,N_15095,N_15980);
nor U16897 (N_16897,N_14884,N_14243);
nand U16898 (N_16898,N_14987,N_15893);
or U16899 (N_16899,N_15047,N_15494);
nor U16900 (N_16900,N_14472,N_14813);
nor U16901 (N_16901,N_14730,N_14517);
nor U16902 (N_16902,N_15197,N_14927);
or U16903 (N_16903,N_14724,N_15037);
or U16904 (N_16904,N_14234,N_14421);
nand U16905 (N_16905,N_15876,N_14753);
or U16906 (N_16906,N_14327,N_15225);
nor U16907 (N_16907,N_15264,N_15314);
xor U16908 (N_16908,N_14726,N_15803);
or U16909 (N_16909,N_14745,N_14130);
nor U16910 (N_16910,N_14496,N_15408);
nand U16911 (N_16911,N_15133,N_14950);
xor U16912 (N_16912,N_14300,N_15353);
nand U16913 (N_16913,N_15563,N_15905);
nor U16914 (N_16914,N_14596,N_14966);
nor U16915 (N_16915,N_14181,N_14592);
nand U16916 (N_16916,N_15712,N_15300);
nor U16917 (N_16917,N_14923,N_15784);
or U16918 (N_16918,N_14361,N_14367);
nand U16919 (N_16919,N_14385,N_15771);
xnor U16920 (N_16920,N_14774,N_14522);
and U16921 (N_16921,N_14487,N_14559);
nor U16922 (N_16922,N_14509,N_14490);
nor U16923 (N_16923,N_15669,N_14949);
nand U16924 (N_16924,N_15102,N_14119);
and U16925 (N_16925,N_14519,N_14240);
xnor U16926 (N_16926,N_14577,N_15894);
nand U16927 (N_16927,N_14614,N_15246);
xor U16928 (N_16928,N_14143,N_14690);
or U16929 (N_16929,N_14238,N_14046);
xor U16930 (N_16930,N_15317,N_15797);
and U16931 (N_16931,N_15516,N_14646);
nor U16932 (N_16932,N_14206,N_15828);
or U16933 (N_16933,N_14236,N_14211);
xnor U16934 (N_16934,N_15156,N_15616);
nor U16935 (N_16935,N_15553,N_14332);
nand U16936 (N_16936,N_14668,N_15903);
nand U16937 (N_16937,N_15379,N_14560);
nand U16938 (N_16938,N_15929,N_14404);
nand U16939 (N_16939,N_14928,N_15250);
and U16940 (N_16940,N_15726,N_14533);
and U16941 (N_16941,N_15231,N_15290);
nor U16942 (N_16942,N_14055,N_14328);
nand U16943 (N_16943,N_14880,N_15548);
and U16944 (N_16944,N_14018,N_15175);
nand U16945 (N_16945,N_14394,N_15422);
nor U16946 (N_16946,N_15998,N_15363);
nand U16947 (N_16947,N_14426,N_15748);
and U16948 (N_16948,N_15170,N_15736);
nand U16949 (N_16949,N_14926,N_15344);
nor U16950 (N_16950,N_15496,N_15253);
and U16951 (N_16951,N_14584,N_14287);
nor U16952 (N_16952,N_15914,N_14104);
or U16953 (N_16953,N_15489,N_14930);
xor U16954 (N_16954,N_14781,N_14742);
and U16955 (N_16955,N_15145,N_14912);
nand U16956 (N_16956,N_15684,N_15324);
or U16957 (N_16957,N_15335,N_15042);
nand U16958 (N_16958,N_15792,N_14214);
and U16959 (N_16959,N_15972,N_15674);
or U16960 (N_16960,N_14454,N_15450);
nor U16961 (N_16961,N_14666,N_15199);
and U16962 (N_16962,N_15068,N_15432);
nand U16963 (N_16963,N_14878,N_14765);
or U16964 (N_16964,N_14276,N_15458);
and U16965 (N_16965,N_15958,N_15459);
or U16966 (N_16966,N_14127,N_15271);
and U16967 (N_16967,N_14871,N_15438);
nand U16968 (N_16968,N_14456,N_14431);
or U16969 (N_16969,N_14916,N_14561);
and U16970 (N_16970,N_15262,N_14502);
nand U16971 (N_16971,N_14185,N_15571);
nand U16972 (N_16972,N_15848,N_15931);
xnor U16973 (N_16973,N_15640,N_14946);
nor U16974 (N_16974,N_15895,N_15965);
nand U16975 (N_16975,N_14292,N_14825);
xor U16976 (N_16976,N_14004,N_15700);
or U16977 (N_16977,N_14764,N_14500);
nor U16978 (N_16978,N_14241,N_14516);
nor U16979 (N_16979,N_15592,N_15846);
and U16980 (N_16980,N_15252,N_14572);
nor U16981 (N_16981,N_15067,N_14486);
or U16982 (N_16982,N_14176,N_15228);
xor U16983 (N_16983,N_14948,N_14334);
nand U16984 (N_16984,N_14786,N_14344);
nor U16985 (N_16985,N_14721,N_14469);
nor U16986 (N_16986,N_15932,N_14639);
and U16987 (N_16987,N_15055,N_15858);
xnor U16988 (N_16988,N_15701,N_15796);
or U16989 (N_16989,N_15948,N_15305);
xnor U16990 (N_16990,N_14457,N_15734);
nor U16991 (N_16991,N_15382,N_14530);
xor U16992 (N_16992,N_14089,N_15676);
nor U16993 (N_16993,N_15292,N_14434);
xnor U16994 (N_16994,N_15242,N_14620);
nor U16995 (N_16995,N_14357,N_14476);
xor U16996 (N_16996,N_14800,N_14613);
or U16997 (N_16997,N_14804,N_15957);
xnor U16998 (N_16998,N_15859,N_14744);
nor U16999 (N_16999,N_14867,N_15757);
nor U17000 (N_17000,N_15013,N_15457);
nor U17001 (N_17001,N_14957,N_14894);
nor U17002 (N_17002,N_14074,N_15399);
xor U17003 (N_17003,N_14881,N_14688);
or U17004 (N_17004,N_14799,N_15189);
nor U17005 (N_17005,N_14239,N_14081);
and U17006 (N_17006,N_14289,N_14137);
and U17007 (N_17007,N_15078,N_14257);
xor U17008 (N_17008,N_15932,N_14685);
and U17009 (N_17009,N_14729,N_14572);
nand U17010 (N_17010,N_15955,N_14556);
nand U17011 (N_17011,N_15170,N_15051);
nor U17012 (N_17012,N_14664,N_15163);
xnor U17013 (N_17013,N_14428,N_15027);
and U17014 (N_17014,N_15780,N_15236);
xor U17015 (N_17015,N_15644,N_15575);
nand U17016 (N_17016,N_15334,N_15366);
nand U17017 (N_17017,N_14108,N_15127);
nand U17018 (N_17018,N_14601,N_14766);
or U17019 (N_17019,N_15685,N_14711);
and U17020 (N_17020,N_15830,N_14099);
and U17021 (N_17021,N_14840,N_14175);
nand U17022 (N_17022,N_15048,N_14187);
nand U17023 (N_17023,N_14452,N_15492);
nor U17024 (N_17024,N_14370,N_15220);
xnor U17025 (N_17025,N_14211,N_15538);
xor U17026 (N_17026,N_15451,N_14381);
nor U17027 (N_17027,N_15955,N_15953);
nor U17028 (N_17028,N_14043,N_15414);
and U17029 (N_17029,N_14745,N_14186);
or U17030 (N_17030,N_14953,N_14918);
or U17031 (N_17031,N_14427,N_15598);
nand U17032 (N_17032,N_15900,N_14651);
and U17033 (N_17033,N_14018,N_15472);
and U17034 (N_17034,N_15551,N_14148);
and U17035 (N_17035,N_14354,N_14181);
xor U17036 (N_17036,N_15461,N_14638);
and U17037 (N_17037,N_14395,N_15657);
nand U17038 (N_17038,N_14996,N_15138);
or U17039 (N_17039,N_14386,N_14480);
nor U17040 (N_17040,N_15583,N_14544);
or U17041 (N_17041,N_14968,N_15506);
xor U17042 (N_17042,N_15505,N_14334);
nor U17043 (N_17043,N_14785,N_14667);
or U17044 (N_17044,N_15422,N_15963);
xnor U17045 (N_17045,N_14291,N_15061);
nor U17046 (N_17046,N_14199,N_15932);
or U17047 (N_17047,N_15657,N_14755);
or U17048 (N_17048,N_14519,N_14842);
nor U17049 (N_17049,N_15508,N_14720);
xor U17050 (N_17050,N_14952,N_15013);
nand U17051 (N_17051,N_14414,N_14599);
nand U17052 (N_17052,N_15243,N_14109);
and U17053 (N_17053,N_14081,N_15769);
xnor U17054 (N_17054,N_15664,N_15508);
or U17055 (N_17055,N_15303,N_15383);
or U17056 (N_17056,N_15221,N_15868);
xor U17057 (N_17057,N_15560,N_15096);
or U17058 (N_17058,N_15684,N_15123);
or U17059 (N_17059,N_14485,N_15656);
nor U17060 (N_17060,N_15358,N_15565);
or U17061 (N_17061,N_14034,N_14741);
nand U17062 (N_17062,N_14588,N_15145);
nand U17063 (N_17063,N_15522,N_14802);
nor U17064 (N_17064,N_14312,N_15588);
or U17065 (N_17065,N_15026,N_15038);
nand U17066 (N_17066,N_15030,N_14382);
or U17067 (N_17067,N_15683,N_14533);
and U17068 (N_17068,N_15988,N_15787);
and U17069 (N_17069,N_14246,N_14908);
or U17070 (N_17070,N_14955,N_14493);
xnor U17071 (N_17071,N_15948,N_15661);
nand U17072 (N_17072,N_14694,N_15089);
and U17073 (N_17073,N_15357,N_14757);
xor U17074 (N_17074,N_14923,N_15338);
xnor U17075 (N_17075,N_14753,N_14582);
and U17076 (N_17076,N_14083,N_15893);
xnor U17077 (N_17077,N_15535,N_14142);
nor U17078 (N_17078,N_15842,N_15569);
xor U17079 (N_17079,N_15875,N_14906);
nand U17080 (N_17080,N_15968,N_14862);
nand U17081 (N_17081,N_15504,N_14202);
nor U17082 (N_17082,N_15346,N_14588);
nor U17083 (N_17083,N_14490,N_14078);
or U17084 (N_17084,N_15409,N_14823);
or U17085 (N_17085,N_14401,N_14934);
and U17086 (N_17086,N_14868,N_14853);
xnor U17087 (N_17087,N_15448,N_14313);
nor U17088 (N_17088,N_14444,N_15466);
nand U17089 (N_17089,N_14868,N_14916);
or U17090 (N_17090,N_15555,N_14864);
and U17091 (N_17091,N_14934,N_14978);
xnor U17092 (N_17092,N_14439,N_14011);
xnor U17093 (N_17093,N_15820,N_14259);
or U17094 (N_17094,N_14607,N_15822);
or U17095 (N_17095,N_14866,N_15286);
nor U17096 (N_17096,N_14987,N_15014);
or U17097 (N_17097,N_14342,N_15860);
and U17098 (N_17098,N_15405,N_15035);
xnor U17099 (N_17099,N_14123,N_15261);
nor U17100 (N_17100,N_15908,N_15018);
nand U17101 (N_17101,N_15205,N_14907);
nor U17102 (N_17102,N_15463,N_14179);
nand U17103 (N_17103,N_15866,N_14887);
nor U17104 (N_17104,N_14239,N_15756);
nand U17105 (N_17105,N_15402,N_14089);
xnor U17106 (N_17106,N_15316,N_15764);
nor U17107 (N_17107,N_14728,N_15784);
nand U17108 (N_17108,N_15731,N_15602);
nand U17109 (N_17109,N_15838,N_14270);
nor U17110 (N_17110,N_15956,N_15994);
xnor U17111 (N_17111,N_15303,N_15654);
nand U17112 (N_17112,N_14931,N_15123);
xnor U17113 (N_17113,N_15488,N_15328);
nor U17114 (N_17114,N_15883,N_14426);
nor U17115 (N_17115,N_14807,N_14673);
nand U17116 (N_17116,N_14478,N_15191);
and U17117 (N_17117,N_14295,N_14374);
xor U17118 (N_17118,N_14609,N_15639);
and U17119 (N_17119,N_14289,N_14032);
xor U17120 (N_17120,N_15574,N_15958);
or U17121 (N_17121,N_15031,N_15941);
nor U17122 (N_17122,N_14496,N_14976);
nor U17123 (N_17123,N_15602,N_14293);
and U17124 (N_17124,N_15256,N_14367);
nand U17125 (N_17125,N_14445,N_14669);
and U17126 (N_17126,N_14059,N_14424);
or U17127 (N_17127,N_15958,N_14248);
or U17128 (N_17128,N_15166,N_15798);
nor U17129 (N_17129,N_15970,N_14025);
nor U17130 (N_17130,N_14085,N_14985);
nor U17131 (N_17131,N_15942,N_14990);
nand U17132 (N_17132,N_14829,N_15444);
nand U17133 (N_17133,N_15808,N_14120);
nand U17134 (N_17134,N_15897,N_14315);
nand U17135 (N_17135,N_14597,N_15381);
xor U17136 (N_17136,N_14315,N_14142);
and U17137 (N_17137,N_15298,N_14406);
xor U17138 (N_17138,N_15412,N_15833);
and U17139 (N_17139,N_15363,N_15214);
or U17140 (N_17140,N_14385,N_15691);
and U17141 (N_17141,N_14769,N_14422);
nand U17142 (N_17142,N_15001,N_15991);
and U17143 (N_17143,N_14424,N_15867);
nand U17144 (N_17144,N_15763,N_14514);
nand U17145 (N_17145,N_15634,N_15011);
xnor U17146 (N_17146,N_15716,N_14978);
and U17147 (N_17147,N_14617,N_14374);
nand U17148 (N_17148,N_15007,N_15629);
nor U17149 (N_17149,N_15561,N_14506);
nor U17150 (N_17150,N_14135,N_15448);
nor U17151 (N_17151,N_14602,N_15373);
or U17152 (N_17152,N_14508,N_15535);
or U17153 (N_17153,N_14321,N_14237);
nand U17154 (N_17154,N_15033,N_15079);
nand U17155 (N_17155,N_15832,N_14708);
nand U17156 (N_17156,N_15127,N_15103);
and U17157 (N_17157,N_15121,N_15623);
nand U17158 (N_17158,N_15500,N_14846);
and U17159 (N_17159,N_15694,N_15669);
xor U17160 (N_17160,N_15985,N_14027);
and U17161 (N_17161,N_14643,N_15253);
or U17162 (N_17162,N_14241,N_15780);
nor U17163 (N_17163,N_14126,N_15435);
nand U17164 (N_17164,N_15075,N_15315);
xnor U17165 (N_17165,N_14046,N_15737);
nand U17166 (N_17166,N_15819,N_14867);
nor U17167 (N_17167,N_15434,N_14023);
xnor U17168 (N_17168,N_15506,N_15789);
or U17169 (N_17169,N_14702,N_15190);
xor U17170 (N_17170,N_15625,N_14397);
nand U17171 (N_17171,N_15983,N_14355);
or U17172 (N_17172,N_15696,N_14690);
nand U17173 (N_17173,N_14748,N_15748);
nand U17174 (N_17174,N_14564,N_14920);
or U17175 (N_17175,N_15321,N_14328);
or U17176 (N_17176,N_14088,N_15388);
nand U17177 (N_17177,N_15773,N_15256);
xnor U17178 (N_17178,N_14001,N_14263);
nor U17179 (N_17179,N_15410,N_15815);
or U17180 (N_17180,N_15326,N_14110);
xnor U17181 (N_17181,N_14665,N_15249);
or U17182 (N_17182,N_14612,N_15046);
and U17183 (N_17183,N_14796,N_14000);
nand U17184 (N_17184,N_14716,N_14813);
or U17185 (N_17185,N_14972,N_14199);
or U17186 (N_17186,N_15936,N_14649);
or U17187 (N_17187,N_14255,N_15941);
nor U17188 (N_17188,N_15106,N_15367);
nand U17189 (N_17189,N_15547,N_15566);
nor U17190 (N_17190,N_14713,N_14501);
xnor U17191 (N_17191,N_14746,N_15238);
and U17192 (N_17192,N_15411,N_14805);
or U17193 (N_17193,N_15994,N_15792);
xor U17194 (N_17194,N_15924,N_14448);
nand U17195 (N_17195,N_15351,N_14934);
and U17196 (N_17196,N_14479,N_14205);
or U17197 (N_17197,N_15346,N_14765);
nand U17198 (N_17198,N_14046,N_14719);
xor U17199 (N_17199,N_14456,N_14531);
or U17200 (N_17200,N_14560,N_15838);
and U17201 (N_17201,N_14664,N_14264);
or U17202 (N_17202,N_14501,N_15929);
and U17203 (N_17203,N_15434,N_15383);
xnor U17204 (N_17204,N_15788,N_15934);
nand U17205 (N_17205,N_15082,N_14243);
nor U17206 (N_17206,N_15705,N_15453);
xor U17207 (N_17207,N_15459,N_15841);
xor U17208 (N_17208,N_15397,N_15859);
nand U17209 (N_17209,N_14798,N_14925);
nor U17210 (N_17210,N_15789,N_14824);
and U17211 (N_17211,N_15438,N_14580);
nand U17212 (N_17212,N_15408,N_15073);
nor U17213 (N_17213,N_14977,N_14402);
or U17214 (N_17214,N_15945,N_15898);
and U17215 (N_17215,N_14365,N_14005);
nor U17216 (N_17216,N_15059,N_14293);
or U17217 (N_17217,N_15547,N_14539);
nor U17218 (N_17218,N_15498,N_15452);
or U17219 (N_17219,N_14709,N_14307);
xnor U17220 (N_17220,N_15545,N_14644);
nor U17221 (N_17221,N_15868,N_14482);
or U17222 (N_17222,N_15490,N_15235);
and U17223 (N_17223,N_14636,N_15127);
or U17224 (N_17224,N_15581,N_14715);
nand U17225 (N_17225,N_15196,N_15892);
nor U17226 (N_17226,N_14926,N_15829);
or U17227 (N_17227,N_15847,N_15497);
nand U17228 (N_17228,N_14783,N_15265);
or U17229 (N_17229,N_15683,N_15088);
or U17230 (N_17230,N_14513,N_14777);
and U17231 (N_17231,N_14517,N_15040);
or U17232 (N_17232,N_14768,N_14286);
nor U17233 (N_17233,N_14399,N_14754);
nor U17234 (N_17234,N_14517,N_14361);
xor U17235 (N_17235,N_14503,N_14944);
and U17236 (N_17236,N_14672,N_15657);
and U17237 (N_17237,N_15474,N_15451);
nand U17238 (N_17238,N_14295,N_15887);
nor U17239 (N_17239,N_15422,N_14955);
xnor U17240 (N_17240,N_14208,N_14757);
or U17241 (N_17241,N_14985,N_14049);
or U17242 (N_17242,N_14263,N_15199);
xor U17243 (N_17243,N_15235,N_14391);
nand U17244 (N_17244,N_14730,N_14932);
xor U17245 (N_17245,N_14602,N_15051);
nand U17246 (N_17246,N_14242,N_15599);
xor U17247 (N_17247,N_14665,N_15814);
nand U17248 (N_17248,N_15353,N_14811);
nor U17249 (N_17249,N_15168,N_15012);
or U17250 (N_17250,N_14054,N_14798);
nand U17251 (N_17251,N_15245,N_14111);
xor U17252 (N_17252,N_14619,N_14661);
nor U17253 (N_17253,N_15037,N_15943);
nand U17254 (N_17254,N_14481,N_15849);
xor U17255 (N_17255,N_14070,N_15560);
or U17256 (N_17256,N_15602,N_15050);
nand U17257 (N_17257,N_15469,N_15169);
or U17258 (N_17258,N_14743,N_15825);
xnor U17259 (N_17259,N_14708,N_14497);
nand U17260 (N_17260,N_14317,N_15987);
nand U17261 (N_17261,N_15918,N_14530);
xnor U17262 (N_17262,N_14313,N_15989);
nor U17263 (N_17263,N_14178,N_14343);
or U17264 (N_17264,N_14935,N_15791);
and U17265 (N_17265,N_14193,N_15843);
and U17266 (N_17266,N_14346,N_15744);
nor U17267 (N_17267,N_14052,N_15717);
or U17268 (N_17268,N_15697,N_14927);
nand U17269 (N_17269,N_15119,N_15769);
xnor U17270 (N_17270,N_15616,N_14929);
nand U17271 (N_17271,N_15273,N_14164);
xor U17272 (N_17272,N_14811,N_15625);
or U17273 (N_17273,N_14302,N_14562);
xor U17274 (N_17274,N_14647,N_15722);
nor U17275 (N_17275,N_14918,N_15975);
nor U17276 (N_17276,N_14319,N_14968);
xor U17277 (N_17277,N_15355,N_15112);
nor U17278 (N_17278,N_15600,N_14645);
and U17279 (N_17279,N_14338,N_15185);
xor U17280 (N_17280,N_14676,N_15604);
nand U17281 (N_17281,N_14296,N_15883);
and U17282 (N_17282,N_14832,N_14839);
xnor U17283 (N_17283,N_14464,N_15254);
or U17284 (N_17284,N_15243,N_14863);
nor U17285 (N_17285,N_15213,N_14325);
nand U17286 (N_17286,N_15241,N_15082);
nand U17287 (N_17287,N_14779,N_15832);
nor U17288 (N_17288,N_15685,N_14750);
nor U17289 (N_17289,N_15187,N_14426);
nor U17290 (N_17290,N_14625,N_14461);
nor U17291 (N_17291,N_14110,N_15247);
xor U17292 (N_17292,N_14290,N_15535);
and U17293 (N_17293,N_14476,N_14889);
nand U17294 (N_17294,N_15822,N_15764);
xnor U17295 (N_17295,N_14133,N_14972);
or U17296 (N_17296,N_15934,N_15504);
or U17297 (N_17297,N_14350,N_15098);
xor U17298 (N_17298,N_15098,N_14315);
and U17299 (N_17299,N_14612,N_15646);
and U17300 (N_17300,N_14943,N_15625);
xnor U17301 (N_17301,N_14617,N_14414);
nand U17302 (N_17302,N_14571,N_15192);
nor U17303 (N_17303,N_14293,N_14004);
or U17304 (N_17304,N_14920,N_14200);
or U17305 (N_17305,N_15892,N_14212);
xor U17306 (N_17306,N_15844,N_14154);
nor U17307 (N_17307,N_15391,N_15594);
or U17308 (N_17308,N_14330,N_14764);
nor U17309 (N_17309,N_15262,N_15740);
or U17310 (N_17310,N_14637,N_14231);
and U17311 (N_17311,N_15322,N_15910);
and U17312 (N_17312,N_14842,N_14014);
nor U17313 (N_17313,N_14356,N_14848);
nand U17314 (N_17314,N_15886,N_14710);
and U17315 (N_17315,N_14137,N_14730);
nor U17316 (N_17316,N_15004,N_15510);
nand U17317 (N_17317,N_14949,N_14516);
nor U17318 (N_17318,N_15844,N_15388);
nand U17319 (N_17319,N_15462,N_15074);
nor U17320 (N_17320,N_15575,N_14977);
nor U17321 (N_17321,N_15199,N_14492);
xor U17322 (N_17322,N_15313,N_14156);
and U17323 (N_17323,N_14168,N_14379);
or U17324 (N_17324,N_15737,N_15443);
or U17325 (N_17325,N_14462,N_15836);
nor U17326 (N_17326,N_14227,N_15473);
nand U17327 (N_17327,N_14047,N_14891);
xor U17328 (N_17328,N_14396,N_15644);
and U17329 (N_17329,N_14474,N_15590);
nor U17330 (N_17330,N_14842,N_15999);
nor U17331 (N_17331,N_15013,N_14600);
and U17332 (N_17332,N_15650,N_14267);
or U17333 (N_17333,N_15962,N_15515);
nor U17334 (N_17334,N_14978,N_15705);
nor U17335 (N_17335,N_15386,N_15156);
nor U17336 (N_17336,N_15383,N_14748);
and U17337 (N_17337,N_14263,N_15693);
or U17338 (N_17338,N_14497,N_14323);
and U17339 (N_17339,N_15736,N_15211);
and U17340 (N_17340,N_15906,N_15055);
nor U17341 (N_17341,N_15841,N_15656);
nand U17342 (N_17342,N_15397,N_14779);
nand U17343 (N_17343,N_14788,N_14487);
nor U17344 (N_17344,N_14369,N_14763);
nand U17345 (N_17345,N_15005,N_15861);
nor U17346 (N_17346,N_15327,N_14354);
nor U17347 (N_17347,N_15784,N_15877);
or U17348 (N_17348,N_15703,N_14835);
and U17349 (N_17349,N_15238,N_15548);
nand U17350 (N_17350,N_14862,N_14044);
or U17351 (N_17351,N_15864,N_15146);
xor U17352 (N_17352,N_15689,N_15186);
or U17353 (N_17353,N_14059,N_15439);
or U17354 (N_17354,N_15283,N_15792);
nand U17355 (N_17355,N_15076,N_14172);
and U17356 (N_17356,N_14089,N_14026);
xnor U17357 (N_17357,N_14095,N_14921);
or U17358 (N_17358,N_15394,N_14900);
nor U17359 (N_17359,N_14496,N_15526);
xnor U17360 (N_17360,N_15487,N_15380);
nor U17361 (N_17361,N_15992,N_14340);
or U17362 (N_17362,N_15195,N_14433);
or U17363 (N_17363,N_15978,N_15201);
xnor U17364 (N_17364,N_15509,N_14836);
nand U17365 (N_17365,N_15347,N_14820);
nand U17366 (N_17366,N_14153,N_14312);
nor U17367 (N_17367,N_15661,N_15810);
nor U17368 (N_17368,N_14136,N_14569);
nor U17369 (N_17369,N_15587,N_14991);
xor U17370 (N_17370,N_14037,N_14734);
and U17371 (N_17371,N_15261,N_14805);
nor U17372 (N_17372,N_15854,N_14535);
xor U17373 (N_17373,N_15276,N_15753);
nand U17374 (N_17374,N_14877,N_15305);
nor U17375 (N_17375,N_15005,N_15050);
or U17376 (N_17376,N_15552,N_15079);
nand U17377 (N_17377,N_14017,N_15335);
nor U17378 (N_17378,N_15657,N_14078);
or U17379 (N_17379,N_14246,N_14296);
nand U17380 (N_17380,N_14193,N_14547);
and U17381 (N_17381,N_14772,N_14968);
xnor U17382 (N_17382,N_15472,N_15273);
nor U17383 (N_17383,N_15234,N_14447);
or U17384 (N_17384,N_15861,N_15790);
and U17385 (N_17385,N_15504,N_15766);
or U17386 (N_17386,N_14695,N_15354);
nor U17387 (N_17387,N_15173,N_15251);
xnor U17388 (N_17388,N_14381,N_15849);
nand U17389 (N_17389,N_15727,N_14279);
xnor U17390 (N_17390,N_15206,N_14257);
and U17391 (N_17391,N_15301,N_14340);
or U17392 (N_17392,N_15999,N_15204);
nand U17393 (N_17393,N_14967,N_14173);
nor U17394 (N_17394,N_14374,N_14026);
nor U17395 (N_17395,N_14610,N_15702);
nand U17396 (N_17396,N_14264,N_14353);
nor U17397 (N_17397,N_14711,N_15174);
nand U17398 (N_17398,N_14317,N_14453);
nor U17399 (N_17399,N_14334,N_14701);
and U17400 (N_17400,N_15011,N_15304);
nand U17401 (N_17401,N_15823,N_15785);
nand U17402 (N_17402,N_14430,N_14093);
xor U17403 (N_17403,N_15576,N_14955);
xor U17404 (N_17404,N_15702,N_15438);
nor U17405 (N_17405,N_15522,N_14537);
xor U17406 (N_17406,N_14363,N_14127);
and U17407 (N_17407,N_15974,N_15384);
and U17408 (N_17408,N_14552,N_15870);
or U17409 (N_17409,N_14163,N_15546);
nand U17410 (N_17410,N_14115,N_14117);
or U17411 (N_17411,N_14641,N_15751);
or U17412 (N_17412,N_15850,N_14803);
and U17413 (N_17413,N_15473,N_15749);
and U17414 (N_17414,N_15510,N_14162);
nor U17415 (N_17415,N_14163,N_15035);
nand U17416 (N_17416,N_14543,N_15072);
nor U17417 (N_17417,N_14542,N_15959);
or U17418 (N_17418,N_14852,N_14091);
or U17419 (N_17419,N_14798,N_15859);
nand U17420 (N_17420,N_14245,N_14349);
or U17421 (N_17421,N_15017,N_15238);
or U17422 (N_17422,N_15202,N_14505);
or U17423 (N_17423,N_15881,N_14560);
nor U17424 (N_17424,N_14666,N_15614);
nor U17425 (N_17425,N_15319,N_15194);
nand U17426 (N_17426,N_14054,N_14805);
and U17427 (N_17427,N_15463,N_14514);
nor U17428 (N_17428,N_14015,N_15432);
nor U17429 (N_17429,N_14217,N_14286);
nor U17430 (N_17430,N_15146,N_14923);
nor U17431 (N_17431,N_15309,N_14096);
or U17432 (N_17432,N_15077,N_14999);
nand U17433 (N_17433,N_15047,N_15810);
nand U17434 (N_17434,N_15787,N_15004);
nor U17435 (N_17435,N_15234,N_15744);
nand U17436 (N_17436,N_14304,N_15193);
nand U17437 (N_17437,N_14426,N_14090);
or U17438 (N_17438,N_15678,N_14080);
nor U17439 (N_17439,N_15611,N_14512);
or U17440 (N_17440,N_15804,N_15397);
or U17441 (N_17441,N_14155,N_15460);
and U17442 (N_17442,N_15462,N_14857);
xor U17443 (N_17443,N_14550,N_15469);
and U17444 (N_17444,N_14896,N_15741);
and U17445 (N_17445,N_14927,N_14168);
xor U17446 (N_17446,N_15529,N_14465);
nor U17447 (N_17447,N_15663,N_15024);
or U17448 (N_17448,N_15948,N_14814);
nor U17449 (N_17449,N_15549,N_15115);
nor U17450 (N_17450,N_14187,N_14595);
nand U17451 (N_17451,N_14441,N_15822);
xnor U17452 (N_17452,N_15677,N_15744);
nand U17453 (N_17453,N_14440,N_15124);
and U17454 (N_17454,N_15191,N_15344);
xnor U17455 (N_17455,N_15966,N_14963);
nor U17456 (N_17456,N_14101,N_15209);
nor U17457 (N_17457,N_14583,N_15317);
nor U17458 (N_17458,N_15370,N_15035);
xnor U17459 (N_17459,N_14393,N_14389);
nand U17460 (N_17460,N_15069,N_14231);
xnor U17461 (N_17461,N_14927,N_14375);
nand U17462 (N_17462,N_15669,N_15109);
nand U17463 (N_17463,N_15285,N_14211);
nor U17464 (N_17464,N_14901,N_15746);
and U17465 (N_17465,N_14423,N_14932);
and U17466 (N_17466,N_15988,N_15438);
nor U17467 (N_17467,N_15915,N_15072);
nor U17468 (N_17468,N_15733,N_14705);
nor U17469 (N_17469,N_14716,N_15336);
or U17470 (N_17470,N_14592,N_15155);
nor U17471 (N_17471,N_15692,N_15505);
nand U17472 (N_17472,N_15171,N_14506);
xor U17473 (N_17473,N_15107,N_15731);
and U17474 (N_17474,N_14692,N_14507);
xor U17475 (N_17475,N_14709,N_15342);
and U17476 (N_17476,N_15911,N_15692);
nor U17477 (N_17477,N_15572,N_14723);
or U17478 (N_17478,N_14499,N_15474);
and U17479 (N_17479,N_14133,N_15015);
nand U17480 (N_17480,N_14784,N_15131);
and U17481 (N_17481,N_15614,N_14299);
or U17482 (N_17482,N_15129,N_14292);
or U17483 (N_17483,N_15366,N_15970);
nand U17484 (N_17484,N_15233,N_15875);
nor U17485 (N_17485,N_14759,N_14999);
xor U17486 (N_17486,N_14072,N_15264);
nand U17487 (N_17487,N_14750,N_15373);
nor U17488 (N_17488,N_14253,N_14113);
nor U17489 (N_17489,N_15637,N_15473);
nand U17490 (N_17490,N_15009,N_14645);
nand U17491 (N_17491,N_15443,N_14194);
xor U17492 (N_17492,N_15027,N_15019);
and U17493 (N_17493,N_14222,N_15701);
nand U17494 (N_17494,N_15647,N_15771);
nor U17495 (N_17495,N_14400,N_15310);
nand U17496 (N_17496,N_15819,N_15272);
nand U17497 (N_17497,N_15733,N_14020);
or U17498 (N_17498,N_14423,N_14822);
xnor U17499 (N_17499,N_15692,N_14221);
nor U17500 (N_17500,N_15619,N_14285);
or U17501 (N_17501,N_14167,N_15855);
nor U17502 (N_17502,N_15444,N_15686);
or U17503 (N_17503,N_15352,N_15961);
xnor U17504 (N_17504,N_15174,N_14458);
or U17505 (N_17505,N_14899,N_14689);
xnor U17506 (N_17506,N_15270,N_14078);
nand U17507 (N_17507,N_15275,N_15646);
nand U17508 (N_17508,N_14102,N_15202);
and U17509 (N_17509,N_14725,N_14101);
and U17510 (N_17510,N_15812,N_15869);
xnor U17511 (N_17511,N_15618,N_14973);
or U17512 (N_17512,N_15183,N_15816);
nand U17513 (N_17513,N_14639,N_15464);
nor U17514 (N_17514,N_14293,N_15038);
nand U17515 (N_17515,N_14849,N_14059);
xor U17516 (N_17516,N_14691,N_15375);
xnor U17517 (N_17517,N_15486,N_15865);
and U17518 (N_17518,N_15693,N_15510);
or U17519 (N_17519,N_15975,N_15715);
and U17520 (N_17520,N_15834,N_15223);
and U17521 (N_17521,N_15499,N_14422);
xnor U17522 (N_17522,N_14254,N_15156);
xnor U17523 (N_17523,N_14759,N_15104);
nor U17524 (N_17524,N_14744,N_15596);
xor U17525 (N_17525,N_14988,N_14522);
nand U17526 (N_17526,N_14140,N_15854);
xnor U17527 (N_17527,N_14744,N_15487);
nand U17528 (N_17528,N_15025,N_15899);
or U17529 (N_17529,N_14170,N_15654);
nor U17530 (N_17530,N_15505,N_15914);
and U17531 (N_17531,N_14472,N_15850);
and U17532 (N_17532,N_14170,N_14007);
nor U17533 (N_17533,N_15526,N_15188);
nand U17534 (N_17534,N_15772,N_15146);
or U17535 (N_17535,N_14092,N_15136);
nand U17536 (N_17536,N_15373,N_14550);
nor U17537 (N_17537,N_15805,N_15445);
nor U17538 (N_17538,N_15775,N_14981);
xnor U17539 (N_17539,N_15529,N_14080);
and U17540 (N_17540,N_14222,N_14989);
nor U17541 (N_17541,N_15774,N_15509);
nand U17542 (N_17542,N_14322,N_14309);
or U17543 (N_17543,N_14442,N_15972);
nor U17544 (N_17544,N_15432,N_14204);
nand U17545 (N_17545,N_14909,N_15922);
nor U17546 (N_17546,N_14642,N_15708);
and U17547 (N_17547,N_14944,N_15485);
or U17548 (N_17548,N_15454,N_14934);
or U17549 (N_17549,N_14297,N_15270);
nand U17550 (N_17550,N_15970,N_14112);
and U17551 (N_17551,N_15809,N_15185);
nor U17552 (N_17552,N_14965,N_14219);
or U17553 (N_17553,N_14191,N_15116);
nand U17554 (N_17554,N_14737,N_14703);
nor U17555 (N_17555,N_15405,N_15918);
or U17556 (N_17556,N_14083,N_14254);
nor U17557 (N_17557,N_14306,N_15685);
xnor U17558 (N_17558,N_15852,N_14993);
nor U17559 (N_17559,N_14808,N_15969);
nor U17560 (N_17560,N_15377,N_15097);
xnor U17561 (N_17561,N_15283,N_15471);
xnor U17562 (N_17562,N_14997,N_15417);
nor U17563 (N_17563,N_15193,N_14072);
and U17564 (N_17564,N_15337,N_15616);
or U17565 (N_17565,N_14419,N_15545);
xor U17566 (N_17566,N_14504,N_15153);
or U17567 (N_17567,N_14692,N_14364);
xor U17568 (N_17568,N_15077,N_14045);
xor U17569 (N_17569,N_15277,N_15316);
nor U17570 (N_17570,N_15585,N_14346);
or U17571 (N_17571,N_15661,N_14037);
xnor U17572 (N_17572,N_15429,N_15918);
and U17573 (N_17573,N_14289,N_14975);
and U17574 (N_17574,N_15974,N_15478);
or U17575 (N_17575,N_14487,N_14979);
nand U17576 (N_17576,N_15533,N_15763);
nor U17577 (N_17577,N_15762,N_14542);
xnor U17578 (N_17578,N_14259,N_14611);
nand U17579 (N_17579,N_14322,N_15611);
and U17580 (N_17580,N_15760,N_14660);
or U17581 (N_17581,N_14512,N_15158);
nor U17582 (N_17582,N_14701,N_14478);
xor U17583 (N_17583,N_14666,N_15730);
xor U17584 (N_17584,N_14738,N_15594);
xor U17585 (N_17585,N_15256,N_14278);
and U17586 (N_17586,N_15940,N_14037);
xor U17587 (N_17587,N_15510,N_14322);
or U17588 (N_17588,N_14683,N_15555);
or U17589 (N_17589,N_15095,N_15199);
xor U17590 (N_17590,N_14876,N_15166);
xnor U17591 (N_17591,N_15887,N_14958);
nor U17592 (N_17592,N_15633,N_14900);
and U17593 (N_17593,N_14834,N_14728);
and U17594 (N_17594,N_14868,N_14624);
nor U17595 (N_17595,N_14894,N_15264);
xnor U17596 (N_17596,N_14353,N_15609);
or U17597 (N_17597,N_15119,N_14436);
nor U17598 (N_17598,N_14666,N_14752);
or U17599 (N_17599,N_14479,N_14233);
nand U17600 (N_17600,N_14500,N_14740);
nor U17601 (N_17601,N_14775,N_14685);
nor U17602 (N_17602,N_15543,N_14667);
xnor U17603 (N_17603,N_15419,N_15956);
xor U17604 (N_17604,N_14984,N_14605);
or U17605 (N_17605,N_15911,N_14057);
or U17606 (N_17606,N_15809,N_14806);
nand U17607 (N_17607,N_14188,N_14342);
and U17608 (N_17608,N_14030,N_14808);
or U17609 (N_17609,N_14700,N_14876);
nand U17610 (N_17610,N_14818,N_14156);
nand U17611 (N_17611,N_15758,N_15108);
nand U17612 (N_17612,N_14527,N_14883);
xor U17613 (N_17613,N_15673,N_14279);
and U17614 (N_17614,N_15905,N_14577);
xor U17615 (N_17615,N_14214,N_14801);
or U17616 (N_17616,N_14975,N_14502);
xnor U17617 (N_17617,N_14420,N_15479);
and U17618 (N_17618,N_15711,N_14369);
nand U17619 (N_17619,N_15139,N_15907);
nand U17620 (N_17620,N_15594,N_14246);
or U17621 (N_17621,N_15664,N_14204);
or U17622 (N_17622,N_14079,N_14479);
or U17623 (N_17623,N_14085,N_14244);
xnor U17624 (N_17624,N_14683,N_15146);
nand U17625 (N_17625,N_14498,N_15545);
xor U17626 (N_17626,N_14711,N_15152);
xor U17627 (N_17627,N_15576,N_15487);
and U17628 (N_17628,N_14532,N_15684);
nor U17629 (N_17629,N_14220,N_15948);
nand U17630 (N_17630,N_14769,N_14894);
or U17631 (N_17631,N_15308,N_14634);
nand U17632 (N_17632,N_15154,N_14740);
or U17633 (N_17633,N_14032,N_15317);
or U17634 (N_17634,N_15725,N_15271);
xnor U17635 (N_17635,N_14277,N_15214);
or U17636 (N_17636,N_14869,N_15922);
nand U17637 (N_17637,N_14798,N_15470);
and U17638 (N_17638,N_15799,N_15308);
xnor U17639 (N_17639,N_15682,N_14807);
xor U17640 (N_17640,N_14492,N_15929);
or U17641 (N_17641,N_14813,N_14393);
or U17642 (N_17642,N_15115,N_14440);
and U17643 (N_17643,N_14726,N_14804);
nor U17644 (N_17644,N_14313,N_15680);
or U17645 (N_17645,N_15564,N_15123);
nor U17646 (N_17646,N_15876,N_15417);
xnor U17647 (N_17647,N_15015,N_14280);
nor U17648 (N_17648,N_15213,N_15347);
nor U17649 (N_17649,N_14843,N_14634);
nand U17650 (N_17650,N_15101,N_14714);
nand U17651 (N_17651,N_14742,N_14916);
xor U17652 (N_17652,N_15447,N_14725);
nand U17653 (N_17653,N_15438,N_14560);
nand U17654 (N_17654,N_15738,N_15114);
nor U17655 (N_17655,N_14446,N_14068);
nand U17656 (N_17656,N_15459,N_14740);
nor U17657 (N_17657,N_14840,N_14839);
xor U17658 (N_17658,N_14353,N_15876);
nor U17659 (N_17659,N_15117,N_15672);
xnor U17660 (N_17660,N_15941,N_14112);
nand U17661 (N_17661,N_14710,N_15709);
or U17662 (N_17662,N_14804,N_14926);
xor U17663 (N_17663,N_14642,N_14170);
and U17664 (N_17664,N_14990,N_14008);
nor U17665 (N_17665,N_15555,N_15787);
nand U17666 (N_17666,N_14941,N_14853);
nor U17667 (N_17667,N_14381,N_15879);
and U17668 (N_17668,N_14595,N_15731);
nand U17669 (N_17669,N_15978,N_14844);
or U17670 (N_17670,N_15897,N_15581);
nand U17671 (N_17671,N_14326,N_14714);
or U17672 (N_17672,N_14528,N_15678);
or U17673 (N_17673,N_15025,N_14492);
nand U17674 (N_17674,N_15212,N_14019);
or U17675 (N_17675,N_15352,N_15541);
and U17676 (N_17676,N_14920,N_15551);
xor U17677 (N_17677,N_15694,N_14949);
or U17678 (N_17678,N_14197,N_14469);
and U17679 (N_17679,N_14820,N_14168);
nand U17680 (N_17680,N_15634,N_14684);
nand U17681 (N_17681,N_15223,N_14282);
nor U17682 (N_17682,N_14544,N_14489);
nor U17683 (N_17683,N_15752,N_14259);
xnor U17684 (N_17684,N_14786,N_15928);
nand U17685 (N_17685,N_14912,N_14958);
and U17686 (N_17686,N_15204,N_15470);
or U17687 (N_17687,N_15237,N_15009);
nand U17688 (N_17688,N_14105,N_15724);
nor U17689 (N_17689,N_14074,N_14609);
xor U17690 (N_17690,N_15574,N_14993);
or U17691 (N_17691,N_14145,N_15458);
and U17692 (N_17692,N_15669,N_15329);
nor U17693 (N_17693,N_15398,N_14931);
and U17694 (N_17694,N_15631,N_15951);
nor U17695 (N_17695,N_14836,N_14454);
nor U17696 (N_17696,N_15613,N_14955);
or U17697 (N_17697,N_14220,N_15582);
or U17698 (N_17698,N_15949,N_14796);
nand U17699 (N_17699,N_15941,N_14552);
xor U17700 (N_17700,N_14207,N_14308);
xor U17701 (N_17701,N_15095,N_14414);
nor U17702 (N_17702,N_15224,N_14258);
xnor U17703 (N_17703,N_15982,N_14257);
and U17704 (N_17704,N_14676,N_14045);
or U17705 (N_17705,N_15324,N_15406);
xnor U17706 (N_17706,N_14375,N_14112);
xor U17707 (N_17707,N_15974,N_14113);
xnor U17708 (N_17708,N_14437,N_14542);
and U17709 (N_17709,N_14649,N_14323);
or U17710 (N_17710,N_14580,N_14540);
and U17711 (N_17711,N_15432,N_15591);
nor U17712 (N_17712,N_15438,N_14506);
nor U17713 (N_17713,N_15111,N_15505);
nand U17714 (N_17714,N_15979,N_15130);
xnor U17715 (N_17715,N_14750,N_14564);
xor U17716 (N_17716,N_15340,N_14499);
or U17717 (N_17717,N_14849,N_14824);
nand U17718 (N_17718,N_14947,N_15379);
xnor U17719 (N_17719,N_15685,N_14085);
xnor U17720 (N_17720,N_15047,N_15860);
nand U17721 (N_17721,N_14696,N_15094);
xnor U17722 (N_17722,N_15662,N_14183);
nor U17723 (N_17723,N_14173,N_15683);
nand U17724 (N_17724,N_15843,N_15091);
and U17725 (N_17725,N_15382,N_15594);
and U17726 (N_17726,N_15449,N_15558);
nor U17727 (N_17727,N_14600,N_15947);
nor U17728 (N_17728,N_15990,N_14092);
or U17729 (N_17729,N_14704,N_14686);
nor U17730 (N_17730,N_14042,N_15468);
or U17731 (N_17731,N_15549,N_15306);
nor U17732 (N_17732,N_15138,N_14892);
nand U17733 (N_17733,N_15768,N_14267);
nand U17734 (N_17734,N_15322,N_15211);
and U17735 (N_17735,N_14059,N_15873);
xnor U17736 (N_17736,N_14874,N_14300);
and U17737 (N_17737,N_15925,N_15308);
or U17738 (N_17738,N_15396,N_15506);
or U17739 (N_17739,N_15794,N_14310);
xor U17740 (N_17740,N_14312,N_14039);
nand U17741 (N_17741,N_14984,N_15479);
nand U17742 (N_17742,N_14100,N_14794);
nor U17743 (N_17743,N_15102,N_14317);
and U17744 (N_17744,N_14731,N_14181);
or U17745 (N_17745,N_14541,N_15650);
or U17746 (N_17746,N_14938,N_14859);
nor U17747 (N_17747,N_15671,N_14292);
nand U17748 (N_17748,N_14374,N_15869);
nand U17749 (N_17749,N_15782,N_14386);
nor U17750 (N_17750,N_14283,N_14541);
and U17751 (N_17751,N_14392,N_15437);
nor U17752 (N_17752,N_14855,N_15139);
and U17753 (N_17753,N_15679,N_15312);
nor U17754 (N_17754,N_15880,N_15971);
xnor U17755 (N_17755,N_15641,N_14894);
xor U17756 (N_17756,N_15703,N_15485);
or U17757 (N_17757,N_14833,N_14910);
nand U17758 (N_17758,N_14083,N_15175);
xor U17759 (N_17759,N_15882,N_15828);
xnor U17760 (N_17760,N_15491,N_15420);
nor U17761 (N_17761,N_14582,N_14214);
nor U17762 (N_17762,N_15155,N_15039);
and U17763 (N_17763,N_15961,N_15802);
or U17764 (N_17764,N_14569,N_14211);
nor U17765 (N_17765,N_15018,N_14274);
nand U17766 (N_17766,N_15412,N_15873);
or U17767 (N_17767,N_14866,N_15774);
or U17768 (N_17768,N_14015,N_14747);
xor U17769 (N_17769,N_15416,N_15610);
or U17770 (N_17770,N_15762,N_14935);
xor U17771 (N_17771,N_14053,N_14441);
xnor U17772 (N_17772,N_14721,N_14221);
nand U17773 (N_17773,N_14646,N_15141);
nor U17774 (N_17774,N_15538,N_15664);
and U17775 (N_17775,N_15173,N_15346);
xnor U17776 (N_17776,N_14860,N_15099);
xnor U17777 (N_17777,N_15490,N_15599);
nor U17778 (N_17778,N_14210,N_14542);
nand U17779 (N_17779,N_14602,N_14732);
nand U17780 (N_17780,N_14757,N_15181);
and U17781 (N_17781,N_14231,N_15787);
or U17782 (N_17782,N_15002,N_14513);
nor U17783 (N_17783,N_15949,N_15003);
nand U17784 (N_17784,N_14484,N_15868);
nand U17785 (N_17785,N_15866,N_15712);
or U17786 (N_17786,N_15521,N_14366);
nand U17787 (N_17787,N_14669,N_15456);
and U17788 (N_17788,N_14023,N_15220);
xnor U17789 (N_17789,N_15874,N_14623);
nand U17790 (N_17790,N_15102,N_15026);
nor U17791 (N_17791,N_15064,N_15062);
xor U17792 (N_17792,N_15077,N_15004);
xor U17793 (N_17793,N_14634,N_15448);
nor U17794 (N_17794,N_14498,N_15451);
and U17795 (N_17795,N_14264,N_15383);
and U17796 (N_17796,N_14030,N_14675);
nor U17797 (N_17797,N_14930,N_15449);
or U17798 (N_17798,N_15722,N_14526);
nand U17799 (N_17799,N_14501,N_14561);
or U17800 (N_17800,N_14614,N_14466);
nand U17801 (N_17801,N_14262,N_14539);
and U17802 (N_17802,N_15150,N_14395);
nand U17803 (N_17803,N_15389,N_14532);
xor U17804 (N_17804,N_14599,N_15710);
nor U17805 (N_17805,N_14535,N_15956);
and U17806 (N_17806,N_14644,N_15397);
nor U17807 (N_17807,N_15916,N_15567);
nor U17808 (N_17808,N_14847,N_15984);
or U17809 (N_17809,N_15227,N_15742);
xnor U17810 (N_17810,N_15559,N_15552);
nand U17811 (N_17811,N_15347,N_14693);
xnor U17812 (N_17812,N_15713,N_14530);
or U17813 (N_17813,N_14439,N_15295);
or U17814 (N_17814,N_15586,N_14850);
nand U17815 (N_17815,N_14244,N_14144);
nor U17816 (N_17816,N_15733,N_15690);
and U17817 (N_17817,N_15776,N_14747);
or U17818 (N_17818,N_15199,N_14385);
or U17819 (N_17819,N_15920,N_14656);
nor U17820 (N_17820,N_14685,N_15405);
nand U17821 (N_17821,N_14927,N_14294);
xor U17822 (N_17822,N_15513,N_15099);
nor U17823 (N_17823,N_14294,N_14020);
and U17824 (N_17824,N_15815,N_15364);
xor U17825 (N_17825,N_14736,N_15250);
and U17826 (N_17826,N_15254,N_15372);
and U17827 (N_17827,N_14408,N_15259);
xor U17828 (N_17828,N_15792,N_15237);
or U17829 (N_17829,N_14663,N_14519);
nand U17830 (N_17830,N_15382,N_14063);
xor U17831 (N_17831,N_14586,N_15927);
nand U17832 (N_17832,N_15963,N_14468);
or U17833 (N_17833,N_14768,N_14504);
xnor U17834 (N_17834,N_15815,N_14491);
nand U17835 (N_17835,N_15101,N_15556);
or U17836 (N_17836,N_14811,N_15990);
nor U17837 (N_17837,N_15735,N_14731);
nand U17838 (N_17838,N_15058,N_15124);
and U17839 (N_17839,N_15043,N_15975);
or U17840 (N_17840,N_14460,N_14226);
and U17841 (N_17841,N_14503,N_14290);
xnor U17842 (N_17842,N_15421,N_14479);
nand U17843 (N_17843,N_15502,N_14091);
xor U17844 (N_17844,N_14931,N_15606);
nor U17845 (N_17845,N_15377,N_14046);
nand U17846 (N_17846,N_15783,N_14737);
nor U17847 (N_17847,N_15785,N_14323);
and U17848 (N_17848,N_14541,N_14657);
nor U17849 (N_17849,N_15864,N_15483);
xnor U17850 (N_17850,N_15326,N_15991);
xor U17851 (N_17851,N_15688,N_14925);
nor U17852 (N_17852,N_14638,N_15825);
nor U17853 (N_17853,N_15780,N_15667);
or U17854 (N_17854,N_14851,N_14642);
and U17855 (N_17855,N_15891,N_14757);
nand U17856 (N_17856,N_15874,N_14362);
nand U17857 (N_17857,N_14833,N_15950);
nand U17858 (N_17858,N_15896,N_15511);
nor U17859 (N_17859,N_14152,N_15782);
nand U17860 (N_17860,N_15347,N_14868);
or U17861 (N_17861,N_15427,N_14165);
and U17862 (N_17862,N_15079,N_15826);
nor U17863 (N_17863,N_14370,N_15525);
xor U17864 (N_17864,N_15790,N_15142);
xnor U17865 (N_17865,N_15417,N_15564);
xor U17866 (N_17866,N_15436,N_14689);
or U17867 (N_17867,N_14027,N_15374);
xnor U17868 (N_17868,N_15300,N_15808);
and U17869 (N_17869,N_15355,N_14352);
nor U17870 (N_17870,N_14086,N_15394);
nor U17871 (N_17871,N_14963,N_14862);
xnor U17872 (N_17872,N_14178,N_14433);
xor U17873 (N_17873,N_15620,N_14807);
xnor U17874 (N_17874,N_14395,N_15645);
xnor U17875 (N_17875,N_14813,N_14466);
or U17876 (N_17876,N_15287,N_15282);
nand U17877 (N_17877,N_14059,N_15049);
or U17878 (N_17878,N_14193,N_14984);
nand U17879 (N_17879,N_15026,N_15570);
nor U17880 (N_17880,N_14821,N_15367);
xor U17881 (N_17881,N_14329,N_15421);
nand U17882 (N_17882,N_15149,N_15537);
and U17883 (N_17883,N_14693,N_15419);
nor U17884 (N_17884,N_14756,N_14937);
nor U17885 (N_17885,N_15180,N_14628);
xor U17886 (N_17886,N_15103,N_14756);
xor U17887 (N_17887,N_15906,N_14739);
or U17888 (N_17888,N_15093,N_15826);
or U17889 (N_17889,N_15187,N_15085);
or U17890 (N_17890,N_15141,N_14478);
nand U17891 (N_17891,N_15595,N_15354);
nor U17892 (N_17892,N_14935,N_15820);
nor U17893 (N_17893,N_15948,N_14904);
xnor U17894 (N_17894,N_14271,N_15989);
xor U17895 (N_17895,N_14582,N_15814);
xnor U17896 (N_17896,N_15189,N_14955);
or U17897 (N_17897,N_15358,N_15329);
nand U17898 (N_17898,N_15452,N_14158);
xnor U17899 (N_17899,N_15003,N_15392);
nand U17900 (N_17900,N_15029,N_14401);
xnor U17901 (N_17901,N_14700,N_14087);
nor U17902 (N_17902,N_14656,N_15967);
nand U17903 (N_17903,N_14544,N_14620);
nand U17904 (N_17904,N_14902,N_14476);
and U17905 (N_17905,N_15028,N_14483);
or U17906 (N_17906,N_15614,N_15373);
xor U17907 (N_17907,N_14323,N_15615);
nand U17908 (N_17908,N_15971,N_15051);
and U17909 (N_17909,N_15125,N_15709);
nor U17910 (N_17910,N_15661,N_14669);
nor U17911 (N_17911,N_15233,N_14941);
and U17912 (N_17912,N_15047,N_14289);
and U17913 (N_17913,N_14608,N_14834);
nand U17914 (N_17914,N_15245,N_15890);
nor U17915 (N_17915,N_14865,N_15939);
or U17916 (N_17916,N_15138,N_14982);
and U17917 (N_17917,N_14992,N_15256);
nand U17918 (N_17918,N_14631,N_14577);
xor U17919 (N_17919,N_14959,N_15067);
and U17920 (N_17920,N_15795,N_14354);
and U17921 (N_17921,N_14209,N_15266);
nand U17922 (N_17922,N_14824,N_14948);
nor U17923 (N_17923,N_14209,N_14859);
and U17924 (N_17924,N_15651,N_15876);
and U17925 (N_17925,N_15836,N_14598);
xnor U17926 (N_17926,N_15167,N_14978);
nand U17927 (N_17927,N_14620,N_14766);
and U17928 (N_17928,N_14619,N_15995);
nor U17929 (N_17929,N_14583,N_15662);
nor U17930 (N_17930,N_15743,N_15938);
xnor U17931 (N_17931,N_15959,N_15496);
nand U17932 (N_17932,N_15925,N_14439);
nand U17933 (N_17933,N_14300,N_15349);
nor U17934 (N_17934,N_15379,N_15359);
nand U17935 (N_17935,N_15212,N_15019);
or U17936 (N_17936,N_15005,N_14546);
nor U17937 (N_17937,N_14969,N_15972);
and U17938 (N_17938,N_14705,N_14424);
or U17939 (N_17939,N_15130,N_15452);
and U17940 (N_17940,N_15833,N_15028);
nand U17941 (N_17941,N_15684,N_14436);
nor U17942 (N_17942,N_14795,N_15844);
nand U17943 (N_17943,N_15498,N_14607);
nand U17944 (N_17944,N_15102,N_15439);
or U17945 (N_17945,N_14136,N_15323);
or U17946 (N_17946,N_15353,N_14100);
nor U17947 (N_17947,N_15012,N_15322);
nand U17948 (N_17948,N_15345,N_15152);
and U17949 (N_17949,N_14618,N_15583);
and U17950 (N_17950,N_14764,N_15949);
nand U17951 (N_17951,N_15901,N_14927);
and U17952 (N_17952,N_14826,N_14673);
nand U17953 (N_17953,N_15164,N_15682);
nor U17954 (N_17954,N_14025,N_14124);
nand U17955 (N_17955,N_14431,N_15082);
and U17956 (N_17956,N_14451,N_15151);
xor U17957 (N_17957,N_15122,N_15940);
or U17958 (N_17958,N_14487,N_14785);
and U17959 (N_17959,N_15079,N_15540);
nor U17960 (N_17960,N_14701,N_15624);
xnor U17961 (N_17961,N_15153,N_15440);
xnor U17962 (N_17962,N_14006,N_15690);
or U17963 (N_17963,N_14075,N_15642);
and U17964 (N_17964,N_15009,N_14995);
nor U17965 (N_17965,N_14553,N_14894);
or U17966 (N_17966,N_15502,N_14878);
nand U17967 (N_17967,N_14224,N_15840);
or U17968 (N_17968,N_14553,N_14875);
and U17969 (N_17969,N_15684,N_14415);
nand U17970 (N_17970,N_15435,N_15617);
nand U17971 (N_17971,N_15699,N_14282);
nand U17972 (N_17972,N_14991,N_15242);
nand U17973 (N_17973,N_15551,N_15510);
nand U17974 (N_17974,N_15656,N_15991);
and U17975 (N_17975,N_14665,N_14400);
nor U17976 (N_17976,N_15026,N_14838);
xnor U17977 (N_17977,N_15586,N_14609);
and U17978 (N_17978,N_14444,N_15680);
xor U17979 (N_17979,N_15358,N_14971);
nand U17980 (N_17980,N_14888,N_15378);
nor U17981 (N_17981,N_15394,N_15719);
and U17982 (N_17982,N_14222,N_15142);
nand U17983 (N_17983,N_14742,N_14683);
and U17984 (N_17984,N_14558,N_14786);
and U17985 (N_17985,N_15932,N_14130);
nor U17986 (N_17986,N_15101,N_15254);
and U17987 (N_17987,N_14277,N_15082);
or U17988 (N_17988,N_15547,N_15854);
nor U17989 (N_17989,N_15176,N_14997);
or U17990 (N_17990,N_15727,N_14267);
and U17991 (N_17991,N_14716,N_14392);
or U17992 (N_17992,N_14645,N_15814);
nor U17993 (N_17993,N_15079,N_15120);
and U17994 (N_17994,N_14916,N_14698);
or U17995 (N_17995,N_15647,N_15411);
and U17996 (N_17996,N_15112,N_14507);
and U17997 (N_17997,N_14025,N_15264);
and U17998 (N_17998,N_14308,N_15721);
nand U17999 (N_17999,N_14760,N_15329);
nand U18000 (N_18000,N_17663,N_16921);
nand U18001 (N_18001,N_17937,N_16621);
xnor U18002 (N_18002,N_16259,N_17322);
nor U18003 (N_18003,N_17085,N_16347);
xnor U18004 (N_18004,N_17630,N_16583);
or U18005 (N_18005,N_17581,N_17224);
nor U18006 (N_18006,N_17132,N_17619);
or U18007 (N_18007,N_17072,N_16391);
nor U18008 (N_18008,N_16443,N_16898);
or U18009 (N_18009,N_17246,N_17609);
nor U18010 (N_18010,N_17133,N_17305);
nand U18011 (N_18011,N_17873,N_16301);
nor U18012 (N_18012,N_16791,N_17101);
nor U18013 (N_18013,N_17153,N_17091);
nor U18014 (N_18014,N_17127,N_17610);
nor U18015 (N_18015,N_16258,N_16668);
xor U18016 (N_18016,N_17177,N_17466);
and U18017 (N_18017,N_17809,N_16177);
nor U18018 (N_18018,N_16433,N_17589);
nand U18019 (N_18019,N_17641,N_16656);
or U18020 (N_18020,N_17108,N_16124);
or U18021 (N_18021,N_17147,N_16874);
nand U18022 (N_18022,N_17154,N_16514);
nand U18023 (N_18023,N_17977,N_16441);
and U18024 (N_18024,N_16011,N_17036);
nand U18025 (N_18025,N_16565,N_17478);
or U18026 (N_18026,N_17171,N_16102);
nand U18027 (N_18027,N_16842,N_16864);
xor U18028 (N_18028,N_17256,N_17999);
nor U18029 (N_18029,N_17754,N_17134);
xor U18030 (N_18030,N_16855,N_17251);
and U18031 (N_18031,N_16046,N_16755);
nor U18032 (N_18032,N_17995,N_16469);
and U18033 (N_18033,N_17897,N_17720);
xor U18034 (N_18034,N_16615,N_17096);
or U18035 (N_18035,N_17751,N_17500);
and U18036 (N_18036,N_17283,N_17302);
and U18037 (N_18037,N_17567,N_17864);
and U18038 (N_18038,N_17923,N_16551);
nand U18039 (N_18039,N_17136,N_17170);
and U18040 (N_18040,N_17038,N_16942);
nor U18041 (N_18041,N_16998,N_16742);
xnor U18042 (N_18042,N_16264,N_17672);
xor U18043 (N_18043,N_16552,N_16138);
nor U18044 (N_18044,N_17932,N_16672);
nand U18045 (N_18045,N_17094,N_16987);
or U18046 (N_18046,N_16269,N_17859);
or U18047 (N_18047,N_17150,N_16032);
or U18048 (N_18048,N_17568,N_16815);
and U18049 (N_18049,N_16848,N_17056);
nand U18050 (N_18050,N_16233,N_17802);
xnor U18051 (N_18051,N_16013,N_17936);
or U18052 (N_18052,N_16705,N_16876);
nor U18053 (N_18053,N_16939,N_17253);
nand U18054 (N_18054,N_16674,N_17240);
nand U18055 (N_18055,N_16053,N_17161);
nor U18056 (N_18056,N_16213,N_17972);
nand U18057 (N_18057,N_17539,N_16206);
nor U18058 (N_18058,N_17647,N_17002);
xor U18059 (N_18059,N_17661,N_17871);
xor U18060 (N_18060,N_17238,N_17390);
xor U18061 (N_18061,N_16450,N_17462);
nor U18062 (N_18062,N_17090,N_17687);
nor U18063 (N_18063,N_16039,N_17214);
nor U18064 (N_18064,N_16048,N_17826);
or U18065 (N_18065,N_16308,N_17047);
nor U18066 (N_18066,N_16750,N_16877);
nor U18067 (N_18067,N_16290,N_16250);
nor U18068 (N_18068,N_16067,N_17503);
xnor U18069 (N_18069,N_17285,N_17039);
nand U18070 (N_18070,N_16334,N_17213);
nor U18071 (N_18071,N_16645,N_16393);
nand U18072 (N_18072,N_16662,N_16811);
and U18073 (N_18073,N_17679,N_17145);
nor U18074 (N_18074,N_17530,N_17703);
nor U18075 (N_18075,N_17388,N_17683);
xor U18076 (N_18076,N_17446,N_16113);
nand U18077 (N_18077,N_16875,N_17645);
nand U18078 (N_18078,N_16818,N_17537);
nor U18079 (N_18079,N_16604,N_16891);
and U18080 (N_18080,N_16316,N_16911);
and U18081 (N_18081,N_16091,N_17655);
xnor U18082 (N_18082,N_17633,N_16817);
and U18083 (N_18083,N_16388,N_16485);
or U18084 (N_18084,N_17823,N_16423);
nand U18085 (N_18085,N_17548,N_16816);
nand U18086 (N_18086,N_17674,N_16295);
xor U18087 (N_18087,N_17768,N_16344);
nand U18088 (N_18088,N_16792,N_16235);
or U18089 (N_18089,N_17287,N_17459);
xnor U18090 (N_18090,N_16822,N_17423);
and U18091 (N_18091,N_17763,N_16663);
nor U18092 (N_18092,N_17340,N_16171);
nand U18093 (N_18093,N_16355,N_16904);
nand U18094 (N_18094,N_17342,N_17863);
nand U18095 (N_18095,N_16991,N_17688);
xnor U18096 (N_18096,N_17190,N_17080);
or U18097 (N_18097,N_17684,N_16505);
or U18098 (N_18098,N_17579,N_16895);
and U18099 (N_18099,N_16731,N_17780);
nand U18100 (N_18100,N_17796,N_16252);
xor U18101 (N_18101,N_17129,N_16439);
or U18102 (N_18102,N_16041,N_16919);
nor U18103 (N_18103,N_16479,N_17824);
xnor U18104 (N_18104,N_17033,N_16691);
nor U18105 (N_18105,N_16140,N_17658);
and U18106 (N_18106,N_17964,N_16541);
and U18107 (N_18107,N_17962,N_16879);
xnor U18108 (N_18108,N_16370,N_16167);
or U18109 (N_18109,N_16926,N_16854);
or U18110 (N_18110,N_17447,N_16924);
nand U18111 (N_18111,N_16180,N_16482);
or U18112 (N_18112,N_16297,N_16150);
or U18113 (N_18113,N_16516,N_17973);
or U18114 (N_18114,N_16289,N_17418);
or U18115 (N_18115,N_16786,N_17901);
nor U18116 (N_18116,N_16785,N_17515);
and U18117 (N_18117,N_17990,N_17612);
nor U18118 (N_18118,N_16456,N_17392);
and U18119 (N_18119,N_16654,N_17781);
and U18120 (N_18120,N_16179,N_17531);
or U18121 (N_18121,N_17829,N_16256);
nor U18122 (N_18122,N_16409,N_16160);
or U18123 (N_18123,N_17842,N_17347);
nor U18124 (N_18124,N_17245,N_17014);
nand U18125 (N_18125,N_16499,N_17680);
xor U18126 (N_18126,N_17350,N_17187);
nand U18127 (N_18127,N_17731,N_17594);
xor U18128 (N_18128,N_17336,N_16120);
or U18129 (N_18129,N_17818,N_17030);
xnor U18130 (N_18130,N_17266,N_17389);
nand U18131 (N_18131,N_17975,N_16064);
nor U18132 (N_18132,N_16631,N_17702);
xor U18133 (N_18133,N_16777,N_16317);
or U18134 (N_18134,N_16520,N_16843);
and U18135 (N_18135,N_17562,N_16165);
xnor U18136 (N_18136,N_17868,N_16835);
or U18137 (N_18137,N_16889,N_16447);
nand U18138 (N_18138,N_16861,N_17698);
xor U18139 (N_18139,N_16502,N_16244);
nor U18140 (N_18140,N_17352,N_16986);
xor U18141 (N_18141,N_17832,N_17095);
and U18142 (N_18142,N_16951,N_17029);
xor U18143 (N_18143,N_17670,N_16519);
nor U18144 (N_18144,N_17373,N_17361);
nand U18145 (N_18145,N_16679,N_16993);
and U18146 (N_18146,N_16477,N_17066);
nand U18147 (N_18147,N_17615,N_16022);
or U18148 (N_18148,N_16737,N_16579);
nand U18149 (N_18149,N_16484,N_17173);
nor U18150 (N_18150,N_16573,N_17560);
xor U18151 (N_18151,N_17757,N_16857);
and U18152 (N_18152,N_16694,N_16943);
or U18153 (N_18153,N_16599,N_17738);
or U18154 (N_18154,N_17149,N_16979);
xor U18155 (N_18155,N_17607,N_16675);
nor U18156 (N_18156,N_16953,N_16436);
or U18157 (N_18157,N_16188,N_17506);
nor U18158 (N_18158,N_16553,N_17559);
nor U18159 (N_18159,N_16827,N_17068);
nand U18160 (N_18160,N_16262,N_16554);
xnor U18161 (N_18161,N_16389,N_16337);
xor U18162 (N_18162,N_16728,N_17800);
nor U18163 (N_18163,N_16714,N_17954);
xor U18164 (N_18164,N_17192,N_17284);
xor U18165 (N_18165,N_16260,N_17370);
and U18166 (N_18166,N_17998,N_17465);
nor U18167 (N_18167,N_17635,N_16532);
nor U18168 (N_18168,N_16030,N_17382);
xor U18169 (N_18169,N_17669,N_17265);
xor U18170 (N_18170,N_17529,N_17541);
xor U18171 (N_18171,N_16868,N_17407);
nor U18172 (N_18172,N_17598,N_16078);
or U18173 (N_18173,N_16133,N_16017);
or U18174 (N_18174,N_16920,N_16760);
xnor U18175 (N_18175,N_16561,N_17102);
and U18176 (N_18176,N_17773,N_17926);
or U18177 (N_18177,N_16493,N_16227);
nand U18178 (N_18178,N_17237,N_16076);
xor U18179 (N_18179,N_17602,N_16710);
nor U18180 (N_18180,N_17605,N_17510);
nand U18181 (N_18181,N_16985,N_16717);
nand U18182 (N_18182,N_16923,N_17303);
xnor U18183 (N_18183,N_17070,N_16384);
or U18184 (N_18184,N_16232,N_17606);
nor U18185 (N_18185,N_17031,N_17480);
or U18186 (N_18186,N_17502,N_17097);
xor U18187 (N_18187,N_16038,N_17379);
nand U18188 (N_18188,N_17421,N_16646);
nand U18189 (N_18189,N_16821,N_17413);
xor U18190 (N_18190,N_17899,N_17384);
xor U18191 (N_18191,N_17601,N_17726);
or U18192 (N_18192,N_16051,N_16435);
xor U18193 (N_18193,N_17337,N_16147);
nor U18194 (N_18194,N_17069,N_16036);
or U18195 (N_18195,N_17062,N_17967);
xor U18196 (N_18196,N_17434,N_16324);
xor U18197 (N_18197,N_17521,N_17550);
or U18198 (N_18198,N_16653,N_16291);
nand U18199 (N_18199,N_16421,N_16172);
nor U18200 (N_18200,N_16130,N_16824);
nand U18201 (N_18201,N_17742,N_16525);
nand U18202 (N_18202,N_16361,N_17053);
and U18203 (N_18203,N_17769,N_16734);
nor U18204 (N_18204,N_17263,N_16747);
nor U18205 (N_18205,N_16066,N_16884);
or U18206 (N_18206,N_16819,N_17578);
nor U18207 (N_18207,N_17712,N_17986);
and U18208 (N_18208,N_16584,N_16853);
xor U18209 (N_18209,N_17920,N_17216);
xnor U18210 (N_18210,N_17783,N_16712);
and U18211 (N_18211,N_17428,N_17089);
and U18212 (N_18212,N_17667,N_17991);
nor U18213 (N_18213,N_16097,N_17314);
nor U18214 (N_18214,N_17533,N_16352);
nand U18215 (N_18215,N_16189,N_16556);
and U18216 (N_18216,N_16144,N_16906);
nand U18217 (N_18217,N_16429,N_16970);
or U18218 (N_18218,N_16320,N_17164);
and U18219 (N_18219,N_16152,N_17599);
nand U18220 (N_18220,N_17715,N_16153);
or U18221 (N_18221,N_17297,N_17179);
or U18222 (N_18222,N_16354,N_17577);
and U18223 (N_18223,N_16859,N_17656);
nand U18224 (N_18224,N_17344,N_17205);
xnor U18225 (N_18225,N_16358,N_17250);
nand U18226 (N_18226,N_16746,N_16830);
or U18227 (N_18227,N_16305,N_16524);
and U18228 (N_18228,N_16123,N_16190);
nand U18229 (N_18229,N_17003,N_16820);
nand U18230 (N_18230,N_17513,N_17834);
or U18231 (N_18231,N_17188,N_16428);
xnor U18232 (N_18232,N_16618,N_17135);
nand U18233 (N_18233,N_16248,N_17831);
or U18234 (N_18234,N_16914,N_17725);
nor U18235 (N_18235,N_16753,N_16600);
and U18236 (N_18236,N_17528,N_17137);
or U18237 (N_18237,N_17126,N_17634);
or U18238 (N_18238,N_17078,N_16501);
xor U18239 (N_18239,N_16945,N_16601);
or U18240 (N_18240,N_17945,N_16897);
and U18241 (N_18241,N_16251,N_17000);
or U18242 (N_18242,N_16950,N_17469);
and U18243 (N_18243,N_16468,N_16964);
nor U18244 (N_18244,N_17570,N_17328);
nor U18245 (N_18245,N_17438,N_17323);
xor U18246 (N_18246,N_16218,N_17678);
nand U18247 (N_18247,N_17121,N_17196);
or U18248 (N_18248,N_17181,N_17339);
or U18249 (N_18249,N_16782,N_17890);
nor U18250 (N_18250,N_17701,N_17957);
nor U18251 (N_18251,N_16744,N_16274);
and U18252 (N_18252,N_17209,N_16548);
xor U18253 (N_18253,N_17608,N_16191);
or U18254 (N_18254,N_16803,N_17772);
xnor U18255 (N_18255,N_17282,N_17919);
nand U18256 (N_18256,N_17182,N_17782);
nand U18257 (N_18257,N_17050,N_16383);
nand U18258 (N_18258,N_17983,N_16687);
and U18259 (N_18259,N_17393,N_17639);
xnor U18260 (N_18260,N_17005,N_17944);
and U18261 (N_18261,N_17792,N_16885);
and U18262 (N_18262,N_16238,N_17113);
nand U18263 (N_18263,N_17477,N_16413);
nand U18264 (N_18264,N_17844,N_17719);
xnor U18265 (N_18265,N_16214,N_17142);
nand U18266 (N_18266,N_17636,N_17996);
or U18267 (N_18267,N_17877,N_16912);
and U18268 (N_18268,N_16764,N_16931);
or U18269 (N_18269,N_16693,N_16922);
or U18270 (N_18270,N_16963,N_16087);
xor U18271 (N_18271,N_16806,N_16692);
or U18272 (N_18272,N_16606,N_16709);
xor U18273 (N_18273,N_17222,N_17067);
nand U18274 (N_18274,N_17507,N_16761);
or U18275 (N_18275,N_17854,N_16356);
and U18276 (N_18276,N_17320,N_17059);
or U18277 (N_18277,N_17160,N_17939);
nor U18278 (N_18278,N_17816,N_17694);
or U18279 (N_18279,N_17843,N_17232);
and U18280 (N_18280,N_16567,N_17898);
xnor U18281 (N_18281,N_17290,N_17243);
xor U18282 (N_18282,N_17774,N_17026);
nor U18283 (N_18283,N_16122,N_16278);
xor U18284 (N_18284,N_16417,N_17316);
xor U18285 (N_18285,N_16340,N_16804);
and U18286 (N_18286,N_17906,N_17318);
or U18287 (N_18287,N_17564,N_17269);
xnor U18288 (N_18288,N_17759,N_16222);
nand U18289 (N_18289,N_17288,N_16425);
xnor U18290 (N_18290,N_16664,N_16476);
xor U18291 (N_18291,N_16104,N_16472);
and U18292 (N_18292,N_17495,N_16159);
xnor U18293 (N_18293,N_17911,N_16292);
xor U18294 (N_18294,N_16156,N_16220);
nand U18295 (N_18295,N_16142,N_17805);
xnor U18296 (N_18296,N_16062,N_17304);
xnor U18297 (N_18297,N_17479,N_16648);
and U18298 (N_18298,N_16330,N_16716);
nor U18299 (N_18299,N_17907,N_17046);
and U18300 (N_18300,N_17184,N_16170);
nor U18301 (N_18301,N_16367,N_16007);
nand U18302 (N_18302,N_17692,N_17985);
xnor U18303 (N_18303,N_16770,N_16281);
nor U18304 (N_18304,N_16173,N_16607);
nand U18305 (N_18305,N_16800,N_17858);
nand U18306 (N_18306,N_17662,N_17885);
nand U18307 (N_18307,N_17012,N_17793);
nor U18308 (N_18308,N_17207,N_17249);
nand U18309 (N_18309,N_16775,N_17399);
xnor U18310 (N_18310,N_16302,N_16808);
xnor U18311 (N_18311,N_17021,N_17894);
nand U18312 (N_18312,N_17387,N_16195);
nor U18313 (N_18313,N_16681,N_16397);
and U18314 (N_18314,N_16415,N_16743);
and U18315 (N_18315,N_16155,N_16504);
and U18316 (N_18316,N_16266,N_16465);
or U18317 (N_18317,N_16410,N_16670);
xor U18318 (N_18318,N_17426,N_16759);
nor U18319 (N_18319,N_17404,N_16910);
nand U18320 (N_18320,N_17042,N_16080);
and U18321 (N_18321,N_17358,N_16570);
nor U18322 (N_18322,N_17227,N_16143);
nand U18323 (N_18323,N_16339,N_16380);
nand U18324 (N_18324,N_16009,N_16946);
nor U18325 (N_18325,N_17354,N_16478);
nor U18326 (N_18326,N_17498,N_16119);
or U18327 (N_18327,N_17378,N_17511);
or U18328 (N_18328,N_17439,N_16839);
nand U18329 (N_18329,N_16589,N_17125);
or U18330 (N_18330,N_16272,N_16515);
and U18331 (N_18331,N_17377,N_16201);
and U18332 (N_18332,N_17105,N_16578);
nor U18333 (N_18333,N_17406,N_16459);
nor U18334 (N_18334,N_17553,N_17155);
nand U18335 (N_18335,N_16245,N_17431);
xnor U18336 (N_18336,N_16503,N_16639);
nor U18337 (N_18337,N_16224,N_16916);
or U18338 (N_18338,N_17355,N_17756);
or U18339 (N_18339,N_17931,N_16497);
nor U18340 (N_18340,N_17968,N_17784);
or U18341 (N_18341,N_17419,N_16765);
nor U18342 (N_18342,N_17023,N_17079);
nand U18343 (N_18343,N_16431,N_17152);
and U18344 (N_18344,N_17924,N_16669);
nor U18345 (N_18345,N_16304,N_16636);
xor U18346 (N_18346,N_17229,N_17686);
nand U18347 (N_18347,N_16902,N_16070);
nor U18348 (N_18348,N_17846,N_17371);
nor U18349 (N_18349,N_16137,N_17411);
and U18350 (N_18350,N_16597,N_17797);
xor U18351 (N_18351,N_17724,N_17312);
nand U18352 (N_18352,N_16762,N_16121);
nand U18353 (N_18353,N_16451,N_16257);
and U18354 (N_18354,N_17799,N_16186);
or U18355 (N_18355,N_16182,N_17082);
or U18356 (N_18356,N_16392,N_16253);
nand U18357 (N_18357,N_17043,N_16569);
nand U18358 (N_18358,N_16933,N_17194);
and U18359 (N_18359,N_17575,N_16293);
or U18360 (N_18360,N_16054,N_17206);
nor U18361 (N_18361,N_16660,N_17275);
nand U18362 (N_18362,N_17013,N_17010);
or U18363 (N_18363,N_16194,N_16586);
nor U18364 (N_18364,N_17252,N_17481);
nand U18365 (N_18365,N_17143,N_16215);
nor U18366 (N_18366,N_16972,N_17364);
or U18367 (N_18367,N_17211,N_17963);
xnor U18368 (N_18368,N_17886,N_17948);
nor U18369 (N_18369,N_17737,N_16061);
xnor U18370 (N_18370,N_16114,N_17953);
or U18371 (N_18371,N_17280,N_17604);
nand U18372 (N_18372,N_17436,N_16027);
or U18373 (N_18373,N_16322,N_17812);
nand U18374 (N_18374,N_16125,N_17801);
nor U18375 (N_18375,N_17261,N_17811);
or U18376 (N_18376,N_16682,N_16825);
xnor U18377 (N_18377,N_16328,N_17632);
nor U18378 (N_18378,N_17928,N_17274);
or U18379 (N_18379,N_16990,N_17435);
nor U18380 (N_18380,N_16065,N_17665);
xnor U18381 (N_18381,N_17007,N_16342);
xnor U18382 (N_18382,N_17821,N_17162);
xnor U18383 (N_18383,N_17117,N_16483);
and U18384 (N_18384,N_17174,N_16956);
or U18385 (N_18385,N_16587,N_16386);
and U18386 (N_18386,N_17074,N_17360);
and U18387 (N_18387,N_17935,N_17257);
nand U18388 (N_18388,N_17084,N_16632);
or U18389 (N_18389,N_16212,N_16852);
nor U18390 (N_18390,N_16141,N_16845);
xnor U18391 (N_18391,N_16627,N_17949);
xnor U18392 (N_18392,N_16312,N_17855);
nand U18393 (N_18393,N_17345,N_16677);
nand U18394 (N_18394,N_17167,N_16040);
nand U18395 (N_18395,N_17348,N_16591);
nand U18396 (N_18396,N_17139,N_17730);
xnor U18397 (N_18397,N_16594,N_17705);
and U18398 (N_18398,N_16457,N_16470);
xnor U18399 (N_18399,N_16458,N_17468);
or U18400 (N_18400,N_17292,N_16767);
xor U18401 (N_18401,N_17119,N_17760);
xor U18402 (N_18402,N_16079,N_17300);
nand U18403 (N_18403,N_17200,N_16338);
xnor U18404 (N_18404,N_16231,N_17707);
nor U18405 (N_18405,N_16239,N_16086);
nor U18406 (N_18406,N_17696,N_16975);
nor U18407 (N_18407,N_17087,N_17482);
or U18408 (N_18408,N_16847,N_17018);
xor U18409 (N_18409,N_16778,N_17111);
nor U18410 (N_18410,N_16241,N_17400);
nand U18411 (N_18411,N_17277,N_17808);
or U18412 (N_18412,N_16807,N_17106);
and U18413 (N_18413,N_17644,N_17158);
nor U18414 (N_18414,N_16050,N_16892);
xnor U18415 (N_18415,N_17351,N_17467);
xor U18416 (N_18416,N_17412,N_17828);
and U18417 (N_18417,N_17526,N_16193);
nor U18418 (N_18418,N_17497,N_16754);
and U18419 (N_18419,N_16265,N_17475);
xor U18420 (N_18420,N_17518,N_16109);
or U18421 (N_18421,N_17422,N_16420);
nand U18422 (N_18422,N_17856,N_16613);
nor U18423 (N_18423,N_17959,N_17603);
xor U18424 (N_18424,N_16058,N_16460);
or U18425 (N_18425,N_16192,N_17100);
xnor U18426 (N_18426,N_16813,N_17375);
or U18427 (N_18427,N_17169,N_16723);
nand U18428 (N_18428,N_17806,N_16560);
nor U18429 (N_18429,N_16683,N_16625);
or U18430 (N_18430,N_16512,N_17989);
or U18431 (N_18431,N_16900,N_16035);
nand U18432 (N_18432,N_16965,N_16696);
and U18433 (N_18433,N_17766,N_16846);
and U18434 (N_18434,N_17118,N_16135);
nor U18435 (N_18435,N_17722,N_16365);
xor U18436 (N_18436,N_16210,N_16486);
nor U18437 (N_18437,N_16836,N_17576);
nor U18438 (N_18438,N_17994,N_17586);
nor U18439 (N_18439,N_16325,N_17307);
and U18440 (N_18440,N_17675,N_17729);
and U18441 (N_18441,N_16890,N_17148);
or U18442 (N_18442,N_17613,N_16666);
and U18443 (N_18443,N_16907,N_17869);
or U18444 (N_18444,N_16204,N_16401);
nand U18445 (N_18445,N_17524,N_17410);
xor U18446 (N_18446,N_17402,N_16684);
or U18447 (N_18447,N_16455,N_17193);
xnor U18448 (N_18448,N_16219,N_16858);
or U18449 (N_18449,N_16357,N_17293);
nor U18450 (N_18450,N_17938,N_17073);
nor U18451 (N_18451,N_17903,N_17547);
xnor U18452 (N_18452,N_16546,N_16043);
nand U18453 (N_18453,N_16650,N_17294);
nand U18454 (N_18454,N_16100,N_17473);
nor U18455 (N_18455,N_17850,N_17444);
nand U18456 (N_18456,N_17460,N_16037);
nor U18457 (N_18457,N_17628,N_17837);
and U18458 (N_18458,N_17176,N_16833);
nor U18459 (N_18459,N_17254,N_17753);
or U18460 (N_18460,N_16111,N_17918);
and U18461 (N_18461,N_16616,N_16562);
xnor U18462 (N_18462,N_17489,N_16937);
xnor U18463 (N_18463,N_16359,N_16015);
nor U18464 (N_18464,N_17723,N_16279);
and U18465 (N_18465,N_17197,N_16812);
and U18466 (N_18466,N_17234,N_17368);
xor U18467 (N_18467,N_16789,N_17470);
or U18468 (N_18468,N_16918,N_17734);
and U18469 (N_18469,N_16074,N_17872);
nand U18470 (N_18470,N_17088,N_16136);
nand U18471 (N_18471,N_17519,N_16867);
nor U18472 (N_18472,N_16448,N_17363);
xnor U18473 (N_18473,N_16480,N_16756);
xor U18474 (N_18474,N_16901,N_17175);
nor U18475 (N_18475,N_17978,N_17588);
or U18476 (N_18476,N_16154,N_17311);
and U18477 (N_18477,N_17075,N_16886);
and U18478 (N_18478,N_16379,N_17278);
nor U18479 (N_18479,N_16196,N_17714);
or U18480 (N_18480,N_17758,N_16318);
or U18481 (N_18481,N_17219,N_16418);
and U18482 (N_18482,N_16905,N_17396);
nand U18483 (N_18483,N_16255,N_16609);
nor U18484 (N_18484,N_16856,N_16406);
or U18485 (N_18485,N_16234,N_17803);
nor U18486 (N_18486,N_16572,N_17353);
xor U18487 (N_18487,N_16680,N_17165);
nand U18488 (N_18488,N_16880,N_16678);
or U18489 (N_18489,N_16657,N_17540);
nor U18490 (N_18490,N_17827,N_16139);
nor U18491 (N_18491,N_17156,N_17346);
and U18492 (N_18492,N_17916,N_17386);
nor U18493 (N_18493,N_16612,N_17777);
xor U18494 (N_18494,N_16373,N_16799);
nand U18495 (N_18495,N_16055,N_17220);
nand U18496 (N_18496,N_17848,N_17425);
xnor U18497 (N_18497,N_17618,N_17092);
and U18498 (N_18498,N_17943,N_17747);
nand U18499 (N_18499,N_16473,N_17584);
xnor U18500 (N_18500,N_16823,N_17883);
nor U18501 (N_18501,N_17851,N_17004);
and U18502 (N_18502,N_17223,N_17866);
and U18503 (N_18503,N_17942,N_16603);
nand U18504 (N_18504,N_16449,N_17319);
nor U18505 (N_18505,N_16313,N_17852);
and U18506 (N_18506,N_16844,N_17921);
and U18507 (N_18507,N_17741,N_17693);
xnor U18508 (N_18508,N_16829,N_16403);
nor U18509 (N_18509,N_16385,N_17657);
or U18510 (N_18510,N_17982,N_17966);
or U18511 (N_18511,N_16108,N_16276);
nor U18512 (N_18512,N_17660,N_16909);
xor U18513 (N_18513,N_16608,N_17381);
and U18514 (N_18514,N_16101,N_16249);
and U18515 (N_18515,N_16863,N_17542);
nand U18516 (N_18516,N_16658,N_17417);
nand U18517 (N_18517,N_16426,N_17372);
nor U18518 (N_18518,N_17201,N_16563);
nand U18519 (N_18519,N_16781,N_16461);
xnor U18520 (N_18520,N_16166,N_17051);
nor U18521 (N_18521,N_17795,N_16810);
nand U18522 (N_18522,N_17454,N_16841);
xor U18523 (N_18523,N_17556,N_16995);
or U18524 (N_18524,N_17086,N_16790);
nand U18525 (N_18525,N_16971,N_17366);
nor U18526 (N_18526,N_16273,N_17081);
or U18527 (N_18527,N_16619,N_17980);
xor U18528 (N_18528,N_16862,N_16726);
nand U18529 (N_18529,N_16277,N_16134);
and U18530 (N_18530,N_16736,N_16327);
nand U18531 (N_18531,N_16713,N_16596);
nor U18532 (N_18532,N_17700,N_16063);
or U18533 (N_18533,N_17652,N_17571);
and U18534 (N_18534,N_16973,N_16208);
xor U18535 (N_18535,N_17840,N_17764);
nand U18536 (N_18536,N_16949,N_17600);
or U18537 (N_18537,N_17739,N_16298);
or U18538 (N_18538,N_16024,N_17833);
nor U18539 (N_18539,N_17514,N_17034);
nand U18540 (N_18540,N_17308,N_17879);
xor U18541 (N_18541,N_16702,N_17597);
xor U18542 (N_18542,N_16346,N_16414);
nand U18543 (N_18543,N_17496,N_17504);
and U18544 (N_18544,N_16335,N_17071);
xor U18545 (N_18545,N_16296,N_17064);
nor U18546 (N_18546,N_17971,N_17791);
nor U18547 (N_18547,N_17534,N_17241);
or U18548 (N_18548,N_17917,N_16535);
nor U18549 (N_18549,N_17189,N_16093);
xor U18550 (N_18550,N_17794,N_17555);
nor U18551 (N_18551,N_16667,N_16209);
and U18552 (N_18552,N_16598,N_17841);
and U18553 (N_18553,N_16112,N_16788);
nand U18554 (N_18554,N_16697,N_16023);
and U18555 (N_18555,N_16992,N_16377);
xor U18556 (N_18556,N_17545,N_17296);
and U18557 (N_18557,N_17970,N_16977);
and U18558 (N_18558,N_16530,N_16787);
and U18559 (N_18559,N_17020,N_16974);
or U18560 (N_18560,N_16199,N_16090);
nor U18561 (N_18561,N_17870,N_17523);
nand U18562 (N_18562,N_17733,N_16270);
and U18563 (N_18563,N_16952,N_17522);
nand U18564 (N_18564,N_17621,N_16703);
or U18565 (N_18565,N_17332,N_17140);
or U18566 (N_18566,N_16887,N_16042);
nand U18567 (N_18567,N_17228,N_16623);
nor U18568 (N_18568,N_17546,N_16733);
or U18569 (N_18569,N_16126,N_16780);
nand U18570 (N_18570,N_17457,N_17329);
nand U18571 (N_18571,N_17517,N_16202);
nand U18572 (N_18572,N_17585,N_17433);
nor U18573 (N_18573,N_16997,N_17486);
or U18574 (N_18574,N_17437,N_16072);
and U18575 (N_18575,N_16968,N_16665);
xnor U18576 (N_18576,N_17380,N_16655);
xor U18577 (N_18577,N_16353,N_16299);
nor U18578 (N_18578,N_17199,N_16960);
nor U18579 (N_18579,N_17049,N_16529);
nor U18580 (N_18580,N_16634,N_16018);
or U18581 (N_18581,N_17019,N_16060);
or U18582 (N_18582,N_16533,N_16522);
nor U18583 (N_18583,N_17558,N_17544);
xnor U18584 (N_18584,N_16588,N_17218);
nor U18585 (N_18585,N_17711,N_16757);
xor U18586 (N_18586,N_16944,N_17273);
nand U18587 (N_18587,N_16784,N_16128);
and U18588 (N_18588,N_17306,N_17960);
or U18589 (N_18589,N_16164,N_16105);
xnor U18590 (N_18590,N_17309,N_17779);
nand U18591 (N_18591,N_17909,N_16633);
or U18592 (N_18592,N_16236,N_17006);
and U18593 (N_18593,N_17958,N_16207);
xor U18594 (N_18594,N_16031,N_17509);
nand U18595 (N_18595,N_16983,N_17403);
or U18596 (N_18596,N_16303,N_17130);
nand U18597 (N_18597,N_17037,N_17659);
or U18598 (N_18598,N_16732,N_17882);
nand U18599 (N_18599,N_17910,N_17453);
nor U18600 (N_18600,N_17017,N_17321);
xnor U18601 (N_18601,N_16081,N_16368);
or U18602 (N_18602,N_17884,N_17109);
xor U18603 (N_18603,N_16246,N_17617);
nand U18604 (N_18604,N_16364,N_16492);
and U18605 (N_18605,N_17706,N_16471);
xnor U18606 (N_18606,N_17203,N_16708);
nand U18607 (N_18607,N_16216,N_17341);
nor U18608 (N_18608,N_16523,N_17272);
xor U18609 (N_18609,N_17776,N_16730);
xnor U18610 (N_18610,N_17732,N_16254);
xnor U18611 (N_18611,N_16151,N_16715);
and U18612 (N_18612,N_16582,N_16893);
or U18613 (N_18613,N_16422,N_17180);
or U18614 (N_18614,N_16851,N_16001);
nand U18615 (N_18615,N_16026,N_16145);
nor U18616 (N_18616,N_17098,N_17146);
and U18617 (N_18617,N_16307,N_17956);
xor U18618 (N_18618,N_16382,N_16568);
nand U18619 (N_18619,N_16430,N_16837);
and U18620 (N_18620,N_16801,N_16617);
nor U18621 (N_18621,N_17895,N_17849);
nand U18622 (N_18622,N_16161,N_16826);
nand U18623 (N_18623,N_17178,N_16381);
or U18624 (N_18624,N_16809,N_16178);
or U18625 (N_18625,N_17573,N_16982);
nand U18626 (N_18626,N_17727,N_17961);
or U18627 (N_18627,N_16940,N_17765);
and U18628 (N_18628,N_16225,N_16962);
nand U18629 (N_18629,N_17157,N_17359);
and U18630 (N_18630,N_16640,N_17424);
nand U18631 (N_18631,N_16059,N_16644);
and U18632 (N_18632,N_16763,N_16739);
nand U18633 (N_18633,N_16506,N_16129);
or U18634 (N_18634,N_17947,N_17474);
or U18635 (N_18635,N_17326,N_17934);
or U18636 (N_18636,N_16375,N_17115);
xor U18637 (N_18637,N_17993,N_16704);
or U18638 (N_18638,N_16869,N_17242);
or U18639 (N_18639,N_16440,N_17596);
or U18640 (N_18640,N_16205,N_17762);
or U18641 (N_18641,N_16649,N_17093);
and U18642 (N_18642,N_17011,N_17231);
nor U18643 (N_18643,N_17367,N_17574);
and U18644 (N_18644,N_17432,N_17409);
nor U18645 (N_18645,N_16424,N_17835);
xnor U18646 (N_18646,N_17061,N_16735);
nor U18647 (N_18647,N_17443,N_16690);
and U18648 (N_18648,N_16174,N_17212);
nand U18649 (N_18649,N_16527,N_16651);
nor U18650 (N_18650,N_16511,N_17035);
and U18651 (N_18651,N_17629,N_16966);
nor U18652 (N_18652,N_16936,N_17464);
or U18653 (N_18653,N_17699,N_16175);
and U18654 (N_18654,N_17259,N_16187);
nand U18655 (N_18655,N_16348,N_16185);
and U18656 (N_18656,N_16127,N_16107);
or U18657 (N_18657,N_16620,N_17915);
or U18658 (N_18658,N_17124,N_16741);
or U18659 (N_18659,N_17822,N_17044);
nor U18660 (N_18660,N_16776,N_16850);
or U18661 (N_18661,N_17952,N_17681);
or U18662 (N_18662,N_16980,N_16282);
nor U18663 (N_18663,N_17429,N_17709);
nor U18664 (N_18664,N_16629,N_16395);
nor U18665 (N_18665,N_17138,N_17925);
xnor U18666 (N_18666,N_16698,N_16610);
and U18667 (N_18667,N_17032,N_17334);
or U18668 (N_18668,N_17969,N_16378);
nor U18669 (N_18669,N_16280,N_17484);
and U18670 (N_18670,N_17582,N_16321);
nor U18671 (N_18671,N_17976,N_17491);
or U18672 (N_18672,N_17324,N_17315);
nand U18673 (N_18673,N_16769,N_16590);
or U18674 (N_18674,N_17476,N_17398);
or U18675 (N_18675,N_17637,N_16774);
nor U18676 (N_18676,N_17449,N_16495);
xnor U18677 (N_18677,N_16542,N_16016);
or U18678 (N_18678,N_16643,N_16407);
and U18679 (N_18679,N_16947,N_16773);
nor U18680 (N_18680,N_16686,N_16118);
nor U18681 (N_18681,N_16462,N_17295);
xnor U18682 (N_18682,N_16574,N_16545);
or U18683 (N_18683,N_16832,N_17913);
or U18684 (N_18684,N_17083,N_17258);
nor U18685 (N_18685,N_17750,N_17463);
nand U18686 (N_18686,N_17058,N_16699);
nand U18687 (N_18687,N_17357,N_16146);
or U18688 (N_18688,N_16345,N_17369);
nand U18689 (N_18689,N_17505,N_16442);
nor U18690 (N_18690,N_17557,N_16203);
nand U18691 (N_18691,N_16411,N_17676);
or U18692 (N_18692,N_16445,N_17493);
and U18693 (N_18693,N_16306,N_16052);
and U18694 (N_18694,N_17244,N_16294);
xnor U18695 (N_18695,N_16103,N_17041);
nor U18696 (N_18696,N_17927,N_17721);
nor U18697 (N_18697,N_17650,N_16350);
and U18698 (N_18698,N_16019,N_16148);
and U18699 (N_18699,N_17362,N_17880);
nand U18700 (N_18700,N_17825,N_17185);
xor U18701 (N_18701,N_16908,N_16870);
and U18702 (N_18702,N_16724,N_17408);
or U18703 (N_18703,N_16332,N_17356);
nand U18704 (N_18704,N_17289,N_17771);
xnor U18705 (N_18705,N_16243,N_17298);
or U18706 (N_18706,N_16917,N_16881);
xnor U18707 (N_18707,N_16957,N_16840);
xor U18708 (N_18708,N_17472,N_16084);
nor U18709 (N_18709,N_17015,N_16550);
and U18710 (N_18710,N_17914,N_17569);
or U18711 (N_18711,N_17668,N_17325);
xor U18712 (N_18712,N_16223,N_16400);
nand U18713 (N_18713,N_16398,N_16575);
nand U18714 (N_18714,N_17343,N_17638);
or U18715 (N_18715,N_16047,N_17501);
and U18716 (N_18716,N_17025,N_17416);
or U18717 (N_18717,N_17536,N_16701);
and U18718 (N_18718,N_16437,N_17440);
or U18719 (N_18719,N_16534,N_16602);
nand U18720 (N_18720,N_16637,N_17626);
and U18721 (N_18721,N_17857,N_17456);
or U18722 (N_18722,N_17445,N_17365);
and U18723 (N_18723,N_16323,N_16967);
nor U18724 (N_18724,N_16622,N_16419);
and U18725 (N_18725,N_16537,N_17448);
nor U18726 (N_18726,N_17902,N_16706);
or U18727 (N_18727,N_17151,N_17875);
and U18728 (N_18728,N_16002,N_16056);
and U18729 (N_18729,N_17767,N_17112);
nand U18730 (N_18730,N_16463,N_16509);
and U18731 (N_18731,N_16498,N_16162);
or U18732 (N_18732,N_17905,N_17166);
nand U18733 (N_18733,N_17268,N_17103);
and U18734 (N_18734,N_16275,N_16157);
nor U18735 (N_18735,N_16834,N_17450);
and U18736 (N_18736,N_16075,N_17697);
or U18737 (N_18737,N_16489,N_16673);
and U18738 (N_18738,N_16115,N_16768);
or U18739 (N_18739,N_16242,N_16828);
nand U18740 (N_18740,N_17746,N_16475);
or U18741 (N_18741,N_16528,N_16286);
xor U18742 (N_18742,N_16508,N_16758);
xor U18743 (N_18743,N_17904,N_17022);
xor U18744 (N_18744,N_16399,N_17163);
or U18745 (N_18745,N_17131,N_16771);
and U18746 (N_18746,N_17865,N_17527);
nor U18747 (N_18747,N_17974,N_17060);
nand U18748 (N_18748,N_16941,N_17236);
or U18749 (N_18749,N_17997,N_17186);
nor U18750 (N_18750,N_16996,N_16000);
nand U18751 (N_18751,N_17648,N_16197);
or U18752 (N_18752,N_17595,N_17144);
and U18753 (N_18753,N_17892,N_17888);
xnor U18754 (N_18754,N_17532,N_17930);
or U18755 (N_18755,N_16517,N_16034);
or U18756 (N_18756,N_17485,N_16434);
nand U18757 (N_18757,N_16200,N_17281);
xor U18758 (N_18758,N_17752,N_16237);
nor U18759 (N_18759,N_17861,N_16329);
and U18760 (N_18760,N_17063,N_16797);
and U18761 (N_18761,N_16131,N_16547);
nor U18762 (N_18762,N_17876,N_16096);
and U18763 (N_18763,N_17716,N_16626);
nor U18764 (N_18764,N_16488,N_16044);
and U18765 (N_18765,N_16149,N_16749);
or U18766 (N_18766,N_17717,N_17516);
and U18767 (N_18767,N_17195,N_16029);
and U18768 (N_18768,N_16376,N_17335);
nand U18769 (N_18769,N_17690,N_16538);
or U18770 (N_18770,N_17116,N_17587);
and U18771 (N_18771,N_16510,N_16752);
xor U18772 (N_18772,N_16446,N_16288);
and U18773 (N_18773,N_17583,N_16671);
and U18774 (N_18774,N_17830,N_16432);
nand U18775 (N_18775,N_17807,N_16831);
nor U18776 (N_18776,N_16183,N_16935);
xor U18777 (N_18777,N_17327,N_17349);
nor U18778 (N_18778,N_16814,N_16496);
xor U18779 (N_18779,N_17271,N_17317);
or U18780 (N_18780,N_16319,N_17427);
or U18781 (N_18781,N_17817,N_16955);
and U18782 (N_18782,N_17385,N_17778);
xor U18783 (N_18783,N_17141,N_16661);
nor U18784 (N_18784,N_17643,N_17755);
and U18785 (N_18785,N_16363,N_16676);
xnor U18786 (N_18786,N_17452,N_17616);
nand U18787 (N_18787,N_16549,N_17535);
or U18788 (N_18788,N_16427,N_16247);
nand U18789 (N_18789,N_16707,N_16896);
and U18790 (N_18790,N_16721,N_17198);
xnor U18791 (N_18791,N_16872,N_16467);
nor U18792 (N_18792,N_17677,N_16795);
nor U18793 (N_18793,N_16555,N_17052);
xor U18794 (N_18794,N_16287,N_17941);
xnor U18795 (N_18795,N_17168,N_17735);
xor U18796 (N_18796,N_17664,N_17631);
or U18797 (N_18797,N_17552,N_17666);
nor U18798 (N_18798,N_16481,N_16311);
xnor U18799 (N_18799,N_16271,N_16849);
nand U18800 (N_18800,N_17770,N_17889);
nor U18801 (N_18801,N_16362,N_16082);
and U18802 (N_18802,N_17814,N_17483);
or U18803 (N_18803,N_16394,N_16695);
nor U18804 (N_18804,N_16025,N_17397);
and U18805 (N_18805,N_16915,N_16932);
nand U18806 (N_18806,N_16794,N_17867);
nand U18807 (N_18807,N_17286,N_17673);
xor U18808 (N_18808,N_17543,N_16878);
or U18809 (N_18809,N_17331,N_16873);
xor U18810 (N_18810,N_16961,N_17247);
xor U18811 (N_18811,N_17009,N_16263);
or U18812 (N_18812,N_17839,N_17225);
nor U18813 (N_18813,N_16088,N_17016);
nor U18814 (N_18814,N_17922,N_16005);
nand U18815 (N_18815,N_16641,N_17775);
and U18816 (N_18816,N_17045,N_16372);
nor U18817 (N_18817,N_16719,N_16360);
or U18818 (N_18818,N_16720,N_17748);
xor U18819 (N_18819,N_16659,N_16745);
nand U18820 (N_18820,N_17987,N_16085);
or U18821 (N_18821,N_16581,N_17950);
nand U18822 (N_18822,N_17651,N_16444);
or U18823 (N_18823,N_16284,N_17860);
nor U18824 (N_18824,N_16559,N_16976);
or U18825 (N_18825,N_16158,N_17819);
xor U18826 (N_18826,N_16903,N_17988);
and U18827 (N_18827,N_16981,N_16988);
or U18828 (N_18828,N_17276,N_16464);
xor U18829 (N_18829,N_16098,N_16487);
nand U18830 (N_18830,N_16116,N_17054);
xnor U18831 (N_18831,N_17520,N_16738);
nor U18832 (N_18832,N_17128,N_16772);
xnor U18833 (N_18833,N_17965,N_16117);
nand U18834 (N_18834,N_16068,N_17900);
nor U18835 (N_18835,N_17183,N_16595);
nor U18836 (N_18836,N_17561,N_17611);
nand U18837 (N_18837,N_16740,N_16543);
or U18838 (N_18838,N_16176,N_16729);
xor U18839 (N_18839,N_16899,N_16711);
xnor U18840 (N_18840,N_16226,N_16396);
nand U18841 (N_18841,N_16198,N_16576);
nand U18842 (N_18842,N_16518,N_17267);
or U18843 (N_18843,N_17191,N_17114);
and U18844 (N_18844,N_17110,N_17210);
nand U18845 (N_18845,N_17401,N_17235);
xor U18846 (N_18846,N_16638,N_17710);
or U18847 (N_18847,N_16315,N_16700);
xor U18848 (N_18848,N_16300,N_16012);
or U18849 (N_18849,N_17099,N_17789);
nand U18850 (N_18850,N_16261,N_17813);
xor U18851 (N_18851,N_17878,N_16490);
nor U18852 (N_18852,N_17490,N_17442);
xnor U18853 (N_18853,N_17736,N_17077);
or U18854 (N_18854,N_17494,N_17291);
and U18855 (N_18855,N_16689,N_16452);
nor U18856 (N_18856,N_17685,N_16635);
nand U18857 (N_18857,N_17622,N_17248);
and U18858 (N_18858,N_17215,N_16106);
nor U18859 (N_18859,N_17992,N_16092);
nand U18860 (N_18860,N_16779,N_17499);
or U18861 (N_18861,N_16557,N_16494);
nand U18862 (N_18862,N_16566,N_17395);
nand U18863 (N_18863,N_16267,N_16184);
nand U18864 (N_18864,N_17159,N_16838);
xor U18865 (N_18865,N_17572,N_17654);
or U18866 (N_18866,N_16387,N_16882);
or U18867 (N_18867,N_17893,N_16934);
or U18868 (N_18868,N_16544,N_17028);
nand U18869 (N_18869,N_16958,N_16685);
nand U18870 (N_18870,N_17301,N_16927);
nor U18871 (N_18871,N_17415,N_16531);
nand U18872 (N_18872,N_17640,N_17441);
xor U18873 (N_18873,N_17120,N_17122);
nand U18874 (N_18874,N_16894,N_16071);
nand U18875 (N_18875,N_16163,N_17590);
or U18876 (N_18876,N_16539,N_16110);
and U18877 (N_18877,N_16630,N_17420);
nor U18878 (N_18878,N_16474,N_16454);
or U18879 (N_18879,N_16624,N_17226);
and U18880 (N_18880,N_17891,N_17979);
nand U18881 (N_18881,N_16010,N_16954);
nand U18882 (N_18882,N_17538,N_17786);
nand U18883 (N_18883,N_17691,N_17623);
xnor U18884 (N_18884,N_17862,N_17614);
xor U18885 (N_18885,N_16959,N_16310);
nor U18886 (N_18886,N_17853,N_16526);
nor U18887 (N_18887,N_16094,N_17815);
xor U18888 (N_18888,N_17798,N_17653);
and U18889 (N_18889,N_17563,N_17566);
and U18890 (N_18890,N_17740,N_16500);
or U18891 (N_18891,N_16647,N_17874);
nand U18892 (N_18892,N_16351,N_16229);
and U18893 (N_18893,N_16466,N_17055);
or U18894 (N_18894,N_16580,N_17264);
nor U18895 (N_18895,N_16558,N_16033);
xor U18896 (N_18896,N_17787,N_17749);
and U18897 (N_18897,N_16083,N_17065);
nor U18898 (N_18898,N_16614,N_17512);
or U18899 (N_18899,N_17671,N_16585);
nand U18900 (N_18900,N_17580,N_17451);
or U18901 (N_18901,N_16336,N_16865);
or U18902 (N_18902,N_17217,N_16331);
or U18903 (N_18903,N_17984,N_17845);
nor U18904 (N_18904,N_17761,N_17008);
nand U18905 (N_18905,N_16507,N_17313);
or U18906 (N_18906,N_17708,N_17788);
xor U18907 (N_18907,N_17104,N_17202);
nand U18908 (N_18908,N_16309,N_16766);
and U18909 (N_18909,N_16089,N_17981);
and U18910 (N_18910,N_17744,N_16285);
nand U18911 (N_18911,N_16984,N_16652);
nand U18912 (N_18912,N_16513,N_16008);
nor U18913 (N_18913,N_16577,N_16268);
xor U18914 (N_18914,N_16540,N_17204);
or U18915 (N_18915,N_16228,N_17804);
or U18916 (N_18916,N_17728,N_16371);
and U18917 (N_18917,N_16722,N_17076);
and U18918 (N_18918,N_16783,N_16802);
nand U18919 (N_18919,N_17230,N_16871);
nand U18920 (N_18920,N_16049,N_16883);
or U18921 (N_18921,N_17887,N_17946);
or U18922 (N_18922,N_17624,N_16564);
nor U18923 (N_18923,N_17172,N_16402);
or U18924 (N_18924,N_17896,N_16003);
or U18925 (N_18925,N_16888,N_16725);
xor U18926 (N_18926,N_17333,N_17330);
and U18927 (N_18927,N_17488,N_16536);
nand U18928 (N_18928,N_17785,N_16798);
or U18929 (N_18929,N_17279,N_17682);
nor U18930 (N_18930,N_17745,N_17508);
nor U18931 (N_18931,N_17525,N_16751);
xor U18932 (N_18932,N_17391,N_17492);
and U18933 (N_18933,N_16748,N_17592);
xor U18934 (N_18934,N_16408,N_17881);
nand U18935 (N_18935,N_16593,N_16642);
xor U18936 (N_18936,N_16628,N_16969);
nand U18937 (N_18937,N_17123,N_17299);
nor U18938 (N_18938,N_16020,N_17718);
xnor U18939 (N_18939,N_17255,N_16796);
xor U18940 (N_18940,N_17394,N_17001);
nor U18941 (N_18941,N_16521,N_16805);
and U18942 (N_18942,N_17057,N_17940);
nand U18943 (N_18943,N_17790,N_16099);
xor U18944 (N_18944,N_16412,N_16366);
xnor U18945 (N_18945,N_17933,N_16077);
or U18946 (N_18946,N_17551,N_16390);
nor U18947 (N_18947,N_17951,N_16913);
nor U18948 (N_18948,N_16405,N_17743);
or U18949 (N_18949,N_17955,N_16341);
and U18950 (N_18950,N_17262,N_16230);
xnor U18951 (N_18951,N_17625,N_17260);
or U18952 (N_18952,N_17376,N_17455);
or U18953 (N_18953,N_16132,N_16592);
and U18954 (N_18954,N_17405,N_16928);
or U18955 (N_18955,N_16240,N_16989);
and U18956 (N_18956,N_16793,N_16211);
nand U18957 (N_18957,N_16095,N_16028);
nand U18958 (N_18958,N_17565,N_17838);
or U18959 (N_18959,N_16491,N_17239);
and U18960 (N_18960,N_17549,N_16349);
nor U18961 (N_18961,N_16006,N_17487);
or U18962 (N_18962,N_16571,N_17912);
nor U18963 (N_18963,N_17107,N_16727);
xor U18964 (N_18964,N_16333,N_16057);
and U18965 (N_18965,N_16605,N_16314);
xnor U18966 (N_18966,N_17338,N_16866);
nand U18967 (N_18967,N_17642,N_17620);
and U18968 (N_18968,N_16283,N_17221);
and U18969 (N_18969,N_16453,N_17048);
nor U18970 (N_18970,N_17461,N_16014);
nand U18971 (N_18971,N_16169,N_16004);
xnor U18972 (N_18972,N_17270,N_16948);
or U18973 (N_18973,N_17929,N_16978);
or U18974 (N_18974,N_16416,N_16045);
and U18975 (N_18975,N_16688,N_16929);
or U18976 (N_18976,N_17233,N_17027);
nand U18977 (N_18977,N_16221,N_16343);
and U18978 (N_18978,N_17627,N_17024);
nor U18979 (N_18979,N_17554,N_17908);
nand U18980 (N_18980,N_16994,N_16860);
or U18981 (N_18981,N_16930,N_16069);
and U18982 (N_18982,N_17713,N_17847);
nor U18983 (N_18983,N_16369,N_17310);
nand U18984 (N_18984,N_16073,N_17649);
or U18985 (N_18985,N_17383,N_17040);
or U18986 (N_18986,N_16718,N_17646);
and U18987 (N_18987,N_17704,N_16611);
xnor U18988 (N_18988,N_16938,N_17689);
nor U18989 (N_18989,N_17836,N_17414);
nand U18990 (N_18990,N_16999,N_16181);
nor U18991 (N_18991,N_17458,N_17810);
xnor U18992 (N_18992,N_16374,N_16925);
xor U18993 (N_18993,N_16217,N_17591);
nand U18994 (N_18994,N_17695,N_16021);
and U18995 (N_18995,N_17820,N_16326);
and U18996 (N_18996,N_17208,N_17593);
or U18997 (N_18997,N_16168,N_16404);
and U18998 (N_18998,N_17430,N_17374);
nor U18999 (N_18999,N_17471,N_16438);
xnor U19000 (N_19000,N_16316,N_17596);
and U19001 (N_19001,N_17225,N_17902);
nor U19002 (N_19002,N_17967,N_16723);
xor U19003 (N_19003,N_16481,N_16723);
or U19004 (N_19004,N_16687,N_17588);
nor U19005 (N_19005,N_17687,N_17566);
or U19006 (N_19006,N_17893,N_16241);
nand U19007 (N_19007,N_16402,N_17117);
nand U19008 (N_19008,N_16967,N_17340);
nor U19009 (N_19009,N_17521,N_16256);
nor U19010 (N_19010,N_16597,N_16179);
and U19011 (N_19011,N_16001,N_16690);
and U19012 (N_19012,N_16784,N_16276);
nor U19013 (N_19013,N_16181,N_16463);
nor U19014 (N_19014,N_17375,N_16352);
xnor U19015 (N_19015,N_16702,N_16013);
nor U19016 (N_19016,N_17032,N_16877);
nor U19017 (N_19017,N_17703,N_16423);
and U19018 (N_19018,N_16263,N_17854);
nand U19019 (N_19019,N_16968,N_17779);
or U19020 (N_19020,N_16384,N_17882);
xor U19021 (N_19021,N_16184,N_17434);
or U19022 (N_19022,N_17290,N_16024);
nand U19023 (N_19023,N_17428,N_16532);
or U19024 (N_19024,N_17483,N_16510);
nor U19025 (N_19025,N_16293,N_16138);
and U19026 (N_19026,N_16796,N_17189);
and U19027 (N_19027,N_17289,N_16916);
and U19028 (N_19028,N_16818,N_17644);
xor U19029 (N_19029,N_16945,N_16764);
nor U19030 (N_19030,N_17809,N_16960);
or U19031 (N_19031,N_17805,N_16673);
nor U19032 (N_19032,N_16169,N_17846);
nand U19033 (N_19033,N_17794,N_17553);
xnor U19034 (N_19034,N_17463,N_17602);
xnor U19035 (N_19035,N_17521,N_16674);
nand U19036 (N_19036,N_17120,N_16854);
and U19037 (N_19037,N_17048,N_16417);
xnor U19038 (N_19038,N_16940,N_17922);
and U19039 (N_19039,N_16886,N_16653);
xnor U19040 (N_19040,N_16990,N_17468);
nand U19041 (N_19041,N_17213,N_16026);
nand U19042 (N_19042,N_16447,N_17377);
and U19043 (N_19043,N_16502,N_17065);
and U19044 (N_19044,N_16061,N_17630);
nand U19045 (N_19045,N_17083,N_17232);
or U19046 (N_19046,N_17370,N_17283);
and U19047 (N_19047,N_17619,N_16052);
xor U19048 (N_19048,N_16748,N_16053);
and U19049 (N_19049,N_17132,N_17975);
and U19050 (N_19050,N_16379,N_17833);
xnor U19051 (N_19051,N_17580,N_16442);
or U19052 (N_19052,N_17275,N_16423);
xor U19053 (N_19053,N_16903,N_17090);
or U19054 (N_19054,N_16918,N_16356);
or U19055 (N_19055,N_16196,N_16083);
or U19056 (N_19056,N_17765,N_16540);
nor U19057 (N_19057,N_16996,N_16453);
nor U19058 (N_19058,N_16167,N_17312);
nand U19059 (N_19059,N_17617,N_16565);
xor U19060 (N_19060,N_17513,N_16877);
and U19061 (N_19061,N_16587,N_16924);
nor U19062 (N_19062,N_17581,N_16946);
or U19063 (N_19063,N_16631,N_16603);
or U19064 (N_19064,N_17284,N_16890);
or U19065 (N_19065,N_16049,N_16847);
nor U19066 (N_19066,N_16148,N_16336);
xor U19067 (N_19067,N_16631,N_17750);
nor U19068 (N_19068,N_17106,N_17271);
nand U19069 (N_19069,N_16193,N_16787);
or U19070 (N_19070,N_16265,N_16758);
nand U19071 (N_19071,N_17281,N_17923);
nor U19072 (N_19072,N_16895,N_16327);
and U19073 (N_19073,N_16762,N_17793);
nand U19074 (N_19074,N_17493,N_16898);
xor U19075 (N_19075,N_17657,N_16191);
nor U19076 (N_19076,N_17866,N_16185);
and U19077 (N_19077,N_16833,N_16098);
and U19078 (N_19078,N_16796,N_16885);
or U19079 (N_19079,N_16373,N_17113);
xor U19080 (N_19080,N_16833,N_17761);
nand U19081 (N_19081,N_17049,N_17079);
and U19082 (N_19082,N_17000,N_17926);
or U19083 (N_19083,N_17591,N_16341);
nor U19084 (N_19084,N_17705,N_16622);
nand U19085 (N_19085,N_16652,N_16683);
and U19086 (N_19086,N_16895,N_16103);
xnor U19087 (N_19087,N_17293,N_16548);
and U19088 (N_19088,N_16140,N_16207);
and U19089 (N_19089,N_17763,N_17933);
or U19090 (N_19090,N_17815,N_17452);
and U19091 (N_19091,N_16864,N_16334);
xnor U19092 (N_19092,N_16785,N_16723);
nor U19093 (N_19093,N_17765,N_17822);
or U19094 (N_19094,N_17567,N_16334);
nor U19095 (N_19095,N_17155,N_16976);
and U19096 (N_19096,N_16505,N_16431);
nor U19097 (N_19097,N_16215,N_17604);
and U19098 (N_19098,N_17852,N_16403);
and U19099 (N_19099,N_17821,N_16109);
or U19100 (N_19100,N_17771,N_16924);
nand U19101 (N_19101,N_17996,N_17270);
nand U19102 (N_19102,N_17772,N_17452);
or U19103 (N_19103,N_17294,N_17651);
or U19104 (N_19104,N_17241,N_17477);
xnor U19105 (N_19105,N_17208,N_17369);
xnor U19106 (N_19106,N_17749,N_16096);
nand U19107 (N_19107,N_17919,N_16747);
and U19108 (N_19108,N_17304,N_16220);
xnor U19109 (N_19109,N_17673,N_17414);
nor U19110 (N_19110,N_16458,N_17360);
or U19111 (N_19111,N_16975,N_17063);
nor U19112 (N_19112,N_17309,N_16166);
and U19113 (N_19113,N_16726,N_17321);
nand U19114 (N_19114,N_16729,N_17266);
nand U19115 (N_19115,N_17842,N_17406);
nor U19116 (N_19116,N_17079,N_17971);
and U19117 (N_19117,N_17658,N_16978);
nand U19118 (N_19118,N_16944,N_17020);
nor U19119 (N_19119,N_17961,N_16853);
and U19120 (N_19120,N_16772,N_16716);
nor U19121 (N_19121,N_17502,N_16487);
nand U19122 (N_19122,N_17023,N_16721);
and U19123 (N_19123,N_17855,N_16987);
nor U19124 (N_19124,N_16568,N_17162);
nand U19125 (N_19125,N_16973,N_17542);
xor U19126 (N_19126,N_16877,N_16624);
and U19127 (N_19127,N_16059,N_16065);
nand U19128 (N_19128,N_16873,N_17504);
and U19129 (N_19129,N_17060,N_16221);
or U19130 (N_19130,N_17198,N_17201);
or U19131 (N_19131,N_17932,N_16254);
nor U19132 (N_19132,N_17602,N_17994);
or U19133 (N_19133,N_16276,N_17966);
or U19134 (N_19134,N_17852,N_16142);
or U19135 (N_19135,N_17361,N_16050);
and U19136 (N_19136,N_16117,N_17329);
or U19137 (N_19137,N_16103,N_17585);
xor U19138 (N_19138,N_17818,N_16796);
xor U19139 (N_19139,N_17733,N_16328);
or U19140 (N_19140,N_16054,N_16333);
or U19141 (N_19141,N_16387,N_16876);
nand U19142 (N_19142,N_16612,N_17538);
nor U19143 (N_19143,N_16358,N_16033);
xnor U19144 (N_19144,N_17368,N_16326);
xor U19145 (N_19145,N_16707,N_16875);
nor U19146 (N_19146,N_17522,N_17067);
and U19147 (N_19147,N_16893,N_16847);
xor U19148 (N_19148,N_17226,N_16445);
or U19149 (N_19149,N_16940,N_17441);
or U19150 (N_19150,N_16557,N_16228);
xnor U19151 (N_19151,N_17514,N_17789);
or U19152 (N_19152,N_17986,N_16440);
nand U19153 (N_19153,N_17051,N_16115);
and U19154 (N_19154,N_17951,N_16445);
nor U19155 (N_19155,N_17995,N_17343);
nand U19156 (N_19156,N_16795,N_17099);
or U19157 (N_19157,N_16758,N_17098);
nand U19158 (N_19158,N_17836,N_17683);
xor U19159 (N_19159,N_17544,N_17219);
nor U19160 (N_19160,N_16367,N_16478);
and U19161 (N_19161,N_17149,N_16480);
nor U19162 (N_19162,N_17646,N_17894);
nor U19163 (N_19163,N_16062,N_16048);
and U19164 (N_19164,N_17102,N_17784);
nand U19165 (N_19165,N_17783,N_17024);
nand U19166 (N_19166,N_16877,N_17072);
nor U19167 (N_19167,N_17819,N_16638);
and U19168 (N_19168,N_16412,N_16876);
and U19169 (N_19169,N_16222,N_17997);
and U19170 (N_19170,N_16279,N_16024);
nand U19171 (N_19171,N_17151,N_16225);
nor U19172 (N_19172,N_16300,N_17985);
xnor U19173 (N_19173,N_17724,N_17765);
or U19174 (N_19174,N_16577,N_16819);
and U19175 (N_19175,N_16780,N_17151);
nand U19176 (N_19176,N_17570,N_17143);
nor U19177 (N_19177,N_17455,N_16059);
nor U19178 (N_19178,N_16815,N_16421);
xnor U19179 (N_19179,N_16381,N_17230);
nor U19180 (N_19180,N_16413,N_17842);
nand U19181 (N_19181,N_16716,N_17373);
and U19182 (N_19182,N_16250,N_17538);
or U19183 (N_19183,N_17698,N_17783);
nand U19184 (N_19184,N_17035,N_17790);
and U19185 (N_19185,N_17877,N_16105);
or U19186 (N_19186,N_17933,N_17532);
xor U19187 (N_19187,N_16933,N_17564);
nor U19188 (N_19188,N_16617,N_17143);
or U19189 (N_19189,N_17350,N_17695);
nand U19190 (N_19190,N_17781,N_17338);
or U19191 (N_19191,N_17782,N_16538);
and U19192 (N_19192,N_17097,N_16453);
and U19193 (N_19193,N_16669,N_16985);
and U19194 (N_19194,N_17881,N_17050);
nand U19195 (N_19195,N_16606,N_16639);
nor U19196 (N_19196,N_16484,N_16165);
and U19197 (N_19197,N_17801,N_17344);
nand U19198 (N_19198,N_17493,N_16433);
nand U19199 (N_19199,N_17947,N_16214);
or U19200 (N_19200,N_16597,N_17937);
nand U19201 (N_19201,N_17876,N_17149);
and U19202 (N_19202,N_16487,N_16161);
and U19203 (N_19203,N_16239,N_17660);
xnor U19204 (N_19204,N_16539,N_17786);
xor U19205 (N_19205,N_17525,N_16542);
nand U19206 (N_19206,N_16951,N_17339);
nor U19207 (N_19207,N_16146,N_16407);
nor U19208 (N_19208,N_16373,N_17163);
xor U19209 (N_19209,N_16335,N_17637);
or U19210 (N_19210,N_16102,N_17464);
and U19211 (N_19211,N_17536,N_16196);
and U19212 (N_19212,N_17513,N_16523);
xor U19213 (N_19213,N_16289,N_16006);
and U19214 (N_19214,N_16878,N_16167);
nor U19215 (N_19215,N_16673,N_16104);
nand U19216 (N_19216,N_17467,N_16912);
nand U19217 (N_19217,N_17782,N_17607);
nor U19218 (N_19218,N_16627,N_17111);
and U19219 (N_19219,N_16429,N_17247);
and U19220 (N_19220,N_17454,N_16498);
or U19221 (N_19221,N_17074,N_16919);
xor U19222 (N_19222,N_17859,N_17641);
nand U19223 (N_19223,N_16801,N_17867);
nand U19224 (N_19224,N_17243,N_17617);
or U19225 (N_19225,N_17724,N_17590);
and U19226 (N_19226,N_17171,N_16761);
nand U19227 (N_19227,N_17888,N_16436);
or U19228 (N_19228,N_17043,N_17948);
xor U19229 (N_19229,N_17985,N_17401);
or U19230 (N_19230,N_17544,N_17723);
and U19231 (N_19231,N_16916,N_17953);
or U19232 (N_19232,N_17956,N_17959);
and U19233 (N_19233,N_16635,N_17173);
nor U19234 (N_19234,N_17386,N_17110);
and U19235 (N_19235,N_17827,N_16570);
xor U19236 (N_19236,N_16253,N_16627);
nor U19237 (N_19237,N_16736,N_17891);
and U19238 (N_19238,N_16942,N_16409);
or U19239 (N_19239,N_16651,N_17608);
and U19240 (N_19240,N_17252,N_17649);
and U19241 (N_19241,N_17161,N_17533);
nor U19242 (N_19242,N_17848,N_16128);
and U19243 (N_19243,N_17862,N_16408);
and U19244 (N_19244,N_16902,N_16377);
nor U19245 (N_19245,N_17666,N_16547);
or U19246 (N_19246,N_16373,N_17532);
nand U19247 (N_19247,N_17270,N_16773);
nand U19248 (N_19248,N_17190,N_17275);
xor U19249 (N_19249,N_17604,N_16070);
or U19250 (N_19250,N_16743,N_17566);
nand U19251 (N_19251,N_17776,N_16915);
nor U19252 (N_19252,N_17705,N_16375);
nand U19253 (N_19253,N_17475,N_16070);
nor U19254 (N_19254,N_17003,N_16166);
nor U19255 (N_19255,N_16830,N_16530);
xnor U19256 (N_19256,N_17932,N_17057);
or U19257 (N_19257,N_17563,N_17961);
or U19258 (N_19258,N_16942,N_17952);
and U19259 (N_19259,N_16311,N_16553);
and U19260 (N_19260,N_16101,N_17263);
and U19261 (N_19261,N_17875,N_16142);
nor U19262 (N_19262,N_17686,N_17216);
nor U19263 (N_19263,N_16649,N_16687);
xnor U19264 (N_19264,N_16828,N_16333);
nand U19265 (N_19265,N_16179,N_16984);
nor U19266 (N_19266,N_16959,N_17835);
nand U19267 (N_19267,N_16768,N_16943);
and U19268 (N_19268,N_16181,N_17556);
nand U19269 (N_19269,N_17856,N_16322);
nand U19270 (N_19270,N_17873,N_16048);
nor U19271 (N_19271,N_17759,N_17092);
or U19272 (N_19272,N_17512,N_17693);
and U19273 (N_19273,N_16722,N_16698);
xor U19274 (N_19274,N_17084,N_17495);
or U19275 (N_19275,N_17194,N_17597);
or U19276 (N_19276,N_17099,N_16255);
xnor U19277 (N_19277,N_17697,N_16538);
xor U19278 (N_19278,N_17695,N_16368);
or U19279 (N_19279,N_16529,N_17101);
nor U19280 (N_19280,N_17848,N_17096);
nor U19281 (N_19281,N_17277,N_16694);
or U19282 (N_19282,N_16306,N_17107);
nand U19283 (N_19283,N_16512,N_17325);
nand U19284 (N_19284,N_16540,N_16107);
nand U19285 (N_19285,N_16040,N_17033);
xor U19286 (N_19286,N_16662,N_17348);
nor U19287 (N_19287,N_17613,N_16400);
xor U19288 (N_19288,N_16901,N_17513);
nor U19289 (N_19289,N_17791,N_16754);
xnor U19290 (N_19290,N_16917,N_17899);
or U19291 (N_19291,N_17229,N_16495);
and U19292 (N_19292,N_16998,N_17912);
or U19293 (N_19293,N_16888,N_16247);
and U19294 (N_19294,N_16666,N_16611);
nand U19295 (N_19295,N_16958,N_17826);
and U19296 (N_19296,N_17984,N_16962);
nand U19297 (N_19297,N_17955,N_17423);
or U19298 (N_19298,N_16659,N_16418);
and U19299 (N_19299,N_17838,N_17986);
or U19300 (N_19300,N_16497,N_17936);
or U19301 (N_19301,N_17512,N_17058);
nand U19302 (N_19302,N_16586,N_17183);
and U19303 (N_19303,N_16216,N_17235);
and U19304 (N_19304,N_16068,N_17384);
nand U19305 (N_19305,N_16619,N_17510);
nand U19306 (N_19306,N_17946,N_17643);
or U19307 (N_19307,N_17613,N_16162);
and U19308 (N_19308,N_17314,N_16517);
or U19309 (N_19309,N_16048,N_17596);
xor U19310 (N_19310,N_17993,N_17077);
xor U19311 (N_19311,N_16151,N_16837);
nor U19312 (N_19312,N_17880,N_17150);
and U19313 (N_19313,N_17901,N_17995);
nand U19314 (N_19314,N_17342,N_16435);
or U19315 (N_19315,N_17075,N_17830);
nand U19316 (N_19316,N_16351,N_17010);
xor U19317 (N_19317,N_17741,N_16800);
xnor U19318 (N_19318,N_16020,N_17449);
xor U19319 (N_19319,N_17561,N_17296);
and U19320 (N_19320,N_17390,N_17182);
xor U19321 (N_19321,N_16470,N_16044);
nand U19322 (N_19322,N_16505,N_17939);
nor U19323 (N_19323,N_16666,N_16456);
nor U19324 (N_19324,N_17259,N_17509);
or U19325 (N_19325,N_16980,N_16559);
and U19326 (N_19326,N_17888,N_17418);
or U19327 (N_19327,N_17325,N_16848);
or U19328 (N_19328,N_17127,N_17303);
or U19329 (N_19329,N_17819,N_17817);
xor U19330 (N_19330,N_17094,N_17633);
or U19331 (N_19331,N_17954,N_16814);
nor U19332 (N_19332,N_16589,N_16269);
or U19333 (N_19333,N_17210,N_16069);
xnor U19334 (N_19334,N_16082,N_17149);
xnor U19335 (N_19335,N_16443,N_16286);
and U19336 (N_19336,N_17963,N_16976);
and U19337 (N_19337,N_16131,N_16093);
and U19338 (N_19338,N_17765,N_16663);
and U19339 (N_19339,N_16266,N_17904);
nand U19340 (N_19340,N_17842,N_17377);
and U19341 (N_19341,N_16670,N_17608);
or U19342 (N_19342,N_16570,N_17219);
or U19343 (N_19343,N_16669,N_17265);
xnor U19344 (N_19344,N_16773,N_17320);
nand U19345 (N_19345,N_17430,N_17057);
or U19346 (N_19346,N_16284,N_17964);
nand U19347 (N_19347,N_17330,N_16827);
and U19348 (N_19348,N_16875,N_17912);
xor U19349 (N_19349,N_16179,N_16720);
and U19350 (N_19350,N_16769,N_16719);
nand U19351 (N_19351,N_16605,N_16975);
xnor U19352 (N_19352,N_17606,N_17801);
nand U19353 (N_19353,N_16940,N_16651);
and U19354 (N_19354,N_16096,N_17599);
and U19355 (N_19355,N_17017,N_16069);
and U19356 (N_19356,N_17164,N_17052);
nand U19357 (N_19357,N_17208,N_16302);
or U19358 (N_19358,N_17470,N_16634);
nor U19359 (N_19359,N_17660,N_17571);
or U19360 (N_19360,N_17037,N_16235);
nor U19361 (N_19361,N_16476,N_16658);
nor U19362 (N_19362,N_17692,N_17832);
nand U19363 (N_19363,N_17212,N_16044);
nand U19364 (N_19364,N_17117,N_17381);
nor U19365 (N_19365,N_16901,N_16613);
or U19366 (N_19366,N_17020,N_16129);
or U19367 (N_19367,N_17812,N_16226);
or U19368 (N_19368,N_16004,N_16278);
nor U19369 (N_19369,N_16404,N_17555);
nand U19370 (N_19370,N_17805,N_16982);
nor U19371 (N_19371,N_17061,N_17257);
xnor U19372 (N_19372,N_16858,N_16382);
xnor U19373 (N_19373,N_16289,N_17841);
or U19374 (N_19374,N_17735,N_17989);
xor U19375 (N_19375,N_16665,N_16905);
and U19376 (N_19376,N_17215,N_16304);
nand U19377 (N_19377,N_16764,N_17337);
and U19378 (N_19378,N_17178,N_16112);
nor U19379 (N_19379,N_16048,N_16343);
or U19380 (N_19380,N_16405,N_17620);
and U19381 (N_19381,N_16818,N_17269);
nand U19382 (N_19382,N_16961,N_17119);
or U19383 (N_19383,N_17691,N_16912);
and U19384 (N_19384,N_16075,N_17221);
nand U19385 (N_19385,N_16991,N_16705);
and U19386 (N_19386,N_16738,N_16935);
nor U19387 (N_19387,N_16671,N_16319);
nand U19388 (N_19388,N_17367,N_17885);
or U19389 (N_19389,N_16586,N_16448);
nand U19390 (N_19390,N_16797,N_17254);
and U19391 (N_19391,N_17263,N_16037);
or U19392 (N_19392,N_16789,N_17219);
nand U19393 (N_19393,N_16463,N_17636);
nor U19394 (N_19394,N_16735,N_16933);
or U19395 (N_19395,N_16332,N_17804);
nand U19396 (N_19396,N_16175,N_17295);
nand U19397 (N_19397,N_16630,N_16784);
nor U19398 (N_19398,N_17465,N_16848);
and U19399 (N_19399,N_17411,N_16067);
or U19400 (N_19400,N_16616,N_17761);
xnor U19401 (N_19401,N_16496,N_17366);
nor U19402 (N_19402,N_17862,N_16110);
nand U19403 (N_19403,N_17125,N_17769);
nor U19404 (N_19404,N_17604,N_17570);
nand U19405 (N_19405,N_16535,N_17429);
or U19406 (N_19406,N_16787,N_16018);
xor U19407 (N_19407,N_16932,N_17178);
nor U19408 (N_19408,N_16993,N_16062);
or U19409 (N_19409,N_16278,N_16303);
nor U19410 (N_19410,N_17466,N_17009);
nor U19411 (N_19411,N_17651,N_16217);
or U19412 (N_19412,N_17852,N_16518);
or U19413 (N_19413,N_17511,N_16199);
nand U19414 (N_19414,N_17916,N_17975);
xnor U19415 (N_19415,N_16823,N_16938);
xnor U19416 (N_19416,N_17515,N_17801);
and U19417 (N_19417,N_17003,N_16659);
and U19418 (N_19418,N_16147,N_17149);
xor U19419 (N_19419,N_16535,N_16599);
xnor U19420 (N_19420,N_17818,N_17094);
nand U19421 (N_19421,N_17006,N_17451);
nand U19422 (N_19422,N_17271,N_16931);
nor U19423 (N_19423,N_17534,N_16045);
xnor U19424 (N_19424,N_17053,N_16072);
and U19425 (N_19425,N_17204,N_16263);
or U19426 (N_19426,N_17712,N_17750);
or U19427 (N_19427,N_16941,N_17093);
nor U19428 (N_19428,N_16602,N_17113);
nor U19429 (N_19429,N_17248,N_17109);
xnor U19430 (N_19430,N_16445,N_17035);
nand U19431 (N_19431,N_17685,N_17823);
xnor U19432 (N_19432,N_16688,N_16542);
or U19433 (N_19433,N_17916,N_17425);
nor U19434 (N_19434,N_16776,N_16308);
and U19435 (N_19435,N_16972,N_16994);
nand U19436 (N_19436,N_16453,N_16179);
nor U19437 (N_19437,N_17527,N_17793);
and U19438 (N_19438,N_17402,N_16058);
and U19439 (N_19439,N_16006,N_17845);
nor U19440 (N_19440,N_17480,N_16323);
nor U19441 (N_19441,N_16985,N_16788);
and U19442 (N_19442,N_17085,N_16176);
nor U19443 (N_19443,N_16033,N_17936);
nor U19444 (N_19444,N_16548,N_16686);
nor U19445 (N_19445,N_16944,N_16784);
and U19446 (N_19446,N_17502,N_16262);
xor U19447 (N_19447,N_16721,N_17796);
nand U19448 (N_19448,N_17793,N_17761);
or U19449 (N_19449,N_16404,N_16582);
xnor U19450 (N_19450,N_16691,N_16379);
or U19451 (N_19451,N_16027,N_17960);
nor U19452 (N_19452,N_17763,N_17975);
nand U19453 (N_19453,N_16527,N_17582);
nor U19454 (N_19454,N_16823,N_17218);
nor U19455 (N_19455,N_17260,N_17440);
nand U19456 (N_19456,N_16249,N_16642);
nor U19457 (N_19457,N_17792,N_16969);
and U19458 (N_19458,N_16577,N_16254);
nor U19459 (N_19459,N_17875,N_17574);
nor U19460 (N_19460,N_17450,N_16081);
nor U19461 (N_19461,N_17860,N_16348);
or U19462 (N_19462,N_16797,N_16778);
nand U19463 (N_19463,N_16535,N_16953);
or U19464 (N_19464,N_17615,N_17129);
nor U19465 (N_19465,N_17610,N_16956);
xor U19466 (N_19466,N_16246,N_16322);
and U19467 (N_19467,N_17020,N_17446);
xnor U19468 (N_19468,N_16499,N_17303);
nand U19469 (N_19469,N_17161,N_16426);
and U19470 (N_19470,N_17732,N_16117);
nor U19471 (N_19471,N_16912,N_16873);
nor U19472 (N_19472,N_16174,N_16633);
nor U19473 (N_19473,N_17045,N_16178);
nor U19474 (N_19474,N_16759,N_17645);
nand U19475 (N_19475,N_17219,N_16300);
nor U19476 (N_19476,N_16509,N_16102);
or U19477 (N_19477,N_16199,N_17015);
nand U19478 (N_19478,N_17118,N_17558);
nor U19479 (N_19479,N_17224,N_17643);
xnor U19480 (N_19480,N_17617,N_17553);
xor U19481 (N_19481,N_17031,N_16277);
and U19482 (N_19482,N_16390,N_17912);
nor U19483 (N_19483,N_17192,N_17466);
or U19484 (N_19484,N_17036,N_16462);
nand U19485 (N_19485,N_16987,N_16892);
or U19486 (N_19486,N_16068,N_16100);
and U19487 (N_19487,N_16195,N_17940);
or U19488 (N_19488,N_16961,N_17877);
xnor U19489 (N_19489,N_16932,N_16457);
nand U19490 (N_19490,N_17475,N_16657);
xor U19491 (N_19491,N_16379,N_16262);
nand U19492 (N_19492,N_17204,N_16234);
nand U19493 (N_19493,N_16730,N_16753);
xor U19494 (N_19494,N_17960,N_16638);
or U19495 (N_19495,N_16785,N_17584);
nor U19496 (N_19496,N_17188,N_16472);
and U19497 (N_19497,N_17399,N_17033);
or U19498 (N_19498,N_16659,N_17086);
xor U19499 (N_19499,N_17181,N_16154);
nor U19500 (N_19500,N_17515,N_17540);
and U19501 (N_19501,N_17215,N_17192);
nor U19502 (N_19502,N_17980,N_16530);
nor U19503 (N_19503,N_16822,N_16343);
nor U19504 (N_19504,N_16486,N_17721);
nand U19505 (N_19505,N_17761,N_16204);
nor U19506 (N_19506,N_17114,N_17815);
nor U19507 (N_19507,N_16468,N_16379);
nand U19508 (N_19508,N_16976,N_17660);
nor U19509 (N_19509,N_16007,N_16031);
xnor U19510 (N_19510,N_16326,N_17080);
nor U19511 (N_19511,N_16430,N_16942);
xor U19512 (N_19512,N_16250,N_17689);
nor U19513 (N_19513,N_16118,N_16133);
nand U19514 (N_19514,N_17953,N_16100);
nor U19515 (N_19515,N_16833,N_16545);
nand U19516 (N_19516,N_17526,N_16708);
and U19517 (N_19517,N_16540,N_17468);
nand U19518 (N_19518,N_17192,N_17292);
or U19519 (N_19519,N_17574,N_16709);
nor U19520 (N_19520,N_17522,N_17198);
and U19521 (N_19521,N_16684,N_17651);
or U19522 (N_19522,N_16887,N_17622);
and U19523 (N_19523,N_16413,N_16333);
or U19524 (N_19524,N_16827,N_17641);
xor U19525 (N_19525,N_17491,N_17303);
and U19526 (N_19526,N_17760,N_16095);
and U19527 (N_19527,N_17342,N_16352);
nor U19528 (N_19528,N_16350,N_16523);
nor U19529 (N_19529,N_17285,N_16856);
and U19530 (N_19530,N_17280,N_17534);
nor U19531 (N_19531,N_17411,N_16197);
and U19532 (N_19532,N_16125,N_16943);
and U19533 (N_19533,N_16294,N_17371);
or U19534 (N_19534,N_17331,N_16890);
or U19535 (N_19535,N_16023,N_17433);
and U19536 (N_19536,N_16069,N_16722);
nand U19537 (N_19537,N_17329,N_17602);
or U19538 (N_19538,N_17414,N_16366);
or U19539 (N_19539,N_17043,N_16246);
xor U19540 (N_19540,N_16481,N_16422);
and U19541 (N_19541,N_17634,N_17085);
nor U19542 (N_19542,N_16281,N_16988);
and U19543 (N_19543,N_17339,N_16807);
xnor U19544 (N_19544,N_17607,N_16968);
xnor U19545 (N_19545,N_16864,N_17630);
nor U19546 (N_19546,N_17462,N_17042);
xnor U19547 (N_19547,N_17276,N_16789);
or U19548 (N_19548,N_17238,N_16981);
nor U19549 (N_19549,N_17839,N_16788);
nand U19550 (N_19550,N_17816,N_16845);
nand U19551 (N_19551,N_17339,N_17253);
nor U19552 (N_19552,N_17733,N_17341);
or U19553 (N_19553,N_16615,N_16155);
nand U19554 (N_19554,N_17275,N_16323);
nand U19555 (N_19555,N_16438,N_16704);
nand U19556 (N_19556,N_16738,N_17173);
nand U19557 (N_19557,N_17143,N_16957);
nand U19558 (N_19558,N_17154,N_16974);
or U19559 (N_19559,N_16069,N_17727);
nor U19560 (N_19560,N_16732,N_16660);
nand U19561 (N_19561,N_17160,N_17006);
nand U19562 (N_19562,N_16139,N_16808);
and U19563 (N_19563,N_17178,N_17769);
nand U19564 (N_19564,N_17857,N_16641);
nand U19565 (N_19565,N_16185,N_16833);
nor U19566 (N_19566,N_16344,N_17673);
and U19567 (N_19567,N_16668,N_17567);
or U19568 (N_19568,N_16712,N_16083);
and U19569 (N_19569,N_16386,N_16315);
nand U19570 (N_19570,N_17554,N_17664);
and U19571 (N_19571,N_17379,N_16424);
xor U19572 (N_19572,N_16798,N_17252);
nor U19573 (N_19573,N_17984,N_16227);
nor U19574 (N_19574,N_16508,N_17567);
nand U19575 (N_19575,N_16810,N_16994);
and U19576 (N_19576,N_16337,N_16162);
and U19577 (N_19577,N_16771,N_17749);
and U19578 (N_19578,N_17017,N_17112);
xor U19579 (N_19579,N_16934,N_16588);
nor U19580 (N_19580,N_17756,N_17697);
xor U19581 (N_19581,N_17413,N_17180);
nor U19582 (N_19582,N_16208,N_17910);
xnor U19583 (N_19583,N_17587,N_17793);
or U19584 (N_19584,N_16453,N_16246);
or U19585 (N_19585,N_16633,N_17757);
or U19586 (N_19586,N_16668,N_16388);
xnor U19587 (N_19587,N_16324,N_17358);
and U19588 (N_19588,N_17304,N_17506);
or U19589 (N_19589,N_16077,N_17642);
and U19590 (N_19590,N_16588,N_16066);
nand U19591 (N_19591,N_16051,N_17230);
nor U19592 (N_19592,N_17427,N_16085);
nand U19593 (N_19593,N_17434,N_17070);
or U19594 (N_19594,N_16930,N_16520);
and U19595 (N_19595,N_16489,N_16443);
nor U19596 (N_19596,N_16777,N_17332);
nor U19597 (N_19597,N_17844,N_16549);
nand U19598 (N_19598,N_17055,N_17669);
and U19599 (N_19599,N_17739,N_16304);
and U19600 (N_19600,N_16891,N_16026);
or U19601 (N_19601,N_17785,N_17994);
or U19602 (N_19602,N_17902,N_17630);
nor U19603 (N_19603,N_17668,N_16288);
nand U19604 (N_19604,N_16113,N_17695);
nand U19605 (N_19605,N_16997,N_16381);
or U19606 (N_19606,N_16184,N_17090);
xnor U19607 (N_19607,N_17312,N_17959);
xor U19608 (N_19608,N_16199,N_17839);
and U19609 (N_19609,N_16910,N_16335);
and U19610 (N_19610,N_17083,N_17639);
nor U19611 (N_19611,N_16841,N_17988);
nand U19612 (N_19612,N_17633,N_17468);
xor U19613 (N_19613,N_17207,N_17959);
nor U19614 (N_19614,N_17671,N_17942);
xnor U19615 (N_19615,N_16248,N_16356);
or U19616 (N_19616,N_17821,N_17752);
and U19617 (N_19617,N_16779,N_17202);
xor U19618 (N_19618,N_17735,N_17893);
or U19619 (N_19619,N_17175,N_17842);
nor U19620 (N_19620,N_16987,N_16807);
and U19621 (N_19621,N_17861,N_16108);
nor U19622 (N_19622,N_16959,N_17686);
nand U19623 (N_19623,N_16952,N_16878);
or U19624 (N_19624,N_17901,N_17877);
nor U19625 (N_19625,N_17182,N_17947);
nor U19626 (N_19626,N_17270,N_16194);
nand U19627 (N_19627,N_16206,N_17292);
nor U19628 (N_19628,N_17262,N_16492);
or U19629 (N_19629,N_16513,N_16144);
or U19630 (N_19630,N_17387,N_17103);
nor U19631 (N_19631,N_17190,N_17442);
nand U19632 (N_19632,N_17398,N_16718);
xor U19633 (N_19633,N_17691,N_17896);
xnor U19634 (N_19634,N_17700,N_17392);
or U19635 (N_19635,N_17724,N_17018);
and U19636 (N_19636,N_17498,N_16520);
or U19637 (N_19637,N_16736,N_16845);
and U19638 (N_19638,N_17345,N_16793);
or U19639 (N_19639,N_17684,N_17766);
nor U19640 (N_19640,N_17278,N_16822);
or U19641 (N_19641,N_17266,N_16087);
xnor U19642 (N_19642,N_17192,N_17173);
nand U19643 (N_19643,N_17110,N_17750);
and U19644 (N_19644,N_17266,N_16765);
nor U19645 (N_19645,N_16530,N_17868);
or U19646 (N_19646,N_16477,N_16178);
or U19647 (N_19647,N_16053,N_16423);
nand U19648 (N_19648,N_17405,N_16402);
or U19649 (N_19649,N_16679,N_16224);
nor U19650 (N_19650,N_16350,N_17819);
nand U19651 (N_19651,N_17514,N_16185);
or U19652 (N_19652,N_17739,N_16156);
xor U19653 (N_19653,N_16710,N_16849);
nand U19654 (N_19654,N_17989,N_17382);
nor U19655 (N_19655,N_16881,N_16635);
nor U19656 (N_19656,N_17115,N_16649);
nand U19657 (N_19657,N_16838,N_16415);
nor U19658 (N_19658,N_17103,N_16045);
or U19659 (N_19659,N_17654,N_17030);
or U19660 (N_19660,N_16502,N_17545);
xnor U19661 (N_19661,N_17145,N_16792);
or U19662 (N_19662,N_17388,N_16045);
xnor U19663 (N_19663,N_17009,N_17803);
nor U19664 (N_19664,N_17503,N_16487);
or U19665 (N_19665,N_17366,N_17277);
nor U19666 (N_19666,N_17981,N_17739);
and U19667 (N_19667,N_17211,N_17462);
nor U19668 (N_19668,N_16829,N_17804);
xor U19669 (N_19669,N_17088,N_17363);
nor U19670 (N_19670,N_16915,N_17643);
nand U19671 (N_19671,N_17623,N_16894);
nor U19672 (N_19672,N_17484,N_17900);
nand U19673 (N_19673,N_16124,N_16348);
nor U19674 (N_19674,N_17324,N_16248);
or U19675 (N_19675,N_16259,N_17872);
or U19676 (N_19676,N_16245,N_17570);
xnor U19677 (N_19677,N_16363,N_16154);
and U19678 (N_19678,N_16776,N_17777);
nor U19679 (N_19679,N_16238,N_17633);
and U19680 (N_19680,N_16241,N_17149);
and U19681 (N_19681,N_16271,N_17486);
and U19682 (N_19682,N_16643,N_17367);
or U19683 (N_19683,N_16928,N_17079);
or U19684 (N_19684,N_17844,N_17005);
or U19685 (N_19685,N_16519,N_17895);
nor U19686 (N_19686,N_17814,N_16732);
nand U19687 (N_19687,N_16897,N_17524);
and U19688 (N_19688,N_16824,N_16535);
nand U19689 (N_19689,N_17443,N_16512);
nor U19690 (N_19690,N_16722,N_16786);
xor U19691 (N_19691,N_16974,N_16252);
and U19692 (N_19692,N_16842,N_16313);
nand U19693 (N_19693,N_16588,N_17833);
xnor U19694 (N_19694,N_16222,N_17207);
nor U19695 (N_19695,N_17947,N_17790);
and U19696 (N_19696,N_16928,N_16627);
or U19697 (N_19697,N_16916,N_17415);
or U19698 (N_19698,N_16391,N_16761);
and U19699 (N_19699,N_17870,N_16830);
or U19700 (N_19700,N_16662,N_17601);
or U19701 (N_19701,N_17235,N_16543);
xor U19702 (N_19702,N_16898,N_16136);
and U19703 (N_19703,N_16601,N_17329);
nand U19704 (N_19704,N_17406,N_16043);
nor U19705 (N_19705,N_16988,N_16889);
or U19706 (N_19706,N_16666,N_16167);
or U19707 (N_19707,N_17752,N_16788);
nor U19708 (N_19708,N_16954,N_17200);
nand U19709 (N_19709,N_16774,N_16355);
or U19710 (N_19710,N_17389,N_17044);
or U19711 (N_19711,N_16354,N_17404);
xor U19712 (N_19712,N_17235,N_16452);
xnor U19713 (N_19713,N_16772,N_17248);
nor U19714 (N_19714,N_17865,N_17089);
or U19715 (N_19715,N_16983,N_17573);
and U19716 (N_19716,N_16081,N_16292);
or U19717 (N_19717,N_17311,N_17879);
or U19718 (N_19718,N_16663,N_16589);
and U19719 (N_19719,N_17027,N_17140);
xor U19720 (N_19720,N_16383,N_17053);
nand U19721 (N_19721,N_17730,N_17986);
or U19722 (N_19722,N_16330,N_17133);
or U19723 (N_19723,N_16498,N_17630);
or U19724 (N_19724,N_17461,N_17832);
and U19725 (N_19725,N_17102,N_17294);
nor U19726 (N_19726,N_17481,N_17511);
nand U19727 (N_19727,N_17529,N_16966);
xnor U19728 (N_19728,N_17477,N_17853);
xor U19729 (N_19729,N_17290,N_17935);
nor U19730 (N_19730,N_17047,N_17543);
and U19731 (N_19731,N_17551,N_17400);
nor U19732 (N_19732,N_16189,N_16978);
or U19733 (N_19733,N_16311,N_17864);
nand U19734 (N_19734,N_16576,N_16887);
nand U19735 (N_19735,N_17346,N_16250);
nand U19736 (N_19736,N_16540,N_16397);
nand U19737 (N_19737,N_16170,N_16479);
nand U19738 (N_19738,N_17832,N_16118);
or U19739 (N_19739,N_17731,N_16857);
nand U19740 (N_19740,N_17459,N_16174);
nor U19741 (N_19741,N_17163,N_16632);
and U19742 (N_19742,N_16568,N_17259);
or U19743 (N_19743,N_16333,N_16679);
and U19744 (N_19744,N_17843,N_16554);
and U19745 (N_19745,N_16340,N_16381);
or U19746 (N_19746,N_17515,N_17433);
nand U19747 (N_19747,N_17542,N_16037);
or U19748 (N_19748,N_17179,N_16953);
or U19749 (N_19749,N_16750,N_16135);
nor U19750 (N_19750,N_17134,N_16767);
xnor U19751 (N_19751,N_17080,N_16162);
xor U19752 (N_19752,N_17429,N_16947);
or U19753 (N_19753,N_17462,N_17884);
nand U19754 (N_19754,N_16088,N_17319);
nand U19755 (N_19755,N_16537,N_16971);
nor U19756 (N_19756,N_16881,N_17949);
nand U19757 (N_19757,N_16252,N_17909);
or U19758 (N_19758,N_17427,N_16627);
and U19759 (N_19759,N_16748,N_16858);
nand U19760 (N_19760,N_17839,N_16961);
xor U19761 (N_19761,N_16858,N_16448);
nand U19762 (N_19762,N_17196,N_16629);
nor U19763 (N_19763,N_16543,N_17394);
nand U19764 (N_19764,N_16406,N_16506);
nor U19765 (N_19765,N_17004,N_16165);
nand U19766 (N_19766,N_16320,N_17469);
nor U19767 (N_19767,N_16154,N_16866);
nor U19768 (N_19768,N_16561,N_16393);
nor U19769 (N_19769,N_17099,N_17058);
and U19770 (N_19770,N_16129,N_17576);
and U19771 (N_19771,N_17178,N_16353);
and U19772 (N_19772,N_17347,N_17397);
nor U19773 (N_19773,N_16768,N_16544);
or U19774 (N_19774,N_16417,N_17899);
or U19775 (N_19775,N_17174,N_17816);
xor U19776 (N_19776,N_16489,N_16299);
and U19777 (N_19777,N_16067,N_16983);
nand U19778 (N_19778,N_16879,N_16972);
and U19779 (N_19779,N_17180,N_16999);
xnor U19780 (N_19780,N_16812,N_17985);
nand U19781 (N_19781,N_17531,N_17438);
nor U19782 (N_19782,N_16547,N_17001);
xor U19783 (N_19783,N_17594,N_17347);
and U19784 (N_19784,N_17864,N_17992);
nand U19785 (N_19785,N_17651,N_16790);
nand U19786 (N_19786,N_17159,N_17837);
and U19787 (N_19787,N_16213,N_17290);
and U19788 (N_19788,N_16349,N_16143);
and U19789 (N_19789,N_16231,N_16813);
nor U19790 (N_19790,N_16943,N_17231);
or U19791 (N_19791,N_16959,N_17566);
nor U19792 (N_19792,N_16846,N_17813);
or U19793 (N_19793,N_17680,N_17282);
nand U19794 (N_19794,N_16205,N_17085);
xor U19795 (N_19795,N_16082,N_17686);
or U19796 (N_19796,N_16915,N_16081);
nor U19797 (N_19797,N_17127,N_17952);
nand U19798 (N_19798,N_16954,N_16020);
xnor U19799 (N_19799,N_17379,N_16893);
xor U19800 (N_19800,N_17916,N_17362);
nand U19801 (N_19801,N_16914,N_16868);
xor U19802 (N_19802,N_17174,N_16737);
nand U19803 (N_19803,N_17513,N_16663);
nor U19804 (N_19804,N_17987,N_16643);
and U19805 (N_19805,N_17848,N_16963);
xnor U19806 (N_19806,N_16404,N_16543);
nor U19807 (N_19807,N_17494,N_16376);
xnor U19808 (N_19808,N_17478,N_16907);
nor U19809 (N_19809,N_16940,N_16279);
nor U19810 (N_19810,N_16468,N_17149);
xnor U19811 (N_19811,N_16559,N_16640);
and U19812 (N_19812,N_16540,N_16944);
and U19813 (N_19813,N_16220,N_16989);
xor U19814 (N_19814,N_16676,N_17289);
and U19815 (N_19815,N_17592,N_16342);
and U19816 (N_19816,N_16296,N_17396);
nor U19817 (N_19817,N_16420,N_17745);
nand U19818 (N_19818,N_16113,N_17011);
xor U19819 (N_19819,N_16569,N_16562);
nor U19820 (N_19820,N_17968,N_16184);
nand U19821 (N_19821,N_17154,N_16202);
or U19822 (N_19822,N_17567,N_17690);
or U19823 (N_19823,N_17425,N_16406);
and U19824 (N_19824,N_17411,N_17540);
xnor U19825 (N_19825,N_17420,N_16301);
xnor U19826 (N_19826,N_17052,N_16644);
or U19827 (N_19827,N_17307,N_17465);
nand U19828 (N_19828,N_16833,N_16419);
nand U19829 (N_19829,N_17336,N_17798);
xnor U19830 (N_19830,N_17342,N_17732);
nand U19831 (N_19831,N_17845,N_17994);
or U19832 (N_19832,N_16783,N_16912);
or U19833 (N_19833,N_17191,N_16871);
and U19834 (N_19834,N_17554,N_17778);
and U19835 (N_19835,N_17815,N_16527);
and U19836 (N_19836,N_16290,N_17685);
nor U19837 (N_19837,N_16719,N_17140);
and U19838 (N_19838,N_16434,N_17471);
or U19839 (N_19839,N_17623,N_17020);
xor U19840 (N_19840,N_17231,N_17879);
xor U19841 (N_19841,N_17222,N_16633);
or U19842 (N_19842,N_17922,N_16077);
or U19843 (N_19843,N_16249,N_16923);
or U19844 (N_19844,N_16258,N_16757);
xnor U19845 (N_19845,N_17240,N_16578);
or U19846 (N_19846,N_17930,N_16106);
and U19847 (N_19847,N_17998,N_16984);
and U19848 (N_19848,N_17765,N_16269);
nand U19849 (N_19849,N_16950,N_16844);
nand U19850 (N_19850,N_16389,N_16723);
or U19851 (N_19851,N_16778,N_17325);
or U19852 (N_19852,N_17509,N_16891);
and U19853 (N_19853,N_17634,N_16715);
and U19854 (N_19854,N_16971,N_17324);
nand U19855 (N_19855,N_17342,N_17288);
and U19856 (N_19856,N_16478,N_17573);
xor U19857 (N_19857,N_17546,N_17479);
and U19858 (N_19858,N_17560,N_17697);
or U19859 (N_19859,N_16334,N_16932);
nor U19860 (N_19860,N_17633,N_16302);
nor U19861 (N_19861,N_17903,N_17181);
xor U19862 (N_19862,N_17649,N_16193);
nor U19863 (N_19863,N_16523,N_16023);
and U19864 (N_19864,N_16474,N_17944);
or U19865 (N_19865,N_17367,N_17992);
or U19866 (N_19866,N_16072,N_17691);
nand U19867 (N_19867,N_16607,N_17713);
nand U19868 (N_19868,N_17215,N_16557);
xor U19869 (N_19869,N_17583,N_16447);
nand U19870 (N_19870,N_16974,N_17096);
or U19871 (N_19871,N_17366,N_17251);
and U19872 (N_19872,N_17192,N_16129);
and U19873 (N_19873,N_16710,N_16756);
nand U19874 (N_19874,N_17589,N_17756);
or U19875 (N_19875,N_16229,N_16432);
nor U19876 (N_19876,N_16624,N_16501);
and U19877 (N_19877,N_17529,N_17497);
xor U19878 (N_19878,N_17112,N_16822);
nor U19879 (N_19879,N_16106,N_16740);
or U19880 (N_19880,N_17696,N_16821);
nor U19881 (N_19881,N_17576,N_17509);
or U19882 (N_19882,N_16016,N_16108);
and U19883 (N_19883,N_16926,N_16021);
and U19884 (N_19884,N_16012,N_17258);
or U19885 (N_19885,N_17627,N_17274);
or U19886 (N_19886,N_16704,N_17218);
and U19887 (N_19887,N_17288,N_17857);
nand U19888 (N_19888,N_17266,N_17633);
or U19889 (N_19889,N_16288,N_17583);
nand U19890 (N_19890,N_17354,N_16183);
xnor U19891 (N_19891,N_17117,N_17994);
nor U19892 (N_19892,N_17977,N_16610);
or U19893 (N_19893,N_17269,N_16786);
or U19894 (N_19894,N_17805,N_17847);
nand U19895 (N_19895,N_17493,N_16831);
and U19896 (N_19896,N_16987,N_16097);
and U19897 (N_19897,N_16900,N_16769);
xor U19898 (N_19898,N_17101,N_16429);
and U19899 (N_19899,N_17813,N_17090);
nand U19900 (N_19900,N_17920,N_17836);
and U19901 (N_19901,N_17263,N_17754);
xnor U19902 (N_19902,N_16044,N_16720);
or U19903 (N_19903,N_16531,N_17576);
nor U19904 (N_19904,N_17853,N_16013);
xor U19905 (N_19905,N_16642,N_16382);
xnor U19906 (N_19906,N_16025,N_17752);
nand U19907 (N_19907,N_16649,N_16246);
nor U19908 (N_19908,N_16989,N_17777);
nand U19909 (N_19909,N_17236,N_16176);
xnor U19910 (N_19910,N_17335,N_17719);
xnor U19911 (N_19911,N_16133,N_16352);
nor U19912 (N_19912,N_16371,N_16886);
xor U19913 (N_19913,N_16273,N_16706);
and U19914 (N_19914,N_17325,N_17249);
nor U19915 (N_19915,N_16801,N_17073);
or U19916 (N_19916,N_16531,N_16810);
nand U19917 (N_19917,N_16155,N_17532);
nor U19918 (N_19918,N_16875,N_17721);
or U19919 (N_19919,N_16485,N_16037);
nor U19920 (N_19920,N_16779,N_17923);
nor U19921 (N_19921,N_17599,N_16511);
xor U19922 (N_19922,N_17790,N_16906);
nand U19923 (N_19923,N_16544,N_16829);
nor U19924 (N_19924,N_16338,N_16762);
nand U19925 (N_19925,N_16317,N_17113);
xor U19926 (N_19926,N_16854,N_17102);
nand U19927 (N_19927,N_16269,N_16199);
xnor U19928 (N_19928,N_16240,N_17228);
nor U19929 (N_19929,N_17779,N_17673);
or U19930 (N_19930,N_16877,N_16418);
xor U19931 (N_19931,N_16506,N_17642);
nor U19932 (N_19932,N_17306,N_17120);
nand U19933 (N_19933,N_16357,N_17594);
nand U19934 (N_19934,N_16451,N_17595);
or U19935 (N_19935,N_16766,N_17415);
or U19936 (N_19936,N_16510,N_16128);
nand U19937 (N_19937,N_17957,N_17582);
nor U19938 (N_19938,N_16972,N_17134);
nand U19939 (N_19939,N_17434,N_16632);
nor U19940 (N_19940,N_16616,N_17725);
nor U19941 (N_19941,N_17383,N_17823);
and U19942 (N_19942,N_16109,N_16725);
and U19943 (N_19943,N_17065,N_17959);
xor U19944 (N_19944,N_16301,N_16913);
and U19945 (N_19945,N_16297,N_17942);
and U19946 (N_19946,N_17650,N_16372);
or U19947 (N_19947,N_17337,N_17258);
xnor U19948 (N_19948,N_17563,N_16398);
nor U19949 (N_19949,N_17060,N_17433);
or U19950 (N_19950,N_17000,N_17757);
nand U19951 (N_19951,N_17904,N_17186);
and U19952 (N_19952,N_17692,N_16050);
xnor U19953 (N_19953,N_16784,N_17848);
xor U19954 (N_19954,N_16745,N_16325);
nand U19955 (N_19955,N_16129,N_16546);
nand U19956 (N_19956,N_17253,N_17755);
nand U19957 (N_19957,N_17475,N_17477);
nand U19958 (N_19958,N_16717,N_17144);
xor U19959 (N_19959,N_16517,N_16816);
and U19960 (N_19960,N_17064,N_17488);
nor U19961 (N_19961,N_16010,N_17036);
nor U19962 (N_19962,N_17776,N_16767);
nor U19963 (N_19963,N_17961,N_16341);
nand U19964 (N_19964,N_17985,N_16333);
and U19965 (N_19965,N_17121,N_17957);
and U19966 (N_19966,N_16127,N_16380);
nor U19967 (N_19967,N_16407,N_17133);
nand U19968 (N_19968,N_16017,N_16156);
or U19969 (N_19969,N_16401,N_17539);
or U19970 (N_19970,N_16249,N_17358);
nor U19971 (N_19971,N_17457,N_17788);
xor U19972 (N_19972,N_17364,N_16394);
and U19973 (N_19973,N_16066,N_16842);
nand U19974 (N_19974,N_16185,N_17406);
nor U19975 (N_19975,N_17859,N_17688);
nor U19976 (N_19976,N_16691,N_16562);
or U19977 (N_19977,N_16546,N_17872);
nor U19978 (N_19978,N_17692,N_16846);
or U19979 (N_19979,N_16828,N_17365);
and U19980 (N_19980,N_16641,N_16507);
nand U19981 (N_19981,N_17217,N_16411);
nor U19982 (N_19982,N_17767,N_17700);
nand U19983 (N_19983,N_16648,N_17148);
or U19984 (N_19984,N_16834,N_16441);
nor U19985 (N_19985,N_17199,N_17780);
nand U19986 (N_19986,N_17683,N_16667);
nand U19987 (N_19987,N_17267,N_17814);
nor U19988 (N_19988,N_17437,N_17130);
and U19989 (N_19989,N_16174,N_17224);
xnor U19990 (N_19990,N_16653,N_17613);
nand U19991 (N_19991,N_17965,N_17903);
nand U19992 (N_19992,N_17225,N_16812);
xnor U19993 (N_19993,N_17315,N_16658);
or U19994 (N_19994,N_17495,N_16280);
nor U19995 (N_19995,N_16550,N_17365);
nor U19996 (N_19996,N_17965,N_17565);
or U19997 (N_19997,N_16090,N_17337);
or U19998 (N_19998,N_16916,N_17943);
and U19999 (N_19999,N_17278,N_16699);
nor UO_0 (O_0,N_19020,N_18726);
nand UO_1 (O_1,N_19422,N_19247);
or UO_2 (O_2,N_18031,N_18837);
xnor UO_3 (O_3,N_18488,N_18101);
xnor UO_4 (O_4,N_19197,N_18772);
or UO_5 (O_5,N_18591,N_18251);
or UO_6 (O_6,N_18344,N_18906);
nor UO_7 (O_7,N_19368,N_19217);
and UO_8 (O_8,N_18197,N_19405);
xor UO_9 (O_9,N_18621,N_18858);
and UO_10 (O_10,N_19187,N_18176);
nor UO_11 (O_11,N_18040,N_19813);
xnor UO_12 (O_12,N_19407,N_19530);
nor UO_13 (O_13,N_18080,N_18972);
nor UO_14 (O_14,N_19550,N_19935);
and UO_15 (O_15,N_18536,N_19005);
nor UO_16 (O_16,N_19641,N_18196);
nor UO_17 (O_17,N_19842,N_18616);
nor UO_18 (O_18,N_19671,N_19763);
nor UO_19 (O_19,N_18375,N_18423);
or UO_20 (O_20,N_19387,N_18125);
xor UO_21 (O_21,N_19992,N_19988);
xnor UO_22 (O_22,N_19209,N_19078);
and UO_23 (O_23,N_19539,N_18180);
xor UO_24 (O_24,N_19127,N_19555);
nand UO_25 (O_25,N_19939,N_19196);
nor UO_26 (O_26,N_19699,N_18129);
and UO_27 (O_27,N_19288,N_18099);
nor UO_28 (O_28,N_18645,N_18851);
nand UO_29 (O_29,N_18059,N_18317);
nand UO_30 (O_30,N_18421,N_18308);
xor UO_31 (O_31,N_18511,N_19451);
nor UO_32 (O_32,N_19309,N_18753);
xor UO_33 (O_33,N_19305,N_19681);
and UO_34 (O_34,N_19154,N_19929);
and UO_35 (O_35,N_18786,N_18212);
xor UO_36 (O_36,N_19706,N_18428);
or UO_37 (O_37,N_19902,N_19468);
or UO_38 (O_38,N_18350,N_19470);
xor UO_39 (O_39,N_19836,N_18311);
or UO_40 (O_40,N_18980,N_18143);
or UO_41 (O_41,N_18495,N_19337);
or UO_42 (O_42,N_19622,N_18496);
or UO_43 (O_43,N_18225,N_19852);
or UO_44 (O_44,N_19172,N_19045);
and UO_45 (O_45,N_18050,N_18657);
or UO_46 (O_46,N_19609,N_18363);
and UO_47 (O_47,N_19921,N_18992);
nand UO_48 (O_48,N_19439,N_19116);
and UO_49 (O_49,N_19794,N_19535);
xor UO_50 (O_50,N_18452,N_18364);
nand UO_51 (O_51,N_19199,N_19185);
nand UO_52 (O_52,N_19460,N_18727);
or UO_53 (O_53,N_19801,N_19653);
nor UO_54 (O_54,N_19354,N_18867);
and UO_55 (O_55,N_19677,N_19096);
xor UO_56 (O_56,N_18417,N_18009);
and UO_57 (O_57,N_19322,N_19263);
nor UO_58 (O_58,N_19300,N_19252);
and UO_59 (O_59,N_19219,N_18969);
and UO_60 (O_60,N_19245,N_18401);
xnor UO_61 (O_61,N_18512,N_18324);
or UO_62 (O_62,N_18289,N_19048);
or UO_63 (O_63,N_19459,N_18169);
xor UO_64 (O_64,N_19546,N_19548);
xnor UO_65 (O_65,N_18988,N_18817);
nor UO_66 (O_66,N_18655,N_19869);
nand UO_67 (O_67,N_18260,N_19983);
nand UO_68 (O_68,N_19824,N_19807);
nand UO_69 (O_69,N_18694,N_19499);
nand UO_70 (O_70,N_18541,N_19188);
or UO_71 (O_71,N_18204,N_19142);
nor UO_72 (O_72,N_18083,N_18704);
or UO_73 (O_73,N_19965,N_19120);
and UO_74 (O_74,N_19849,N_18661);
or UO_75 (O_75,N_18079,N_19355);
nor UO_76 (O_76,N_19634,N_19118);
and UO_77 (O_77,N_19229,N_19558);
or UO_78 (O_78,N_19596,N_18662);
or UO_79 (O_79,N_19950,N_18192);
nand UO_80 (O_80,N_19338,N_19254);
xor UO_81 (O_81,N_18893,N_19086);
nor UO_82 (O_82,N_18041,N_19533);
xnor UO_83 (O_83,N_18241,N_19186);
or UO_84 (O_84,N_19620,N_18530);
or UO_85 (O_85,N_18901,N_19746);
nand UO_86 (O_86,N_19532,N_18303);
nand UO_87 (O_87,N_19287,N_19081);
nand UO_88 (O_88,N_19053,N_18049);
and UO_89 (O_89,N_18022,N_18320);
xnor UO_90 (O_90,N_18791,N_18834);
or UO_91 (O_91,N_19203,N_18957);
xor UO_92 (O_92,N_19388,N_19315);
and UO_93 (O_93,N_18414,N_18798);
or UO_94 (O_94,N_19421,N_19665);
or UO_95 (O_95,N_19833,N_18730);
and UO_96 (O_96,N_19614,N_18577);
and UO_97 (O_97,N_19011,N_18744);
nand UO_98 (O_98,N_18675,N_19115);
nand UO_99 (O_99,N_19456,N_18234);
nand UO_100 (O_100,N_19313,N_18047);
or UO_101 (O_101,N_19095,N_18356);
xor UO_102 (O_102,N_18956,N_18250);
or UO_103 (O_103,N_19790,N_19717);
and UO_104 (O_104,N_19832,N_18390);
xor UO_105 (O_105,N_18658,N_19625);
xnor UO_106 (O_106,N_18590,N_18546);
nand UO_107 (O_107,N_19751,N_19231);
or UO_108 (O_108,N_19168,N_18291);
nand UO_109 (O_109,N_18127,N_18701);
nor UO_110 (O_110,N_18416,N_19789);
nand UO_111 (O_111,N_19701,N_19960);
nor UO_112 (O_112,N_18751,N_19381);
nand UO_113 (O_113,N_18776,N_18869);
nand UO_114 (O_114,N_19099,N_19075);
xnor UO_115 (O_115,N_19289,N_18014);
nor UO_116 (O_116,N_19870,N_18315);
or UO_117 (O_117,N_18912,N_18134);
and UO_118 (O_118,N_19759,N_19526);
and UO_119 (O_119,N_19705,N_19332);
or UO_120 (O_120,N_19258,N_19396);
nand UO_121 (O_121,N_18908,N_19403);
nand UO_122 (O_122,N_19781,N_19292);
or UO_123 (O_123,N_19787,N_18807);
and UO_124 (O_124,N_19382,N_19108);
xnor UO_125 (O_125,N_19176,N_18497);
xnor UO_126 (O_126,N_19017,N_18777);
and UO_127 (O_127,N_18220,N_18809);
nor UO_128 (O_128,N_18270,N_18264);
or UO_129 (O_129,N_19624,N_18028);
nand UO_130 (O_130,N_19933,N_18240);
xor UO_131 (O_131,N_18248,N_18115);
nand UO_132 (O_132,N_18432,N_19452);
or UO_133 (O_133,N_19371,N_18567);
and UO_134 (O_134,N_19386,N_18671);
and UO_135 (O_135,N_18935,N_19628);
and UO_136 (O_136,N_19964,N_18709);
and UO_137 (O_137,N_19588,N_18319);
or UO_138 (O_138,N_19385,N_18337);
xnor UO_139 (O_139,N_18140,N_19942);
or UO_140 (O_140,N_19238,N_18411);
or UO_141 (O_141,N_18454,N_18610);
nand UO_142 (O_142,N_19586,N_18903);
nor UO_143 (O_143,N_19205,N_19006);
xnor UO_144 (O_144,N_19718,N_19672);
nor UO_145 (O_145,N_19283,N_18941);
or UO_146 (O_146,N_19331,N_18019);
nand UO_147 (O_147,N_18642,N_18879);
nand UO_148 (O_148,N_19366,N_19211);
or UO_149 (O_149,N_19136,N_18237);
or UO_150 (O_150,N_19675,N_18024);
nand UO_151 (O_151,N_18729,N_18557);
or UO_152 (O_152,N_19919,N_18669);
xor UO_153 (O_153,N_18659,N_19682);
xor UO_154 (O_154,N_19685,N_19952);
or UO_155 (O_155,N_19028,N_19777);
nand UO_156 (O_156,N_19733,N_18529);
nor UO_157 (O_157,N_18789,N_19834);
nand UO_158 (O_158,N_18396,N_18293);
xnor UO_159 (O_159,N_18299,N_18412);
nor UO_160 (O_160,N_18921,N_18975);
nor UO_161 (O_161,N_18819,N_19246);
nor UO_162 (O_162,N_19450,N_18711);
xnor UO_163 (O_163,N_19339,N_19150);
nor UO_164 (O_164,N_19394,N_19074);
nand UO_165 (O_165,N_19798,N_19893);
xor UO_166 (O_166,N_19092,N_19156);
xnor UO_167 (O_167,N_19709,N_18145);
nand UO_168 (O_168,N_18932,N_18164);
nand UO_169 (O_169,N_18058,N_19696);
and UO_170 (O_170,N_18934,N_19866);
nor UO_171 (O_171,N_18501,N_19481);
or UO_172 (O_172,N_18021,N_19666);
and UO_173 (O_173,N_19523,N_19037);
or UO_174 (O_174,N_19103,N_18314);
and UO_175 (O_175,N_18780,N_19559);
and UO_176 (O_176,N_19910,N_19743);
nand UO_177 (O_177,N_18369,N_18861);
xnor UO_178 (O_178,N_19494,N_19419);
and UO_179 (O_179,N_19298,N_19432);
xor UO_180 (O_180,N_19811,N_19365);
nand UO_181 (O_181,N_18628,N_18153);
and UO_182 (O_182,N_19930,N_18779);
xnor UO_183 (O_183,N_18526,N_18468);
nand UO_184 (O_184,N_19629,N_19433);
and UO_185 (O_185,N_19577,N_19537);
nor UO_186 (O_186,N_19175,N_18632);
or UO_187 (O_187,N_19390,N_18995);
and UO_188 (O_188,N_18110,N_18137);
or UO_189 (O_189,N_18576,N_18760);
and UO_190 (O_190,N_19969,N_19324);
or UO_191 (O_191,N_18651,N_19585);
and UO_192 (O_192,N_18706,N_18967);
and UO_193 (O_193,N_18409,N_19241);
nand UO_194 (O_194,N_19391,N_19441);
nand UO_195 (O_195,N_18207,N_18046);
xnor UO_196 (O_196,N_19151,N_19016);
xor UO_197 (O_197,N_18962,N_18702);
xnor UO_198 (O_198,N_19655,N_18441);
and UO_199 (O_199,N_18533,N_19650);
nor UO_200 (O_200,N_19761,N_19589);
or UO_201 (O_201,N_19525,N_19491);
or UO_202 (O_202,N_19991,N_19265);
xnor UO_203 (O_203,N_19621,N_19444);
and UO_204 (O_204,N_18928,N_19707);
nor UO_205 (O_205,N_19540,N_19610);
or UO_206 (O_206,N_19000,N_19465);
or UO_207 (O_207,N_19236,N_19512);
xnor UO_208 (O_208,N_19141,N_18377);
and UO_209 (O_209,N_18721,N_19233);
or UO_210 (O_210,N_19818,N_18784);
nand UO_211 (O_211,N_19778,N_19956);
and UO_212 (O_212,N_19259,N_18588);
nor UO_213 (O_213,N_19959,N_19035);
nor UO_214 (O_214,N_19947,N_18647);
xnor UO_215 (O_215,N_19080,N_19941);
xnor UO_216 (O_216,N_18684,N_19731);
or UO_217 (O_217,N_19690,N_18551);
and UO_218 (O_218,N_19018,N_18355);
nor UO_219 (O_219,N_18128,N_19061);
or UO_220 (O_220,N_19106,N_19047);
or UO_221 (O_221,N_18518,N_18609);
nand UO_222 (O_222,N_18818,N_18746);
nand UO_223 (O_223,N_19090,N_18783);
xor UO_224 (O_224,N_18097,N_18348);
xor UO_225 (O_225,N_19534,N_18894);
xor UO_226 (O_226,N_18193,N_19180);
nand UO_227 (O_227,N_18177,N_18224);
xnor UO_228 (O_228,N_18810,N_19125);
nand UO_229 (O_229,N_19033,N_19311);
nor UO_230 (O_230,N_19282,N_19167);
or UO_231 (O_231,N_19580,N_18823);
and UO_232 (O_232,N_19206,N_19483);
and UO_233 (O_233,N_18071,N_18833);
and UO_234 (O_234,N_19242,N_19886);
or UO_235 (O_235,N_18318,N_19198);
and UO_236 (O_236,N_18800,N_19130);
and UO_237 (O_237,N_18082,N_18135);
xnor UO_238 (O_238,N_19587,N_19021);
nor UO_239 (O_239,N_18687,N_18279);
or UO_240 (O_240,N_19519,N_18506);
or UO_241 (O_241,N_18742,N_18309);
or UO_242 (O_242,N_19520,N_18078);
nor UO_243 (O_243,N_18829,N_19771);
and UO_244 (O_244,N_19883,N_19235);
nor UO_245 (O_245,N_19182,N_19592);
nand UO_246 (O_246,N_18924,N_18508);
and UO_247 (O_247,N_19595,N_18963);
xnor UO_248 (O_248,N_19341,N_18252);
or UO_249 (O_249,N_19788,N_19498);
xor UO_250 (O_250,N_18987,N_18007);
or UO_251 (O_251,N_19318,N_18208);
and UO_252 (O_252,N_18682,N_18882);
nand UO_253 (O_253,N_18144,N_19511);
and UO_254 (O_254,N_18563,N_19556);
xnor UO_255 (O_255,N_18615,N_18371);
nand UO_256 (O_256,N_19384,N_19213);
xor UO_257 (O_257,N_19924,N_18166);
nand UO_258 (O_258,N_19604,N_18302);
or UO_259 (O_259,N_19662,N_19361);
and UO_260 (O_260,N_18648,N_18313);
nand UO_261 (O_261,N_19104,N_18068);
nand UO_262 (O_262,N_19266,N_19899);
or UO_263 (O_263,N_18464,N_18354);
nand UO_264 (O_264,N_19170,N_19515);
nand UO_265 (O_265,N_18275,N_18516);
xnor UO_266 (O_266,N_19190,N_18267);
or UO_267 (O_267,N_19827,N_18827);
nor UO_268 (O_268,N_19776,N_18568);
nor UO_269 (O_269,N_19748,N_18262);
or UO_270 (O_270,N_18604,N_18623);
xor UO_271 (O_271,N_18334,N_18582);
and UO_272 (O_272,N_18538,N_19109);
and UO_273 (O_273,N_18971,N_19750);
and UO_274 (O_274,N_18718,N_19226);
nor UO_275 (O_275,N_18639,N_19200);
and UO_276 (O_276,N_18277,N_18855);
nor UO_277 (O_277,N_18612,N_18089);
and UO_278 (O_278,N_19193,N_19766);
xor UO_279 (O_279,N_18030,N_18304);
and UO_280 (O_280,N_18806,N_18206);
nor UO_281 (O_281,N_19412,N_18649);
xor UO_282 (O_282,N_19635,N_19256);
nor UO_283 (O_283,N_19358,N_18184);
or UO_284 (O_284,N_18133,N_19431);
nor UO_285 (O_285,N_19314,N_18722);
and UO_286 (O_286,N_19907,N_18764);
xor UO_287 (O_287,N_19729,N_19100);
nand UO_288 (O_288,N_19846,N_18010);
xnor UO_289 (O_289,N_18902,N_19144);
xnor UO_290 (O_290,N_18054,N_19202);
and UO_291 (O_291,N_19274,N_19928);
nor UO_292 (O_292,N_19296,N_18449);
or UO_293 (O_293,N_19079,N_19885);
or UO_294 (O_294,N_19440,N_19476);
or UO_295 (O_295,N_18832,N_18725);
or UO_296 (O_296,N_19906,N_19216);
and UO_297 (O_297,N_19514,N_19069);
nand UO_298 (O_298,N_19521,N_19607);
or UO_299 (O_299,N_19327,N_18247);
xor UO_300 (O_300,N_19058,N_18871);
or UO_301 (O_301,N_18660,N_18710);
nand UO_302 (O_302,N_18794,N_18425);
xor UO_303 (O_303,N_18678,N_18976);
xnor UO_304 (O_304,N_18700,N_19303);
xnor UO_305 (O_305,N_18084,N_18636);
nand UO_306 (O_306,N_18094,N_18802);
nor UO_307 (O_307,N_18575,N_19101);
nor UO_308 (O_308,N_18981,N_18347);
or UO_309 (O_309,N_19453,N_18258);
and UO_310 (O_310,N_18160,N_18974);
xnor UO_311 (O_311,N_19775,N_19333);
xor UO_312 (O_312,N_18219,N_18653);
xnor UO_313 (O_313,N_18483,N_19575);
xor UO_314 (O_314,N_18062,N_18820);
or UO_315 (O_315,N_18221,N_19619);
xnor UO_316 (O_316,N_18695,N_18044);
xnor UO_317 (O_317,N_18297,N_18189);
nor UO_318 (O_318,N_18514,N_18559);
nand UO_319 (O_319,N_18067,N_18051);
or UO_320 (O_320,N_18946,N_18599);
nor UO_321 (O_321,N_19486,N_18433);
or UO_322 (O_322,N_18142,N_18544);
nand UO_323 (O_323,N_18598,N_19593);
xnor UO_324 (O_324,N_18171,N_19986);
nand UO_325 (O_325,N_19493,N_18646);
nand UO_326 (O_326,N_19978,N_18378);
and UO_327 (O_327,N_19207,N_19372);
nand UO_328 (O_328,N_18923,N_19937);
and UO_329 (O_329,N_18292,N_19711);
xnor UO_330 (O_330,N_18435,N_19085);
nor UO_331 (O_331,N_19401,N_18732);
nand UO_332 (O_332,N_18715,N_19067);
nor UO_333 (O_333,N_19544,N_19812);
nor UO_334 (O_334,N_19113,N_18228);
and UO_335 (O_335,N_19411,N_19326);
nand UO_336 (O_336,N_18927,N_18523);
and UO_337 (O_337,N_19554,N_19572);
nor UO_338 (O_338,N_18719,N_19565);
nor UO_339 (O_339,N_18170,N_19830);
xor UO_340 (O_340,N_19317,N_18217);
xnor UO_341 (O_341,N_18929,N_19214);
xor UO_342 (O_342,N_19336,N_18190);
xor UO_343 (O_343,N_19398,N_18349);
or UO_344 (O_344,N_19615,N_19809);
nand UO_345 (O_345,N_19414,N_18060);
nand UO_346 (O_346,N_18973,N_19474);
nand UO_347 (O_347,N_18922,N_18614);
or UO_348 (O_348,N_18589,N_19027);
or UO_349 (O_349,N_18307,N_19268);
or UO_350 (O_350,N_19631,N_18606);
nor UO_351 (O_351,N_18004,N_19880);
or UO_352 (O_352,N_19590,N_18970);
and UO_353 (O_353,N_18203,N_19423);
and UO_354 (O_354,N_19121,N_18061);
nor UO_355 (O_355,N_18092,N_18688);
nor UO_356 (O_356,N_19944,N_19562);
and UO_357 (O_357,N_18410,N_19260);
nor UO_358 (O_358,N_19728,N_19557);
nand UO_359 (O_359,N_18052,N_18448);
and UO_360 (O_360,N_19210,N_18857);
xnor UO_361 (O_361,N_18964,N_18816);
xor UO_362 (O_362,N_18280,N_18186);
nor UO_363 (O_363,N_18728,N_19645);
or UO_364 (O_364,N_18255,N_18391);
and UO_365 (O_365,N_18185,N_18795);
and UO_366 (O_366,N_19143,N_18244);
nor UO_367 (O_367,N_18545,N_18521);
and UO_368 (O_368,N_19510,N_18571);
or UO_369 (O_369,N_18522,N_18141);
nand UO_370 (O_370,N_19767,N_19408);
xor UO_371 (O_371,N_19803,N_19715);
or UO_372 (O_372,N_19457,N_18382);
xnor UO_373 (O_373,N_18057,N_19221);
nand UO_374 (O_374,N_18911,N_18269);
and UO_375 (O_375,N_18025,N_18999);
nor UO_376 (O_376,N_18285,N_19022);
and UO_377 (O_377,N_18667,N_19397);
nor UO_378 (O_378,N_19495,N_19598);
nor UO_379 (O_379,N_19377,N_18930);
or UO_380 (O_380,N_18803,N_18288);
or UO_381 (O_381,N_19009,N_19997);
and UO_382 (O_382,N_18380,N_18006);
and UO_383 (O_383,N_19500,N_18895);
xnor UO_384 (O_384,N_18278,N_19968);
nor UO_385 (O_385,N_18982,N_18897);
nor UO_386 (O_386,N_19471,N_18331);
and UO_387 (O_387,N_19529,N_18741);
nand UO_388 (O_388,N_19461,N_19779);
and UO_389 (O_389,N_19135,N_18294);
or UO_390 (O_390,N_18644,N_19255);
or UO_391 (O_391,N_18365,N_19741);
nor UO_392 (O_392,N_19984,N_18676);
nor UO_393 (O_393,N_19912,N_19579);
nor UO_394 (O_394,N_19742,N_18951);
xor UO_395 (O_395,N_19132,N_19882);
or UO_396 (O_396,N_19862,N_18513);
xnor UO_397 (O_397,N_18515,N_19083);
nor UO_398 (O_398,N_19379,N_18617);
nor UO_399 (O_399,N_19990,N_19062);
and UO_400 (O_400,N_19026,N_18393);
xor UO_401 (O_401,N_19019,N_19147);
xor UO_402 (O_402,N_18948,N_19905);
or UO_403 (O_403,N_19972,N_19612);
or UO_404 (O_404,N_18835,N_19249);
xnor UO_405 (O_405,N_18261,N_19814);
and UO_406 (O_406,N_19369,N_18398);
nand UO_407 (O_407,N_19864,N_18996);
or UO_408 (O_408,N_18230,N_18778);
xor UO_409 (O_409,N_19039,N_19458);
or UO_410 (O_410,N_18805,N_19153);
xnor UO_411 (O_411,N_19228,N_19674);
nand UO_412 (O_412,N_18766,N_18451);
and UO_413 (O_413,N_19097,N_18287);
nand UO_414 (O_414,N_19804,N_19884);
nand UO_415 (O_415,N_18899,N_19449);
nand UO_416 (O_416,N_18553,N_19128);
xnor UO_417 (O_417,N_18625,N_18707);
and UO_418 (O_418,N_19363,N_19957);
xnor UO_419 (O_419,N_18717,N_18271);
nor UO_420 (O_420,N_18400,N_19603);
nand UO_421 (O_421,N_18864,N_18130);
nand UO_422 (O_422,N_18005,N_18535);
or UO_423 (O_423,N_18476,N_18274);
nand UO_424 (O_424,N_19410,N_18579);
nand UO_425 (O_425,N_18358,N_18329);
xnor UO_426 (O_426,N_19373,N_18856);
xnor UO_427 (O_427,N_19908,N_19111);
xor UO_428 (O_428,N_19646,N_19816);
nor UO_429 (O_429,N_19126,N_18573);
xnor UO_430 (O_430,N_19976,N_18201);
nor UO_431 (O_431,N_19591,N_18001);
nand UO_432 (O_432,N_19914,N_19687);
nor UO_433 (O_433,N_18211,N_18146);
nand UO_434 (O_434,N_19760,N_19567);
xor UO_435 (O_435,N_18443,N_18105);
nor UO_436 (O_436,N_18183,N_19889);
xnor UO_437 (O_437,N_18032,N_18462);
xnor UO_438 (O_438,N_19043,N_19497);
xor UO_439 (O_439,N_18017,N_19736);
nand UO_440 (O_440,N_18265,N_19443);
or UO_441 (O_441,N_18540,N_18222);
or UO_442 (O_442,N_19578,N_18322);
xnor UO_443 (O_443,N_19349,N_18427);
and UO_444 (O_444,N_19155,N_19334);
or UO_445 (O_445,N_18442,N_18527);
nor UO_446 (O_446,N_19719,N_19858);
and UO_447 (O_447,N_18181,N_18828);
nand UO_448 (O_448,N_18238,N_19999);
nor UO_449 (O_449,N_18830,N_19561);
nor UO_450 (O_450,N_19797,N_18738);
and UO_451 (O_451,N_18752,N_19770);
nand UO_452 (O_452,N_18782,N_18876);
nand UO_453 (O_453,N_18395,N_19581);
nor UO_454 (O_454,N_18120,N_19693);
nand UO_455 (O_455,N_19989,N_19189);
nor UO_456 (O_456,N_18942,N_18799);
or UO_457 (O_457,N_18853,N_19668);
or UO_458 (O_458,N_18979,N_19279);
nor UO_459 (O_459,N_18860,N_19538);
nand UO_460 (O_460,N_19485,N_18747);
nor UO_461 (O_461,N_18066,N_18822);
xor UO_462 (O_462,N_19823,N_19139);
and UO_463 (O_463,N_18703,N_19077);
and UO_464 (O_464,N_19124,N_19034);
nor UO_465 (O_465,N_18473,N_19010);
nor UO_466 (O_466,N_18471,N_18013);
and UO_467 (O_467,N_18446,N_18438);
or UO_468 (O_468,N_19654,N_19088);
xnor UO_469 (O_469,N_18670,N_19949);
nor UO_470 (O_470,N_18503,N_18692);
xnor UO_471 (O_471,N_19223,N_19758);
xnor UO_472 (O_472,N_18070,N_19089);
xnor UO_473 (O_473,N_19826,N_18566);
xor UO_474 (O_474,N_18223,N_18459);
nand UO_475 (O_475,N_19865,N_19277);
nand UO_476 (O_476,N_18788,N_18104);
nor UO_477 (O_477,N_18194,N_18968);
xnor UO_478 (O_478,N_19087,N_18330);
nor UO_479 (O_479,N_18811,N_19898);
or UO_480 (O_480,N_19031,N_18664);
nor UO_481 (O_481,N_18215,N_18774);
or UO_482 (O_482,N_19680,N_18015);
nor UO_483 (O_483,N_18997,N_18680);
nor UO_484 (O_484,N_19040,N_18900);
nand UO_485 (O_485,N_19564,N_18520);
xnor UO_486 (O_486,N_18804,N_18198);
and UO_487 (O_487,N_19212,N_19963);
or UO_488 (O_488,N_18117,N_18403);
nand UO_489 (O_489,N_18163,N_18295);
nand UO_490 (O_490,N_19566,N_18273);
or UO_491 (O_491,N_19806,N_18074);
and UO_492 (O_492,N_19897,N_18790);
nor UO_493 (O_493,N_18504,N_18213);
and UO_494 (O_494,N_18755,N_18826);
or UO_495 (O_495,N_19340,N_19446);
nand UO_496 (O_496,N_19716,N_18392);
and UO_497 (O_497,N_18114,N_18584);
xor UO_498 (O_498,N_18843,N_19420);
nand UO_499 (O_499,N_18543,N_19726);
nor UO_500 (O_500,N_18555,N_18808);
xor UO_501 (O_501,N_19608,N_19735);
or UO_502 (O_502,N_18654,N_18431);
and UO_503 (O_503,N_18090,N_18524);
or UO_504 (O_504,N_18175,N_18787);
and UO_505 (O_505,N_19734,N_18075);
nor UO_506 (O_506,N_18959,N_18157);
or UO_507 (O_507,N_19054,N_19875);
nor UO_508 (O_508,N_18824,N_18147);
and UO_509 (O_509,N_19723,N_18402);
nand UO_510 (O_510,N_18681,N_18159);
xor UO_511 (O_511,N_19119,N_18990);
or UO_512 (O_512,N_18202,N_18539);
or UO_513 (O_513,N_18600,N_18888);
nand UO_514 (O_514,N_18603,N_18910);
nor UO_515 (O_515,N_19102,N_19599);
nand UO_516 (O_516,N_19417,N_18088);
xnor UO_517 (O_517,N_19903,N_18761);
nand UO_518 (O_518,N_18306,N_19896);
and UO_519 (O_519,N_19688,N_19513);
and UO_520 (O_520,N_18713,N_18896);
nor UO_521 (O_521,N_18413,N_19643);
and UO_522 (O_522,N_18939,N_19996);
nand UO_523 (O_523,N_18583,N_19320);
xnor UO_524 (O_524,N_18534,N_18619);
nor UO_525 (O_525,N_19934,N_19297);
xor UO_526 (O_526,N_19478,N_19744);
and UO_527 (O_527,N_19669,N_18862);
or UO_528 (O_528,N_18466,N_18913);
and UO_529 (O_529,N_18890,N_19248);
xor UO_530 (O_530,N_19304,N_19425);
nand UO_531 (O_531,N_18510,N_19808);
xnor UO_532 (O_532,N_18622,N_18408);
xor UO_533 (O_533,N_18042,N_19007);
nor UO_534 (O_534,N_18672,N_19644);
nand UO_535 (O_535,N_19295,N_18859);
xnor UO_536 (O_536,N_18064,N_19725);
nand UO_537 (O_537,N_18938,N_19541);
and UO_538 (O_538,N_19046,N_18626);
or UO_539 (O_539,N_18581,N_18038);
xnor UO_540 (O_540,N_18276,N_18793);
and UO_541 (O_541,N_18769,N_18737);
or UO_542 (O_542,N_18961,N_18429);
nand UO_543 (O_543,N_19721,N_19430);
or UO_544 (O_544,N_19946,N_18674);
nor UO_545 (O_545,N_19887,N_18043);
and UO_546 (O_546,N_18564,N_18362);
or UO_547 (O_547,N_18989,N_19492);
or UO_548 (O_548,N_19967,N_18310);
or UO_549 (O_549,N_18447,N_19308);
nor UO_550 (O_550,N_19065,N_18771);
nand UO_551 (O_551,N_18056,N_18445);
or UO_552 (O_552,N_18756,N_19378);
nor UO_553 (O_553,N_19570,N_19301);
nor UO_554 (O_554,N_18003,N_18884);
and UO_555 (O_555,N_18918,N_18096);
xnor UO_556 (O_556,N_19890,N_18305);
nand UO_557 (O_557,N_18205,N_19793);
or UO_558 (O_558,N_19253,N_18458);
or UO_559 (O_559,N_19413,N_19374);
and UO_560 (O_560,N_18149,N_19070);
nor UO_561 (O_561,N_19505,N_19094);
nor UO_562 (O_562,N_18487,N_18282);
xor UO_563 (O_563,N_18955,N_19689);
xnor UO_564 (O_564,N_18685,N_19302);
nand UO_565 (O_565,N_18011,N_19522);
or UO_566 (O_566,N_19392,N_18161);
nand UO_567 (O_567,N_19795,N_19051);
nor UO_568 (O_568,N_19975,N_18477);
and UO_569 (O_569,N_18627,N_18841);
xor UO_570 (O_570,N_18572,N_19041);
nor UO_571 (O_571,N_19310,N_18345);
or UO_572 (O_572,N_19877,N_18107);
xnor UO_573 (O_573,N_18465,N_18239);
xnor UO_574 (O_574,N_19184,N_19714);
nand UO_575 (O_575,N_18775,N_19847);
xnor UO_576 (O_576,N_18420,N_19837);
nand UO_577 (O_577,N_18650,N_18940);
or UO_578 (O_578,N_18150,N_18374);
or UO_579 (O_579,N_18242,N_18815);
nor UO_580 (O_580,N_19024,N_18668);
nand UO_581 (O_581,N_19066,N_18677);
and UO_582 (O_582,N_18455,N_18123);
and UO_583 (O_583,N_18846,N_18404);
nor UO_584 (O_584,N_19059,N_19250);
nor UO_585 (O_585,N_18785,N_19161);
or UO_586 (O_586,N_18630,N_18863);
or UO_587 (O_587,N_19755,N_19490);
nand UO_588 (O_588,N_18881,N_19117);
and UO_589 (O_589,N_18943,N_18326);
xor UO_590 (O_590,N_18993,N_19036);
or UO_591 (O_591,N_18148,N_19166);
nand UO_592 (O_592,N_18953,N_19574);
nand UO_593 (O_593,N_18831,N_18870);
nand UO_594 (O_594,N_19477,N_19445);
xor UO_595 (O_595,N_19159,N_19800);
or UO_596 (O_596,N_18792,N_19239);
and UO_597 (O_597,N_19306,N_18087);
and UO_598 (O_598,N_18960,N_18643);
xnor UO_599 (O_599,N_18994,N_19399);
or UO_600 (O_600,N_19700,N_18492);
nor UO_601 (O_601,N_18173,N_18229);
nor UO_602 (O_602,N_18595,N_18698);
nor UO_603 (O_603,N_19571,N_19215);
xor UO_604 (O_604,N_19762,N_19918);
or UO_605 (O_605,N_18370,N_19507);
xnor UO_606 (O_606,N_19791,N_19264);
and UO_607 (O_607,N_18735,N_19627);
or UO_608 (O_608,N_19664,N_19563);
xnor UO_609 (O_609,N_19879,N_19290);
xnor UO_610 (O_610,N_19518,N_18958);
or UO_611 (O_611,N_18977,N_18399);
or UO_612 (O_612,N_19853,N_19171);
nand UO_613 (O_613,N_19370,N_19822);
or UO_614 (O_614,N_19855,N_19082);
or UO_615 (O_615,N_18475,N_18405);
nand UO_616 (O_616,N_18284,N_18696);
xor UO_617 (O_617,N_18565,N_18801);
nand UO_618 (O_618,N_19482,N_18020);
xnor UO_619 (O_619,N_19861,N_19527);
xor UO_620 (O_620,N_18434,N_18586);
xor UO_621 (O_621,N_18256,N_18366);
nand UO_622 (O_622,N_19840,N_19025);
nor UO_623 (O_623,N_19901,N_18124);
nand UO_624 (O_624,N_18023,N_19774);
nand UO_625 (O_625,N_18359,N_19321);
or UO_626 (O_626,N_18949,N_19740);
nor UO_627 (O_627,N_19138,N_19697);
and UO_628 (O_628,N_19426,N_18950);
xnor UO_629 (O_629,N_18907,N_19909);
and UO_630 (O_630,N_19484,N_19931);
xnor UO_631 (O_631,N_18108,N_19848);
nor UO_632 (O_632,N_18231,N_19936);
and UO_633 (O_633,N_18316,N_18027);
nor UO_634 (O_634,N_18407,N_19359);
and UO_635 (O_635,N_19945,N_19971);
or UO_636 (O_636,N_18012,N_18880);
nand UO_637 (O_637,N_18560,N_18323);
and UO_638 (O_638,N_18069,N_19269);
nor UO_639 (O_639,N_18965,N_19325);
xor UO_640 (O_640,N_19691,N_19829);
or UO_641 (O_641,N_19395,N_18550);
xnor UO_642 (O_642,N_18387,N_19549);
and UO_643 (O_643,N_18360,N_19133);
and UO_644 (O_644,N_18986,N_18768);
or UO_645 (O_645,N_18850,N_19042);
and UO_646 (O_646,N_18482,N_18086);
xor UO_647 (O_647,N_19594,N_19192);
nor UO_648 (O_648,N_19165,N_18406);
or UO_649 (O_649,N_19319,N_19400);
xnor UO_650 (O_650,N_19071,N_18554);
and UO_651 (O_651,N_19970,N_19543);
xnor UO_652 (O_652,N_19783,N_19973);
or UO_653 (O_653,N_18686,N_18773);
or UO_654 (O_654,N_19642,N_19922);
or UO_655 (O_655,N_18925,N_19469);
and UO_656 (O_656,N_18936,N_18341);
xnor UO_657 (O_657,N_19084,N_18926);
nor UO_658 (O_658,N_19244,N_19434);
xor UO_659 (O_659,N_18679,N_19569);
nand UO_660 (O_660,N_19517,N_18245);
xor UO_661 (O_661,N_19632,N_18765);
and UO_662 (O_662,N_18376,N_18343);
nand UO_663 (O_663,N_18767,N_18381);
nand UO_664 (O_664,N_18168,N_19545);
nor UO_665 (O_665,N_18509,N_18734);
nand UO_666 (O_666,N_18342,N_18733);
or UO_667 (O_667,N_18666,N_18484);
nor UO_668 (O_668,N_18154,N_19772);
xnor UO_669 (O_669,N_19844,N_18714);
nand UO_670 (O_670,N_18891,N_19350);
nand UO_671 (O_671,N_18689,N_19055);
or UO_672 (O_672,N_19353,N_19149);
xnor UO_673 (O_673,N_18840,N_19851);
or UO_674 (O_674,N_18500,N_19064);
nand UO_675 (O_675,N_18035,N_19448);
or UO_676 (O_676,N_19162,N_18739);
or UO_677 (O_677,N_19954,N_19049);
nand UO_678 (O_678,N_18629,N_18081);
nor UO_679 (O_679,N_19276,N_19129);
nand UO_680 (O_680,N_19416,N_18167);
or UO_681 (O_681,N_18367,N_18485);
xor UO_682 (O_682,N_19195,N_19488);
xor UO_683 (O_683,N_19280,N_18570);
nand UO_684 (O_684,N_18909,N_18635);
nand UO_685 (O_685,N_18077,N_18966);
xnor UO_686 (O_686,N_18537,N_19821);
and UO_687 (O_687,N_19286,N_19072);
or UO_688 (O_688,N_18098,N_18821);
or UO_689 (O_689,N_19730,N_19764);
or UO_690 (O_690,N_19915,N_18029);
nand UO_691 (O_691,N_19980,N_18758);
nand UO_692 (O_692,N_18898,N_18836);
and UO_693 (O_693,N_18952,N_19786);
or UO_694 (O_694,N_18716,N_19843);
nand UO_695 (O_695,N_19611,N_18873);
or UO_696 (O_696,N_19163,N_18418);
or UO_697 (O_697,N_18426,N_19375);
nand UO_698 (O_698,N_18558,N_19769);
and UO_699 (O_699,N_19597,N_18905);
nor UO_700 (O_700,N_18547,N_18033);
and UO_701 (O_701,N_18574,N_18914);
or UO_702 (O_702,N_18383,N_18450);
or UO_703 (O_703,N_19839,N_19878);
or UO_704 (O_704,N_19261,N_19076);
nand UO_705 (O_705,N_19501,N_18656);
and UO_706 (O_706,N_18770,N_18562);
xnor UO_707 (O_707,N_19148,N_19029);
or UO_708 (O_708,N_18351,N_18076);
nor UO_709 (O_709,N_18607,N_19782);
xnor UO_710 (O_710,N_18132,N_18983);
and UO_711 (O_711,N_18602,N_19820);
nand UO_712 (O_712,N_18397,N_19467);
nand UO_713 (O_713,N_19222,N_18548);
nand UO_714 (O_714,N_18638,N_18720);
and UO_715 (O_715,N_19352,N_19335);
nor UO_716 (O_716,N_18226,N_19489);
and UO_717 (O_717,N_19134,N_19553);
nor UO_718 (O_718,N_18422,N_18415);
xnor UO_719 (O_719,N_18813,N_19982);
and UO_720 (O_720,N_19651,N_18440);
nand UO_721 (O_721,N_19536,N_19475);
xnor UO_722 (O_722,N_19868,N_18743);
or UO_723 (O_723,N_18444,N_19169);
or UO_724 (O_724,N_19050,N_19686);
or UO_725 (O_725,N_19647,N_18298);
or UO_726 (O_726,N_19345,N_19091);
nand UO_727 (O_727,N_18618,N_18210);
and UO_728 (O_728,N_18708,N_19995);
and UO_729 (O_729,N_18045,N_18048);
and UO_730 (O_730,N_18394,N_18640);
nor UO_731 (O_731,N_18608,N_18493);
and UO_732 (O_732,N_19406,N_19278);
xor UO_733 (O_733,N_19551,N_18745);
or UO_734 (O_734,N_19356,N_19859);
xnor UO_735 (O_735,N_19140,N_19583);
nor UO_736 (O_736,N_18587,N_18121);
and UO_737 (O_737,N_18138,N_18325);
nand UO_738 (O_738,N_19617,N_18187);
and UO_739 (O_739,N_18209,N_18736);
xnor UO_740 (O_740,N_19900,N_18102);
or UO_741 (O_741,N_18542,N_18156);
or UO_742 (O_742,N_18152,N_18236);
or UO_743 (O_743,N_18683,N_18593);
xor UO_744 (O_744,N_19201,N_19857);
nand UO_745 (O_745,N_18457,N_19346);
and UO_746 (O_746,N_19605,N_19661);
xor UO_747 (O_747,N_18472,N_19825);
xor UO_748 (O_748,N_19001,N_18249);
nand UO_749 (O_749,N_18266,N_18486);
and UO_750 (O_750,N_18456,N_19676);
xnor UO_751 (O_751,N_19904,N_18991);
nor UO_752 (O_752,N_19815,N_19961);
nor UO_753 (O_753,N_18385,N_19658);
and UO_754 (O_754,N_18933,N_19472);
and UO_755 (O_755,N_18200,N_19925);
or UO_756 (O_756,N_19576,N_19098);
and UO_757 (O_757,N_19722,N_19873);
nand UO_758 (O_758,N_19616,N_19785);
and UO_759 (O_759,N_19618,N_19953);
or UO_760 (O_760,N_18634,N_19724);
nor UO_761 (O_761,N_18182,N_18162);
xor UO_762 (O_762,N_18368,N_18916);
nand UO_763 (O_763,N_18312,N_18065);
xnor UO_764 (O_764,N_18158,N_18754);
nand UO_765 (O_765,N_19145,N_18797);
and UO_766 (O_766,N_18885,N_18259);
and UO_767 (O_767,N_19582,N_18848);
nand UO_768 (O_768,N_19638,N_19503);
and UO_769 (O_769,N_19784,N_19330);
nand UO_770 (O_770,N_18613,N_18931);
nor UO_771 (O_771,N_18361,N_19738);
nand UO_772 (O_772,N_19657,N_18878);
nor UO_773 (O_773,N_19856,N_19547);
and UO_774 (O_774,N_18008,N_19275);
xnor UO_775 (O_775,N_19060,N_19323);
or UO_776 (O_776,N_18596,N_18111);
or UO_777 (O_777,N_18072,N_18232);
nor UO_778 (O_778,N_18489,N_18673);
xor UO_779 (O_779,N_18723,N_18759);
or UO_780 (O_780,N_19473,N_19920);
nand UO_781 (O_781,N_19123,N_19294);
nand UO_782 (O_782,N_18842,N_18998);
and UO_783 (O_783,N_18243,N_19218);
nor UO_784 (O_784,N_19389,N_19981);
or UO_785 (O_785,N_19796,N_18227);
xor UO_786 (O_786,N_19131,N_19673);
xnor UO_787 (O_787,N_19753,N_18340);
or UO_788 (O_788,N_19240,N_19955);
and UO_789 (O_789,N_19146,N_19601);
or UO_790 (O_790,N_18286,N_19828);
xnor UO_791 (O_791,N_19860,N_18631);
xor UO_792 (O_792,N_18388,N_19281);
nor UO_793 (O_793,N_18191,N_18122);
xnor UO_794 (O_794,N_19237,N_19948);
and UO_795 (O_795,N_19876,N_19683);
nand UO_796 (O_796,N_19958,N_18116);
and UO_797 (O_797,N_19845,N_18601);
xnor UO_798 (O_798,N_19251,N_18384);
nor UO_799 (O_799,N_18093,N_18053);
or UO_800 (O_800,N_18531,N_18460);
and UO_801 (O_801,N_18174,N_18796);
nand UO_802 (O_802,N_18886,N_19480);
and UO_803 (O_803,N_18346,N_19177);
and UO_804 (O_804,N_19173,N_19835);
nand UO_805 (O_805,N_19623,N_19951);
or UO_806 (O_806,N_18257,N_18505);
nand UO_807 (O_807,N_18195,N_19927);
nor UO_808 (O_808,N_19409,N_18063);
nand UO_809 (O_809,N_18073,N_18178);
and UO_810 (O_810,N_18263,N_19913);
or UO_811 (O_811,N_19002,N_19291);
and UO_812 (O_812,N_19703,N_19932);
and UO_813 (O_813,N_19438,N_19917);
xor UO_814 (O_814,N_18592,N_19891);
xor UO_815 (O_815,N_19737,N_18491);
and UO_816 (O_816,N_18016,N_18494);
nand UO_817 (O_817,N_19093,N_19639);
and UO_818 (O_818,N_18915,N_18597);
nor UO_819 (O_819,N_19105,N_19692);
xnor UO_820 (O_820,N_18283,N_18026);
nand UO_821 (O_821,N_18281,N_19179);
xor UO_822 (O_822,N_19380,N_18724);
nand UO_823 (O_823,N_19799,N_18937);
and UO_824 (O_824,N_18430,N_18000);
and UO_825 (O_825,N_19044,N_18165);
and UO_826 (O_826,N_19348,N_19038);
nand UO_827 (O_827,N_18437,N_19768);
or UO_828 (O_828,N_18139,N_18002);
or UO_829 (O_829,N_18731,N_18757);
and UO_830 (O_830,N_19393,N_19888);
nor UO_831 (O_831,N_18480,N_19817);
nand UO_832 (O_832,N_18461,N_19923);
nor UO_833 (O_833,N_18690,N_18268);
nor UO_834 (O_834,N_18352,N_18235);
xnor UO_835 (O_835,N_19602,N_19107);
nor UO_836 (O_836,N_19293,N_18155);
xor UO_837 (O_837,N_19911,N_19987);
nand UO_838 (O_838,N_18749,N_18113);
nor UO_839 (O_839,N_19752,N_18849);
nand UO_840 (O_840,N_18373,N_18218);
xnor UO_841 (O_841,N_19110,N_19008);
xnor UO_842 (O_842,N_19739,N_18920);
nand UO_843 (O_843,N_18357,N_19998);
xor UO_844 (O_844,N_18532,N_19152);
nand UO_845 (O_845,N_18889,N_19164);
xnor UO_846 (O_846,N_19660,N_18637);
xor UO_847 (O_847,N_18919,N_19013);
and UO_848 (O_848,N_19442,N_19516);
and UO_849 (O_849,N_19600,N_19916);
nand UO_850 (O_850,N_19158,N_19383);
or UO_851 (O_851,N_19867,N_18478);
nor UO_852 (O_852,N_19157,N_19985);
xor UO_853 (O_853,N_18917,N_18333);
xnor UO_854 (O_854,N_19208,N_19463);
nand UO_855 (O_855,N_18525,N_18978);
xor UO_856 (O_856,N_19679,N_18419);
and UO_857 (O_857,N_19506,N_19504);
xnor UO_858 (O_858,N_18290,N_19694);
or UO_859 (O_859,N_19892,N_19531);
and UO_860 (O_860,N_18838,N_18034);
xnor UO_861 (O_861,N_19670,N_19342);
or UO_862 (O_862,N_19757,N_19606);
xor UO_863 (O_863,N_18131,N_18781);
and UO_864 (O_864,N_19977,N_18868);
xor UO_865 (O_865,N_19183,N_19966);
or UO_866 (O_866,N_19613,N_18847);
and UO_867 (O_867,N_19940,N_19267);
nor UO_868 (O_868,N_18296,N_18519);
and UO_869 (O_869,N_19805,N_19926);
xnor UO_870 (O_870,N_18039,N_18246);
xor UO_871 (O_871,N_19307,N_19659);
nand UO_872 (O_872,N_18877,N_18954);
nor UO_873 (O_873,N_19272,N_18172);
nand UO_874 (O_874,N_18036,N_19056);
nor UO_875 (O_875,N_19376,N_18335);
xnor UO_876 (O_876,N_19630,N_19284);
xor UO_877 (O_877,N_19943,N_19792);
and UO_878 (O_878,N_18470,N_19243);
or UO_879 (O_879,N_19227,N_18055);
xor UO_880 (O_880,N_19351,N_18463);
or UO_881 (O_881,N_19684,N_19114);
and UO_882 (O_882,N_19648,N_19708);
nor UO_883 (O_883,N_19831,N_19542);
or UO_884 (O_884,N_19802,N_18254);
nand UO_885 (O_885,N_18100,N_19328);
or UO_886 (O_886,N_18844,N_18126);
and UO_887 (O_887,N_19270,N_19720);
and UO_888 (O_888,N_19032,N_19012);
nand UO_889 (O_889,N_19194,N_19068);
nor UO_890 (O_890,N_19584,N_19667);
and UO_891 (O_891,N_19698,N_18578);
and UO_892 (O_892,N_19636,N_19649);
and UO_893 (O_893,N_18118,N_19568);
nand UO_894 (O_894,N_19895,N_19052);
or UO_895 (O_895,N_19508,N_19466);
nor UO_896 (O_896,N_18332,N_19633);
nor UO_897 (O_897,N_18439,N_18499);
nand UO_898 (O_898,N_18328,N_19841);
and UO_899 (O_899,N_19181,N_18327);
xnor UO_900 (O_900,N_19160,N_19230);
nor UO_901 (O_901,N_18944,N_19712);
nor UO_902 (O_902,N_18762,N_18865);
nand UO_903 (O_903,N_19347,N_19191);
nor UO_904 (O_904,N_18389,N_19178);
and UO_905 (O_905,N_19754,N_19312);
nand UO_906 (O_906,N_18112,N_19745);
xor UO_907 (O_907,N_18663,N_18561);
xnor UO_908 (O_908,N_19427,N_18091);
xnor UO_909 (O_909,N_19810,N_19063);
nor UO_910 (O_910,N_19626,N_18109);
nor UO_911 (O_911,N_18338,N_19224);
nor UO_912 (O_912,N_19938,N_19487);
and UO_913 (O_913,N_19418,N_18854);
nand UO_914 (O_914,N_19732,N_19713);
or UO_915 (O_915,N_19863,N_19455);
nor UO_916 (O_916,N_18507,N_18825);
nand UO_917 (O_917,N_18037,N_19727);
and UO_918 (O_918,N_19436,N_18697);
and UO_919 (O_919,N_18151,N_19871);
and UO_920 (O_920,N_19962,N_19509);
and UO_921 (O_921,N_19030,N_19057);
and UO_922 (O_922,N_19560,N_18665);
nand UO_923 (O_923,N_19299,N_18605);
nor UO_924 (O_924,N_18424,N_19415);
xor UO_925 (O_925,N_18712,N_18272);
nand UO_926 (O_926,N_18549,N_19174);
xor UO_927 (O_927,N_19004,N_18216);
xnor UO_928 (O_928,N_18552,N_19424);
nand UO_929 (O_929,N_19015,N_18436);
nand UO_930 (O_930,N_19854,N_19765);
nand UO_931 (O_931,N_18339,N_18699);
or UO_932 (O_932,N_19014,N_18095);
nand UO_933 (O_933,N_19435,N_18528);
xnor UO_934 (O_934,N_18874,N_19702);
xor UO_935 (O_935,N_18336,N_18136);
xnor UO_936 (O_936,N_19023,N_18611);
xor UO_937 (O_937,N_19993,N_19454);
xor UO_938 (O_938,N_19881,N_18652);
or UO_939 (O_939,N_19464,N_18641);
nor UO_940 (O_940,N_18585,N_19819);
and UO_941 (O_941,N_18947,N_19872);
nor UO_942 (O_942,N_19112,N_19663);
nor UO_943 (O_943,N_18750,N_19747);
nand UO_944 (O_944,N_18945,N_18106);
and UO_945 (O_945,N_19271,N_18705);
nand UO_946 (O_946,N_18748,N_19232);
xnor UO_947 (O_947,N_19979,N_19894);
or UO_948 (O_948,N_19003,N_18845);
nand UO_949 (O_949,N_19838,N_19756);
or UO_950 (O_950,N_18469,N_18321);
and UO_951 (O_951,N_19367,N_18502);
xor UO_952 (O_952,N_19994,N_18763);
xnor UO_953 (O_953,N_19360,N_18199);
nand UO_954 (O_954,N_18892,N_19220);
nor UO_955 (O_955,N_18984,N_19678);
nor UO_956 (O_956,N_19364,N_19344);
nand UO_957 (O_957,N_18386,N_19552);
and UO_958 (O_958,N_18904,N_18214);
nand UO_959 (O_959,N_18887,N_19695);
and UO_960 (O_960,N_18372,N_19462);
and UO_961 (O_961,N_19502,N_19524);
nand UO_962 (O_962,N_18253,N_18119);
nor UO_963 (O_963,N_19343,N_19262);
nor UO_964 (O_964,N_19329,N_18300);
nor UO_965 (O_965,N_19640,N_19710);
nor UO_966 (O_966,N_19204,N_18467);
xnor UO_967 (O_967,N_18103,N_18453);
and UO_968 (O_968,N_18633,N_18353);
nand UO_969 (O_969,N_19234,N_19773);
xor UO_970 (O_970,N_19974,N_18875);
xnor UO_971 (O_971,N_19122,N_19073);
nand UO_972 (O_972,N_18474,N_18814);
and UO_973 (O_973,N_18620,N_18883);
xnor UO_974 (O_974,N_18594,N_19850);
xor UO_975 (O_975,N_18479,N_18740);
or UO_976 (O_976,N_18517,N_18498);
and UO_977 (O_977,N_18693,N_19273);
and UO_978 (O_978,N_18872,N_19137);
xnor UO_979 (O_979,N_18556,N_18985);
xnor UO_980 (O_980,N_19357,N_18490);
xnor UO_981 (O_981,N_18852,N_18018);
xnor UO_982 (O_982,N_18379,N_18301);
nand UO_983 (O_983,N_19573,N_19316);
and UO_984 (O_984,N_19429,N_19637);
or UO_985 (O_985,N_19749,N_18188);
and UO_986 (O_986,N_18233,N_18812);
xnor UO_987 (O_987,N_19652,N_19780);
nand UO_988 (O_988,N_18624,N_18866);
nor UO_989 (O_989,N_19362,N_18179);
and UO_990 (O_990,N_19428,N_19257);
xnor UO_991 (O_991,N_19447,N_19874);
nand UO_992 (O_992,N_19285,N_19404);
and UO_993 (O_993,N_19496,N_18085);
and UO_994 (O_994,N_19225,N_18839);
xor UO_995 (O_995,N_19528,N_18569);
and UO_996 (O_996,N_19704,N_19437);
nand UO_997 (O_997,N_19402,N_19656);
and UO_998 (O_998,N_18481,N_18691);
nand UO_999 (O_999,N_19479,N_18580);
and UO_1000 (O_1000,N_18054,N_18289);
nand UO_1001 (O_1001,N_18064,N_19513);
nand UO_1002 (O_1002,N_19721,N_18346);
nor UO_1003 (O_1003,N_18000,N_18100);
nand UO_1004 (O_1004,N_18425,N_18621);
or UO_1005 (O_1005,N_19630,N_19985);
or UO_1006 (O_1006,N_18072,N_18011);
and UO_1007 (O_1007,N_19909,N_18811);
nor UO_1008 (O_1008,N_18397,N_18937);
and UO_1009 (O_1009,N_18520,N_18332);
or UO_1010 (O_1010,N_19270,N_18273);
xnor UO_1011 (O_1011,N_18093,N_19514);
or UO_1012 (O_1012,N_19975,N_18818);
and UO_1013 (O_1013,N_19918,N_19933);
and UO_1014 (O_1014,N_19159,N_19396);
nor UO_1015 (O_1015,N_18088,N_19666);
xor UO_1016 (O_1016,N_18887,N_18933);
nand UO_1017 (O_1017,N_18777,N_19233);
and UO_1018 (O_1018,N_19317,N_18210);
nor UO_1019 (O_1019,N_18702,N_18722);
and UO_1020 (O_1020,N_19883,N_18412);
nor UO_1021 (O_1021,N_18627,N_19494);
and UO_1022 (O_1022,N_18427,N_19003);
nor UO_1023 (O_1023,N_19182,N_18115);
xor UO_1024 (O_1024,N_19292,N_18723);
nor UO_1025 (O_1025,N_19890,N_19888);
nand UO_1026 (O_1026,N_18706,N_18883);
nand UO_1027 (O_1027,N_18371,N_19903);
or UO_1028 (O_1028,N_18739,N_19338);
nor UO_1029 (O_1029,N_18408,N_19313);
or UO_1030 (O_1030,N_19019,N_18990);
and UO_1031 (O_1031,N_19800,N_19455);
xor UO_1032 (O_1032,N_19501,N_18398);
nand UO_1033 (O_1033,N_19365,N_18075);
nor UO_1034 (O_1034,N_18983,N_18937);
nor UO_1035 (O_1035,N_18905,N_18105);
nor UO_1036 (O_1036,N_18523,N_19370);
and UO_1037 (O_1037,N_19850,N_19210);
nand UO_1038 (O_1038,N_18445,N_19905);
or UO_1039 (O_1039,N_19317,N_18277);
and UO_1040 (O_1040,N_19802,N_19345);
or UO_1041 (O_1041,N_19356,N_18428);
and UO_1042 (O_1042,N_19932,N_19138);
or UO_1043 (O_1043,N_19839,N_18883);
nor UO_1044 (O_1044,N_18834,N_19867);
nand UO_1045 (O_1045,N_19689,N_18846);
or UO_1046 (O_1046,N_19380,N_19062);
nor UO_1047 (O_1047,N_19802,N_19983);
or UO_1048 (O_1048,N_19538,N_18526);
or UO_1049 (O_1049,N_18199,N_19169);
nor UO_1050 (O_1050,N_19196,N_18412);
and UO_1051 (O_1051,N_19932,N_18543);
or UO_1052 (O_1052,N_18596,N_18765);
and UO_1053 (O_1053,N_19229,N_19091);
nand UO_1054 (O_1054,N_19025,N_18184);
and UO_1055 (O_1055,N_19823,N_19780);
nor UO_1056 (O_1056,N_18035,N_18466);
and UO_1057 (O_1057,N_18950,N_19641);
nor UO_1058 (O_1058,N_19507,N_18474);
nand UO_1059 (O_1059,N_18634,N_19958);
or UO_1060 (O_1060,N_18119,N_18590);
or UO_1061 (O_1061,N_19071,N_18062);
nor UO_1062 (O_1062,N_19683,N_18028);
or UO_1063 (O_1063,N_19672,N_18162);
or UO_1064 (O_1064,N_19520,N_19806);
and UO_1065 (O_1065,N_19050,N_18379);
xnor UO_1066 (O_1066,N_18800,N_19799);
nor UO_1067 (O_1067,N_18323,N_19232);
nand UO_1068 (O_1068,N_19948,N_18280);
nand UO_1069 (O_1069,N_19022,N_19145);
nand UO_1070 (O_1070,N_19814,N_18245);
xnor UO_1071 (O_1071,N_19380,N_18662);
nor UO_1072 (O_1072,N_18862,N_19604);
or UO_1073 (O_1073,N_19780,N_19051);
nor UO_1074 (O_1074,N_19309,N_19031);
xor UO_1075 (O_1075,N_19095,N_18828);
and UO_1076 (O_1076,N_18229,N_19613);
and UO_1077 (O_1077,N_19813,N_19725);
nor UO_1078 (O_1078,N_18567,N_19653);
or UO_1079 (O_1079,N_19665,N_19066);
or UO_1080 (O_1080,N_18823,N_19794);
nand UO_1081 (O_1081,N_19681,N_18524);
nand UO_1082 (O_1082,N_18373,N_18321);
nand UO_1083 (O_1083,N_18508,N_18541);
nand UO_1084 (O_1084,N_18668,N_18118);
or UO_1085 (O_1085,N_18909,N_19454);
or UO_1086 (O_1086,N_18960,N_19629);
and UO_1087 (O_1087,N_18427,N_18844);
nand UO_1088 (O_1088,N_19253,N_19191);
or UO_1089 (O_1089,N_19615,N_19644);
xnor UO_1090 (O_1090,N_19280,N_18834);
or UO_1091 (O_1091,N_19811,N_18598);
nand UO_1092 (O_1092,N_18979,N_18938);
and UO_1093 (O_1093,N_18359,N_18124);
xor UO_1094 (O_1094,N_19360,N_18124);
nor UO_1095 (O_1095,N_18067,N_19565);
nand UO_1096 (O_1096,N_18768,N_18246);
nand UO_1097 (O_1097,N_19704,N_19064);
or UO_1098 (O_1098,N_19866,N_19376);
and UO_1099 (O_1099,N_19675,N_19491);
and UO_1100 (O_1100,N_19469,N_19544);
xnor UO_1101 (O_1101,N_19598,N_18181);
xor UO_1102 (O_1102,N_19523,N_18865);
and UO_1103 (O_1103,N_18848,N_19071);
and UO_1104 (O_1104,N_18775,N_18374);
xor UO_1105 (O_1105,N_18293,N_18646);
xor UO_1106 (O_1106,N_18114,N_18476);
or UO_1107 (O_1107,N_18985,N_19569);
or UO_1108 (O_1108,N_19261,N_19138);
xor UO_1109 (O_1109,N_19441,N_19660);
or UO_1110 (O_1110,N_19149,N_18630);
or UO_1111 (O_1111,N_19301,N_19868);
nand UO_1112 (O_1112,N_18543,N_18465);
and UO_1113 (O_1113,N_18133,N_18004);
xor UO_1114 (O_1114,N_19516,N_18390);
and UO_1115 (O_1115,N_19061,N_18806);
nand UO_1116 (O_1116,N_19052,N_19012);
or UO_1117 (O_1117,N_18923,N_19090);
xor UO_1118 (O_1118,N_18289,N_18554);
and UO_1119 (O_1119,N_19789,N_19230);
xor UO_1120 (O_1120,N_18743,N_19371);
and UO_1121 (O_1121,N_19557,N_18353);
xnor UO_1122 (O_1122,N_19124,N_19735);
nor UO_1123 (O_1123,N_19573,N_19274);
nand UO_1124 (O_1124,N_19044,N_19148);
xnor UO_1125 (O_1125,N_18000,N_19034);
nor UO_1126 (O_1126,N_19616,N_19047);
nand UO_1127 (O_1127,N_18210,N_19826);
xnor UO_1128 (O_1128,N_18841,N_19081);
nor UO_1129 (O_1129,N_19360,N_18196);
nor UO_1130 (O_1130,N_19487,N_18572);
nand UO_1131 (O_1131,N_19040,N_18263);
xnor UO_1132 (O_1132,N_19491,N_19555);
nor UO_1133 (O_1133,N_19868,N_19308);
nor UO_1134 (O_1134,N_18582,N_18716);
and UO_1135 (O_1135,N_19310,N_19012);
or UO_1136 (O_1136,N_19142,N_18748);
or UO_1137 (O_1137,N_18968,N_18329);
or UO_1138 (O_1138,N_18725,N_19200);
or UO_1139 (O_1139,N_18891,N_19140);
xnor UO_1140 (O_1140,N_18425,N_18686);
and UO_1141 (O_1141,N_18113,N_18734);
nand UO_1142 (O_1142,N_18143,N_18697);
xnor UO_1143 (O_1143,N_18033,N_18021);
or UO_1144 (O_1144,N_18072,N_18545);
and UO_1145 (O_1145,N_19838,N_19766);
or UO_1146 (O_1146,N_18228,N_19915);
or UO_1147 (O_1147,N_19803,N_18371);
and UO_1148 (O_1148,N_18712,N_18567);
xnor UO_1149 (O_1149,N_19117,N_19552);
nor UO_1150 (O_1150,N_19350,N_18691);
and UO_1151 (O_1151,N_18059,N_18204);
or UO_1152 (O_1152,N_18852,N_19861);
nand UO_1153 (O_1153,N_19456,N_19319);
and UO_1154 (O_1154,N_19808,N_19441);
nor UO_1155 (O_1155,N_19939,N_19008);
nand UO_1156 (O_1156,N_18616,N_19783);
nand UO_1157 (O_1157,N_18611,N_18787);
and UO_1158 (O_1158,N_18304,N_18595);
or UO_1159 (O_1159,N_18752,N_19541);
nor UO_1160 (O_1160,N_19572,N_19055);
and UO_1161 (O_1161,N_18482,N_18578);
nor UO_1162 (O_1162,N_19671,N_18838);
nor UO_1163 (O_1163,N_18011,N_19366);
xor UO_1164 (O_1164,N_18693,N_18110);
nand UO_1165 (O_1165,N_19586,N_18612);
or UO_1166 (O_1166,N_19615,N_19378);
xnor UO_1167 (O_1167,N_19750,N_18998);
nor UO_1168 (O_1168,N_19322,N_19488);
nor UO_1169 (O_1169,N_19106,N_18119);
and UO_1170 (O_1170,N_18713,N_19687);
nand UO_1171 (O_1171,N_18574,N_19365);
nor UO_1172 (O_1172,N_19957,N_19171);
xnor UO_1173 (O_1173,N_19608,N_19013);
nand UO_1174 (O_1174,N_18226,N_18315);
or UO_1175 (O_1175,N_18230,N_19195);
and UO_1176 (O_1176,N_19387,N_18089);
xor UO_1177 (O_1177,N_19566,N_19713);
nor UO_1178 (O_1178,N_19027,N_19219);
nor UO_1179 (O_1179,N_19221,N_19306);
nand UO_1180 (O_1180,N_19708,N_19765);
and UO_1181 (O_1181,N_19083,N_18044);
or UO_1182 (O_1182,N_18967,N_19614);
and UO_1183 (O_1183,N_19011,N_19019);
or UO_1184 (O_1184,N_18214,N_18339);
nand UO_1185 (O_1185,N_19354,N_18404);
xor UO_1186 (O_1186,N_19999,N_18314);
nand UO_1187 (O_1187,N_18402,N_19981);
and UO_1188 (O_1188,N_19102,N_19724);
and UO_1189 (O_1189,N_19334,N_19501);
nor UO_1190 (O_1190,N_19171,N_18710);
xnor UO_1191 (O_1191,N_19645,N_19466);
nor UO_1192 (O_1192,N_18353,N_19763);
nor UO_1193 (O_1193,N_18010,N_18336);
xnor UO_1194 (O_1194,N_19267,N_18746);
xnor UO_1195 (O_1195,N_19450,N_19633);
nand UO_1196 (O_1196,N_18121,N_19796);
nand UO_1197 (O_1197,N_19945,N_19731);
and UO_1198 (O_1198,N_19419,N_18739);
nor UO_1199 (O_1199,N_18848,N_18660);
and UO_1200 (O_1200,N_18409,N_18379);
or UO_1201 (O_1201,N_18646,N_18531);
xor UO_1202 (O_1202,N_18410,N_19784);
and UO_1203 (O_1203,N_18430,N_18673);
xor UO_1204 (O_1204,N_19992,N_18646);
or UO_1205 (O_1205,N_18684,N_19619);
or UO_1206 (O_1206,N_18797,N_18924);
nand UO_1207 (O_1207,N_19751,N_18572);
nand UO_1208 (O_1208,N_19307,N_19915);
nor UO_1209 (O_1209,N_18735,N_19450);
xnor UO_1210 (O_1210,N_19247,N_18297);
or UO_1211 (O_1211,N_19940,N_18399);
xor UO_1212 (O_1212,N_18264,N_18265);
xor UO_1213 (O_1213,N_19234,N_18650);
nand UO_1214 (O_1214,N_19933,N_19027);
nand UO_1215 (O_1215,N_18595,N_19617);
nand UO_1216 (O_1216,N_18504,N_18699);
xor UO_1217 (O_1217,N_19161,N_18535);
nor UO_1218 (O_1218,N_19326,N_18675);
or UO_1219 (O_1219,N_18682,N_19155);
nand UO_1220 (O_1220,N_19716,N_18201);
xor UO_1221 (O_1221,N_18678,N_18874);
nand UO_1222 (O_1222,N_18878,N_19341);
nor UO_1223 (O_1223,N_19779,N_18030);
and UO_1224 (O_1224,N_19729,N_19959);
and UO_1225 (O_1225,N_18267,N_18152);
xnor UO_1226 (O_1226,N_18727,N_19032);
nand UO_1227 (O_1227,N_19055,N_19495);
or UO_1228 (O_1228,N_19803,N_18843);
and UO_1229 (O_1229,N_18770,N_18613);
or UO_1230 (O_1230,N_19752,N_18395);
xnor UO_1231 (O_1231,N_18202,N_19589);
or UO_1232 (O_1232,N_18572,N_19122);
or UO_1233 (O_1233,N_18699,N_19505);
and UO_1234 (O_1234,N_18622,N_19949);
or UO_1235 (O_1235,N_18892,N_19966);
xnor UO_1236 (O_1236,N_18512,N_19872);
or UO_1237 (O_1237,N_19357,N_18900);
or UO_1238 (O_1238,N_18553,N_18537);
nor UO_1239 (O_1239,N_18447,N_19798);
or UO_1240 (O_1240,N_18232,N_19078);
nand UO_1241 (O_1241,N_19615,N_18739);
xor UO_1242 (O_1242,N_18141,N_18545);
or UO_1243 (O_1243,N_19500,N_19084);
or UO_1244 (O_1244,N_19427,N_19423);
or UO_1245 (O_1245,N_19568,N_18637);
and UO_1246 (O_1246,N_19345,N_18971);
or UO_1247 (O_1247,N_19356,N_18077);
xnor UO_1248 (O_1248,N_18379,N_18228);
nand UO_1249 (O_1249,N_18639,N_19364);
nand UO_1250 (O_1250,N_18406,N_19856);
xor UO_1251 (O_1251,N_19961,N_18945);
and UO_1252 (O_1252,N_18237,N_18855);
nand UO_1253 (O_1253,N_18939,N_18149);
nor UO_1254 (O_1254,N_19671,N_18568);
xnor UO_1255 (O_1255,N_19469,N_18251);
or UO_1256 (O_1256,N_19290,N_18653);
nand UO_1257 (O_1257,N_18821,N_19585);
xor UO_1258 (O_1258,N_18615,N_18669);
and UO_1259 (O_1259,N_18644,N_18041);
nand UO_1260 (O_1260,N_19217,N_18951);
nor UO_1261 (O_1261,N_18912,N_19251);
nand UO_1262 (O_1262,N_19228,N_19574);
or UO_1263 (O_1263,N_18454,N_19060);
nand UO_1264 (O_1264,N_18456,N_18491);
nand UO_1265 (O_1265,N_19793,N_18212);
nor UO_1266 (O_1266,N_19311,N_18259);
nor UO_1267 (O_1267,N_18973,N_18180);
and UO_1268 (O_1268,N_19783,N_18542);
or UO_1269 (O_1269,N_18454,N_19011);
xor UO_1270 (O_1270,N_18571,N_18434);
nor UO_1271 (O_1271,N_18545,N_18126);
or UO_1272 (O_1272,N_19957,N_18277);
nor UO_1273 (O_1273,N_18341,N_18883);
and UO_1274 (O_1274,N_18406,N_19831);
nand UO_1275 (O_1275,N_18218,N_18156);
nand UO_1276 (O_1276,N_18076,N_19137);
nand UO_1277 (O_1277,N_19590,N_19177);
or UO_1278 (O_1278,N_19672,N_19894);
nor UO_1279 (O_1279,N_19007,N_19159);
nor UO_1280 (O_1280,N_19679,N_18557);
xor UO_1281 (O_1281,N_19522,N_19263);
and UO_1282 (O_1282,N_18743,N_19207);
and UO_1283 (O_1283,N_18072,N_18328);
nor UO_1284 (O_1284,N_18098,N_19277);
nor UO_1285 (O_1285,N_19482,N_19428);
or UO_1286 (O_1286,N_19079,N_19604);
or UO_1287 (O_1287,N_18574,N_18791);
and UO_1288 (O_1288,N_18214,N_19670);
xor UO_1289 (O_1289,N_19679,N_18379);
or UO_1290 (O_1290,N_19992,N_18530);
nand UO_1291 (O_1291,N_18262,N_19397);
nand UO_1292 (O_1292,N_19575,N_18195);
xor UO_1293 (O_1293,N_18285,N_18593);
xor UO_1294 (O_1294,N_18786,N_18986);
nor UO_1295 (O_1295,N_18589,N_18884);
nand UO_1296 (O_1296,N_18789,N_18364);
xor UO_1297 (O_1297,N_19210,N_19116);
nand UO_1298 (O_1298,N_19408,N_18351);
or UO_1299 (O_1299,N_19603,N_18039);
nand UO_1300 (O_1300,N_19322,N_18215);
nor UO_1301 (O_1301,N_18165,N_18925);
nand UO_1302 (O_1302,N_18392,N_19487);
or UO_1303 (O_1303,N_18047,N_18525);
or UO_1304 (O_1304,N_18430,N_19153);
xor UO_1305 (O_1305,N_19713,N_19761);
nor UO_1306 (O_1306,N_19043,N_18121);
and UO_1307 (O_1307,N_19147,N_19808);
and UO_1308 (O_1308,N_19512,N_19650);
or UO_1309 (O_1309,N_18866,N_18317);
or UO_1310 (O_1310,N_18401,N_18369);
nand UO_1311 (O_1311,N_19404,N_18714);
xor UO_1312 (O_1312,N_18379,N_19644);
nand UO_1313 (O_1313,N_19845,N_19768);
or UO_1314 (O_1314,N_19581,N_18613);
nand UO_1315 (O_1315,N_19249,N_18996);
and UO_1316 (O_1316,N_18693,N_18882);
nand UO_1317 (O_1317,N_19870,N_19696);
xnor UO_1318 (O_1318,N_18874,N_18234);
xor UO_1319 (O_1319,N_19500,N_18113);
and UO_1320 (O_1320,N_18918,N_19599);
nand UO_1321 (O_1321,N_19967,N_19706);
or UO_1322 (O_1322,N_19728,N_18262);
nand UO_1323 (O_1323,N_18932,N_18639);
xor UO_1324 (O_1324,N_18883,N_19522);
or UO_1325 (O_1325,N_18033,N_18517);
xnor UO_1326 (O_1326,N_19470,N_19381);
xor UO_1327 (O_1327,N_18495,N_18475);
nor UO_1328 (O_1328,N_19028,N_19870);
nor UO_1329 (O_1329,N_18268,N_18062);
or UO_1330 (O_1330,N_18403,N_18243);
nor UO_1331 (O_1331,N_19110,N_18861);
nand UO_1332 (O_1332,N_18327,N_19047);
or UO_1333 (O_1333,N_18686,N_19456);
and UO_1334 (O_1334,N_19164,N_18200);
and UO_1335 (O_1335,N_18550,N_19304);
or UO_1336 (O_1336,N_18182,N_18183);
xnor UO_1337 (O_1337,N_18877,N_18414);
nand UO_1338 (O_1338,N_19365,N_18483);
xnor UO_1339 (O_1339,N_19833,N_19588);
and UO_1340 (O_1340,N_18512,N_19876);
nand UO_1341 (O_1341,N_18962,N_19062);
nand UO_1342 (O_1342,N_18286,N_18695);
and UO_1343 (O_1343,N_19703,N_18410);
or UO_1344 (O_1344,N_19687,N_18608);
nor UO_1345 (O_1345,N_19097,N_18872);
nand UO_1346 (O_1346,N_18459,N_19760);
nor UO_1347 (O_1347,N_19248,N_18986);
nor UO_1348 (O_1348,N_18150,N_18112);
nor UO_1349 (O_1349,N_19693,N_18677);
and UO_1350 (O_1350,N_18288,N_19483);
xor UO_1351 (O_1351,N_18617,N_18132);
and UO_1352 (O_1352,N_18530,N_18565);
xnor UO_1353 (O_1353,N_18380,N_18231);
nand UO_1354 (O_1354,N_18833,N_19837);
xor UO_1355 (O_1355,N_19369,N_18373);
nor UO_1356 (O_1356,N_19273,N_18201);
nor UO_1357 (O_1357,N_19370,N_18271);
nand UO_1358 (O_1358,N_19624,N_19934);
xnor UO_1359 (O_1359,N_19387,N_19262);
xnor UO_1360 (O_1360,N_18322,N_18289);
xnor UO_1361 (O_1361,N_18753,N_19453);
nor UO_1362 (O_1362,N_18781,N_18571);
nor UO_1363 (O_1363,N_19464,N_19917);
and UO_1364 (O_1364,N_18251,N_19673);
or UO_1365 (O_1365,N_18244,N_18458);
and UO_1366 (O_1366,N_18812,N_18331);
or UO_1367 (O_1367,N_18900,N_19768);
xnor UO_1368 (O_1368,N_18158,N_19812);
and UO_1369 (O_1369,N_19272,N_19038);
or UO_1370 (O_1370,N_18483,N_18847);
or UO_1371 (O_1371,N_18267,N_18141);
and UO_1372 (O_1372,N_19516,N_19958);
and UO_1373 (O_1373,N_19658,N_19638);
and UO_1374 (O_1374,N_19130,N_19315);
nand UO_1375 (O_1375,N_18401,N_18603);
xnor UO_1376 (O_1376,N_18096,N_18166);
or UO_1377 (O_1377,N_19601,N_18760);
nor UO_1378 (O_1378,N_19804,N_19988);
xnor UO_1379 (O_1379,N_18541,N_19217);
or UO_1380 (O_1380,N_19627,N_19686);
nor UO_1381 (O_1381,N_18174,N_18483);
and UO_1382 (O_1382,N_18233,N_19514);
xnor UO_1383 (O_1383,N_19874,N_18354);
xnor UO_1384 (O_1384,N_19307,N_18537);
or UO_1385 (O_1385,N_18949,N_19390);
xnor UO_1386 (O_1386,N_19112,N_18915);
or UO_1387 (O_1387,N_18580,N_19164);
and UO_1388 (O_1388,N_18717,N_19587);
xor UO_1389 (O_1389,N_19875,N_18793);
xor UO_1390 (O_1390,N_19446,N_19109);
nand UO_1391 (O_1391,N_19321,N_19173);
and UO_1392 (O_1392,N_19826,N_18711);
or UO_1393 (O_1393,N_18581,N_18822);
xnor UO_1394 (O_1394,N_19502,N_19386);
or UO_1395 (O_1395,N_18834,N_18277);
nand UO_1396 (O_1396,N_19198,N_19738);
or UO_1397 (O_1397,N_19014,N_18675);
and UO_1398 (O_1398,N_18216,N_18944);
or UO_1399 (O_1399,N_19680,N_19622);
nand UO_1400 (O_1400,N_19816,N_18160);
nor UO_1401 (O_1401,N_18882,N_19286);
xnor UO_1402 (O_1402,N_19393,N_19570);
and UO_1403 (O_1403,N_19930,N_19612);
xor UO_1404 (O_1404,N_19342,N_19154);
nor UO_1405 (O_1405,N_19356,N_19468);
nand UO_1406 (O_1406,N_18995,N_18330);
or UO_1407 (O_1407,N_19777,N_18211);
xor UO_1408 (O_1408,N_18246,N_18541);
or UO_1409 (O_1409,N_18669,N_18201);
or UO_1410 (O_1410,N_19443,N_18831);
and UO_1411 (O_1411,N_19891,N_18460);
xnor UO_1412 (O_1412,N_19261,N_19417);
nor UO_1413 (O_1413,N_18929,N_19993);
nand UO_1414 (O_1414,N_19468,N_18916);
nor UO_1415 (O_1415,N_19971,N_19383);
xnor UO_1416 (O_1416,N_19372,N_18802);
or UO_1417 (O_1417,N_19171,N_19654);
xnor UO_1418 (O_1418,N_19877,N_19350);
nor UO_1419 (O_1419,N_18355,N_18802);
nand UO_1420 (O_1420,N_18266,N_19666);
and UO_1421 (O_1421,N_18983,N_19704);
nand UO_1422 (O_1422,N_19406,N_18494);
nand UO_1423 (O_1423,N_19239,N_18122);
and UO_1424 (O_1424,N_18076,N_18024);
nand UO_1425 (O_1425,N_19501,N_19263);
xor UO_1426 (O_1426,N_18103,N_18122);
and UO_1427 (O_1427,N_18136,N_18137);
and UO_1428 (O_1428,N_19747,N_19009);
xor UO_1429 (O_1429,N_19027,N_19270);
xnor UO_1430 (O_1430,N_18437,N_19002);
nor UO_1431 (O_1431,N_18223,N_18673);
xor UO_1432 (O_1432,N_18531,N_19778);
nand UO_1433 (O_1433,N_18412,N_19080);
or UO_1434 (O_1434,N_18783,N_18224);
and UO_1435 (O_1435,N_19053,N_18410);
nand UO_1436 (O_1436,N_18065,N_18915);
xnor UO_1437 (O_1437,N_19770,N_19087);
nand UO_1438 (O_1438,N_19227,N_19104);
nand UO_1439 (O_1439,N_19116,N_18877);
nor UO_1440 (O_1440,N_19724,N_19986);
xnor UO_1441 (O_1441,N_19651,N_18872);
and UO_1442 (O_1442,N_19871,N_19759);
and UO_1443 (O_1443,N_18221,N_19753);
nand UO_1444 (O_1444,N_18943,N_19879);
or UO_1445 (O_1445,N_18528,N_18970);
nand UO_1446 (O_1446,N_18732,N_19043);
xnor UO_1447 (O_1447,N_18713,N_18129);
nor UO_1448 (O_1448,N_18510,N_19942);
or UO_1449 (O_1449,N_18932,N_19073);
and UO_1450 (O_1450,N_19447,N_18291);
nor UO_1451 (O_1451,N_19349,N_19008);
and UO_1452 (O_1452,N_18269,N_18230);
or UO_1453 (O_1453,N_18971,N_18734);
xor UO_1454 (O_1454,N_19671,N_18082);
nor UO_1455 (O_1455,N_18397,N_18231);
or UO_1456 (O_1456,N_18830,N_18996);
or UO_1457 (O_1457,N_18025,N_19646);
or UO_1458 (O_1458,N_19663,N_19670);
nor UO_1459 (O_1459,N_18606,N_18422);
or UO_1460 (O_1460,N_18170,N_18617);
nor UO_1461 (O_1461,N_18498,N_18030);
and UO_1462 (O_1462,N_18387,N_18213);
xor UO_1463 (O_1463,N_18325,N_18708);
nand UO_1464 (O_1464,N_18618,N_18262);
and UO_1465 (O_1465,N_18035,N_19358);
nor UO_1466 (O_1466,N_19884,N_18204);
nor UO_1467 (O_1467,N_19360,N_19013);
or UO_1468 (O_1468,N_19566,N_18211);
or UO_1469 (O_1469,N_18180,N_19788);
nor UO_1470 (O_1470,N_19143,N_18959);
or UO_1471 (O_1471,N_19389,N_18199);
or UO_1472 (O_1472,N_18175,N_18157);
nor UO_1473 (O_1473,N_18140,N_18539);
nor UO_1474 (O_1474,N_18183,N_19470);
and UO_1475 (O_1475,N_19705,N_18259);
nand UO_1476 (O_1476,N_19128,N_18746);
nand UO_1477 (O_1477,N_18220,N_19480);
and UO_1478 (O_1478,N_18168,N_18301);
nand UO_1479 (O_1479,N_19623,N_19646);
nor UO_1480 (O_1480,N_19109,N_19261);
and UO_1481 (O_1481,N_18235,N_19485);
nor UO_1482 (O_1482,N_18864,N_18569);
xor UO_1483 (O_1483,N_19414,N_18628);
nor UO_1484 (O_1484,N_19223,N_19729);
xnor UO_1485 (O_1485,N_18566,N_19781);
xnor UO_1486 (O_1486,N_18373,N_19509);
nor UO_1487 (O_1487,N_18792,N_19116);
nand UO_1488 (O_1488,N_18126,N_19400);
nor UO_1489 (O_1489,N_19586,N_18786);
xor UO_1490 (O_1490,N_19519,N_19824);
or UO_1491 (O_1491,N_18741,N_19816);
and UO_1492 (O_1492,N_19732,N_18095);
xor UO_1493 (O_1493,N_19370,N_18089);
xor UO_1494 (O_1494,N_19864,N_18285);
xnor UO_1495 (O_1495,N_18999,N_19048);
nand UO_1496 (O_1496,N_19040,N_18793);
or UO_1497 (O_1497,N_18228,N_18954);
nor UO_1498 (O_1498,N_19214,N_18586);
nor UO_1499 (O_1499,N_18371,N_19708);
or UO_1500 (O_1500,N_19511,N_19365);
or UO_1501 (O_1501,N_18796,N_18799);
nand UO_1502 (O_1502,N_19505,N_18972);
xor UO_1503 (O_1503,N_19452,N_19497);
xor UO_1504 (O_1504,N_19920,N_18615);
nor UO_1505 (O_1505,N_19446,N_19919);
nor UO_1506 (O_1506,N_18547,N_18497);
and UO_1507 (O_1507,N_19246,N_18366);
and UO_1508 (O_1508,N_18342,N_19743);
xor UO_1509 (O_1509,N_18638,N_18456);
and UO_1510 (O_1510,N_18194,N_19409);
and UO_1511 (O_1511,N_19906,N_19609);
nor UO_1512 (O_1512,N_18717,N_19998);
and UO_1513 (O_1513,N_18591,N_19654);
nand UO_1514 (O_1514,N_18989,N_18900);
or UO_1515 (O_1515,N_18073,N_19190);
nor UO_1516 (O_1516,N_19083,N_19609);
xor UO_1517 (O_1517,N_19406,N_18905);
nand UO_1518 (O_1518,N_19483,N_18117);
xnor UO_1519 (O_1519,N_19572,N_19856);
nand UO_1520 (O_1520,N_18441,N_19153);
nor UO_1521 (O_1521,N_18597,N_18985);
nor UO_1522 (O_1522,N_19602,N_18912);
and UO_1523 (O_1523,N_18019,N_18552);
and UO_1524 (O_1524,N_18221,N_18909);
xnor UO_1525 (O_1525,N_18157,N_18160);
nor UO_1526 (O_1526,N_19206,N_19740);
nor UO_1527 (O_1527,N_19376,N_18804);
xor UO_1528 (O_1528,N_19278,N_18109);
xnor UO_1529 (O_1529,N_18937,N_19886);
or UO_1530 (O_1530,N_18424,N_19800);
nor UO_1531 (O_1531,N_18959,N_18476);
xnor UO_1532 (O_1532,N_19812,N_18850);
xor UO_1533 (O_1533,N_18970,N_18688);
xor UO_1534 (O_1534,N_18311,N_18316);
xor UO_1535 (O_1535,N_19789,N_18210);
or UO_1536 (O_1536,N_18855,N_18426);
nand UO_1537 (O_1537,N_19885,N_19609);
nand UO_1538 (O_1538,N_19813,N_18785);
or UO_1539 (O_1539,N_19740,N_19068);
nor UO_1540 (O_1540,N_18112,N_18932);
xnor UO_1541 (O_1541,N_19505,N_18516);
nor UO_1542 (O_1542,N_18103,N_19125);
nand UO_1543 (O_1543,N_18314,N_19175);
or UO_1544 (O_1544,N_18190,N_19147);
and UO_1545 (O_1545,N_19392,N_18935);
or UO_1546 (O_1546,N_19812,N_18757);
and UO_1547 (O_1547,N_19620,N_18774);
nor UO_1548 (O_1548,N_19939,N_18649);
or UO_1549 (O_1549,N_18586,N_19195);
or UO_1550 (O_1550,N_18967,N_19955);
and UO_1551 (O_1551,N_19091,N_19332);
nor UO_1552 (O_1552,N_19268,N_19207);
and UO_1553 (O_1553,N_18566,N_19446);
nand UO_1554 (O_1554,N_18670,N_18053);
or UO_1555 (O_1555,N_18128,N_19033);
xor UO_1556 (O_1556,N_18497,N_19921);
and UO_1557 (O_1557,N_19660,N_19805);
xnor UO_1558 (O_1558,N_19873,N_18865);
xor UO_1559 (O_1559,N_18033,N_19918);
nor UO_1560 (O_1560,N_18335,N_18455);
xnor UO_1561 (O_1561,N_18632,N_19374);
or UO_1562 (O_1562,N_19271,N_18970);
or UO_1563 (O_1563,N_19487,N_18499);
and UO_1564 (O_1564,N_18458,N_19222);
nor UO_1565 (O_1565,N_19852,N_18853);
or UO_1566 (O_1566,N_19204,N_19173);
and UO_1567 (O_1567,N_18219,N_18290);
or UO_1568 (O_1568,N_19572,N_19888);
and UO_1569 (O_1569,N_18355,N_19277);
nor UO_1570 (O_1570,N_18887,N_18738);
xor UO_1571 (O_1571,N_18773,N_19597);
xor UO_1572 (O_1572,N_19117,N_19105);
nand UO_1573 (O_1573,N_18618,N_19959);
nor UO_1574 (O_1574,N_19725,N_19589);
xnor UO_1575 (O_1575,N_19013,N_18864);
or UO_1576 (O_1576,N_19488,N_18429);
and UO_1577 (O_1577,N_19389,N_18347);
nor UO_1578 (O_1578,N_18609,N_18856);
xnor UO_1579 (O_1579,N_18438,N_18552);
nand UO_1580 (O_1580,N_19361,N_18073);
nor UO_1581 (O_1581,N_18349,N_18655);
and UO_1582 (O_1582,N_19326,N_18771);
or UO_1583 (O_1583,N_19656,N_18945);
and UO_1584 (O_1584,N_19274,N_18394);
nor UO_1585 (O_1585,N_19577,N_18893);
nand UO_1586 (O_1586,N_19669,N_19470);
xor UO_1587 (O_1587,N_18141,N_19552);
or UO_1588 (O_1588,N_18827,N_19946);
nand UO_1589 (O_1589,N_18576,N_18966);
nor UO_1590 (O_1590,N_18369,N_18070);
or UO_1591 (O_1591,N_18114,N_19127);
xnor UO_1592 (O_1592,N_19143,N_18525);
nor UO_1593 (O_1593,N_19393,N_19705);
or UO_1594 (O_1594,N_18926,N_19654);
xor UO_1595 (O_1595,N_19581,N_19060);
and UO_1596 (O_1596,N_19311,N_18720);
nor UO_1597 (O_1597,N_18139,N_18897);
and UO_1598 (O_1598,N_19800,N_18397);
nor UO_1599 (O_1599,N_19119,N_18084);
xor UO_1600 (O_1600,N_18052,N_18130);
xnor UO_1601 (O_1601,N_19777,N_18204);
nor UO_1602 (O_1602,N_19479,N_18353);
or UO_1603 (O_1603,N_18490,N_18449);
xnor UO_1604 (O_1604,N_19040,N_19497);
xnor UO_1605 (O_1605,N_18879,N_18194);
or UO_1606 (O_1606,N_18968,N_18838);
nand UO_1607 (O_1607,N_19000,N_19313);
or UO_1608 (O_1608,N_19368,N_18011);
xnor UO_1609 (O_1609,N_18124,N_19127);
nand UO_1610 (O_1610,N_19811,N_18187);
and UO_1611 (O_1611,N_19082,N_19276);
or UO_1612 (O_1612,N_19831,N_18509);
xor UO_1613 (O_1613,N_19402,N_19322);
nor UO_1614 (O_1614,N_19541,N_19308);
or UO_1615 (O_1615,N_18003,N_18142);
xnor UO_1616 (O_1616,N_18769,N_19084);
and UO_1617 (O_1617,N_19094,N_19865);
and UO_1618 (O_1618,N_18934,N_18718);
nor UO_1619 (O_1619,N_19770,N_19619);
xor UO_1620 (O_1620,N_18310,N_18369);
nor UO_1621 (O_1621,N_18862,N_18865);
and UO_1622 (O_1622,N_19746,N_18842);
xor UO_1623 (O_1623,N_19423,N_18896);
xor UO_1624 (O_1624,N_18581,N_18311);
or UO_1625 (O_1625,N_19335,N_18626);
nand UO_1626 (O_1626,N_19594,N_18458);
xor UO_1627 (O_1627,N_18396,N_19499);
and UO_1628 (O_1628,N_18424,N_18529);
and UO_1629 (O_1629,N_18719,N_19760);
or UO_1630 (O_1630,N_19605,N_19850);
and UO_1631 (O_1631,N_19326,N_18890);
and UO_1632 (O_1632,N_18933,N_18389);
xnor UO_1633 (O_1633,N_18877,N_19281);
or UO_1634 (O_1634,N_18049,N_18703);
nand UO_1635 (O_1635,N_19560,N_18777);
nand UO_1636 (O_1636,N_19916,N_19260);
and UO_1637 (O_1637,N_18428,N_19614);
or UO_1638 (O_1638,N_18116,N_19605);
nor UO_1639 (O_1639,N_18012,N_19081);
nor UO_1640 (O_1640,N_19302,N_18748);
xor UO_1641 (O_1641,N_19856,N_19264);
nand UO_1642 (O_1642,N_18168,N_18668);
or UO_1643 (O_1643,N_18997,N_18935);
nand UO_1644 (O_1644,N_19124,N_18722);
and UO_1645 (O_1645,N_18574,N_18098);
and UO_1646 (O_1646,N_18204,N_18075);
nand UO_1647 (O_1647,N_19257,N_19763);
xor UO_1648 (O_1648,N_19515,N_19572);
nand UO_1649 (O_1649,N_19414,N_19005);
nand UO_1650 (O_1650,N_18390,N_19396);
nand UO_1651 (O_1651,N_19222,N_19601);
nand UO_1652 (O_1652,N_19776,N_19696);
xnor UO_1653 (O_1653,N_18236,N_19117);
or UO_1654 (O_1654,N_18091,N_19100);
xor UO_1655 (O_1655,N_18056,N_19011);
or UO_1656 (O_1656,N_18319,N_19206);
xor UO_1657 (O_1657,N_19376,N_18323);
nand UO_1658 (O_1658,N_19207,N_19894);
nand UO_1659 (O_1659,N_18410,N_19844);
nand UO_1660 (O_1660,N_19348,N_18393);
and UO_1661 (O_1661,N_18988,N_18214);
nand UO_1662 (O_1662,N_18549,N_18479);
and UO_1663 (O_1663,N_18483,N_18438);
nor UO_1664 (O_1664,N_19402,N_19771);
nand UO_1665 (O_1665,N_19572,N_19945);
xor UO_1666 (O_1666,N_19784,N_18555);
or UO_1667 (O_1667,N_19252,N_19296);
xnor UO_1668 (O_1668,N_19202,N_19028);
nor UO_1669 (O_1669,N_18861,N_18412);
nand UO_1670 (O_1670,N_19614,N_19490);
nand UO_1671 (O_1671,N_19287,N_18367);
nand UO_1672 (O_1672,N_18334,N_19578);
or UO_1673 (O_1673,N_18027,N_18044);
nor UO_1674 (O_1674,N_19035,N_19217);
or UO_1675 (O_1675,N_19202,N_18523);
or UO_1676 (O_1676,N_19299,N_18800);
nor UO_1677 (O_1677,N_19480,N_19976);
and UO_1678 (O_1678,N_19222,N_19830);
and UO_1679 (O_1679,N_18470,N_18508);
xor UO_1680 (O_1680,N_19358,N_19411);
nor UO_1681 (O_1681,N_19681,N_18713);
nor UO_1682 (O_1682,N_19520,N_19935);
xnor UO_1683 (O_1683,N_19905,N_19030);
nand UO_1684 (O_1684,N_19874,N_19213);
and UO_1685 (O_1685,N_19198,N_18835);
or UO_1686 (O_1686,N_19691,N_18926);
nor UO_1687 (O_1687,N_18562,N_19030);
nand UO_1688 (O_1688,N_18224,N_18438);
xor UO_1689 (O_1689,N_18491,N_19401);
and UO_1690 (O_1690,N_18501,N_19316);
nor UO_1691 (O_1691,N_18708,N_18350);
or UO_1692 (O_1692,N_19686,N_19067);
and UO_1693 (O_1693,N_19749,N_18948);
or UO_1694 (O_1694,N_19806,N_18387);
xnor UO_1695 (O_1695,N_18589,N_19270);
or UO_1696 (O_1696,N_19656,N_19424);
xnor UO_1697 (O_1697,N_19052,N_18861);
and UO_1698 (O_1698,N_19441,N_18039);
nor UO_1699 (O_1699,N_19458,N_19396);
or UO_1700 (O_1700,N_19115,N_18534);
and UO_1701 (O_1701,N_19938,N_18828);
or UO_1702 (O_1702,N_18042,N_18581);
or UO_1703 (O_1703,N_19970,N_19507);
or UO_1704 (O_1704,N_18063,N_19165);
or UO_1705 (O_1705,N_19219,N_18416);
nand UO_1706 (O_1706,N_18077,N_19032);
and UO_1707 (O_1707,N_19539,N_18844);
and UO_1708 (O_1708,N_19076,N_18020);
xor UO_1709 (O_1709,N_19933,N_19476);
and UO_1710 (O_1710,N_19567,N_19538);
xor UO_1711 (O_1711,N_19233,N_18388);
nand UO_1712 (O_1712,N_18872,N_18504);
xnor UO_1713 (O_1713,N_18615,N_18241);
nand UO_1714 (O_1714,N_18379,N_19582);
and UO_1715 (O_1715,N_19924,N_19257);
nor UO_1716 (O_1716,N_18683,N_18642);
xnor UO_1717 (O_1717,N_19573,N_19614);
and UO_1718 (O_1718,N_19649,N_19362);
xor UO_1719 (O_1719,N_19929,N_18792);
or UO_1720 (O_1720,N_19814,N_19243);
and UO_1721 (O_1721,N_18135,N_18046);
xor UO_1722 (O_1722,N_18439,N_19754);
or UO_1723 (O_1723,N_18898,N_19697);
nor UO_1724 (O_1724,N_19622,N_18913);
xnor UO_1725 (O_1725,N_18832,N_19779);
xnor UO_1726 (O_1726,N_18470,N_19035);
and UO_1727 (O_1727,N_18419,N_18666);
nand UO_1728 (O_1728,N_19628,N_19694);
xor UO_1729 (O_1729,N_19776,N_19576);
or UO_1730 (O_1730,N_19082,N_19334);
nor UO_1731 (O_1731,N_19444,N_18309);
nor UO_1732 (O_1732,N_19194,N_18566);
xor UO_1733 (O_1733,N_19706,N_18434);
and UO_1734 (O_1734,N_18360,N_19734);
nand UO_1735 (O_1735,N_19863,N_18902);
nand UO_1736 (O_1736,N_19718,N_19539);
and UO_1737 (O_1737,N_19678,N_19305);
nor UO_1738 (O_1738,N_19587,N_18555);
nor UO_1739 (O_1739,N_19277,N_19002);
and UO_1740 (O_1740,N_18675,N_18366);
nor UO_1741 (O_1741,N_18236,N_18954);
nand UO_1742 (O_1742,N_18657,N_18764);
nand UO_1743 (O_1743,N_19306,N_19088);
and UO_1744 (O_1744,N_19341,N_19488);
or UO_1745 (O_1745,N_18623,N_19313);
xor UO_1746 (O_1746,N_19116,N_19862);
nand UO_1747 (O_1747,N_18758,N_18988);
nand UO_1748 (O_1748,N_18623,N_19767);
nor UO_1749 (O_1749,N_19979,N_19198);
or UO_1750 (O_1750,N_18239,N_18244);
or UO_1751 (O_1751,N_19248,N_18156);
xnor UO_1752 (O_1752,N_19179,N_19659);
and UO_1753 (O_1753,N_18620,N_18469);
and UO_1754 (O_1754,N_19699,N_18791);
nor UO_1755 (O_1755,N_19160,N_18592);
nand UO_1756 (O_1756,N_19237,N_18774);
or UO_1757 (O_1757,N_18479,N_19507);
or UO_1758 (O_1758,N_19486,N_18027);
and UO_1759 (O_1759,N_19916,N_19055);
nor UO_1760 (O_1760,N_18535,N_18870);
or UO_1761 (O_1761,N_19096,N_18926);
xor UO_1762 (O_1762,N_19247,N_18293);
nor UO_1763 (O_1763,N_19563,N_19052);
and UO_1764 (O_1764,N_19572,N_18452);
or UO_1765 (O_1765,N_19355,N_18074);
xor UO_1766 (O_1766,N_18090,N_19688);
and UO_1767 (O_1767,N_19209,N_18072);
nand UO_1768 (O_1768,N_19426,N_19440);
nor UO_1769 (O_1769,N_19512,N_18167);
and UO_1770 (O_1770,N_19864,N_18035);
nor UO_1771 (O_1771,N_18669,N_18301);
and UO_1772 (O_1772,N_19346,N_19453);
and UO_1773 (O_1773,N_19357,N_19451);
and UO_1774 (O_1774,N_18043,N_18649);
or UO_1775 (O_1775,N_19075,N_18302);
xnor UO_1776 (O_1776,N_19256,N_18472);
or UO_1777 (O_1777,N_19100,N_18796);
and UO_1778 (O_1778,N_18174,N_18263);
nand UO_1779 (O_1779,N_18302,N_18365);
or UO_1780 (O_1780,N_18375,N_19076);
nand UO_1781 (O_1781,N_18490,N_19385);
or UO_1782 (O_1782,N_19232,N_19648);
or UO_1783 (O_1783,N_19604,N_18083);
nor UO_1784 (O_1784,N_18833,N_19049);
and UO_1785 (O_1785,N_19972,N_18913);
or UO_1786 (O_1786,N_19428,N_19953);
or UO_1787 (O_1787,N_19260,N_19685);
xor UO_1788 (O_1788,N_19300,N_18839);
nor UO_1789 (O_1789,N_19068,N_18411);
nor UO_1790 (O_1790,N_19765,N_18269);
and UO_1791 (O_1791,N_19699,N_18276);
xor UO_1792 (O_1792,N_19210,N_18628);
nand UO_1793 (O_1793,N_19488,N_19974);
nand UO_1794 (O_1794,N_18375,N_18089);
xor UO_1795 (O_1795,N_19863,N_18186);
nor UO_1796 (O_1796,N_19359,N_18591);
and UO_1797 (O_1797,N_18562,N_19609);
and UO_1798 (O_1798,N_18877,N_18422);
xnor UO_1799 (O_1799,N_19246,N_19557);
nand UO_1800 (O_1800,N_19628,N_19473);
nor UO_1801 (O_1801,N_18998,N_18434);
or UO_1802 (O_1802,N_18311,N_18850);
nor UO_1803 (O_1803,N_19892,N_19555);
or UO_1804 (O_1804,N_19266,N_18878);
nand UO_1805 (O_1805,N_18441,N_19868);
or UO_1806 (O_1806,N_19448,N_18317);
and UO_1807 (O_1807,N_18549,N_19727);
nor UO_1808 (O_1808,N_18346,N_18337);
xnor UO_1809 (O_1809,N_18080,N_19497);
or UO_1810 (O_1810,N_18733,N_19531);
and UO_1811 (O_1811,N_19583,N_19277);
and UO_1812 (O_1812,N_18396,N_19537);
and UO_1813 (O_1813,N_19679,N_18706);
and UO_1814 (O_1814,N_18783,N_18833);
nor UO_1815 (O_1815,N_19683,N_18861);
xnor UO_1816 (O_1816,N_19828,N_18993);
and UO_1817 (O_1817,N_18706,N_19667);
and UO_1818 (O_1818,N_19444,N_18576);
and UO_1819 (O_1819,N_18574,N_19953);
nand UO_1820 (O_1820,N_18701,N_18984);
or UO_1821 (O_1821,N_18536,N_19364);
or UO_1822 (O_1822,N_19922,N_18858);
or UO_1823 (O_1823,N_19526,N_19633);
and UO_1824 (O_1824,N_19352,N_19543);
or UO_1825 (O_1825,N_19428,N_19746);
xor UO_1826 (O_1826,N_18625,N_18342);
or UO_1827 (O_1827,N_18378,N_19194);
and UO_1828 (O_1828,N_19044,N_19403);
and UO_1829 (O_1829,N_18631,N_18463);
xor UO_1830 (O_1830,N_18321,N_19883);
nand UO_1831 (O_1831,N_19357,N_18026);
or UO_1832 (O_1832,N_19955,N_19126);
and UO_1833 (O_1833,N_19007,N_18373);
or UO_1834 (O_1834,N_18775,N_19951);
and UO_1835 (O_1835,N_19130,N_18481);
or UO_1836 (O_1836,N_19839,N_19214);
nor UO_1837 (O_1837,N_18782,N_18742);
nand UO_1838 (O_1838,N_19409,N_18160);
nor UO_1839 (O_1839,N_18226,N_18734);
and UO_1840 (O_1840,N_19851,N_19765);
nor UO_1841 (O_1841,N_19834,N_19369);
nor UO_1842 (O_1842,N_18877,N_19667);
xor UO_1843 (O_1843,N_18765,N_18328);
and UO_1844 (O_1844,N_18089,N_18129);
and UO_1845 (O_1845,N_18981,N_19720);
and UO_1846 (O_1846,N_18918,N_19445);
xnor UO_1847 (O_1847,N_19517,N_18777);
or UO_1848 (O_1848,N_19225,N_18709);
nand UO_1849 (O_1849,N_18071,N_18572);
nor UO_1850 (O_1850,N_18849,N_18556);
and UO_1851 (O_1851,N_18551,N_18827);
nand UO_1852 (O_1852,N_19814,N_19712);
nand UO_1853 (O_1853,N_18820,N_18101);
nor UO_1854 (O_1854,N_19151,N_18403);
nand UO_1855 (O_1855,N_19286,N_19262);
nand UO_1856 (O_1856,N_19457,N_19315);
nor UO_1857 (O_1857,N_19913,N_19436);
nor UO_1858 (O_1858,N_19788,N_18693);
nand UO_1859 (O_1859,N_18048,N_19819);
and UO_1860 (O_1860,N_18090,N_19234);
nor UO_1861 (O_1861,N_19102,N_19003);
nand UO_1862 (O_1862,N_19172,N_18158);
or UO_1863 (O_1863,N_18028,N_19972);
nand UO_1864 (O_1864,N_19731,N_19267);
and UO_1865 (O_1865,N_18252,N_19245);
nor UO_1866 (O_1866,N_18816,N_19434);
xnor UO_1867 (O_1867,N_18908,N_18843);
or UO_1868 (O_1868,N_19245,N_19243);
xnor UO_1869 (O_1869,N_19815,N_19599);
nand UO_1870 (O_1870,N_19962,N_19980);
xnor UO_1871 (O_1871,N_19716,N_19212);
and UO_1872 (O_1872,N_18644,N_19479);
xor UO_1873 (O_1873,N_19830,N_19633);
nand UO_1874 (O_1874,N_18967,N_19088);
nor UO_1875 (O_1875,N_19029,N_19323);
and UO_1876 (O_1876,N_19856,N_18360);
and UO_1877 (O_1877,N_19597,N_19990);
or UO_1878 (O_1878,N_18031,N_18056);
xnor UO_1879 (O_1879,N_18723,N_18860);
xnor UO_1880 (O_1880,N_19378,N_18211);
nor UO_1881 (O_1881,N_18191,N_18697);
nor UO_1882 (O_1882,N_19517,N_18873);
nand UO_1883 (O_1883,N_18243,N_18653);
or UO_1884 (O_1884,N_18315,N_19591);
nor UO_1885 (O_1885,N_18078,N_19915);
xor UO_1886 (O_1886,N_18176,N_19441);
xor UO_1887 (O_1887,N_18969,N_19251);
or UO_1888 (O_1888,N_18405,N_18046);
or UO_1889 (O_1889,N_18718,N_19766);
and UO_1890 (O_1890,N_19717,N_18362);
nor UO_1891 (O_1891,N_18491,N_18884);
nor UO_1892 (O_1892,N_19582,N_18510);
xnor UO_1893 (O_1893,N_19771,N_19523);
or UO_1894 (O_1894,N_19209,N_18016);
nor UO_1895 (O_1895,N_18600,N_19377);
nor UO_1896 (O_1896,N_19883,N_19600);
nand UO_1897 (O_1897,N_19725,N_19480);
xor UO_1898 (O_1898,N_19339,N_18021);
nor UO_1899 (O_1899,N_19949,N_19543);
nor UO_1900 (O_1900,N_19209,N_18544);
or UO_1901 (O_1901,N_18364,N_19085);
nand UO_1902 (O_1902,N_19432,N_19099);
and UO_1903 (O_1903,N_19082,N_19866);
xor UO_1904 (O_1904,N_18827,N_19134);
nand UO_1905 (O_1905,N_18382,N_18236);
or UO_1906 (O_1906,N_18033,N_19333);
and UO_1907 (O_1907,N_18171,N_19059);
and UO_1908 (O_1908,N_19972,N_18064);
nor UO_1909 (O_1909,N_18244,N_19854);
xor UO_1910 (O_1910,N_19196,N_18425);
nor UO_1911 (O_1911,N_19693,N_19476);
nand UO_1912 (O_1912,N_18928,N_19716);
xor UO_1913 (O_1913,N_19446,N_19821);
and UO_1914 (O_1914,N_19823,N_19305);
nor UO_1915 (O_1915,N_18359,N_19807);
nand UO_1916 (O_1916,N_19145,N_18055);
nand UO_1917 (O_1917,N_19531,N_19344);
xor UO_1918 (O_1918,N_19466,N_18573);
nand UO_1919 (O_1919,N_18095,N_18594);
nor UO_1920 (O_1920,N_18441,N_18495);
or UO_1921 (O_1921,N_19836,N_18257);
xor UO_1922 (O_1922,N_19382,N_18052);
nand UO_1923 (O_1923,N_18055,N_18532);
or UO_1924 (O_1924,N_19006,N_18885);
and UO_1925 (O_1925,N_19454,N_19055);
or UO_1926 (O_1926,N_18703,N_19857);
or UO_1927 (O_1927,N_19956,N_18203);
xnor UO_1928 (O_1928,N_18207,N_19175);
nand UO_1929 (O_1929,N_18683,N_18672);
nor UO_1930 (O_1930,N_19936,N_19968);
and UO_1931 (O_1931,N_18987,N_19927);
and UO_1932 (O_1932,N_18560,N_19403);
nand UO_1933 (O_1933,N_18987,N_19776);
and UO_1934 (O_1934,N_19897,N_18051);
or UO_1935 (O_1935,N_19765,N_18634);
or UO_1936 (O_1936,N_18474,N_19179);
and UO_1937 (O_1937,N_18312,N_18146);
and UO_1938 (O_1938,N_18726,N_19726);
xnor UO_1939 (O_1939,N_18368,N_18402);
nand UO_1940 (O_1940,N_19183,N_18623);
nor UO_1941 (O_1941,N_19649,N_18524);
and UO_1942 (O_1942,N_18504,N_18848);
nor UO_1943 (O_1943,N_18860,N_19156);
or UO_1944 (O_1944,N_19400,N_19977);
or UO_1945 (O_1945,N_19329,N_18844);
xor UO_1946 (O_1946,N_19712,N_18313);
and UO_1947 (O_1947,N_18018,N_19747);
nor UO_1948 (O_1948,N_19202,N_18032);
nor UO_1949 (O_1949,N_19157,N_19156);
or UO_1950 (O_1950,N_18944,N_18443);
nand UO_1951 (O_1951,N_19193,N_18607);
or UO_1952 (O_1952,N_18579,N_18596);
nor UO_1953 (O_1953,N_18743,N_18374);
and UO_1954 (O_1954,N_19923,N_18316);
xor UO_1955 (O_1955,N_18728,N_18415);
nand UO_1956 (O_1956,N_18775,N_18377);
and UO_1957 (O_1957,N_18396,N_19263);
or UO_1958 (O_1958,N_19909,N_18902);
and UO_1959 (O_1959,N_18343,N_19604);
nor UO_1960 (O_1960,N_19167,N_18587);
or UO_1961 (O_1961,N_19330,N_18229);
or UO_1962 (O_1962,N_18021,N_18344);
or UO_1963 (O_1963,N_19474,N_18898);
nand UO_1964 (O_1964,N_18772,N_18387);
or UO_1965 (O_1965,N_19002,N_18367);
xnor UO_1966 (O_1966,N_18241,N_18205);
xor UO_1967 (O_1967,N_18974,N_19824);
nand UO_1968 (O_1968,N_19059,N_19610);
nor UO_1969 (O_1969,N_19936,N_19064);
and UO_1970 (O_1970,N_19466,N_18571);
or UO_1971 (O_1971,N_18202,N_18925);
or UO_1972 (O_1972,N_19294,N_19966);
or UO_1973 (O_1973,N_19284,N_18859);
nand UO_1974 (O_1974,N_18015,N_18915);
nor UO_1975 (O_1975,N_19996,N_18957);
and UO_1976 (O_1976,N_19230,N_18317);
or UO_1977 (O_1977,N_19724,N_18536);
nand UO_1978 (O_1978,N_18509,N_18675);
nand UO_1979 (O_1979,N_18031,N_19569);
xor UO_1980 (O_1980,N_18963,N_18024);
nand UO_1981 (O_1981,N_19240,N_19308);
nor UO_1982 (O_1982,N_19031,N_18262);
or UO_1983 (O_1983,N_19567,N_19996);
nor UO_1984 (O_1984,N_19155,N_18844);
nor UO_1985 (O_1985,N_18354,N_19032);
nor UO_1986 (O_1986,N_19873,N_19958);
and UO_1987 (O_1987,N_19854,N_18547);
nor UO_1988 (O_1988,N_19004,N_19862);
and UO_1989 (O_1989,N_18713,N_19353);
nand UO_1990 (O_1990,N_18603,N_19042);
or UO_1991 (O_1991,N_19487,N_18789);
nand UO_1992 (O_1992,N_19042,N_18780);
nor UO_1993 (O_1993,N_19045,N_18867);
xnor UO_1994 (O_1994,N_18232,N_18957);
xor UO_1995 (O_1995,N_18111,N_18680);
xor UO_1996 (O_1996,N_18899,N_19683);
nand UO_1997 (O_1997,N_18756,N_18495);
xor UO_1998 (O_1998,N_19047,N_18875);
nor UO_1999 (O_1999,N_19575,N_18784);
xnor UO_2000 (O_2000,N_18939,N_18851);
xor UO_2001 (O_2001,N_18349,N_19536);
xnor UO_2002 (O_2002,N_18112,N_18263);
or UO_2003 (O_2003,N_19644,N_19258);
xor UO_2004 (O_2004,N_19375,N_18710);
or UO_2005 (O_2005,N_18796,N_19825);
or UO_2006 (O_2006,N_19976,N_18006);
nand UO_2007 (O_2007,N_18219,N_19847);
xnor UO_2008 (O_2008,N_18103,N_18318);
and UO_2009 (O_2009,N_18690,N_18453);
and UO_2010 (O_2010,N_19465,N_19828);
nor UO_2011 (O_2011,N_18903,N_19703);
nor UO_2012 (O_2012,N_18941,N_19235);
nand UO_2013 (O_2013,N_18022,N_19357);
xnor UO_2014 (O_2014,N_19091,N_18175);
nand UO_2015 (O_2015,N_18443,N_19665);
xnor UO_2016 (O_2016,N_18167,N_18185);
or UO_2017 (O_2017,N_19384,N_19230);
and UO_2018 (O_2018,N_18405,N_18782);
xnor UO_2019 (O_2019,N_19743,N_18362);
nor UO_2020 (O_2020,N_19879,N_18642);
nor UO_2021 (O_2021,N_19086,N_18370);
nand UO_2022 (O_2022,N_19812,N_18733);
and UO_2023 (O_2023,N_18933,N_19601);
or UO_2024 (O_2024,N_19523,N_19799);
xnor UO_2025 (O_2025,N_19455,N_19714);
nand UO_2026 (O_2026,N_19514,N_18785);
xnor UO_2027 (O_2027,N_18971,N_18764);
and UO_2028 (O_2028,N_18591,N_19475);
xnor UO_2029 (O_2029,N_18849,N_19528);
and UO_2030 (O_2030,N_19552,N_19220);
nand UO_2031 (O_2031,N_18216,N_18737);
nand UO_2032 (O_2032,N_18754,N_19234);
xor UO_2033 (O_2033,N_19945,N_19519);
nand UO_2034 (O_2034,N_19852,N_19001);
xnor UO_2035 (O_2035,N_19205,N_19380);
nand UO_2036 (O_2036,N_18251,N_18971);
xnor UO_2037 (O_2037,N_19745,N_19630);
and UO_2038 (O_2038,N_18967,N_19669);
and UO_2039 (O_2039,N_18699,N_19263);
or UO_2040 (O_2040,N_18917,N_18940);
or UO_2041 (O_2041,N_19773,N_18533);
or UO_2042 (O_2042,N_19522,N_19947);
nand UO_2043 (O_2043,N_19876,N_18019);
or UO_2044 (O_2044,N_19051,N_18667);
nor UO_2045 (O_2045,N_19248,N_18429);
and UO_2046 (O_2046,N_18531,N_19506);
or UO_2047 (O_2047,N_18748,N_19366);
and UO_2048 (O_2048,N_18176,N_19537);
nor UO_2049 (O_2049,N_18826,N_18722);
nor UO_2050 (O_2050,N_18087,N_19235);
xnor UO_2051 (O_2051,N_18480,N_19140);
xor UO_2052 (O_2052,N_18510,N_18813);
nor UO_2053 (O_2053,N_18942,N_19332);
nand UO_2054 (O_2054,N_18452,N_19472);
or UO_2055 (O_2055,N_18829,N_19973);
and UO_2056 (O_2056,N_18638,N_19573);
and UO_2057 (O_2057,N_19996,N_19081);
nor UO_2058 (O_2058,N_18918,N_18937);
nor UO_2059 (O_2059,N_19924,N_18635);
xnor UO_2060 (O_2060,N_18293,N_19716);
nor UO_2061 (O_2061,N_18127,N_18644);
xor UO_2062 (O_2062,N_18231,N_19039);
xor UO_2063 (O_2063,N_19454,N_18367);
nand UO_2064 (O_2064,N_18540,N_18535);
nand UO_2065 (O_2065,N_18800,N_18965);
xnor UO_2066 (O_2066,N_18946,N_18276);
or UO_2067 (O_2067,N_19905,N_18968);
xor UO_2068 (O_2068,N_19368,N_19759);
nor UO_2069 (O_2069,N_18079,N_19824);
nor UO_2070 (O_2070,N_19447,N_18944);
or UO_2071 (O_2071,N_19753,N_18754);
nand UO_2072 (O_2072,N_18744,N_18750);
xor UO_2073 (O_2073,N_18722,N_18213);
nor UO_2074 (O_2074,N_19985,N_19709);
and UO_2075 (O_2075,N_19579,N_19675);
or UO_2076 (O_2076,N_19507,N_18292);
nand UO_2077 (O_2077,N_18651,N_19861);
and UO_2078 (O_2078,N_18870,N_18097);
xor UO_2079 (O_2079,N_19964,N_19300);
nor UO_2080 (O_2080,N_18919,N_18384);
nand UO_2081 (O_2081,N_19816,N_18774);
or UO_2082 (O_2082,N_18024,N_19485);
or UO_2083 (O_2083,N_18063,N_19449);
nand UO_2084 (O_2084,N_18524,N_18643);
or UO_2085 (O_2085,N_18132,N_19513);
xnor UO_2086 (O_2086,N_19148,N_18720);
or UO_2087 (O_2087,N_18547,N_18417);
and UO_2088 (O_2088,N_18663,N_19183);
nand UO_2089 (O_2089,N_18212,N_19302);
and UO_2090 (O_2090,N_19913,N_19667);
nand UO_2091 (O_2091,N_19570,N_19206);
nand UO_2092 (O_2092,N_19031,N_19464);
and UO_2093 (O_2093,N_19302,N_18521);
xor UO_2094 (O_2094,N_18276,N_19484);
or UO_2095 (O_2095,N_18518,N_18626);
and UO_2096 (O_2096,N_18160,N_19709);
nand UO_2097 (O_2097,N_19823,N_18808);
or UO_2098 (O_2098,N_19950,N_18032);
or UO_2099 (O_2099,N_18084,N_18896);
xor UO_2100 (O_2100,N_18774,N_19381);
xor UO_2101 (O_2101,N_18000,N_18352);
and UO_2102 (O_2102,N_18970,N_19535);
and UO_2103 (O_2103,N_18534,N_18712);
nand UO_2104 (O_2104,N_19990,N_19989);
xnor UO_2105 (O_2105,N_19915,N_18119);
or UO_2106 (O_2106,N_19630,N_18815);
nor UO_2107 (O_2107,N_19554,N_19821);
xnor UO_2108 (O_2108,N_18904,N_19026);
and UO_2109 (O_2109,N_18979,N_18324);
and UO_2110 (O_2110,N_19286,N_18683);
xor UO_2111 (O_2111,N_18955,N_19075);
and UO_2112 (O_2112,N_19868,N_19173);
or UO_2113 (O_2113,N_18670,N_19387);
nor UO_2114 (O_2114,N_19588,N_19682);
nand UO_2115 (O_2115,N_19240,N_19152);
or UO_2116 (O_2116,N_19975,N_18880);
and UO_2117 (O_2117,N_19532,N_19512);
and UO_2118 (O_2118,N_18809,N_18153);
or UO_2119 (O_2119,N_18923,N_19907);
nand UO_2120 (O_2120,N_18474,N_18505);
and UO_2121 (O_2121,N_18497,N_19111);
xor UO_2122 (O_2122,N_19263,N_19735);
nand UO_2123 (O_2123,N_19632,N_19475);
nand UO_2124 (O_2124,N_18266,N_19882);
nor UO_2125 (O_2125,N_18161,N_18692);
or UO_2126 (O_2126,N_18966,N_19163);
and UO_2127 (O_2127,N_19625,N_18264);
nand UO_2128 (O_2128,N_19717,N_18882);
xor UO_2129 (O_2129,N_18741,N_19575);
nand UO_2130 (O_2130,N_19997,N_18250);
xnor UO_2131 (O_2131,N_18774,N_18600);
or UO_2132 (O_2132,N_18571,N_19276);
nor UO_2133 (O_2133,N_18316,N_18881);
or UO_2134 (O_2134,N_18465,N_18833);
xnor UO_2135 (O_2135,N_18347,N_18921);
nand UO_2136 (O_2136,N_19769,N_18081);
xnor UO_2137 (O_2137,N_18795,N_19885);
nor UO_2138 (O_2138,N_19774,N_18982);
nor UO_2139 (O_2139,N_18687,N_19220);
or UO_2140 (O_2140,N_18428,N_18980);
nand UO_2141 (O_2141,N_19851,N_18378);
xor UO_2142 (O_2142,N_19273,N_19434);
nand UO_2143 (O_2143,N_19485,N_19575);
and UO_2144 (O_2144,N_18143,N_18836);
nand UO_2145 (O_2145,N_19069,N_19976);
or UO_2146 (O_2146,N_19857,N_18299);
or UO_2147 (O_2147,N_19096,N_19574);
or UO_2148 (O_2148,N_18918,N_19973);
and UO_2149 (O_2149,N_19562,N_18842);
or UO_2150 (O_2150,N_18623,N_18489);
and UO_2151 (O_2151,N_18032,N_18379);
and UO_2152 (O_2152,N_18154,N_19875);
xor UO_2153 (O_2153,N_18375,N_18668);
nor UO_2154 (O_2154,N_19040,N_19767);
and UO_2155 (O_2155,N_19604,N_18295);
nand UO_2156 (O_2156,N_18901,N_18870);
xor UO_2157 (O_2157,N_19226,N_18831);
nor UO_2158 (O_2158,N_18183,N_19183);
or UO_2159 (O_2159,N_18659,N_18057);
or UO_2160 (O_2160,N_19566,N_19598);
or UO_2161 (O_2161,N_19646,N_19051);
nand UO_2162 (O_2162,N_19913,N_19400);
or UO_2163 (O_2163,N_19556,N_18830);
xor UO_2164 (O_2164,N_19838,N_19758);
nor UO_2165 (O_2165,N_19399,N_19435);
and UO_2166 (O_2166,N_18700,N_18028);
xor UO_2167 (O_2167,N_19848,N_18760);
nor UO_2168 (O_2168,N_18212,N_19055);
nand UO_2169 (O_2169,N_18609,N_19096);
nand UO_2170 (O_2170,N_19690,N_18624);
or UO_2171 (O_2171,N_18198,N_19418);
xor UO_2172 (O_2172,N_19095,N_19740);
nand UO_2173 (O_2173,N_18667,N_18565);
xnor UO_2174 (O_2174,N_19116,N_19647);
and UO_2175 (O_2175,N_19087,N_19842);
nand UO_2176 (O_2176,N_18213,N_19284);
xnor UO_2177 (O_2177,N_18365,N_18479);
nand UO_2178 (O_2178,N_18757,N_19803);
xor UO_2179 (O_2179,N_18616,N_19405);
nor UO_2180 (O_2180,N_18244,N_18578);
nand UO_2181 (O_2181,N_18869,N_19615);
and UO_2182 (O_2182,N_18506,N_19902);
xnor UO_2183 (O_2183,N_19218,N_18453);
and UO_2184 (O_2184,N_18301,N_18964);
xnor UO_2185 (O_2185,N_18375,N_18453);
nand UO_2186 (O_2186,N_18344,N_18147);
and UO_2187 (O_2187,N_18741,N_18956);
nand UO_2188 (O_2188,N_19011,N_18161);
xnor UO_2189 (O_2189,N_19820,N_19845);
and UO_2190 (O_2190,N_19703,N_19964);
xor UO_2191 (O_2191,N_18213,N_18711);
nand UO_2192 (O_2192,N_19880,N_18550);
and UO_2193 (O_2193,N_18305,N_18580);
nor UO_2194 (O_2194,N_19012,N_18550);
or UO_2195 (O_2195,N_18992,N_18122);
or UO_2196 (O_2196,N_19167,N_19268);
nand UO_2197 (O_2197,N_19532,N_18005);
nand UO_2198 (O_2198,N_18095,N_18795);
nand UO_2199 (O_2199,N_19100,N_18570);
xor UO_2200 (O_2200,N_19267,N_18759);
xnor UO_2201 (O_2201,N_18955,N_19082);
nor UO_2202 (O_2202,N_18961,N_18797);
or UO_2203 (O_2203,N_18434,N_19337);
nand UO_2204 (O_2204,N_19819,N_18926);
and UO_2205 (O_2205,N_19132,N_19077);
xnor UO_2206 (O_2206,N_18040,N_18185);
nor UO_2207 (O_2207,N_18435,N_18175);
nand UO_2208 (O_2208,N_18018,N_19151);
nor UO_2209 (O_2209,N_19127,N_19659);
and UO_2210 (O_2210,N_18733,N_18696);
nand UO_2211 (O_2211,N_18400,N_19629);
nand UO_2212 (O_2212,N_18644,N_18339);
xnor UO_2213 (O_2213,N_18983,N_19026);
and UO_2214 (O_2214,N_19051,N_18165);
or UO_2215 (O_2215,N_19085,N_18991);
or UO_2216 (O_2216,N_19189,N_18076);
nor UO_2217 (O_2217,N_18633,N_19624);
nor UO_2218 (O_2218,N_18263,N_18593);
nand UO_2219 (O_2219,N_18018,N_18470);
or UO_2220 (O_2220,N_18247,N_18543);
nor UO_2221 (O_2221,N_18356,N_18096);
or UO_2222 (O_2222,N_19291,N_18621);
and UO_2223 (O_2223,N_18410,N_18751);
or UO_2224 (O_2224,N_19692,N_19615);
nand UO_2225 (O_2225,N_18515,N_18006);
xor UO_2226 (O_2226,N_18204,N_18862);
xnor UO_2227 (O_2227,N_18809,N_18101);
nor UO_2228 (O_2228,N_19691,N_19049);
nor UO_2229 (O_2229,N_18332,N_19102);
nand UO_2230 (O_2230,N_19113,N_19823);
and UO_2231 (O_2231,N_18963,N_18088);
or UO_2232 (O_2232,N_18664,N_18697);
or UO_2233 (O_2233,N_18026,N_19128);
and UO_2234 (O_2234,N_19737,N_18459);
nand UO_2235 (O_2235,N_19021,N_19621);
and UO_2236 (O_2236,N_19085,N_19474);
xor UO_2237 (O_2237,N_19886,N_18970);
nor UO_2238 (O_2238,N_18468,N_19778);
xnor UO_2239 (O_2239,N_18016,N_19412);
nor UO_2240 (O_2240,N_19487,N_19587);
xnor UO_2241 (O_2241,N_18810,N_18595);
and UO_2242 (O_2242,N_18033,N_19922);
nand UO_2243 (O_2243,N_18022,N_18597);
xnor UO_2244 (O_2244,N_18178,N_18366);
nor UO_2245 (O_2245,N_19182,N_18305);
or UO_2246 (O_2246,N_18418,N_19850);
xor UO_2247 (O_2247,N_19582,N_18189);
nand UO_2248 (O_2248,N_18884,N_19287);
and UO_2249 (O_2249,N_19810,N_18361);
and UO_2250 (O_2250,N_18692,N_19102);
nor UO_2251 (O_2251,N_18963,N_19329);
or UO_2252 (O_2252,N_19555,N_18738);
nor UO_2253 (O_2253,N_19547,N_18182);
nand UO_2254 (O_2254,N_19201,N_18716);
nand UO_2255 (O_2255,N_18981,N_18387);
nor UO_2256 (O_2256,N_19784,N_18608);
and UO_2257 (O_2257,N_18906,N_19874);
or UO_2258 (O_2258,N_18473,N_18358);
and UO_2259 (O_2259,N_19348,N_19067);
or UO_2260 (O_2260,N_19074,N_18128);
nand UO_2261 (O_2261,N_18246,N_19061);
nor UO_2262 (O_2262,N_19898,N_18091);
and UO_2263 (O_2263,N_19568,N_19460);
or UO_2264 (O_2264,N_18088,N_19477);
and UO_2265 (O_2265,N_19655,N_18501);
and UO_2266 (O_2266,N_18318,N_18763);
xor UO_2267 (O_2267,N_18128,N_19423);
nor UO_2268 (O_2268,N_19395,N_19282);
xor UO_2269 (O_2269,N_19954,N_18935);
and UO_2270 (O_2270,N_19248,N_18859);
nand UO_2271 (O_2271,N_18070,N_19065);
nand UO_2272 (O_2272,N_19007,N_18778);
nand UO_2273 (O_2273,N_18298,N_18467);
xor UO_2274 (O_2274,N_18282,N_19275);
xor UO_2275 (O_2275,N_18050,N_18512);
xor UO_2276 (O_2276,N_19920,N_19175);
xnor UO_2277 (O_2277,N_19138,N_19507);
or UO_2278 (O_2278,N_18534,N_19283);
nand UO_2279 (O_2279,N_18994,N_18023);
or UO_2280 (O_2280,N_18069,N_18970);
xnor UO_2281 (O_2281,N_19839,N_19548);
nand UO_2282 (O_2282,N_19100,N_19670);
nor UO_2283 (O_2283,N_19593,N_19934);
nor UO_2284 (O_2284,N_18664,N_18183);
xor UO_2285 (O_2285,N_18644,N_18854);
and UO_2286 (O_2286,N_19784,N_19882);
nand UO_2287 (O_2287,N_18995,N_19447);
nand UO_2288 (O_2288,N_18215,N_18113);
or UO_2289 (O_2289,N_19237,N_18251);
nor UO_2290 (O_2290,N_19648,N_18806);
and UO_2291 (O_2291,N_18461,N_19589);
or UO_2292 (O_2292,N_18626,N_19508);
xnor UO_2293 (O_2293,N_19825,N_19376);
xnor UO_2294 (O_2294,N_19597,N_19644);
nor UO_2295 (O_2295,N_18593,N_18354);
and UO_2296 (O_2296,N_18815,N_18379);
or UO_2297 (O_2297,N_18036,N_19133);
or UO_2298 (O_2298,N_19302,N_18381);
nor UO_2299 (O_2299,N_18082,N_19804);
or UO_2300 (O_2300,N_18697,N_18201);
and UO_2301 (O_2301,N_18344,N_19570);
or UO_2302 (O_2302,N_18991,N_19464);
nand UO_2303 (O_2303,N_19581,N_19158);
nand UO_2304 (O_2304,N_18434,N_18405);
nor UO_2305 (O_2305,N_18914,N_19625);
or UO_2306 (O_2306,N_18466,N_19395);
and UO_2307 (O_2307,N_19722,N_18628);
or UO_2308 (O_2308,N_19767,N_18982);
or UO_2309 (O_2309,N_18626,N_19817);
or UO_2310 (O_2310,N_18504,N_18708);
nand UO_2311 (O_2311,N_19873,N_18654);
nor UO_2312 (O_2312,N_18992,N_18406);
xor UO_2313 (O_2313,N_19306,N_19196);
xor UO_2314 (O_2314,N_18024,N_19179);
or UO_2315 (O_2315,N_18305,N_19385);
nor UO_2316 (O_2316,N_19670,N_19126);
nor UO_2317 (O_2317,N_18520,N_19893);
or UO_2318 (O_2318,N_19199,N_19398);
xor UO_2319 (O_2319,N_19208,N_19663);
xor UO_2320 (O_2320,N_19435,N_18069);
and UO_2321 (O_2321,N_19360,N_18236);
or UO_2322 (O_2322,N_19720,N_19257);
nor UO_2323 (O_2323,N_19562,N_18878);
nand UO_2324 (O_2324,N_18885,N_19259);
nand UO_2325 (O_2325,N_19856,N_18056);
nor UO_2326 (O_2326,N_19527,N_19372);
nor UO_2327 (O_2327,N_18931,N_18348);
nand UO_2328 (O_2328,N_18138,N_18823);
nand UO_2329 (O_2329,N_19378,N_19702);
nor UO_2330 (O_2330,N_18103,N_18891);
nand UO_2331 (O_2331,N_19609,N_19061);
xor UO_2332 (O_2332,N_18902,N_19212);
nand UO_2333 (O_2333,N_19938,N_19642);
xnor UO_2334 (O_2334,N_18011,N_18496);
or UO_2335 (O_2335,N_19380,N_19083);
nand UO_2336 (O_2336,N_18093,N_18686);
nand UO_2337 (O_2337,N_19777,N_18038);
xnor UO_2338 (O_2338,N_18350,N_19369);
or UO_2339 (O_2339,N_19288,N_19098);
nand UO_2340 (O_2340,N_18852,N_19956);
xor UO_2341 (O_2341,N_18238,N_18414);
or UO_2342 (O_2342,N_19894,N_19856);
nor UO_2343 (O_2343,N_18960,N_19045);
nor UO_2344 (O_2344,N_18244,N_18079);
or UO_2345 (O_2345,N_19965,N_18595);
or UO_2346 (O_2346,N_19259,N_18577);
nand UO_2347 (O_2347,N_18837,N_19144);
xor UO_2348 (O_2348,N_19176,N_19011);
nand UO_2349 (O_2349,N_19306,N_19992);
or UO_2350 (O_2350,N_18523,N_18020);
xnor UO_2351 (O_2351,N_18781,N_18422);
nand UO_2352 (O_2352,N_18636,N_19795);
and UO_2353 (O_2353,N_19650,N_19860);
xor UO_2354 (O_2354,N_18877,N_18849);
or UO_2355 (O_2355,N_18181,N_18316);
or UO_2356 (O_2356,N_19349,N_19935);
and UO_2357 (O_2357,N_18385,N_19875);
or UO_2358 (O_2358,N_18255,N_19808);
or UO_2359 (O_2359,N_18370,N_18436);
or UO_2360 (O_2360,N_18489,N_19014);
nor UO_2361 (O_2361,N_18616,N_18986);
nor UO_2362 (O_2362,N_18212,N_18269);
and UO_2363 (O_2363,N_19000,N_18440);
xnor UO_2364 (O_2364,N_18738,N_18154);
and UO_2365 (O_2365,N_18314,N_18615);
or UO_2366 (O_2366,N_18823,N_18324);
xnor UO_2367 (O_2367,N_18709,N_18905);
xor UO_2368 (O_2368,N_19726,N_18172);
nand UO_2369 (O_2369,N_18324,N_19570);
nor UO_2370 (O_2370,N_19389,N_19233);
nor UO_2371 (O_2371,N_18646,N_19324);
and UO_2372 (O_2372,N_18582,N_18123);
and UO_2373 (O_2373,N_19654,N_18853);
nand UO_2374 (O_2374,N_19769,N_18923);
xor UO_2375 (O_2375,N_19444,N_19666);
xnor UO_2376 (O_2376,N_19899,N_18622);
and UO_2377 (O_2377,N_19865,N_19431);
xnor UO_2378 (O_2378,N_18962,N_19920);
and UO_2379 (O_2379,N_18264,N_18387);
nor UO_2380 (O_2380,N_19695,N_19197);
nand UO_2381 (O_2381,N_18391,N_18166);
and UO_2382 (O_2382,N_19507,N_18204);
xnor UO_2383 (O_2383,N_19174,N_18538);
and UO_2384 (O_2384,N_19971,N_19912);
or UO_2385 (O_2385,N_18649,N_18609);
and UO_2386 (O_2386,N_19629,N_19519);
nand UO_2387 (O_2387,N_18045,N_18299);
nor UO_2388 (O_2388,N_19572,N_18796);
nor UO_2389 (O_2389,N_18334,N_18752);
xor UO_2390 (O_2390,N_18551,N_18171);
and UO_2391 (O_2391,N_19476,N_18775);
xor UO_2392 (O_2392,N_19611,N_19828);
nand UO_2393 (O_2393,N_19466,N_19722);
and UO_2394 (O_2394,N_19670,N_19593);
nand UO_2395 (O_2395,N_18920,N_18445);
nor UO_2396 (O_2396,N_18762,N_19554);
nand UO_2397 (O_2397,N_19966,N_19869);
and UO_2398 (O_2398,N_19638,N_19958);
and UO_2399 (O_2399,N_18191,N_18909);
or UO_2400 (O_2400,N_18934,N_18865);
xor UO_2401 (O_2401,N_19848,N_19496);
or UO_2402 (O_2402,N_19484,N_19290);
xor UO_2403 (O_2403,N_18116,N_19073);
and UO_2404 (O_2404,N_19967,N_18383);
nor UO_2405 (O_2405,N_18130,N_19833);
xor UO_2406 (O_2406,N_18715,N_19584);
nand UO_2407 (O_2407,N_19084,N_19998);
nand UO_2408 (O_2408,N_19550,N_19110);
and UO_2409 (O_2409,N_18541,N_19259);
xor UO_2410 (O_2410,N_18930,N_18519);
nor UO_2411 (O_2411,N_19464,N_19771);
nand UO_2412 (O_2412,N_19163,N_18315);
nand UO_2413 (O_2413,N_18374,N_19001);
nand UO_2414 (O_2414,N_19429,N_18848);
xor UO_2415 (O_2415,N_19149,N_18874);
nand UO_2416 (O_2416,N_19200,N_19486);
nand UO_2417 (O_2417,N_18833,N_19065);
and UO_2418 (O_2418,N_19841,N_18611);
nand UO_2419 (O_2419,N_18047,N_19503);
nor UO_2420 (O_2420,N_18760,N_18339);
nor UO_2421 (O_2421,N_19183,N_19418);
nand UO_2422 (O_2422,N_18874,N_19106);
nor UO_2423 (O_2423,N_19972,N_18470);
xor UO_2424 (O_2424,N_18357,N_19990);
or UO_2425 (O_2425,N_19881,N_18044);
or UO_2426 (O_2426,N_19289,N_18954);
nor UO_2427 (O_2427,N_19242,N_18655);
nand UO_2428 (O_2428,N_19926,N_18738);
and UO_2429 (O_2429,N_18770,N_19853);
and UO_2430 (O_2430,N_19879,N_18118);
nand UO_2431 (O_2431,N_18483,N_18072);
or UO_2432 (O_2432,N_18143,N_19587);
xor UO_2433 (O_2433,N_19411,N_18836);
and UO_2434 (O_2434,N_18899,N_18024);
nand UO_2435 (O_2435,N_18495,N_18546);
xnor UO_2436 (O_2436,N_19662,N_19221);
and UO_2437 (O_2437,N_18879,N_18793);
xor UO_2438 (O_2438,N_19571,N_19709);
xor UO_2439 (O_2439,N_19282,N_18475);
nand UO_2440 (O_2440,N_19448,N_18351);
xor UO_2441 (O_2441,N_18229,N_19745);
or UO_2442 (O_2442,N_18902,N_18339);
and UO_2443 (O_2443,N_19540,N_18014);
and UO_2444 (O_2444,N_18486,N_18888);
or UO_2445 (O_2445,N_19926,N_19041);
nor UO_2446 (O_2446,N_19560,N_18349);
xor UO_2447 (O_2447,N_19263,N_19697);
or UO_2448 (O_2448,N_19866,N_19107);
nand UO_2449 (O_2449,N_19273,N_18627);
xnor UO_2450 (O_2450,N_19259,N_19467);
nand UO_2451 (O_2451,N_18651,N_18729);
and UO_2452 (O_2452,N_19524,N_18739);
xor UO_2453 (O_2453,N_19146,N_18625);
or UO_2454 (O_2454,N_19078,N_18981);
nor UO_2455 (O_2455,N_18678,N_18673);
and UO_2456 (O_2456,N_18810,N_18692);
or UO_2457 (O_2457,N_18834,N_18575);
nor UO_2458 (O_2458,N_19576,N_18353);
nor UO_2459 (O_2459,N_18545,N_19304);
or UO_2460 (O_2460,N_18619,N_19750);
nor UO_2461 (O_2461,N_19170,N_19308);
nand UO_2462 (O_2462,N_19342,N_19585);
and UO_2463 (O_2463,N_19657,N_19968);
xor UO_2464 (O_2464,N_19177,N_18696);
xor UO_2465 (O_2465,N_19501,N_18421);
nor UO_2466 (O_2466,N_18469,N_18304);
and UO_2467 (O_2467,N_18757,N_18915);
and UO_2468 (O_2468,N_19700,N_19877);
nand UO_2469 (O_2469,N_19715,N_19484);
xor UO_2470 (O_2470,N_19803,N_19428);
nor UO_2471 (O_2471,N_19084,N_19611);
or UO_2472 (O_2472,N_19520,N_18325);
or UO_2473 (O_2473,N_19199,N_19855);
xnor UO_2474 (O_2474,N_18816,N_19499);
or UO_2475 (O_2475,N_18488,N_18502);
and UO_2476 (O_2476,N_18400,N_19451);
nand UO_2477 (O_2477,N_19119,N_18286);
and UO_2478 (O_2478,N_18930,N_18409);
nor UO_2479 (O_2479,N_18932,N_18654);
or UO_2480 (O_2480,N_18489,N_18036);
nor UO_2481 (O_2481,N_19817,N_18489);
nand UO_2482 (O_2482,N_18888,N_18013);
or UO_2483 (O_2483,N_18581,N_18361);
nor UO_2484 (O_2484,N_19593,N_19680);
or UO_2485 (O_2485,N_18206,N_19473);
and UO_2486 (O_2486,N_19875,N_18787);
or UO_2487 (O_2487,N_19829,N_18897);
and UO_2488 (O_2488,N_19987,N_18433);
xor UO_2489 (O_2489,N_19698,N_19016);
xor UO_2490 (O_2490,N_18379,N_19666);
nand UO_2491 (O_2491,N_19085,N_19035);
xnor UO_2492 (O_2492,N_19790,N_18203);
nor UO_2493 (O_2493,N_19515,N_19098);
xnor UO_2494 (O_2494,N_19810,N_18278);
nor UO_2495 (O_2495,N_19163,N_19098);
nor UO_2496 (O_2496,N_18809,N_19532);
or UO_2497 (O_2497,N_18469,N_18939);
nor UO_2498 (O_2498,N_18245,N_18669);
and UO_2499 (O_2499,N_19948,N_18505);
endmodule