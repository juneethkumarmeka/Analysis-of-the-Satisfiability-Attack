module basic_1000_10000_1500_5_levels_2xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nand U0 (N_0,In_740,In_708);
nor U1 (N_1,In_553,In_6);
or U2 (N_2,In_790,In_774);
nor U3 (N_3,In_683,In_654);
or U4 (N_4,In_437,In_552);
nor U5 (N_5,In_45,In_797);
nand U6 (N_6,In_153,In_501);
and U7 (N_7,In_17,In_756);
nand U8 (N_8,In_559,In_825);
or U9 (N_9,In_281,In_180);
or U10 (N_10,In_784,In_27);
and U11 (N_11,In_212,In_700);
nor U12 (N_12,In_758,In_389);
and U13 (N_13,In_912,In_21);
and U14 (N_14,In_283,In_253);
nor U15 (N_15,In_833,In_210);
and U16 (N_16,In_342,In_584);
nand U17 (N_17,In_38,In_331);
or U18 (N_18,In_175,In_427);
nor U19 (N_19,In_47,In_676);
or U20 (N_20,In_960,In_117);
and U21 (N_21,In_773,In_159);
nand U22 (N_22,In_977,In_177);
or U23 (N_23,In_375,In_338);
nor U24 (N_24,In_981,In_674);
and U25 (N_25,In_793,In_333);
or U26 (N_26,In_271,In_964);
nor U27 (N_27,In_927,In_255);
nand U28 (N_28,In_258,In_318);
nor U29 (N_29,In_938,In_532);
nor U30 (N_30,In_818,In_934);
and U31 (N_31,In_109,In_178);
and U32 (N_32,In_777,In_989);
and U33 (N_33,In_902,In_138);
nand U34 (N_34,In_441,In_165);
and U35 (N_35,In_382,In_174);
nand U36 (N_36,In_79,In_594);
or U37 (N_37,In_666,In_794);
nand U38 (N_38,In_30,In_800);
or U39 (N_39,In_328,In_839);
and U40 (N_40,In_209,In_298);
nand U41 (N_41,In_768,In_761);
and U42 (N_42,In_639,In_698);
nand U43 (N_43,In_324,In_963);
and U44 (N_44,In_668,In_837);
nor U45 (N_45,In_918,In_411);
nand U46 (N_46,In_134,In_414);
or U47 (N_47,In_861,In_597);
and U48 (N_48,In_786,In_107);
nand U49 (N_49,In_645,In_815);
or U50 (N_50,In_471,In_518);
and U51 (N_51,In_403,In_944);
nor U52 (N_52,In_882,In_785);
and U53 (N_53,In_408,In_326);
or U54 (N_54,In_57,In_462);
or U55 (N_55,In_200,In_713);
nand U56 (N_56,In_937,In_863);
nand U57 (N_57,In_737,In_536);
and U58 (N_58,In_776,In_633);
nor U59 (N_59,In_73,In_940);
and U60 (N_60,In_739,In_859);
and U61 (N_61,In_933,In_978);
nor U62 (N_62,In_686,In_280);
nor U63 (N_63,In_868,In_161);
nand U64 (N_64,In_976,In_923);
or U65 (N_65,In_231,In_359);
or U66 (N_66,In_315,In_80);
nand U67 (N_67,In_75,In_354);
nor U68 (N_68,In_631,In_448);
or U69 (N_69,In_916,In_580);
nor U70 (N_70,In_391,In_337);
or U71 (N_71,In_495,In_906);
nand U72 (N_72,In_856,In_910);
and U73 (N_73,In_77,In_339);
nor U74 (N_74,In_541,In_755);
nand U75 (N_75,In_903,In_702);
nor U76 (N_76,In_945,In_742);
nand U77 (N_77,In_751,In_491);
nor U78 (N_78,In_808,In_929);
and U79 (N_79,In_44,In_40);
or U80 (N_80,In_424,In_274);
nor U81 (N_81,In_162,In_406);
nor U82 (N_82,In_4,In_886);
nor U83 (N_83,In_156,In_309);
nor U84 (N_84,In_572,In_879);
nor U85 (N_85,In_19,In_596);
or U86 (N_86,In_419,In_197);
or U87 (N_87,In_465,In_121);
nand U88 (N_88,In_582,In_360);
or U89 (N_89,In_704,In_176);
nand U90 (N_90,In_904,In_148);
xnor U91 (N_91,In_781,In_997);
nand U92 (N_92,In_726,In_529);
nand U93 (N_93,In_993,In_642);
or U94 (N_94,In_621,In_190);
or U95 (N_95,In_105,In_681);
xnor U96 (N_96,In_504,In_191);
nand U97 (N_97,In_377,In_822);
and U98 (N_98,In_196,In_507);
and U99 (N_99,In_242,In_72);
and U100 (N_100,In_962,In_990);
nand U101 (N_101,In_523,In_450);
or U102 (N_102,In_98,In_358);
or U103 (N_103,In_843,In_587);
nor U104 (N_104,In_18,In_249);
nand U105 (N_105,In_136,In_239);
or U106 (N_106,In_278,In_476);
xnor U107 (N_107,In_772,In_519);
or U108 (N_108,In_458,In_24);
nand U109 (N_109,In_583,In_764);
nor U110 (N_110,In_444,In_889);
and U111 (N_111,In_881,In_157);
or U112 (N_112,In_376,In_59);
nor U113 (N_113,In_703,In_928);
nand U114 (N_114,In_853,In_97);
or U115 (N_115,In_67,In_567);
nor U116 (N_116,In_623,In_284);
nor U117 (N_117,In_82,In_41);
and U118 (N_118,In_449,In_343);
nand U119 (N_119,In_132,In_538);
or U120 (N_120,In_693,In_12);
nor U121 (N_121,In_247,In_464);
nor U122 (N_122,In_512,In_958);
or U123 (N_123,In_22,In_617);
nand U124 (N_124,In_113,In_514);
nor U125 (N_125,In_561,In_468);
nand U126 (N_126,In_168,In_540);
or U127 (N_127,In_206,In_480);
nor U128 (N_128,In_380,In_695);
or U129 (N_129,In_723,In_469);
or U130 (N_130,In_463,In_876);
or U131 (N_131,In_240,In_615);
and U132 (N_132,In_96,In_675);
or U133 (N_133,In_575,In_943);
nor U134 (N_134,In_460,In_854);
or U135 (N_135,In_942,In_544);
nor U136 (N_136,In_586,In_126);
nand U137 (N_137,In_51,In_81);
and U138 (N_138,In_423,In_896);
nand U139 (N_139,In_515,In_361);
and U140 (N_140,In_619,In_749);
and U141 (N_141,In_558,In_763);
and U142 (N_142,In_48,In_579);
or U143 (N_143,In_33,In_849);
nand U144 (N_144,In_50,In_946);
nand U145 (N_145,In_277,In_806);
and U146 (N_146,In_771,In_517);
nand U147 (N_147,In_133,In_895);
nand U148 (N_148,In_577,In_202);
nand U149 (N_149,In_101,In_497);
nand U150 (N_150,In_84,In_248);
nor U151 (N_151,In_110,In_474);
nor U152 (N_152,In_643,In_418);
or U153 (N_153,In_778,In_791);
nand U154 (N_154,In_893,In_201);
or U155 (N_155,In_730,In_400);
and U156 (N_156,In_883,In_754);
and U157 (N_157,In_139,In_744);
or U158 (N_158,In_263,In_104);
nor U159 (N_159,In_917,In_959);
nor U160 (N_160,In_349,In_769);
nor U161 (N_161,In_690,In_61);
nand U162 (N_162,In_919,In_598);
and U163 (N_163,In_647,In_446);
nor U164 (N_164,In_119,In_262);
nand U165 (N_165,In_115,In_860);
or U166 (N_166,In_238,In_312);
nor U167 (N_167,In_485,In_844);
or U168 (N_168,In_106,In_346);
or U169 (N_169,In_76,In_53);
nor U170 (N_170,In_43,In_957);
or U171 (N_171,In_295,In_630);
or U172 (N_172,In_653,In_847);
and U173 (N_173,In_569,In_166);
nand U174 (N_174,In_762,In_838);
nand U175 (N_175,In_649,In_272);
nor U176 (N_176,In_486,In_885);
nor U177 (N_177,In_520,In_691);
nor U178 (N_178,In_546,In_760);
or U179 (N_179,In_306,In_116);
nor U180 (N_180,In_32,In_842);
nand U181 (N_181,In_807,In_875);
and U182 (N_182,In_369,In_734);
nor U183 (N_183,In_15,In_454);
or U184 (N_184,In_588,In_398);
nor U185 (N_185,In_214,In_827);
or U186 (N_186,In_69,In_371);
or U187 (N_187,In_207,In_429);
nand U188 (N_188,In_143,In_11);
or U189 (N_189,In_221,In_974);
or U190 (N_190,In_128,In_140);
and U191 (N_191,In_28,In_409);
nand U192 (N_192,In_564,In_129);
nor U193 (N_193,In_144,In_951);
nand U194 (N_194,In_287,In_732);
or U195 (N_195,In_600,In_9);
or U196 (N_196,In_415,In_325);
nand U197 (N_197,In_152,In_370);
nand U198 (N_198,In_194,In_864);
or U199 (N_199,In_641,In_692);
nand U200 (N_200,In_788,In_801);
and U201 (N_201,In_810,In_330);
nor U202 (N_202,In_817,In_372);
nor U203 (N_203,In_770,In_884);
or U204 (N_204,In_646,In_605);
and U205 (N_205,In_31,In_273);
nand U206 (N_206,In_672,In_150);
nor U207 (N_207,In_706,In_952);
or U208 (N_208,In_440,In_521);
nand U209 (N_209,In_809,In_921);
and U210 (N_210,In_319,In_767);
nand U211 (N_211,In_846,In_393);
or U212 (N_212,In_955,In_688);
or U213 (N_213,In_738,In_871);
or U214 (N_214,In_112,In_385);
and U215 (N_215,In_932,In_498);
nand U216 (N_216,In_114,In_867);
nor U217 (N_217,In_717,In_604);
nor U218 (N_218,In_589,In_612);
nand U219 (N_219,In_877,In_215);
nor U220 (N_220,In_673,In_897);
nand U221 (N_221,In_595,In_980);
nand U222 (N_222,In_716,In_765);
or U223 (N_223,In_223,In_0);
nand U224 (N_224,In_805,In_386);
or U225 (N_225,In_626,In_147);
nand U226 (N_226,In_823,In_865);
or U227 (N_227,In_551,In_236);
nand U228 (N_228,In_489,In_430);
nand U229 (N_229,In_968,In_873);
nand U230 (N_230,In_443,In_122);
nand U231 (N_231,In_227,In_611);
nand U232 (N_232,In_137,In_205);
nor U233 (N_233,In_14,In_267);
or U234 (N_234,In_718,In_590);
nor U235 (N_235,In_426,In_379);
nand U236 (N_236,In_746,In_5);
or U237 (N_237,In_701,In_811);
nor U238 (N_238,In_91,In_986);
nor U239 (N_239,In_949,In_591);
nand U240 (N_240,In_678,In_145);
nor U241 (N_241,In_752,In_696);
or U242 (N_242,In_317,In_270);
or U243 (N_243,In_282,In_42);
nor U244 (N_244,In_336,In_650);
nand U245 (N_245,In_250,In_340);
and U246 (N_246,In_783,In_365);
nand U247 (N_247,In_658,In_571);
and U248 (N_248,In_260,In_939);
and U249 (N_249,In_813,In_614);
nand U250 (N_250,In_357,In_94);
nand U251 (N_251,In_640,In_728);
xor U252 (N_252,In_92,In_301);
nor U253 (N_253,In_729,In_494);
or U254 (N_254,In_83,In_473);
or U255 (N_255,In_313,In_417);
nand U256 (N_256,In_627,In_715);
nand U257 (N_257,In_870,In_131);
nand U258 (N_258,In_350,In_276);
nor U259 (N_259,In_7,In_830);
nand U260 (N_260,In_511,In_635);
nor U261 (N_261,In_85,In_648);
and U262 (N_262,In_233,In_714);
nor U263 (N_263,In_508,In_130);
and U264 (N_264,In_362,In_931);
and U265 (N_265,In_905,In_432);
and U266 (N_266,In_172,In_509);
and U267 (N_267,In_438,In_186);
or U268 (N_268,In_505,In_736);
nand U269 (N_269,In_181,In_188);
nand U270 (N_270,In_163,In_36);
and U271 (N_271,In_593,In_279);
or U272 (N_272,In_499,In_108);
and U273 (N_273,In_345,In_911);
nand U274 (N_274,In_164,In_506);
and U275 (N_275,In_71,In_599);
nand U276 (N_276,In_545,In_891);
nand U277 (N_277,In_55,In_447);
and U278 (N_278,In_62,In_971);
or U279 (N_279,In_405,In_20);
nand U280 (N_280,In_433,In_251);
nand U281 (N_281,In_522,In_327);
nor U282 (N_282,In_965,In_457);
and U283 (N_283,In_219,In_234);
nand U284 (N_284,In_887,In_435);
nor U285 (N_285,In_568,In_404);
and U286 (N_286,In_490,In_332);
nand U287 (N_287,In_821,In_845);
nor U288 (N_288,In_195,In_824);
and U289 (N_289,In_149,In_347);
nand U290 (N_290,In_265,In_620);
or U291 (N_291,In_973,In_743);
nor U292 (N_292,In_733,In_314);
and U293 (N_293,In_747,In_256);
and U294 (N_294,In_70,In_413);
or U295 (N_295,In_235,In_442);
nand U296 (N_296,In_982,In_302);
nand U297 (N_297,In_320,In_218);
nand U298 (N_298,In_991,In_3);
and U299 (N_299,In_554,In_697);
and U300 (N_300,In_228,In_607);
nor U301 (N_301,In_23,In_213);
nor U302 (N_302,In_890,In_657);
nand U303 (N_303,In_920,In_914);
nand U304 (N_304,In_851,In_211);
nand U305 (N_305,In_880,In_95);
or U306 (N_306,In_812,In_34);
nor U307 (N_307,In_539,In_60);
nor U308 (N_308,In_828,In_748);
and U309 (N_309,In_637,In_798);
nor U310 (N_310,In_470,In_574);
nand U311 (N_311,In_608,In_585);
or U312 (N_312,In_225,In_322);
and U313 (N_313,In_556,In_226);
nand U314 (N_314,In_563,In_745);
nand U315 (N_315,In_461,In_930);
nor U316 (N_316,In_609,In_988);
nand U317 (N_317,In_992,In_570);
nand U318 (N_318,In_158,In_364);
or U319 (N_319,In_90,In_802);
nand U320 (N_320,In_995,In_689);
and U321 (N_321,In_455,In_775);
nand U322 (N_322,In_296,In_682);
or U323 (N_323,In_52,In_146);
nand U324 (N_324,In_664,In_819);
nand U325 (N_325,In_516,In_266);
or U326 (N_326,In_118,In_560);
nand U327 (N_327,In_54,In_453);
nor U328 (N_328,In_155,In_535);
or U329 (N_329,In_220,In_628);
nand U330 (N_330,In_492,In_548);
or U331 (N_331,In_624,In_581);
nand U332 (N_332,In_8,In_954);
nor U333 (N_333,In_759,In_387);
and U334 (N_334,In_638,In_335);
nor U335 (N_335,In_410,In_757);
and U336 (N_336,In_294,In_305);
nor U337 (N_337,In_99,In_245);
nand U338 (N_338,In_392,In_334);
and U339 (N_339,In_709,In_680);
and U340 (N_340,In_451,In_779);
or U341 (N_341,In_669,In_618);
nand U342 (N_342,In_852,In_994);
nand U343 (N_343,In_479,In_151);
or U344 (N_344,In_987,In_431);
or U345 (N_345,In_1,In_789);
and U346 (N_346,In_254,In_719);
nor U347 (N_347,In_374,In_894);
nor U348 (N_348,In_803,In_16);
nand U349 (N_349,In_656,In_537);
and U350 (N_350,In_950,In_241);
or U351 (N_351,In_29,In_565);
nand U352 (N_352,In_169,In_420);
nand U353 (N_353,In_292,In_383);
nand U354 (N_354,In_592,In_304);
and U355 (N_355,In_753,In_183);
and U356 (N_356,In_125,In_780);
nor U357 (N_357,In_766,In_244);
nand U358 (N_358,In_86,In_711);
nor U359 (N_359,In_731,In_829);
and U360 (N_360,In_983,In_232);
or U361 (N_361,In_401,In_834);
nor U362 (N_362,In_500,In_268);
and U363 (N_363,In_351,In_722);
nor U364 (N_364,In_124,In_64);
and U365 (N_365,In_578,In_100);
nor U366 (N_366,In_475,In_625);
nand U367 (N_367,In_542,In_229);
or U368 (N_368,In_66,In_549);
and U369 (N_369,In_310,In_291);
or U370 (N_370,In_869,In_198);
and U371 (N_371,In_493,In_308);
nor U372 (N_372,In_230,In_841);
nand U373 (N_373,In_452,In_900);
nor U374 (N_374,In_550,In_353);
or U375 (N_375,In_872,In_961);
nand U376 (N_376,In_685,In_329);
or U377 (N_377,In_56,In_46);
and U378 (N_378,In_727,In_792);
or U379 (N_379,In_68,In_533);
nor U380 (N_380,In_366,In_513);
and U381 (N_381,In_297,In_356);
or U382 (N_382,In_384,In_710);
nand U383 (N_383,In_472,In_381);
nand U384 (N_384,In_120,In_246);
nand U385 (N_385,In_913,In_78);
and U386 (N_386,In_321,In_217);
nor U387 (N_387,In_93,In_243);
nor U388 (N_388,In_699,In_445);
or U389 (N_389,In_831,In_275);
and U390 (N_390,In_526,In_257);
xor U391 (N_391,In_679,In_288);
and U392 (N_392,In_835,In_316);
or U393 (N_393,In_502,In_855);
and U394 (N_394,In_103,In_483);
and U395 (N_395,In_557,In_179);
or U396 (N_396,In_111,In_832);
nand U397 (N_397,In_467,In_850);
and U398 (N_398,In_300,In_299);
and U399 (N_399,In_503,In_208);
nor U400 (N_400,In_947,In_488);
nor U401 (N_401,In_555,In_456);
nand U402 (N_402,In_707,In_799);
nor U403 (N_403,In_979,In_787);
and U404 (N_404,In_936,In_795);
or U405 (N_405,In_355,In_915);
nor U406 (N_406,In_665,In_684);
or U407 (N_407,In_524,In_264);
nand U408 (N_408,In_397,In_636);
nand U409 (N_409,In_394,In_428);
nor U410 (N_410,In_694,In_422);
and U411 (N_411,In_935,In_848);
nand U412 (N_412,In_712,In_661);
nand U413 (N_413,In_65,In_286);
nand U414 (N_414,In_127,In_725);
nand U415 (N_415,In_613,In_416);
nand U416 (N_416,In_237,In_434);
xnor U417 (N_417,In_412,In_368);
and U418 (N_418,In_193,In_204);
and U419 (N_419,In_290,In_459);
nand U420 (N_420,In_189,In_816);
nand U421 (N_421,In_750,In_13);
and U422 (N_422,In_363,In_285);
and U423 (N_423,In_953,In_820);
or U424 (N_424,In_926,In_622);
and U425 (N_425,In_466,In_970);
nor U426 (N_426,In_123,In_814);
or U427 (N_427,In_606,In_396);
xnor U428 (N_428,In_135,In_252);
nor U429 (N_429,In_601,In_909);
nor U430 (N_430,In_141,In_173);
nor U431 (N_431,In_25,In_348);
nand U432 (N_432,In_941,In_184);
nor U433 (N_433,In_74,In_222);
nand U434 (N_434,In_187,In_956);
or U435 (N_435,In_667,In_610);
nand U436 (N_436,In_858,In_436);
and U437 (N_437,In_857,In_259);
nand U438 (N_438,In_655,In_477);
nand U439 (N_439,In_487,In_402);
nor U440 (N_440,In_677,In_63);
nand U441 (N_441,In_660,In_407);
and U442 (N_442,In_311,In_167);
nand U443 (N_443,In_439,In_566);
nand U444 (N_444,In_373,In_616);
nand U445 (N_445,In_88,In_2);
nand U446 (N_446,In_878,In_293);
nor U447 (N_447,In_874,In_87);
and U448 (N_448,In_528,In_199);
xor U449 (N_449,In_659,In_662);
nor U450 (N_450,In_948,In_898);
or U451 (N_451,In_352,In_826);
or U452 (N_452,In_573,In_721);
nand U453 (N_453,In_999,In_323);
nand U454 (N_454,In_344,In_525);
or U455 (N_455,In_289,In_527);
and U456 (N_456,In_261,In_367);
nor U457 (N_457,In_972,In_154);
or U458 (N_458,In_862,In_705);
nor U459 (N_459,In_303,In_496);
and U460 (N_460,In_530,In_171);
nand U461 (N_461,In_170,In_741);
and U462 (N_462,In_924,In_576);
or U463 (N_463,In_603,In_35);
or U464 (N_464,In_142,In_378);
nor U465 (N_465,In_644,In_421);
and U466 (N_466,In_866,In_203);
and U467 (N_467,In_39,In_836);
and U468 (N_468,In_804,In_484);
nand U469 (N_469,In_269,In_796);
nand U470 (N_470,In_602,In_984);
nor U471 (N_471,In_562,In_975);
or U472 (N_472,In_735,In_388);
nand U473 (N_473,In_26,In_224);
and U474 (N_474,In_89,In_998);
or U475 (N_475,In_996,In_724);
or U476 (N_476,In_481,In_37);
nand U477 (N_477,In_922,In_969);
nand U478 (N_478,In_892,In_341);
or U479 (N_479,In_888,In_907);
and U480 (N_480,In_925,In_840);
and U481 (N_481,In_192,In_307);
nand U482 (N_482,In_671,In_102);
nor U483 (N_483,In_216,In_510);
nand U484 (N_484,In_49,In_901);
and U485 (N_485,In_652,In_543);
or U486 (N_486,In_632,In_547);
or U487 (N_487,In_182,In_531);
and U488 (N_488,In_399,In_651);
or U489 (N_489,In_687,In_10);
or U490 (N_490,In_670,In_482);
nand U491 (N_491,In_425,In_720);
nor U492 (N_492,In_899,In_395);
nand U493 (N_493,In_782,In_185);
nand U494 (N_494,In_985,In_629);
nor U495 (N_495,In_160,In_908);
or U496 (N_496,In_58,In_534);
or U497 (N_497,In_663,In_966);
or U498 (N_498,In_634,In_967);
or U499 (N_499,In_478,In_390);
nand U500 (N_500,In_874,In_100);
or U501 (N_501,In_608,In_723);
nand U502 (N_502,In_204,In_822);
xor U503 (N_503,In_35,In_31);
or U504 (N_504,In_767,In_567);
nand U505 (N_505,In_637,In_333);
nor U506 (N_506,In_593,In_873);
or U507 (N_507,In_82,In_140);
or U508 (N_508,In_58,In_750);
nand U509 (N_509,In_357,In_320);
or U510 (N_510,In_400,In_610);
or U511 (N_511,In_165,In_394);
or U512 (N_512,In_857,In_874);
nand U513 (N_513,In_635,In_364);
or U514 (N_514,In_114,In_939);
and U515 (N_515,In_220,In_767);
or U516 (N_516,In_709,In_309);
nand U517 (N_517,In_80,In_65);
and U518 (N_518,In_513,In_569);
or U519 (N_519,In_236,In_411);
or U520 (N_520,In_871,In_233);
or U521 (N_521,In_7,In_46);
and U522 (N_522,In_242,In_705);
nand U523 (N_523,In_515,In_341);
nand U524 (N_524,In_212,In_951);
nor U525 (N_525,In_870,In_741);
nor U526 (N_526,In_381,In_546);
nand U527 (N_527,In_317,In_691);
nand U528 (N_528,In_994,In_160);
nand U529 (N_529,In_572,In_316);
or U530 (N_530,In_499,In_619);
or U531 (N_531,In_717,In_856);
nand U532 (N_532,In_593,In_364);
nand U533 (N_533,In_280,In_364);
or U534 (N_534,In_832,In_411);
or U535 (N_535,In_952,In_853);
nand U536 (N_536,In_844,In_334);
nand U537 (N_537,In_692,In_33);
nand U538 (N_538,In_17,In_175);
and U539 (N_539,In_680,In_688);
and U540 (N_540,In_680,In_842);
or U541 (N_541,In_26,In_31);
nor U542 (N_542,In_891,In_130);
nand U543 (N_543,In_567,In_876);
and U544 (N_544,In_965,In_316);
and U545 (N_545,In_91,In_314);
nand U546 (N_546,In_596,In_185);
and U547 (N_547,In_526,In_743);
nand U548 (N_548,In_458,In_589);
xnor U549 (N_549,In_564,In_482);
nor U550 (N_550,In_159,In_429);
or U551 (N_551,In_436,In_81);
or U552 (N_552,In_755,In_743);
and U553 (N_553,In_383,In_395);
nor U554 (N_554,In_573,In_246);
nand U555 (N_555,In_593,In_148);
and U556 (N_556,In_130,In_109);
nor U557 (N_557,In_568,In_197);
nor U558 (N_558,In_183,In_19);
and U559 (N_559,In_161,In_706);
or U560 (N_560,In_304,In_605);
and U561 (N_561,In_359,In_95);
nand U562 (N_562,In_655,In_127);
xnor U563 (N_563,In_471,In_291);
nand U564 (N_564,In_375,In_497);
nand U565 (N_565,In_371,In_873);
nor U566 (N_566,In_658,In_993);
or U567 (N_567,In_997,In_192);
nor U568 (N_568,In_411,In_707);
nand U569 (N_569,In_356,In_526);
nand U570 (N_570,In_470,In_391);
and U571 (N_571,In_763,In_406);
and U572 (N_572,In_973,In_797);
nand U573 (N_573,In_971,In_650);
nor U574 (N_574,In_734,In_44);
xor U575 (N_575,In_150,In_277);
or U576 (N_576,In_241,In_890);
nand U577 (N_577,In_502,In_812);
nor U578 (N_578,In_602,In_328);
or U579 (N_579,In_161,In_209);
nand U580 (N_580,In_828,In_87);
nand U581 (N_581,In_140,In_538);
or U582 (N_582,In_453,In_854);
nand U583 (N_583,In_723,In_293);
and U584 (N_584,In_598,In_580);
and U585 (N_585,In_830,In_177);
and U586 (N_586,In_857,In_489);
and U587 (N_587,In_470,In_376);
nand U588 (N_588,In_333,In_812);
nor U589 (N_589,In_715,In_854);
or U590 (N_590,In_919,In_309);
nand U591 (N_591,In_559,In_16);
or U592 (N_592,In_215,In_331);
and U593 (N_593,In_904,In_85);
and U594 (N_594,In_863,In_328);
nor U595 (N_595,In_352,In_468);
and U596 (N_596,In_601,In_581);
and U597 (N_597,In_687,In_848);
nand U598 (N_598,In_64,In_154);
nand U599 (N_599,In_748,In_977);
and U600 (N_600,In_855,In_439);
nand U601 (N_601,In_912,In_111);
nor U602 (N_602,In_825,In_106);
or U603 (N_603,In_885,In_774);
nor U604 (N_604,In_265,In_447);
nand U605 (N_605,In_651,In_878);
nand U606 (N_606,In_931,In_975);
or U607 (N_607,In_11,In_85);
and U608 (N_608,In_441,In_389);
or U609 (N_609,In_745,In_743);
and U610 (N_610,In_853,In_988);
nor U611 (N_611,In_939,In_66);
xnor U612 (N_612,In_761,In_312);
nand U613 (N_613,In_697,In_101);
and U614 (N_614,In_950,In_692);
and U615 (N_615,In_262,In_572);
and U616 (N_616,In_732,In_691);
xor U617 (N_617,In_645,In_226);
nand U618 (N_618,In_604,In_459);
nand U619 (N_619,In_89,In_349);
and U620 (N_620,In_823,In_275);
and U621 (N_621,In_575,In_468);
and U622 (N_622,In_650,In_132);
nor U623 (N_623,In_477,In_32);
nor U624 (N_624,In_449,In_980);
xor U625 (N_625,In_654,In_519);
nor U626 (N_626,In_963,In_464);
or U627 (N_627,In_473,In_976);
nand U628 (N_628,In_825,In_853);
xor U629 (N_629,In_398,In_701);
nand U630 (N_630,In_543,In_538);
nand U631 (N_631,In_140,In_604);
and U632 (N_632,In_116,In_173);
or U633 (N_633,In_396,In_978);
nor U634 (N_634,In_102,In_786);
xor U635 (N_635,In_983,In_427);
or U636 (N_636,In_791,In_876);
and U637 (N_637,In_146,In_791);
nor U638 (N_638,In_884,In_142);
or U639 (N_639,In_451,In_984);
and U640 (N_640,In_948,In_719);
and U641 (N_641,In_585,In_899);
and U642 (N_642,In_464,In_954);
nor U643 (N_643,In_698,In_901);
or U644 (N_644,In_332,In_817);
and U645 (N_645,In_688,In_218);
nor U646 (N_646,In_126,In_654);
or U647 (N_647,In_175,In_847);
nand U648 (N_648,In_109,In_37);
nor U649 (N_649,In_947,In_788);
or U650 (N_650,In_872,In_568);
nand U651 (N_651,In_144,In_373);
and U652 (N_652,In_685,In_140);
nand U653 (N_653,In_379,In_230);
or U654 (N_654,In_958,In_604);
and U655 (N_655,In_788,In_633);
nor U656 (N_656,In_390,In_436);
nand U657 (N_657,In_458,In_332);
nand U658 (N_658,In_691,In_313);
nand U659 (N_659,In_528,In_147);
and U660 (N_660,In_977,In_12);
nor U661 (N_661,In_902,In_657);
nand U662 (N_662,In_312,In_199);
nor U663 (N_663,In_878,In_798);
or U664 (N_664,In_55,In_957);
or U665 (N_665,In_783,In_568);
xnor U666 (N_666,In_192,In_825);
nor U667 (N_667,In_969,In_160);
and U668 (N_668,In_378,In_457);
and U669 (N_669,In_50,In_157);
or U670 (N_670,In_688,In_731);
or U671 (N_671,In_723,In_383);
nand U672 (N_672,In_74,In_688);
nor U673 (N_673,In_439,In_259);
and U674 (N_674,In_901,In_267);
nand U675 (N_675,In_854,In_426);
nor U676 (N_676,In_116,In_480);
or U677 (N_677,In_404,In_62);
nor U678 (N_678,In_828,In_968);
nor U679 (N_679,In_497,In_976);
or U680 (N_680,In_876,In_602);
nor U681 (N_681,In_390,In_673);
xnor U682 (N_682,In_547,In_853);
nor U683 (N_683,In_94,In_510);
and U684 (N_684,In_220,In_618);
and U685 (N_685,In_342,In_359);
or U686 (N_686,In_130,In_708);
and U687 (N_687,In_500,In_428);
and U688 (N_688,In_849,In_581);
nor U689 (N_689,In_756,In_868);
nor U690 (N_690,In_192,In_144);
nor U691 (N_691,In_142,In_230);
nor U692 (N_692,In_912,In_515);
or U693 (N_693,In_963,In_247);
and U694 (N_694,In_781,In_794);
nor U695 (N_695,In_305,In_581);
and U696 (N_696,In_901,In_363);
nor U697 (N_697,In_447,In_465);
and U698 (N_698,In_322,In_942);
xor U699 (N_699,In_940,In_471);
nor U700 (N_700,In_203,In_114);
or U701 (N_701,In_983,In_562);
or U702 (N_702,In_128,In_14);
nor U703 (N_703,In_914,In_142);
and U704 (N_704,In_322,In_680);
or U705 (N_705,In_342,In_83);
or U706 (N_706,In_373,In_400);
and U707 (N_707,In_624,In_547);
nor U708 (N_708,In_739,In_52);
or U709 (N_709,In_91,In_640);
or U710 (N_710,In_429,In_749);
or U711 (N_711,In_781,In_156);
and U712 (N_712,In_855,In_707);
nor U713 (N_713,In_942,In_941);
nor U714 (N_714,In_118,In_807);
nand U715 (N_715,In_945,In_155);
nor U716 (N_716,In_33,In_947);
xor U717 (N_717,In_567,In_647);
nor U718 (N_718,In_439,In_37);
or U719 (N_719,In_9,In_531);
or U720 (N_720,In_66,In_95);
nand U721 (N_721,In_636,In_757);
or U722 (N_722,In_216,In_691);
nor U723 (N_723,In_369,In_336);
or U724 (N_724,In_577,In_334);
xnor U725 (N_725,In_867,In_611);
or U726 (N_726,In_952,In_869);
and U727 (N_727,In_425,In_874);
and U728 (N_728,In_817,In_28);
nor U729 (N_729,In_942,In_454);
nor U730 (N_730,In_267,In_310);
nor U731 (N_731,In_919,In_116);
nand U732 (N_732,In_466,In_726);
or U733 (N_733,In_986,In_360);
nor U734 (N_734,In_159,In_633);
nand U735 (N_735,In_288,In_320);
nor U736 (N_736,In_68,In_45);
or U737 (N_737,In_618,In_892);
or U738 (N_738,In_960,In_296);
nand U739 (N_739,In_527,In_419);
or U740 (N_740,In_652,In_327);
nor U741 (N_741,In_300,In_790);
or U742 (N_742,In_840,In_563);
or U743 (N_743,In_33,In_628);
and U744 (N_744,In_70,In_177);
nor U745 (N_745,In_533,In_51);
or U746 (N_746,In_1,In_97);
nand U747 (N_747,In_893,In_361);
or U748 (N_748,In_481,In_333);
and U749 (N_749,In_875,In_760);
or U750 (N_750,In_804,In_970);
and U751 (N_751,In_639,In_669);
nor U752 (N_752,In_364,In_189);
or U753 (N_753,In_247,In_837);
or U754 (N_754,In_568,In_347);
nand U755 (N_755,In_766,In_959);
xor U756 (N_756,In_400,In_147);
and U757 (N_757,In_929,In_821);
or U758 (N_758,In_243,In_876);
nand U759 (N_759,In_975,In_419);
nor U760 (N_760,In_668,In_42);
nor U761 (N_761,In_81,In_434);
nand U762 (N_762,In_431,In_728);
xor U763 (N_763,In_205,In_592);
nor U764 (N_764,In_930,In_775);
and U765 (N_765,In_152,In_210);
and U766 (N_766,In_274,In_558);
or U767 (N_767,In_951,In_862);
or U768 (N_768,In_655,In_502);
or U769 (N_769,In_631,In_409);
and U770 (N_770,In_967,In_784);
and U771 (N_771,In_861,In_552);
or U772 (N_772,In_548,In_804);
or U773 (N_773,In_25,In_999);
or U774 (N_774,In_259,In_70);
and U775 (N_775,In_883,In_13);
nor U776 (N_776,In_921,In_234);
or U777 (N_777,In_508,In_103);
and U778 (N_778,In_608,In_707);
or U779 (N_779,In_183,In_129);
nand U780 (N_780,In_884,In_0);
and U781 (N_781,In_862,In_719);
or U782 (N_782,In_113,In_297);
nor U783 (N_783,In_151,In_56);
xor U784 (N_784,In_456,In_637);
or U785 (N_785,In_53,In_688);
nand U786 (N_786,In_887,In_994);
nand U787 (N_787,In_818,In_822);
or U788 (N_788,In_862,In_139);
and U789 (N_789,In_34,In_893);
or U790 (N_790,In_575,In_848);
and U791 (N_791,In_247,In_750);
or U792 (N_792,In_439,In_580);
xnor U793 (N_793,In_720,In_823);
nand U794 (N_794,In_294,In_810);
nor U795 (N_795,In_122,In_827);
nor U796 (N_796,In_482,In_283);
and U797 (N_797,In_660,In_522);
or U798 (N_798,In_529,In_94);
xnor U799 (N_799,In_172,In_422);
nor U800 (N_800,In_962,In_702);
nor U801 (N_801,In_812,In_708);
or U802 (N_802,In_496,In_966);
and U803 (N_803,In_312,In_621);
and U804 (N_804,In_648,In_852);
nor U805 (N_805,In_292,In_393);
or U806 (N_806,In_871,In_289);
or U807 (N_807,In_786,In_411);
and U808 (N_808,In_765,In_926);
nand U809 (N_809,In_183,In_278);
and U810 (N_810,In_111,In_441);
and U811 (N_811,In_959,In_445);
nand U812 (N_812,In_193,In_305);
nand U813 (N_813,In_876,In_823);
nor U814 (N_814,In_202,In_399);
nand U815 (N_815,In_851,In_669);
nor U816 (N_816,In_391,In_612);
nand U817 (N_817,In_527,In_187);
nand U818 (N_818,In_119,In_407);
or U819 (N_819,In_993,In_224);
or U820 (N_820,In_89,In_316);
nor U821 (N_821,In_423,In_767);
and U822 (N_822,In_951,In_623);
and U823 (N_823,In_697,In_215);
or U824 (N_824,In_833,In_296);
or U825 (N_825,In_519,In_449);
or U826 (N_826,In_171,In_192);
or U827 (N_827,In_879,In_73);
nand U828 (N_828,In_34,In_28);
and U829 (N_829,In_821,In_915);
nor U830 (N_830,In_761,In_34);
and U831 (N_831,In_791,In_748);
or U832 (N_832,In_451,In_251);
nor U833 (N_833,In_775,In_29);
nand U834 (N_834,In_15,In_88);
nor U835 (N_835,In_655,In_491);
or U836 (N_836,In_758,In_40);
nand U837 (N_837,In_73,In_293);
nand U838 (N_838,In_591,In_316);
nand U839 (N_839,In_608,In_754);
nand U840 (N_840,In_610,In_242);
nor U841 (N_841,In_334,In_711);
nand U842 (N_842,In_613,In_65);
and U843 (N_843,In_644,In_438);
nor U844 (N_844,In_226,In_328);
nand U845 (N_845,In_637,In_571);
or U846 (N_846,In_446,In_903);
and U847 (N_847,In_759,In_65);
nand U848 (N_848,In_597,In_787);
and U849 (N_849,In_273,In_490);
xnor U850 (N_850,In_298,In_378);
or U851 (N_851,In_37,In_490);
or U852 (N_852,In_650,In_134);
nand U853 (N_853,In_298,In_590);
or U854 (N_854,In_969,In_257);
nand U855 (N_855,In_869,In_73);
nand U856 (N_856,In_287,In_569);
or U857 (N_857,In_620,In_854);
nor U858 (N_858,In_622,In_56);
nor U859 (N_859,In_40,In_51);
and U860 (N_860,In_446,In_871);
nor U861 (N_861,In_224,In_788);
or U862 (N_862,In_96,In_874);
nor U863 (N_863,In_193,In_257);
nand U864 (N_864,In_887,In_464);
nand U865 (N_865,In_909,In_971);
nor U866 (N_866,In_824,In_833);
nor U867 (N_867,In_625,In_920);
nor U868 (N_868,In_652,In_93);
nor U869 (N_869,In_235,In_736);
nand U870 (N_870,In_623,In_850);
and U871 (N_871,In_724,In_543);
nor U872 (N_872,In_38,In_636);
nand U873 (N_873,In_532,In_7);
or U874 (N_874,In_37,In_645);
nand U875 (N_875,In_228,In_723);
and U876 (N_876,In_489,In_123);
nor U877 (N_877,In_114,In_213);
or U878 (N_878,In_697,In_746);
nand U879 (N_879,In_822,In_540);
and U880 (N_880,In_204,In_494);
nor U881 (N_881,In_252,In_223);
and U882 (N_882,In_166,In_738);
nor U883 (N_883,In_297,In_225);
nor U884 (N_884,In_285,In_943);
nor U885 (N_885,In_309,In_585);
nor U886 (N_886,In_43,In_364);
nor U887 (N_887,In_384,In_449);
nor U888 (N_888,In_3,In_117);
or U889 (N_889,In_289,In_616);
and U890 (N_890,In_674,In_732);
nor U891 (N_891,In_65,In_711);
and U892 (N_892,In_304,In_549);
nand U893 (N_893,In_919,In_466);
xnor U894 (N_894,In_77,In_521);
and U895 (N_895,In_988,In_450);
nand U896 (N_896,In_908,In_960);
nor U897 (N_897,In_47,In_729);
and U898 (N_898,In_798,In_444);
or U899 (N_899,In_25,In_525);
and U900 (N_900,In_78,In_486);
nand U901 (N_901,In_204,In_902);
or U902 (N_902,In_66,In_551);
and U903 (N_903,In_83,In_573);
or U904 (N_904,In_285,In_196);
or U905 (N_905,In_809,In_380);
nor U906 (N_906,In_786,In_876);
and U907 (N_907,In_323,In_498);
or U908 (N_908,In_295,In_109);
nand U909 (N_909,In_826,In_189);
nand U910 (N_910,In_663,In_197);
nand U911 (N_911,In_328,In_621);
nand U912 (N_912,In_622,In_187);
xnor U913 (N_913,In_944,In_132);
nand U914 (N_914,In_818,In_923);
nand U915 (N_915,In_271,In_842);
nand U916 (N_916,In_423,In_549);
nand U917 (N_917,In_544,In_403);
and U918 (N_918,In_780,In_621);
nor U919 (N_919,In_83,In_849);
and U920 (N_920,In_610,In_541);
nand U921 (N_921,In_48,In_695);
xor U922 (N_922,In_732,In_339);
or U923 (N_923,In_543,In_797);
xor U924 (N_924,In_646,In_754);
nor U925 (N_925,In_78,In_663);
and U926 (N_926,In_165,In_864);
and U927 (N_927,In_341,In_199);
nor U928 (N_928,In_730,In_395);
nor U929 (N_929,In_847,In_141);
and U930 (N_930,In_939,In_950);
and U931 (N_931,In_434,In_514);
nor U932 (N_932,In_677,In_717);
nand U933 (N_933,In_662,In_65);
nand U934 (N_934,In_173,In_201);
and U935 (N_935,In_587,In_714);
and U936 (N_936,In_334,In_52);
nand U937 (N_937,In_346,In_21);
or U938 (N_938,In_596,In_713);
or U939 (N_939,In_511,In_698);
nand U940 (N_940,In_565,In_993);
xor U941 (N_941,In_572,In_566);
or U942 (N_942,In_848,In_548);
nand U943 (N_943,In_451,In_29);
and U944 (N_944,In_523,In_16);
or U945 (N_945,In_347,In_270);
nor U946 (N_946,In_630,In_413);
nor U947 (N_947,In_67,In_799);
xor U948 (N_948,In_181,In_933);
xor U949 (N_949,In_616,In_819);
xnor U950 (N_950,In_40,In_168);
or U951 (N_951,In_358,In_552);
and U952 (N_952,In_736,In_335);
nor U953 (N_953,In_876,In_863);
and U954 (N_954,In_776,In_499);
nand U955 (N_955,In_545,In_768);
nand U956 (N_956,In_778,In_144);
nor U957 (N_957,In_389,In_314);
nor U958 (N_958,In_292,In_682);
or U959 (N_959,In_578,In_860);
and U960 (N_960,In_355,In_599);
or U961 (N_961,In_936,In_543);
nor U962 (N_962,In_706,In_159);
nand U963 (N_963,In_263,In_680);
and U964 (N_964,In_803,In_551);
nor U965 (N_965,In_21,In_588);
and U966 (N_966,In_843,In_549);
nor U967 (N_967,In_373,In_634);
nand U968 (N_968,In_688,In_702);
or U969 (N_969,In_971,In_921);
nand U970 (N_970,In_255,In_709);
or U971 (N_971,In_583,In_775);
nor U972 (N_972,In_217,In_328);
and U973 (N_973,In_299,In_49);
xor U974 (N_974,In_856,In_345);
and U975 (N_975,In_94,In_19);
nand U976 (N_976,In_550,In_120);
xnor U977 (N_977,In_753,In_425);
and U978 (N_978,In_497,In_303);
nor U979 (N_979,In_629,In_213);
nand U980 (N_980,In_141,In_908);
nor U981 (N_981,In_318,In_475);
nor U982 (N_982,In_481,In_175);
nand U983 (N_983,In_866,In_55);
nor U984 (N_984,In_798,In_125);
and U985 (N_985,In_574,In_728);
or U986 (N_986,In_257,In_448);
xor U987 (N_987,In_75,In_733);
or U988 (N_988,In_929,In_659);
xor U989 (N_989,In_204,In_549);
nor U990 (N_990,In_930,In_348);
or U991 (N_991,In_141,In_423);
nand U992 (N_992,In_459,In_289);
or U993 (N_993,In_554,In_464);
or U994 (N_994,In_172,In_205);
or U995 (N_995,In_239,In_222);
or U996 (N_996,In_693,In_788);
nor U997 (N_997,In_807,In_46);
nor U998 (N_998,In_738,In_828);
nand U999 (N_999,In_370,In_284);
and U1000 (N_1000,In_696,In_246);
nor U1001 (N_1001,In_834,In_621);
or U1002 (N_1002,In_219,In_578);
and U1003 (N_1003,In_738,In_173);
or U1004 (N_1004,In_403,In_619);
nand U1005 (N_1005,In_310,In_298);
and U1006 (N_1006,In_740,In_643);
nor U1007 (N_1007,In_747,In_217);
and U1008 (N_1008,In_90,In_516);
nand U1009 (N_1009,In_316,In_291);
nor U1010 (N_1010,In_867,In_87);
or U1011 (N_1011,In_837,In_954);
and U1012 (N_1012,In_334,In_185);
and U1013 (N_1013,In_775,In_727);
and U1014 (N_1014,In_964,In_274);
and U1015 (N_1015,In_234,In_108);
nand U1016 (N_1016,In_791,In_98);
and U1017 (N_1017,In_921,In_727);
nand U1018 (N_1018,In_577,In_643);
nor U1019 (N_1019,In_574,In_442);
or U1020 (N_1020,In_689,In_202);
nand U1021 (N_1021,In_442,In_328);
and U1022 (N_1022,In_893,In_348);
nor U1023 (N_1023,In_136,In_915);
and U1024 (N_1024,In_561,In_575);
or U1025 (N_1025,In_65,In_381);
nor U1026 (N_1026,In_917,In_831);
or U1027 (N_1027,In_843,In_908);
nand U1028 (N_1028,In_230,In_901);
and U1029 (N_1029,In_344,In_544);
nor U1030 (N_1030,In_63,In_661);
or U1031 (N_1031,In_165,In_884);
and U1032 (N_1032,In_679,In_475);
and U1033 (N_1033,In_256,In_960);
xnor U1034 (N_1034,In_433,In_729);
nand U1035 (N_1035,In_164,In_500);
or U1036 (N_1036,In_805,In_381);
nand U1037 (N_1037,In_711,In_817);
or U1038 (N_1038,In_666,In_178);
or U1039 (N_1039,In_230,In_679);
nor U1040 (N_1040,In_364,In_771);
or U1041 (N_1041,In_191,In_210);
or U1042 (N_1042,In_987,In_251);
or U1043 (N_1043,In_367,In_382);
or U1044 (N_1044,In_506,In_900);
nand U1045 (N_1045,In_556,In_536);
xnor U1046 (N_1046,In_516,In_195);
nor U1047 (N_1047,In_557,In_204);
nand U1048 (N_1048,In_90,In_289);
or U1049 (N_1049,In_849,In_860);
or U1050 (N_1050,In_318,In_238);
and U1051 (N_1051,In_504,In_840);
or U1052 (N_1052,In_29,In_370);
xnor U1053 (N_1053,In_488,In_248);
xnor U1054 (N_1054,In_385,In_598);
nor U1055 (N_1055,In_901,In_725);
nand U1056 (N_1056,In_506,In_364);
and U1057 (N_1057,In_765,In_948);
or U1058 (N_1058,In_495,In_42);
nand U1059 (N_1059,In_657,In_659);
and U1060 (N_1060,In_530,In_997);
nand U1061 (N_1061,In_805,In_885);
and U1062 (N_1062,In_224,In_943);
nand U1063 (N_1063,In_385,In_428);
nor U1064 (N_1064,In_671,In_604);
and U1065 (N_1065,In_826,In_532);
nor U1066 (N_1066,In_928,In_727);
and U1067 (N_1067,In_236,In_775);
and U1068 (N_1068,In_769,In_395);
nor U1069 (N_1069,In_217,In_975);
nor U1070 (N_1070,In_8,In_804);
or U1071 (N_1071,In_424,In_876);
nand U1072 (N_1072,In_832,In_824);
nor U1073 (N_1073,In_964,In_97);
nor U1074 (N_1074,In_468,In_985);
or U1075 (N_1075,In_800,In_735);
and U1076 (N_1076,In_208,In_924);
and U1077 (N_1077,In_984,In_904);
and U1078 (N_1078,In_579,In_957);
nor U1079 (N_1079,In_323,In_991);
nor U1080 (N_1080,In_997,In_12);
or U1081 (N_1081,In_897,In_695);
or U1082 (N_1082,In_341,In_47);
nand U1083 (N_1083,In_980,In_584);
or U1084 (N_1084,In_335,In_492);
nand U1085 (N_1085,In_259,In_558);
nand U1086 (N_1086,In_290,In_984);
or U1087 (N_1087,In_387,In_134);
nand U1088 (N_1088,In_125,In_107);
nand U1089 (N_1089,In_239,In_508);
xnor U1090 (N_1090,In_133,In_882);
or U1091 (N_1091,In_691,In_326);
and U1092 (N_1092,In_142,In_868);
or U1093 (N_1093,In_759,In_453);
or U1094 (N_1094,In_351,In_418);
and U1095 (N_1095,In_229,In_985);
or U1096 (N_1096,In_421,In_803);
or U1097 (N_1097,In_666,In_86);
xnor U1098 (N_1098,In_894,In_599);
and U1099 (N_1099,In_723,In_292);
and U1100 (N_1100,In_116,In_647);
and U1101 (N_1101,In_418,In_992);
and U1102 (N_1102,In_690,In_448);
nor U1103 (N_1103,In_71,In_190);
or U1104 (N_1104,In_976,In_385);
or U1105 (N_1105,In_47,In_253);
and U1106 (N_1106,In_866,In_612);
or U1107 (N_1107,In_46,In_976);
nand U1108 (N_1108,In_95,In_116);
or U1109 (N_1109,In_209,In_694);
or U1110 (N_1110,In_89,In_253);
nor U1111 (N_1111,In_765,In_69);
or U1112 (N_1112,In_518,In_629);
or U1113 (N_1113,In_799,In_953);
and U1114 (N_1114,In_817,In_757);
nor U1115 (N_1115,In_165,In_784);
and U1116 (N_1116,In_110,In_464);
nor U1117 (N_1117,In_979,In_459);
nand U1118 (N_1118,In_18,In_495);
nand U1119 (N_1119,In_813,In_491);
nand U1120 (N_1120,In_237,In_499);
and U1121 (N_1121,In_232,In_30);
and U1122 (N_1122,In_735,In_552);
and U1123 (N_1123,In_664,In_838);
nand U1124 (N_1124,In_783,In_440);
nand U1125 (N_1125,In_897,In_875);
nand U1126 (N_1126,In_694,In_362);
nand U1127 (N_1127,In_780,In_710);
nor U1128 (N_1128,In_582,In_571);
nand U1129 (N_1129,In_78,In_281);
xor U1130 (N_1130,In_434,In_901);
nor U1131 (N_1131,In_6,In_352);
nand U1132 (N_1132,In_625,In_177);
or U1133 (N_1133,In_260,In_295);
xnor U1134 (N_1134,In_403,In_105);
nand U1135 (N_1135,In_426,In_790);
xnor U1136 (N_1136,In_980,In_414);
nor U1137 (N_1137,In_970,In_352);
or U1138 (N_1138,In_153,In_316);
or U1139 (N_1139,In_405,In_792);
or U1140 (N_1140,In_770,In_579);
or U1141 (N_1141,In_698,In_476);
or U1142 (N_1142,In_767,In_594);
nand U1143 (N_1143,In_408,In_953);
or U1144 (N_1144,In_750,In_815);
nand U1145 (N_1145,In_230,In_58);
nand U1146 (N_1146,In_84,In_743);
or U1147 (N_1147,In_445,In_70);
nand U1148 (N_1148,In_240,In_899);
or U1149 (N_1149,In_748,In_342);
or U1150 (N_1150,In_559,In_157);
nand U1151 (N_1151,In_909,In_108);
nand U1152 (N_1152,In_858,In_523);
and U1153 (N_1153,In_832,In_990);
or U1154 (N_1154,In_826,In_565);
nand U1155 (N_1155,In_96,In_40);
and U1156 (N_1156,In_414,In_0);
xnor U1157 (N_1157,In_556,In_347);
and U1158 (N_1158,In_94,In_755);
nand U1159 (N_1159,In_833,In_38);
xor U1160 (N_1160,In_171,In_392);
or U1161 (N_1161,In_773,In_753);
nor U1162 (N_1162,In_467,In_233);
nor U1163 (N_1163,In_560,In_61);
or U1164 (N_1164,In_306,In_206);
nand U1165 (N_1165,In_898,In_977);
nor U1166 (N_1166,In_459,In_894);
or U1167 (N_1167,In_738,In_445);
or U1168 (N_1168,In_560,In_710);
and U1169 (N_1169,In_857,In_566);
xnor U1170 (N_1170,In_620,In_246);
or U1171 (N_1171,In_517,In_450);
or U1172 (N_1172,In_276,In_851);
nand U1173 (N_1173,In_674,In_282);
nand U1174 (N_1174,In_347,In_478);
and U1175 (N_1175,In_347,In_941);
and U1176 (N_1176,In_486,In_523);
or U1177 (N_1177,In_899,In_82);
xnor U1178 (N_1178,In_652,In_766);
nor U1179 (N_1179,In_783,In_789);
nor U1180 (N_1180,In_739,In_5);
and U1181 (N_1181,In_256,In_613);
or U1182 (N_1182,In_910,In_67);
and U1183 (N_1183,In_745,In_188);
or U1184 (N_1184,In_276,In_451);
and U1185 (N_1185,In_722,In_331);
and U1186 (N_1186,In_852,In_806);
nand U1187 (N_1187,In_629,In_493);
nor U1188 (N_1188,In_224,In_997);
or U1189 (N_1189,In_974,In_726);
or U1190 (N_1190,In_812,In_731);
nor U1191 (N_1191,In_334,In_255);
and U1192 (N_1192,In_882,In_938);
nand U1193 (N_1193,In_801,In_1);
nand U1194 (N_1194,In_272,In_907);
xnor U1195 (N_1195,In_497,In_697);
nor U1196 (N_1196,In_226,In_293);
nor U1197 (N_1197,In_954,In_807);
nor U1198 (N_1198,In_458,In_938);
and U1199 (N_1199,In_973,In_318);
and U1200 (N_1200,In_214,In_708);
and U1201 (N_1201,In_467,In_445);
nor U1202 (N_1202,In_644,In_562);
or U1203 (N_1203,In_977,In_710);
nor U1204 (N_1204,In_474,In_606);
nor U1205 (N_1205,In_700,In_552);
nor U1206 (N_1206,In_668,In_599);
or U1207 (N_1207,In_845,In_627);
nor U1208 (N_1208,In_352,In_863);
and U1209 (N_1209,In_221,In_307);
nand U1210 (N_1210,In_923,In_74);
or U1211 (N_1211,In_467,In_872);
nand U1212 (N_1212,In_164,In_156);
nor U1213 (N_1213,In_262,In_789);
nor U1214 (N_1214,In_718,In_561);
xor U1215 (N_1215,In_553,In_503);
and U1216 (N_1216,In_763,In_673);
nor U1217 (N_1217,In_73,In_881);
and U1218 (N_1218,In_344,In_921);
xor U1219 (N_1219,In_85,In_666);
xor U1220 (N_1220,In_711,In_214);
or U1221 (N_1221,In_955,In_769);
nand U1222 (N_1222,In_255,In_260);
nor U1223 (N_1223,In_797,In_826);
and U1224 (N_1224,In_851,In_245);
nand U1225 (N_1225,In_371,In_958);
or U1226 (N_1226,In_968,In_151);
nand U1227 (N_1227,In_476,In_183);
and U1228 (N_1228,In_330,In_106);
nand U1229 (N_1229,In_762,In_111);
or U1230 (N_1230,In_44,In_437);
nor U1231 (N_1231,In_68,In_548);
nand U1232 (N_1232,In_339,In_574);
and U1233 (N_1233,In_977,In_150);
or U1234 (N_1234,In_968,In_675);
and U1235 (N_1235,In_403,In_690);
and U1236 (N_1236,In_746,In_633);
nand U1237 (N_1237,In_200,In_930);
nand U1238 (N_1238,In_933,In_613);
and U1239 (N_1239,In_222,In_220);
nor U1240 (N_1240,In_210,In_270);
nor U1241 (N_1241,In_284,In_474);
or U1242 (N_1242,In_544,In_905);
nor U1243 (N_1243,In_471,In_402);
nor U1244 (N_1244,In_366,In_736);
or U1245 (N_1245,In_663,In_447);
nor U1246 (N_1246,In_993,In_915);
nand U1247 (N_1247,In_928,In_594);
and U1248 (N_1248,In_700,In_308);
and U1249 (N_1249,In_273,In_132);
nand U1250 (N_1250,In_20,In_120);
nand U1251 (N_1251,In_377,In_586);
nand U1252 (N_1252,In_418,In_293);
nand U1253 (N_1253,In_785,In_525);
or U1254 (N_1254,In_324,In_66);
xor U1255 (N_1255,In_388,In_444);
nand U1256 (N_1256,In_14,In_747);
nand U1257 (N_1257,In_40,In_354);
xnor U1258 (N_1258,In_218,In_377);
nand U1259 (N_1259,In_776,In_197);
or U1260 (N_1260,In_815,In_466);
and U1261 (N_1261,In_270,In_123);
xor U1262 (N_1262,In_266,In_15);
and U1263 (N_1263,In_272,In_952);
xnor U1264 (N_1264,In_273,In_503);
or U1265 (N_1265,In_908,In_594);
and U1266 (N_1266,In_987,In_556);
nor U1267 (N_1267,In_32,In_422);
or U1268 (N_1268,In_875,In_104);
xnor U1269 (N_1269,In_347,In_33);
and U1270 (N_1270,In_387,In_952);
xnor U1271 (N_1271,In_551,In_496);
and U1272 (N_1272,In_747,In_200);
nor U1273 (N_1273,In_866,In_51);
nor U1274 (N_1274,In_888,In_860);
and U1275 (N_1275,In_413,In_838);
nand U1276 (N_1276,In_393,In_370);
nor U1277 (N_1277,In_305,In_695);
or U1278 (N_1278,In_437,In_181);
or U1279 (N_1279,In_83,In_245);
or U1280 (N_1280,In_667,In_528);
nand U1281 (N_1281,In_440,In_324);
or U1282 (N_1282,In_85,In_392);
nand U1283 (N_1283,In_107,In_681);
or U1284 (N_1284,In_545,In_378);
and U1285 (N_1285,In_873,In_308);
and U1286 (N_1286,In_487,In_374);
nand U1287 (N_1287,In_503,In_459);
and U1288 (N_1288,In_277,In_453);
or U1289 (N_1289,In_846,In_437);
nor U1290 (N_1290,In_827,In_307);
nor U1291 (N_1291,In_805,In_148);
xor U1292 (N_1292,In_937,In_368);
nor U1293 (N_1293,In_10,In_608);
or U1294 (N_1294,In_191,In_378);
nor U1295 (N_1295,In_47,In_456);
or U1296 (N_1296,In_975,In_101);
or U1297 (N_1297,In_357,In_351);
or U1298 (N_1298,In_10,In_973);
and U1299 (N_1299,In_857,In_536);
or U1300 (N_1300,In_656,In_180);
nor U1301 (N_1301,In_974,In_586);
or U1302 (N_1302,In_34,In_391);
or U1303 (N_1303,In_452,In_487);
and U1304 (N_1304,In_820,In_818);
nor U1305 (N_1305,In_316,In_927);
and U1306 (N_1306,In_89,In_823);
nor U1307 (N_1307,In_867,In_350);
nor U1308 (N_1308,In_992,In_953);
nor U1309 (N_1309,In_236,In_684);
or U1310 (N_1310,In_734,In_464);
or U1311 (N_1311,In_999,In_390);
nor U1312 (N_1312,In_660,In_384);
or U1313 (N_1313,In_724,In_538);
nor U1314 (N_1314,In_478,In_553);
or U1315 (N_1315,In_547,In_398);
and U1316 (N_1316,In_404,In_945);
nand U1317 (N_1317,In_925,In_526);
nand U1318 (N_1318,In_611,In_887);
nor U1319 (N_1319,In_628,In_398);
nor U1320 (N_1320,In_271,In_637);
or U1321 (N_1321,In_57,In_100);
and U1322 (N_1322,In_653,In_674);
or U1323 (N_1323,In_426,In_764);
or U1324 (N_1324,In_750,In_97);
nor U1325 (N_1325,In_367,In_993);
nor U1326 (N_1326,In_225,In_101);
and U1327 (N_1327,In_407,In_153);
or U1328 (N_1328,In_701,In_782);
nand U1329 (N_1329,In_569,In_249);
and U1330 (N_1330,In_787,In_259);
and U1331 (N_1331,In_782,In_8);
or U1332 (N_1332,In_341,In_720);
xnor U1333 (N_1333,In_944,In_178);
or U1334 (N_1334,In_880,In_709);
or U1335 (N_1335,In_445,In_449);
or U1336 (N_1336,In_426,In_29);
nand U1337 (N_1337,In_850,In_636);
nor U1338 (N_1338,In_555,In_932);
nand U1339 (N_1339,In_137,In_185);
xor U1340 (N_1340,In_497,In_793);
nor U1341 (N_1341,In_502,In_192);
or U1342 (N_1342,In_690,In_560);
xor U1343 (N_1343,In_645,In_283);
or U1344 (N_1344,In_346,In_973);
and U1345 (N_1345,In_742,In_563);
or U1346 (N_1346,In_678,In_346);
nand U1347 (N_1347,In_275,In_968);
nor U1348 (N_1348,In_204,In_991);
and U1349 (N_1349,In_116,In_501);
nand U1350 (N_1350,In_387,In_360);
nor U1351 (N_1351,In_561,In_957);
or U1352 (N_1352,In_672,In_950);
or U1353 (N_1353,In_231,In_701);
and U1354 (N_1354,In_380,In_18);
nor U1355 (N_1355,In_7,In_54);
xnor U1356 (N_1356,In_484,In_738);
or U1357 (N_1357,In_788,In_103);
nor U1358 (N_1358,In_151,In_355);
and U1359 (N_1359,In_544,In_88);
or U1360 (N_1360,In_772,In_785);
and U1361 (N_1361,In_286,In_292);
nand U1362 (N_1362,In_365,In_902);
and U1363 (N_1363,In_811,In_784);
or U1364 (N_1364,In_978,In_892);
nor U1365 (N_1365,In_659,In_425);
or U1366 (N_1366,In_582,In_367);
and U1367 (N_1367,In_797,In_134);
nor U1368 (N_1368,In_516,In_207);
nand U1369 (N_1369,In_906,In_769);
nor U1370 (N_1370,In_819,In_698);
xnor U1371 (N_1371,In_650,In_494);
nor U1372 (N_1372,In_36,In_259);
nand U1373 (N_1373,In_973,In_950);
nor U1374 (N_1374,In_702,In_352);
nor U1375 (N_1375,In_812,In_105);
and U1376 (N_1376,In_742,In_531);
nand U1377 (N_1377,In_372,In_870);
or U1378 (N_1378,In_696,In_812);
nor U1379 (N_1379,In_86,In_975);
xor U1380 (N_1380,In_896,In_368);
nor U1381 (N_1381,In_965,In_304);
xor U1382 (N_1382,In_685,In_655);
and U1383 (N_1383,In_316,In_98);
nand U1384 (N_1384,In_213,In_67);
xnor U1385 (N_1385,In_216,In_86);
nor U1386 (N_1386,In_521,In_132);
nand U1387 (N_1387,In_665,In_443);
xor U1388 (N_1388,In_136,In_268);
nor U1389 (N_1389,In_337,In_997);
or U1390 (N_1390,In_760,In_516);
nor U1391 (N_1391,In_593,In_977);
nor U1392 (N_1392,In_137,In_402);
nor U1393 (N_1393,In_596,In_273);
and U1394 (N_1394,In_820,In_3);
nand U1395 (N_1395,In_313,In_711);
nor U1396 (N_1396,In_327,In_699);
and U1397 (N_1397,In_734,In_415);
or U1398 (N_1398,In_730,In_850);
or U1399 (N_1399,In_454,In_62);
and U1400 (N_1400,In_257,In_261);
and U1401 (N_1401,In_338,In_534);
and U1402 (N_1402,In_174,In_246);
xor U1403 (N_1403,In_31,In_697);
and U1404 (N_1404,In_305,In_677);
or U1405 (N_1405,In_908,In_229);
and U1406 (N_1406,In_419,In_302);
and U1407 (N_1407,In_577,In_735);
or U1408 (N_1408,In_818,In_466);
or U1409 (N_1409,In_581,In_766);
or U1410 (N_1410,In_30,In_38);
or U1411 (N_1411,In_132,In_942);
and U1412 (N_1412,In_351,In_286);
nor U1413 (N_1413,In_665,In_671);
and U1414 (N_1414,In_418,In_788);
nor U1415 (N_1415,In_93,In_952);
nand U1416 (N_1416,In_185,In_697);
or U1417 (N_1417,In_73,In_141);
or U1418 (N_1418,In_519,In_643);
or U1419 (N_1419,In_498,In_833);
and U1420 (N_1420,In_57,In_9);
nand U1421 (N_1421,In_426,In_243);
or U1422 (N_1422,In_945,In_98);
nor U1423 (N_1423,In_137,In_246);
nand U1424 (N_1424,In_923,In_160);
and U1425 (N_1425,In_80,In_927);
nor U1426 (N_1426,In_854,In_986);
and U1427 (N_1427,In_459,In_552);
or U1428 (N_1428,In_735,In_64);
xnor U1429 (N_1429,In_625,In_655);
nor U1430 (N_1430,In_738,In_427);
nor U1431 (N_1431,In_453,In_367);
nor U1432 (N_1432,In_998,In_178);
nand U1433 (N_1433,In_588,In_837);
xor U1434 (N_1434,In_225,In_827);
nand U1435 (N_1435,In_415,In_332);
nor U1436 (N_1436,In_156,In_837);
and U1437 (N_1437,In_631,In_847);
xor U1438 (N_1438,In_407,In_531);
and U1439 (N_1439,In_33,In_74);
nor U1440 (N_1440,In_733,In_942);
nand U1441 (N_1441,In_446,In_484);
nor U1442 (N_1442,In_463,In_765);
or U1443 (N_1443,In_715,In_497);
and U1444 (N_1444,In_627,In_51);
or U1445 (N_1445,In_714,In_991);
nor U1446 (N_1446,In_747,In_290);
and U1447 (N_1447,In_778,In_520);
nand U1448 (N_1448,In_269,In_424);
nor U1449 (N_1449,In_273,In_46);
and U1450 (N_1450,In_288,In_698);
nand U1451 (N_1451,In_435,In_614);
or U1452 (N_1452,In_240,In_904);
or U1453 (N_1453,In_990,In_714);
and U1454 (N_1454,In_890,In_612);
nand U1455 (N_1455,In_165,In_879);
and U1456 (N_1456,In_663,In_808);
and U1457 (N_1457,In_686,In_887);
and U1458 (N_1458,In_483,In_332);
nor U1459 (N_1459,In_580,In_82);
nor U1460 (N_1460,In_512,In_177);
or U1461 (N_1461,In_706,In_135);
nor U1462 (N_1462,In_523,In_632);
and U1463 (N_1463,In_11,In_565);
nand U1464 (N_1464,In_886,In_713);
or U1465 (N_1465,In_629,In_878);
or U1466 (N_1466,In_648,In_685);
nand U1467 (N_1467,In_602,In_685);
and U1468 (N_1468,In_366,In_75);
xor U1469 (N_1469,In_269,In_260);
and U1470 (N_1470,In_525,In_856);
and U1471 (N_1471,In_798,In_139);
nand U1472 (N_1472,In_789,In_702);
nand U1473 (N_1473,In_168,In_220);
nand U1474 (N_1474,In_345,In_484);
or U1475 (N_1475,In_928,In_870);
and U1476 (N_1476,In_131,In_125);
nand U1477 (N_1477,In_112,In_782);
xnor U1478 (N_1478,In_456,In_713);
and U1479 (N_1479,In_752,In_190);
nor U1480 (N_1480,In_602,In_443);
nand U1481 (N_1481,In_192,In_205);
nand U1482 (N_1482,In_45,In_665);
and U1483 (N_1483,In_235,In_51);
or U1484 (N_1484,In_264,In_591);
and U1485 (N_1485,In_114,In_709);
nand U1486 (N_1486,In_133,In_249);
or U1487 (N_1487,In_568,In_62);
or U1488 (N_1488,In_532,In_570);
nand U1489 (N_1489,In_885,In_138);
or U1490 (N_1490,In_536,In_202);
nand U1491 (N_1491,In_271,In_448);
and U1492 (N_1492,In_132,In_81);
nor U1493 (N_1493,In_715,In_130);
nand U1494 (N_1494,In_530,In_576);
nand U1495 (N_1495,In_529,In_739);
or U1496 (N_1496,In_913,In_675);
or U1497 (N_1497,In_877,In_612);
or U1498 (N_1498,In_326,In_543);
and U1499 (N_1499,In_613,In_457);
and U1500 (N_1500,In_863,In_506);
or U1501 (N_1501,In_667,In_508);
and U1502 (N_1502,In_616,In_1);
or U1503 (N_1503,In_10,In_229);
nor U1504 (N_1504,In_583,In_475);
or U1505 (N_1505,In_683,In_505);
and U1506 (N_1506,In_258,In_685);
or U1507 (N_1507,In_446,In_43);
nor U1508 (N_1508,In_645,In_935);
nor U1509 (N_1509,In_340,In_887);
and U1510 (N_1510,In_579,In_712);
nor U1511 (N_1511,In_381,In_106);
nor U1512 (N_1512,In_801,In_986);
and U1513 (N_1513,In_240,In_280);
nor U1514 (N_1514,In_961,In_316);
or U1515 (N_1515,In_957,In_466);
or U1516 (N_1516,In_636,In_87);
and U1517 (N_1517,In_500,In_799);
or U1518 (N_1518,In_606,In_742);
and U1519 (N_1519,In_744,In_573);
nor U1520 (N_1520,In_635,In_763);
and U1521 (N_1521,In_997,In_496);
or U1522 (N_1522,In_789,In_843);
nor U1523 (N_1523,In_432,In_580);
nor U1524 (N_1524,In_693,In_426);
or U1525 (N_1525,In_969,In_763);
or U1526 (N_1526,In_273,In_180);
nand U1527 (N_1527,In_684,In_530);
and U1528 (N_1528,In_588,In_365);
nor U1529 (N_1529,In_777,In_458);
nor U1530 (N_1530,In_346,In_703);
nand U1531 (N_1531,In_254,In_935);
and U1532 (N_1532,In_449,In_509);
and U1533 (N_1533,In_351,In_54);
nand U1534 (N_1534,In_517,In_411);
or U1535 (N_1535,In_342,In_106);
and U1536 (N_1536,In_252,In_340);
nand U1537 (N_1537,In_184,In_382);
or U1538 (N_1538,In_517,In_505);
or U1539 (N_1539,In_336,In_14);
nand U1540 (N_1540,In_688,In_614);
or U1541 (N_1541,In_96,In_94);
nand U1542 (N_1542,In_388,In_670);
xnor U1543 (N_1543,In_807,In_368);
or U1544 (N_1544,In_650,In_739);
and U1545 (N_1545,In_70,In_81);
or U1546 (N_1546,In_835,In_803);
nand U1547 (N_1547,In_862,In_285);
xor U1548 (N_1548,In_160,In_47);
or U1549 (N_1549,In_567,In_938);
and U1550 (N_1550,In_511,In_874);
or U1551 (N_1551,In_596,In_884);
and U1552 (N_1552,In_834,In_737);
and U1553 (N_1553,In_805,In_167);
or U1554 (N_1554,In_902,In_910);
xnor U1555 (N_1555,In_623,In_403);
or U1556 (N_1556,In_78,In_731);
or U1557 (N_1557,In_819,In_977);
or U1558 (N_1558,In_182,In_777);
or U1559 (N_1559,In_862,In_144);
nand U1560 (N_1560,In_711,In_58);
and U1561 (N_1561,In_472,In_132);
or U1562 (N_1562,In_316,In_939);
or U1563 (N_1563,In_628,In_734);
or U1564 (N_1564,In_749,In_338);
or U1565 (N_1565,In_49,In_471);
nor U1566 (N_1566,In_986,In_79);
nor U1567 (N_1567,In_702,In_470);
or U1568 (N_1568,In_241,In_285);
or U1569 (N_1569,In_583,In_334);
nor U1570 (N_1570,In_723,In_684);
nor U1571 (N_1571,In_621,In_730);
nor U1572 (N_1572,In_655,In_799);
nand U1573 (N_1573,In_84,In_284);
or U1574 (N_1574,In_516,In_341);
nor U1575 (N_1575,In_126,In_281);
or U1576 (N_1576,In_692,In_673);
and U1577 (N_1577,In_613,In_282);
or U1578 (N_1578,In_873,In_947);
and U1579 (N_1579,In_744,In_504);
nor U1580 (N_1580,In_288,In_874);
nand U1581 (N_1581,In_90,In_448);
and U1582 (N_1582,In_7,In_888);
and U1583 (N_1583,In_798,In_704);
and U1584 (N_1584,In_416,In_724);
or U1585 (N_1585,In_370,In_246);
nor U1586 (N_1586,In_288,In_536);
or U1587 (N_1587,In_997,In_628);
and U1588 (N_1588,In_705,In_389);
nand U1589 (N_1589,In_862,In_63);
or U1590 (N_1590,In_451,In_765);
and U1591 (N_1591,In_298,In_337);
or U1592 (N_1592,In_371,In_5);
and U1593 (N_1593,In_151,In_448);
nor U1594 (N_1594,In_16,In_721);
nor U1595 (N_1595,In_158,In_360);
nand U1596 (N_1596,In_485,In_223);
nor U1597 (N_1597,In_117,In_85);
or U1598 (N_1598,In_473,In_669);
and U1599 (N_1599,In_461,In_520);
or U1600 (N_1600,In_898,In_110);
nor U1601 (N_1601,In_455,In_306);
nor U1602 (N_1602,In_42,In_297);
or U1603 (N_1603,In_832,In_294);
nor U1604 (N_1604,In_378,In_34);
and U1605 (N_1605,In_910,In_906);
nand U1606 (N_1606,In_558,In_25);
and U1607 (N_1607,In_690,In_513);
or U1608 (N_1608,In_799,In_566);
or U1609 (N_1609,In_337,In_598);
or U1610 (N_1610,In_610,In_457);
nor U1611 (N_1611,In_792,In_50);
nor U1612 (N_1612,In_950,In_476);
nand U1613 (N_1613,In_686,In_437);
nor U1614 (N_1614,In_66,In_275);
nor U1615 (N_1615,In_624,In_230);
nor U1616 (N_1616,In_165,In_669);
or U1617 (N_1617,In_429,In_270);
nor U1618 (N_1618,In_857,In_483);
nand U1619 (N_1619,In_369,In_618);
nand U1620 (N_1620,In_341,In_604);
and U1621 (N_1621,In_352,In_275);
and U1622 (N_1622,In_392,In_73);
nor U1623 (N_1623,In_573,In_423);
or U1624 (N_1624,In_70,In_203);
and U1625 (N_1625,In_800,In_518);
and U1626 (N_1626,In_599,In_48);
or U1627 (N_1627,In_871,In_132);
nand U1628 (N_1628,In_693,In_73);
xnor U1629 (N_1629,In_674,In_777);
nor U1630 (N_1630,In_928,In_645);
or U1631 (N_1631,In_229,In_626);
nand U1632 (N_1632,In_849,In_45);
or U1633 (N_1633,In_156,In_877);
and U1634 (N_1634,In_6,In_538);
or U1635 (N_1635,In_2,In_462);
nand U1636 (N_1636,In_471,In_597);
nand U1637 (N_1637,In_94,In_292);
nand U1638 (N_1638,In_490,In_746);
xnor U1639 (N_1639,In_257,In_470);
or U1640 (N_1640,In_620,In_972);
and U1641 (N_1641,In_486,In_809);
nor U1642 (N_1642,In_347,In_827);
and U1643 (N_1643,In_208,In_373);
nand U1644 (N_1644,In_869,In_804);
or U1645 (N_1645,In_851,In_595);
nor U1646 (N_1646,In_79,In_609);
or U1647 (N_1647,In_609,In_338);
or U1648 (N_1648,In_86,In_180);
nand U1649 (N_1649,In_443,In_424);
and U1650 (N_1650,In_103,In_386);
or U1651 (N_1651,In_368,In_154);
nand U1652 (N_1652,In_668,In_6);
and U1653 (N_1653,In_2,In_765);
and U1654 (N_1654,In_965,In_564);
nor U1655 (N_1655,In_374,In_757);
nand U1656 (N_1656,In_453,In_741);
nor U1657 (N_1657,In_96,In_621);
or U1658 (N_1658,In_654,In_0);
nor U1659 (N_1659,In_267,In_227);
or U1660 (N_1660,In_14,In_295);
and U1661 (N_1661,In_404,In_699);
nand U1662 (N_1662,In_423,In_850);
nand U1663 (N_1663,In_388,In_666);
or U1664 (N_1664,In_933,In_816);
nor U1665 (N_1665,In_79,In_831);
and U1666 (N_1666,In_82,In_693);
or U1667 (N_1667,In_771,In_561);
and U1668 (N_1668,In_611,In_750);
or U1669 (N_1669,In_891,In_800);
nor U1670 (N_1670,In_119,In_412);
or U1671 (N_1671,In_387,In_159);
nand U1672 (N_1672,In_212,In_602);
nor U1673 (N_1673,In_513,In_575);
or U1674 (N_1674,In_308,In_444);
nor U1675 (N_1675,In_664,In_990);
or U1676 (N_1676,In_44,In_989);
nand U1677 (N_1677,In_411,In_137);
or U1678 (N_1678,In_834,In_689);
nor U1679 (N_1679,In_912,In_45);
and U1680 (N_1680,In_816,In_909);
and U1681 (N_1681,In_90,In_597);
nor U1682 (N_1682,In_252,In_824);
and U1683 (N_1683,In_771,In_929);
xor U1684 (N_1684,In_274,In_623);
nand U1685 (N_1685,In_183,In_514);
or U1686 (N_1686,In_542,In_134);
nand U1687 (N_1687,In_73,In_647);
nand U1688 (N_1688,In_446,In_855);
or U1689 (N_1689,In_793,In_588);
or U1690 (N_1690,In_567,In_587);
or U1691 (N_1691,In_760,In_598);
and U1692 (N_1692,In_305,In_107);
or U1693 (N_1693,In_883,In_570);
nor U1694 (N_1694,In_15,In_898);
or U1695 (N_1695,In_108,In_993);
xor U1696 (N_1696,In_313,In_247);
nand U1697 (N_1697,In_17,In_949);
and U1698 (N_1698,In_777,In_606);
and U1699 (N_1699,In_285,In_989);
or U1700 (N_1700,In_72,In_585);
nor U1701 (N_1701,In_806,In_744);
or U1702 (N_1702,In_779,In_542);
and U1703 (N_1703,In_802,In_546);
nand U1704 (N_1704,In_843,In_617);
xor U1705 (N_1705,In_648,In_228);
and U1706 (N_1706,In_894,In_910);
nand U1707 (N_1707,In_228,In_583);
or U1708 (N_1708,In_896,In_408);
and U1709 (N_1709,In_944,In_445);
and U1710 (N_1710,In_560,In_439);
and U1711 (N_1711,In_300,In_927);
nor U1712 (N_1712,In_917,In_859);
and U1713 (N_1713,In_641,In_750);
or U1714 (N_1714,In_665,In_660);
and U1715 (N_1715,In_832,In_611);
nor U1716 (N_1716,In_772,In_546);
and U1717 (N_1717,In_617,In_669);
or U1718 (N_1718,In_349,In_118);
and U1719 (N_1719,In_978,In_711);
and U1720 (N_1720,In_434,In_303);
or U1721 (N_1721,In_515,In_541);
nor U1722 (N_1722,In_877,In_861);
and U1723 (N_1723,In_760,In_399);
or U1724 (N_1724,In_956,In_355);
or U1725 (N_1725,In_433,In_581);
nor U1726 (N_1726,In_66,In_441);
or U1727 (N_1727,In_313,In_866);
and U1728 (N_1728,In_96,In_572);
nor U1729 (N_1729,In_279,In_778);
nand U1730 (N_1730,In_202,In_116);
or U1731 (N_1731,In_548,In_118);
or U1732 (N_1732,In_688,In_419);
or U1733 (N_1733,In_237,In_759);
or U1734 (N_1734,In_119,In_169);
nand U1735 (N_1735,In_215,In_904);
nor U1736 (N_1736,In_740,In_524);
and U1737 (N_1737,In_369,In_860);
or U1738 (N_1738,In_65,In_284);
or U1739 (N_1739,In_350,In_230);
and U1740 (N_1740,In_454,In_482);
nor U1741 (N_1741,In_922,In_33);
nand U1742 (N_1742,In_778,In_560);
or U1743 (N_1743,In_743,In_318);
nand U1744 (N_1744,In_8,In_533);
nand U1745 (N_1745,In_328,In_846);
nand U1746 (N_1746,In_622,In_380);
and U1747 (N_1747,In_657,In_930);
or U1748 (N_1748,In_500,In_243);
and U1749 (N_1749,In_541,In_944);
nor U1750 (N_1750,In_956,In_460);
or U1751 (N_1751,In_820,In_38);
nand U1752 (N_1752,In_246,In_655);
and U1753 (N_1753,In_215,In_854);
or U1754 (N_1754,In_607,In_700);
nor U1755 (N_1755,In_540,In_954);
and U1756 (N_1756,In_38,In_588);
nand U1757 (N_1757,In_192,In_773);
nand U1758 (N_1758,In_77,In_820);
nor U1759 (N_1759,In_109,In_392);
nand U1760 (N_1760,In_310,In_369);
xor U1761 (N_1761,In_277,In_639);
and U1762 (N_1762,In_444,In_690);
nand U1763 (N_1763,In_209,In_855);
nor U1764 (N_1764,In_725,In_6);
nor U1765 (N_1765,In_511,In_937);
nor U1766 (N_1766,In_332,In_768);
or U1767 (N_1767,In_432,In_126);
and U1768 (N_1768,In_336,In_454);
or U1769 (N_1769,In_981,In_3);
or U1770 (N_1770,In_436,In_278);
or U1771 (N_1771,In_199,In_455);
and U1772 (N_1772,In_826,In_128);
nor U1773 (N_1773,In_345,In_158);
nand U1774 (N_1774,In_148,In_149);
and U1775 (N_1775,In_141,In_974);
nor U1776 (N_1776,In_831,In_272);
or U1777 (N_1777,In_203,In_31);
or U1778 (N_1778,In_787,In_958);
nor U1779 (N_1779,In_882,In_711);
nand U1780 (N_1780,In_87,In_751);
nand U1781 (N_1781,In_941,In_975);
nand U1782 (N_1782,In_768,In_91);
nand U1783 (N_1783,In_601,In_715);
nor U1784 (N_1784,In_609,In_584);
and U1785 (N_1785,In_616,In_760);
and U1786 (N_1786,In_657,In_270);
nand U1787 (N_1787,In_684,In_533);
or U1788 (N_1788,In_10,In_947);
nand U1789 (N_1789,In_34,In_630);
nor U1790 (N_1790,In_369,In_621);
and U1791 (N_1791,In_82,In_221);
and U1792 (N_1792,In_881,In_247);
or U1793 (N_1793,In_137,In_947);
or U1794 (N_1794,In_84,In_397);
nor U1795 (N_1795,In_999,In_631);
nand U1796 (N_1796,In_832,In_146);
nand U1797 (N_1797,In_755,In_151);
nand U1798 (N_1798,In_892,In_814);
nand U1799 (N_1799,In_374,In_729);
and U1800 (N_1800,In_804,In_510);
nor U1801 (N_1801,In_262,In_364);
or U1802 (N_1802,In_684,In_837);
and U1803 (N_1803,In_24,In_863);
nand U1804 (N_1804,In_512,In_881);
or U1805 (N_1805,In_40,In_85);
nor U1806 (N_1806,In_717,In_36);
or U1807 (N_1807,In_188,In_437);
and U1808 (N_1808,In_64,In_148);
or U1809 (N_1809,In_398,In_917);
nor U1810 (N_1810,In_751,In_53);
nand U1811 (N_1811,In_836,In_548);
or U1812 (N_1812,In_729,In_604);
nand U1813 (N_1813,In_210,In_570);
nor U1814 (N_1814,In_991,In_224);
nand U1815 (N_1815,In_827,In_270);
and U1816 (N_1816,In_790,In_392);
and U1817 (N_1817,In_399,In_514);
nor U1818 (N_1818,In_810,In_718);
nand U1819 (N_1819,In_31,In_560);
nor U1820 (N_1820,In_989,In_253);
nand U1821 (N_1821,In_477,In_949);
or U1822 (N_1822,In_115,In_181);
and U1823 (N_1823,In_242,In_86);
and U1824 (N_1824,In_555,In_478);
or U1825 (N_1825,In_218,In_318);
and U1826 (N_1826,In_537,In_39);
and U1827 (N_1827,In_916,In_540);
nand U1828 (N_1828,In_640,In_591);
nand U1829 (N_1829,In_57,In_25);
xor U1830 (N_1830,In_29,In_128);
nor U1831 (N_1831,In_863,In_921);
and U1832 (N_1832,In_281,In_108);
and U1833 (N_1833,In_783,In_29);
nand U1834 (N_1834,In_413,In_119);
nand U1835 (N_1835,In_121,In_812);
nor U1836 (N_1836,In_406,In_713);
and U1837 (N_1837,In_999,In_208);
and U1838 (N_1838,In_632,In_145);
nand U1839 (N_1839,In_309,In_559);
nand U1840 (N_1840,In_645,In_281);
and U1841 (N_1841,In_973,In_110);
nand U1842 (N_1842,In_886,In_414);
nand U1843 (N_1843,In_407,In_206);
nor U1844 (N_1844,In_274,In_841);
or U1845 (N_1845,In_918,In_394);
nor U1846 (N_1846,In_80,In_88);
and U1847 (N_1847,In_431,In_983);
nand U1848 (N_1848,In_553,In_56);
nand U1849 (N_1849,In_546,In_15);
or U1850 (N_1850,In_181,In_134);
or U1851 (N_1851,In_875,In_749);
or U1852 (N_1852,In_976,In_227);
or U1853 (N_1853,In_841,In_818);
or U1854 (N_1854,In_97,In_299);
nand U1855 (N_1855,In_404,In_673);
xor U1856 (N_1856,In_920,In_586);
or U1857 (N_1857,In_804,In_962);
xnor U1858 (N_1858,In_738,In_425);
or U1859 (N_1859,In_788,In_740);
nand U1860 (N_1860,In_241,In_516);
or U1861 (N_1861,In_942,In_311);
or U1862 (N_1862,In_43,In_543);
or U1863 (N_1863,In_101,In_673);
and U1864 (N_1864,In_236,In_278);
nand U1865 (N_1865,In_610,In_884);
or U1866 (N_1866,In_736,In_611);
nor U1867 (N_1867,In_51,In_80);
and U1868 (N_1868,In_934,In_714);
nand U1869 (N_1869,In_240,In_563);
or U1870 (N_1870,In_822,In_902);
nor U1871 (N_1871,In_489,In_998);
nand U1872 (N_1872,In_494,In_934);
and U1873 (N_1873,In_890,In_121);
and U1874 (N_1874,In_332,In_351);
nor U1875 (N_1875,In_848,In_507);
and U1876 (N_1876,In_801,In_794);
nand U1877 (N_1877,In_436,In_34);
nand U1878 (N_1878,In_63,In_104);
and U1879 (N_1879,In_716,In_44);
and U1880 (N_1880,In_87,In_417);
nor U1881 (N_1881,In_784,In_96);
and U1882 (N_1882,In_558,In_165);
or U1883 (N_1883,In_964,In_181);
or U1884 (N_1884,In_713,In_600);
nor U1885 (N_1885,In_770,In_889);
nand U1886 (N_1886,In_832,In_65);
nand U1887 (N_1887,In_712,In_225);
nor U1888 (N_1888,In_410,In_351);
nor U1889 (N_1889,In_502,In_890);
or U1890 (N_1890,In_106,In_870);
nand U1891 (N_1891,In_812,In_645);
or U1892 (N_1892,In_435,In_245);
or U1893 (N_1893,In_379,In_535);
and U1894 (N_1894,In_327,In_677);
and U1895 (N_1895,In_468,In_829);
and U1896 (N_1896,In_360,In_823);
or U1897 (N_1897,In_980,In_339);
or U1898 (N_1898,In_934,In_89);
nor U1899 (N_1899,In_728,In_907);
or U1900 (N_1900,In_993,In_0);
and U1901 (N_1901,In_957,In_14);
or U1902 (N_1902,In_858,In_169);
nor U1903 (N_1903,In_336,In_745);
nand U1904 (N_1904,In_606,In_584);
and U1905 (N_1905,In_945,In_333);
and U1906 (N_1906,In_846,In_314);
nand U1907 (N_1907,In_766,In_568);
nor U1908 (N_1908,In_527,In_737);
or U1909 (N_1909,In_788,In_236);
or U1910 (N_1910,In_807,In_415);
and U1911 (N_1911,In_748,In_489);
and U1912 (N_1912,In_784,In_444);
or U1913 (N_1913,In_131,In_501);
nand U1914 (N_1914,In_327,In_137);
and U1915 (N_1915,In_592,In_299);
nor U1916 (N_1916,In_84,In_716);
nor U1917 (N_1917,In_651,In_473);
and U1918 (N_1918,In_649,In_619);
nor U1919 (N_1919,In_998,In_57);
nand U1920 (N_1920,In_410,In_577);
and U1921 (N_1921,In_515,In_563);
or U1922 (N_1922,In_540,In_972);
nor U1923 (N_1923,In_196,In_264);
xor U1924 (N_1924,In_175,In_632);
or U1925 (N_1925,In_662,In_370);
nor U1926 (N_1926,In_346,In_970);
nor U1927 (N_1927,In_547,In_678);
nand U1928 (N_1928,In_122,In_666);
or U1929 (N_1929,In_297,In_244);
nor U1930 (N_1930,In_42,In_740);
nor U1931 (N_1931,In_714,In_124);
nand U1932 (N_1932,In_207,In_493);
or U1933 (N_1933,In_829,In_506);
or U1934 (N_1934,In_901,In_771);
nor U1935 (N_1935,In_208,In_501);
or U1936 (N_1936,In_847,In_533);
and U1937 (N_1937,In_157,In_678);
nor U1938 (N_1938,In_935,In_349);
and U1939 (N_1939,In_476,In_363);
nand U1940 (N_1940,In_180,In_270);
nor U1941 (N_1941,In_317,In_350);
and U1942 (N_1942,In_62,In_492);
or U1943 (N_1943,In_716,In_255);
or U1944 (N_1944,In_378,In_105);
and U1945 (N_1945,In_866,In_136);
and U1946 (N_1946,In_784,In_730);
and U1947 (N_1947,In_989,In_430);
nor U1948 (N_1948,In_716,In_959);
or U1949 (N_1949,In_604,In_680);
or U1950 (N_1950,In_914,In_451);
nor U1951 (N_1951,In_283,In_509);
and U1952 (N_1952,In_2,In_402);
nand U1953 (N_1953,In_627,In_664);
nand U1954 (N_1954,In_491,In_735);
or U1955 (N_1955,In_146,In_748);
nand U1956 (N_1956,In_960,In_991);
nor U1957 (N_1957,In_100,In_4);
and U1958 (N_1958,In_855,In_983);
and U1959 (N_1959,In_820,In_573);
nand U1960 (N_1960,In_171,In_981);
nand U1961 (N_1961,In_898,In_321);
and U1962 (N_1962,In_998,In_82);
and U1963 (N_1963,In_55,In_759);
and U1964 (N_1964,In_77,In_434);
nand U1965 (N_1965,In_851,In_725);
nand U1966 (N_1966,In_88,In_755);
xor U1967 (N_1967,In_239,In_62);
and U1968 (N_1968,In_302,In_0);
nor U1969 (N_1969,In_818,In_706);
and U1970 (N_1970,In_611,In_432);
nand U1971 (N_1971,In_317,In_121);
nand U1972 (N_1972,In_569,In_656);
and U1973 (N_1973,In_684,In_785);
and U1974 (N_1974,In_971,In_368);
nor U1975 (N_1975,In_737,In_375);
or U1976 (N_1976,In_769,In_492);
or U1977 (N_1977,In_130,In_393);
or U1978 (N_1978,In_569,In_603);
or U1979 (N_1979,In_588,In_430);
nor U1980 (N_1980,In_591,In_186);
and U1981 (N_1981,In_407,In_958);
xnor U1982 (N_1982,In_813,In_643);
nand U1983 (N_1983,In_492,In_367);
xor U1984 (N_1984,In_259,In_287);
or U1985 (N_1985,In_680,In_391);
nor U1986 (N_1986,In_873,In_486);
or U1987 (N_1987,In_622,In_836);
and U1988 (N_1988,In_730,In_577);
and U1989 (N_1989,In_557,In_675);
nand U1990 (N_1990,In_316,In_668);
or U1991 (N_1991,In_674,In_426);
nor U1992 (N_1992,In_498,In_594);
nand U1993 (N_1993,In_245,In_314);
nand U1994 (N_1994,In_797,In_652);
nor U1995 (N_1995,In_616,In_454);
nand U1996 (N_1996,In_982,In_415);
nand U1997 (N_1997,In_89,In_975);
or U1998 (N_1998,In_385,In_266);
nand U1999 (N_1999,In_49,In_630);
nor U2000 (N_2000,N_1743,N_866);
or U2001 (N_2001,N_1993,N_1148);
and U2002 (N_2002,N_1955,N_1238);
nand U2003 (N_2003,N_1417,N_1939);
nand U2004 (N_2004,N_1801,N_4);
and U2005 (N_2005,N_1609,N_82);
and U2006 (N_2006,N_371,N_195);
or U2007 (N_2007,N_1235,N_1927);
nor U2008 (N_2008,N_149,N_309);
and U2009 (N_2009,N_1740,N_1626);
nor U2010 (N_2010,N_1206,N_406);
and U2011 (N_2011,N_842,N_36);
and U2012 (N_2012,N_1281,N_709);
nor U2013 (N_2013,N_1461,N_347);
and U2014 (N_2014,N_443,N_490);
nor U2015 (N_2015,N_224,N_227);
and U2016 (N_2016,N_1604,N_783);
nor U2017 (N_2017,N_1180,N_806);
nor U2018 (N_2018,N_365,N_179);
or U2019 (N_2019,N_1698,N_805);
nand U2020 (N_2020,N_1845,N_1284);
and U2021 (N_2021,N_37,N_1713);
nand U2022 (N_2022,N_1804,N_995);
nor U2023 (N_2023,N_1791,N_1203);
nor U2024 (N_2024,N_959,N_1314);
nand U2025 (N_2025,N_1077,N_1857);
or U2026 (N_2026,N_73,N_1156);
or U2027 (N_2027,N_379,N_780);
nor U2028 (N_2028,N_15,N_1997);
nand U2029 (N_2029,N_507,N_751);
nand U2030 (N_2030,N_1871,N_785);
nand U2031 (N_2031,N_606,N_577);
or U2032 (N_2032,N_90,N_337);
and U2033 (N_2033,N_967,N_311);
and U2034 (N_2034,N_1049,N_448);
and U2035 (N_2035,N_1310,N_703);
xor U2036 (N_2036,N_1442,N_468);
nor U2037 (N_2037,N_279,N_171);
or U2038 (N_2038,N_1233,N_1839);
or U2039 (N_2039,N_1289,N_217);
nor U2040 (N_2040,N_887,N_612);
and U2041 (N_2041,N_839,N_1759);
nor U2042 (N_2042,N_794,N_84);
nand U2043 (N_2043,N_871,N_289);
nand U2044 (N_2044,N_412,N_1229);
and U2045 (N_2045,N_450,N_1918);
and U2046 (N_2046,N_109,N_1470);
nor U2047 (N_2047,N_91,N_668);
xor U2048 (N_2048,N_1559,N_1989);
and U2049 (N_2049,N_1981,N_1856);
and U2050 (N_2050,N_1533,N_188);
nand U2051 (N_2051,N_1798,N_1455);
nand U2052 (N_2052,N_315,N_1015);
or U2053 (N_2053,N_342,N_1732);
nand U2054 (N_2054,N_1551,N_620);
nor U2055 (N_2055,N_387,N_1968);
or U2056 (N_2056,N_1560,N_1902);
nor U2057 (N_2057,N_62,N_1007);
or U2058 (N_2058,N_128,N_1087);
or U2059 (N_2059,N_1762,N_457);
nor U2060 (N_2060,N_1367,N_1772);
nand U2061 (N_2061,N_994,N_303);
and U2062 (N_2062,N_1598,N_1612);
and U2063 (N_2063,N_1773,N_334);
nand U2064 (N_2064,N_1123,N_1276);
or U2065 (N_2065,N_661,N_398);
nor U2066 (N_2066,N_576,N_1805);
nor U2067 (N_2067,N_25,N_1429);
nand U2068 (N_2068,N_1402,N_1568);
or U2069 (N_2069,N_1122,N_597);
nand U2070 (N_2070,N_1127,N_1465);
or U2071 (N_2071,N_1980,N_990);
nor U2072 (N_2072,N_755,N_1374);
nor U2073 (N_2073,N_1887,N_1843);
nor U2074 (N_2074,N_1877,N_1253);
nor U2075 (N_2075,N_79,N_1269);
or U2076 (N_2076,N_1034,N_833);
nand U2077 (N_2077,N_393,N_1022);
nand U2078 (N_2078,N_1178,N_446);
and U2079 (N_2079,N_1701,N_1216);
and U2080 (N_2080,N_556,N_300);
nand U2081 (N_2081,N_1308,N_459);
nand U2082 (N_2082,N_1225,N_1948);
nor U2083 (N_2083,N_1489,N_472);
nor U2084 (N_2084,N_123,N_1067);
nand U2085 (N_2085,N_1564,N_939);
or U2086 (N_2086,N_1386,N_1357);
nor U2087 (N_2087,N_1135,N_242);
or U2088 (N_2088,N_1230,N_759);
nor U2089 (N_2089,N_110,N_1690);
nand U2090 (N_2090,N_376,N_1545);
or U2091 (N_2091,N_918,N_72);
and U2092 (N_2092,N_138,N_438);
nand U2093 (N_2093,N_103,N_87);
nor U2094 (N_2094,N_595,N_1193);
and U2095 (N_2095,N_1614,N_1524);
or U2096 (N_2096,N_182,N_1247);
or U2097 (N_2097,N_1864,N_1058);
or U2098 (N_2098,N_470,N_161);
xor U2099 (N_2099,N_1766,N_1624);
and U2100 (N_2100,N_466,N_697);
and U2101 (N_2101,N_861,N_875);
or U2102 (N_2102,N_1358,N_813);
and U2103 (N_2103,N_1011,N_1344);
or U2104 (N_2104,N_276,N_167);
nor U2105 (N_2105,N_904,N_1466);
nand U2106 (N_2106,N_1395,N_1050);
or U2107 (N_2107,N_1115,N_1953);
nand U2108 (N_2108,N_1498,N_894);
or U2109 (N_2109,N_1616,N_1542);
nor U2110 (N_2110,N_1544,N_692);
or U2111 (N_2111,N_1280,N_1248);
and U2112 (N_2112,N_1549,N_1271);
nand U2113 (N_2113,N_1913,N_7);
xnor U2114 (N_2114,N_1320,N_1454);
nor U2115 (N_2115,N_1337,N_679);
nor U2116 (N_2116,N_847,N_1899);
nor U2117 (N_2117,N_44,N_1543);
and U2118 (N_2118,N_296,N_1033);
and U2119 (N_2119,N_1062,N_822);
and U2120 (N_2120,N_302,N_1673);
and U2121 (N_2121,N_1041,N_1069);
and U2122 (N_2122,N_1586,N_1240);
nor U2123 (N_2123,N_1605,N_1052);
and U2124 (N_2124,N_793,N_69);
and U2125 (N_2125,N_1671,N_1005);
and U2126 (N_2126,N_392,N_1014);
nor U2127 (N_2127,N_1095,N_1736);
and U2128 (N_2128,N_488,N_1644);
or U2129 (N_2129,N_530,N_405);
nor U2130 (N_2130,N_1046,N_1456);
nor U2131 (N_2131,N_1438,N_629);
nand U2132 (N_2132,N_1194,N_1029);
nand U2133 (N_2133,N_1497,N_747);
or U2134 (N_2134,N_1929,N_622);
nor U2135 (N_2135,N_1189,N_1141);
and U2136 (N_2136,N_665,N_1922);
nand U2137 (N_2137,N_16,N_433);
nor U2138 (N_2138,N_732,N_854);
nand U2139 (N_2139,N_153,N_1567);
or U2140 (N_2140,N_89,N_1200);
xnor U2141 (N_2141,N_1841,N_1728);
nand U2142 (N_2142,N_1629,N_441);
nor U2143 (N_2143,N_28,N_632);
and U2144 (N_2144,N_966,N_1341);
and U2145 (N_2145,N_796,N_808);
and U2146 (N_2146,N_343,N_1602);
nor U2147 (N_2147,N_1878,N_624);
or U2148 (N_2148,N_1219,N_583);
nand U2149 (N_2149,N_1053,N_341);
nor U2150 (N_2150,N_156,N_115);
nand U2151 (N_2151,N_1696,N_504);
and U2152 (N_2152,N_1943,N_71);
nor U2153 (N_2153,N_1622,N_493);
nand U2154 (N_2154,N_1170,N_1484);
and U2155 (N_2155,N_338,N_1304);
or U2156 (N_2156,N_559,N_225);
or U2157 (N_2157,N_201,N_1411);
nand U2158 (N_2158,N_418,N_1583);
nor U2159 (N_2159,N_1196,N_529);
nor U2160 (N_2160,N_1969,N_723);
or U2161 (N_2161,N_1302,N_718);
xor U2162 (N_2162,N_1630,N_1517);
nor U2163 (N_2163,N_545,N_1645);
nor U2164 (N_2164,N_1316,N_618);
nor U2165 (N_2165,N_1361,N_1575);
and U2166 (N_2166,N_155,N_810);
or U2167 (N_2167,N_1255,N_193);
nor U2168 (N_2168,N_215,N_971);
and U2169 (N_2169,N_667,N_1990);
nor U2170 (N_2170,N_125,N_1243);
and U2171 (N_2171,N_672,N_210);
or U2172 (N_2172,N_1160,N_141);
or U2173 (N_2173,N_1432,N_1802);
nor U2174 (N_2174,N_1717,N_584);
nand U2175 (N_2175,N_1515,N_1824);
nor U2176 (N_2176,N_340,N_586);
nor U2177 (N_2177,N_1708,N_38);
and U2178 (N_2178,N_1163,N_1472);
nor U2179 (N_2179,N_795,N_1075);
or U2180 (N_2180,N_1526,N_758);
or U2181 (N_2181,N_1844,N_851);
and U2182 (N_2182,N_1486,N_1);
and U2183 (N_2183,N_106,N_476);
nand U2184 (N_2184,N_1827,N_250);
xnor U2185 (N_2185,N_230,N_693);
and U2186 (N_2186,N_1114,N_497);
nor U2187 (N_2187,N_708,N_88);
nand U2188 (N_2188,N_688,N_626);
nor U2189 (N_2189,N_1781,N_605);
or U2190 (N_2190,N_190,N_982);
nand U2191 (N_2191,N_1719,N_915);
nand U2192 (N_2192,N_1474,N_1352);
and U2193 (N_2193,N_1680,N_993);
nor U2194 (N_2194,N_734,N_878);
nor U2195 (N_2195,N_1169,N_1735);
or U2196 (N_2196,N_1172,N_820);
or U2197 (N_2197,N_1836,N_409);
nand U2198 (N_2198,N_1443,N_389);
nor U2199 (N_2199,N_328,N_998);
or U2200 (N_2200,N_1511,N_1829);
nor U2201 (N_2201,N_1168,N_1419);
nand U2202 (N_2202,N_1152,N_237);
or U2203 (N_2203,N_1082,N_211);
nor U2204 (N_2204,N_360,N_677);
nand U2205 (N_2205,N_701,N_1978);
and U2206 (N_2206,N_1848,N_295);
nand U2207 (N_2207,N_940,N_1900);
and U2208 (N_2208,N_938,N_1600);
and U2209 (N_2209,N_1938,N_1648);
nor U2210 (N_2210,N_401,N_953);
or U2211 (N_2211,N_1108,N_837);
nand U2212 (N_2212,N_1322,N_272);
and U2213 (N_2213,N_1699,N_5);
nand U2214 (N_2214,N_1942,N_1146);
and U2215 (N_2215,N_1550,N_163);
nor U2216 (N_2216,N_565,N_1928);
nand U2217 (N_2217,N_160,N_1555);
nor U2218 (N_2218,N_453,N_56);
or U2219 (N_2219,N_893,N_1822);
nand U2220 (N_2220,N_1558,N_891);
or U2221 (N_2221,N_1202,N_1868);
or U2222 (N_2222,N_1319,N_1399);
nor U2223 (N_2223,N_977,N_1599);
or U2224 (N_2224,N_1998,N_1339);
nand U2225 (N_2225,N_1334,N_1991);
or U2226 (N_2226,N_521,N_293);
and U2227 (N_2227,N_102,N_526);
and U2228 (N_2228,N_1979,N_1274);
nor U2229 (N_2229,N_1278,N_1950);
nor U2230 (N_2230,N_1256,N_479);
or U2231 (N_2231,N_1045,N_706);
xnor U2232 (N_2232,N_1579,N_1338);
or U2233 (N_2233,N_1394,N_18);
and U2234 (N_2234,N_1907,N_856);
or U2235 (N_2235,N_763,N_542);
or U2236 (N_2236,N_1724,N_1966);
and U2237 (N_2237,N_1407,N_435);
and U2238 (N_2238,N_1227,N_1353);
nor U2239 (N_2239,N_1557,N_55);
nand U2240 (N_2240,N_419,N_651);
or U2241 (N_2241,N_1705,N_1273);
or U2242 (N_2242,N_1679,N_1783);
and U2243 (N_2243,N_455,N_1342);
or U2244 (N_2244,N_6,N_1422);
nand U2245 (N_2245,N_275,N_650);
and U2246 (N_2246,N_1300,N_996);
nand U2247 (N_2247,N_738,N_528);
nor U2248 (N_2248,N_34,N_273);
nor U2249 (N_2249,N_1885,N_1576);
and U2250 (N_2250,N_588,N_1686);
or U2251 (N_2251,N_1984,N_580);
or U2252 (N_2252,N_463,N_614);
nand U2253 (N_2253,N_1056,N_817);
nand U2254 (N_2254,N_277,N_807);
or U2255 (N_2255,N_1987,N_1157);
nor U2256 (N_2256,N_1179,N_1329);
and U2257 (N_2257,N_284,N_1912);
and U2258 (N_2258,N_546,N_963);
or U2259 (N_2259,N_579,N_257);
and U2260 (N_2260,N_176,N_930);
nor U2261 (N_2261,N_669,N_1716);
and U2262 (N_2262,N_321,N_1584);
and U2263 (N_2263,N_1167,N_1875);
and U2264 (N_2264,N_1734,N_178);
xor U2265 (N_2265,N_634,N_1574);
nor U2266 (N_2266,N_999,N_183);
nor U2267 (N_2267,N_1646,N_1129);
nor U2268 (N_2268,N_1946,N_846);
xnor U2269 (N_2269,N_370,N_946);
nor U2270 (N_2270,N_1267,N_1910);
nor U2271 (N_2271,N_1427,N_1682);
nand U2272 (N_2272,N_1529,N_481);
nand U2273 (N_2273,N_675,N_1016);
nand U2274 (N_2274,N_881,N_1116);
nor U2275 (N_2275,N_263,N_1873);
nor U2276 (N_2276,N_567,N_451);
or U2277 (N_2277,N_663,N_1239);
or U2278 (N_2278,N_883,N_494);
and U2279 (N_2279,N_1400,N_327);
or U2280 (N_2280,N_400,N_863);
and U2281 (N_2281,N_762,N_424);
and U2282 (N_2282,N_462,N_749);
and U2283 (N_2283,N_1591,N_1720);
or U2284 (N_2284,N_1711,N_269);
and U2285 (N_2285,N_322,N_1659);
or U2286 (N_2286,N_613,N_59);
nor U2287 (N_2287,N_53,N_460);
or U2288 (N_2288,N_169,N_245);
nor U2289 (N_2289,N_205,N_1217);
nor U2290 (N_2290,N_1897,N_148);
and U2291 (N_2291,N_757,N_864);
and U2292 (N_2292,N_484,N_702);
and U2293 (N_2293,N_301,N_524);
nand U2294 (N_2294,N_1042,N_1688);
and U2295 (N_2295,N_168,N_635);
nand U2296 (N_2296,N_1261,N_126);
or U2297 (N_2297,N_1272,N_1293);
nor U2298 (N_2298,N_827,N_386);
or U2299 (N_2299,N_974,N_222);
nor U2300 (N_2300,N_1351,N_1265);
and U2301 (N_2301,N_391,N_94);
and U2302 (N_2302,N_666,N_1488);
or U2303 (N_2303,N_1401,N_1870);
or U2304 (N_2304,N_1136,N_1995);
and U2305 (N_2305,N_477,N_495);
nand U2306 (N_2306,N_243,N_20);
and U2307 (N_2307,N_1816,N_234);
nand U2308 (N_2308,N_1371,N_748);
nand U2309 (N_2309,N_778,N_388);
nand U2310 (N_2310,N_1949,N_882);
and U2311 (N_2311,N_1769,N_1643);
and U2312 (N_2312,N_1933,N_951);
and U2313 (N_2313,N_1161,N_304);
and U2314 (N_2314,N_905,N_766);
nand U2315 (N_2315,N_1974,N_417);
and U2316 (N_2316,N_1828,N_1865);
and U2317 (N_2317,N_403,N_1467);
or U2318 (N_2318,N_1012,N_1428);
nand U2319 (N_2319,N_1635,N_1986);
nor U2320 (N_2320,N_1785,N_870);
and U2321 (N_2321,N_1538,N_544);
nand U2322 (N_2322,N_1722,N_1296);
and U2323 (N_2323,N_1318,N_1074);
or U2324 (N_2324,N_465,N_578);
and U2325 (N_2325,N_180,N_1208);
nor U2326 (N_2326,N_478,N_1668);
nand U2327 (N_2327,N_1889,N_1071);
xor U2328 (N_2328,N_1301,N_1391);
nor U2329 (N_2329,N_1960,N_727);
nand U2330 (N_2330,N_1295,N_1177);
xnor U2331 (N_2331,N_114,N_1651);
nor U2332 (N_2332,N_120,N_592);
and U2333 (N_2333,N_884,N_1655);
nor U2334 (N_2334,N_1424,N_1633);
and U2335 (N_2335,N_714,N_1493);
nand U2336 (N_2336,N_814,N_744);
nand U2337 (N_2337,N_1096,N_1081);
or U2338 (N_2338,N_609,N_278);
nand U2339 (N_2339,N_1796,N_533);
nand U2340 (N_2340,N_306,N_1752);
nor U2341 (N_2341,N_1185,N_1530);
nor U2342 (N_2342,N_538,N_8);
or U2343 (N_2343,N_1657,N_710);
nand U2344 (N_2344,N_1259,N_1628);
and U2345 (N_2345,N_662,N_1468);
or U2346 (N_2346,N_218,N_850);
and U2347 (N_2347,N_261,N_1749);
and U2348 (N_2348,N_1704,N_1669);
and U2349 (N_2349,N_1482,N_1617);
and U2350 (N_2350,N_925,N_1692);
nor U2351 (N_2351,N_313,N_1967);
or U2352 (N_2352,N_1649,N_829);
nand U2353 (N_2353,N_64,N_202);
nor U2354 (N_2354,N_911,N_1171);
or U2355 (N_2355,N_654,N_442);
and U2356 (N_2356,N_1092,N_1840);
nand U2357 (N_2357,N_1057,N_1154);
and U2358 (N_2358,N_921,N_444);
or U2359 (N_2359,N_185,N_1744);
xnor U2360 (N_2360,N_1436,N_906);
nand U2361 (N_2361,N_562,N_139);
xnor U2362 (N_2362,N_1770,N_962);
nor U2363 (N_2363,N_857,N_1106);
nand U2364 (N_2364,N_1001,N_1742);
nand U2365 (N_2365,N_181,N_75);
nor U2366 (N_2366,N_888,N_1354);
and U2367 (N_2367,N_671,N_1257);
nand U2368 (N_2368,N_1309,N_1676);
nand U2369 (N_2369,N_124,N_536);
nor U2370 (N_2370,N_1416,N_791);
xor U2371 (N_2371,N_1457,N_652);
and U2372 (N_2372,N_281,N_825);
or U2373 (N_2373,N_320,N_1712);
and U2374 (N_2374,N_235,N_118);
nor U2375 (N_2375,N_1126,N_1390);
and U2376 (N_2376,N_1697,N_283);
nand U2377 (N_2377,N_367,N_1027);
nor U2378 (N_2378,N_1317,N_98);
or U2379 (N_2379,N_876,N_601);
or U2380 (N_2380,N_502,N_1187);
nor U2381 (N_2381,N_1565,N_687);
or U2382 (N_2382,N_1502,N_240);
and U2383 (N_2383,N_1547,N_9);
and U2384 (N_2384,N_375,N_1691);
nor U2385 (N_2385,N_1729,N_1348);
and U2386 (N_2386,N_700,N_792);
nor U2387 (N_2387,N_1774,N_655);
nand U2388 (N_2388,N_1408,N_816);
or U2389 (N_2389,N_1174,N_1483);
or U2390 (N_2390,N_1364,N_1250);
or U2391 (N_2391,N_1144,N_1509);
and U2392 (N_2392,N_1236,N_19);
nand U2393 (N_2393,N_838,N_162);
nand U2394 (N_2394,N_177,N_362);
nand U2395 (N_2395,N_383,N_1055);
nand U2396 (N_2396,N_191,N_1621);
nor U2397 (N_2397,N_127,N_1919);
or U2398 (N_2398,N_889,N_725);
and U2399 (N_2399,N_1283,N_831);
or U2400 (N_2400,N_599,N_901);
and U2401 (N_2401,N_143,N_1365);
nand U2402 (N_2402,N_1937,N_1715);
nor U2403 (N_2403,N_518,N_726);
and U2404 (N_2404,N_947,N_1009);
and U2405 (N_2405,N_512,N_39);
or U2406 (N_2406,N_1125,N_2);
and U2407 (N_2407,N_1748,N_1477);
and U2408 (N_2408,N_522,N_927);
or U2409 (N_2409,N_426,N_1406);
and U2410 (N_2410,N_552,N_1776);
or U2411 (N_2411,N_1932,N_1287);
or U2412 (N_2412,N_1113,N_1833);
and U2413 (N_2413,N_1858,N_855);
or U2414 (N_2414,N_1037,N_449);
and U2415 (N_2415,N_743,N_1355);
and U2416 (N_2416,N_1039,N_1448);
and U2417 (N_2417,N_253,N_975);
xor U2418 (N_2418,N_683,N_1531);
nor U2419 (N_2419,N_1940,N_213);
or U2420 (N_2420,N_61,N_1331);
and U2421 (N_2421,N_48,N_698);
nand U2422 (N_2422,N_1909,N_571);
or U2423 (N_2423,N_1755,N_1571);
and U2424 (N_2424,N_1879,N_1464);
and U2425 (N_2425,N_603,N_1388);
xor U2426 (N_2426,N_1514,N_122);
and U2427 (N_2427,N_1479,N_540);
or U2428 (N_2428,N_228,N_1445);
or U2429 (N_2429,N_413,N_1996);
or U2430 (N_2430,N_1925,N_1539);
or U2431 (N_2431,N_1028,N_1186);
and U2432 (N_2432,N_731,N_1820);
nor U2433 (N_2433,N_745,N_395);
or U2434 (N_2434,N_437,N_1880);
and U2435 (N_2435,N_1393,N_1917);
nand U2436 (N_2436,N_991,N_531);
nor U2437 (N_2437,N_789,N_1220);
and U2438 (N_2438,N_802,N_722);
nor U2439 (N_2439,N_226,N_1963);
xnor U2440 (N_2440,N_1204,N_616);
and U2441 (N_2441,N_1312,N_1094);
or U2442 (N_2442,N_1473,N_1527);
or U2443 (N_2443,N_117,N_937);
or U2444 (N_2444,N_374,N_1916);
or U2445 (N_2445,N_1205,N_1849);
and U2446 (N_2446,N_354,N_1176);
and U2447 (N_2447,N_1131,N_1876);
or U2448 (N_2448,N_608,N_1241);
or U2449 (N_2449,N_135,N_1377);
xor U2450 (N_2450,N_355,N_916);
and U2451 (N_2451,N_421,N_93);
nor U2452 (N_2452,N_1100,N_694);
nor U2453 (N_2453,N_335,N_648);
and U2454 (N_2454,N_1852,N_1546);
nor U2455 (N_2455,N_330,N_933);
nor U2456 (N_2456,N_316,N_1786);
nor U2457 (N_2457,N_1258,N_619);
nor U2458 (N_2458,N_569,N_547);
or U2459 (N_2459,N_339,N_1961);
and U2460 (N_2460,N_1634,N_454);
and U2461 (N_2461,N_1260,N_644);
and U2462 (N_2462,N_945,N_843);
and U2463 (N_2463,N_1693,N_903);
and U2464 (N_2464,N_1494,N_769);
nand U2465 (N_2465,N_845,N_1359);
and U2466 (N_2466,N_853,N_1590);
nand U2467 (N_2467,N_452,N_1866);
nand U2468 (N_2468,N_1199,N_189);
and U2469 (N_2469,N_509,N_1703);
nand U2470 (N_2470,N_910,N_95);
and U2471 (N_2471,N_1104,N_832);
or U2472 (N_2472,N_862,N_57);
nand U2473 (N_2473,N_359,N_63);
or U2474 (N_2474,N_1660,N_1751);
nand U2475 (N_2475,N_49,N_645);
and U2476 (N_2476,N_1155,N_1487);
or U2477 (N_2477,N_1895,N_1418);
nor U2478 (N_2478,N_1362,N_611);
nand U2479 (N_2479,N_27,N_146);
and U2480 (N_2480,N_1971,N_1982);
nand U2481 (N_2481,N_1387,N_1678);
and U2482 (N_2482,N_1327,N_1097);
nor U2483 (N_2483,N_1972,N_1663);
nor U2484 (N_2484,N_0,N_1279);
or U2485 (N_2485,N_271,N_416);
and U2486 (N_2486,N_1638,N_372);
nor U2487 (N_2487,N_458,N_978);
nor U2488 (N_2488,N_828,N_407);
or U2489 (N_2489,N_1935,N_1745);
or U2490 (N_2490,N_1110,N_1190);
or U2491 (N_2491,N_384,N_377);
and U2492 (N_2492,N_1882,N_1434);
nor U2493 (N_2493,N_1573,N_184);
or U2494 (N_2494,N_1587,N_1893);
nand U2495 (N_2495,N_630,N_811);
nand U2496 (N_2496,N_23,N_1288);
nand U2497 (N_2497,N_1166,N_1409);
nand U2498 (N_2498,N_724,N_174);
or U2499 (N_2499,N_404,N_1924);
or U2500 (N_2500,N_657,N_1784);
and U2501 (N_2501,N_1505,N_1750);
nand U2502 (N_2502,N_1681,N_775);
nand U2503 (N_2503,N_1631,N_638);
nand U2504 (N_2504,N_1814,N_505);
nand U2505 (N_2505,N_1218,N_1811);
and U2506 (N_2506,N_1025,N_1051);
xnor U2507 (N_2507,N_1452,N_1192);
nand U2508 (N_2508,N_1132,N_886);
or U2509 (N_2509,N_267,N_525);
nor U2510 (N_2510,N_517,N_1021);
or U2511 (N_2511,N_1210,N_1119);
or U2512 (N_2512,N_501,N_1290);
or U2513 (N_2513,N_65,N_285);
and U2514 (N_2514,N_575,N_765);
and U2515 (N_2515,N_1731,N_1201);
or U2516 (N_2516,N_41,N_1469);
and U2517 (N_2517,N_594,N_1263);
nand U2518 (N_2518,N_1000,N_969);
or U2519 (N_2519,N_840,N_643);
and U2520 (N_2520,N_952,N_1164);
or U2521 (N_2521,N_1026,N_1817);
nand U2522 (N_2522,N_1398,N_844);
xnor U2523 (N_2523,N_76,N_1262);
and U2524 (N_2524,N_976,N_1884);
nor U2525 (N_2525,N_1444,N_1091);
and U2526 (N_2526,N_1725,N_1458);
and U2527 (N_2527,N_1777,N_768);
or U2528 (N_2528,N_1085,N_1003);
and U2529 (N_2529,N_582,N_907);
nand U2530 (N_2530,N_1675,N_394);
or U2531 (N_2531,N_1345,N_349);
and U2532 (N_2532,N_430,N_1992);
and U2533 (N_2533,N_1637,N_673);
nand U2534 (N_2534,N_1117,N_67);
and U2535 (N_2535,N_1874,N_1107);
nand U2536 (N_2536,N_137,N_1439);
and U2537 (N_2537,N_209,N_11);
nand U2538 (N_2538,N_1449,N_1385);
and U2539 (N_2539,N_314,N_591);
nor U2540 (N_2540,N_1898,N_572);
or U2541 (N_2541,N_231,N_1032);
nor U2542 (N_2542,N_782,N_1410);
and U2543 (N_2543,N_539,N_24);
nand U2544 (N_2544,N_1632,N_1471);
nand U2545 (N_2545,N_1554,N_848);
nand U2546 (N_2546,N_1883,N_134);
or U2547 (N_2547,N_1294,N_500);
nor U2548 (N_2548,N_1459,N_1491);
and U2549 (N_2549,N_1595,N_1739);
nand U2550 (N_2550,N_1596,N_1862);
nand U2551 (N_2551,N_923,N_682);
or U2552 (N_2552,N_1023,N_1321);
or U2553 (N_2553,N_1608,N_239);
or U2554 (N_2554,N_898,N_1232);
and U2555 (N_2555,N_1797,N_1881);
and U2556 (N_2556,N_173,N_908);
or U2557 (N_2557,N_1249,N_553);
nor U2558 (N_2558,N_986,N_487);
and U2559 (N_2559,N_108,N_1589);
and U2560 (N_2560,N_873,N_1767);
nand U2561 (N_2561,N_194,N_116);
nor U2562 (N_2562,N_1142,N_212);
nor U2563 (N_2563,N_1794,N_1658);
nand U2564 (N_2564,N_865,N_81);
or U2565 (N_2565,N_1112,N_1872);
nand U2566 (N_2566,N_1672,N_784);
xor U2567 (N_2567,N_1140,N_610);
xnor U2568 (N_2568,N_1209,N_600);
and U2569 (N_2569,N_1674,N_1368);
nor U2570 (N_2570,N_1832,N_1702);
nor U2571 (N_2571,N_80,N_260);
and U2572 (N_2572,N_968,N_1420);
nand U2573 (N_2573,N_1476,N_877);
and U2574 (N_2574,N_1809,N_589);
or U2575 (N_2575,N_111,N_1561);
or U2576 (N_2576,N_914,N_1346);
nand U2577 (N_2577,N_199,N_1747);
nand U2578 (N_2578,N_97,N_1709);
nor U2579 (N_2579,N_1004,N_642);
nor U2580 (N_2580,N_1510,N_1453);
nor U2581 (N_2581,N_1830,N_506);
nor U2582 (N_2582,N_1437,N_639);
nand U2583 (N_2583,N_988,N_1431);
or U2584 (N_2584,N_874,N_568);
and U2585 (N_2585,N_381,N_1286);
and U2586 (N_2586,N_1006,N_13);
or U2587 (N_2587,N_1277,N_779);
nor U2588 (N_2588,N_1381,N_1184);
or U2589 (N_2589,N_1532,N_107);
or U2590 (N_2590,N_890,N_1723);
nand U2591 (N_2591,N_436,N_944);
and U2592 (N_2592,N_198,N_70);
nand U2593 (N_2593,N_985,N_729);
nor U2594 (N_2594,N_1291,N_1807);
nor U2595 (N_2595,N_196,N_1315);
or U2596 (N_2596,N_1519,N_598);
nor U2597 (N_2597,N_1297,N_1450);
or U2598 (N_2598,N_40,N_1661);
and U2599 (N_2599,N_428,N_913);
or U2600 (N_2600,N_411,N_1552);
nor U2601 (N_2601,N_1423,N_204);
nand U2602 (N_2602,N_532,N_1562);
nand U2603 (N_2603,N_1372,N_989);
xor U2604 (N_2604,N_77,N_399);
nor U2605 (N_2605,N_319,N_51);
xnor U2606 (N_2606,N_1079,N_772);
or U2607 (N_2607,N_1954,N_647);
nand U2608 (N_2608,N_761,N_1415);
nand U2609 (N_2609,N_236,N_26);
or U2610 (N_2610,N_818,N_1855);
nor U2611 (N_2611,N_909,N_1780);
or U2612 (N_2612,N_1480,N_307);
and U2613 (N_2613,N_207,N_1516);
or U2614 (N_2614,N_1414,N_535);
and U2615 (N_2615,N_860,N_1109);
and U2616 (N_2616,N_86,N_471);
nor U2617 (N_2617,N_1306,N_1463);
xor U2618 (N_2618,N_1447,N_473);
nand U2619 (N_2619,N_1754,N_1335);
nand U2620 (N_2620,N_965,N_1815);
nor U2621 (N_2621,N_364,N_1008);
and U2622 (N_2622,N_1268,N_158);
or U2623 (N_2623,N_1044,N_821);
or U2624 (N_2624,N_824,N_1541);
and U2625 (N_2625,N_1741,N_1641);
and U2626 (N_2626,N_1799,N_972);
or U2627 (N_2627,N_1093,N_297);
nor U2628 (N_2628,N_1689,N_920);
or U2629 (N_2629,N_46,N_17);
nor U2630 (N_2630,N_1506,N_423);
xor U2631 (N_2631,N_1298,N_1650);
or U2632 (N_2632,N_1061,N_564);
and U2633 (N_2633,N_144,N_247);
or U2634 (N_2634,N_197,N_1513);
nand U2635 (N_2635,N_1603,N_1083);
and U2636 (N_2636,N_711,N_1496);
or U2637 (N_2637,N_1501,N_1894);
and U2638 (N_2638,N_1588,N_1834);
nand U2639 (N_2639,N_1404,N_1695);
nor U2640 (N_2640,N_1890,N_646);
or U2641 (N_2641,N_1066,N_456);
and U2642 (N_2642,N_561,N_1507);
and U2643 (N_2643,N_1610,N_684);
or U2644 (N_2644,N_1242,N_308);
nor U2645 (N_2645,N_514,N_604);
or U2646 (N_2646,N_941,N_804);
nor U2647 (N_2647,N_262,N_1389);
or U2648 (N_2648,N_1305,N_1592);
or U2649 (N_2649,N_1010,N_705);
and U2650 (N_2650,N_1072,N_819);
xor U2651 (N_2651,N_1782,N_1700);
and U2652 (N_2652,N_216,N_803);
nand U2653 (N_2653,N_1973,N_1647);
or U2654 (N_2654,N_58,N_1373);
nand U2655 (N_2655,N_1653,N_1964);
and U2656 (N_2656,N_291,N_1903);
and U2657 (N_2657,N_1627,N_1165);
xor U2658 (N_2658,N_1183,N_299);
nand U2659 (N_2659,N_510,N_131);
and U2660 (N_2660,N_1518,N_997);
nand U2661 (N_2661,N_1182,N_492);
or U2662 (N_2662,N_934,N_721);
and U2663 (N_2663,N_1764,N_1383);
nand U2664 (N_2664,N_754,N_1837);
and U2665 (N_2665,N_1756,N_823);
nor U2666 (N_2666,N_47,N_1325);
nand U2667 (N_2667,N_3,N_690);
nand U2668 (N_2668,N_1825,N_499);
nand U2669 (N_2669,N_1906,N_1787);
nor U2670 (N_2670,N_223,N_736);
and U2671 (N_2671,N_1888,N_469);
or U2672 (N_2672,N_429,N_1490);
xnor U2673 (N_2673,N_1369,N_1002);
nor U2674 (N_2674,N_1613,N_1252);
nand U2675 (N_2675,N_573,N_1694);
nand U2676 (N_2676,N_658,N_1636);
nand U2677 (N_2677,N_689,N_1570);
nand U2678 (N_2678,N_1036,N_660);
or U2679 (N_2679,N_1585,N_1435);
and U2680 (N_2680,N_631,N_1492);
nor U2681 (N_2681,N_1396,N_1721);
and U2682 (N_2682,N_113,N_1640);
nor U2683 (N_2683,N_1330,N_558);
and U2684 (N_2684,N_1556,N_1500);
nand U2685 (N_2685,N_602,N_14);
or U2686 (N_2686,N_1664,N_1965);
nor U2687 (N_2687,N_1800,N_1956);
and U2688 (N_2688,N_1475,N_563);
nand U2689 (N_2689,N_713,N_1215);
or U2690 (N_2690,N_1677,N_1111);
nor U2691 (N_2691,N_841,N_331);
and U2692 (N_2692,N_159,N_756);
nand U2693 (N_2693,N_1040,N_1958);
and U2694 (N_2694,N_286,N_96);
and U2695 (N_2695,N_251,N_809);
or U2696 (N_2696,N_10,N_317);
and U2697 (N_2697,N_1324,N_1826);
nor U2698 (N_2698,N_1124,N_636);
or U2699 (N_2699,N_422,N_943);
and U2700 (N_2700,N_764,N_1508);
or U2701 (N_2701,N_1606,N_1896);
nand U2702 (N_2702,N_397,N_129);
and U2703 (N_2703,N_1535,N_935);
nand U2704 (N_2704,N_1860,N_753);
or U2705 (N_2705,N_1838,N_554);
nand U2706 (N_2706,N_593,N_1652);
and U2707 (N_2707,N_485,N_1941);
nand U2708 (N_2708,N_1191,N_1099);
nor U2709 (N_2709,N_1080,N_742);
or U2710 (N_2710,N_1303,N_318);
xnor U2711 (N_2711,N_1019,N_1195);
or U2712 (N_2712,N_1266,N_192);
xor U2713 (N_2713,N_681,N_1118);
nor U2714 (N_2714,N_1718,N_895);
nand U2715 (N_2715,N_1460,N_1485);
and U2716 (N_2716,N_1264,N_154);
nand U2717 (N_2717,N_979,N_1911);
and U2718 (N_2718,N_1380,N_1376);
or U2719 (N_2719,N_704,N_987);
or U2720 (N_2720,N_885,N_1581);
nand U2721 (N_2721,N_834,N_922);
and U2722 (N_2722,N_801,N_1043);
nor U2723 (N_2723,N_740,N_1285);
and U2724 (N_2724,N_352,N_1806);
and U2725 (N_2725,N_1378,N_425);
or U2726 (N_2726,N_348,N_800);
and U2727 (N_2727,N_1433,N_1921);
and U2728 (N_2728,N_170,N_746);
or U2729 (N_2729,N_798,N_1133);
and U2730 (N_2730,N_942,N_1020);
and U2731 (N_2731,N_385,N_1730);
nor U2732 (N_2732,N_696,N_1597);
or U2733 (N_2733,N_992,N_924);
nor U2734 (N_2734,N_912,N_1771);
nor U2735 (N_2735,N_100,N_1384);
and U2736 (N_2736,N_265,N_1038);
and U2737 (N_2737,N_771,N_368);
or U2738 (N_2738,N_637,N_1854);
and U2739 (N_2739,N_259,N_541);
and U2740 (N_2740,N_66,N_22);
nor U2741 (N_2741,N_1753,N_140);
nand U2742 (N_2742,N_1625,N_166);
and U2743 (N_2743,N_699,N_799);
or U2744 (N_2744,N_1211,N_1425);
nor U2745 (N_2745,N_12,N_1687);
nand U2746 (N_2746,N_1810,N_35);
nor U2747 (N_2747,N_1328,N_1379);
or U2748 (N_2748,N_1370,N_1098);
or U2749 (N_2749,N_513,N_919);
nor U2750 (N_2750,N_1665,N_1540);
xnor U2751 (N_2751,N_345,N_1145);
or U2752 (N_2752,N_382,N_574);
nor U2753 (N_2753,N_1254,N_1582);
and U2754 (N_2754,N_1332,N_1985);
nand U2755 (N_2755,N_515,N_254);
nand U2756 (N_2756,N_1959,N_1947);
or U2757 (N_2757,N_1580,N_1915);
and U2758 (N_2758,N_587,N_1363);
nand U2759 (N_2759,N_1528,N_1563);
and U2760 (N_2760,N_555,N_233);
nor U2761 (N_2761,N_33,N_21);
and U2762 (N_2762,N_511,N_615);
nor U2763 (N_2763,N_165,N_1988);
and U2764 (N_2764,N_1143,N_486);
or U2765 (N_2765,N_1392,N_835);
nor U2766 (N_2766,N_773,N_1537);
and U2767 (N_2767,N_1931,N_52);
or U2768 (N_2768,N_1024,N_695);
nand U2769 (N_2769,N_852,N_483);
nand U2770 (N_2770,N_1495,N_1951);
nand U2771 (N_2771,N_121,N_232);
or U2772 (N_2772,N_266,N_739);
and U2773 (N_2773,N_720,N_1930);
nand U2774 (N_2774,N_244,N_973);
nand U2775 (N_2775,N_1013,N_305);
xnor U2776 (N_2776,N_132,N_674);
nor U2777 (N_2777,N_1246,N_607);
and U2778 (N_2778,N_1763,N_447);
nor U2779 (N_2779,N_1221,N_187);
nand U2780 (N_2780,N_560,N_1105);
and U2781 (N_2781,N_78,N_797);
or U2782 (N_2782,N_957,N_1823);
nor U2783 (N_2783,N_1977,N_1137);
xor U2784 (N_2784,N_929,N_1863);
or U2785 (N_2785,N_1440,N_712);
and U2786 (N_2786,N_1207,N_350);
and U2787 (N_2787,N_1710,N_1760);
and U2788 (N_2788,N_1212,N_776);
or U2789 (N_2789,N_1088,N_43);
nor U2790 (N_2790,N_252,N_1162);
xor U2791 (N_2791,N_105,N_691);
or U2792 (N_2792,N_50,N_1430);
and U2793 (N_2793,N_1134,N_229);
nor U2794 (N_2794,N_1901,N_981);
nand U2795 (N_2795,N_1121,N_241);
or U2796 (N_2796,N_294,N_104);
xnor U2797 (N_2797,N_440,N_1523);
and U2798 (N_2798,N_1999,N_1223);
nand U2799 (N_2799,N_1601,N_408);
or U2800 (N_2800,N_1150,N_1788);
nand U2801 (N_2801,N_92,N_206);
nor U2802 (N_2802,N_461,N_498);
nand U2803 (N_2803,N_1578,N_445);
and U2804 (N_2804,N_1792,N_788);
nor U2805 (N_2805,N_737,N_678);
and U2806 (N_2806,N_1224,N_357);
nor U2807 (N_2807,N_145,N_1188);
nor U2808 (N_2808,N_410,N_958);
nand U2809 (N_2809,N_786,N_1994);
xor U2810 (N_2810,N_1017,N_1812);
or U2811 (N_2811,N_1451,N_516);
and U2812 (N_2812,N_1299,N_1795);
or U2813 (N_2813,N_1738,N_1356);
and U2814 (N_2814,N_949,N_312);
or U2815 (N_2815,N_750,N_101);
or U2816 (N_2816,N_336,N_1793);
and U2817 (N_2817,N_1031,N_1765);
and U2818 (N_2818,N_1397,N_68);
or U2819 (N_2819,N_1405,N_287);
and U2820 (N_2820,N_1642,N_1685);
and U2821 (N_2821,N_1270,N_1102);
or U2822 (N_2822,N_1727,N_1343);
nor U2823 (N_2823,N_475,N_363);
nor U2824 (N_2824,N_147,N_649);
nor U2825 (N_2825,N_1733,N_1173);
or U2826 (N_2826,N_332,N_220);
nor U2827 (N_2827,N_152,N_1821);
nor U2828 (N_2828,N_1761,N_523);
nor U2829 (N_2829,N_1934,N_1446);
or U2830 (N_2830,N_1983,N_1779);
or U2831 (N_2831,N_491,N_954);
nand U2832 (N_2832,N_1048,N_1462);
and U2833 (N_2833,N_717,N_760);
nand U2834 (N_2834,N_527,N_60);
nand U2835 (N_2835,N_770,N_427);
or U2836 (N_2836,N_1070,N_136);
nor U2837 (N_2837,N_325,N_480);
and U2838 (N_2838,N_329,N_557);
xor U2839 (N_2839,N_1670,N_1349);
nor U2840 (N_2840,N_520,N_200);
and U2841 (N_2841,N_292,N_256);
and U2842 (N_2842,N_581,N_1926);
nor U2843 (N_2843,N_1861,N_280);
and U2844 (N_2844,N_879,N_1054);
or U2845 (N_2845,N_1326,N_932);
nand U2846 (N_2846,N_1175,N_1128);
or U2847 (N_2847,N_1962,N_1819);
or U2848 (N_2848,N_1313,N_1835);
nor U2849 (N_2849,N_1153,N_621);
nor U2850 (N_2850,N_1251,N_1292);
xnor U2851 (N_2851,N_248,N_1244);
nand U2852 (N_2852,N_777,N_1521);
or U2853 (N_2853,N_970,N_1886);
and U2854 (N_2854,N_790,N_1914);
nand U2855 (N_2855,N_1891,N_1375);
and U2856 (N_2856,N_268,N_1867);
or U2857 (N_2857,N_625,N_390);
xor U2858 (N_2858,N_151,N_767);
or U2859 (N_2859,N_112,N_208);
and U2860 (N_2860,N_1403,N_551);
nor U2861 (N_2861,N_1512,N_290);
or U2862 (N_2862,N_1726,N_1620);
or U2863 (N_2863,N_716,N_508);
and U2864 (N_2864,N_414,N_1904);
nand U2865 (N_2865,N_172,N_1534);
and U2866 (N_2866,N_826,N_464);
nand U2867 (N_2867,N_1522,N_896);
nor U2868 (N_2868,N_1594,N_1593);
nor U2869 (N_2869,N_282,N_150);
nand U2870 (N_2870,N_752,N_264);
nand U2871 (N_2871,N_1758,N_917);
nand U2872 (N_2872,N_219,N_214);
and U2873 (N_2873,N_1619,N_1707);
nand U2874 (N_2874,N_1222,N_1656);
or U2875 (N_2875,N_142,N_715);
or U2876 (N_2876,N_869,N_1073);
nor U2877 (N_2877,N_1149,N_956);
or U2878 (N_2878,N_326,N_1101);
and U2879 (N_2879,N_203,N_1499);
or U2880 (N_2880,N_1197,N_830);
or U2881 (N_2881,N_1350,N_570);
nand U2882 (N_2882,N_373,N_489);
xnor U2883 (N_2883,N_984,N_1018);
and U2884 (N_2884,N_358,N_849);
nor U2885 (N_2885,N_366,N_186);
nor U2886 (N_2886,N_1234,N_1198);
and U2887 (N_2887,N_1525,N_1569);
nor U2888 (N_2888,N_119,N_1311);
nor U2889 (N_2889,N_333,N_787);
nor U2890 (N_2890,N_1181,N_1228);
and U2891 (N_2891,N_1086,N_1035);
and U2892 (N_2892,N_246,N_1607);
and U2893 (N_2893,N_1572,N_1944);
nor U2894 (N_2894,N_1340,N_899);
nand U2895 (N_2895,N_623,N_29);
nand U2896 (N_2896,N_1078,N_1970);
nand U2897 (N_2897,N_880,N_1076);
or U2898 (N_2898,N_482,N_964);
nand U2899 (N_2899,N_900,N_640);
nor U2900 (N_2900,N_31,N_664);
nor U2901 (N_2901,N_1548,N_519);
and U2902 (N_2902,N_344,N_730);
nor U2903 (N_2903,N_936,N_641);
nand U2904 (N_2904,N_1566,N_432);
nand U2905 (N_2905,N_707,N_1957);
and U2906 (N_2906,N_1768,N_590);
and U2907 (N_2907,N_42,N_1089);
nor U2908 (N_2908,N_897,N_1778);
or U2909 (N_2909,N_467,N_380);
or U2910 (N_2910,N_361,N_836);
or U2911 (N_2911,N_815,N_1412);
nand U2912 (N_2912,N_1847,N_503);
nand U2913 (N_2913,N_549,N_346);
nor U2914 (N_2914,N_627,N_1757);
and U2915 (N_2915,N_1553,N_434);
nand U2916 (N_2916,N_1936,N_130);
nand U2917 (N_2917,N_1063,N_928);
or U2918 (N_2918,N_1952,N_858);
or U2919 (N_2919,N_1103,N_420);
or U2920 (N_2920,N_1333,N_617);
and U2921 (N_2921,N_1159,N_1130);
and U2922 (N_2922,N_356,N_537);
nor U2923 (N_2923,N_659,N_1120);
nand U2924 (N_2924,N_1892,N_1842);
or U2925 (N_2925,N_868,N_396);
nand U2926 (N_2926,N_585,N_351);
or U2927 (N_2927,N_950,N_548);
nor U2928 (N_2928,N_1047,N_1275);
nand U2929 (N_2929,N_1503,N_1945);
and U2930 (N_2930,N_1851,N_1226);
or U2931 (N_2931,N_867,N_719);
and U2932 (N_2932,N_1905,N_99);
nor U2933 (N_2933,N_1504,N_670);
or U2934 (N_2934,N_1853,N_653);
nand U2935 (N_2935,N_1147,N_1068);
nor U2936 (N_2936,N_859,N_948);
or U2937 (N_2937,N_534,N_85);
nor U2938 (N_2938,N_628,N_1151);
nand U2939 (N_2939,N_1059,N_680);
nand U2940 (N_2940,N_812,N_324);
nand U2941 (N_2941,N_164,N_1790);
nor U2942 (N_2942,N_1060,N_1231);
or U2943 (N_2943,N_54,N_74);
xor U2944 (N_2944,N_1850,N_596);
nor U2945 (N_2945,N_931,N_926);
or U2946 (N_2946,N_439,N_369);
nor U2947 (N_2947,N_1737,N_1382);
nor U2948 (N_2948,N_310,N_1413);
nand U2949 (N_2949,N_1065,N_1667);
nand U2950 (N_2950,N_1714,N_431);
nor U2951 (N_2951,N_1618,N_83);
or U2952 (N_2952,N_902,N_1158);
nand U2953 (N_2953,N_1869,N_402);
nor U2954 (N_2954,N_1623,N_288);
or U2955 (N_2955,N_1662,N_1360);
nand U2956 (N_2956,N_238,N_1639);
nor U2957 (N_2957,N_1214,N_1064);
nor U2958 (N_2958,N_1481,N_298);
or U2959 (N_2959,N_30,N_550);
or U2960 (N_2960,N_1307,N_1789);
or U2961 (N_2961,N_474,N_1746);
and U2962 (N_2962,N_1426,N_1213);
nand U2963 (N_2963,N_1808,N_1976);
nand U2964 (N_2964,N_1706,N_872);
nor U2965 (N_2965,N_1478,N_175);
xor U2966 (N_2966,N_741,N_1347);
nand U2967 (N_2967,N_892,N_157);
nor U2968 (N_2968,N_728,N_1803);
or U2969 (N_2969,N_685,N_1831);
and U2970 (N_2970,N_733,N_1336);
nor U2971 (N_2971,N_378,N_1441);
nor U2972 (N_2972,N_1282,N_1920);
or U2973 (N_2973,N_1245,N_1323);
and U2974 (N_2974,N_258,N_656);
or U2975 (N_2975,N_955,N_1683);
nand U2976 (N_2976,N_32,N_735);
and U2977 (N_2977,N_1611,N_1684);
or U2978 (N_2978,N_1859,N_1520);
or U2979 (N_2979,N_1138,N_543);
nand U2980 (N_2980,N_1139,N_1818);
nand U2981 (N_2981,N_980,N_1813);
nor U2982 (N_2982,N_781,N_221);
nor U2983 (N_2983,N_255,N_1366);
nor U2984 (N_2984,N_566,N_633);
nand U2985 (N_2985,N_676,N_1421);
and U2986 (N_2986,N_1923,N_1536);
nand U2987 (N_2987,N_1030,N_1084);
nand U2988 (N_2988,N_274,N_774);
or U2989 (N_2989,N_960,N_1237);
nor U2990 (N_2990,N_323,N_270);
nor U2991 (N_2991,N_1846,N_1775);
or U2992 (N_2992,N_1666,N_496);
or U2993 (N_2993,N_353,N_983);
and U2994 (N_2994,N_133,N_686);
and U2995 (N_2995,N_1615,N_1577);
and U2996 (N_2996,N_415,N_45);
and U2997 (N_2997,N_1654,N_961);
or U2998 (N_2998,N_1908,N_249);
and U2999 (N_2999,N_1975,N_1090);
or U3000 (N_3000,N_1896,N_1277);
and U3001 (N_3001,N_1837,N_1960);
or U3002 (N_3002,N_37,N_140);
nand U3003 (N_3003,N_1743,N_1862);
nand U3004 (N_3004,N_903,N_34);
nand U3005 (N_3005,N_54,N_899);
or U3006 (N_3006,N_1533,N_1805);
nand U3007 (N_3007,N_1176,N_1824);
nand U3008 (N_3008,N_1934,N_1621);
and U3009 (N_3009,N_1612,N_526);
or U3010 (N_3010,N_63,N_1400);
nand U3011 (N_3011,N_1384,N_793);
nor U3012 (N_3012,N_924,N_105);
and U3013 (N_3013,N_1808,N_953);
or U3014 (N_3014,N_37,N_677);
nand U3015 (N_3015,N_1835,N_1472);
and U3016 (N_3016,N_965,N_1634);
and U3017 (N_3017,N_386,N_399);
nand U3018 (N_3018,N_204,N_721);
or U3019 (N_3019,N_1811,N_428);
nor U3020 (N_3020,N_624,N_1288);
nand U3021 (N_3021,N_659,N_281);
nand U3022 (N_3022,N_353,N_1878);
and U3023 (N_3023,N_1087,N_1138);
nor U3024 (N_3024,N_1193,N_912);
nand U3025 (N_3025,N_159,N_1140);
or U3026 (N_3026,N_1844,N_1197);
or U3027 (N_3027,N_1732,N_614);
or U3028 (N_3028,N_51,N_1018);
nor U3029 (N_3029,N_1423,N_1144);
and U3030 (N_3030,N_873,N_356);
nor U3031 (N_3031,N_735,N_710);
and U3032 (N_3032,N_1338,N_1410);
nor U3033 (N_3033,N_402,N_1362);
or U3034 (N_3034,N_850,N_1090);
nand U3035 (N_3035,N_1965,N_521);
or U3036 (N_3036,N_1137,N_299);
nand U3037 (N_3037,N_1305,N_1293);
nor U3038 (N_3038,N_980,N_43);
nand U3039 (N_3039,N_1437,N_414);
and U3040 (N_3040,N_442,N_1348);
or U3041 (N_3041,N_1316,N_1130);
nand U3042 (N_3042,N_469,N_447);
nor U3043 (N_3043,N_483,N_157);
nand U3044 (N_3044,N_1525,N_1765);
or U3045 (N_3045,N_429,N_15);
and U3046 (N_3046,N_839,N_105);
or U3047 (N_3047,N_302,N_1396);
nor U3048 (N_3048,N_902,N_1796);
nor U3049 (N_3049,N_1220,N_459);
or U3050 (N_3050,N_1025,N_961);
or U3051 (N_3051,N_722,N_337);
or U3052 (N_3052,N_535,N_224);
nor U3053 (N_3053,N_963,N_1048);
nand U3054 (N_3054,N_1751,N_51);
nor U3055 (N_3055,N_1511,N_792);
xor U3056 (N_3056,N_847,N_1012);
or U3057 (N_3057,N_631,N_1070);
or U3058 (N_3058,N_503,N_1939);
and U3059 (N_3059,N_512,N_1610);
nand U3060 (N_3060,N_1224,N_1424);
nor U3061 (N_3061,N_220,N_980);
nand U3062 (N_3062,N_893,N_355);
or U3063 (N_3063,N_1184,N_1611);
nand U3064 (N_3064,N_1364,N_421);
xnor U3065 (N_3065,N_577,N_97);
nor U3066 (N_3066,N_1731,N_684);
nor U3067 (N_3067,N_636,N_1190);
nand U3068 (N_3068,N_265,N_426);
and U3069 (N_3069,N_1905,N_464);
nand U3070 (N_3070,N_1046,N_150);
nand U3071 (N_3071,N_1970,N_540);
nand U3072 (N_3072,N_1467,N_1338);
or U3073 (N_3073,N_1885,N_241);
nand U3074 (N_3074,N_1357,N_287);
nor U3075 (N_3075,N_1941,N_1926);
and U3076 (N_3076,N_1579,N_1539);
or U3077 (N_3077,N_1648,N_448);
and U3078 (N_3078,N_1339,N_693);
nand U3079 (N_3079,N_836,N_959);
nand U3080 (N_3080,N_1010,N_1012);
and U3081 (N_3081,N_1278,N_242);
nor U3082 (N_3082,N_67,N_991);
nor U3083 (N_3083,N_525,N_158);
or U3084 (N_3084,N_1944,N_653);
or U3085 (N_3085,N_1008,N_1044);
nand U3086 (N_3086,N_1753,N_181);
and U3087 (N_3087,N_1520,N_849);
and U3088 (N_3088,N_1352,N_1580);
or U3089 (N_3089,N_320,N_1453);
nor U3090 (N_3090,N_373,N_1170);
and U3091 (N_3091,N_180,N_18);
or U3092 (N_3092,N_49,N_402);
nor U3093 (N_3093,N_1584,N_1745);
nand U3094 (N_3094,N_291,N_65);
nand U3095 (N_3095,N_1615,N_1694);
nand U3096 (N_3096,N_435,N_1216);
nand U3097 (N_3097,N_1364,N_347);
or U3098 (N_3098,N_1917,N_406);
and U3099 (N_3099,N_48,N_1493);
nor U3100 (N_3100,N_1532,N_629);
or U3101 (N_3101,N_1681,N_101);
or U3102 (N_3102,N_290,N_1519);
nor U3103 (N_3103,N_1534,N_688);
or U3104 (N_3104,N_987,N_1781);
and U3105 (N_3105,N_28,N_881);
nor U3106 (N_3106,N_1354,N_749);
nor U3107 (N_3107,N_1933,N_1179);
and U3108 (N_3108,N_1377,N_1403);
and U3109 (N_3109,N_762,N_345);
or U3110 (N_3110,N_322,N_251);
and U3111 (N_3111,N_1725,N_250);
nor U3112 (N_3112,N_480,N_1153);
nand U3113 (N_3113,N_1472,N_1941);
or U3114 (N_3114,N_546,N_910);
nand U3115 (N_3115,N_345,N_376);
and U3116 (N_3116,N_972,N_1671);
nand U3117 (N_3117,N_1102,N_238);
nor U3118 (N_3118,N_703,N_1221);
and U3119 (N_3119,N_1548,N_655);
and U3120 (N_3120,N_1245,N_973);
nor U3121 (N_3121,N_1041,N_1574);
and U3122 (N_3122,N_520,N_1242);
nand U3123 (N_3123,N_1644,N_1912);
and U3124 (N_3124,N_1842,N_1519);
nor U3125 (N_3125,N_434,N_1910);
nor U3126 (N_3126,N_951,N_204);
nor U3127 (N_3127,N_559,N_578);
nor U3128 (N_3128,N_1974,N_94);
and U3129 (N_3129,N_1148,N_818);
nor U3130 (N_3130,N_1141,N_952);
or U3131 (N_3131,N_1137,N_139);
nor U3132 (N_3132,N_507,N_1189);
nand U3133 (N_3133,N_1156,N_1996);
nor U3134 (N_3134,N_688,N_1106);
and U3135 (N_3135,N_999,N_243);
and U3136 (N_3136,N_690,N_894);
or U3137 (N_3137,N_1002,N_1837);
and U3138 (N_3138,N_1861,N_1650);
or U3139 (N_3139,N_149,N_1574);
or U3140 (N_3140,N_584,N_1002);
nor U3141 (N_3141,N_803,N_1290);
and U3142 (N_3142,N_1437,N_938);
and U3143 (N_3143,N_189,N_696);
nand U3144 (N_3144,N_1207,N_91);
and U3145 (N_3145,N_728,N_809);
and U3146 (N_3146,N_619,N_811);
nand U3147 (N_3147,N_1520,N_285);
nor U3148 (N_3148,N_85,N_1096);
and U3149 (N_3149,N_880,N_1742);
and U3150 (N_3150,N_750,N_1243);
or U3151 (N_3151,N_1020,N_1348);
nand U3152 (N_3152,N_76,N_1705);
and U3153 (N_3153,N_651,N_1197);
and U3154 (N_3154,N_1462,N_1211);
xnor U3155 (N_3155,N_1586,N_424);
or U3156 (N_3156,N_1334,N_1313);
and U3157 (N_3157,N_740,N_417);
nor U3158 (N_3158,N_607,N_1443);
and U3159 (N_3159,N_218,N_215);
and U3160 (N_3160,N_1886,N_1490);
or U3161 (N_3161,N_6,N_1448);
or U3162 (N_3162,N_764,N_332);
and U3163 (N_3163,N_440,N_145);
nand U3164 (N_3164,N_1476,N_36);
xor U3165 (N_3165,N_1345,N_196);
or U3166 (N_3166,N_1081,N_1667);
nand U3167 (N_3167,N_782,N_1737);
nand U3168 (N_3168,N_1589,N_846);
nand U3169 (N_3169,N_131,N_536);
xnor U3170 (N_3170,N_547,N_1787);
and U3171 (N_3171,N_322,N_1867);
and U3172 (N_3172,N_1026,N_760);
or U3173 (N_3173,N_1350,N_1165);
nor U3174 (N_3174,N_518,N_14);
nand U3175 (N_3175,N_579,N_337);
or U3176 (N_3176,N_1444,N_1148);
nor U3177 (N_3177,N_839,N_1091);
or U3178 (N_3178,N_616,N_1937);
nand U3179 (N_3179,N_703,N_534);
and U3180 (N_3180,N_1644,N_1520);
nor U3181 (N_3181,N_1924,N_628);
nor U3182 (N_3182,N_645,N_1182);
or U3183 (N_3183,N_1442,N_1942);
nor U3184 (N_3184,N_402,N_1822);
nor U3185 (N_3185,N_1836,N_218);
nor U3186 (N_3186,N_789,N_906);
or U3187 (N_3187,N_235,N_1776);
nand U3188 (N_3188,N_715,N_1009);
nor U3189 (N_3189,N_184,N_742);
and U3190 (N_3190,N_1285,N_1805);
or U3191 (N_3191,N_1907,N_769);
nand U3192 (N_3192,N_1823,N_922);
nand U3193 (N_3193,N_192,N_1023);
and U3194 (N_3194,N_1366,N_877);
and U3195 (N_3195,N_1097,N_1824);
nor U3196 (N_3196,N_1154,N_1280);
nand U3197 (N_3197,N_46,N_854);
and U3198 (N_3198,N_230,N_741);
nand U3199 (N_3199,N_880,N_975);
nor U3200 (N_3200,N_409,N_1129);
xnor U3201 (N_3201,N_420,N_1802);
nor U3202 (N_3202,N_1412,N_1603);
nand U3203 (N_3203,N_1987,N_870);
and U3204 (N_3204,N_554,N_1701);
nor U3205 (N_3205,N_177,N_1085);
or U3206 (N_3206,N_1565,N_391);
or U3207 (N_3207,N_473,N_1030);
nor U3208 (N_3208,N_1456,N_462);
and U3209 (N_3209,N_1256,N_1323);
nand U3210 (N_3210,N_859,N_186);
nor U3211 (N_3211,N_805,N_1228);
nor U3212 (N_3212,N_181,N_1203);
nand U3213 (N_3213,N_1958,N_1737);
nand U3214 (N_3214,N_226,N_1440);
nand U3215 (N_3215,N_379,N_389);
or U3216 (N_3216,N_502,N_1970);
and U3217 (N_3217,N_1506,N_729);
xor U3218 (N_3218,N_1063,N_288);
nor U3219 (N_3219,N_385,N_1721);
nand U3220 (N_3220,N_141,N_1125);
nand U3221 (N_3221,N_498,N_210);
and U3222 (N_3222,N_231,N_1864);
or U3223 (N_3223,N_1795,N_419);
and U3224 (N_3224,N_440,N_97);
and U3225 (N_3225,N_895,N_19);
nand U3226 (N_3226,N_1105,N_594);
nor U3227 (N_3227,N_186,N_21);
nand U3228 (N_3228,N_109,N_973);
or U3229 (N_3229,N_517,N_978);
or U3230 (N_3230,N_1284,N_958);
nor U3231 (N_3231,N_1361,N_452);
and U3232 (N_3232,N_1152,N_990);
nor U3233 (N_3233,N_1042,N_1010);
nor U3234 (N_3234,N_1047,N_465);
nand U3235 (N_3235,N_1601,N_964);
nor U3236 (N_3236,N_530,N_538);
nor U3237 (N_3237,N_1030,N_914);
or U3238 (N_3238,N_1003,N_242);
and U3239 (N_3239,N_1851,N_1048);
or U3240 (N_3240,N_1292,N_1148);
and U3241 (N_3241,N_1742,N_227);
nor U3242 (N_3242,N_507,N_1552);
xor U3243 (N_3243,N_1186,N_974);
nor U3244 (N_3244,N_1931,N_365);
and U3245 (N_3245,N_1793,N_878);
or U3246 (N_3246,N_937,N_642);
or U3247 (N_3247,N_1653,N_960);
or U3248 (N_3248,N_1245,N_1049);
or U3249 (N_3249,N_900,N_972);
nor U3250 (N_3250,N_1848,N_1049);
nand U3251 (N_3251,N_1251,N_714);
and U3252 (N_3252,N_1937,N_256);
and U3253 (N_3253,N_483,N_353);
and U3254 (N_3254,N_1649,N_356);
or U3255 (N_3255,N_483,N_1355);
nor U3256 (N_3256,N_1724,N_309);
or U3257 (N_3257,N_266,N_819);
nor U3258 (N_3258,N_1280,N_347);
nor U3259 (N_3259,N_911,N_700);
or U3260 (N_3260,N_99,N_922);
nor U3261 (N_3261,N_29,N_1453);
or U3262 (N_3262,N_607,N_232);
or U3263 (N_3263,N_856,N_141);
and U3264 (N_3264,N_790,N_609);
nand U3265 (N_3265,N_879,N_338);
nor U3266 (N_3266,N_1785,N_901);
nand U3267 (N_3267,N_485,N_518);
nand U3268 (N_3268,N_950,N_239);
or U3269 (N_3269,N_80,N_342);
or U3270 (N_3270,N_296,N_1557);
nand U3271 (N_3271,N_1273,N_1335);
nand U3272 (N_3272,N_623,N_233);
or U3273 (N_3273,N_556,N_1938);
nand U3274 (N_3274,N_877,N_958);
nor U3275 (N_3275,N_1271,N_1548);
or U3276 (N_3276,N_276,N_380);
nor U3277 (N_3277,N_1643,N_943);
nand U3278 (N_3278,N_1784,N_1097);
nand U3279 (N_3279,N_534,N_1653);
or U3280 (N_3280,N_1553,N_1546);
nor U3281 (N_3281,N_1697,N_111);
nor U3282 (N_3282,N_1081,N_344);
and U3283 (N_3283,N_1236,N_935);
xnor U3284 (N_3284,N_1344,N_539);
or U3285 (N_3285,N_125,N_1919);
or U3286 (N_3286,N_1740,N_721);
or U3287 (N_3287,N_1615,N_1103);
nor U3288 (N_3288,N_1541,N_402);
xor U3289 (N_3289,N_1291,N_564);
nand U3290 (N_3290,N_1202,N_1216);
nand U3291 (N_3291,N_1265,N_1034);
or U3292 (N_3292,N_1847,N_666);
and U3293 (N_3293,N_608,N_398);
and U3294 (N_3294,N_488,N_573);
xor U3295 (N_3295,N_1431,N_1717);
nand U3296 (N_3296,N_731,N_670);
or U3297 (N_3297,N_565,N_1622);
or U3298 (N_3298,N_1108,N_130);
and U3299 (N_3299,N_1870,N_1650);
nor U3300 (N_3300,N_1640,N_146);
nor U3301 (N_3301,N_93,N_1168);
nand U3302 (N_3302,N_276,N_1197);
nor U3303 (N_3303,N_87,N_369);
and U3304 (N_3304,N_1407,N_597);
or U3305 (N_3305,N_192,N_811);
nor U3306 (N_3306,N_51,N_497);
nor U3307 (N_3307,N_1294,N_1544);
and U3308 (N_3308,N_1728,N_739);
and U3309 (N_3309,N_1144,N_115);
nand U3310 (N_3310,N_178,N_1144);
and U3311 (N_3311,N_190,N_933);
nand U3312 (N_3312,N_998,N_1402);
and U3313 (N_3313,N_1085,N_1790);
and U3314 (N_3314,N_567,N_1196);
and U3315 (N_3315,N_1175,N_1708);
or U3316 (N_3316,N_732,N_1804);
and U3317 (N_3317,N_168,N_373);
nor U3318 (N_3318,N_1943,N_1198);
nor U3319 (N_3319,N_765,N_1985);
nand U3320 (N_3320,N_484,N_989);
or U3321 (N_3321,N_807,N_137);
and U3322 (N_3322,N_1553,N_158);
nor U3323 (N_3323,N_1638,N_855);
or U3324 (N_3324,N_1579,N_1914);
or U3325 (N_3325,N_1946,N_229);
and U3326 (N_3326,N_1531,N_1806);
or U3327 (N_3327,N_486,N_771);
or U3328 (N_3328,N_1917,N_1878);
nor U3329 (N_3329,N_1997,N_1760);
nand U3330 (N_3330,N_1591,N_1347);
nor U3331 (N_3331,N_47,N_992);
and U3332 (N_3332,N_589,N_1949);
or U3333 (N_3333,N_359,N_1260);
nor U3334 (N_3334,N_594,N_765);
nand U3335 (N_3335,N_1903,N_838);
nor U3336 (N_3336,N_388,N_1116);
and U3337 (N_3337,N_627,N_1904);
or U3338 (N_3338,N_269,N_284);
nor U3339 (N_3339,N_290,N_744);
nor U3340 (N_3340,N_591,N_196);
and U3341 (N_3341,N_1308,N_85);
and U3342 (N_3342,N_241,N_317);
or U3343 (N_3343,N_1785,N_1959);
nor U3344 (N_3344,N_1746,N_632);
or U3345 (N_3345,N_1445,N_1997);
or U3346 (N_3346,N_1302,N_838);
and U3347 (N_3347,N_113,N_498);
nor U3348 (N_3348,N_1827,N_616);
and U3349 (N_3349,N_57,N_1280);
or U3350 (N_3350,N_1222,N_1523);
nand U3351 (N_3351,N_1928,N_885);
and U3352 (N_3352,N_1774,N_1688);
nand U3353 (N_3353,N_1089,N_203);
or U3354 (N_3354,N_262,N_895);
nand U3355 (N_3355,N_422,N_1346);
or U3356 (N_3356,N_557,N_1509);
nor U3357 (N_3357,N_1142,N_328);
nand U3358 (N_3358,N_1366,N_1556);
nand U3359 (N_3359,N_753,N_336);
and U3360 (N_3360,N_1658,N_1632);
xnor U3361 (N_3361,N_746,N_1575);
and U3362 (N_3362,N_789,N_1951);
nor U3363 (N_3363,N_1807,N_602);
nor U3364 (N_3364,N_1057,N_164);
nand U3365 (N_3365,N_1065,N_741);
or U3366 (N_3366,N_1586,N_920);
and U3367 (N_3367,N_555,N_1246);
and U3368 (N_3368,N_117,N_991);
nor U3369 (N_3369,N_138,N_1729);
or U3370 (N_3370,N_627,N_1690);
nor U3371 (N_3371,N_703,N_1882);
nand U3372 (N_3372,N_1639,N_322);
nand U3373 (N_3373,N_6,N_169);
and U3374 (N_3374,N_1799,N_1273);
or U3375 (N_3375,N_1853,N_40);
or U3376 (N_3376,N_1759,N_367);
and U3377 (N_3377,N_896,N_1632);
or U3378 (N_3378,N_288,N_1513);
nand U3379 (N_3379,N_274,N_1001);
nand U3380 (N_3380,N_1915,N_560);
nand U3381 (N_3381,N_1726,N_1565);
or U3382 (N_3382,N_1901,N_1834);
and U3383 (N_3383,N_837,N_1318);
nor U3384 (N_3384,N_1101,N_1426);
xnor U3385 (N_3385,N_1261,N_1199);
nand U3386 (N_3386,N_1660,N_118);
or U3387 (N_3387,N_1193,N_498);
or U3388 (N_3388,N_1484,N_161);
and U3389 (N_3389,N_1134,N_1768);
nor U3390 (N_3390,N_985,N_1473);
nand U3391 (N_3391,N_1613,N_1798);
or U3392 (N_3392,N_1647,N_967);
nor U3393 (N_3393,N_172,N_309);
and U3394 (N_3394,N_322,N_1743);
and U3395 (N_3395,N_455,N_1915);
and U3396 (N_3396,N_1053,N_686);
nand U3397 (N_3397,N_216,N_1311);
and U3398 (N_3398,N_1288,N_372);
nand U3399 (N_3399,N_1359,N_1732);
nand U3400 (N_3400,N_1882,N_589);
and U3401 (N_3401,N_1505,N_1934);
and U3402 (N_3402,N_1370,N_1103);
or U3403 (N_3403,N_1973,N_348);
or U3404 (N_3404,N_1185,N_652);
nand U3405 (N_3405,N_555,N_264);
and U3406 (N_3406,N_1273,N_741);
nand U3407 (N_3407,N_1588,N_1888);
nand U3408 (N_3408,N_1406,N_1842);
and U3409 (N_3409,N_620,N_398);
nand U3410 (N_3410,N_444,N_652);
and U3411 (N_3411,N_934,N_596);
nor U3412 (N_3412,N_679,N_1574);
nor U3413 (N_3413,N_1137,N_1783);
and U3414 (N_3414,N_265,N_157);
or U3415 (N_3415,N_174,N_285);
and U3416 (N_3416,N_291,N_505);
nand U3417 (N_3417,N_1055,N_858);
nand U3418 (N_3418,N_85,N_974);
nand U3419 (N_3419,N_129,N_1445);
nand U3420 (N_3420,N_744,N_1740);
or U3421 (N_3421,N_1552,N_1296);
and U3422 (N_3422,N_1862,N_348);
or U3423 (N_3423,N_1016,N_1375);
nand U3424 (N_3424,N_1660,N_1907);
nor U3425 (N_3425,N_1893,N_1699);
and U3426 (N_3426,N_574,N_1917);
and U3427 (N_3427,N_750,N_966);
nand U3428 (N_3428,N_1012,N_1439);
and U3429 (N_3429,N_1831,N_323);
nand U3430 (N_3430,N_732,N_1037);
nor U3431 (N_3431,N_207,N_45);
nor U3432 (N_3432,N_1357,N_219);
nor U3433 (N_3433,N_1112,N_1783);
nor U3434 (N_3434,N_424,N_1217);
or U3435 (N_3435,N_1980,N_14);
nor U3436 (N_3436,N_1675,N_1814);
or U3437 (N_3437,N_1921,N_898);
nor U3438 (N_3438,N_189,N_1294);
or U3439 (N_3439,N_1372,N_698);
nand U3440 (N_3440,N_904,N_1394);
or U3441 (N_3441,N_1320,N_800);
nand U3442 (N_3442,N_1085,N_640);
or U3443 (N_3443,N_277,N_928);
and U3444 (N_3444,N_1050,N_1128);
nor U3445 (N_3445,N_1712,N_1365);
nand U3446 (N_3446,N_531,N_1067);
nor U3447 (N_3447,N_978,N_712);
or U3448 (N_3448,N_514,N_489);
nor U3449 (N_3449,N_1252,N_727);
nand U3450 (N_3450,N_706,N_816);
or U3451 (N_3451,N_1546,N_1465);
xnor U3452 (N_3452,N_473,N_155);
and U3453 (N_3453,N_315,N_1562);
nand U3454 (N_3454,N_1919,N_1798);
and U3455 (N_3455,N_651,N_1778);
nand U3456 (N_3456,N_1257,N_1114);
nor U3457 (N_3457,N_1357,N_1929);
and U3458 (N_3458,N_359,N_601);
or U3459 (N_3459,N_293,N_1655);
or U3460 (N_3460,N_1625,N_244);
or U3461 (N_3461,N_110,N_1127);
or U3462 (N_3462,N_1712,N_1864);
and U3463 (N_3463,N_1584,N_1532);
xor U3464 (N_3464,N_862,N_1793);
or U3465 (N_3465,N_1969,N_1844);
nor U3466 (N_3466,N_1566,N_738);
and U3467 (N_3467,N_320,N_446);
and U3468 (N_3468,N_433,N_625);
nand U3469 (N_3469,N_1017,N_256);
nand U3470 (N_3470,N_1417,N_1576);
or U3471 (N_3471,N_75,N_792);
or U3472 (N_3472,N_708,N_422);
nor U3473 (N_3473,N_1285,N_428);
or U3474 (N_3474,N_167,N_1933);
and U3475 (N_3475,N_15,N_501);
nor U3476 (N_3476,N_1724,N_1058);
or U3477 (N_3477,N_163,N_1271);
and U3478 (N_3478,N_177,N_1189);
or U3479 (N_3479,N_524,N_433);
nand U3480 (N_3480,N_381,N_212);
or U3481 (N_3481,N_1786,N_1839);
and U3482 (N_3482,N_1076,N_51);
nand U3483 (N_3483,N_1190,N_520);
and U3484 (N_3484,N_963,N_1800);
and U3485 (N_3485,N_1472,N_1123);
nor U3486 (N_3486,N_1499,N_875);
nor U3487 (N_3487,N_1360,N_1899);
and U3488 (N_3488,N_1906,N_1560);
and U3489 (N_3489,N_467,N_935);
nor U3490 (N_3490,N_1670,N_452);
or U3491 (N_3491,N_1016,N_1207);
nand U3492 (N_3492,N_1959,N_79);
nand U3493 (N_3493,N_1582,N_376);
or U3494 (N_3494,N_1681,N_811);
and U3495 (N_3495,N_1262,N_48);
nand U3496 (N_3496,N_1781,N_814);
and U3497 (N_3497,N_663,N_700);
nand U3498 (N_3498,N_541,N_898);
nand U3499 (N_3499,N_1622,N_1324);
and U3500 (N_3500,N_519,N_772);
and U3501 (N_3501,N_305,N_1735);
and U3502 (N_3502,N_1681,N_882);
nand U3503 (N_3503,N_1453,N_446);
nand U3504 (N_3504,N_777,N_1998);
nand U3505 (N_3505,N_1579,N_1315);
nand U3506 (N_3506,N_1458,N_1277);
nand U3507 (N_3507,N_1194,N_345);
and U3508 (N_3508,N_508,N_618);
and U3509 (N_3509,N_988,N_787);
and U3510 (N_3510,N_1450,N_126);
nand U3511 (N_3511,N_386,N_1335);
nand U3512 (N_3512,N_684,N_1253);
nand U3513 (N_3513,N_1704,N_368);
or U3514 (N_3514,N_780,N_35);
nor U3515 (N_3515,N_777,N_747);
and U3516 (N_3516,N_817,N_1466);
nand U3517 (N_3517,N_1584,N_492);
nand U3518 (N_3518,N_1622,N_56);
or U3519 (N_3519,N_1360,N_1756);
nor U3520 (N_3520,N_1634,N_287);
nand U3521 (N_3521,N_1823,N_1637);
or U3522 (N_3522,N_354,N_696);
or U3523 (N_3523,N_1939,N_1183);
or U3524 (N_3524,N_1363,N_1742);
nor U3525 (N_3525,N_1088,N_1190);
nor U3526 (N_3526,N_547,N_1222);
or U3527 (N_3527,N_1762,N_539);
nand U3528 (N_3528,N_1512,N_1511);
nor U3529 (N_3529,N_1396,N_1923);
or U3530 (N_3530,N_690,N_1809);
and U3531 (N_3531,N_1430,N_554);
or U3532 (N_3532,N_1931,N_1234);
and U3533 (N_3533,N_590,N_455);
or U3534 (N_3534,N_1357,N_1485);
nand U3535 (N_3535,N_1948,N_442);
or U3536 (N_3536,N_1021,N_1237);
nor U3537 (N_3537,N_1479,N_534);
or U3538 (N_3538,N_1757,N_1372);
or U3539 (N_3539,N_1849,N_458);
nand U3540 (N_3540,N_1420,N_878);
nor U3541 (N_3541,N_621,N_199);
or U3542 (N_3542,N_117,N_676);
nand U3543 (N_3543,N_851,N_924);
nor U3544 (N_3544,N_390,N_1541);
or U3545 (N_3545,N_1337,N_235);
nand U3546 (N_3546,N_1638,N_689);
and U3547 (N_3547,N_1278,N_1437);
nor U3548 (N_3548,N_1698,N_660);
and U3549 (N_3549,N_370,N_1551);
and U3550 (N_3550,N_1247,N_1516);
nor U3551 (N_3551,N_22,N_794);
nand U3552 (N_3552,N_1279,N_824);
nand U3553 (N_3553,N_1963,N_665);
or U3554 (N_3554,N_530,N_401);
nand U3555 (N_3555,N_1923,N_780);
or U3556 (N_3556,N_126,N_175);
nor U3557 (N_3557,N_611,N_372);
and U3558 (N_3558,N_521,N_249);
and U3559 (N_3559,N_1899,N_702);
or U3560 (N_3560,N_1723,N_1628);
and U3561 (N_3561,N_1644,N_1140);
nand U3562 (N_3562,N_119,N_1219);
or U3563 (N_3563,N_1802,N_165);
and U3564 (N_3564,N_647,N_250);
nor U3565 (N_3565,N_1797,N_702);
nand U3566 (N_3566,N_513,N_1328);
and U3567 (N_3567,N_161,N_1715);
nor U3568 (N_3568,N_1446,N_1590);
or U3569 (N_3569,N_1631,N_770);
and U3570 (N_3570,N_147,N_1695);
or U3571 (N_3571,N_1149,N_1231);
or U3572 (N_3572,N_1988,N_1862);
nor U3573 (N_3573,N_1917,N_637);
or U3574 (N_3574,N_1783,N_1223);
nand U3575 (N_3575,N_1685,N_1794);
or U3576 (N_3576,N_1911,N_639);
nand U3577 (N_3577,N_1051,N_349);
nand U3578 (N_3578,N_14,N_1858);
or U3579 (N_3579,N_220,N_630);
nor U3580 (N_3580,N_1187,N_1183);
and U3581 (N_3581,N_692,N_406);
and U3582 (N_3582,N_878,N_973);
or U3583 (N_3583,N_1389,N_1725);
and U3584 (N_3584,N_1721,N_1241);
nor U3585 (N_3585,N_202,N_142);
nand U3586 (N_3586,N_1551,N_494);
nand U3587 (N_3587,N_1849,N_1797);
and U3588 (N_3588,N_669,N_375);
nor U3589 (N_3589,N_1616,N_1745);
or U3590 (N_3590,N_793,N_1747);
and U3591 (N_3591,N_1570,N_1181);
nor U3592 (N_3592,N_882,N_1021);
and U3593 (N_3593,N_634,N_1630);
or U3594 (N_3594,N_52,N_1372);
nor U3595 (N_3595,N_1271,N_1246);
and U3596 (N_3596,N_1926,N_680);
nand U3597 (N_3597,N_1486,N_1235);
and U3598 (N_3598,N_778,N_883);
and U3599 (N_3599,N_1836,N_1018);
and U3600 (N_3600,N_1515,N_1096);
and U3601 (N_3601,N_1278,N_1682);
nand U3602 (N_3602,N_1584,N_498);
or U3603 (N_3603,N_766,N_38);
and U3604 (N_3604,N_523,N_57);
nand U3605 (N_3605,N_493,N_985);
or U3606 (N_3606,N_1981,N_494);
and U3607 (N_3607,N_1472,N_1209);
and U3608 (N_3608,N_429,N_1392);
and U3609 (N_3609,N_501,N_853);
nand U3610 (N_3610,N_1847,N_286);
nor U3611 (N_3611,N_1449,N_644);
nand U3612 (N_3612,N_895,N_373);
or U3613 (N_3613,N_384,N_1418);
nor U3614 (N_3614,N_1405,N_737);
or U3615 (N_3615,N_978,N_1107);
or U3616 (N_3616,N_1215,N_1022);
and U3617 (N_3617,N_1396,N_1979);
nand U3618 (N_3618,N_1612,N_1175);
or U3619 (N_3619,N_1792,N_1669);
xnor U3620 (N_3620,N_1424,N_681);
nand U3621 (N_3621,N_1462,N_1180);
nor U3622 (N_3622,N_649,N_1751);
nand U3623 (N_3623,N_1527,N_1206);
nand U3624 (N_3624,N_23,N_1565);
and U3625 (N_3625,N_1004,N_191);
and U3626 (N_3626,N_1962,N_1884);
nor U3627 (N_3627,N_1236,N_819);
and U3628 (N_3628,N_982,N_319);
and U3629 (N_3629,N_584,N_1593);
and U3630 (N_3630,N_1352,N_527);
nand U3631 (N_3631,N_148,N_245);
or U3632 (N_3632,N_272,N_15);
nor U3633 (N_3633,N_1954,N_905);
and U3634 (N_3634,N_1534,N_1727);
nor U3635 (N_3635,N_518,N_1801);
nor U3636 (N_3636,N_1100,N_1522);
nand U3637 (N_3637,N_1590,N_189);
and U3638 (N_3638,N_1162,N_508);
xor U3639 (N_3639,N_1118,N_773);
nor U3640 (N_3640,N_82,N_1213);
or U3641 (N_3641,N_1669,N_1868);
and U3642 (N_3642,N_1067,N_1967);
nor U3643 (N_3643,N_1310,N_182);
or U3644 (N_3644,N_845,N_888);
nor U3645 (N_3645,N_1993,N_40);
or U3646 (N_3646,N_1426,N_464);
and U3647 (N_3647,N_362,N_1712);
nand U3648 (N_3648,N_1618,N_572);
xor U3649 (N_3649,N_352,N_635);
and U3650 (N_3650,N_177,N_1406);
and U3651 (N_3651,N_1545,N_989);
or U3652 (N_3652,N_115,N_1602);
nand U3653 (N_3653,N_123,N_141);
xor U3654 (N_3654,N_257,N_759);
and U3655 (N_3655,N_1291,N_1143);
xor U3656 (N_3656,N_89,N_1747);
and U3657 (N_3657,N_1413,N_705);
nor U3658 (N_3658,N_403,N_923);
nor U3659 (N_3659,N_1136,N_1348);
and U3660 (N_3660,N_1538,N_726);
and U3661 (N_3661,N_1706,N_463);
and U3662 (N_3662,N_311,N_1086);
nand U3663 (N_3663,N_992,N_1840);
or U3664 (N_3664,N_219,N_1679);
or U3665 (N_3665,N_852,N_1506);
nor U3666 (N_3666,N_452,N_1941);
nand U3667 (N_3667,N_399,N_80);
and U3668 (N_3668,N_1105,N_1145);
nor U3669 (N_3669,N_453,N_639);
or U3670 (N_3670,N_550,N_412);
or U3671 (N_3671,N_1581,N_464);
nor U3672 (N_3672,N_1635,N_1014);
and U3673 (N_3673,N_1036,N_1074);
nor U3674 (N_3674,N_981,N_518);
nor U3675 (N_3675,N_1087,N_919);
nor U3676 (N_3676,N_815,N_372);
or U3677 (N_3677,N_1261,N_592);
and U3678 (N_3678,N_1844,N_1428);
and U3679 (N_3679,N_778,N_571);
nand U3680 (N_3680,N_750,N_771);
nor U3681 (N_3681,N_1186,N_980);
and U3682 (N_3682,N_1055,N_686);
and U3683 (N_3683,N_302,N_521);
nor U3684 (N_3684,N_1359,N_818);
or U3685 (N_3685,N_1846,N_1602);
nand U3686 (N_3686,N_1886,N_151);
nand U3687 (N_3687,N_973,N_1221);
or U3688 (N_3688,N_224,N_825);
nor U3689 (N_3689,N_986,N_733);
nor U3690 (N_3690,N_170,N_1322);
nor U3691 (N_3691,N_1132,N_541);
and U3692 (N_3692,N_1090,N_666);
nor U3693 (N_3693,N_646,N_1427);
and U3694 (N_3694,N_109,N_320);
nand U3695 (N_3695,N_71,N_1760);
nand U3696 (N_3696,N_429,N_1951);
or U3697 (N_3697,N_102,N_798);
or U3698 (N_3698,N_525,N_593);
nand U3699 (N_3699,N_348,N_1212);
and U3700 (N_3700,N_411,N_407);
nor U3701 (N_3701,N_1593,N_1633);
nand U3702 (N_3702,N_474,N_1123);
or U3703 (N_3703,N_1213,N_444);
nor U3704 (N_3704,N_142,N_1780);
or U3705 (N_3705,N_347,N_383);
or U3706 (N_3706,N_1097,N_1558);
nand U3707 (N_3707,N_1752,N_820);
nand U3708 (N_3708,N_1728,N_771);
nor U3709 (N_3709,N_836,N_1554);
and U3710 (N_3710,N_622,N_1059);
nand U3711 (N_3711,N_1555,N_1867);
nor U3712 (N_3712,N_1192,N_1591);
or U3713 (N_3713,N_141,N_96);
nand U3714 (N_3714,N_1097,N_1362);
nand U3715 (N_3715,N_1754,N_432);
and U3716 (N_3716,N_311,N_1944);
and U3717 (N_3717,N_1459,N_919);
or U3718 (N_3718,N_151,N_1829);
xor U3719 (N_3719,N_1917,N_1643);
and U3720 (N_3720,N_972,N_981);
and U3721 (N_3721,N_961,N_1109);
nand U3722 (N_3722,N_1232,N_73);
nor U3723 (N_3723,N_802,N_395);
nand U3724 (N_3724,N_203,N_1955);
and U3725 (N_3725,N_1663,N_289);
or U3726 (N_3726,N_1022,N_1162);
and U3727 (N_3727,N_1551,N_976);
nand U3728 (N_3728,N_384,N_1563);
nor U3729 (N_3729,N_1,N_551);
nor U3730 (N_3730,N_1879,N_1445);
and U3731 (N_3731,N_807,N_1699);
nand U3732 (N_3732,N_1080,N_126);
or U3733 (N_3733,N_596,N_18);
nand U3734 (N_3734,N_833,N_213);
nand U3735 (N_3735,N_1437,N_1785);
nor U3736 (N_3736,N_1757,N_950);
and U3737 (N_3737,N_1139,N_903);
and U3738 (N_3738,N_1523,N_1502);
nand U3739 (N_3739,N_1342,N_1891);
nor U3740 (N_3740,N_254,N_492);
or U3741 (N_3741,N_788,N_1021);
xnor U3742 (N_3742,N_746,N_206);
nand U3743 (N_3743,N_678,N_1347);
nor U3744 (N_3744,N_1780,N_279);
nor U3745 (N_3745,N_1188,N_165);
and U3746 (N_3746,N_1450,N_347);
and U3747 (N_3747,N_818,N_607);
or U3748 (N_3748,N_1311,N_1537);
nor U3749 (N_3749,N_639,N_214);
or U3750 (N_3750,N_1739,N_113);
and U3751 (N_3751,N_1006,N_834);
nand U3752 (N_3752,N_1402,N_1468);
or U3753 (N_3753,N_901,N_1764);
or U3754 (N_3754,N_1082,N_87);
nor U3755 (N_3755,N_334,N_466);
nand U3756 (N_3756,N_614,N_1046);
and U3757 (N_3757,N_628,N_408);
xnor U3758 (N_3758,N_170,N_419);
nor U3759 (N_3759,N_1288,N_824);
and U3760 (N_3760,N_1851,N_1947);
nand U3761 (N_3761,N_233,N_1151);
nand U3762 (N_3762,N_793,N_792);
or U3763 (N_3763,N_778,N_1678);
or U3764 (N_3764,N_1496,N_49);
and U3765 (N_3765,N_1708,N_1120);
and U3766 (N_3766,N_1719,N_522);
and U3767 (N_3767,N_961,N_706);
and U3768 (N_3768,N_414,N_1073);
or U3769 (N_3769,N_892,N_418);
and U3770 (N_3770,N_1329,N_396);
and U3771 (N_3771,N_789,N_1805);
nand U3772 (N_3772,N_747,N_678);
nor U3773 (N_3773,N_1104,N_130);
nor U3774 (N_3774,N_1054,N_399);
and U3775 (N_3775,N_1656,N_605);
or U3776 (N_3776,N_338,N_1811);
xnor U3777 (N_3777,N_205,N_945);
nand U3778 (N_3778,N_1314,N_524);
nor U3779 (N_3779,N_178,N_403);
nand U3780 (N_3780,N_1475,N_1065);
nor U3781 (N_3781,N_1755,N_1295);
or U3782 (N_3782,N_773,N_1777);
nor U3783 (N_3783,N_1211,N_1703);
or U3784 (N_3784,N_607,N_1471);
nand U3785 (N_3785,N_568,N_1295);
nor U3786 (N_3786,N_1284,N_534);
nand U3787 (N_3787,N_99,N_1312);
nand U3788 (N_3788,N_1822,N_1364);
xnor U3789 (N_3789,N_1094,N_305);
or U3790 (N_3790,N_1871,N_1345);
nor U3791 (N_3791,N_1342,N_105);
nand U3792 (N_3792,N_391,N_1107);
and U3793 (N_3793,N_1961,N_805);
and U3794 (N_3794,N_1438,N_1364);
or U3795 (N_3795,N_45,N_1059);
nand U3796 (N_3796,N_76,N_1468);
and U3797 (N_3797,N_1209,N_1460);
nand U3798 (N_3798,N_581,N_520);
or U3799 (N_3799,N_866,N_1118);
and U3800 (N_3800,N_886,N_1502);
nand U3801 (N_3801,N_685,N_1911);
and U3802 (N_3802,N_977,N_1067);
and U3803 (N_3803,N_90,N_1230);
and U3804 (N_3804,N_1054,N_370);
nor U3805 (N_3805,N_195,N_1120);
nand U3806 (N_3806,N_1902,N_1433);
and U3807 (N_3807,N_601,N_1185);
and U3808 (N_3808,N_571,N_1494);
nand U3809 (N_3809,N_561,N_1391);
xor U3810 (N_3810,N_1610,N_1799);
or U3811 (N_3811,N_787,N_72);
and U3812 (N_3812,N_1191,N_1546);
nand U3813 (N_3813,N_1574,N_822);
and U3814 (N_3814,N_559,N_843);
xnor U3815 (N_3815,N_1798,N_1410);
nor U3816 (N_3816,N_1610,N_1156);
nand U3817 (N_3817,N_12,N_978);
and U3818 (N_3818,N_1710,N_1783);
or U3819 (N_3819,N_1011,N_1845);
nor U3820 (N_3820,N_734,N_452);
and U3821 (N_3821,N_233,N_55);
nand U3822 (N_3822,N_1217,N_758);
and U3823 (N_3823,N_1082,N_1348);
and U3824 (N_3824,N_957,N_513);
or U3825 (N_3825,N_632,N_24);
nor U3826 (N_3826,N_1699,N_214);
and U3827 (N_3827,N_1193,N_1775);
nor U3828 (N_3828,N_413,N_1817);
xnor U3829 (N_3829,N_1003,N_1681);
nor U3830 (N_3830,N_1275,N_1364);
xor U3831 (N_3831,N_440,N_688);
nor U3832 (N_3832,N_254,N_176);
nand U3833 (N_3833,N_313,N_1787);
nor U3834 (N_3834,N_152,N_1658);
or U3835 (N_3835,N_377,N_1453);
or U3836 (N_3836,N_1711,N_621);
or U3837 (N_3837,N_1164,N_629);
and U3838 (N_3838,N_533,N_876);
or U3839 (N_3839,N_862,N_679);
or U3840 (N_3840,N_1285,N_399);
nor U3841 (N_3841,N_1131,N_1321);
and U3842 (N_3842,N_1887,N_26);
and U3843 (N_3843,N_1996,N_58);
nand U3844 (N_3844,N_1812,N_953);
and U3845 (N_3845,N_1532,N_1558);
nand U3846 (N_3846,N_880,N_1710);
nand U3847 (N_3847,N_1955,N_1703);
and U3848 (N_3848,N_1131,N_851);
nand U3849 (N_3849,N_131,N_777);
nor U3850 (N_3850,N_1401,N_1602);
and U3851 (N_3851,N_1054,N_300);
nor U3852 (N_3852,N_1964,N_1676);
nor U3853 (N_3853,N_155,N_1982);
nand U3854 (N_3854,N_1324,N_1529);
nand U3855 (N_3855,N_585,N_1907);
and U3856 (N_3856,N_1613,N_939);
and U3857 (N_3857,N_1671,N_1803);
xnor U3858 (N_3858,N_776,N_1656);
and U3859 (N_3859,N_209,N_922);
and U3860 (N_3860,N_1865,N_1125);
nand U3861 (N_3861,N_1052,N_1583);
nor U3862 (N_3862,N_1269,N_1295);
nand U3863 (N_3863,N_1855,N_1084);
or U3864 (N_3864,N_1819,N_575);
or U3865 (N_3865,N_1386,N_483);
xnor U3866 (N_3866,N_1241,N_1566);
and U3867 (N_3867,N_128,N_812);
nor U3868 (N_3868,N_565,N_862);
nor U3869 (N_3869,N_1815,N_1104);
nor U3870 (N_3870,N_412,N_1095);
and U3871 (N_3871,N_1792,N_1466);
nand U3872 (N_3872,N_1225,N_27);
and U3873 (N_3873,N_863,N_1666);
nor U3874 (N_3874,N_1587,N_1582);
or U3875 (N_3875,N_655,N_1230);
or U3876 (N_3876,N_21,N_468);
nand U3877 (N_3877,N_328,N_768);
or U3878 (N_3878,N_1551,N_30);
and U3879 (N_3879,N_800,N_1045);
nand U3880 (N_3880,N_642,N_1604);
nor U3881 (N_3881,N_829,N_1874);
nand U3882 (N_3882,N_938,N_1533);
or U3883 (N_3883,N_222,N_546);
nand U3884 (N_3884,N_1070,N_1773);
or U3885 (N_3885,N_416,N_1546);
and U3886 (N_3886,N_1598,N_1962);
nor U3887 (N_3887,N_300,N_1561);
and U3888 (N_3888,N_1152,N_475);
nor U3889 (N_3889,N_1637,N_1667);
nand U3890 (N_3890,N_1811,N_397);
nand U3891 (N_3891,N_243,N_1223);
and U3892 (N_3892,N_1248,N_1456);
nor U3893 (N_3893,N_210,N_703);
nor U3894 (N_3894,N_886,N_325);
or U3895 (N_3895,N_1021,N_1342);
or U3896 (N_3896,N_225,N_1577);
and U3897 (N_3897,N_8,N_1722);
or U3898 (N_3898,N_1565,N_501);
or U3899 (N_3899,N_1669,N_1908);
and U3900 (N_3900,N_472,N_24);
nand U3901 (N_3901,N_1598,N_1366);
xor U3902 (N_3902,N_563,N_731);
or U3903 (N_3903,N_121,N_1276);
nor U3904 (N_3904,N_1739,N_622);
or U3905 (N_3905,N_906,N_1470);
or U3906 (N_3906,N_388,N_671);
or U3907 (N_3907,N_525,N_811);
nand U3908 (N_3908,N_207,N_496);
nor U3909 (N_3909,N_1794,N_1079);
or U3910 (N_3910,N_1842,N_274);
nor U3911 (N_3911,N_1132,N_507);
or U3912 (N_3912,N_1225,N_849);
or U3913 (N_3913,N_1570,N_1145);
and U3914 (N_3914,N_1774,N_1137);
nand U3915 (N_3915,N_1290,N_1786);
nand U3916 (N_3916,N_980,N_817);
nor U3917 (N_3917,N_874,N_169);
or U3918 (N_3918,N_1122,N_1751);
and U3919 (N_3919,N_225,N_1310);
and U3920 (N_3920,N_1252,N_1564);
nand U3921 (N_3921,N_577,N_650);
and U3922 (N_3922,N_1884,N_1157);
and U3923 (N_3923,N_212,N_1958);
or U3924 (N_3924,N_342,N_757);
nand U3925 (N_3925,N_1488,N_30);
nor U3926 (N_3926,N_258,N_1542);
and U3927 (N_3927,N_280,N_1726);
or U3928 (N_3928,N_1365,N_846);
and U3929 (N_3929,N_232,N_178);
nand U3930 (N_3930,N_1568,N_191);
or U3931 (N_3931,N_281,N_49);
nand U3932 (N_3932,N_1784,N_996);
or U3933 (N_3933,N_1066,N_1654);
nor U3934 (N_3934,N_604,N_459);
nand U3935 (N_3935,N_42,N_40);
and U3936 (N_3936,N_335,N_1568);
or U3937 (N_3937,N_1165,N_1011);
and U3938 (N_3938,N_257,N_691);
nand U3939 (N_3939,N_31,N_1580);
and U3940 (N_3940,N_503,N_1903);
or U3941 (N_3941,N_541,N_1126);
nand U3942 (N_3942,N_1531,N_1254);
nand U3943 (N_3943,N_17,N_78);
nor U3944 (N_3944,N_15,N_1700);
nor U3945 (N_3945,N_1835,N_157);
or U3946 (N_3946,N_1450,N_1275);
xnor U3947 (N_3947,N_1476,N_1741);
nor U3948 (N_3948,N_1798,N_920);
nand U3949 (N_3949,N_44,N_516);
and U3950 (N_3950,N_328,N_1842);
nor U3951 (N_3951,N_1847,N_1678);
or U3952 (N_3952,N_1756,N_177);
and U3953 (N_3953,N_1440,N_1587);
or U3954 (N_3954,N_1791,N_287);
nor U3955 (N_3955,N_132,N_1207);
nand U3956 (N_3956,N_15,N_842);
xnor U3957 (N_3957,N_1004,N_683);
or U3958 (N_3958,N_1953,N_216);
nor U3959 (N_3959,N_1584,N_228);
and U3960 (N_3960,N_533,N_312);
nand U3961 (N_3961,N_1177,N_882);
and U3962 (N_3962,N_19,N_143);
and U3963 (N_3963,N_895,N_1935);
nor U3964 (N_3964,N_1068,N_166);
nand U3965 (N_3965,N_1498,N_1695);
and U3966 (N_3966,N_1912,N_1899);
nor U3967 (N_3967,N_1640,N_872);
nand U3968 (N_3968,N_1508,N_1935);
and U3969 (N_3969,N_1517,N_1112);
nand U3970 (N_3970,N_1867,N_956);
or U3971 (N_3971,N_663,N_613);
nor U3972 (N_3972,N_1297,N_158);
nor U3973 (N_3973,N_352,N_1949);
and U3974 (N_3974,N_230,N_321);
or U3975 (N_3975,N_1945,N_1882);
or U3976 (N_3976,N_1115,N_1449);
nor U3977 (N_3977,N_602,N_147);
nor U3978 (N_3978,N_199,N_532);
or U3979 (N_3979,N_1891,N_603);
nand U3980 (N_3980,N_226,N_1496);
nand U3981 (N_3981,N_263,N_1163);
and U3982 (N_3982,N_221,N_1291);
and U3983 (N_3983,N_1782,N_1960);
and U3984 (N_3984,N_814,N_1380);
and U3985 (N_3985,N_971,N_167);
and U3986 (N_3986,N_281,N_507);
and U3987 (N_3987,N_1177,N_692);
or U3988 (N_3988,N_1509,N_242);
nor U3989 (N_3989,N_1183,N_1962);
or U3990 (N_3990,N_932,N_1425);
nand U3991 (N_3991,N_840,N_86);
or U3992 (N_3992,N_1047,N_520);
and U3993 (N_3993,N_1497,N_449);
and U3994 (N_3994,N_1893,N_1187);
or U3995 (N_3995,N_1247,N_1862);
or U3996 (N_3996,N_1065,N_1596);
and U3997 (N_3997,N_1798,N_152);
nand U3998 (N_3998,N_1552,N_1939);
or U3999 (N_3999,N_10,N_961);
nor U4000 (N_4000,N_3182,N_2782);
or U4001 (N_4001,N_3075,N_2175);
nor U4002 (N_4002,N_2933,N_2253);
nand U4003 (N_4003,N_3045,N_3165);
nand U4004 (N_4004,N_2455,N_3366);
xor U4005 (N_4005,N_2660,N_2234);
and U4006 (N_4006,N_3328,N_3871);
or U4007 (N_4007,N_2796,N_3210);
nor U4008 (N_4008,N_2707,N_2907);
and U4009 (N_4009,N_3826,N_3434);
and U4010 (N_4010,N_2497,N_2541);
or U4011 (N_4011,N_3715,N_3428);
or U4012 (N_4012,N_2565,N_2518);
or U4013 (N_4013,N_3270,N_3954);
nand U4014 (N_4014,N_2107,N_2795);
or U4015 (N_4015,N_3556,N_3734);
nand U4016 (N_4016,N_3299,N_2240);
nor U4017 (N_4017,N_2005,N_2526);
nand U4018 (N_4018,N_3236,N_2028);
and U4019 (N_4019,N_3418,N_3787);
nor U4020 (N_4020,N_2901,N_2978);
or U4021 (N_4021,N_2010,N_3049);
nand U4022 (N_4022,N_2668,N_2197);
nand U4023 (N_4023,N_2679,N_2231);
nor U4024 (N_4024,N_3143,N_3334);
or U4025 (N_4025,N_3613,N_2764);
and U4026 (N_4026,N_3400,N_2603);
nand U4027 (N_4027,N_2325,N_3998);
and U4028 (N_4028,N_2025,N_3385);
nor U4029 (N_4029,N_3872,N_3372);
and U4030 (N_4030,N_3078,N_3470);
nand U4031 (N_4031,N_2693,N_3444);
nand U4032 (N_4032,N_3692,N_3408);
nand U4033 (N_4033,N_3716,N_3948);
and U4034 (N_4034,N_2773,N_3067);
and U4035 (N_4035,N_2881,N_3909);
and U4036 (N_4036,N_3922,N_3336);
and U4037 (N_4037,N_2094,N_3901);
nand U4038 (N_4038,N_2689,N_2636);
or U4039 (N_4039,N_3166,N_2628);
and U4040 (N_4040,N_3647,N_3240);
or U4041 (N_4041,N_3212,N_2586);
and U4042 (N_4042,N_3534,N_3294);
nand U4043 (N_4043,N_2752,N_3395);
or U4044 (N_4044,N_2997,N_3174);
nand U4045 (N_4045,N_3256,N_2295);
and U4046 (N_4046,N_3151,N_2601);
and U4047 (N_4047,N_2629,N_2258);
nor U4048 (N_4048,N_3357,N_2362);
nand U4049 (N_4049,N_3131,N_2973);
or U4050 (N_4050,N_2806,N_3474);
or U4051 (N_4051,N_2033,N_3278);
or U4052 (N_4052,N_3409,N_3015);
and U4053 (N_4053,N_2211,N_3417);
nor U4054 (N_4054,N_2101,N_2132);
or U4055 (N_4055,N_2056,N_3019);
nand U4056 (N_4056,N_3185,N_2963);
nor U4057 (N_4057,N_2675,N_2554);
and U4058 (N_4058,N_3047,N_3358);
nand U4059 (N_4059,N_3897,N_2366);
nand U4060 (N_4060,N_2567,N_2999);
nor U4061 (N_4061,N_2673,N_2616);
nor U4062 (N_4062,N_3624,N_3806);
nand U4063 (N_4063,N_3322,N_2169);
nand U4064 (N_4064,N_3489,N_3359);
or U4065 (N_4065,N_2535,N_3773);
nor U4066 (N_4066,N_2082,N_3644);
nand U4067 (N_4067,N_3247,N_2584);
nand U4068 (N_4068,N_2369,N_3490);
nor U4069 (N_4069,N_2161,N_2407);
nor U4070 (N_4070,N_2392,N_2484);
or U4071 (N_4071,N_3803,N_3241);
nand U4072 (N_4072,N_2867,N_3452);
or U4073 (N_4073,N_3094,N_2371);
and U4074 (N_4074,N_3029,N_3371);
nor U4075 (N_4075,N_3375,N_3632);
and U4076 (N_4076,N_2207,N_2388);
nor U4077 (N_4077,N_3581,N_3096);
nand U4078 (N_4078,N_2179,N_2265);
nand U4079 (N_4079,N_2247,N_3112);
nor U4080 (N_4080,N_2469,N_2364);
or U4081 (N_4081,N_3955,N_2780);
nor U4082 (N_4082,N_3337,N_3656);
or U4083 (N_4083,N_2958,N_2411);
nor U4084 (N_4084,N_2448,N_2530);
xnor U4085 (N_4085,N_3219,N_2694);
nand U4086 (N_4086,N_3022,N_3913);
xor U4087 (N_4087,N_2343,N_3439);
nand U4088 (N_4088,N_2236,N_3223);
nor U4089 (N_4089,N_2092,N_2509);
nand U4090 (N_4090,N_3881,N_2739);
or U4091 (N_4091,N_3972,N_3851);
and U4092 (N_4092,N_2375,N_3422);
nand U4093 (N_4093,N_3124,N_2154);
nand U4094 (N_4094,N_3462,N_3627);
nor U4095 (N_4095,N_3370,N_2548);
or U4096 (N_4096,N_2142,N_2290);
and U4097 (N_4097,N_2964,N_3283);
nor U4098 (N_4098,N_3501,N_2130);
nand U4099 (N_4099,N_3616,N_2012);
nor U4100 (N_4100,N_3480,N_2007);
or U4101 (N_4101,N_2453,N_2182);
or U4102 (N_4102,N_3544,N_3595);
nand U4103 (N_4103,N_3947,N_3840);
xor U4104 (N_4104,N_2318,N_2850);
nand U4105 (N_4105,N_3532,N_3429);
nand U4106 (N_4106,N_3011,N_3658);
and U4107 (N_4107,N_2564,N_3579);
nor U4108 (N_4108,N_2073,N_2023);
xnor U4109 (N_4109,N_3473,N_3583);
nand U4110 (N_4110,N_2767,N_3754);
and U4111 (N_4111,N_3245,N_2651);
or U4112 (N_4112,N_3515,N_2048);
or U4113 (N_4113,N_3708,N_3288);
or U4114 (N_4114,N_2786,N_3760);
or U4115 (N_4115,N_2755,N_2902);
and U4116 (N_4116,N_3073,N_3438);
and U4117 (N_4117,N_2003,N_3214);
nor U4118 (N_4118,N_3817,N_2864);
or U4119 (N_4119,N_3351,N_3244);
or U4120 (N_4120,N_2488,N_3399);
and U4121 (N_4121,N_2176,N_3957);
nor U4122 (N_4122,N_3320,N_3013);
nor U4123 (N_4123,N_2647,N_2361);
xnor U4124 (N_4124,N_3999,N_3394);
nand U4125 (N_4125,N_3483,N_3771);
and U4126 (N_4126,N_3653,N_2861);
nand U4127 (N_4127,N_2426,N_3828);
nand U4128 (N_4128,N_3114,N_3421);
or U4129 (N_4129,N_3309,N_3977);
or U4130 (N_4130,N_3195,N_2572);
xnor U4131 (N_4131,N_3393,N_3929);
xor U4132 (N_4132,N_2662,N_2969);
or U4133 (N_4133,N_3237,N_3028);
nand U4134 (N_4134,N_3102,N_3844);
nor U4135 (N_4135,N_3514,N_3904);
nor U4136 (N_4136,N_2198,N_3589);
nor U4137 (N_4137,N_3722,N_2346);
or U4138 (N_4138,N_2804,N_2674);
or U4139 (N_4139,N_3782,N_3042);
nand U4140 (N_4140,N_3058,N_2127);
nor U4141 (N_4141,N_3946,N_3891);
and U4142 (N_4142,N_3598,N_2740);
nand U4143 (N_4143,N_2008,N_3784);
or U4144 (N_4144,N_3874,N_2529);
nand U4145 (N_4145,N_2264,N_3744);
and U4146 (N_4146,N_2981,N_3920);
nor U4147 (N_4147,N_3976,N_3208);
nand U4148 (N_4148,N_3111,N_2681);
and U4149 (N_4149,N_3146,N_3565);
nor U4150 (N_4150,N_2924,N_3170);
or U4151 (N_4151,N_3362,N_2695);
nand U4152 (N_4152,N_2738,N_2133);
nor U4153 (N_4153,N_2344,N_3985);
and U4154 (N_4154,N_2550,N_3537);
and U4155 (N_4155,N_2878,N_3933);
and U4156 (N_4156,N_3861,N_2514);
nor U4157 (N_4157,N_2756,N_3227);
and U4158 (N_4158,N_3493,N_3367);
nor U4159 (N_4159,N_3883,N_2456);
xnor U4160 (N_4160,N_2291,N_2523);
and U4161 (N_4161,N_2957,N_3035);
nor U4162 (N_4162,N_2229,N_3816);
nor U4163 (N_4163,N_2019,N_2687);
or U4164 (N_4164,N_3477,N_3369);
and U4165 (N_4165,N_3413,N_2128);
and U4166 (N_4166,N_2091,N_2474);
or U4167 (N_4167,N_3390,N_3009);
nand U4168 (N_4168,N_2429,N_2063);
nand U4169 (N_4169,N_3994,N_2285);
and U4170 (N_4170,N_3533,N_2947);
and U4171 (N_4171,N_3794,N_2083);
nor U4172 (N_4172,N_3043,N_2174);
nor U4173 (N_4173,N_3020,N_2734);
or U4174 (N_4174,N_2750,N_3238);
nor U4175 (N_4175,N_3354,N_2663);
nand U4176 (N_4176,N_2613,N_3695);
nand U4177 (N_4177,N_2465,N_2437);
or U4178 (N_4178,N_3125,N_3885);
and U4179 (N_4179,N_3486,N_3295);
nand U4180 (N_4180,N_2097,N_3276);
nand U4181 (N_4181,N_3451,N_2931);
and U4182 (N_4182,N_3785,N_3608);
nand U4183 (N_4183,N_2417,N_2959);
and U4184 (N_4184,N_2753,N_3266);
nand U4185 (N_4185,N_3655,N_3520);
nor U4186 (N_4186,N_3100,N_3242);
nand U4187 (N_4187,N_2862,N_3416);
nor U4188 (N_4188,N_2099,N_3352);
nand U4189 (N_4189,N_2528,N_2288);
nor U4190 (N_4190,N_3916,N_3696);
nand U4191 (N_4191,N_3542,N_2877);
and U4192 (N_4192,N_3681,N_3700);
and U4193 (N_4193,N_2146,N_2200);
nor U4194 (N_4194,N_2577,N_3196);
or U4195 (N_4195,N_2823,N_2042);
nor U4196 (N_4196,N_3932,N_2697);
nor U4197 (N_4197,N_3081,N_3126);
or U4198 (N_4198,N_2057,N_2827);
nor U4199 (N_4199,N_2113,N_3113);
or U4200 (N_4200,N_3942,N_2754);
nor U4201 (N_4201,N_3825,N_3694);
or U4202 (N_4202,N_3732,N_3604);
or U4203 (N_4203,N_2208,N_2071);
nand U4204 (N_4204,N_2269,N_3342);
and U4205 (N_4205,N_2404,N_3997);
nor U4206 (N_4206,N_2106,N_3723);
and U4207 (N_4207,N_3870,N_3169);
nand U4208 (N_4208,N_2451,N_3878);
nor U4209 (N_4209,N_3203,N_3445);
nor U4210 (N_4210,N_2916,N_2140);
nand U4211 (N_4211,N_2201,N_3064);
and U4212 (N_4212,N_3566,N_3471);
nand U4213 (N_4213,N_2031,N_2972);
xor U4214 (N_4214,N_2490,N_2139);
nand U4215 (N_4215,N_3088,N_3181);
nand U4216 (N_4216,N_3882,N_3391);
and U4217 (N_4217,N_3667,N_2081);
nor U4218 (N_4218,N_3800,N_3202);
nand U4219 (N_4219,N_2301,N_3683);
and U4220 (N_4220,N_3802,N_3024);
and U4221 (N_4221,N_3341,N_3211);
and U4222 (N_4222,N_2164,N_2922);
nand U4223 (N_4223,N_2173,N_3699);
xor U4224 (N_4224,N_3160,N_2566);
or U4225 (N_4225,N_2499,N_3951);
nor U4226 (N_4226,N_2270,N_2946);
nand U4227 (N_4227,N_2180,N_3569);
or U4228 (N_4228,N_2832,N_2618);
or U4229 (N_4229,N_3318,N_2875);
nor U4230 (N_4230,N_2563,N_3750);
nand U4231 (N_4231,N_2966,N_2148);
or U4232 (N_4232,N_2519,N_2661);
nand U4233 (N_4233,N_2108,N_3652);
and U4234 (N_4234,N_2225,N_2928);
nor U4235 (N_4235,N_3980,N_3496);
and U4236 (N_4236,N_3292,N_2276);
nor U4237 (N_4237,N_2701,N_3426);
xnor U4238 (N_4238,N_2228,N_3260);
and U4239 (N_4239,N_2249,N_3264);
nand U4240 (N_4240,N_2976,N_2955);
nor U4241 (N_4241,N_2272,N_3105);
nor U4242 (N_4242,N_2266,N_2400);
nor U4243 (N_4243,N_3739,N_3475);
or U4244 (N_4244,N_3665,N_3122);
and U4245 (N_4245,N_2461,N_2432);
nor U4246 (N_4246,N_3407,N_3827);
nor U4247 (N_4247,N_3258,N_3780);
or U4248 (N_4248,N_3691,N_2310);
nor U4249 (N_4249,N_3635,N_3025);
or U4250 (N_4250,N_3988,N_2084);
or U4251 (N_4251,N_2079,N_2599);
or U4252 (N_4252,N_2781,N_2398);
xnor U4253 (N_4253,N_3865,N_3823);
nand U4254 (N_4254,N_2116,N_3476);
and U4255 (N_4255,N_3465,N_3335);
and U4256 (N_4256,N_3841,N_2095);
and U4257 (N_4257,N_3459,N_3662);
and U4258 (N_4258,N_3559,N_2252);
nand U4259 (N_4259,N_3919,N_2579);
or U4260 (N_4260,N_2510,N_3085);
nor U4261 (N_4261,N_2335,N_2606);
and U4262 (N_4262,N_2306,N_2365);
or U4263 (N_4263,N_3497,N_3279);
and U4264 (N_4264,N_3846,N_3661);
or U4265 (N_4265,N_2965,N_2984);
or U4266 (N_4266,N_3619,N_2975);
and U4267 (N_4267,N_2297,N_3996);
and U4268 (N_4268,N_3360,N_3066);
nand U4269 (N_4269,N_3140,N_3233);
and U4270 (N_4270,N_2076,N_3839);
or U4271 (N_4271,N_3848,N_2822);
nand U4272 (N_4272,N_3059,N_2941);
and U4273 (N_4273,N_3729,N_2570);
and U4274 (N_4274,N_3941,N_3324);
nand U4275 (N_4275,N_3228,N_3973);
nor U4276 (N_4276,N_2477,N_2517);
and U4277 (N_4277,N_3461,N_3083);
or U4278 (N_4278,N_2480,N_2552);
and U4279 (N_4279,N_2527,N_3858);
nor U4280 (N_4280,N_3164,N_2585);
nand U4281 (N_4281,N_2214,N_2038);
and U4282 (N_4282,N_2016,N_2467);
and U4283 (N_4283,N_3755,N_2657);
nand U4284 (N_4284,N_3873,N_3134);
and U4285 (N_4285,N_2558,N_2360);
nor U4286 (N_4286,N_3859,N_2814);
and U4287 (N_4287,N_2302,N_3725);
or U4288 (N_4288,N_2708,N_3044);
and U4289 (N_4289,N_3198,N_3697);
nand U4290 (N_4290,N_2985,N_2103);
or U4291 (N_4291,N_2612,N_3669);
and U4292 (N_4292,N_2553,N_2784);
or U4293 (N_4293,N_2655,N_2724);
xnor U4294 (N_4294,N_3611,N_3648);
or U4295 (N_4295,N_3961,N_2713);
nor U4296 (N_4296,N_3205,N_2876);
and U4297 (N_4297,N_2122,N_2086);
xor U4298 (N_4298,N_3610,N_3055);
and U4299 (N_4299,N_3726,N_3824);
nor U4300 (N_4300,N_2900,N_2135);
nand U4301 (N_4301,N_3504,N_2706);
nand U4302 (N_4302,N_3835,N_2515);
or U4303 (N_4303,N_2096,N_3731);
nor U4304 (N_4304,N_2858,N_3117);
and U4305 (N_4305,N_3641,N_2696);
or U4306 (N_4306,N_3646,N_2645);
or U4307 (N_4307,N_2995,N_2102);
xnor U4308 (N_4308,N_2654,N_3261);
and U4309 (N_4309,N_3629,N_3289);
or U4310 (N_4310,N_2359,N_2328);
nand U4311 (N_4311,N_2222,N_2615);
nand U4312 (N_4312,N_2195,N_2233);
and U4313 (N_4313,N_3511,N_3796);
xor U4314 (N_4314,N_2934,N_3150);
nand U4315 (N_4315,N_3030,N_2383);
xor U4316 (N_4316,N_3617,N_2380);
and U4317 (N_4317,N_2298,N_2637);
and U4318 (N_4318,N_2431,N_3424);
or U4319 (N_4319,N_3061,N_2703);
nor U4320 (N_4320,N_2436,N_3041);
or U4321 (N_4321,N_3072,N_2605);
and U4322 (N_4322,N_3781,N_3547);
and U4323 (N_4323,N_2652,N_2891);
and U4324 (N_4324,N_2089,N_2368);
nor U4325 (N_4325,N_2304,N_2742);
nand U4326 (N_4326,N_3222,N_2341);
and U4327 (N_4327,N_2275,N_3312);
nor U4328 (N_4328,N_3381,N_2866);
nor U4329 (N_4329,N_2575,N_3555);
nor U4330 (N_4330,N_2791,N_2960);
nand U4331 (N_4331,N_3963,N_2882);
or U4332 (N_4332,N_3855,N_2165);
nand U4333 (N_4333,N_2838,N_2243);
nand U4334 (N_4334,N_2351,N_2982);
nor U4335 (N_4335,N_2593,N_2373);
and U4336 (N_4336,N_3597,N_3050);
xor U4337 (N_4337,N_3206,N_2935);
and U4338 (N_4338,N_3778,N_3079);
nor U4339 (N_4339,N_2017,N_2774);
and U4340 (N_4340,N_3163,N_2716);
and U4341 (N_4341,N_2143,N_3675);
or U4342 (N_4342,N_2379,N_3580);
nand U4343 (N_4343,N_2493,N_3770);
and U4344 (N_4344,N_3344,N_3767);
and U4345 (N_4345,N_2549,N_3423);
xor U4346 (N_4346,N_3801,N_3609);
nor U4347 (N_4347,N_3343,N_3678);
nand U4348 (N_4348,N_3054,N_2705);
or U4349 (N_4349,N_3271,N_3006);
or U4350 (N_4350,N_2539,N_2559);
nor U4351 (N_4351,N_2337,N_3593);
nand U4352 (N_4352,N_3090,N_2908);
and U4353 (N_4353,N_2513,N_3194);
and U4354 (N_4354,N_3690,N_3888);
nor U4355 (N_4355,N_2452,N_2930);
xnor U4356 (N_4356,N_3526,N_3502);
and U4357 (N_4357,N_3435,N_2619);
or U4358 (N_4358,N_3698,N_3805);
and U4359 (N_4359,N_2691,N_3162);
and U4360 (N_4360,N_3201,N_3121);
nor U4361 (N_4361,N_2410,N_2415);
nor U4362 (N_4362,N_2378,N_2803);
nor U4363 (N_4363,N_2193,N_2171);
nand U4364 (N_4364,N_3226,N_3590);
or U4365 (N_4365,N_2659,N_3192);
nor U4366 (N_4366,N_2909,N_2594);
nor U4367 (N_4367,N_2798,N_2066);
and U4368 (N_4368,N_2376,N_3176);
or U4369 (N_4369,N_2851,N_2951);
nor U4370 (N_4370,N_3880,N_2896);
nor U4371 (N_4371,N_3106,N_3255);
nand U4372 (N_4372,N_3101,N_2873);
and U4373 (N_4373,N_2303,N_2669);
nor U4374 (N_4374,N_3177,N_2797);
nor U4375 (N_4375,N_2709,N_3524);
nor U4376 (N_4376,N_3152,N_3230);
or U4377 (N_4377,N_2671,N_2970);
nor U4378 (N_4378,N_3852,N_3495);
nand U4379 (N_4379,N_2075,N_3097);
and U4380 (N_4380,N_3587,N_3602);
and U4381 (N_4381,N_2993,N_3376);
nand U4382 (N_4382,N_3735,N_3257);
or U4383 (N_4383,N_2151,N_3832);
nand U4384 (N_4384,N_2444,N_3906);
nor U4385 (N_4385,N_2641,N_2137);
nor U4386 (N_4386,N_2206,N_2672);
xnor U4387 (N_4387,N_2185,N_3759);
or U4388 (N_4388,N_3348,N_2634);
nor U4389 (N_4389,N_2869,N_2653);
nand U4390 (N_4390,N_2865,N_3762);
or U4391 (N_4391,N_3745,N_2109);
nand U4392 (N_4392,N_3068,N_3115);
or U4393 (N_4393,N_2492,N_3625);
nand U4394 (N_4394,N_2807,N_2255);
nor U4395 (N_4395,N_2913,N_3069);
or U4396 (N_4396,N_2961,N_2611);
nand U4397 (N_4397,N_3269,N_3962);
nand U4398 (N_4398,N_3720,N_2824);
nor U4399 (N_4399,N_3968,N_2494);
nor U4400 (N_4400,N_2329,N_2943);
nand U4401 (N_4401,N_3217,N_3943);
xnor U4402 (N_4402,N_3758,N_3728);
or U4403 (N_4403,N_3631,N_3172);
nand U4404 (N_4404,N_2733,N_3017);
xnor U4405 (N_4405,N_2203,N_3310);
and U4406 (N_4406,N_3186,N_3837);
or U4407 (N_4407,N_2544,N_2846);
and U4408 (N_4408,N_2481,N_3159);
nor U4409 (N_4409,N_2726,N_3792);
and U4410 (N_4410,N_2598,N_3554);
and U4411 (N_4411,N_3949,N_2333);
or U4412 (N_4412,N_3250,N_2863);
nor U4413 (N_4413,N_3747,N_3535);
or U4414 (N_4414,N_2087,N_3761);
nand U4415 (N_4415,N_2962,N_2036);
or U4416 (N_4416,N_2906,N_2817);
or U4417 (N_4417,N_3937,N_2188);
or U4418 (N_4418,N_3464,N_3905);
and U4419 (N_4419,N_2785,N_3636);
or U4420 (N_4420,N_3512,N_3670);
nand U4421 (N_4421,N_2792,N_2254);
and U4422 (N_4422,N_2639,N_2447);
and U4423 (N_4423,N_3879,N_2013);
nand U4424 (N_4424,N_2473,N_3812);
and U4425 (N_4425,N_2423,N_2910);
and U4426 (N_4426,N_2980,N_3207);
or U4427 (N_4427,N_3516,N_3903);
or U4428 (N_4428,N_3651,N_3065);
nor U4429 (N_4429,N_2261,N_2021);
xnor U4430 (N_4430,N_2177,N_2915);
nand U4431 (N_4431,N_2058,N_3529);
and U4432 (N_4432,N_2646,N_2090);
nor U4433 (N_4433,N_3300,N_3314);
nand U4434 (N_4434,N_3703,N_2720);
and U4435 (N_4435,N_3315,N_2401);
nand U4436 (N_4436,N_3831,N_2434);
and U4437 (N_4437,N_2986,N_3912);
and U4438 (N_4438,N_3743,N_3330);
or U4439 (N_4439,N_2219,N_3282);
or U4440 (N_4440,N_3265,N_3016);
nand U4441 (N_4441,N_3711,N_2583);
or U4442 (N_4442,N_2402,N_3221);
nand U4443 (N_4443,N_3586,N_2608);
nor U4444 (N_4444,N_3676,N_2888);
nor U4445 (N_4445,N_2027,N_3021);
or U4446 (N_4446,N_3506,N_3564);
and U4447 (N_4447,N_3702,N_3014);
nand U4448 (N_4448,N_2443,N_3436);
nor U4449 (N_4449,N_2617,N_3389);
and U4450 (N_4450,N_3612,N_3074);
nand U4451 (N_4451,N_2289,N_2610);
and U4452 (N_4452,N_3740,N_2293);
nor U4453 (N_4453,N_3239,N_3517);
or U4454 (N_4454,N_2745,N_2316);
and U4455 (N_4455,N_3965,N_3978);
and U4456 (N_4456,N_2018,N_2370);
nor U4457 (N_4457,N_3974,N_2884);
nand U4458 (N_4458,N_3129,N_3910);
nand U4459 (N_4459,N_3430,N_2837);
xnor U4460 (N_4460,N_2039,N_3523);
or U4461 (N_4461,N_2592,N_2748);
or U4462 (N_4462,N_3967,N_2658);
xnor U4463 (N_4463,N_2438,N_3373);
nor U4464 (N_4464,N_3406,N_2897);
or U4465 (N_4465,N_2799,N_3432);
and U4466 (N_4466,N_2256,N_3650);
or U4467 (N_4467,N_3287,N_3446);
or U4468 (N_4468,N_3374,N_3705);
nand U4469 (N_4469,N_2595,N_2352);
nor U4470 (N_4470,N_3304,N_2723);
nor U4471 (N_4471,N_3147,N_2347);
and U4472 (N_4472,N_3688,N_3981);
and U4473 (N_4473,N_2698,N_2296);
nand U4474 (N_4474,N_2131,N_3663);
and U4475 (N_4475,N_2309,N_3145);
and U4476 (N_4476,N_2852,N_2805);
nor U4477 (N_4477,N_2987,N_2160);
nand U4478 (N_4478,N_3290,N_3706);
or U4479 (N_4479,N_2842,N_3543);
nand U4480 (N_4480,N_3442,N_3737);
nand U4481 (N_4481,N_3660,N_3232);
nor U4482 (N_4482,N_2011,N_3457);
or U4483 (N_4483,N_3254,N_2377);
nor U4484 (N_4484,N_3037,N_2495);
and U4485 (N_4485,N_2470,N_3628);
nand U4486 (N_4486,N_2126,N_3763);
or U4487 (N_4487,N_3293,N_3479);
and U4488 (N_4488,N_2118,N_3911);
or U4489 (N_4489,N_2573,N_3349);
and U4490 (N_4490,N_2825,N_3630);
or U4491 (N_4491,N_3482,N_3599);
nor U4492 (N_4492,N_2855,N_3926);
xnor U4493 (N_4493,N_2883,N_3591);
and U4494 (N_4494,N_2677,N_3275);
nand U4495 (N_4495,N_2656,N_2504);
nand U4496 (N_4496,N_3229,N_2604);
nand U4497 (N_4497,N_2524,N_2561);
or U4498 (N_4498,N_3645,N_2421);
nand U4499 (N_4499,N_2170,N_3766);
nor U4500 (N_4500,N_3838,N_3607);
or U4501 (N_4501,N_2845,N_2684);
nand U4502 (N_4502,N_3989,N_3005);
and U4503 (N_4503,N_3057,N_2808);
or U4504 (N_4504,N_3189,N_2257);
and U4505 (N_4505,N_3798,N_3829);
or U4506 (N_4506,N_3321,N_3808);
nand U4507 (N_4507,N_3756,N_3118);
nor U4508 (N_4508,N_2562,N_2543);
or U4509 (N_4509,N_3188,N_2224);
nor U4510 (N_4510,N_2050,N_2667);
nand U4511 (N_4511,N_2516,N_2839);
and U4512 (N_4512,N_3538,N_3353);
nor U4513 (N_4513,N_2396,N_3052);
nand U4514 (N_4514,N_2609,N_2152);
nand U4515 (N_4515,N_3605,N_3709);
nor U4516 (N_4516,N_2600,N_3107);
nand U4517 (N_4517,N_2110,N_3783);
and U4518 (N_4518,N_2542,N_2196);
nand U4519 (N_4519,N_3235,N_2299);
and U4520 (N_4520,N_2070,N_3272);
nand U4521 (N_4521,N_3876,N_3984);
or U4522 (N_4522,N_3959,N_2189);
and U4523 (N_4523,N_3087,N_2123);
and U4524 (N_4524,N_3887,N_2427);
nand U4525 (N_4525,N_3795,N_2487);
and U4526 (N_4526,N_3769,N_2194);
or U4527 (N_4527,N_2537,N_3730);
and U4528 (N_4528,N_3777,N_3718);
nor U4529 (N_4529,N_3899,N_3398);
nand U4530 (N_4530,N_3940,N_2267);
nor U4531 (N_4531,N_2047,N_3527);
and U4532 (N_4532,N_2489,N_3086);
nor U4533 (N_4533,N_2046,N_2853);
nor U4534 (N_4534,N_2326,N_3713);
nor U4535 (N_4535,N_3945,N_3133);
nand U4536 (N_4536,N_3031,N_2769);
nor U4537 (N_4537,N_3500,N_3053);
and U4538 (N_4538,N_3281,N_2271);
or U4539 (N_4539,N_3018,N_3187);
xor U4540 (N_4540,N_3522,N_3116);
nand U4541 (N_4541,N_3886,N_2239);
or U4542 (N_4542,N_2744,N_2835);
nor U4543 (N_4543,N_2953,N_2202);
xor U4544 (N_4544,N_3727,N_2787);
or U4545 (N_4545,N_2037,N_3637);
or U4546 (N_4546,N_3986,N_2760);
and U4547 (N_4547,N_2190,N_2068);
nand U4548 (N_4548,N_2942,N_3956);
nand U4549 (N_4549,N_3869,N_3403);
nor U4550 (N_4550,N_3818,N_3809);
or U4551 (N_4551,N_3302,N_2433);
or U4552 (N_4552,N_2279,N_2121);
nor U4553 (N_4553,N_3062,N_3026);
nor U4554 (N_4554,N_3384,N_2308);
nor U4555 (N_4555,N_2642,N_3157);
nor U4556 (N_4556,N_3466,N_3259);
nand U4557 (N_4557,N_2717,N_2728);
nor U4558 (N_4558,N_3833,N_2349);
nor U4559 (N_4559,N_2625,N_3204);
or U4560 (N_4560,N_3285,N_3907);
or U4561 (N_4561,N_2967,N_2576);
nor U4562 (N_4562,N_3900,N_2676);
or U4563 (N_4563,N_3173,N_3076);
nand U4564 (N_4564,N_3386,N_2692);
or U4565 (N_4565,N_2849,N_3267);
and U4566 (N_4566,N_2428,N_2664);
or U4567 (N_4567,N_2630,N_3993);
nand U4568 (N_4568,N_2040,N_3674);
nand U4569 (N_4569,N_2927,N_2623);
or U4570 (N_4570,N_3966,N_3333);
and U4571 (N_4571,N_3051,N_2859);
nor U4572 (N_4572,N_3148,N_2330);
and U4573 (N_4573,N_3253,N_2334);
xnor U4574 (N_4574,N_2551,N_3070);
and U4575 (N_4575,N_3578,N_2080);
and U4576 (N_4576,N_2751,N_3797);
or U4577 (N_4577,N_2885,N_2105);
nor U4578 (N_4578,N_3775,N_3953);
or U4579 (N_4579,N_3584,N_2227);
or U4580 (N_4580,N_3274,N_2950);
nand U4581 (N_4581,N_2812,N_2460);
or U4582 (N_4582,N_3412,N_2472);
or U4583 (N_4583,N_3622,N_3930);
and U4584 (N_4584,N_2077,N_3487);
and U4585 (N_4585,N_2442,N_3135);
nor U4586 (N_4586,N_2034,N_3200);
and U4587 (N_4587,N_2363,N_2125);
nor U4588 (N_4588,N_3469,N_3558);
and U4589 (N_4589,N_3693,N_3092);
or U4590 (N_4590,N_2336,N_3724);
nor U4591 (N_4591,N_3472,N_2938);
and U4592 (N_4592,N_3819,N_3546);
and U4593 (N_4593,N_2793,N_3918);
nor U4594 (N_4594,N_2119,N_3215);
nor U4595 (N_4595,N_3640,N_3184);
nor U4596 (N_4596,N_2940,N_3915);
or U4597 (N_4597,N_2145,N_2893);
or U4598 (N_4598,N_2992,N_2422);
nor U4599 (N_4599,N_2060,N_2844);
xor U4600 (N_4600,N_2991,N_3449);
and U4601 (N_4601,N_2115,N_2918);
nor U4602 (N_4602,N_2525,N_3350);
and U4603 (N_4603,N_2763,N_3103);
or U4604 (N_4604,N_3329,N_3468);
or U4605 (N_4605,N_2929,N_2059);
nor U4606 (N_4606,N_2589,N_3082);
nand U4607 (N_4607,N_3071,N_3856);
and U4608 (N_4608,N_3036,N_3528);
nand U4609 (N_4609,N_2425,N_3220);
nor U4610 (N_4610,N_3218,N_2638);
nand U4611 (N_4611,N_2098,N_3594);
nand U4612 (N_4612,N_3541,N_3643);
nor U4613 (N_4613,N_3091,N_3668);
nor U4614 (N_4614,N_2714,N_3491);
nand U4615 (N_4615,N_2749,N_3199);
and U4616 (N_4616,N_3751,N_3454);
nor U4617 (N_4617,N_2282,N_2802);
and U4618 (N_4618,N_2284,N_2331);
or U4619 (N_4619,N_3519,N_2905);
or U4620 (N_4620,N_2345,N_3392);
or U4621 (N_4621,N_3789,N_3815);
and U4622 (N_4622,N_3317,N_2468);
or U4623 (N_4623,N_2320,N_2324);
nor U4624 (N_4624,N_2830,N_2014);
and U4625 (N_4625,N_3327,N_2847);
nor U4626 (N_4626,N_3167,N_3243);
nor U4627 (N_4627,N_3753,N_3786);
or U4628 (N_4628,N_3216,N_3156);
nor U4629 (N_4629,N_3925,N_2685);
or U4630 (N_4630,N_3405,N_3938);
or U4631 (N_4631,N_2372,N_3620);
xor U4632 (N_4632,N_2209,N_2508);
or U4633 (N_4633,N_3427,N_3460);
or U4634 (N_4634,N_3433,N_3982);
nand U4635 (N_4635,N_2024,N_2536);
or U4636 (N_4636,N_3563,N_3896);
nand U4637 (N_4637,N_2828,N_2732);
or U4638 (N_4638,N_3023,N_3849);
nand U4639 (N_4639,N_3862,N_3450);
nand U4640 (N_4640,N_2217,N_2277);
or U4641 (N_4641,N_3550,N_2800);
nand U4642 (N_4642,N_3056,N_3765);
or U4643 (N_4643,N_2597,N_2722);
nand U4644 (N_4644,N_3225,N_2578);
and U4645 (N_4645,N_2104,N_2533);
and U4646 (N_4646,N_2220,N_3027);
or U4647 (N_4647,N_3251,N_3388);
and U4648 (N_4648,N_3736,N_3467);
and U4649 (N_4649,N_3788,N_2571);
or U4650 (N_4650,N_2307,N_2020);
and U4651 (N_4651,N_2053,N_3346);
or U4652 (N_4652,N_3099,N_2887);
nor U4653 (N_4653,N_2030,N_2816);
or U4654 (N_4654,N_2412,N_2503);
nand U4655 (N_4655,N_2829,N_3415);
nand U4656 (N_4656,N_3821,N_3377);
and U4657 (N_4657,N_3448,N_3813);
or U4658 (N_4658,N_2890,N_2914);
nand U4659 (N_4659,N_2479,N_3132);
or U4660 (N_4660,N_2466,N_3084);
and U4661 (N_4661,N_2582,N_2983);
or U4662 (N_4662,N_3682,N_3742);
or U4663 (N_4663,N_3168,N_3000);
nand U4664 (N_4664,N_2172,N_3864);
or U4665 (N_4665,N_3685,N_3884);
or U4666 (N_4666,N_3822,N_3714);
nand U4667 (N_4667,N_2191,N_2644);
nand U4668 (N_4668,N_3562,N_2731);
and U4669 (N_4669,N_3380,N_3684);
nand U4670 (N_4670,N_2052,N_2840);
or U4671 (N_4671,N_3790,N_2163);
and U4672 (N_4672,N_2759,N_2280);
or U4673 (N_4673,N_3191,N_3860);
or U4674 (N_4674,N_3895,N_2144);
nor U4675 (N_4675,N_2649,N_2044);
or U4676 (N_4676,N_2766,N_2178);
or U4677 (N_4677,N_3179,N_2424);
nor U4678 (N_4678,N_2274,N_2218);
and U4679 (N_4679,N_2587,N_2556);
and U4680 (N_4680,N_3575,N_3440);
and U4681 (N_4681,N_2602,N_2245);
or U4682 (N_4682,N_2153,N_3799);
nand U4683 (N_4683,N_2356,N_2199);
and U4684 (N_4684,N_3811,N_3306);
and U4685 (N_4685,N_2311,N_2314);
and U4686 (N_4686,N_2226,N_3093);
nand U4687 (N_4687,N_3582,N_2416);
or U4688 (N_4688,N_3379,N_3396);
and U4689 (N_4689,N_3231,N_2879);
nor U4690 (N_4690,N_3262,N_2819);
nor U4691 (N_4691,N_2439,N_2062);
or U4692 (N_4692,N_2156,N_3772);
and U4693 (N_4693,N_3443,N_2166);
or U4694 (N_4694,N_3549,N_3987);
nor U4695 (N_4695,N_3513,N_2880);
nor U4696 (N_4696,N_2626,N_3128);
and U4697 (N_4697,N_3877,N_2482);
nor U4698 (N_4698,N_2971,N_2278);
or U4699 (N_4699,N_3224,N_2735);
nand U4700 (N_4700,N_2281,N_3268);
and U4701 (N_4701,N_3991,N_3137);
nor U4702 (N_4702,N_2332,N_3530);
or U4703 (N_4703,N_2323,N_2357);
nor U4704 (N_4704,N_3046,N_3332);
and U4705 (N_4705,N_2511,N_3975);
or U4706 (N_4706,N_3387,N_2353);
or U4707 (N_4707,N_2159,N_3291);
or U4708 (N_4708,N_2768,N_3606);
or U4709 (N_4709,N_2032,N_3577);
nor U4710 (N_4710,N_2064,N_3331);
or U4711 (N_4711,N_2783,N_3508);
nor U4712 (N_4712,N_2454,N_3752);
nor U4713 (N_4713,N_2815,N_2393);
nor U4714 (N_4714,N_2794,N_2287);
nor U4715 (N_4715,N_3356,N_2996);
nand U4716 (N_4716,N_2496,N_3992);
and U4717 (N_4717,N_3567,N_2831);
xnor U4718 (N_4718,N_2540,N_2730);
nand U4719 (N_4719,N_3531,N_3894);
nor U4720 (N_4720,N_2167,N_3175);
or U4721 (N_4721,N_2384,N_3935);
or U4722 (N_4722,N_2546,N_2157);
nor U4723 (N_4723,N_3867,N_2093);
nand U4724 (N_4724,N_2015,N_3130);
nand U4725 (N_4725,N_2936,N_2462);
nor U4726 (N_4726,N_2486,N_3814);
xor U4727 (N_4727,N_3425,N_3923);
nor U4728 (N_4728,N_2666,N_2242);
and U4729 (N_4729,N_2522,N_3420);
nor U4730 (N_4730,N_2358,N_2391);
nor U4731 (N_4731,N_2367,N_2757);
or U4732 (N_4732,N_3048,N_2665);
or U4733 (N_4733,N_3401,N_3010);
nor U4734 (N_4734,N_3364,N_2312);
and U4735 (N_4735,N_3654,N_3507);
nand U4736 (N_4736,N_3931,N_2843);
and U4737 (N_4737,N_3863,N_3666);
xor U4738 (N_4738,N_2322,N_2181);
and U4739 (N_4739,N_2051,N_2230);
nand U4740 (N_4740,N_2259,N_2834);
or U4741 (N_4741,N_2342,N_3089);
nor U4742 (N_4742,N_2237,N_2710);
nand U4743 (N_4743,N_3893,N_3095);
nor U4744 (N_4744,N_2483,N_3853);
or U4745 (N_4745,N_2871,N_3190);
nor U4746 (N_4746,N_2263,N_2811);
nand U4747 (N_4747,N_2860,N_2262);
or U4748 (N_4748,N_3626,N_3303);
nor U4749 (N_4749,N_2979,N_3286);
and U4750 (N_4750,N_2778,N_2678);
nor U4751 (N_4751,N_2643,N_3453);
or U4752 (N_4752,N_3834,N_2990);
or U4753 (N_4753,N_3924,N_2988);
and U4754 (N_4754,N_2009,N_2450);
and U4755 (N_4755,N_3921,N_2925);
nor U4756 (N_4756,N_3437,N_2445);
nand U4757 (N_4757,N_3615,N_2989);
nand U4758 (N_4758,N_3488,N_3701);
and U4759 (N_4759,N_2574,N_2374);
nor U4760 (N_4760,N_3677,N_3969);
or U4761 (N_4761,N_3639,N_3952);
or U4762 (N_4762,N_2397,N_2250);
and U4763 (N_4763,N_3307,N_3764);
and U4764 (N_4764,N_3779,N_3008);
xor U4765 (N_4765,N_2413,N_2868);
nand U4766 (N_4766,N_3741,N_2463);
nand U4767 (N_4767,N_2607,N_2779);
nand U4768 (N_4768,N_3733,N_3458);
and U4769 (N_4769,N_3447,N_2117);
or U4770 (N_4770,N_2841,N_2491);
or U4771 (N_4771,N_2903,N_3518);
and U4772 (N_4772,N_3119,N_2313);
or U4773 (N_4773,N_2471,N_3308);
and U4774 (N_4774,N_2507,N_2789);
nor U4775 (N_4775,N_3402,N_3875);
and U4776 (N_4776,N_2761,N_2022);
nor U4777 (N_4777,N_2029,N_2718);
nand U4778 (N_4778,N_2520,N_2836);
and U4779 (N_4779,N_2478,N_3180);
nor U4780 (N_4780,N_2205,N_2633);
and U4781 (N_4781,N_2632,N_3481);
nand U4782 (N_4782,N_3990,N_2149);
and U4783 (N_4783,N_3478,N_2441);
and U4784 (N_4784,N_2580,N_3503);
and U4785 (N_4785,N_2591,N_2339);
nand U4786 (N_4786,N_3738,N_3123);
nand U4787 (N_4787,N_2770,N_2919);
xor U4788 (N_4788,N_2818,N_2485);
or U4789 (N_4789,N_2821,N_3964);
nor U4790 (N_4790,N_3441,N_3548);
and U4791 (N_4791,N_2952,N_3007);
nor U4792 (N_4792,N_2640,N_2801);
nor U4793 (N_4793,N_2305,N_3614);
xnor U4794 (N_4794,N_2788,N_3463);
nor U4795 (N_4795,N_3355,N_2506);
or U4796 (N_4796,N_2385,N_2420);
nand U4797 (N_4797,N_3305,N_2215);
or U4798 (N_4798,N_2894,N_2624);
and U4799 (N_4799,N_2810,N_2596);
and U4800 (N_4800,N_3934,N_2414);
nor U4801 (N_4801,N_2035,N_3914);
nand U4802 (N_4802,N_3039,N_2409);
and U4803 (N_4803,N_3557,N_2238);
or U4804 (N_4804,N_2746,N_3158);
nand U4805 (N_4805,N_2390,N_3033);
xnor U4806 (N_4806,N_3712,N_3136);
nor U4807 (N_4807,N_3034,N_3618);
nor U4808 (N_4808,N_3361,N_3363);
and U4809 (N_4809,N_2260,N_2045);
or U4810 (N_4810,N_2502,N_3551);
and U4811 (N_4811,N_2419,N_2283);
nand U4812 (N_4812,N_2622,N_2809);
nor U4813 (N_4813,N_2614,N_2244);
or U4814 (N_4814,N_3277,N_3671);
nor U4815 (N_4815,N_2688,N_2631);
and U4816 (N_4816,N_3971,N_3983);
and U4817 (N_4817,N_2389,N_3323);
nand U4818 (N_4818,N_2568,N_3012);
or U4819 (N_4819,N_3845,N_3521);
nor U4820 (N_4820,N_3525,N_2512);
and U4821 (N_4821,N_2061,N_3704);
nor U4822 (N_4822,N_2968,N_2771);
and U4823 (N_4823,N_2926,N_2292);
nor U4824 (N_4824,N_3144,N_2235);
and U4825 (N_4825,N_2854,N_3142);
and U4826 (N_4826,N_2870,N_2700);
and U4827 (N_4827,N_2394,N_3536);
xor U4828 (N_4828,N_3746,N_3153);
or U4829 (N_4829,N_2069,N_2403);
and U4830 (N_4830,N_2327,N_2974);
nand U4831 (N_4831,N_3485,N_2475);
nor U4832 (N_4832,N_3183,N_3063);
nand U4833 (N_4833,N_2026,N_3455);
and U4834 (N_4834,N_3032,N_3576);
or U4835 (N_4835,N_3368,N_2680);
nor U4836 (N_4836,N_2945,N_3154);
nor U4837 (N_4837,N_2775,N_2300);
nor U4838 (N_4838,N_2204,N_2790);
xnor U4839 (N_4839,N_3890,N_3248);
nor U4840 (N_4840,N_3719,N_2405);
nor U4841 (N_4841,N_3807,N_2534);
nor U4842 (N_4842,N_2686,N_2319);
nand U4843 (N_4843,N_3621,N_2124);
nand U4844 (N_4844,N_2538,N_2772);
or U4845 (N_4845,N_2350,N_3296);
or U4846 (N_4846,N_2702,N_2168);
and U4847 (N_4847,N_3995,N_3679);
nand U4848 (N_4848,N_3338,N_3298);
nor U4849 (N_4849,N_2054,N_2911);
nor U4850 (N_4850,N_2355,N_3252);
nor U4851 (N_4851,N_2682,N_3494);
nand U4852 (N_4852,N_3171,N_3979);
or U4853 (N_4853,N_2588,N_3553);
and U4854 (N_4854,N_2857,N_3098);
nand U4855 (N_4855,N_3687,N_3139);
xor U4856 (N_4856,N_3545,N_2338);
or U4857 (N_4857,N_2547,N_3672);
and U4858 (N_4858,N_2719,N_2777);
or U4859 (N_4859,N_3768,N_2650);
and U4860 (N_4860,N_3484,N_2590);
or U4861 (N_4861,N_3657,N_3209);
nand U4862 (N_4862,N_3970,N_2221);
nor U4863 (N_4863,N_3060,N_2848);
xnor U4864 (N_4864,N_3585,N_3378);
nand U4865 (N_4865,N_3950,N_3311);
and U4866 (N_4866,N_3498,N_2136);
nor U4867 (N_4867,N_2112,N_2889);
or U4868 (N_4868,N_3109,N_3002);
nor U4869 (N_4869,N_2886,N_3004);
nor U4870 (N_4870,N_2670,N_3908);
nor U4871 (N_4871,N_3540,N_2956);
nor U4872 (N_4872,N_2435,N_3138);
nor U4873 (N_4873,N_2904,N_3492);
and U4874 (N_4874,N_2387,N_2004);
nor U4875 (N_4875,N_3326,N_3120);
and U4876 (N_4876,N_3411,N_3280);
and U4877 (N_4877,N_3689,N_2949);
nand U4878 (N_4878,N_2476,N_2505);
or U4879 (N_4879,N_2743,N_2162);
nor U4880 (N_4880,N_3804,N_3301);
or U4881 (N_4881,N_2043,N_2000);
and U4882 (N_4882,N_3710,N_2317);
nand U4883 (N_4883,N_3561,N_2418);
or U4884 (N_4884,N_2241,N_2895);
and U4885 (N_4885,N_2704,N_3038);
nor U4886 (N_4886,N_2621,N_2994);
nand U4887 (N_4887,N_3898,N_2348);
nand U4888 (N_4888,N_2557,N_3820);
and U4889 (N_4889,N_2440,N_3917);
nand U4890 (N_4890,N_2937,N_3776);
and U4891 (N_4891,N_3003,N_3836);
nor U4892 (N_4892,N_2727,N_3213);
and U4893 (N_4893,N_2758,N_2998);
and U4894 (N_4894,N_3847,N_3414);
and U4895 (N_4895,N_3596,N_3552);
and U4896 (N_4896,N_2813,N_2381);
nor U4897 (N_4897,N_2041,N_2856);
nand U4898 (N_4898,N_3659,N_2273);
xor U4899 (N_4899,N_3600,N_3892);
or U4900 (N_4900,N_2049,N_3560);
or U4901 (N_4901,N_3345,N_2158);
nor U4902 (N_4902,N_3431,N_2899);
nand U4903 (N_4903,N_2100,N_3686);
nor U4904 (N_4904,N_3623,N_2315);
or U4905 (N_4905,N_3273,N_2939);
or U4906 (N_4906,N_2531,N_3397);
and U4907 (N_4907,N_3339,N_2074);
nand U4908 (N_4908,N_2501,N_2408);
nand U4909 (N_4909,N_2948,N_2464);
nor U4910 (N_4910,N_3410,N_3383);
or U4911 (N_4911,N_2223,N_3001);
nor U4912 (N_4912,N_3588,N_3539);
or U4913 (N_4913,N_3603,N_2747);
nand U4914 (N_4914,N_3161,N_3749);
nor U4915 (N_4915,N_2183,N_2114);
nor U4916 (N_4916,N_2459,N_3633);
nor U4917 (N_4917,N_2294,N_3080);
nand U4918 (N_4918,N_2395,N_3104);
or U4919 (N_4919,N_2446,N_2129);
or U4920 (N_4920,N_2690,N_3570);
nor U4921 (N_4921,N_3592,N_3717);
xnor U4922 (N_4922,N_2184,N_2340);
nand U4923 (N_4923,N_3707,N_3791);
nand U4924 (N_4924,N_2826,N_2741);
or U4925 (N_4925,N_2134,N_2699);
nor U4926 (N_4926,N_3649,N_3572);
nor U4927 (N_4927,N_3110,N_2765);
and U4928 (N_4928,N_2833,N_3927);
or U4929 (N_4929,N_2683,N_2192);
nand U4930 (N_4930,N_3944,N_2923);
or U4931 (N_4931,N_3721,N_3601);
nor U4932 (N_4932,N_2555,N_2498);
nand U4933 (N_4933,N_2251,N_2627);
and U4934 (N_4934,N_2268,N_3664);
or U4935 (N_4935,N_3830,N_2065);
nand U4936 (N_4936,N_3960,N_3077);
and U4937 (N_4937,N_2067,N_2406);
nor U4938 (N_4938,N_2210,N_2286);
and U4939 (N_4939,N_3843,N_3404);
and U4940 (N_4940,N_2055,N_3127);
or U4941 (N_4941,N_3149,N_2944);
or U4942 (N_4942,N_2776,N_2729);
nor U4943 (N_4943,N_3857,N_2430);
and U4944 (N_4944,N_2141,N_3325);
xor U4945 (N_4945,N_2072,N_2820);
nand U4946 (N_4946,N_2248,N_3040);
nand U4947 (N_4947,N_2898,N_2213);
or U4948 (N_4948,N_2399,N_3793);
and U4949 (N_4949,N_3850,N_2648);
and U4950 (N_4950,N_2921,N_3574);
and U4951 (N_4951,N_2085,N_3810);
nand U4952 (N_4952,N_3902,N_3263);
nor U4953 (N_4953,N_2521,N_3854);
or U4954 (N_4954,N_2721,N_2088);
or U4955 (N_4955,N_3842,N_3889);
and U4956 (N_4956,N_2912,N_3748);
nand U4957 (N_4957,N_3340,N_3313);
or U4958 (N_4958,N_2212,N_2382);
nand U4959 (N_4959,N_3193,N_2715);
xnor U4960 (N_4960,N_3347,N_3673);
nand U4961 (N_4961,N_3510,N_3365);
or U4962 (N_4962,N_3958,N_2620);
and U4963 (N_4963,N_2736,N_3939);
and U4964 (N_4964,N_2216,N_2532);
nor U4965 (N_4965,N_2138,N_2500);
and U4966 (N_4966,N_2002,N_2120);
and U4967 (N_4967,N_3505,N_3499);
or U4968 (N_4968,N_2147,N_2954);
nor U4969 (N_4969,N_3419,N_2635);
nor U4970 (N_4970,N_3246,N_3571);
nor U4971 (N_4971,N_3297,N_2232);
or U4972 (N_4972,N_2457,N_2449);
and U4973 (N_4973,N_2186,N_3197);
or U4974 (N_4974,N_2932,N_2917);
nor U4975 (N_4975,N_3568,N_2737);
nor U4976 (N_4976,N_2078,N_3284);
nand U4977 (N_4977,N_3774,N_2111);
nor U4978 (N_4978,N_2874,N_2569);
nor U4979 (N_4979,N_3757,N_2872);
and U4980 (N_4980,N_2150,N_3234);
nand U4981 (N_4981,N_2458,N_3456);
nand U4982 (N_4982,N_3178,N_3634);
nor U4983 (N_4983,N_3928,N_3316);
or U4984 (N_4984,N_3638,N_2321);
nor U4985 (N_4985,N_3642,N_2386);
and U4986 (N_4986,N_2155,N_3866);
or U4987 (N_4987,N_2246,N_2560);
or U4988 (N_4988,N_2711,N_2725);
nand U4989 (N_4989,N_3141,N_3680);
nor U4990 (N_4990,N_3319,N_3108);
and U4991 (N_4991,N_2920,N_3868);
nor U4992 (N_4992,N_2354,N_2892);
nor U4993 (N_4993,N_2187,N_2581);
nand U4994 (N_4994,N_3155,N_3249);
or U4995 (N_4995,N_2762,N_3509);
nand U4996 (N_4996,N_3936,N_3382);
and U4997 (N_4997,N_2001,N_2712);
nand U4998 (N_4998,N_2977,N_2006);
and U4999 (N_4999,N_3573,N_2545);
nor U5000 (N_5000,N_3915,N_3714);
nor U5001 (N_5001,N_3583,N_3587);
and U5002 (N_5002,N_2742,N_3495);
nand U5003 (N_5003,N_3431,N_2745);
or U5004 (N_5004,N_2234,N_2553);
nand U5005 (N_5005,N_2156,N_3511);
nand U5006 (N_5006,N_2591,N_3432);
and U5007 (N_5007,N_2327,N_2951);
and U5008 (N_5008,N_2477,N_2545);
nor U5009 (N_5009,N_3324,N_3594);
or U5010 (N_5010,N_3940,N_2328);
nor U5011 (N_5011,N_2993,N_2499);
or U5012 (N_5012,N_2642,N_3333);
xor U5013 (N_5013,N_3756,N_2041);
and U5014 (N_5014,N_2617,N_2515);
nand U5015 (N_5015,N_2128,N_2220);
nand U5016 (N_5016,N_2578,N_2001);
nand U5017 (N_5017,N_3866,N_2373);
nor U5018 (N_5018,N_2123,N_3153);
or U5019 (N_5019,N_2880,N_3256);
and U5020 (N_5020,N_3017,N_2579);
or U5021 (N_5021,N_3386,N_3574);
nand U5022 (N_5022,N_2195,N_2176);
nand U5023 (N_5023,N_3416,N_2763);
nor U5024 (N_5024,N_3590,N_2161);
and U5025 (N_5025,N_2897,N_3517);
and U5026 (N_5026,N_2935,N_3769);
and U5027 (N_5027,N_3110,N_2467);
nor U5028 (N_5028,N_3671,N_2962);
nor U5029 (N_5029,N_3571,N_3551);
nand U5030 (N_5030,N_3856,N_2040);
nand U5031 (N_5031,N_3814,N_2836);
or U5032 (N_5032,N_2886,N_2312);
and U5033 (N_5033,N_3254,N_2352);
nand U5034 (N_5034,N_3550,N_3956);
and U5035 (N_5035,N_2721,N_3143);
and U5036 (N_5036,N_3447,N_3993);
and U5037 (N_5037,N_3895,N_2203);
and U5038 (N_5038,N_2366,N_2772);
nor U5039 (N_5039,N_2364,N_2555);
or U5040 (N_5040,N_2559,N_2781);
nor U5041 (N_5041,N_3172,N_3805);
and U5042 (N_5042,N_2026,N_3689);
or U5043 (N_5043,N_2178,N_2014);
and U5044 (N_5044,N_2194,N_2449);
nand U5045 (N_5045,N_2810,N_2714);
nand U5046 (N_5046,N_2841,N_3023);
nor U5047 (N_5047,N_3376,N_2379);
or U5048 (N_5048,N_3845,N_3175);
or U5049 (N_5049,N_3987,N_2260);
or U5050 (N_5050,N_2265,N_3551);
or U5051 (N_5051,N_2156,N_3158);
nand U5052 (N_5052,N_3871,N_2086);
nor U5053 (N_5053,N_2023,N_3621);
nand U5054 (N_5054,N_3199,N_3620);
nand U5055 (N_5055,N_2482,N_3995);
and U5056 (N_5056,N_3259,N_2956);
or U5057 (N_5057,N_2537,N_3345);
and U5058 (N_5058,N_2611,N_2908);
or U5059 (N_5059,N_2252,N_3957);
nand U5060 (N_5060,N_2157,N_2030);
nand U5061 (N_5061,N_3915,N_2335);
and U5062 (N_5062,N_2725,N_2840);
nand U5063 (N_5063,N_3319,N_3250);
and U5064 (N_5064,N_3616,N_3798);
nand U5065 (N_5065,N_3374,N_3048);
nand U5066 (N_5066,N_3244,N_3751);
nand U5067 (N_5067,N_3736,N_3655);
nand U5068 (N_5068,N_2887,N_3021);
nand U5069 (N_5069,N_2551,N_3501);
and U5070 (N_5070,N_3325,N_2676);
and U5071 (N_5071,N_3424,N_2443);
and U5072 (N_5072,N_3947,N_3148);
and U5073 (N_5073,N_3662,N_3163);
nor U5074 (N_5074,N_2168,N_3358);
nor U5075 (N_5075,N_3651,N_2722);
nand U5076 (N_5076,N_3885,N_2823);
or U5077 (N_5077,N_3162,N_3021);
nor U5078 (N_5078,N_2528,N_3785);
nand U5079 (N_5079,N_3047,N_3764);
and U5080 (N_5080,N_2003,N_3015);
nor U5081 (N_5081,N_3679,N_2771);
nand U5082 (N_5082,N_2133,N_3554);
or U5083 (N_5083,N_2081,N_2553);
nor U5084 (N_5084,N_3860,N_3445);
nand U5085 (N_5085,N_3087,N_3580);
nor U5086 (N_5086,N_2594,N_2112);
and U5087 (N_5087,N_3519,N_3417);
or U5088 (N_5088,N_3445,N_3823);
nor U5089 (N_5089,N_2734,N_2051);
and U5090 (N_5090,N_3370,N_3230);
nand U5091 (N_5091,N_2684,N_2124);
and U5092 (N_5092,N_2281,N_3435);
and U5093 (N_5093,N_2289,N_2747);
nor U5094 (N_5094,N_3042,N_3129);
nand U5095 (N_5095,N_2253,N_2242);
nor U5096 (N_5096,N_2982,N_3254);
or U5097 (N_5097,N_2561,N_3016);
nor U5098 (N_5098,N_2713,N_3130);
nor U5099 (N_5099,N_3155,N_3135);
nand U5100 (N_5100,N_2662,N_2888);
or U5101 (N_5101,N_2386,N_3974);
nor U5102 (N_5102,N_2738,N_3806);
or U5103 (N_5103,N_2058,N_3066);
or U5104 (N_5104,N_2773,N_3092);
nor U5105 (N_5105,N_3549,N_2010);
nand U5106 (N_5106,N_2316,N_3930);
nor U5107 (N_5107,N_3678,N_2053);
nand U5108 (N_5108,N_2818,N_3816);
nand U5109 (N_5109,N_2886,N_3767);
nor U5110 (N_5110,N_3892,N_2369);
and U5111 (N_5111,N_3543,N_3128);
nor U5112 (N_5112,N_3385,N_3122);
and U5113 (N_5113,N_3730,N_2774);
nand U5114 (N_5114,N_2851,N_3586);
nor U5115 (N_5115,N_2901,N_3637);
nand U5116 (N_5116,N_2942,N_2140);
and U5117 (N_5117,N_3420,N_3215);
nor U5118 (N_5118,N_2222,N_2497);
nand U5119 (N_5119,N_2598,N_2324);
or U5120 (N_5120,N_3103,N_3757);
or U5121 (N_5121,N_3878,N_2492);
and U5122 (N_5122,N_2577,N_3148);
nor U5123 (N_5123,N_3928,N_3302);
and U5124 (N_5124,N_3892,N_2031);
nor U5125 (N_5125,N_3078,N_2704);
nand U5126 (N_5126,N_2681,N_2272);
nand U5127 (N_5127,N_2701,N_3483);
nand U5128 (N_5128,N_2254,N_2375);
nand U5129 (N_5129,N_2469,N_3796);
or U5130 (N_5130,N_3270,N_2253);
or U5131 (N_5131,N_2167,N_2855);
nand U5132 (N_5132,N_2275,N_3253);
nand U5133 (N_5133,N_2971,N_2306);
xor U5134 (N_5134,N_2203,N_3821);
nand U5135 (N_5135,N_2024,N_3337);
or U5136 (N_5136,N_2233,N_3024);
nor U5137 (N_5137,N_3905,N_3549);
or U5138 (N_5138,N_2519,N_3440);
nor U5139 (N_5139,N_2021,N_2360);
and U5140 (N_5140,N_2912,N_2428);
or U5141 (N_5141,N_3782,N_2108);
nor U5142 (N_5142,N_2853,N_2258);
or U5143 (N_5143,N_3818,N_2302);
nor U5144 (N_5144,N_2464,N_2946);
nor U5145 (N_5145,N_3786,N_2700);
or U5146 (N_5146,N_3112,N_2976);
or U5147 (N_5147,N_3196,N_2797);
and U5148 (N_5148,N_3282,N_3801);
nor U5149 (N_5149,N_3363,N_3892);
and U5150 (N_5150,N_3021,N_3799);
or U5151 (N_5151,N_2467,N_2149);
nor U5152 (N_5152,N_2459,N_3215);
xnor U5153 (N_5153,N_2141,N_3029);
and U5154 (N_5154,N_3531,N_3082);
or U5155 (N_5155,N_2422,N_3771);
or U5156 (N_5156,N_2642,N_2695);
nor U5157 (N_5157,N_2894,N_3080);
nor U5158 (N_5158,N_3792,N_2595);
and U5159 (N_5159,N_3393,N_3454);
and U5160 (N_5160,N_2506,N_2667);
or U5161 (N_5161,N_2753,N_2775);
nand U5162 (N_5162,N_2403,N_3126);
nand U5163 (N_5163,N_2959,N_2302);
nor U5164 (N_5164,N_3234,N_2917);
nand U5165 (N_5165,N_2540,N_3791);
nor U5166 (N_5166,N_2708,N_3211);
or U5167 (N_5167,N_3202,N_3872);
nand U5168 (N_5168,N_3045,N_3389);
and U5169 (N_5169,N_2375,N_3968);
nor U5170 (N_5170,N_2343,N_3317);
or U5171 (N_5171,N_2421,N_2375);
or U5172 (N_5172,N_3836,N_3675);
nand U5173 (N_5173,N_2019,N_3622);
and U5174 (N_5174,N_2276,N_3625);
nor U5175 (N_5175,N_3377,N_3167);
nor U5176 (N_5176,N_2887,N_2723);
or U5177 (N_5177,N_3367,N_2283);
nor U5178 (N_5178,N_3685,N_2487);
and U5179 (N_5179,N_3301,N_2564);
nand U5180 (N_5180,N_3465,N_2057);
or U5181 (N_5181,N_2193,N_3093);
or U5182 (N_5182,N_3869,N_3375);
nor U5183 (N_5183,N_2910,N_3849);
and U5184 (N_5184,N_2709,N_3555);
nor U5185 (N_5185,N_3727,N_2820);
or U5186 (N_5186,N_3100,N_3742);
and U5187 (N_5187,N_2420,N_2984);
nand U5188 (N_5188,N_2741,N_3034);
nand U5189 (N_5189,N_2697,N_3523);
nand U5190 (N_5190,N_2175,N_3113);
nor U5191 (N_5191,N_3297,N_2396);
nor U5192 (N_5192,N_2731,N_3815);
and U5193 (N_5193,N_2082,N_2484);
nand U5194 (N_5194,N_2701,N_3883);
nand U5195 (N_5195,N_3886,N_2483);
nor U5196 (N_5196,N_2515,N_2311);
nand U5197 (N_5197,N_2879,N_3306);
or U5198 (N_5198,N_2361,N_3509);
and U5199 (N_5199,N_3288,N_3183);
nand U5200 (N_5200,N_3809,N_3770);
nor U5201 (N_5201,N_2435,N_2854);
xnor U5202 (N_5202,N_2140,N_3409);
and U5203 (N_5203,N_3564,N_2243);
and U5204 (N_5204,N_3734,N_2132);
and U5205 (N_5205,N_2759,N_2304);
or U5206 (N_5206,N_3445,N_3784);
and U5207 (N_5207,N_3868,N_2276);
and U5208 (N_5208,N_3387,N_3241);
nor U5209 (N_5209,N_2728,N_3414);
nor U5210 (N_5210,N_3101,N_3861);
or U5211 (N_5211,N_2123,N_3539);
or U5212 (N_5212,N_2034,N_2903);
or U5213 (N_5213,N_2324,N_2698);
nor U5214 (N_5214,N_3195,N_2328);
or U5215 (N_5215,N_2044,N_3163);
and U5216 (N_5216,N_2471,N_2296);
and U5217 (N_5217,N_3279,N_2775);
nand U5218 (N_5218,N_2617,N_3470);
and U5219 (N_5219,N_3299,N_2535);
and U5220 (N_5220,N_3003,N_2341);
nor U5221 (N_5221,N_3442,N_2770);
nand U5222 (N_5222,N_3225,N_2275);
and U5223 (N_5223,N_2356,N_2714);
or U5224 (N_5224,N_2108,N_2425);
nand U5225 (N_5225,N_2723,N_3998);
nor U5226 (N_5226,N_3709,N_3966);
nand U5227 (N_5227,N_2168,N_3560);
nor U5228 (N_5228,N_3808,N_3253);
and U5229 (N_5229,N_3347,N_2613);
nand U5230 (N_5230,N_3229,N_3345);
nor U5231 (N_5231,N_2732,N_3468);
or U5232 (N_5232,N_2649,N_3462);
nor U5233 (N_5233,N_2836,N_2795);
or U5234 (N_5234,N_3177,N_3501);
nand U5235 (N_5235,N_3613,N_3973);
nor U5236 (N_5236,N_2942,N_3320);
nor U5237 (N_5237,N_2821,N_3857);
or U5238 (N_5238,N_2871,N_2609);
or U5239 (N_5239,N_2377,N_3939);
nand U5240 (N_5240,N_3130,N_2042);
or U5241 (N_5241,N_3224,N_2349);
or U5242 (N_5242,N_2862,N_2431);
and U5243 (N_5243,N_3722,N_2592);
or U5244 (N_5244,N_3010,N_3724);
nand U5245 (N_5245,N_3507,N_3828);
nand U5246 (N_5246,N_3784,N_2963);
or U5247 (N_5247,N_2515,N_3375);
and U5248 (N_5248,N_3010,N_2438);
xnor U5249 (N_5249,N_3483,N_3265);
or U5250 (N_5250,N_3827,N_3300);
nor U5251 (N_5251,N_3017,N_2901);
and U5252 (N_5252,N_3674,N_2919);
and U5253 (N_5253,N_3268,N_3741);
xor U5254 (N_5254,N_3008,N_3111);
nor U5255 (N_5255,N_2035,N_2972);
and U5256 (N_5256,N_3266,N_3296);
nor U5257 (N_5257,N_2198,N_2506);
nor U5258 (N_5258,N_2455,N_3404);
nand U5259 (N_5259,N_3811,N_3518);
nor U5260 (N_5260,N_2618,N_3235);
nor U5261 (N_5261,N_3666,N_3060);
nor U5262 (N_5262,N_3432,N_2986);
nand U5263 (N_5263,N_2981,N_3296);
and U5264 (N_5264,N_3828,N_3546);
nor U5265 (N_5265,N_2314,N_2365);
and U5266 (N_5266,N_3617,N_2526);
and U5267 (N_5267,N_3221,N_2498);
and U5268 (N_5268,N_3415,N_2041);
nor U5269 (N_5269,N_2769,N_2137);
nand U5270 (N_5270,N_3440,N_2842);
nand U5271 (N_5271,N_2817,N_2265);
and U5272 (N_5272,N_3977,N_2076);
and U5273 (N_5273,N_3077,N_2408);
or U5274 (N_5274,N_3895,N_3110);
nand U5275 (N_5275,N_2559,N_2122);
and U5276 (N_5276,N_2648,N_3422);
or U5277 (N_5277,N_2378,N_2584);
nand U5278 (N_5278,N_2157,N_2308);
and U5279 (N_5279,N_3951,N_3697);
nor U5280 (N_5280,N_3505,N_2873);
and U5281 (N_5281,N_2476,N_3785);
xor U5282 (N_5282,N_2065,N_3648);
nor U5283 (N_5283,N_2958,N_2229);
and U5284 (N_5284,N_3065,N_3331);
or U5285 (N_5285,N_3875,N_2303);
or U5286 (N_5286,N_3876,N_2405);
nor U5287 (N_5287,N_3802,N_3892);
nor U5288 (N_5288,N_2234,N_3830);
or U5289 (N_5289,N_3826,N_2495);
nor U5290 (N_5290,N_2089,N_3576);
and U5291 (N_5291,N_3507,N_2100);
and U5292 (N_5292,N_3262,N_2689);
nand U5293 (N_5293,N_2734,N_3283);
or U5294 (N_5294,N_2592,N_2063);
nor U5295 (N_5295,N_2719,N_2050);
or U5296 (N_5296,N_2720,N_2678);
and U5297 (N_5297,N_2095,N_2583);
nand U5298 (N_5298,N_2809,N_3512);
nor U5299 (N_5299,N_3076,N_2135);
nor U5300 (N_5300,N_3167,N_2576);
nand U5301 (N_5301,N_3052,N_2497);
or U5302 (N_5302,N_2990,N_3157);
or U5303 (N_5303,N_2581,N_2556);
nand U5304 (N_5304,N_2019,N_2029);
or U5305 (N_5305,N_3795,N_2538);
or U5306 (N_5306,N_2918,N_2581);
or U5307 (N_5307,N_2324,N_2024);
nand U5308 (N_5308,N_2299,N_2751);
or U5309 (N_5309,N_2084,N_2653);
nor U5310 (N_5310,N_2203,N_2622);
nor U5311 (N_5311,N_2436,N_2115);
xnor U5312 (N_5312,N_2831,N_3302);
nand U5313 (N_5313,N_2003,N_2841);
nor U5314 (N_5314,N_2850,N_2337);
and U5315 (N_5315,N_3504,N_2525);
nor U5316 (N_5316,N_2472,N_3257);
or U5317 (N_5317,N_3948,N_2245);
and U5318 (N_5318,N_2422,N_3534);
nand U5319 (N_5319,N_2669,N_3363);
nand U5320 (N_5320,N_2811,N_3633);
nand U5321 (N_5321,N_2991,N_3135);
and U5322 (N_5322,N_3407,N_3732);
and U5323 (N_5323,N_2670,N_2329);
nor U5324 (N_5324,N_2871,N_2288);
or U5325 (N_5325,N_2440,N_2750);
xnor U5326 (N_5326,N_2419,N_3731);
nand U5327 (N_5327,N_2707,N_2563);
nor U5328 (N_5328,N_3523,N_2725);
nand U5329 (N_5329,N_3852,N_3413);
or U5330 (N_5330,N_3655,N_2586);
and U5331 (N_5331,N_2681,N_2871);
or U5332 (N_5332,N_2583,N_3524);
nand U5333 (N_5333,N_3620,N_2327);
nand U5334 (N_5334,N_3825,N_2928);
and U5335 (N_5335,N_2378,N_3800);
and U5336 (N_5336,N_2841,N_2730);
and U5337 (N_5337,N_2300,N_2013);
and U5338 (N_5338,N_2103,N_3985);
and U5339 (N_5339,N_3460,N_2631);
nor U5340 (N_5340,N_2878,N_3278);
nor U5341 (N_5341,N_2645,N_2308);
or U5342 (N_5342,N_2167,N_3089);
and U5343 (N_5343,N_3250,N_3750);
nor U5344 (N_5344,N_3659,N_3695);
and U5345 (N_5345,N_3997,N_3280);
or U5346 (N_5346,N_3347,N_2040);
or U5347 (N_5347,N_2413,N_3141);
nor U5348 (N_5348,N_2915,N_3888);
nor U5349 (N_5349,N_2605,N_3378);
nor U5350 (N_5350,N_2622,N_3285);
or U5351 (N_5351,N_3064,N_2716);
or U5352 (N_5352,N_3200,N_2696);
nand U5353 (N_5353,N_3457,N_2069);
or U5354 (N_5354,N_3210,N_2739);
or U5355 (N_5355,N_3070,N_2938);
or U5356 (N_5356,N_3472,N_2348);
nor U5357 (N_5357,N_3400,N_2883);
nor U5358 (N_5358,N_3390,N_2948);
nand U5359 (N_5359,N_3345,N_3414);
or U5360 (N_5360,N_2101,N_2606);
nor U5361 (N_5361,N_3573,N_3540);
or U5362 (N_5362,N_2272,N_3515);
nand U5363 (N_5363,N_3569,N_2641);
nand U5364 (N_5364,N_3084,N_3080);
or U5365 (N_5365,N_3823,N_3781);
nor U5366 (N_5366,N_2762,N_2297);
and U5367 (N_5367,N_2300,N_2117);
and U5368 (N_5368,N_3801,N_3516);
nand U5369 (N_5369,N_2139,N_3405);
nand U5370 (N_5370,N_2359,N_2140);
nand U5371 (N_5371,N_3230,N_3837);
nand U5372 (N_5372,N_2048,N_2008);
nand U5373 (N_5373,N_2623,N_3308);
or U5374 (N_5374,N_2620,N_3532);
nand U5375 (N_5375,N_3703,N_3789);
or U5376 (N_5376,N_2036,N_2226);
or U5377 (N_5377,N_3467,N_2126);
nand U5378 (N_5378,N_2707,N_2270);
nor U5379 (N_5379,N_2099,N_2491);
or U5380 (N_5380,N_2023,N_3185);
nor U5381 (N_5381,N_3681,N_2936);
or U5382 (N_5382,N_3644,N_3202);
or U5383 (N_5383,N_3193,N_2471);
nor U5384 (N_5384,N_2068,N_2283);
nand U5385 (N_5385,N_2963,N_3351);
or U5386 (N_5386,N_2389,N_3195);
nor U5387 (N_5387,N_2351,N_3193);
nor U5388 (N_5388,N_2048,N_3047);
xnor U5389 (N_5389,N_2355,N_2125);
nand U5390 (N_5390,N_3208,N_3982);
nor U5391 (N_5391,N_2445,N_3462);
nor U5392 (N_5392,N_3472,N_3861);
or U5393 (N_5393,N_2792,N_2034);
and U5394 (N_5394,N_2708,N_2232);
and U5395 (N_5395,N_3693,N_3924);
nand U5396 (N_5396,N_2509,N_3666);
nor U5397 (N_5397,N_2286,N_2311);
or U5398 (N_5398,N_2745,N_2901);
nor U5399 (N_5399,N_3923,N_3816);
nor U5400 (N_5400,N_3851,N_3417);
nand U5401 (N_5401,N_3788,N_3344);
and U5402 (N_5402,N_3761,N_3304);
or U5403 (N_5403,N_2601,N_2921);
or U5404 (N_5404,N_2084,N_3631);
and U5405 (N_5405,N_3264,N_2154);
and U5406 (N_5406,N_2862,N_3840);
or U5407 (N_5407,N_3028,N_3975);
nand U5408 (N_5408,N_2585,N_3579);
or U5409 (N_5409,N_2980,N_3349);
or U5410 (N_5410,N_3237,N_3723);
and U5411 (N_5411,N_2294,N_3465);
nand U5412 (N_5412,N_3771,N_2746);
and U5413 (N_5413,N_2134,N_3823);
and U5414 (N_5414,N_2524,N_3514);
nand U5415 (N_5415,N_2630,N_3656);
nand U5416 (N_5416,N_3213,N_2210);
or U5417 (N_5417,N_2931,N_2445);
and U5418 (N_5418,N_3563,N_3669);
nor U5419 (N_5419,N_3645,N_3204);
or U5420 (N_5420,N_3227,N_3584);
nor U5421 (N_5421,N_3727,N_3218);
nand U5422 (N_5422,N_2347,N_2459);
and U5423 (N_5423,N_2631,N_3658);
nor U5424 (N_5424,N_2168,N_3659);
and U5425 (N_5425,N_3612,N_3174);
and U5426 (N_5426,N_2525,N_2776);
nand U5427 (N_5427,N_2852,N_3350);
nand U5428 (N_5428,N_3664,N_2269);
nor U5429 (N_5429,N_3703,N_3348);
nand U5430 (N_5430,N_3640,N_3302);
nand U5431 (N_5431,N_3296,N_3057);
nor U5432 (N_5432,N_3127,N_3959);
and U5433 (N_5433,N_3895,N_2189);
nor U5434 (N_5434,N_3152,N_3256);
nor U5435 (N_5435,N_3061,N_2435);
nor U5436 (N_5436,N_2839,N_2538);
nand U5437 (N_5437,N_2748,N_3708);
nand U5438 (N_5438,N_2607,N_3756);
and U5439 (N_5439,N_2297,N_2135);
nand U5440 (N_5440,N_3951,N_2071);
nand U5441 (N_5441,N_3782,N_2910);
or U5442 (N_5442,N_3601,N_3492);
or U5443 (N_5443,N_2433,N_2389);
nand U5444 (N_5444,N_2537,N_2778);
nand U5445 (N_5445,N_3282,N_2953);
or U5446 (N_5446,N_2802,N_3768);
nor U5447 (N_5447,N_2614,N_2366);
or U5448 (N_5448,N_3702,N_2217);
nand U5449 (N_5449,N_2960,N_2825);
nor U5450 (N_5450,N_2923,N_2087);
and U5451 (N_5451,N_3653,N_2272);
or U5452 (N_5452,N_3259,N_3568);
and U5453 (N_5453,N_2212,N_3136);
or U5454 (N_5454,N_3142,N_3413);
or U5455 (N_5455,N_3437,N_3483);
or U5456 (N_5456,N_3728,N_3942);
or U5457 (N_5457,N_2969,N_2422);
nor U5458 (N_5458,N_3491,N_2487);
or U5459 (N_5459,N_2758,N_3841);
xnor U5460 (N_5460,N_3057,N_2083);
nor U5461 (N_5461,N_2386,N_2927);
nor U5462 (N_5462,N_2933,N_3759);
and U5463 (N_5463,N_2424,N_2047);
and U5464 (N_5464,N_2525,N_3274);
nand U5465 (N_5465,N_3431,N_3199);
nand U5466 (N_5466,N_2745,N_3470);
or U5467 (N_5467,N_3171,N_2251);
or U5468 (N_5468,N_2174,N_2708);
or U5469 (N_5469,N_3385,N_2511);
and U5470 (N_5470,N_2878,N_2328);
nand U5471 (N_5471,N_2727,N_2666);
nor U5472 (N_5472,N_3919,N_2165);
nand U5473 (N_5473,N_2225,N_3514);
or U5474 (N_5474,N_3587,N_2420);
nor U5475 (N_5475,N_2143,N_3009);
xor U5476 (N_5476,N_3932,N_3964);
nand U5477 (N_5477,N_3073,N_2994);
nand U5478 (N_5478,N_3814,N_3309);
nor U5479 (N_5479,N_2135,N_3558);
nand U5480 (N_5480,N_3772,N_3707);
and U5481 (N_5481,N_3082,N_3414);
or U5482 (N_5482,N_2638,N_3909);
nor U5483 (N_5483,N_2545,N_2599);
or U5484 (N_5484,N_3407,N_3946);
nor U5485 (N_5485,N_2314,N_2526);
or U5486 (N_5486,N_2189,N_3424);
or U5487 (N_5487,N_2645,N_2188);
and U5488 (N_5488,N_3766,N_3278);
nand U5489 (N_5489,N_2379,N_3599);
and U5490 (N_5490,N_2512,N_3922);
nor U5491 (N_5491,N_2078,N_3016);
or U5492 (N_5492,N_2719,N_2029);
and U5493 (N_5493,N_3446,N_3380);
xor U5494 (N_5494,N_3260,N_3929);
and U5495 (N_5495,N_3813,N_2884);
nor U5496 (N_5496,N_3484,N_2505);
nor U5497 (N_5497,N_2776,N_2170);
or U5498 (N_5498,N_3240,N_2480);
nand U5499 (N_5499,N_3455,N_2402);
and U5500 (N_5500,N_2997,N_3097);
nand U5501 (N_5501,N_2368,N_2239);
or U5502 (N_5502,N_3765,N_2373);
or U5503 (N_5503,N_3958,N_2926);
or U5504 (N_5504,N_3373,N_2534);
nor U5505 (N_5505,N_3383,N_3779);
nor U5506 (N_5506,N_2686,N_3962);
or U5507 (N_5507,N_2540,N_2562);
nor U5508 (N_5508,N_3080,N_3258);
or U5509 (N_5509,N_3923,N_2111);
and U5510 (N_5510,N_2079,N_3628);
or U5511 (N_5511,N_3934,N_2231);
nor U5512 (N_5512,N_2958,N_2120);
nor U5513 (N_5513,N_2032,N_3240);
or U5514 (N_5514,N_3678,N_2838);
nand U5515 (N_5515,N_3901,N_3578);
and U5516 (N_5516,N_3393,N_2955);
xor U5517 (N_5517,N_3142,N_3746);
and U5518 (N_5518,N_2488,N_3284);
nand U5519 (N_5519,N_3003,N_3518);
and U5520 (N_5520,N_3763,N_3426);
or U5521 (N_5521,N_3615,N_2663);
or U5522 (N_5522,N_3093,N_3653);
nand U5523 (N_5523,N_3080,N_2896);
nand U5524 (N_5524,N_2665,N_3992);
nor U5525 (N_5525,N_3759,N_2466);
or U5526 (N_5526,N_3862,N_3058);
xnor U5527 (N_5527,N_3250,N_2272);
nand U5528 (N_5528,N_3885,N_3868);
nor U5529 (N_5529,N_3864,N_3676);
nor U5530 (N_5530,N_2119,N_3400);
or U5531 (N_5531,N_3441,N_3011);
nor U5532 (N_5532,N_2304,N_2477);
nand U5533 (N_5533,N_2433,N_3572);
nor U5534 (N_5534,N_3813,N_2078);
or U5535 (N_5535,N_3812,N_2502);
and U5536 (N_5536,N_3159,N_3339);
xor U5537 (N_5537,N_3448,N_3328);
and U5538 (N_5538,N_2038,N_2275);
and U5539 (N_5539,N_2804,N_2331);
xor U5540 (N_5540,N_2869,N_3003);
and U5541 (N_5541,N_3188,N_3571);
or U5542 (N_5542,N_2080,N_2635);
or U5543 (N_5543,N_3844,N_3975);
or U5544 (N_5544,N_2293,N_2357);
nand U5545 (N_5545,N_2332,N_3716);
or U5546 (N_5546,N_3456,N_2148);
nor U5547 (N_5547,N_3697,N_2836);
and U5548 (N_5548,N_3803,N_2222);
nand U5549 (N_5549,N_3416,N_2150);
or U5550 (N_5550,N_3190,N_3380);
xnor U5551 (N_5551,N_3575,N_3251);
nor U5552 (N_5552,N_3797,N_2796);
or U5553 (N_5553,N_2805,N_3388);
nor U5554 (N_5554,N_3280,N_3775);
nor U5555 (N_5555,N_2738,N_2884);
nor U5556 (N_5556,N_3265,N_2684);
or U5557 (N_5557,N_2648,N_3618);
or U5558 (N_5558,N_3737,N_2315);
and U5559 (N_5559,N_2374,N_3309);
and U5560 (N_5560,N_2872,N_2083);
nor U5561 (N_5561,N_2738,N_3520);
nand U5562 (N_5562,N_2750,N_2442);
nand U5563 (N_5563,N_2289,N_3982);
nand U5564 (N_5564,N_3701,N_3537);
xor U5565 (N_5565,N_2355,N_3007);
nor U5566 (N_5566,N_2886,N_3478);
and U5567 (N_5567,N_3637,N_2740);
xor U5568 (N_5568,N_3685,N_3985);
and U5569 (N_5569,N_2472,N_2988);
nand U5570 (N_5570,N_3883,N_3799);
nand U5571 (N_5571,N_3167,N_3276);
nand U5572 (N_5572,N_2178,N_2719);
nand U5573 (N_5573,N_2231,N_2743);
or U5574 (N_5574,N_3525,N_2476);
nand U5575 (N_5575,N_2258,N_2654);
and U5576 (N_5576,N_3760,N_2844);
nor U5577 (N_5577,N_2857,N_2630);
and U5578 (N_5578,N_3717,N_3333);
and U5579 (N_5579,N_3968,N_2177);
nor U5580 (N_5580,N_3533,N_2072);
nor U5581 (N_5581,N_2458,N_3429);
and U5582 (N_5582,N_2481,N_3965);
nor U5583 (N_5583,N_2083,N_2679);
nor U5584 (N_5584,N_3877,N_2679);
nor U5585 (N_5585,N_3214,N_3097);
xnor U5586 (N_5586,N_3553,N_2741);
or U5587 (N_5587,N_2708,N_3992);
or U5588 (N_5588,N_2526,N_2819);
nor U5589 (N_5589,N_2822,N_2138);
and U5590 (N_5590,N_2532,N_3542);
nand U5591 (N_5591,N_2572,N_3589);
nand U5592 (N_5592,N_3708,N_3879);
nor U5593 (N_5593,N_2308,N_2849);
nor U5594 (N_5594,N_3156,N_2357);
or U5595 (N_5595,N_3876,N_3455);
or U5596 (N_5596,N_3294,N_2732);
nor U5597 (N_5597,N_3413,N_2855);
and U5598 (N_5598,N_3779,N_2995);
and U5599 (N_5599,N_3262,N_3685);
or U5600 (N_5600,N_3559,N_3242);
nand U5601 (N_5601,N_3762,N_2122);
or U5602 (N_5602,N_3806,N_2942);
nand U5603 (N_5603,N_3479,N_3436);
nand U5604 (N_5604,N_3658,N_2042);
or U5605 (N_5605,N_2526,N_2626);
and U5606 (N_5606,N_2922,N_2291);
and U5607 (N_5607,N_3686,N_2078);
nand U5608 (N_5608,N_2789,N_2942);
nand U5609 (N_5609,N_2906,N_2905);
or U5610 (N_5610,N_3126,N_2715);
nand U5611 (N_5611,N_3506,N_3632);
and U5612 (N_5612,N_2988,N_2001);
xnor U5613 (N_5613,N_2433,N_3837);
nor U5614 (N_5614,N_2061,N_3275);
or U5615 (N_5615,N_2222,N_3911);
nand U5616 (N_5616,N_2126,N_2796);
nor U5617 (N_5617,N_2309,N_2990);
and U5618 (N_5618,N_2964,N_3664);
nand U5619 (N_5619,N_2036,N_2954);
xnor U5620 (N_5620,N_3143,N_2276);
and U5621 (N_5621,N_2182,N_3474);
nand U5622 (N_5622,N_2314,N_2143);
and U5623 (N_5623,N_3808,N_3587);
nor U5624 (N_5624,N_3619,N_2029);
and U5625 (N_5625,N_3154,N_2559);
or U5626 (N_5626,N_3841,N_2522);
xor U5627 (N_5627,N_2252,N_3401);
nand U5628 (N_5628,N_2857,N_3380);
nor U5629 (N_5629,N_2128,N_3123);
and U5630 (N_5630,N_2418,N_3612);
nor U5631 (N_5631,N_2489,N_2502);
nand U5632 (N_5632,N_3811,N_2198);
and U5633 (N_5633,N_2456,N_3200);
or U5634 (N_5634,N_3512,N_2915);
and U5635 (N_5635,N_2245,N_3151);
nand U5636 (N_5636,N_2731,N_3246);
nand U5637 (N_5637,N_3495,N_3278);
and U5638 (N_5638,N_3327,N_3833);
nor U5639 (N_5639,N_3514,N_3622);
and U5640 (N_5640,N_2432,N_2954);
and U5641 (N_5641,N_3946,N_2886);
and U5642 (N_5642,N_3365,N_3236);
or U5643 (N_5643,N_3250,N_3371);
and U5644 (N_5644,N_2759,N_3625);
nor U5645 (N_5645,N_2984,N_2656);
nor U5646 (N_5646,N_3282,N_2151);
nand U5647 (N_5647,N_3058,N_3577);
and U5648 (N_5648,N_3920,N_2597);
nand U5649 (N_5649,N_2581,N_3255);
nand U5650 (N_5650,N_3333,N_2645);
nand U5651 (N_5651,N_2875,N_2715);
or U5652 (N_5652,N_3899,N_2958);
or U5653 (N_5653,N_3891,N_3552);
nor U5654 (N_5654,N_2100,N_3196);
nor U5655 (N_5655,N_2992,N_3915);
nand U5656 (N_5656,N_3847,N_3422);
nand U5657 (N_5657,N_3933,N_3214);
or U5658 (N_5658,N_3194,N_2968);
or U5659 (N_5659,N_2392,N_2762);
nor U5660 (N_5660,N_3678,N_2726);
or U5661 (N_5661,N_3120,N_3841);
or U5662 (N_5662,N_3137,N_3765);
and U5663 (N_5663,N_2116,N_2387);
nand U5664 (N_5664,N_2365,N_2025);
nor U5665 (N_5665,N_2609,N_2389);
and U5666 (N_5666,N_3343,N_3014);
nand U5667 (N_5667,N_3978,N_2497);
nand U5668 (N_5668,N_2947,N_3048);
and U5669 (N_5669,N_2523,N_3999);
or U5670 (N_5670,N_3124,N_2285);
or U5671 (N_5671,N_3868,N_2019);
nand U5672 (N_5672,N_2554,N_3843);
or U5673 (N_5673,N_3093,N_3400);
xnor U5674 (N_5674,N_3631,N_2201);
nor U5675 (N_5675,N_2192,N_2127);
nand U5676 (N_5676,N_2387,N_3739);
nand U5677 (N_5677,N_3441,N_2601);
and U5678 (N_5678,N_2015,N_2311);
nor U5679 (N_5679,N_2602,N_3293);
and U5680 (N_5680,N_2183,N_2040);
xor U5681 (N_5681,N_3975,N_3610);
xor U5682 (N_5682,N_2038,N_3819);
and U5683 (N_5683,N_3044,N_3165);
or U5684 (N_5684,N_3763,N_2297);
nor U5685 (N_5685,N_2079,N_2434);
or U5686 (N_5686,N_2383,N_3863);
or U5687 (N_5687,N_3024,N_2551);
nor U5688 (N_5688,N_2118,N_2842);
nand U5689 (N_5689,N_3407,N_2537);
nor U5690 (N_5690,N_3274,N_3487);
nand U5691 (N_5691,N_2209,N_2357);
nand U5692 (N_5692,N_2267,N_3571);
or U5693 (N_5693,N_3492,N_3308);
or U5694 (N_5694,N_2633,N_3054);
nor U5695 (N_5695,N_3094,N_3066);
and U5696 (N_5696,N_2126,N_3745);
and U5697 (N_5697,N_3804,N_3627);
and U5698 (N_5698,N_2156,N_2496);
and U5699 (N_5699,N_3083,N_3021);
nand U5700 (N_5700,N_3575,N_3443);
nand U5701 (N_5701,N_3567,N_3474);
or U5702 (N_5702,N_3674,N_2627);
nand U5703 (N_5703,N_3511,N_2590);
nand U5704 (N_5704,N_3049,N_3233);
nand U5705 (N_5705,N_2791,N_3539);
and U5706 (N_5706,N_3712,N_2431);
nand U5707 (N_5707,N_2019,N_2574);
nand U5708 (N_5708,N_3598,N_2278);
nor U5709 (N_5709,N_3993,N_3656);
nor U5710 (N_5710,N_3935,N_3434);
and U5711 (N_5711,N_3359,N_3138);
and U5712 (N_5712,N_2526,N_2681);
or U5713 (N_5713,N_3627,N_2401);
and U5714 (N_5714,N_2356,N_2780);
or U5715 (N_5715,N_2367,N_2724);
nand U5716 (N_5716,N_3808,N_3937);
xor U5717 (N_5717,N_2945,N_3608);
and U5718 (N_5718,N_3147,N_2955);
nor U5719 (N_5719,N_3651,N_2162);
or U5720 (N_5720,N_3808,N_3009);
nand U5721 (N_5721,N_2454,N_2887);
and U5722 (N_5722,N_3596,N_2541);
nand U5723 (N_5723,N_2810,N_2014);
nand U5724 (N_5724,N_3503,N_2604);
nand U5725 (N_5725,N_3146,N_2516);
xor U5726 (N_5726,N_2703,N_3520);
or U5727 (N_5727,N_2989,N_2065);
or U5728 (N_5728,N_3987,N_2922);
and U5729 (N_5729,N_3148,N_2200);
nor U5730 (N_5730,N_3631,N_3951);
nand U5731 (N_5731,N_3929,N_2087);
nor U5732 (N_5732,N_2968,N_3486);
nand U5733 (N_5733,N_3409,N_2192);
nor U5734 (N_5734,N_2291,N_3902);
or U5735 (N_5735,N_2927,N_2956);
nor U5736 (N_5736,N_3979,N_3228);
nand U5737 (N_5737,N_2304,N_2205);
nor U5738 (N_5738,N_3172,N_2081);
and U5739 (N_5739,N_3603,N_3510);
nand U5740 (N_5740,N_2481,N_3816);
nor U5741 (N_5741,N_2817,N_2944);
and U5742 (N_5742,N_3360,N_3519);
and U5743 (N_5743,N_3553,N_3823);
nand U5744 (N_5744,N_3478,N_2325);
or U5745 (N_5745,N_3187,N_3319);
or U5746 (N_5746,N_2819,N_2872);
or U5747 (N_5747,N_2863,N_3118);
and U5748 (N_5748,N_3415,N_3919);
or U5749 (N_5749,N_2169,N_2297);
or U5750 (N_5750,N_3415,N_3972);
nor U5751 (N_5751,N_2306,N_2962);
nand U5752 (N_5752,N_2729,N_3367);
nand U5753 (N_5753,N_3876,N_3847);
or U5754 (N_5754,N_3834,N_2121);
nand U5755 (N_5755,N_2762,N_3527);
and U5756 (N_5756,N_3027,N_3932);
and U5757 (N_5757,N_2329,N_2498);
or U5758 (N_5758,N_2788,N_2609);
or U5759 (N_5759,N_2634,N_2667);
nand U5760 (N_5760,N_3172,N_3361);
xor U5761 (N_5761,N_2432,N_2896);
or U5762 (N_5762,N_3454,N_3677);
and U5763 (N_5763,N_2100,N_2058);
or U5764 (N_5764,N_2773,N_2792);
and U5765 (N_5765,N_3901,N_2620);
and U5766 (N_5766,N_2458,N_2376);
nor U5767 (N_5767,N_2803,N_3342);
and U5768 (N_5768,N_3998,N_3200);
nor U5769 (N_5769,N_2233,N_3604);
and U5770 (N_5770,N_2714,N_2922);
nand U5771 (N_5771,N_3780,N_2595);
or U5772 (N_5772,N_3437,N_2722);
or U5773 (N_5773,N_3031,N_2134);
nor U5774 (N_5774,N_3660,N_2622);
nor U5775 (N_5775,N_3513,N_3586);
or U5776 (N_5776,N_2062,N_2735);
nand U5777 (N_5777,N_2614,N_2256);
nand U5778 (N_5778,N_3326,N_2556);
nor U5779 (N_5779,N_3324,N_3793);
nand U5780 (N_5780,N_3057,N_2009);
nor U5781 (N_5781,N_3664,N_2164);
nor U5782 (N_5782,N_3933,N_2222);
or U5783 (N_5783,N_2901,N_3675);
or U5784 (N_5784,N_2292,N_3975);
or U5785 (N_5785,N_3647,N_2325);
or U5786 (N_5786,N_2738,N_3236);
nand U5787 (N_5787,N_3394,N_3924);
xnor U5788 (N_5788,N_2794,N_2143);
and U5789 (N_5789,N_3887,N_2890);
or U5790 (N_5790,N_3569,N_3000);
nand U5791 (N_5791,N_2372,N_3079);
and U5792 (N_5792,N_3907,N_2448);
nor U5793 (N_5793,N_2454,N_2493);
or U5794 (N_5794,N_2860,N_3976);
nand U5795 (N_5795,N_2349,N_2363);
xor U5796 (N_5796,N_3563,N_2146);
or U5797 (N_5797,N_2320,N_2209);
nand U5798 (N_5798,N_2630,N_3179);
and U5799 (N_5799,N_3307,N_2144);
or U5800 (N_5800,N_3831,N_2333);
nor U5801 (N_5801,N_3853,N_2524);
and U5802 (N_5802,N_3131,N_3184);
and U5803 (N_5803,N_2176,N_3170);
and U5804 (N_5804,N_3314,N_3550);
and U5805 (N_5805,N_3554,N_3177);
or U5806 (N_5806,N_3750,N_3116);
and U5807 (N_5807,N_3309,N_3294);
or U5808 (N_5808,N_2740,N_2251);
and U5809 (N_5809,N_3680,N_3371);
and U5810 (N_5810,N_2368,N_3046);
or U5811 (N_5811,N_2211,N_2314);
nor U5812 (N_5812,N_2015,N_2763);
and U5813 (N_5813,N_3366,N_2579);
and U5814 (N_5814,N_3671,N_3755);
nor U5815 (N_5815,N_3908,N_2472);
nor U5816 (N_5816,N_2313,N_2234);
and U5817 (N_5817,N_2061,N_3386);
and U5818 (N_5818,N_3385,N_3864);
or U5819 (N_5819,N_3386,N_3703);
and U5820 (N_5820,N_2689,N_3263);
and U5821 (N_5821,N_2380,N_3936);
and U5822 (N_5822,N_2611,N_2986);
and U5823 (N_5823,N_3336,N_3304);
xor U5824 (N_5824,N_3637,N_3069);
nor U5825 (N_5825,N_3081,N_3964);
nand U5826 (N_5826,N_2460,N_3087);
or U5827 (N_5827,N_3938,N_2587);
nand U5828 (N_5828,N_2609,N_2213);
and U5829 (N_5829,N_3921,N_3776);
and U5830 (N_5830,N_3646,N_2810);
and U5831 (N_5831,N_2077,N_2964);
and U5832 (N_5832,N_2224,N_2211);
and U5833 (N_5833,N_3931,N_2752);
nand U5834 (N_5834,N_3267,N_2016);
nor U5835 (N_5835,N_3911,N_2082);
xnor U5836 (N_5836,N_2448,N_3366);
or U5837 (N_5837,N_2653,N_2372);
nand U5838 (N_5838,N_2928,N_2954);
xnor U5839 (N_5839,N_2631,N_2259);
and U5840 (N_5840,N_3564,N_3328);
or U5841 (N_5841,N_2340,N_3837);
and U5842 (N_5842,N_3601,N_3105);
or U5843 (N_5843,N_3479,N_3910);
nand U5844 (N_5844,N_3945,N_2181);
and U5845 (N_5845,N_2002,N_2122);
nor U5846 (N_5846,N_2722,N_2713);
or U5847 (N_5847,N_3563,N_2759);
nor U5848 (N_5848,N_3096,N_2190);
or U5849 (N_5849,N_2172,N_2569);
nor U5850 (N_5850,N_2924,N_3431);
or U5851 (N_5851,N_2865,N_2814);
nor U5852 (N_5852,N_2135,N_2097);
nand U5853 (N_5853,N_2107,N_2019);
or U5854 (N_5854,N_3122,N_2987);
or U5855 (N_5855,N_3777,N_3652);
nor U5856 (N_5856,N_3321,N_2101);
or U5857 (N_5857,N_3478,N_3578);
nor U5858 (N_5858,N_2238,N_3450);
nor U5859 (N_5859,N_3464,N_3049);
nand U5860 (N_5860,N_3880,N_2664);
or U5861 (N_5861,N_2522,N_2491);
or U5862 (N_5862,N_3417,N_2029);
or U5863 (N_5863,N_3618,N_3821);
nor U5864 (N_5864,N_3075,N_3278);
nor U5865 (N_5865,N_2784,N_2392);
nor U5866 (N_5866,N_3033,N_2126);
nand U5867 (N_5867,N_2587,N_2063);
nand U5868 (N_5868,N_2702,N_2169);
nor U5869 (N_5869,N_3711,N_3747);
or U5870 (N_5870,N_2186,N_3045);
nand U5871 (N_5871,N_2299,N_2485);
nor U5872 (N_5872,N_2074,N_3885);
nor U5873 (N_5873,N_2397,N_2263);
and U5874 (N_5874,N_3770,N_2800);
or U5875 (N_5875,N_2962,N_2025);
or U5876 (N_5876,N_2012,N_3803);
nor U5877 (N_5877,N_2228,N_3756);
nor U5878 (N_5878,N_3215,N_2457);
or U5879 (N_5879,N_2222,N_3935);
or U5880 (N_5880,N_2058,N_2486);
or U5881 (N_5881,N_2208,N_2936);
nor U5882 (N_5882,N_2811,N_2501);
nor U5883 (N_5883,N_3880,N_2640);
and U5884 (N_5884,N_3106,N_2870);
or U5885 (N_5885,N_3709,N_2692);
or U5886 (N_5886,N_2848,N_3457);
or U5887 (N_5887,N_2787,N_3711);
nand U5888 (N_5888,N_3059,N_2148);
and U5889 (N_5889,N_2687,N_3947);
xor U5890 (N_5890,N_3869,N_3259);
or U5891 (N_5891,N_2007,N_3130);
nor U5892 (N_5892,N_2522,N_2680);
or U5893 (N_5893,N_3439,N_3522);
nand U5894 (N_5894,N_3418,N_3232);
nor U5895 (N_5895,N_2303,N_2984);
nand U5896 (N_5896,N_2512,N_2613);
and U5897 (N_5897,N_3639,N_2733);
or U5898 (N_5898,N_2347,N_2281);
nor U5899 (N_5899,N_2603,N_2092);
or U5900 (N_5900,N_3945,N_2925);
nand U5901 (N_5901,N_3295,N_2774);
and U5902 (N_5902,N_3187,N_3217);
or U5903 (N_5903,N_2343,N_2213);
nor U5904 (N_5904,N_2279,N_3892);
or U5905 (N_5905,N_2830,N_2611);
or U5906 (N_5906,N_3435,N_3073);
or U5907 (N_5907,N_3775,N_2402);
or U5908 (N_5908,N_2909,N_3909);
nor U5909 (N_5909,N_2807,N_2314);
and U5910 (N_5910,N_2074,N_2687);
nand U5911 (N_5911,N_2721,N_2434);
or U5912 (N_5912,N_2344,N_2823);
nand U5913 (N_5913,N_2255,N_2794);
nor U5914 (N_5914,N_3217,N_2653);
or U5915 (N_5915,N_2461,N_2852);
xnor U5916 (N_5916,N_2448,N_3259);
or U5917 (N_5917,N_2571,N_2003);
nand U5918 (N_5918,N_2776,N_2767);
or U5919 (N_5919,N_2147,N_2351);
or U5920 (N_5920,N_2922,N_3631);
and U5921 (N_5921,N_2066,N_3342);
nor U5922 (N_5922,N_2833,N_3876);
or U5923 (N_5923,N_3075,N_2261);
nor U5924 (N_5924,N_2720,N_2782);
or U5925 (N_5925,N_3737,N_3762);
nand U5926 (N_5926,N_2535,N_3903);
nand U5927 (N_5927,N_2075,N_2852);
or U5928 (N_5928,N_2376,N_3929);
nor U5929 (N_5929,N_2941,N_2231);
and U5930 (N_5930,N_3665,N_3177);
xor U5931 (N_5931,N_3401,N_2247);
nand U5932 (N_5932,N_3797,N_3217);
nor U5933 (N_5933,N_2084,N_3768);
nor U5934 (N_5934,N_3563,N_2139);
or U5935 (N_5935,N_2489,N_3556);
nand U5936 (N_5936,N_3114,N_2968);
or U5937 (N_5937,N_2875,N_3757);
nand U5938 (N_5938,N_2380,N_3309);
nand U5939 (N_5939,N_2489,N_2109);
nor U5940 (N_5940,N_3064,N_3691);
or U5941 (N_5941,N_2494,N_3340);
and U5942 (N_5942,N_3503,N_2865);
or U5943 (N_5943,N_2017,N_3134);
nand U5944 (N_5944,N_2847,N_3854);
nand U5945 (N_5945,N_2592,N_2579);
xnor U5946 (N_5946,N_2174,N_2984);
nand U5947 (N_5947,N_2279,N_3156);
or U5948 (N_5948,N_3071,N_2184);
or U5949 (N_5949,N_3190,N_3252);
xnor U5950 (N_5950,N_3279,N_2571);
and U5951 (N_5951,N_2522,N_3812);
nand U5952 (N_5952,N_2161,N_3508);
and U5953 (N_5953,N_2043,N_3778);
nor U5954 (N_5954,N_3149,N_2622);
and U5955 (N_5955,N_2226,N_2994);
and U5956 (N_5956,N_3378,N_2596);
or U5957 (N_5957,N_2036,N_3981);
nor U5958 (N_5958,N_2594,N_3331);
nand U5959 (N_5959,N_2733,N_2618);
and U5960 (N_5960,N_3754,N_2477);
or U5961 (N_5961,N_2222,N_2738);
nor U5962 (N_5962,N_3613,N_2385);
xor U5963 (N_5963,N_2107,N_2439);
and U5964 (N_5964,N_2633,N_3877);
and U5965 (N_5965,N_2599,N_2733);
and U5966 (N_5966,N_2977,N_3482);
or U5967 (N_5967,N_2478,N_2092);
nor U5968 (N_5968,N_2510,N_2755);
nand U5969 (N_5969,N_3194,N_3836);
nand U5970 (N_5970,N_3141,N_2849);
nor U5971 (N_5971,N_2164,N_2078);
and U5972 (N_5972,N_3957,N_3266);
and U5973 (N_5973,N_3190,N_2669);
nor U5974 (N_5974,N_3001,N_3688);
or U5975 (N_5975,N_3789,N_2641);
nor U5976 (N_5976,N_3505,N_3720);
or U5977 (N_5977,N_2120,N_3626);
nand U5978 (N_5978,N_2211,N_2495);
or U5979 (N_5979,N_3546,N_2829);
nor U5980 (N_5980,N_2743,N_2986);
nor U5981 (N_5981,N_3127,N_2583);
or U5982 (N_5982,N_2860,N_2957);
or U5983 (N_5983,N_3674,N_3747);
or U5984 (N_5984,N_2169,N_2658);
or U5985 (N_5985,N_2988,N_2444);
or U5986 (N_5986,N_3677,N_2559);
nand U5987 (N_5987,N_2120,N_2456);
nand U5988 (N_5988,N_3408,N_2357);
nor U5989 (N_5989,N_3640,N_3349);
nand U5990 (N_5990,N_2428,N_2423);
or U5991 (N_5991,N_2815,N_2573);
or U5992 (N_5992,N_2704,N_3625);
and U5993 (N_5993,N_2677,N_2868);
or U5994 (N_5994,N_2558,N_2601);
nand U5995 (N_5995,N_3322,N_2930);
and U5996 (N_5996,N_2556,N_3132);
or U5997 (N_5997,N_2860,N_2768);
and U5998 (N_5998,N_2468,N_2622);
nand U5999 (N_5999,N_2214,N_2470);
or U6000 (N_6000,N_5949,N_4923);
nand U6001 (N_6001,N_4638,N_5292);
xnor U6002 (N_6002,N_4349,N_5867);
or U6003 (N_6003,N_5023,N_4740);
or U6004 (N_6004,N_5696,N_4594);
xnor U6005 (N_6005,N_4366,N_4512);
nand U6006 (N_6006,N_5664,N_4924);
nor U6007 (N_6007,N_4336,N_4585);
nand U6008 (N_6008,N_4211,N_5250);
nand U6009 (N_6009,N_4816,N_5524);
or U6010 (N_6010,N_5813,N_4720);
nor U6011 (N_6011,N_5054,N_4610);
nand U6012 (N_6012,N_5434,N_4750);
or U6013 (N_6013,N_5122,N_4818);
nand U6014 (N_6014,N_4734,N_4363);
and U6015 (N_6015,N_4298,N_4866);
or U6016 (N_6016,N_4985,N_5565);
or U6017 (N_6017,N_4667,N_4094);
nand U6018 (N_6018,N_4814,N_5936);
nand U6019 (N_6019,N_5723,N_5608);
nor U6020 (N_6020,N_5454,N_5266);
nor U6021 (N_6021,N_5844,N_5814);
nor U6022 (N_6022,N_4346,N_5263);
nand U6023 (N_6023,N_5339,N_5010);
or U6024 (N_6024,N_4883,N_4412);
and U6025 (N_6025,N_4255,N_5417);
xor U6026 (N_6026,N_4119,N_5712);
and U6027 (N_6027,N_5981,N_5052);
and U6028 (N_6028,N_5077,N_5633);
nand U6029 (N_6029,N_4803,N_4464);
or U6030 (N_6030,N_4025,N_5420);
nor U6031 (N_6031,N_5815,N_4143);
and U6032 (N_6032,N_5610,N_5069);
or U6033 (N_6033,N_4632,N_5540);
nand U6034 (N_6034,N_4786,N_4327);
nor U6035 (N_6035,N_5729,N_4198);
nand U6036 (N_6036,N_5105,N_5297);
or U6037 (N_6037,N_4636,N_5687);
nor U6038 (N_6038,N_4314,N_5175);
and U6039 (N_6039,N_5967,N_5165);
xor U6040 (N_6040,N_4686,N_4468);
and U6041 (N_6041,N_4268,N_4582);
nor U6042 (N_6042,N_4491,N_5660);
or U6043 (N_6043,N_5973,N_4355);
or U6044 (N_6044,N_4142,N_4552);
nor U6045 (N_6045,N_5935,N_4890);
nor U6046 (N_6046,N_5634,N_4932);
and U6047 (N_6047,N_5317,N_4533);
nor U6048 (N_6048,N_4335,N_4205);
nor U6049 (N_6049,N_5380,N_4398);
nand U6050 (N_6050,N_5431,N_4093);
nand U6051 (N_6051,N_4972,N_4828);
nand U6052 (N_6052,N_4792,N_4567);
and U6053 (N_6053,N_5835,N_5549);
nor U6054 (N_6054,N_5133,N_4015);
nand U6055 (N_6055,N_4584,N_5327);
nand U6056 (N_6056,N_4337,N_4243);
or U6057 (N_6057,N_5436,N_4852);
or U6058 (N_6058,N_5385,N_5659);
or U6059 (N_6059,N_5360,N_4414);
and U6060 (N_6060,N_5612,N_4450);
nand U6061 (N_6061,N_4428,N_5253);
and U6062 (N_6062,N_4113,N_5242);
xnor U6063 (N_6063,N_4045,N_5167);
and U6064 (N_6064,N_4528,N_4879);
or U6065 (N_6065,N_4504,N_5346);
and U6066 (N_6066,N_5617,N_5087);
nor U6067 (N_6067,N_5068,N_4794);
and U6068 (N_6068,N_5162,N_4445);
nand U6069 (N_6069,N_5070,N_4189);
and U6070 (N_6070,N_5822,N_5238);
nand U6071 (N_6071,N_5650,N_4150);
nor U6072 (N_6072,N_4739,N_4315);
or U6073 (N_6073,N_5585,N_5232);
or U6074 (N_6074,N_5745,N_5990);
and U6075 (N_6075,N_4313,N_5163);
nand U6076 (N_6076,N_5316,N_5320);
and U6077 (N_6077,N_4531,N_5923);
and U6078 (N_6078,N_4571,N_5948);
nand U6079 (N_6079,N_4766,N_4643);
nor U6080 (N_6080,N_5917,N_5334);
nor U6081 (N_6081,N_4523,N_5830);
and U6082 (N_6082,N_4622,N_5697);
nand U6083 (N_6083,N_4703,N_5587);
nor U6084 (N_6084,N_4755,N_5440);
nor U6085 (N_6085,N_4707,N_5479);
and U6086 (N_6086,N_4410,N_4275);
nand U6087 (N_6087,N_4770,N_4303);
nor U6088 (N_6088,N_4185,N_4352);
and U6089 (N_6089,N_4112,N_5571);
nor U6090 (N_6090,N_5333,N_5839);
nand U6091 (N_6091,N_5210,N_4057);
or U6092 (N_6092,N_4694,N_4833);
or U6093 (N_6093,N_5314,N_5090);
or U6094 (N_6094,N_4449,N_5290);
nor U6095 (N_6095,N_5742,N_4058);
and U6096 (N_6096,N_4279,N_4272);
nand U6097 (N_6097,N_4863,N_4152);
nand U6098 (N_6098,N_5202,N_4161);
xor U6099 (N_6099,N_5455,N_5159);
and U6100 (N_6100,N_4043,N_4873);
nand U6101 (N_6101,N_4124,N_5776);
or U6102 (N_6102,N_4849,N_4305);
nand U6103 (N_6103,N_4100,N_5136);
or U6104 (N_6104,N_5195,N_5843);
or U6105 (N_6105,N_4541,N_4962);
nor U6106 (N_6106,N_5592,N_5944);
and U6107 (N_6107,N_4598,N_5880);
xnor U6108 (N_6108,N_4300,N_5583);
and U6109 (N_6109,N_5473,N_5925);
xnor U6110 (N_6110,N_5130,N_4477);
nand U6111 (N_6111,N_4576,N_4870);
or U6112 (N_6112,N_5625,N_5366);
nor U6113 (N_6113,N_4155,N_4730);
nand U6114 (N_6114,N_5688,N_5536);
or U6115 (N_6115,N_5627,N_5930);
nor U6116 (N_6116,N_4371,N_4467);
and U6117 (N_6117,N_4262,N_5858);
nand U6118 (N_6118,N_4714,N_5469);
and U6119 (N_6119,N_4490,N_5313);
nand U6120 (N_6120,N_5663,N_4999);
nand U6121 (N_6121,N_4178,N_5017);
nand U6122 (N_6122,N_5638,N_4601);
or U6123 (N_6123,N_4577,N_4283);
nand U6124 (N_6124,N_4173,N_5429);
or U6125 (N_6125,N_5555,N_4805);
or U6126 (N_6126,N_4399,N_4286);
nor U6127 (N_6127,N_5433,N_5151);
nor U6128 (N_6128,N_5271,N_4783);
nand U6129 (N_6129,N_5287,N_4560);
nor U6130 (N_6130,N_5272,N_5189);
nor U6131 (N_6131,N_4354,N_4735);
or U6132 (N_6132,N_5877,N_4245);
and U6133 (N_6133,N_5185,N_4778);
nor U6134 (N_6134,N_5889,N_5645);
nand U6135 (N_6135,N_5522,N_5075);
or U6136 (N_6136,N_5169,N_4758);
nand U6137 (N_6137,N_4745,N_5009);
and U6138 (N_6138,N_4613,N_5104);
or U6139 (N_6139,N_5997,N_4804);
and U6140 (N_6140,N_5037,N_4997);
or U6141 (N_6141,N_5894,N_4955);
nor U6142 (N_6142,N_5464,N_4511);
or U6143 (N_6143,N_4953,N_4098);
or U6144 (N_6144,N_4628,N_5040);
and U6145 (N_6145,N_5643,N_5827);
nand U6146 (N_6146,N_5355,N_4695);
nor U6147 (N_6147,N_4673,N_5057);
or U6148 (N_6148,N_4527,N_4159);
and U6149 (N_6149,N_5616,N_4407);
and U6150 (N_6150,N_4774,N_5763);
nor U6151 (N_6151,N_4421,N_4498);
nor U6152 (N_6152,N_4030,N_5506);
nand U6153 (N_6153,N_4950,N_5442);
or U6154 (N_6154,N_4789,N_5305);
nor U6155 (N_6155,N_4326,N_5875);
and U6156 (N_6156,N_5280,N_4242);
nand U6157 (N_6157,N_5968,N_5324);
nand U6158 (N_6158,N_4811,N_5237);
nand U6159 (N_6159,N_4370,N_4761);
or U6160 (N_6160,N_4517,N_5012);
or U6161 (N_6161,N_5512,N_5890);
nor U6162 (N_6162,N_5582,N_5100);
or U6163 (N_6163,N_4312,N_5132);
and U6164 (N_6164,N_4682,N_5032);
or U6165 (N_6165,N_5779,N_5294);
nand U6166 (N_6166,N_5979,N_4182);
or U6167 (N_6167,N_4088,N_4543);
xor U6168 (N_6168,N_4223,N_5603);
nand U6169 (N_6169,N_4221,N_4549);
nand U6170 (N_6170,N_5938,N_4338);
and U6171 (N_6171,N_4765,N_5517);
nand U6172 (N_6172,N_4383,N_4961);
or U6173 (N_6173,N_5533,N_5089);
nand U6174 (N_6174,N_5093,N_4318);
xor U6175 (N_6175,N_4539,N_4797);
nor U6176 (N_6176,N_4017,N_4146);
and U6177 (N_6177,N_4499,N_5359);
or U6178 (N_6178,N_5124,N_4201);
and U6179 (N_6179,N_5353,N_4603);
nor U6180 (N_6180,N_5515,N_4053);
nand U6181 (N_6181,N_4590,N_5138);
or U6182 (N_6182,N_5443,N_4718);
nor U6183 (N_6183,N_5092,N_5193);
nor U6184 (N_6184,N_4855,N_4966);
nor U6185 (N_6185,N_5128,N_4894);
nor U6186 (N_6186,N_4080,N_5183);
and U6187 (N_6187,N_5681,N_4526);
or U6188 (N_6188,N_5422,N_5720);
and U6189 (N_6189,N_5080,N_4202);
or U6190 (N_6190,N_5363,N_5846);
nor U6191 (N_6191,N_5811,N_4965);
or U6192 (N_6192,N_4438,N_4246);
nand U6193 (N_6193,N_4538,N_5800);
nor U6194 (N_6194,N_5399,N_5851);
nand U6195 (N_6195,N_5841,N_5600);
and U6196 (N_6196,N_5866,N_4705);
and U6197 (N_6197,N_4031,N_5834);
or U6198 (N_6198,N_4501,N_5386);
nor U6199 (N_6199,N_5229,N_4458);
nor U6200 (N_6200,N_5435,N_4285);
nor U6201 (N_6201,N_4505,N_5766);
or U6202 (N_6202,N_4029,N_4977);
nor U6203 (N_6203,N_4630,N_4476);
or U6204 (N_6204,N_4391,N_4564);
nor U6205 (N_6205,N_5771,N_4889);
nor U6206 (N_6206,N_5821,N_5146);
and U6207 (N_6207,N_4406,N_4558);
and U6208 (N_6208,N_5476,N_5387);
nor U6209 (N_6209,N_5013,N_5496);
and U6210 (N_6210,N_5283,N_5853);
or U6211 (N_6211,N_5022,N_4036);
nor U6212 (N_6212,N_5807,N_5437);
and U6213 (N_6213,N_4068,N_4236);
or U6214 (N_6214,N_4599,N_4680);
nand U6215 (N_6215,N_5511,N_4258);
nand U6216 (N_6216,N_4954,N_5769);
nand U6217 (N_6217,N_5942,N_5629);
nor U6218 (N_6218,N_5135,N_4812);
nor U6219 (N_6219,N_4915,N_5791);
nor U6220 (N_6220,N_4126,N_5596);
xor U6221 (N_6221,N_4583,N_5717);
nor U6222 (N_6222,N_4465,N_4308);
nor U6223 (N_6223,N_4557,N_5589);
nor U6224 (N_6224,N_4665,N_5118);
and U6225 (N_6225,N_5929,N_4838);
nor U6226 (N_6226,N_4649,N_5256);
nand U6227 (N_6227,N_4678,N_5502);
and U6228 (N_6228,N_5934,N_5076);
nand U6229 (N_6229,N_5505,N_4779);
nor U6230 (N_6230,N_4569,N_5641);
nor U6231 (N_6231,N_5099,N_4016);
or U6232 (N_6232,N_4076,N_4012);
nand U6233 (N_6233,N_5341,N_4799);
and U6234 (N_6234,N_5624,N_5554);
nor U6235 (N_6235,N_4518,N_4469);
nand U6236 (N_6236,N_5172,N_4418);
or U6237 (N_6237,N_4933,N_5495);
and U6238 (N_6238,N_5457,N_5028);
nand U6239 (N_6239,N_5489,N_5622);
nor U6240 (N_6240,N_5969,N_4020);
nor U6241 (N_6241,N_5906,N_4168);
nor U6242 (N_6242,N_4282,N_5321);
nand U6243 (N_6243,N_5686,N_4843);
xnor U6244 (N_6244,N_4166,N_4460);
or U6245 (N_6245,N_4046,N_4815);
and U6246 (N_6246,N_4690,N_4145);
nor U6247 (N_6247,N_5326,N_4026);
xor U6248 (N_6248,N_5231,N_4897);
nand U6249 (N_6249,N_5330,N_4484);
xor U6250 (N_6250,N_4573,N_4840);
nor U6251 (N_6251,N_4149,N_4942);
or U6252 (N_6252,N_5390,N_5078);
or U6253 (N_6253,N_5221,N_5155);
nor U6254 (N_6254,N_5953,N_4893);
and U6255 (N_6255,N_4929,N_5874);
nor U6256 (N_6256,N_4325,N_5996);
and U6257 (N_6257,N_5142,N_4916);
nor U6258 (N_6258,N_4782,N_4704);
and U6259 (N_6259,N_5668,N_4139);
or U6260 (N_6260,N_5993,N_5567);
and U6261 (N_6261,N_5863,N_5816);
nand U6262 (N_6262,N_5394,N_4448);
nand U6263 (N_6263,N_5050,N_5995);
nand U6264 (N_6264,N_5262,N_5094);
nor U6265 (N_6265,N_4944,N_5736);
and U6266 (N_6266,N_5989,N_5180);
and U6267 (N_6267,N_4565,N_4579);
nor U6268 (N_6268,N_4963,N_4519);
and U6269 (N_6269,N_5487,N_4381);
xor U6270 (N_6270,N_5557,N_4620);
nand U6271 (N_6271,N_4751,N_5873);
nand U6272 (N_6272,N_5369,N_5726);
nor U6273 (N_6273,N_5086,N_5019);
or U6274 (N_6274,N_4022,N_4669);
and U6275 (N_6275,N_5601,N_5750);
and U6276 (N_6276,N_5905,N_4127);
nor U6277 (N_6277,N_5558,N_5613);
and U6278 (N_6278,N_5458,N_4713);
nand U6279 (N_6279,N_4172,N_5992);
or U6280 (N_6280,N_5245,N_4290);
and U6281 (N_6281,N_4600,N_5885);
nor U6282 (N_6282,N_5240,N_5868);
and U6283 (N_6283,N_5578,N_4050);
or U6284 (N_6284,N_5514,N_4203);
xor U6285 (N_6285,N_5538,N_5082);
and U6286 (N_6286,N_5260,N_4712);
nand U6287 (N_6287,N_4230,N_4960);
nor U6288 (N_6288,N_4374,N_4247);
xnor U6289 (N_6289,N_5900,N_5892);
and U6290 (N_6290,N_5637,N_4359);
or U6291 (N_6291,N_4388,N_4070);
and U6292 (N_6292,N_5038,N_4589);
nand U6293 (N_6293,N_4362,N_4864);
nor U6294 (N_6294,N_5907,N_4895);
xor U6295 (N_6295,N_4027,N_4534);
nor U6296 (N_6296,N_5849,N_5295);
or U6297 (N_6297,N_5404,N_5715);
or U6298 (N_6298,N_5241,N_4235);
and U6299 (N_6299,N_5154,N_5225);
nor U6300 (N_6300,N_4905,N_4231);
nor U6301 (N_6301,N_4981,N_5071);
nand U6302 (N_6302,N_5005,N_5338);
nor U6303 (N_6303,N_4424,N_5590);
nand U6304 (N_6304,N_4776,N_5854);
nand U6305 (N_6305,N_5658,N_5466);
or U6306 (N_6306,N_4400,N_4967);
nor U6307 (N_6307,N_5510,N_5739);
or U6308 (N_6308,N_5552,N_5083);
and U6309 (N_6309,N_5484,N_5584);
nor U6310 (N_6310,N_4208,N_4241);
nor U6311 (N_6311,N_4191,N_4914);
and U6312 (N_6312,N_4748,N_5129);
or U6313 (N_6313,N_4545,N_4763);
nand U6314 (N_6314,N_4684,N_5065);
and U6315 (N_6315,N_5423,N_4976);
nand U6316 (N_6316,N_4200,N_4105);
nand U6317 (N_6317,N_5051,N_4696);
or U6318 (N_6318,N_4461,N_5301);
nor U6319 (N_6319,N_5192,N_5449);
xnor U6320 (N_6320,N_5203,N_5621);
and U6321 (N_6321,N_4618,N_5724);
or U6322 (N_6322,N_4555,N_4801);
and U6323 (N_6323,N_5539,N_4456);
and U6324 (N_6324,N_4948,N_5409);
and U6325 (N_6325,N_4034,N_4280);
nand U6326 (N_6326,N_5456,N_4664);
nor U6327 (N_6327,N_5020,N_4825);
nand U6328 (N_6328,N_4524,N_4463);
and U6329 (N_6329,N_5413,N_4451);
nor U6330 (N_6330,N_4767,N_5679);
nand U6331 (N_6331,N_4377,N_4441);
nor U6332 (N_6332,N_4394,N_4344);
nand U6333 (N_6333,N_4423,N_4532);
nor U6334 (N_6334,N_4685,N_4369);
or U6335 (N_6335,N_4073,N_5323);
and U6336 (N_6336,N_5218,N_5752);
and U6337 (N_6337,N_4250,N_4546);
nor U6338 (N_6338,N_5345,N_5852);
nand U6339 (N_6339,N_5626,N_5415);
nand U6340 (N_6340,N_5230,N_4257);
nand U6341 (N_6341,N_5783,N_5680);
nor U6342 (N_6342,N_5756,N_5566);
nand U6343 (N_6343,N_5462,N_5795);
nor U6344 (N_6344,N_4074,N_4040);
nand U6345 (N_6345,N_4844,N_4485);
or U6346 (N_6346,N_5117,N_5212);
and U6347 (N_6347,N_5403,N_4741);
nand U6348 (N_6348,N_4443,N_5699);
and U6349 (N_6349,N_4514,N_4837);
nand U6350 (N_6350,N_4648,N_4486);
xnor U6351 (N_6351,N_5528,N_5044);
and U6352 (N_6352,N_4970,N_5447);
or U6353 (N_6353,N_4084,N_4727);
nor U6354 (N_6354,N_5694,N_5899);
nor U6355 (N_6355,N_4771,N_4578);
and U6356 (N_6356,N_4856,N_4540);
and U6357 (N_6357,N_5101,N_4429);
and U6358 (N_6358,N_4404,N_4506);
and U6359 (N_6359,N_5053,N_5248);
and U6360 (N_6360,N_4850,N_5609);
or U6361 (N_6361,N_4591,N_5375);
nor U6362 (N_6362,N_4516,N_5770);
and U6363 (N_6363,N_4008,N_4759);
nor U6364 (N_6364,N_4787,N_4984);
nor U6365 (N_6365,N_5432,N_4835);
xor U6366 (N_6366,N_5312,N_4321);
nor U6367 (N_6367,N_5598,N_4442);
and U6368 (N_6368,N_5526,N_5418);
nand U6369 (N_6369,N_4785,N_5733);
and U6370 (N_6370,N_4273,N_4368);
and U6371 (N_6371,N_5812,N_4522);
nand U6372 (N_6372,N_4570,N_5111);
and U6373 (N_6373,N_4973,N_4858);
nand U6374 (N_6374,N_5937,N_5714);
and U6375 (N_6375,N_5430,N_4439);
xor U6376 (N_6376,N_5214,N_4219);
or U6377 (N_6377,N_5490,N_5414);
and U6378 (N_6378,N_5755,N_4360);
nand U6379 (N_6379,N_4508,N_4722);
nor U6380 (N_6380,N_4662,N_4329);
or U6381 (N_6381,N_5818,N_4481);
nor U6382 (N_6382,N_5709,N_5467);
and U6383 (N_6383,N_5368,N_5887);
or U6384 (N_6384,N_5309,N_4306);
and U6385 (N_6385,N_4064,N_5927);
nand U6386 (N_6386,N_5021,N_4206);
nor U6387 (N_6387,N_4331,N_5491);
or U6388 (N_6388,N_4762,N_5778);
nor U6389 (N_6389,N_4715,N_5097);
xor U6390 (N_6390,N_4256,N_4559);
nand U6391 (N_6391,N_4611,N_5140);
and U6392 (N_6392,N_5329,N_4433);
or U6393 (N_6393,N_5194,N_5693);
nor U6394 (N_6394,N_4121,N_5182);
or U6395 (N_6395,N_4033,N_4887);
nor U6396 (N_6396,N_5173,N_4302);
and U6397 (N_6397,N_4507,N_4938);
or U6398 (N_6398,N_4078,N_5731);
and U6399 (N_6399,N_4666,N_5149);
and U6400 (N_6400,N_5775,N_5499);
nand U6401 (N_6401,N_5888,N_5014);
nor U6402 (N_6402,N_5980,N_4220);
and U6403 (N_6403,N_5235,N_4091);
nand U6404 (N_6404,N_5655,N_5452);
and U6405 (N_6405,N_4723,N_4260);
nor U6406 (N_6406,N_5131,N_5107);
or U6407 (N_6407,N_4470,N_4642);
or U6408 (N_6408,N_5274,N_5026);
and U6409 (N_6409,N_4568,N_5342);
or U6410 (N_6410,N_4188,N_4876);
nor U6411 (N_6411,N_5036,N_4634);
or U6412 (N_6412,N_4244,N_5817);
and U6413 (N_6413,N_4710,N_5063);
or U6414 (N_6414,N_4077,N_5673);
nor U6415 (N_6415,N_5448,N_4154);
and U6416 (N_6416,N_5809,N_4446);
nor U6417 (N_6417,N_4291,N_5691);
nor U6418 (N_6418,N_4083,N_4288);
and U6419 (N_6419,N_5216,N_4348);
and U6420 (N_6420,N_5698,N_5190);
xnor U6421 (N_6421,N_4365,N_5033);
nor U6422 (N_6422,N_5982,N_5605);
and U6423 (N_6423,N_4553,N_4865);
and U6424 (N_6424,N_4807,N_5573);
and U6425 (N_6425,N_5170,N_5760);
and U6426 (N_6426,N_4940,N_4996);
or U6427 (N_6427,N_5757,N_5544);
and U6428 (N_6428,N_4798,N_4906);
nor U6429 (N_6429,N_4660,N_4222);
and U6430 (N_6430,N_5630,N_4911);
and U6431 (N_6431,N_5667,N_4688);
and U6432 (N_6432,N_4322,N_5672);
and U6433 (N_6433,N_5962,N_5966);
nor U6434 (N_6434,N_5397,N_4270);
nand U6435 (N_6435,N_5897,N_4904);
nor U6436 (N_6436,N_4081,N_5184);
or U6437 (N_6437,N_5494,N_4683);
nand U6438 (N_6438,N_4772,N_5029);
or U6439 (N_6439,N_5347,N_4174);
nor U6440 (N_6440,N_5181,N_4655);
nor U6441 (N_6441,N_4644,N_5870);
and U6442 (N_6442,N_4003,N_4005);
or U6443 (N_6443,N_4276,N_4658);
or U6444 (N_6444,N_4503,N_4744);
nor U6445 (N_6445,N_5396,N_4006);
or U6446 (N_6446,N_5306,N_4132);
or U6447 (N_6447,N_4123,N_5407);
and U6448 (N_6448,N_4452,N_5904);
nand U6449 (N_6449,N_4878,N_5903);
nand U6450 (N_6450,N_4651,N_5956);
and U6451 (N_6451,N_5239,N_5265);
and U6452 (N_6452,N_4425,N_4002);
nand U6453 (N_6453,N_4580,N_4547);
nor U6454 (N_6454,N_4676,N_4378);
or U6455 (N_6455,N_5902,N_5060);
nand U6456 (N_6456,N_5516,N_5761);
and U6457 (N_6457,N_5500,N_4147);
nor U6458 (N_6458,N_5459,N_4278);
and U6459 (N_6459,N_5940,N_4156);
or U6460 (N_6460,N_5651,N_4925);
and U6461 (N_6461,N_5521,N_4769);
or U6462 (N_6462,N_4809,N_5706);
or U6463 (N_6463,N_4384,N_4606);
and U6464 (N_6464,N_4459,N_5357);
nor U6465 (N_6465,N_5998,N_4581);
nand U6466 (N_6466,N_5226,N_5048);
or U6467 (N_6467,N_4373,N_4431);
nand U6468 (N_6468,N_4125,N_5493);
and U6469 (N_6469,N_5416,N_4054);
nand U6470 (N_6470,N_5842,N_5523);
nand U6471 (N_6471,N_4753,N_4982);
nand U6472 (N_6472,N_5143,N_4509);
and U6473 (N_6473,N_5134,N_4138);
nor U6474 (N_6474,N_4047,N_5653);
or U6475 (N_6475,N_5606,N_5782);
and U6476 (N_6476,N_5802,N_4515);
nand U6477 (N_6477,N_5288,N_5919);
nor U6478 (N_6478,N_4310,N_5300);
nand U6479 (N_6479,N_5319,N_4204);
and U6480 (N_6480,N_5110,N_5371);
or U6481 (N_6481,N_5144,N_4708);
or U6482 (N_6482,N_5258,N_4382);
and U6483 (N_6483,N_5145,N_4781);
nand U6484 (N_6484,N_4263,N_4214);
nor U6485 (N_6485,N_4989,N_5788);
and U6486 (N_6486,N_5402,N_5308);
nor U6487 (N_6487,N_4148,N_5468);
nand U6488 (N_6488,N_5632,N_5377);
or U6489 (N_6489,N_5168,N_4724);
nor U6490 (N_6490,N_4072,N_4042);
and U6491 (N_6491,N_5577,N_5351);
or U6492 (N_6492,N_4875,N_4808);
nor U6493 (N_6493,N_5648,N_4930);
and U6494 (N_6494,N_4921,N_4760);
nor U6495 (N_6495,N_4011,N_4817);
and U6496 (N_6496,N_4861,N_5007);
and U6497 (N_6497,N_4831,N_5450);
nand U6498 (N_6498,N_5108,N_5615);
nand U6499 (N_6499,N_5400,N_5518);
and U6500 (N_6500,N_5066,N_5166);
nand U6501 (N_6501,N_5964,N_4544);
or U6502 (N_6502,N_4375,N_5391);
and U6503 (N_6503,N_5527,N_5508);
xnor U6504 (N_6504,N_5411,N_4419);
and U6505 (N_6505,N_5498,N_4862);
and U6506 (N_6506,N_5639,N_4328);
or U6507 (N_6507,N_5958,N_5121);
nor U6508 (N_6508,N_4248,N_4586);
nand U6509 (N_6509,N_5164,N_5798);
nand U6510 (N_6510,N_5910,N_5525);
or U6511 (N_6511,N_4343,N_4502);
nor U6512 (N_6512,N_4992,N_5799);
or U6513 (N_6513,N_4417,N_5674);
and U6514 (N_6514,N_5829,N_5365);
or U6515 (N_6515,N_4457,N_4111);
and U6516 (N_6516,N_5716,N_5545);
nor U6517 (N_6517,N_4434,N_5753);
nand U6518 (N_6518,N_5158,N_5692);
xnor U6519 (N_6519,N_5532,N_4788);
and U6520 (N_6520,N_4180,N_4971);
xor U6521 (N_6521,N_5025,N_4289);
nand U6522 (N_6522,N_5677,N_4239);
nor U6523 (N_6523,N_4192,N_4332);
and U6524 (N_6524,N_5881,N_5808);
and U6525 (N_6525,N_4937,N_4654);
nor U6526 (N_6526,N_4525,N_5971);
or U6527 (N_6527,N_5862,N_4115);
nand U6528 (N_6528,N_4884,N_4689);
nor U6529 (N_6529,N_4489,N_4846);
and U6530 (N_6530,N_5485,N_4086);
or U6531 (N_6531,N_4311,N_5217);
or U6532 (N_6532,N_4874,N_5056);
and U6533 (N_6533,N_4635,N_5580);
nand U6534 (N_6534,N_4736,N_4646);
nor U6535 (N_6535,N_4281,N_4389);
nor U6536 (N_6536,N_4561,N_4096);
and U6537 (N_6537,N_4823,N_4109);
or U6538 (N_6538,N_5482,N_5654);
nand U6539 (N_6539,N_5568,N_4408);
nor U6540 (N_6540,N_5497,N_5825);
or U6541 (N_6541,N_4251,N_4677);
nor U6542 (N_6542,N_5656,N_5067);
and U6543 (N_6543,N_4627,N_5547);
nor U6544 (N_6544,N_5901,N_5299);
and U6545 (N_6545,N_4550,N_4176);
and U6546 (N_6546,N_4347,N_4537);
nand U6547 (N_6547,N_4304,N_4877);
or U6548 (N_6548,N_4854,N_5804);
or U6549 (N_6549,N_4324,N_4520);
and U6550 (N_6550,N_5261,N_5991);
or U6551 (N_6551,N_5307,N_5379);
and U6552 (N_6552,N_4212,N_5161);
nand U6553 (N_6553,N_5188,N_5570);
or U6554 (N_6554,N_5665,N_4892);
nand U6555 (N_6555,N_5354,N_5551);
and U6556 (N_6556,N_5529,N_5304);
nand U6557 (N_6557,N_5085,N_4746);
and U6558 (N_6558,N_5471,N_5220);
and U6559 (N_6559,N_5279,N_5932);
or U6560 (N_6560,N_4896,N_5833);
nor U6561 (N_6561,N_4140,N_4116);
nor U6562 (N_6562,N_5303,N_5201);
or U6563 (N_6563,N_5572,N_4657);
nand U6564 (N_6564,N_4396,N_5254);
nand U6565 (N_6565,N_5574,N_4194);
nor U6566 (N_6566,N_5480,N_4385);
or U6567 (N_6567,N_5157,N_4001);
or U6568 (N_6568,N_5628,N_5553);
nand U6569 (N_6569,N_4482,N_4021);
nor U6570 (N_6570,N_4562,N_5503);
or U6571 (N_6571,N_5859,N_5747);
nand U6572 (N_6572,N_5461,N_4796);
nor U6573 (N_6573,N_5780,N_5920);
and U6574 (N_6574,N_4768,N_4240);
and U6575 (N_6575,N_5797,N_5318);
and U6576 (N_6576,N_4913,N_5777);
nor U6577 (N_6577,N_4044,N_4475);
nand U6578 (N_6578,N_5340,N_4625);
and U6579 (N_6579,N_4640,N_4701);
and U6580 (N_6580,N_4227,N_4233);
or U6581 (N_6581,N_5749,N_4157);
nand U6582 (N_6582,N_5618,N_4259);
nand U6583 (N_6583,N_5611,N_5125);
nand U6584 (N_6584,N_5762,N_5267);
nand U6585 (N_6585,N_4958,N_4092);
or U6586 (N_6586,N_4721,N_4826);
nand U6587 (N_6587,N_4616,N_4162);
nand U6588 (N_6588,N_4415,N_5174);
nand U6589 (N_6589,N_4108,N_4728);
and U6590 (N_6590,N_4411,N_5865);
and U6591 (N_6591,N_5884,N_5358);
nand U6592 (N_6592,N_4069,N_4409);
or U6593 (N_6593,N_5914,N_5999);
nor U6594 (N_6594,N_4014,N_5120);
nand U6595 (N_6595,N_4738,N_5509);
nand U6596 (N_6596,N_4656,N_4061);
nand U6597 (N_6597,N_5564,N_5882);
nor U6598 (N_6598,N_4493,N_4401);
and U6599 (N_6599,N_4402,N_5176);
nor U6600 (N_6600,N_4853,N_5039);
and U6601 (N_6601,N_5640,N_5200);
nand U6602 (N_6602,N_5095,N_5002);
nand U6603 (N_6603,N_4888,N_4842);
nand U6604 (N_6604,N_4462,N_4133);
nand U6605 (N_6605,N_5972,N_4186);
and U6606 (N_6606,N_4294,N_5569);
and U6607 (N_6607,N_4709,N_4060);
nor U6608 (N_6608,N_5088,N_5614);
or U6609 (N_6609,N_4216,N_4117);
or U6610 (N_6610,N_5513,N_4988);
and U6611 (N_6611,N_4454,N_5119);
and U6612 (N_6612,N_4548,N_5361);
or U6613 (N_6613,N_4187,N_4829);
or U6614 (N_6614,N_5302,N_4979);
and U6615 (N_6615,N_5792,N_4190);
nand U6616 (N_6616,N_5344,N_5541);
or U6617 (N_6617,N_4647,N_5244);
nand U6618 (N_6618,N_4037,N_5198);
nand U6619 (N_6619,N_4492,N_4183);
and U6620 (N_6620,N_4292,N_5861);
or U6621 (N_6621,N_5255,N_4872);
or U6622 (N_6622,N_4010,N_4293);
nor U6623 (N_6623,N_4134,N_4158);
and U6624 (N_6624,N_5918,N_5043);
nor U6625 (N_6625,N_4177,N_5737);
and U6626 (N_6626,N_4089,N_5259);
and U6627 (N_6627,N_4049,N_4624);
nor U6628 (N_6628,N_5913,N_5349);
nand U6629 (N_6629,N_5042,N_4536);
and U6630 (N_6630,N_5719,N_4128);
nand U6631 (N_6631,N_5635,N_4716);
nor U6632 (N_6632,N_4102,N_4488);
nand U6633 (N_6633,N_4943,N_4777);
nand U6634 (N_6634,N_4024,N_5983);
and U6635 (N_6635,N_4065,N_5951);
nor U6636 (N_6636,N_5072,N_5520);
or U6637 (N_6637,N_5768,N_5024);
xor U6638 (N_6638,N_4902,N_4672);
nor U6639 (N_6639,N_4706,N_5560);
and U6640 (N_6640,N_5593,N_5049);
nand U6641 (N_6641,N_5223,N_5591);
nor U6642 (N_6642,N_5335,N_4051);
nand U6643 (N_6643,N_5337,N_5790);
nor U6644 (N_6644,N_5909,N_5343);
or U6645 (N_6645,N_5247,N_4009);
and U6646 (N_6646,N_5784,N_4614);
or U6647 (N_6647,N_4164,N_5233);
or U6648 (N_6648,N_4048,N_4032);
nand U6649 (N_6649,N_5678,N_5793);
nor U6650 (N_6650,N_5296,N_5001);
or U6651 (N_6651,N_5045,N_4144);
nand U6652 (N_6652,N_4731,N_4494);
or U6653 (N_6653,N_4479,N_4309);
and U6654 (N_6654,N_4195,N_5926);
or U6655 (N_6655,N_5789,N_4103);
nor U6656 (N_6656,N_4857,N_4217);
or U6657 (N_6657,N_4612,N_4197);
nor U6658 (N_6658,N_4700,N_5109);
or U6659 (N_6659,N_4593,N_4668);
nor U6660 (N_6660,N_4104,N_5563);
nand U6661 (N_6661,N_5098,N_4775);
nand U6662 (N_6662,N_4320,N_4733);
or U6663 (N_6663,N_5126,N_5507);
nor U6664 (N_6664,N_5389,N_4453);
or U6665 (N_6665,N_5199,N_4478);
xnor U6666 (N_6666,N_4041,N_5102);
nand U6667 (N_6667,N_5061,N_5475);
nor U6668 (N_6668,N_5684,N_4427);
or U6669 (N_6669,N_4341,N_4588);
nand U6670 (N_6670,N_5939,N_4968);
or U6671 (N_6671,N_5631,N_4237);
xor U6672 (N_6672,N_5015,N_4592);
nor U6673 (N_6673,N_4252,N_4171);
nor U6674 (N_6674,N_4471,N_4670);
nor U6675 (N_6675,N_4296,N_5732);
nor U6676 (N_6676,N_4082,N_4379);
nand U6677 (N_6677,N_4107,N_5059);
or U6678 (N_6678,N_5249,N_4087);
or U6679 (N_6679,N_4681,N_4563);
nand U6680 (N_6680,N_4860,N_5224);
or U6681 (N_6681,N_4004,N_5311);
nor U6682 (N_6682,N_4234,N_4000);
and U6683 (N_6683,N_4307,N_5446);
or U6684 (N_6684,N_4742,N_4097);
or U6685 (N_6685,N_5362,N_4274);
nor U6686 (N_6686,N_4629,N_5838);
nor U6687 (N_6687,N_5211,N_4075);
xnor U6688 (N_6688,N_5711,N_4551);
nand U6689 (N_6689,N_4287,N_4110);
and U6690 (N_6690,N_4405,N_4218);
nand U6691 (N_6691,N_4934,N_5826);
or U6692 (N_6692,N_4213,N_5227);
and U6693 (N_6693,N_4645,N_4974);
and U6694 (N_6694,N_4927,N_5604);
nand U6695 (N_6695,N_4135,N_5278);
and U6696 (N_6696,N_4085,N_5445);
nor U6697 (N_6697,N_5550,N_4342);
nand U6698 (N_6698,N_4416,N_5011);
and U6699 (N_6699,N_4907,N_5410);
nor U6700 (N_6700,N_4743,N_5581);
or U6701 (N_6701,N_4153,N_5519);
or U6702 (N_6702,N_5405,N_5504);
or U6703 (N_6703,N_5251,N_4995);
nor U6704 (N_6704,N_4639,N_4918);
nand U6705 (N_6705,N_4754,N_5856);
nor U6706 (N_6706,N_5928,N_4993);
or U6707 (N_6707,N_4356,N_4726);
and U6708 (N_6708,N_5425,N_5730);
and U6709 (N_6709,N_4926,N_5392);
xnor U6710 (N_6710,N_5246,N_5728);
or U6711 (N_6711,N_4380,N_5786);
and U6712 (N_6712,N_5352,N_5428);
and U6713 (N_6713,N_5035,N_5735);
nand U6714 (N_6714,N_4299,N_4729);
nand U6715 (N_6715,N_4019,N_5754);
nor U6716 (N_6716,N_4834,N_4095);
nor U6717 (N_6717,N_4899,N_4529);
nor U6718 (N_6718,N_4998,N_4964);
or U6719 (N_6719,N_4238,N_4617);
nand U6720 (N_6720,N_5963,N_4390);
nor U6721 (N_6721,N_5898,N_5847);
nor U6722 (N_6722,N_5062,N_4602);
nor U6723 (N_6723,N_5741,N_4986);
nand U6724 (N_6724,N_4059,N_5207);
nor U6725 (N_6725,N_4752,N_4891);
or U6726 (N_6726,N_4910,N_4773);
nor U6727 (N_6727,N_4056,N_5556);
and U6728 (N_6728,N_5767,N_5041);
nand U6729 (N_6729,N_4692,N_4170);
nor U6730 (N_6730,N_5855,N_5374);
nor U6731 (N_6731,N_5016,N_4900);
or U6732 (N_6732,N_5921,N_4351);
nand U6733 (N_6733,N_5662,N_5781);
or U6734 (N_6734,N_4055,N_4780);
nor U6735 (N_6735,N_4496,N_5562);
nand U6736 (N_6736,N_5602,N_4440);
nor U6737 (N_6737,N_4444,N_5501);
nand U6738 (N_6738,N_5003,N_4137);
nand U6739 (N_6739,N_4334,N_4122);
xnor U6740 (N_6740,N_5976,N_5535);
nand U6741 (N_6741,N_4663,N_4226);
nor U6742 (N_6742,N_4922,N_4487);
nand U6743 (N_6743,N_5772,N_4939);
nand U6744 (N_6744,N_5367,N_5738);
nor U6745 (N_6745,N_4028,N_4269);
nand U6746 (N_6746,N_5718,N_5922);
nor U6747 (N_6747,N_4264,N_5419);
and U6748 (N_6748,N_5298,N_4802);
or U6749 (N_6749,N_5666,N_4413);
and U6750 (N_6750,N_5727,N_5336);
nand U6751 (N_6751,N_5810,N_4671);
nor U6752 (N_6752,N_4868,N_4983);
nand U6753 (N_6753,N_5824,N_4886);
or U6754 (N_6754,N_5671,N_4013);
nor U6755 (N_6755,N_5213,N_4130);
and U6756 (N_6756,N_5426,N_5806);
nand U6757 (N_6757,N_5096,N_4295);
nand U6758 (N_6758,N_4497,N_5141);
nand U6759 (N_6759,N_4756,N_4039);
and U6760 (N_6760,N_5383,N_5328);
nor U6761 (N_6761,N_4691,N_5222);
nand U6762 (N_6762,N_5912,N_4062);
or U6763 (N_6763,N_5764,N_4353);
nand U6764 (N_6764,N_5831,N_4791);
and U6765 (N_6765,N_4254,N_5986);
or U6766 (N_6766,N_5488,N_4959);
or U6767 (N_6767,N_4106,N_4167);
nand U6768 (N_6768,N_5965,N_4575);
and U6769 (N_6769,N_5370,N_5113);
and U6770 (N_6770,N_5695,N_4990);
and U6771 (N_6771,N_4882,N_5289);
and U6772 (N_6772,N_4480,N_4810);
nand U6773 (N_6773,N_4129,N_5945);
nor U6774 (N_6774,N_4023,N_5470);
nand U6775 (N_6775,N_4623,N_4376);
nor U6776 (N_6776,N_5620,N_5486);
or U6777 (N_6777,N_4193,N_5438);
or U6778 (N_6778,N_4845,N_5751);
or U6779 (N_6779,N_5408,N_5127);
or U6780 (N_6780,N_4483,N_5441);
and U6781 (N_6781,N_4038,N_4908);
and U6782 (N_6782,N_4793,N_5576);
and U6783 (N_6783,N_5046,N_5178);
or U6784 (N_6784,N_4447,N_4626);
nand U6785 (N_6785,N_5186,N_5690);
nor U6786 (N_6786,N_4909,N_5058);
and U6787 (N_6787,N_5748,N_5710);
nor U6788 (N_6788,N_4466,N_5725);
and U6789 (N_6789,N_5322,N_5594);
nand U6790 (N_6790,N_4747,N_4165);
or U6791 (N_6791,N_5924,N_5084);
or U6792 (N_6792,N_4956,N_5208);
nor U6793 (N_6793,N_5785,N_5243);
and U6794 (N_6794,N_4795,N_5950);
or U6795 (N_6795,N_5008,N_4637);
nor U6796 (N_6796,N_4836,N_5878);
or U6797 (N_6797,N_5682,N_5378);
and U6798 (N_6798,N_5115,N_5137);
and U6799 (N_6799,N_5836,N_4757);
and U6800 (N_6800,N_5376,N_4392);
nand U6801 (N_6801,N_5543,N_5876);
or U6802 (N_6802,N_5286,N_5970);
nor U6803 (N_6803,N_5147,N_4697);
nor U6804 (N_6804,N_4358,N_5091);
and U6805 (N_6805,N_4530,N_5801);
nor U6806 (N_6806,N_5743,N_4319);
or U6807 (N_6807,N_5740,N_5276);
or U6808 (N_6808,N_5477,N_5364);
and U6809 (N_6809,N_5759,N_4717);
or U6810 (N_6810,N_4437,N_4253);
or U6811 (N_6811,N_5444,N_5988);
and U6812 (N_6812,N_4957,N_4574);
xor U6813 (N_6813,N_4395,N_5474);
or U6814 (N_6814,N_5384,N_4928);
nor U6815 (N_6815,N_4066,N_4869);
or U6816 (N_6816,N_5139,N_4572);
nor U6817 (N_6817,N_5206,N_4650);
and U6818 (N_6818,N_5463,N_5961);
nor U6819 (N_6819,N_5685,N_5828);
or U6820 (N_6820,N_5708,N_5081);
nor U6821 (N_6821,N_5805,N_5196);
nand U6822 (N_6822,N_5160,N_5879);
nor U6823 (N_6823,N_4587,N_4737);
or U6824 (N_6824,N_5412,N_4403);
nand U6825 (N_6825,N_5534,N_4951);
nand U6826 (N_6826,N_4513,N_4175);
xor U6827 (N_6827,N_4609,N_4422);
nor U6828 (N_6828,N_5197,N_5869);
nor U6829 (N_6829,N_4912,N_4372);
nor U6830 (N_6830,N_4969,N_4118);
and U6831 (N_6831,N_5177,N_4063);
nand U6832 (N_6832,N_4566,N_5191);
and U6833 (N_6833,N_5943,N_4554);
nand U6834 (N_6834,N_5886,N_5332);
nor U6835 (N_6835,N_5837,N_4898);
or U6836 (N_6836,N_5974,N_4827);
nor U6837 (N_6837,N_5234,N_4607);
nor U6838 (N_6838,N_4271,N_4880);
nand U6839 (N_6839,N_4131,N_4455);
nand U6840 (N_6840,N_5669,N_4542);
nor U6841 (N_6841,N_5252,N_4946);
nand U6842 (N_6842,N_5388,N_4267);
or U6843 (N_6843,N_5955,N_4435);
or U6844 (N_6844,N_4764,N_5542);
nand U6845 (N_6845,N_5112,N_4361);
nor U6846 (N_6846,N_4919,N_5285);
and U6847 (N_6847,N_4641,N_5106);
and U6848 (N_6848,N_5721,N_5872);
nand U6849 (N_6849,N_5978,N_5348);
nand U6850 (N_6850,N_5382,N_5959);
and U6851 (N_6851,N_5701,N_4071);
nor U6852 (N_6852,N_5787,N_5018);
nor U6853 (N_6853,N_5623,N_5264);
nor U6854 (N_6854,N_4702,N_4980);
nor U6855 (N_6855,N_4277,N_5401);
xor U6856 (N_6856,N_4790,N_5406);
nand U6857 (N_6857,N_4249,N_4196);
nor U6858 (N_6858,N_4608,N_5607);
or U6859 (N_6859,N_5424,N_5034);
and U6860 (N_6860,N_4675,N_5773);
or U6861 (N_6861,N_5453,N_5646);
or U6862 (N_6862,N_5373,N_4474);
and U6863 (N_6863,N_5123,N_5722);
or U6864 (N_6864,N_4301,N_5530);
and U6865 (N_6865,N_5975,N_5642);
and U6866 (N_6866,N_4661,N_4393);
or U6867 (N_6867,N_4821,N_4357);
or U6868 (N_6868,N_4364,N_4719);
nand U6869 (N_6869,N_5215,N_5152);
and U6870 (N_6870,N_5871,N_5257);
nand U6871 (N_6871,N_4674,N_4653);
or U6872 (N_6872,N_5599,N_4284);
and U6873 (N_6873,N_5908,N_4367);
or U6874 (N_6874,N_4619,N_5803);
nor U6875 (N_6875,N_5954,N_5848);
or U6876 (N_6876,N_4987,N_5179);
or U6877 (N_6877,N_4215,N_4345);
or U6878 (N_6878,N_4099,N_4847);
and U6879 (N_6879,N_5823,N_5114);
nand U6880 (N_6880,N_4885,N_5845);
nand U6881 (N_6881,N_4397,N_5393);
nand U6882 (N_6882,N_4830,N_4749);
or U6883 (N_6883,N_5171,N_4867);
and U6884 (N_6884,N_4430,N_5713);
xnor U6885 (N_6885,N_5031,N_4991);
nand U6886 (N_6886,N_5670,N_4163);
and U6887 (N_6887,N_5647,N_4232);
and U6888 (N_6888,N_5481,N_5704);
xnor U6889 (N_6889,N_5734,N_5891);
and U6890 (N_6890,N_5689,N_4813);
and U6891 (N_6891,N_4975,N_5269);
nand U6892 (N_6892,N_4521,N_5325);
nand U6893 (N_6893,N_5588,N_5911);
nand U6894 (N_6894,N_4931,N_5676);
and U6895 (N_6895,N_5004,N_4949);
nor U6896 (N_6896,N_4079,N_4261);
nor U6897 (N_6897,N_5652,N_5774);
nor U6898 (N_6898,N_5561,N_5947);
and U6899 (N_6899,N_4495,N_5758);
xnor U6900 (N_6900,N_5006,N_4297);
and U6901 (N_6901,N_5746,N_5478);
nand U6902 (N_6902,N_4316,N_4711);
xor U6903 (N_6903,N_4207,N_5398);
nand U6904 (N_6904,N_5820,N_5703);
or U6905 (N_6905,N_5579,N_5275);
and U6906 (N_6906,N_5472,N_4018);
nand U6907 (N_6907,N_4330,N_5860);
nor U6908 (N_6908,N_5644,N_5586);
and U6909 (N_6909,N_4114,N_5933);
and U6910 (N_6910,N_4317,N_5277);
or U6911 (N_6911,N_5074,N_5597);
or U6912 (N_6912,N_5840,N_4535);
nor U6913 (N_6913,N_5819,N_5228);
nand U6914 (N_6914,N_4596,N_5079);
and U6915 (N_6915,N_5559,N_5916);
and U6916 (N_6916,N_4052,N_5187);
nand U6917 (N_6917,N_5439,N_5204);
or U6918 (N_6918,N_4920,N_5984);
and U6919 (N_6919,N_4848,N_4621);
nand U6920 (N_6920,N_5707,N_5209);
and U6921 (N_6921,N_4229,N_5952);
and U6922 (N_6922,N_5941,N_4136);
nand U6923 (N_6923,N_4500,N_4323);
or U6924 (N_6924,N_4179,N_5850);
nor U6925 (N_6925,N_5236,N_5575);
nor U6926 (N_6926,N_5293,N_4333);
and U6927 (N_6927,N_5946,N_5649);
nand U6928 (N_6928,N_5985,N_5700);
or U6929 (N_6929,N_5977,N_4605);
xor U6930 (N_6930,N_5268,N_5150);
nand U6931 (N_6931,N_4699,N_5284);
and U6932 (N_6932,N_5282,N_4387);
nand U6933 (N_6933,N_4340,N_4941);
and U6934 (N_6934,N_4822,N_4693);
nor U6935 (N_6935,N_4151,N_4432);
and U6936 (N_6936,N_4199,N_5960);
nand U6937 (N_6937,N_5273,N_5148);
nand U6938 (N_6938,N_5483,N_4687);
nand U6939 (N_6939,N_4339,N_4120);
nor U6940 (N_6940,N_4917,N_4209);
and U6941 (N_6941,N_5657,N_4472);
nand U6942 (N_6942,N_5310,N_4436);
nand U6943 (N_6943,N_4228,N_4819);
xor U6944 (N_6944,N_5427,N_4903);
or U6945 (N_6945,N_4784,N_5270);
or U6946 (N_6946,N_4556,N_5705);
and U6947 (N_6947,N_5381,N_5315);
nor U6948 (N_6948,N_5465,N_5156);
or U6949 (N_6949,N_5421,N_4595);
or U6950 (N_6950,N_5537,N_5047);
nor U6951 (N_6951,N_4090,N_5281);
and U6952 (N_6952,N_5000,N_5636);
nor U6953 (N_6953,N_4851,N_5794);
or U6954 (N_6954,N_4698,N_5451);
and U6955 (N_6955,N_5055,N_4679);
and U6956 (N_6956,N_4732,N_4947);
and U6957 (N_6957,N_4184,N_4631);
nand U6958 (N_6958,N_5531,N_5896);
nand U6959 (N_6959,N_4265,N_5832);
nand U6960 (N_6960,N_4859,N_4473);
nand U6961 (N_6961,N_5765,N_5915);
nor U6962 (N_6962,N_5460,N_4978);
nand U6963 (N_6963,N_5219,N_4420);
nor U6964 (N_6964,N_4901,N_4160);
nand U6965 (N_6965,N_4141,N_4181);
nand U6966 (N_6966,N_4386,N_5661);
xnor U6967 (N_6967,N_5895,N_4597);
nand U6968 (N_6968,N_4101,N_5492);
and U6969 (N_6969,N_4725,N_5675);
nor U6970 (N_6970,N_5350,N_5994);
and U6971 (N_6971,N_5356,N_5548);
nand U6972 (N_6972,N_5864,N_5103);
nor U6973 (N_6973,N_4820,N_5027);
or U6974 (N_6974,N_4800,N_5893);
and U6975 (N_6975,N_4952,N_4945);
nand U6976 (N_6976,N_4615,N_5595);
nor U6977 (N_6977,N_4824,N_5395);
nor U6978 (N_6978,N_4067,N_5931);
nor U6979 (N_6979,N_5153,N_5744);
nand U6980 (N_6980,N_4936,N_4871);
nand U6981 (N_6981,N_4604,N_4841);
and U6982 (N_6982,N_4169,N_5683);
nor U6983 (N_6983,N_5987,N_4224);
nor U6984 (N_6984,N_4225,N_5857);
nand U6985 (N_6985,N_4832,N_5546);
and U6986 (N_6986,N_4035,N_4350);
and U6987 (N_6987,N_5883,N_5331);
and U6988 (N_6988,N_5030,N_4652);
nor U6989 (N_6989,N_4994,N_4510);
nor U6990 (N_6990,N_5073,N_4426);
nor U6991 (N_6991,N_5116,N_5205);
and U6992 (N_6992,N_4266,N_4007);
nand U6993 (N_6993,N_4659,N_5957);
nand U6994 (N_6994,N_5372,N_4839);
nor U6995 (N_6995,N_4633,N_4935);
or U6996 (N_6996,N_4881,N_5702);
nand U6997 (N_6997,N_4806,N_5064);
nor U6998 (N_6998,N_5291,N_5619);
nor U6999 (N_6999,N_4210,N_5796);
nor U7000 (N_7000,N_5515,N_4839);
and U7001 (N_7001,N_4082,N_5399);
nor U7002 (N_7002,N_4207,N_4293);
or U7003 (N_7003,N_5622,N_4980);
nand U7004 (N_7004,N_5753,N_5572);
nor U7005 (N_7005,N_5701,N_4887);
nand U7006 (N_7006,N_4352,N_4184);
and U7007 (N_7007,N_5761,N_4172);
nor U7008 (N_7008,N_5316,N_4462);
nor U7009 (N_7009,N_4271,N_4082);
and U7010 (N_7010,N_4573,N_4679);
nor U7011 (N_7011,N_4375,N_5438);
nand U7012 (N_7012,N_5450,N_5332);
or U7013 (N_7013,N_5360,N_4080);
xor U7014 (N_7014,N_4400,N_5131);
nand U7015 (N_7015,N_4552,N_5489);
or U7016 (N_7016,N_5925,N_4885);
nand U7017 (N_7017,N_5564,N_5874);
nor U7018 (N_7018,N_4601,N_4173);
and U7019 (N_7019,N_4829,N_4196);
nor U7020 (N_7020,N_4336,N_5544);
nor U7021 (N_7021,N_5870,N_4622);
nand U7022 (N_7022,N_4333,N_4942);
nand U7023 (N_7023,N_5267,N_4866);
or U7024 (N_7024,N_5526,N_4130);
and U7025 (N_7025,N_4625,N_5805);
nand U7026 (N_7026,N_5500,N_5528);
nand U7027 (N_7027,N_4941,N_4639);
nand U7028 (N_7028,N_5657,N_4492);
and U7029 (N_7029,N_4854,N_4762);
nor U7030 (N_7030,N_4951,N_5383);
nor U7031 (N_7031,N_5251,N_4072);
nor U7032 (N_7032,N_5368,N_5806);
nor U7033 (N_7033,N_5864,N_5975);
and U7034 (N_7034,N_4575,N_4338);
or U7035 (N_7035,N_5893,N_5179);
and U7036 (N_7036,N_4572,N_5932);
nand U7037 (N_7037,N_4456,N_5321);
nor U7038 (N_7038,N_5547,N_4224);
or U7039 (N_7039,N_5053,N_5075);
nor U7040 (N_7040,N_4400,N_5375);
or U7041 (N_7041,N_5236,N_5083);
and U7042 (N_7042,N_5726,N_5811);
nor U7043 (N_7043,N_4746,N_5814);
and U7044 (N_7044,N_4571,N_5143);
nand U7045 (N_7045,N_4095,N_4010);
nand U7046 (N_7046,N_4091,N_4112);
nor U7047 (N_7047,N_4553,N_5177);
nand U7048 (N_7048,N_4044,N_5168);
or U7049 (N_7049,N_5154,N_4632);
or U7050 (N_7050,N_4344,N_4566);
nand U7051 (N_7051,N_5397,N_4054);
and U7052 (N_7052,N_5211,N_4217);
xnor U7053 (N_7053,N_4432,N_4833);
or U7054 (N_7054,N_5179,N_5839);
or U7055 (N_7055,N_4062,N_4944);
nand U7056 (N_7056,N_4946,N_5470);
or U7057 (N_7057,N_5997,N_5190);
and U7058 (N_7058,N_5705,N_4272);
or U7059 (N_7059,N_5434,N_4462);
or U7060 (N_7060,N_5125,N_5851);
nor U7061 (N_7061,N_5259,N_4787);
or U7062 (N_7062,N_4549,N_5203);
or U7063 (N_7063,N_4210,N_5962);
nor U7064 (N_7064,N_5086,N_4718);
and U7065 (N_7065,N_5148,N_4104);
nor U7066 (N_7066,N_4987,N_4780);
or U7067 (N_7067,N_5114,N_5778);
nand U7068 (N_7068,N_5900,N_4787);
and U7069 (N_7069,N_4830,N_5707);
or U7070 (N_7070,N_4805,N_4563);
nor U7071 (N_7071,N_4919,N_5824);
and U7072 (N_7072,N_5394,N_5235);
and U7073 (N_7073,N_5032,N_5577);
and U7074 (N_7074,N_4664,N_4549);
or U7075 (N_7075,N_5755,N_5759);
or U7076 (N_7076,N_4707,N_5811);
or U7077 (N_7077,N_4958,N_5361);
nand U7078 (N_7078,N_5885,N_4585);
nand U7079 (N_7079,N_5635,N_5568);
nand U7080 (N_7080,N_4051,N_4136);
nand U7081 (N_7081,N_4573,N_5558);
and U7082 (N_7082,N_5767,N_4971);
or U7083 (N_7083,N_4721,N_4046);
and U7084 (N_7084,N_4915,N_4699);
nand U7085 (N_7085,N_5805,N_4866);
nand U7086 (N_7086,N_4813,N_5638);
nand U7087 (N_7087,N_5397,N_5022);
and U7088 (N_7088,N_5744,N_4426);
nor U7089 (N_7089,N_4080,N_5268);
nand U7090 (N_7090,N_5033,N_4255);
nand U7091 (N_7091,N_4941,N_4563);
nand U7092 (N_7092,N_4353,N_5210);
nand U7093 (N_7093,N_4072,N_5031);
or U7094 (N_7094,N_5971,N_4405);
nand U7095 (N_7095,N_4343,N_4490);
and U7096 (N_7096,N_5717,N_5878);
and U7097 (N_7097,N_5528,N_5302);
nor U7098 (N_7098,N_5567,N_4971);
nor U7099 (N_7099,N_5409,N_4368);
nand U7100 (N_7100,N_5852,N_4240);
nor U7101 (N_7101,N_5296,N_5352);
nor U7102 (N_7102,N_4388,N_5062);
or U7103 (N_7103,N_5656,N_4834);
nor U7104 (N_7104,N_5346,N_5550);
nor U7105 (N_7105,N_5408,N_4957);
or U7106 (N_7106,N_5327,N_4383);
and U7107 (N_7107,N_4112,N_4667);
nor U7108 (N_7108,N_4544,N_4184);
or U7109 (N_7109,N_4527,N_4924);
or U7110 (N_7110,N_5939,N_5366);
nor U7111 (N_7111,N_4927,N_5974);
nor U7112 (N_7112,N_4361,N_5114);
nor U7113 (N_7113,N_4622,N_4732);
and U7114 (N_7114,N_5825,N_4056);
nand U7115 (N_7115,N_4750,N_5709);
and U7116 (N_7116,N_4777,N_5670);
or U7117 (N_7117,N_5083,N_5611);
nand U7118 (N_7118,N_5706,N_5409);
and U7119 (N_7119,N_4224,N_5798);
nor U7120 (N_7120,N_5395,N_5890);
or U7121 (N_7121,N_5709,N_4756);
or U7122 (N_7122,N_4839,N_5108);
nand U7123 (N_7123,N_5335,N_4501);
and U7124 (N_7124,N_4171,N_5209);
nor U7125 (N_7125,N_4680,N_4295);
nand U7126 (N_7126,N_5263,N_5987);
nand U7127 (N_7127,N_5813,N_4304);
nand U7128 (N_7128,N_4911,N_4734);
and U7129 (N_7129,N_4498,N_4145);
and U7130 (N_7130,N_5945,N_5711);
or U7131 (N_7131,N_5801,N_4652);
nor U7132 (N_7132,N_5629,N_4584);
nor U7133 (N_7133,N_4761,N_5112);
or U7134 (N_7134,N_4589,N_4315);
nor U7135 (N_7135,N_5994,N_4099);
nor U7136 (N_7136,N_4023,N_5649);
and U7137 (N_7137,N_4294,N_4575);
nand U7138 (N_7138,N_4497,N_4665);
nor U7139 (N_7139,N_5262,N_4550);
or U7140 (N_7140,N_5139,N_4597);
and U7141 (N_7141,N_4890,N_4373);
and U7142 (N_7142,N_5695,N_4266);
and U7143 (N_7143,N_5972,N_5472);
or U7144 (N_7144,N_4780,N_5493);
or U7145 (N_7145,N_5710,N_5847);
nor U7146 (N_7146,N_4766,N_5937);
or U7147 (N_7147,N_4311,N_5175);
or U7148 (N_7148,N_4495,N_5430);
nand U7149 (N_7149,N_5581,N_4243);
and U7150 (N_7150,N_4152,N_5997);
nand U7151 (N_7151,N_4143,N_5087);
nor U7152 (N_7152,N_5942,N_5512);
nand U7153 (N_7153,N_4456,N_4759);
nor U7154 (N_7154,N_5803,N_4443);
nor U7155 (N_7155,N_5604,N_4229);
nor U7156 (N_7156,N_4799,N_5956);
and U7157 (N_7157,N_5602,N_4031);
nand U7158 (N_7158,N_4265,N_5304);
and U7159 (N_7159,N_4357,N_5786);
and U7160 (N_7160,N_4015,N_4040);
and U7161 (N_7161,N_5832,N_5690);
and U7162 (N_7162,N_4195,N_4163);
or U7163 (N_7163,N_5229,N_5344);
and U7164 (N_7164,N_4868,N_4536);
nor U7165 (N_7165,N_5069,N_4269);
xnor U7166 (N_7166,N_5486,N_5120);
nor U7167 (N_7167,N_4580,N_5098);
or U7168 (N_7168,N_4576,N_5145);
nand U7169 (N_7169,N_4757,N_5451);
nand U7170 (N_7170,N_5102,N_5668);
and U7171 (N_7171,N_4590,N_4917);
nor U7172 (N_7172,N_5815,N_4873);
nor U7173 (N_7173,N_5140,N_4204);
or U7174 (N_7174,N_5234,N_5221);
and U7175 (N_7175,N_4228,N_5791);
nand U7176 (N_7176,N_4507,N_5114);
nor U7177 (N_7177,N_5064,N_5026);
or U7178 (N_7178,N_4456,N_4464);
nand U7179 (N_7179,N_5132,N_5714);
and U7180 (N_7180,N_4110,N_4130);
nor U7181 (N_7181,N_5521,N_5023);
nor U7182 (N_7182,N_5555,N_4002);
nor U7183 (N_7183,N_5173,N_5829);
nand U7184 (N_7184,N_4065,N_5223);
nand U7185 (N_7185,N_4405,N_5132);
nor U7186 (N_7186,N_4233,N_4002);
and U7187 (N_7187,N_4465,N_5699);
nand U7188 (N_7188,N_4381,N_4724);
nor U7189 (N_7189,N_4325,N_5583);
or U7190 (N_7190,N_4786,N_4603);
nor U7191 (N_7191,N_4660,N_4844);
nand U7192 (N_7192,N_5838,N_4665);
nand U7193 (N_7193,N_4648,N_4548);
nand U7194 (N_7194,N_4165,N_5860);
nor U7195 (N_7195,N_4072,N_5474);
nand U7196 (N_7196,N_4363,N_5182);
nand U7197 (N_7197,N_4174,N_5936);
nor U7198 (N_7198,N_5341,N_4361);
nand U7199 (N_7199,N_5966,N_4437);
and U7200 (N_7200,N_4264,N_4539);
nand U7201 (N_7201,N_5208,N_5888);
nand U7202 (N_7202,N_4648,N_5886);
nor U7203 (N_7203,N_4415,N_4785);
nor U7204 (N_7204,N_4614,N_5964);
and U7205 (N_7205,N_4856,N_5682);
or U7206 (N_7206,N_4246,N_5128);
nor U7207 (N_7207,N_4371,N_4293);
or U7208 (N_7208,N_5231,N_4541);
and U7209 (N_7209,N_4556,N_4369);
nor U7210 (N_7210,N_4995,N_5368);
and U7211 (N_7211,N_4275,N_5555);
nand U7212 (N_7212,N_4278,N_5329);
nand U7213 (N_7213,N_5775,N_5714);
and U7214 (N_7214,N_5823,N_5478);
nor U7215 (N_7215,N_5826,N_4336);
or U7216 (N_7216,N_5662,N_4160);
or U7217 (N_7217,N_4466,N_4779);
or U7218 (N_7218,N_5013,N_5614);
nand U7219 (N_7219,N_5652,N_5630);
nand U7220 (N_7220,N_5800,N_4666);
nor U7221 (N_7221,N_5455,N_4350);
xnor U7222 (N_7222,N_5934,N_5815);
nand U7223 (N_7223,N_5014,N_5156);
xor U7224 (N_7224,N_4688,N_5048);
or U7225 (N_7225,N_4567,N_5358);
or U7226 (N_7226,N_4419,N_5662);
nor U7227 (N_7227,N_5515,N_4177);
nor U7228 (N_7228,N_4400,N_5004);
nor U7229 (N_7229,N_5435,N_4226);
nand U7230 (N_7230,N_5043,N_4330);
xor U7231 (N_7231,N_4828,N_5518);
or U7232 (N_7232,N_5190,N_5876);
nand U7233 (N_7233,N_5321,N_4219);
or U7234 (N_7234,N_4259,N_4402);
nor U7235 (N_7235,N_4091,N_4186);
nand U7236 (N_7236,N_4596,N_5837);
or U7237 (N_7237,N_5199,N_5054);
nand U7238 (N_7238,N_5456,N_5675);
nand U7239 (N_7239,N_5573,N_4287);
nand U7240 (N_7240,N_4273,N_5697);
nor U7241 (N_7241,N_5907,N_4322);
and U7242 (N_7242,N_5330,N_5795);
nand U7243 (N_7243,N_4019,N_5158);
or U7244 (N_7244,N_5614,N_5405);
nand U7245 (N_7245,N_5290,N_4298);
or U7246 (N_7246,N_4738,N_5531);
nand U7247 (N_7247,N_5576,N_5463);
and U7248 (N_7248,N_4816,N_5754);
or U7249 (N_7249,N_4455,N_5898);
and U7250 (N_7250,N_4652,N_4103);
or U7251 (N_7251,N_4536,N_5612);
or U7252 (N_7252,N_4916,N_5931);
or U7253 (N_7253,N_4195,N_4904);
nand U7254 (N_7254,N_4388,N_5048);
nor U7255 (N_7255,N_4398,N_4768);
and U7256 (N_7256,N_5223,N_4741);
nor U7257 (N_7257,N_5073,N_5818);
nor U7258 (N_7258,N_5611,N_4200);
and U7259 (N_7259,N_5722,N_4022);
nor U7260 (N_7260,N_4907,N_5459);
nand U7261 (N_7261,N_4763,N_4782);
and U7262 (N_7262,N_4090,N_4979);
nor U7263 (N_7263,N_5370,N_5759);
nor U7264 (N_7264,N_4260,N_4447);
and U7265 (N_7265,N_4321,N_4420);
nand U7266 (N_7266,N_5347,N_5247);
nand U7267 (N_7267,N_5252,N_4365);
and U7268 (N_7268,N_5746,N_5567);
nor U7269 (N_7269,N_5098,N_4857);
or U7270 (N_7270,N_4864,N_5260);
xnor U7271 (N_7271,N_4049,N_5989);
nor U7272 (N_7272,N_5633,N_5169);
nor U7273 (N_7273,N_4420,N_4117);
nand U7274 (N_7274,N_4600,N_4748);
and U7275 (N_7275,N_5804,N_4953);
xnor U7276 (N_7276,N_4141,N_4244);
nand U7277 (N_7277,N_4269,N_4718);
and U7278 (N_7278,N_5643,N_5791);
xor U7279 (N_7279,N_5013,N_5042);
and U7280 (N_7280,N_4383,N_4251);
xnor U7281 (N_7281,N_5881,N_5083);
nor U7282 (N_7282,N_4501,N_4692);
nand U7283 (N_7283,N_4674,N_4842);
or U7284 (N_7284,N_4909,N_5012);
nor U7285 (N_7285,N_5051,N_4216);
nor U7286 (N_7286,N_5741,N_4600);
or U7287 (N_7287,N_5432,N_4903);
nor U7288 (N_7288,N_5511,N_4809);
and U7289 (N_7289,N_5164,N_5082);
and U7290 (N_7290,N_5435,N_4253);
or U7291 (N_7291,N_4931,N_5551);
or U7292 (N_7292,N_4502,N_4993);
or U7293 (N_7293,N_4719,N_5143);
or U7294 (N_7294,N_5862,N_5997);
and U7295 (N_7295,N_4754,N_4267);
or U7296 (N_7296,N_4728,N_4335);
nor U7297 (N_7297,N_5841,N_5155);
or U7298 (N_7298,N_5993,N_5103);
and U7299 (N_7299,N_5909,N_5878);
nand U7300 (N_7300,N_4862,N_5811);
nor U7301 (N_7301,N_4047,N_5841);
and U7302 (N_7302,N_4677,N_5670);
nor U7303 (N_7303,N_5792,N_4609);
and U7304 (N_7304,N_5762,N_5649);
and U7305 (N_7305,N_4803,N_4037);
and U7306 (N_7306,N_5524,N_4982);
nor U7307 (N_7307,N_4035,N_5570);
or U7308 (N_7308,N_5607,N_5972);
and U7309 (N_7309,N_4837,N_4017);
nand U7310 (N_7310,N_4797,N_4847);
nand U7311 (N_7311,N_4730,N_5920);
and U7312 (N_7312,N_4816,N_4571);
nor U7313 (N_7313,N_4425,N_4524);
nor U7314 (N_7314,N_4698,N_5719);
and U7315 (N_7315,N_4429,N_5693);
nor U7316 (N_7316,N_4160,N_5598);
nand U7317 (N_7317,N_5869,N_4024);
and U7318 (N_7318,N_5835,N_5222);
and U7319 (N_7319,N_4278,N_5181);
nor U7320 (N_7320,N_4748,N_4847);
nor U7321 (N_7321,N_4441,N_4862);
or U7322 (N_7322,N_5805,N_5827);
and U7323 (N_7323,N_4410,N_4749);
nor U7324 (N_7324,N_4580,N_4405);
nand U7325 (N_7325,N_4167,N_4607);
or U7326 (N_7326,N_5643,N_4667);
and U7327 (N_7327,N_5222,N_5672);
and U7328 (N_7328,N_5772,N_5161);
nand U7329 (N_7329,N_5645,N_4770);
xnor U7330 (N_7330,N_4736,N_4773);
nand U7331 (N_7331,N_4603,N_4196);
or U7332 (N_7332,N_4140,N_4263);
or U7333 (N_7333,N_5197,N_5544);
nand U7334 (N_7334,N_4952,N_5393);
nor U7335 (N_7335,N_4177,N_5767);
nor U7336 (N_7336,N_4622,N_5328);
and U7337 (N_7337,N_4716,N_4180);
nand U7338 (N_7338,N_5106,N_4436);
nor U7339 (N_7339,N_4263,N_4595);
and U7340 (N_7340,N_5143,N_4077);
nand U7341 (N_7341,N_4199,N_4971);
and U7342 (N_7342,N_4049,N_4016);
nand U7343 (N_7343,N_4434,N_5480);
nor U7344 (N_7344,N_4058,N_4676);
nor U7345 (N_7345,N_5127,N_5323);
xor U7346 (N_7346,N_5570,N_5023);
or U7347 (N_7347,N_4073,N_4899);
and U7348 (N_7348,N_4182,N_5222);
nor U7349 (N_7349,N_5816,N_5996);
and U7350 (N_7350,N_5522,N_4473);
nor U7351 (N_7351,N_5684,N_5830);
or U7352 (N_7352,N_4048,N_4076);
or U7353 (N_7353,N_4033,N_5626);
nor U7354 (N_7354,N_4473,N_4650);
or U7355 (N_7355,N_4933,N_5153);
and U7356 (N_7356,N_5569,N_4755);
nand U7357 (N_7357,N_4523,N_4128);
nand U7358 (N_7358,N_5025,N_4736);
and U7359 (N_7359,N_5159,N_4155);
and U7360 (N_7360,N_5834,N_5602);
and U7361 (N_7361,N_5104,N_5788);
xor U7362 (N_7362,N_5991,N_5280);
nand U7363 (N_7363,N_4398,N_4430);
nor U7364 (N_7364,N_4377,N_5291);
nor U7365 (N_7365,N_4792,N_5922);
and U7366 (N_7366,N_4091,N_4109);
nor U7367 (N_7367,N_5880,N_4922);
and U7368 (N_7368,N_4016,N_5885);
xnor U7369 (N_7369,N_4318,N_5789);
nor U7370 (N_7370,N_5041,N_5737);
or U7371 (N_7371,N_5422,N_5412);
nor U7372 (N_7372,N_5627,N_4672);
nor U7373 (N_7373,N_4003,N_5657);
nand U7374 (N_7374,N_4191,N_5167);
or U7375 (N_7375,N_4161,N_4715);
nor U7376 (N_7376,N_5938,N_4069);
or U7377 (N_7377,N_4520,N_5894);
and U7378 (N_7378,N_4260,N_4140);
or U7379 (N_7379,N_4679,N_5690);
or U7380 (N_7380,N_4261,N_4602);
nand U7381 (N_7381,N_5248,N_4429);
and U7382 (N_7382,N_4764,N_5927);
and U7383 (N_7383,N_4772,N_4093);
and U7384 (N_7384,N_5915,N_5362);
nor U7385 (N_7385,N_5076,N_5634);
nor U7386 (N_7386,N_4174,N_5355);
or U7387 (N_7387,N_5402,N_5131);
xnor U7388 (N_7388,N_5774,N_4050);
nor U7389 (N_7389,N_5061,N_5944);
nor U7390 (N_7390,N_5480,N_4660);
nor U7391 (N_7391,N_4527,N_5266);
nand U7392 (N_7392,N_5463,N_5212);
nand U7393 (N_7393,N_5592,N_4556);
nand U7394 (N_7394,N_5374,N_4478);
and U7395 (N_7395,N_4650,N_5393);
nand U7396 (N_7396,N_5181,N_4011);
or U7397 (N_7397,N_4890,N_5322);
or U7398 (N_7398,N_5159,N_4375);
or U7399 (N_7399,N_4325,N_4029);
or U7400 (N_7400,N_4542,N_5664);
nand U7401 (N_7401,N_5448,N_4520);
nor U7402 (N_7402,N_5100,N_5153);
and U7403 (N_7403,N_4501,N_4301);
nor U7404 (N_7404,N_5650,N_4107);
and U7405 (N_7405,N_5217,N_4373);
nor U7406 (N_7406,N_5279,N_4110);
or U7407 (N_7407,N_4408,N_4323);
nor U7408 (N_7408,N_4193,N_5029);
and U7409 (N_7409,N_5900,N_5453);
and U7410 (N_7410,N_5215,N_5621);
nand U7411 (N_7411,N_4267,N_5836);
nand U7412 (N_7412,N_5697,N_4447);
nand U7413 (N_7413,N_5686,N_4610);
nor U7414 (N_7414,N_4316,N_4597);
nor U7415 (N_7415,N_4139,N_4698);
xnor U7416 (N_7416,N_5601,N_5363);
nor U7417 (N_7417,N_4157,N_4033);
and U7418 (N_7418,N_5523,N_5016);
xnor U7419 (N_7419,N_5721,N_4430);
nor U7420 (N_7420,N_4787,N_4465);
nand U7421 (N_7421,N_4667,N_4222);
and U7422 (N_7422,N_4084,N_4117);
nor U7423 (N_7423,N_5671,N_4713);
nor U7424 (N_7424,N_4839,N_4300);
nand U7425 (N_7425,N_4299,N_5585);
or U7426 (N_7426,N_4695,N_4179);
nand U7427 (N_7427,N_5587,N_5015);
and U7428 (N_7428,N_4761,N_5158);
nand U7429 (N_7429,N_5890,N_4577);
and U7430 (N_7430,N_4636,N_4410);
or U7431 (N_7431,N_4368,N_4049);
and U7432 (N_7432,N_4875,N_5432);
or U7433 (N_7433,N_4900,N_5597);
xor U7434 (N_7434,N_5151,N_5821);
nand U7435 (N_7435,N_5758,N_4039);
or U7436 (N_7436,N_4247,N_4064);
or U7437 (N_7437,N_5402,N_4916);
or U7438 (N_7438,N_4280,N_5886);
and U7439 (N_7439,N_4278,N_4507);
nor U7440 (N_7440,N_5870,N_4412);
or U7441 (N_7441,N_4990,N_5120);
and U7442 (N_7442,N_4573,N_4865);
nor U7443 (N_7443,N_4873,N_4761);
nand U7444 (N_7444,N_5089,N_4059);
or U7445 (N_7445,N_4784,N_5739);
or U7446 (N_7446,N_5862,N_5579);
and U7447 (N_7447,N_4613,N_5320);
nand U7448 (N_7448,N_4155,N_5425);
nor U7449 (N_7449,N_5619,N_4128);
and U7450 (N_7450,N_5767,N_5775);
nand U7451 (N_7451,N_4703,N_5995);
xor U7452 (N_7452,N_4703,N_4466);
nor U7453 (N_7453,N_5935,N_4292);
xnor U7454 (N_7454,N_4549,N_5759);
nand U7455 (N_7455,N_5182,N_5071);
nand U7456 (N_7456,N_5066,N_5157);
or U7457 (N_7457,N_4851,N_4183);
nand U7458 (N_7458,N_5181,N_4106);
or U7459 (N_7459,N_4505,N_4440);
and U7460 (N_7460,N_5706,N_5353);
nor U7461 (N_7461,N_4824,N_5176);
or U7462 (N_7462,N_4039,N_4046);
nor U7463 (N_7463,N_5011,N_4183);
or U7464 (N_7464,N_5442,N_5626);
or U7465 (N_7465,N_5614,N_5057);
nand U7466 (N_7466,N_4157,N_4076);
and U7467 (N_7467,N_5799,N_4407);
nand U7468 (N_7468,N_5109,N_5544);
xnor U7469 (N_7469,N_5940,N_4713);
nand U7470 (N_7470,N_4905,N_5434);
and U7471 (N_7471,N_4763,N_5934);
or U7472 (N_7472,N_4892,N_4441);
xor U7473 (N_7473,N_5596,N_4923);
or U7474 (N_7474,N_5341,N_5899);
nand U7475 (N_7475,N_4613,N_5562);
nand U7476 (N_7476,N_5755,N_4557);
xor U7477 (N_7477,N_5040,N_4353);
nor U7478 (N_7478,N_5216,N_5104);
nor U7479 (N_7479,N_5108,N_4402);
and U7480 (N_7480,N_4743,N_4517);
nor U7481 (N_7481,N_5072,N_5078);
or U7482 (N_7482,N_5828,N_5000);
nor U7483 (N_7483,N_5620,N_5360);
nor U7484 (N_7484,N_5877,N_5509);
and U7485 (N_7485,N_4646,N_4706);
nor U7486 (N_7486,N_5848,N_5431);
nand U7487 (N_7487,N_4455,N_5224);
nand U7488 (N_7488,N_4208,N_4823);
or U7489 (N_7489,N_4919,N_5277);
nand U7490 (N_7490,N_4351,N_5224);
or U7491 (N_7491,N_4013,N_4920);
nand U7492 (N_7492,N_5095,N_5056);
nand U7493 (N_7493,N_5925,N_5500);
and U7494 (N_7494,N_4156,N_5323);
or U7495 (N_7495,N_5179,N_4525);
or U7496 (N_7496,N_5648,N_5073);
nor U7497 (N_7497,N_4508,N_4986);
nand U7498 (N_7498,N_5534,N_5669);
and U7499 (N_7499,N_5023,N_4513);
nor U7500 (N_7500,N_5449,N_4530);
and U7501 (N_7501,N_5497,N_5464);
nand U7502 (N_7502,N_5870,N_4537);
nor U7503 (N_7503,N_5863,N_5129);
nand U7504 (N_7504,N_4464,N_5556);
nor U7505 (N_7505,N_5352,N_5954);
nor U7506 (N_7506,N_4620,N_4731);
xor U7507 (N_7507,N_5987,N_4552);
and U7508 (N_7508,N_5896,N_5796);
and U7509 (N_7509,N_5828,N_4055);
nor U7510 (N_7510,N_4441,N_4195);
nand U7511 (N_7511,N_4161,N_4090);
or U7512 (N_7512,N_4192,N_4681);
nand U7513 (N_7513,N_5289,N_5060);
or U7514 (N_7514,N_4799,N_4098);
nand U7515 (N_7515,N_4215,N_5300);
or U7516 (N_7516,N_4288,N_5623);
and U7517 (N_7517,N_4247,N_5606);
or U7518 (N_7518,N_5786,N_5774);
nor U7519 (N_7519,N_5768,N_4148);
and U7520 (N_7520,N_4697,N_4893);
nor U7521 (N_7521,N_5607,N_5578);
nand U7522 (N_7522,N_4944,N_4859);
nand U7523 (N_7523,N_5811,N_5019);
nand U7524 (N_7524,N_5291,N_5478);
nand U7525 (N_7525,N_5140,N_5652);
or U7526 (N_7526,N_5700,N_4451);
nor U7527 (N_7527,N_5774,N_4881);
nor U7528 (N_7528,N_4826,N_5609);
nand U7529 (N_7529,N_4574,N_5929);
and U7530 (N_7530,N_4394,N_4662);
nor U7531 (N_7531,N_5171,N_4596);
nand U7532 (N_7532,N_4769,N_5470);
nand U7533 (N_7533,N_5776,N_5653);
nand U7534 (N_7534,N_4313,N_5078);
nand U7535 (N_7535,N_4846,N_5141);
nand U7536 (N_7536,N_5902,N_5600);
nor U7537 (N_7537,N_4994,N_5955);
or U7538 (N_7538,N_5335,N_4930);
nand U7539 (N_7539,N_4200,N_5454);
and U7540 (N_7540,N_5244,N_5605);
and U7541 (N_7541,N_5476,N_5790);
and U7542 (N_7542,N_5131,N_4727);
xor U7543 (N_7543,N_4791,N_5757);
nor U7544 (N_7544,N_4203,N_5475);
nand U7545 (N_7545,N_4528,N_5259);
nor U7546 (N_7546,N_4814,N_4894);
nor U7547 (N_7547,N_5700,N_5662);
nor U7548 (N_7548,N_5917,N_4973);
nor U7549 (N_7549,N_5825,N_5376);
nand U7550 (N_7550,N_4411,N_5554);
nor U7551 (N_7551,N_4440,N_4676);
or U7552 (N_7552,N_4654,N_4423);
and U7553 (N_7553,N_5998,N_4433);
nand U7554 (N_7554,N_5543,N_4665);
nor U7555 (N_7555,N_4537,N_4601);
nor U7556 (N_7556,N_5674,N_4369);
nand U7557 (N_7557,N_5314,N_4338);
and U7558 (N_7558,N_5512,N_4805);
or U7559 (N_7559,N_5699,N_5353);
or U7560 (N_7560,N_4924,N_4506);
and U7561 (N_7561,N_5057,N_5357);
and U7562 (N_7562,N_4788,N_4157);
and U7563 (N_7563,N_4034,N_4755);
or U7564 (N_7564,N_5092,N_4145);
or U7565 (N_7565,N_5551,N_5514);
nor U7566 (N_7566,N_4948,N_4106);
or U7567 (N_7567,N_5570,N_4782);
and U7568 (N_7568,N_4359,N_5302);
and U7569 (N_7569,N_4119,N_4625);
nand U7570 (N_7570,N_4318,N_5575);
and U7571 (N_7571,N_4555,N_5213);
nor U7572 (N_7572,N_5195,N_4942);
nor U7573 (N_7573,N_5428,N_5084);
nor U7574 (N_7574,N_4685,N_5707);
nand U7575 (N_7575,N_4286,N_5765);
or U7576 (N_7576,N_5457,N_4441);
nand U7577 (N_7577,N_5504,N_5907);
and U7578 (N_7578,N_4992,N_5380);
nor U7579 (N_7579,N_4939,N_5312);
nor U7580 (N_7580,N_5524,N_5716);
xnor U7581 (N_7581,N_4995,N_5320);
nand U7582 (N_7582,N_4530,N_5779);
or U7583 (N_7583,N_5576,N_4336);
nand U7584 (N_7584,N_4240,N_5634);
nand U7585 (N_7585,N_5260,N_5776);
nor U7586 (N_7586,N_4333,N_4382);
nand U7587 (N_7587,N_5447,N_5992);
nand U7588 (N_7588,N_4242,N_5762);
xnor U7589 (N_7589,N_5447,N_5621);
and U7590 (N_7590,N_4457,N_5505);
or U7591 (N_7591,N_4385,N_5555);
and U7592 (N_7592,N_5919,N_5087);
or U7593 (N_7593,N_5473,N_5117);
xnor U7594 (N_7594,N_4234,N_5005);
and U7595 (N_7595,N_5069,N_5062);
or U7596 (N_7596,N_5797,N_4915);
nand U7597 (N_7597,N_5360,N_4230);
nand U7598 (N_7598,N_4471,N_4395);
and U7599 (N_7599,N_4613,N_4310);
or U7600 (N_7600,N_5776,N_4780);
nand U7601 (N_7601,N_5187,N_4977);
or U7602 (N_7602,N_4057,N_4666);
and U7603 (N_7603,N_4505,N_5194);
or U7604 (N_7604,N_4809,N_4824);
nand U7605 (N_7605,N_5109,N_5710);
xnor U7606 (N_7606,N_5488,N_4244);
nor U7607 (N_7607,N_5709,N_4691);
nor U7608 (N_7608,N_4461,N_5216);
nor U7609 (N_7609,N_5945,N_5471);
xnor U7610 (N_7610,N_5027,N_4953);
nor U7611 (N_7611,N_5420,N_4217);
or U7612 (N_7612,N_5886,N_5059);
and U7613 (N_7613,N_5499,N_5539);
nor U7614 (N_7614,N_4966,N_5112);
or U7615 (N_7615,N_4215,N_5849);
and U7616 (N_7616,N_5037,N_4981);
nor U7617 (N_7617,N_5701,N_5658);
or U7618 (N_7618,N_4551,N_4881);
nand U7619 (N_7619,N_5289,N_4516);
nor U7620 (N_7620,N_4281,N_5683);
and U7621 (N_7621,N_5345,N_4513);
nor U7622 (N_7622,N_4205,N_4170);
or U7623 (N_7623,N_4484,N_4139);
and U7624 (N_7624,N_5915,N_5447);
or U7625 (N_7625,N_5920,N_5280);
and U7626 (N_7626,N_4250,N_5098);
nand U7627 (N_7627,N_5772,N_4171);
or U7628 (N_7628,N_5730,N_5567);
nor U7629 (N_7629,N_4380,N_4904);
or U7630 (N_7630,N_5825,N_4733);
and U7631 (N_7631,N_5825,N_5220);
and U7632 (N_7632,N_5031,N_4394);
and U7633 (N_7633,N_4140,N_4355);
and U7634 (N_7634,N_4936,N_5492);
nor U7635 (N_7635,N_5746,N_4879);
or U7636 (N_7636,N_5210,N_4014);
and U7637 (N_7637,N_5433,N_4257);
or U7638 (N_7638,N_4864,N_4417);
or U7639 (N_7639,N_5102,N_5776);
and U7640 (N_7640,N_4309,N_5762);
nand U7641 (N_7641,N_5470,N_5613);
xnor U7642 (N_7642,N_4771,N_4545);
and U7643 (N_7643,N_5426,N_5672);
and U7644 (N_7644,N_5233,N_4198);
nand U7645 (N_7645,N_4010,N_5126);
nand U7646 (N_7646,N_5713,N_5935);
or U7647 (N_7647,N_5137,N_4291);
or U7648 (N_7648,N_5871,N_4987);
or U7649 (N_7649,N_4026,N_4273);
or U7650 (N_7650,N_5123,N_4376);
or U7651 (N_7651,N_5149,N_5954);
and U7652 (N_7652,N_4530,N_4159);
or U7653 (N_7653,N_5825,N_5712);
or U7654 (N_7654,N_5169,N_4549);
nor U7655 (N_7655,N_4116,N_4358);
and U7656 (N_7656,N_4344,N_4497);
nand U7657 (N_7657,N_5290,N_5425);
nand U7658 (N_7658,N_5067,N_4137);
and U7659 (N_7659,N_5970,N_5437);
or U7660 (N_7660,N_5153,N_5936);
and U7661 (N_7661,N_4589,N_5546);
nand U7662 (N_7662,N_5973,N_5862);
or U7663 (N_7663,N_5998,N_5622);
nor U7664 (N_7664,N_5415,N_5293);
nor U7665 (N_7665,N_4540,N_4990);
and U7666 (N_7666,N_4034,N_4896);
xor U7667 (N_7667,N_5025,N_4883);
or U7668 (N_7668,N_4940,N_5611);
and U7669 (N_7669,N_5722,N_5995);
nor U7670 (N_7670,N_5065,N_4276);
or U7671 (N_7671,N_4095,N_4136);
or U7672 (N_7672,N_5417,N_5305);
or U7673 (N_7673,N_4325,N_4006);
nor U7674 (N_7674,N_5472,N_4298);
nor U7675 (N_7675,N_5887,N_4380);
nand U7676 (N_7676,N_5698,N_5285);
or U7677 (N_7677,N_4909,N_5550);
nand U7678 (N_7678,N_4490,N_4482);
or U7679 (N_7679,N_4042,N_5515);
xor U7680 (N_7680,N_4206,N_5031);
and U7681 (N_7681,N_4946,N_4787);
and U7682 (N_7682,N_5364,N_5501);
xor U7683 (N_7683,N_5717,N_5832);
or U7684 (N_7684,N_5766,N_5664);
or U7685 (N_7685,N_5550,N_4706);
xnor U7686 (N_7686,N_4423,N_5470);
nor U7687 (N_7687,N_5142,N_5242);
and U7688 (N_7688,N_4511,N_5227);
xnor U7689 (N_7689,N_5636,N_5439);
nand U7690 (N_7690,N_4432,N_4184);
and U7691 (N_7691,N_4605,N_5725);
or U7692 (N_7692,N_5968,N_5738);
or U7693 (N_7693,N_5537,N_5232);
nand U7694 (N_7694,N_4056,N_4925);
nand U7695 (N_7695,N_4010,N_5333);
nor U7696 (N_7696,N_5212,N_5740);
or U7697 (N_7697,N_5796,N_5161);
or U7698 (N_7698,N_4787,N_5215);
and U7699 (N_7699,N_4254,N_4228);
nor U7700 (N_7700,N_5091,N_4373);
or U7701 (N_7701,N_4580,N_5084);
and U7702 (N_7702,N_4127,N_4082);
and U7703 (N_7703,N_5896,N_4434);
nand U7704 (N_7704,N_4710,N_5017);
or U7705 (N_7705,N_5857,N_4443);
and U7706 (N_7706,N_5958,N_4098);
and U7707 (N_7707,N_4118,N_4127);
and U7708 (N_7708,N_4476,N_4643);
and U7709 (N_7709,N_4210,N_4522);
nand U7710 (N_7710,N_4694,N_4541);
or U7711 (N_7711,N_5446,N_5147);
and U7712 (N_7712,N_4476,N_5574);
xor U7713 (N_7713,N_4143,N_4260);
and U7714 (N_7714,N_4480,N_4506);
nand U7715 (N_7715,N_5601,N_4111);
or U7716 (N_7716,N_5845,N_4473);
nand U7717 (N_7717,N_5193,N_5847);
nor U7718 (N_7718,N_5586,N_4896);
xor U7719 (N_7719,N_4318,N_5809);
or U7720 (N_7720,N_4774,N_4293);
nor U7721 (N_7721,N_4176,N_4843);
and U7722 (N_7722,N_4013,N_5882);
or U7723 (N_7723,N_5542,N_5589);
and U7724 (N_7724,N_5305,N_5569);
nor U7725 (N_7725,N_4465,N_5618);
nand U7726 (N_7726,N_4340,N_4232);
nand U7727 (N_7727,N_5921,N_5201);
nor U7728 (N_7728,N_4165,N_4030);
or U7729 (N_7729,N_5806,N_5295);
nor U7730 (N_7730,N_5064,N_5048);
xnor U7731 (N_7731,N_5930,N_4840);
and U7732 (N_7732,N_5084,N_5259);
nor U7733 (N_7733,N_4860,N_5193);
nor U7734 (N_7734,N_4384,N_5623);
nor U7735 (N_7735,N_5055,N_5540);
or U7736 (N_7736,N_4214,N_5695);
nand U7737 (N_7737,N_5927,N_4875);
nor U7738 (N_7738,N_4098,N_5462);
nand U7739 (N_7739,N_4937,N_5663);
or U7740 (N_7740,N_4846,N_5687);
nor U7741 (N_7741,N_4203,N_4085);
nor U7742 (N_7742,N_5639,N_5174);
or U7743 (N_7743,N_5863,N_4062);
or U7744 (N_7744,N_4890,N_5908);
or U7745 (N_7745,N_4769,N_4553);
nor U7746 (N_7746,N_5843,N_5113);
or U7747 (N_7747,N_5508,N_4720);
and U7748 (N_7748,N_5515,N_4068);
and U7749 (N_7749,N_4192,N_4997);
and U7750 (N_7750,N_5320,N_5539);
nor U7751 (N_7751,N_5851,N_5106);
or U7752 (N_7752,N_4367,N_4202);
and U7753 (N_7753,N_5640,N_4729);
or U7754 (N_7754,N_4898,N_4209);
and U7755 (N_7755,N_4158,N_4924);
nand U7756 (N_7756,N_5681,N_5698);
or U7757 (N_7757,N_5226,N_5882);
and U7758 (N_7758,N_5488,N_4146);
and U7759 (N_7759,N_5899,N_5583);
and U7760 (N_7760,N_4567,N_5355);
nand U7761 (N_7761,N_5620,N_5819);
and U7762 (N_7762,N_4105,N_5973);
nor U7763 (N_7763,N_5554,N_4562);
and U7764 (N_7764,N_4423,N_5117);
nand U7765 (N_7765,N_5675,N_4979);
or U7766 (N_7766,N_5711,N_5450);
nand U7767 (N_7767,N_5792,N_5416);
or U7768 (N_7768,N_4038,N_4401);
and U7769 (N_7769,N_4205,N_5041);
nand U7770 (N_7770,N_4508,N_5702);
nand U7771 (N_7771,N_5736,N_4721);
nand U7772 (N_7772,N_4325,N_4480);
or U7773 (N_7773,N_5462,N_4356);
nand U7774 (N_7774,N_4344,N_4181);
and U7775 (N_7775,N_5452,N_5910);
and U7776 (N_7776,N_4484,N_5628);
nor U7777 (N_7777,N_5697,N_4281);
and U7778 (N_7778,N_5237,N_5290);
nor U7779 (N_7779,N_4264,N_5219);
or U7780 (N_7780,N_5835,N_5780);
nand U7781 (N_7781,N_5070,N_5063);
nand U7782 (N_7782,N_5996,N_5069);
and U7783 (N_7783,N_5777,N_5318);
and U7784 (N_7784,N_4095,N_4301);
nand U7785 (N_7785,N_4942,N_4857);
and U7786 (N_7786,N_4027,N_4820);
or U7787 (N_7787,N_4822,N_4700);
and U7788 (N_7788,N_5124,N_4287);
and U7789 (N_7789,N_4437,N_5437);
xor U7790 (N_7790,N_4604,N_5818);
and U7791 (N_7791,N_5342,N_5728);
nand U7792 (N_7792,N_5850,N_5891);
or U7793 (N_7793,N_5929,N_5353);
or U7794 (N_7794,N_5066,N_5930);
and U7795 (N_7795,N_5805,N_4674);
and U7796 (N_7796,N_4020,N_5387);
nor U7797 (N_7797,N_4231,N_4312);
nor U7798 (N_7798,N_5400,N_5555);
nand U7799 (N_7799,N_4114,N_5451);
nand U7800 (N_7800,N_4276,N_5482);
and U7801 (N_7801,N_5358,N_5605);
or U7802 (N_7802,N_5219,N_5331);
or U7803 (N_7803,N_4453,N_4594);
or U7804 (N_7804,N_5683,N_4853);
and U7805 (N_7805,N_5175,N_4110);
nor U7806 (N_7806,N_4160,N_5193);
and U7807 (N_7807,N_4841,N_5753);
nor U7808 (N_7808,N_4829,N_4257);
or U7809 (N_7809,N_5064,N_4125);
nor U7810 (N_7810,N_4692,N_5368);
and U7811 (N_7811,N_4200,N_4723);
or U7812 (N_7812,N_4950,N_5647);
nor U7813 (N_7813,N_5511,N_4073);
xnor U7814 (N_7814,N_4416,N_4045);
nor U7815 (N_7815,N_4787,N_5165);
nand U7816 (N_7816,N_4479,N_5902);
or U7817 (N_7817,N_4828,N_4229);
nor U7818 (N_7818,N_5561,N_5874);
nor U7819 (N_7819,N_5392,N_5899);
or U7820 (N_7820,N_4693,N_4524);
and U7821 (N_7821,N_5802,N_5783);
nor U7822 (N_7822,N_5179,N_4605);
nand U7823 (N_7823,N_4391,N_5328);
or U7824 (N_7824,N_4600,N_4425);
and U7825 (N_7825,N_4697,N_5160);
nand U7826 (N_7826,N_4729,N_5579);
and U7827 (N_7827,N_5494,N_5500);
nand U7828 (N_7828,N_4319,N_5748);
or U7829 (N_7829,N_4333,N_5877);
and U7830 (N_7830,N_4381,N_4147);
or U7831 (N_7831,N_4331,N_5859);
nand U7832 (N_7832,N_4616,N_4355);
and U7833 (N_7833,N_5881,N_5710);
or U7834 (N_7834,N_4991,N_5918);
or U7835 (N_7835,N_4133,N_4963);
or U7836 (N_7836,N_4521,N_4998);
and U7837 (N_7837,N_4258,N_5689);
or U7838 (N_7838,N_5868,N_4435);
or U7839 (N_7839,N_5356,N_5881);
nor U7840 (N_7840,N_4251,N_5893);
nand U7841 (N_7841,N_4950,N_5846);
nand U7842 (N_7842,N_5066,N_5251);
and U7843 (N_7843,N_5219,N_5657);
and U7844 (N_7844,N_4779,N_5755);
and U7845 (N_7845,N_5356,N_5162);
or U7846 (N_7846,N_4621,N_4044);
and U7847 (N_7847,N_4331,N_5590);
nand U7848 (N_7848,N_5360,N_4506);
and U7849 (N_7849,N_4882,N_5021);
xor U7850 (N_7850,N_5984,N_5996);
nor U7851 (N_7851,N_5136,N_4060);
and U7852 (N_7852,N_4240,N_5217);
or U7853 (N_7853,N_5914,N_4567);
nand U7854 (N_7854,N_5797,N_4129);
nand U7855 (N_7855,N_5207,N_4548);
nand U7856 (N_7856,N_4513,N_5177);
or U7857 (N_7857,N_5421,N_4601);
nand U7858 (N_7858,N_5744,N_5550);
and U7859 (N_7859,N_4931,N_5153);
nand U7860 (N_7860,N_5692,N_5212);
and U7861 (N_7861,N_4006,N_5364);
nor U7862 (N_7862,N_5712,N_5615);
and U7863 (N_7863,N_4389,N_4703);
and U7864 (N_7864,N_4320,N_4084);
and U7865 (N_7865,N_4633,N_5475);
nor U7866 (N_7866,N_4694,N_4618);
or U7867 (N_7867,N_4687,N_4286);
and U7868 (N_7868,N_5206,N_5520);
or U7869 (N_7869,N_4575,N_5309);
nor U7870 (N_7870,N_5082,N_5333);
or U7871 (N_7871,N_4049,N_4053);
nand U7872 (N_7872,N_5770,N_4667);
nor U7873 (N_7873,N_4663,N_4239);
or U7874 (N_7874,N_4839,N_5949);
or U7875 (N_7875,N_5570,N_4631);
and U7876 (N_7876,N_5950,N_4019);
and U7877 (N_7877,N_5032,N_4144);
and U7878 (N_7878,N_4731,N_5623);
and U7879 (N_7879,N_4941,N_5510);
nor U7880 (N_7880,N_5737,N_4530);
nor U7881 (N_7881,N_5663,N_4466);
and U7882 (N_7882,N_5460,N_5163);
and U7883 (N_7883,N_4582,N_4363);
and U7884 (N_7884,N_4417,N_5742);
nand U7885 (N_7885,N_4800,N_4913);
or U7886 (N_7886,N_5559,N_5131);
and U7887 (N_7887,N_4488,N_5368);
or U7888 (N_7888,N_4022,N_5128);
nand U7889 (N_7889,N_4081,N_4777);
nand U7890 (N_7890,N_4590,N_5961);
nand U7891 (N_7891,N_5563,N_4928);
nor U7892 (N_7892,N_4170,N_5315);
nand U7893 (N_7893,N_5600,N_5388);
or U7894 (N_7894,N_4204,N_4626);
and U7895 (N_7895,N_4597,N_4905);
nor U7896 (N_7896,N_4991,N_4489);
or U7897 (N_7897,N_5733,N_5703);
nand U7898 (N_7898,N_5750,N_5609);
nor U7899 (N_7899,N_4263,N_4549);
nor U7900 (N_7900,N_5905,N_5671);
nand U7901 (N_7901,N_4240,N_5103);
nor U7902 (N_7902,N_4975,N_5273);
or U7903 (N_7903,N_4741,N_4662);
nand U7904 (N_7904,N_4083,N_4959);
nand U7905 (N_7905,N_5340,N_5663);
or U7906 (N_7906,N_5954,N_4265);
nand U7907 (N_7907,N_5845,N_4043);
xnor U7908 (N_7908,N_5950,N_5104);
nor U7909 (N_7909,N_4363,N_4508);
nand U7910 (N_7910,N_4584,N_5598);
nand U7911 (N_7911,N_4605,N_4861);
and U7912 (N_7912,N_4003,N_5820);
nand U7913 (N_7913,N_5262,N_4891);
and U7914 (N_7914,N_4165,N_5727);
nor U7915 (N_7915,N_5214,N_4357);
and U7916 (N_7916,N_5362,N_4030);
nand U7917 (N_7917,N_5454,N_5142);
nor U7918 (N_7918,N_4607,N_5195);
or U7919 (N_7919,N_5972,N_5593);
nor U7920 (N_7920,N_4399,N_4035);
nor U7921 (N_7921,N_5995,N_4815);
nand U7922 (N_7922,N_4530,N_5377);
or U7923 (N_7923,N_4589,N_4057);
nand U7924 (N_7924,N_5474,N_4652);
nor U7925 (N_7925,N_5775,N_5408);
nand U7926 (N_7926,N_5991,N_4335);
xor U7927 (N_7927,N_4162,N_4175);
nand U7928 (N_7928,N_5147,N_4070);
xnor U7929 (N_7929,N_5553,N_4236);
nand U7930 (N_7930,N_4014,N_4419);
nor U7931 (N_7931,N_4601,N_4763);
nand U7932 (N_7932,N_5651,N_5439);
or U7933 (N_7933,N_4918,N_4200);
or U7934 (N_7934,N_4599,N_4211);
or U7935 (N_7935,N_4086,N_5388);
and U7936 (N_7936,N_5947,N_5524);
or U7937 (N_7937,N_4041,N_4869);
or U7938 (N_7938,N_5741,N_5072);
and U7939 (N_7939,N_4492,N_4328);
nand U7940 (N_7940,N_5774,N_4004);
nor U7941 (N_7941,N_5565,N_5029);
xor U7942 (N_7942,N_5615,N_4251);
and U7943 (N_7943,N_5325,N_5806);
nor U7944 (N_7944,N_4481,N_4874);
xnor U7945 (N_7945,N_5039,N_4746);
or U7946 (N_7946,N_5594,N_5018);
and U7947 (N_7947,N_5364,N_4135);
nor U7948 (N_7948,N_5939,N_5383);
nor U7949 (N_7949,N_4489,N_5777);
xnor U7950 (N_7950,N_5531,N_5961);
nand U7951 (N_7951,N_4789,N_4949);
and U7952 (N_7952,N_5082,N_5654);
nor U7953 (N_7953,N_5254,N_5439);
nor U7954 (N_7954,N_5272,N_5113);
nand U7955 (N_7955,N_4869,N_4750);
nor U7956 (N_7956,N_4844,N_5017);
and U7957 (N_7957,N_4324,N_4199);
nor U7958 (N_7958,N_5368,N_5981);
nand U7959 (N_7959,N_4317,N_4850);
nand U7960 (N_7960,N_5739,N_5579);
and U7961 (N_7961,N_5663,N_5188);
nand U7962 (N_7962,N_4670,N_4121);
xnor U7963 (N_7963,N_4891,N_4730);
nor U7964 (N_7964,N_5060,N_4874);
nand U7965 (N_7965,N_4362,N_4931);
or U7966 (N_7966,N_4613,N_4844);
nand U7967 (N_7967,N_5416,N_4223);
nand U7968 (N_7968,N_4955,N_4264);
or U7969 (N_7969,N_4055,N_5703);
nand U7970 (N_7970,N_4467,N_5292);
and U7971 (N_7971,N_5842,N_5066);
and U7972 (N_7972,N_4324,N_5817);
and U7973 (N_7973,N_5033,N_5690);
or U7974 (N_7974,N_4935,N_5166);
nor U7975 (N_7975,N_5500,N_5346);
or U7976 (N_7976,N_5426,N_5667);
nor U7977 (N_7977,N_5103,N_5496);
nor U7978 (N_7978,N_4395,N_5361);
nor U7979 (N_7979,N_5859,N_5610);
and U7980 (N_7980,N_5120,N_4351);
nor U7981 (N_7981,N_5042,N_4599);
nand U7982 (N_7982,N_4197,N_5242);
nand U7983 (N_7983,N_4550,N_4412);
and U7984 (N_7984,N_4437,N_4456);
and U7985 (N_7985,N_5901,N_5268);
nor U7986 (N_7986,N_5179,N_5399);
nand U7987 (N_7987,N_5268,N_5217);
nand U7988 (N_7988,N_5875,N_4880);
or U7989 (N_7989,N_4952,N_4689);
nor U7990 (N_7990,N_5080,N_5391);
or U7991 (N_7991,N_5917,N_5138);
nand U7992 (N_7992,N_5420,N_5669);
and U7993 (N_7993,N_5800,N_5390);
or U7994 (N_7994,N_4248,N_5791);
and U7995 (N_7995,N_4591,N_4681);
or U7996 (N_7996,N_4433,N_5157);
nand U7997 (N_7997,N_4557,N_5332);
nand U7998 (N_7998,N_5557,N_5643);
nor U7999 (N_7999,N_4921,N_4025);
nor U8000 (N_8000,N_7002,N_6044);
nor U8001 (N_8001,N_6667,N_6917);
nand U8002 (N_8002,N_6347,N_6449);
xor U8003 (N_8003,N_6642,N_7797);
xor U8004 (N_8004,N_7321,N_7165);
and U8005 (N_8005,N_7056,N_7956);
or U8006 (N_8006,N_7319,N_6016);
and U8007 (N_8007,N_7869,N_6930);
and U8008 (N_8008,N_7040,N_6839);
nand U8009 (N_8009,N_7825,N_7025);
nand U8010 (N_8010,N_7877,N_6544);
nor U8011 (N_8011,N_6268,N_6977);
nand U8012 (N_8012,N_7140,N_6180);
nor U8013 (N_8013,N_7172,N_6330);
nor U8014 (N_8014,N_6192,N_7324);
and U8015 (N_8015,N_6368,N_6351);
xnor U8016 (N_8016,N_7176,N_6688);
nor U8017 (N_8017,N_7828,N_6235);
or U8018 (N_8018,N_6836,N_7686);
nand U8019 (N_8019,N_6079,N_6286);
nand U8020 (N_8020,N_6003,N_7417);
nand U8021 (N_8021,N_6559,N_6308);
and U8022 (N_8022,N_6143,N_7382);
nor U8023 (N_8023,N_6628,N_6554);
nand U8024 (N_8024,N_6501,N_6035);
and U8025 (N_8025,N_6096,N_6332);
or U8026 (N_8026,N_7404,N_6461);
nor U8027 (N_8027,N_6526,N_7611);
or U8028 (N_8028,N_6965,N_6979);
or U8029 (N_8029,N_6795,N_6078);
nand U8030 (N_8030,N_7096,N_6209);
and U8031 (N_8031,N_6263,N_7383);
nand U8032 (N_8032,N_6104,N_6426);
nor U8033 (N_8033,N_7166,N_7440);
or U8034 (N_8034,N_6764,N_7352);
or U8035 (N_8035,N_6729,N_6592);
nand U8036 (N_8036,N_7816,N_7862);
nand U8037 (N_8037,N_6829,N_7203);
nor U8038 (N_8038,N_6799,N_6200);
nand U8039 (N_8039,N_7663,N_7568);
nor U8040 (N_8040,N_7334,N_7061);
or U8041 (N_8041,N_7708,N_6737);
nand U8042 (N_8042,N_6166,N_7488);
or U8043 (N_8043,N_7345,N_7895);
and U8044 (N_8044,N_6086,N_7831);
or U8045 (N_8045,N_6924,N_6512);
nand U8046 (N_8046,N_7270,N_6521);
nor U8047 (N_8047,N_6456,N_6144);
nand U8048 (N_8048,N_7048,N_7662);
nor U8049 (N_8049,N_7434,N_6099);
nand U8050 (N_8050,N_7150,N_7766);
or U8051 (N_8051,N_7433,N_7677);
nand U8052 (N_8052,N_6788,N_7067);
nand U8053 (N_8053,N_7667,N_6274);
or U8054 (N_8054,N_6430,N_7259);
or U8055 (N_8055,N_7944,N_6840);
or U8056 (N_8056,N_6303,N_7551);
nor U8057 (N_8057,N_7225,N_7521);
nor U8058 (N_8058,N_6478,N_6241);
nand U8059 (N_8059,N_7108,N_6765);
or U8060 (N_8060,N_7118,N_7999);
nand U8061 (N_8061,N_7156,N_7634);
nand U8062 (N_8062,N_7294,N_6606);
or U8063 (N_8063,N_7759,N_6171);
and U8064 (N_8064,N_6328,N_6157);
or U8065 (N_8065,N_6293,N_7757);
nand U8066 (N_8066,N_7720,N_6670);
or U8067 (N_8067,N_7325,N_7145);
and U8068 (N_8068,N_7137,N_7813);
nor U8069 (N_8069,N_6149,N_6355);
and U8070 (N_8070,N_7102,N_7457);
nand U8071 (N_8071,N_6348,N_7262);
nor U8072 (N_8072,N_7886,N_7028);
and U8073 (N_8073,N_7548,N_6111);
or U8074 (N_8074,N_7599,N_7798);
or U8075 (N_8075,N_6060,N_6307);
nand U8076 (N_8076,N_6946,N_7495);
nand U8077 (N_8077,N_6254,N_6847);
and U8078 (N_8078,N_6550,N_7550);
nand U8079 (N_8079,N_7251,N_7822);
xnor U8080 (N_8080,N_7955,N_6615);
or U8081 (N_8081,N_6784,N_6305);
and U8082 (N_8082,N_7498,N_7017);
nand U8083 (N_8083,N_6094,N_6383);
or U8084 (N_8084,N_7562,N_6363);
or U8085 (N_8085,N_6935,N_6122);
and U8086 (N_8086,N_6984,N_6871);
or U8087 (N_8087,N_6980,N_7763);
nand U8088 (N_8088,N_6433,N_7516);
and U8089 (N_8089,N_7504,N_6500);
nand U8090 (N_8090,N_6311,N_6830);
and U8091 (N_8091,N_6341,N_7748);
nor U8092 (N_8092,N_6580,N_7904);
or U8093 (N_8093,N_7399,N_6425);
or U8094 (N_8094,N_6561,N_7103);
nor U8095 (N_8095,N_7706,N_7094);
or U8096 (N_8096,N_6159,N_7384);
or U8097 (N_8097,N_7182,N_7450);
or U8098 (N_8098,N_7966,N_6174);
and U8099 (N_8099,N_7249,N_6443);
or U8100 (N_8100,N_6966,N_6732);
or U8101 (N_8101,N_6158,N_6712);
nand U8102 (N_8102,N_6813,N_7122);
or U8103 (N_8103,N_7778,N_7756);
and U8104 (N_8104,N_6922,N_7246);
or U8105 (N_8105,N_6611,N_7692);
nor U8106 (N_8106,N_7809,N_6806);
or U8107 (N_8107,N_7934,N_6523);
nor U8108 (N_8108,N_7059,N_7970);
or U8109 (N_8109,N_7962,N_6359);
nor U8110 (N_8110,N_6109,N_6066);
nand U8111 (N_8111,N_7728,N_6517);
xnor U8112 (N_8112,N_6023,N_7529);
nor U8113 (N_8113,N_6334,N_7295);
and U8114 (N_8114,N_6233,N_6413);
nor U8115 (N_8115,N_7731,N_6696);
nor U8116 (N_8116,N_7751,N_7189);
and U8117 (N_8117,N_7681,N_6375);
nand U8118 (N_8118,N_7930,N_7296);
nand U8119 (N_8119,N_7416,N_7605);
nand U8120 (N_8120,N_7774,N_7621);
nor U8121 (N_8121,N_6113,N_7051);
or U8122 (N_8122,N_7231,N_7979);
nand U8123 (N_8123,N_7049,N_7485);
or U8124 (N_8124,N_7771,N_7596);
or U8125 (N_8125,N_6976,N_7866);
and U8126 (N_8126,N_6914,N_6970);
or U8127 (N_8127,N_7707,N_6001);
and U8128 (N_8128,N_7694,N_6912);
nor U8129 (N_8129,N_7218,N_6895);
nand U8130 (N_8130,N_7491,N_6778);
nor U8131 (N_8131,N_6211,N_7330);
or U8132 (N_8132,N_6605,N_6154);
nor U8133 (N_8133,N_6119,N_7486);
and U8134 (N_8134,N_7467,N_6071);
or U8135 (N_8135,N_7147,N_6537);
nand U8136 (N_8136,N_6316,N_6578);
nor U8137 (N_8137,N_6193,N_7315);
nor U8138 (N_8138,N_7972,N_7777);
nand U8139 (N_8139,N_7060,N_6779);
or U8140 (N_8140,N_6740,N_6306);
nor U8141 (N_8141,N_7505,N_6748);
nor U8142 (N_8142,N_7331,N_6403);
and U8143 (N_8143,N_7957,N_6491);
nand U8144 (N_8144,N_7541,N_7524);
and U8145 (N_8145,N_7292,N_6089);
xor U8146 (N_8146,N_6596,N_7196);
or U8147 (N_8147,N_6133,N_6777);
and U8148 (N_8148,N_7187,N_6278);
nor U8149 (N_8149,N_7847,N_7312);
xnor U8150 (N_8150,N_7987,N_7205);
nand U8151 (N_8151,N_6487,N_6843);
nor U8152 (N_8152,N_7713,N_7607);
or U8153 (N_8153,N_6785,N_6655);
nand U8154 (N_8154,N_6088,N_6352);
and U8155 (N_8155,N_7046,N_6881);
nand U8156 (N_8156,N_6220,N_6898);
or U8157 (N_8157,N_6954,N_7159);
nand U8158 (N_8158,N_7938,N_6804);
nand U8159 (N_8159,N_6705,N_7650);
and U8160 (N_8160,N_7811,N_7202);
nand U8161 (N_8161,N_7597,N_7628);
and U8162 (N_8162,N_7685,N_6602);
nor U8163 (N_8163,N_6167,N_6195);
nor U8164 (N_8164,N_6480,N_7640);
nand U8165 (N_8165,N_7794,N_6736);
nand U8166 (N_8166,N_7229,N_6676);
nor U8167 (N_8167,N_6039,N_6470);
nor U8168 (N_8168,N_6369,N_6796);
and U8169 (N_8169,N_6107,N_7418);
nand U8170 (N_8170,N_7492,N_6128);
xnor U8171 (N_8171,N_7240,N_7919);
nor U8172 (N_8172,N_7965,N_7244);
or U8173 (N_8173,N_7690,N_6678);
or U8174 (N_8174,N_7552,N_7594);
or U8175 (N_8175,N_6838,N_7188);
and U8176 (N_8176,N_6029,N_6077);
nor U8177 (N_8177,N_6315,N_6072);
nor U8178 (N_8178,N_6477,N_6189);
or U8179 (N_8179,N_6656,N_7472);
nor U8180 (N_8180,N_6265,N_6995);
nor U8181 (N_8181,N_7958,N_6604);
and U8182 (N_8182,N_7378,N_7004);
nand U8183 (N_8183,N_7932,N_7887);
nand U8184 (N_8184,N_6713,N_7063);
nor U8185 (N_8185,N_7647,N_6693);
nor U8186 (N_8186,N_7081,N_6923);
nand U8187 (N_8187,N_6400,N_6774);
or U8188 (N_8188,N_7126,N_7307);
or U8189 (N_8189,N_7642,N_6673);
and U8190 (N_8190,N_6669,N_6026);
nand U8191 (N_8191,N_7793,N_7769);
nor U8192 (N_8192,N_7408,N_7986);
and U8193 (N_8193,N_6994,N_6885);
nor U8194 (N_8194,N_7925,N_6223);
nor U8195 (N_8195,N_6507,N_6474);
nand U8196 (N_8196,N_6882,N_7022);
nor U8197 (N_8197,N_7302,N_7554);
or U8198 (N_8198,N_7850,N_7781);
and U8199 (N_8199,N_7845,N_7380);
nand U8200 (N_8200,N_7304,N_7671);
nor U8201 (N_8201,N_7317,N_6878);
or U8202 (N_8202,N_7560,N_7035);
nor U8203 (N_8203,N_6279,N_6131);
nor U8204 (N_8204,N_7158,N_6992);
nor U8205 (N_8205,N_7990,N_7899);
or U8206 (N_8206,N_7186,N_6985);
nand U8207 (N_8207,N_7007,N_7608);
nor U8208 (N_8208,N_6273,N_7428);
nor U8209 (N_8209,N_6508,N_7803);
nand U8210 (N_8210,N_7726,N_7217);
or U8211 (N_8211,N_7574,N_6187);
nand U8212 (N_8212,N_6803,N_6962);
and U8213 (N_8213,N_7870,N_7837);
and U8214 (N_8214,N_6983,N_7897);
or U8215 (N_8215,N_6116,N_7752);
nand U8216 (N_8216,N_6731,N_7068);
xor U8217 (N_8217,N_7664,N_6218);
nand U8218 (N_8218,N_6668,N_7791);
nor U8219 (N_8219,N_6455,N_6793);
and U8220 (N_8220,N_6894,N_6841);
or U8221 (N_8221,N_7506,N_6152);
nor U8222 (N_8222,N_6753,N_6909);
nand U8223 (N_8223,N_6451,N_6130);
nand U8224 (N_8224,N_6025,N_6317);
nand U8225 (N_8225,N_7501,N_6548);
or U8226 (N_8226,N_7374,N_7687);
and U8227 (N_8227,N_7144,N_6190);
or U8228 (N_8228,N_6849,N_6468);
or U8229 (N_8229,N_7714,N_6744);
nor U8230 (N_8230,N_6565,N_6742);
nand U8231 (N_8231,N_6862,N_7660);
or U8232 (N_8232,N_6046,N_7442);
nor U8233 (N_8233,N_6627,N_6905);
or U8234 (N_8234,N_6476,N_6636);
nor U8235 (N_8235,N_6996,N_6951);
or U8236 (N_8236,N_6257,N_6340);
nor U8237 (N_8237,N_7168,N_7151);
xnor U8238 (N_8238,N_7026,N_7091);
or U8239 (N_8239,N_7271,N_6769);
nor U8240 (N_8240,N_6416,N_6019);
or U8241 (N_8241,N_6791,N_6529);
nor U8242 (N_8242,N_6665,N_6524);
and U8243 (N_8243,N_7132,N_6699);
and U8244 (N_8244,N_6350,N_7466);
and U8245 (N_8245,N_7518,N_7053);
and U8246 (N_8246,N_6084,N_6030);
nand U8247 (N_8247,N_7274,N_6835);
xnor U8248 (N_8248,N_7377,N_6250);
nor U8249 (N_8249,N_7092,N_7570);
or U8250 (N_8250,N_7609,N_6323);
nand U8251 (N_8251,N_7848,N_7015);
nand U8252 (N_8252,N_6267,N_7749);
and U8253 (N_8253,N_7572,N_7812);
nor U8254 (N_8254,N_6567,N_6423);
nand U8255 (N_8255,N_6011,N_7738);
and U8256 (N_8256,N_7849,N_7583);
nor U8257 (N_8257,N_7213,N_6822);
nor U8258 (N_8258,N_7426,N_7929);
or U8259 (N_8259,N_7859,N_6600);
nor U8260 (N_8260,N_6239,N_6421);
nand U8261 (N_8261,N_7148,N_7499);
or U8262 (N_8262,N_7358,N_7047);
nand U8263 (N_8263,N_7741,N_7942);
and U8264 (N_8264,N_7069,N_7475);
or U8265 (N_8265,N_7981,N_7914);
and U8266 (N_8266,N_6955,N_7030);
nor U8267 (N_8267,N_6420,N_6204);
or U8268 (N_8268,N_7306,N_6610);
or U8269 (N_8269,N_6182,N_7208);
nor U8270 (N_8270,N_7441,N_7299);
and U8271 (N_8271,N_7101,N_7890);
nand U8272 (N_8272,N_6199,N_6022);
nor U8273 (N_8273,N_6509,N_7398);
nor U8274 (N_8274,N_6063,N_6743);
or U8275 (N_8275,N_6690,N_7902);
or U8276 (N_8276,N_7127,N_7577);
nand U8277 (N_8277,N_6684,N_7160);
and U8278 (N_8278,N_6103,N_6043);
nor U8279 (N_8279,N_7489,N_7373);
nand U8280 (N_8280,N_6540,N_7697);
or U8281 (N_8281,N_7335,N_6772);
or U8282 (N_8282,N_7459,N_7376);
nand U8283 (N_8283,N_7547,N_6591);
and U8284 (N_8284,N_6762,N_7971);
and U8285 (N_8285,N_6815,N_6619);
nand U8286 (N_8286,N_7917,N_6272);
nand U8287 (N_8287,N_7242,N_6117);
and U8288 (N_8288,N_6963,N_7636);
xor U8289 (N_8289,N_6974,N_6380);
nor U8290 (N_8290,N_6302,N_7268);
nor U8291 (N_8291,N_7776,N_6597);
nor U8292 (N_8292,N_7194,N_7522);
nor U8293 (N_8293,N_7349,N_6042);
or U8294 (N_8294,N_6446,N_7922);
and U8295 (N_8295,N_6653,N_6502);
and U8296 (N_8296,N_7065,N_6296);
nor U8297 (N_8297,N_7273,N_6720);
nand U8298 (N_8298,N_7964,N_6018);
nor U8299 (N_8299,N_7832,N_7420);
or U8300 (N_8300,N_6041,N_6346);
nand U8301 (N_8301,N_6625,N_6313);
and U8302 (N_8302,N_7753,N_6014);
nand U8303 (N_8303,N_6747,N_6417);
and U8304 (N_8304,N_7629,N_6552);
nand U8305 (N_8305,N_7199,N_7689);
nor U8306 (N_8306,N_7107,N_6013);
or U8307 (N_8307,N_7410,N_6435);
and U8308 (N_8308,N_7834,N_6134);
nor U8309 (N_8309,N_7737,N_6297);
or U8310 (N_8310,N_7566,N_6343);
and U8311 (N_8311,N_7293,N_6698);
and U8312 (N_8312,N_7614,N_6718);
nand U8313 (N_8313,N_6920,N_6310);
or U8314 (N_8314,N_7604,N_6652);
or U8315 (N_8315,N_6728,N_7308);
nand U8316 (N_8316,N_7994,N_6087);
and U8317 (N_8317,N_6826,N_6759);
and U8318 (N_8318,N_6177,N_7314);
and U8319 (N_8319,N_6365,N_7645);
or U8320 (N_8320,N_6399,N_7054);
nor U8321 (N_8321,N_7393,N_6515);
nand U8322 (N_8322,N_7537,N_6719);
xor U8323 (N_8323,N_7874,N_7184);
and U8324 (N_8324,N_6854,N_7260);
nor U8325 (N_8325,N_6208,N_7180);
and U8326 (N_8326,N_6371,N_7672);
nand U8327 (N_8327,N_6427,N_6183);
xnor U8328 (N_8328,N_7588,N_6378);
nor U8329 (N_8329,N_6522,N_7333);
nand U8330 (N_8330,N_7531,N_7619);
nand U8331 (N_8331,N_6581,N_6110);
and U8332 (N_8332,N_7185,N_6738);
nand U8333 (N_8333,N_7950,N_7973);
nor U8334 (N_8334,N_6650,N_6339);
nand U8335 (N_8335,N_6138,N_7041);
nand U8336 (N_8336,N_6010,N_7578);
xnor U8337 (N_8337,N_7880,N_6216);
nand U8338 (N_8338,N_6875,N_7086);
and U8339 (N_8339,N_7646,N_6558);
or U8340 (N_8340,N_6880,N_6902);
xnor U8341 (N_8341,N_6292,N_7718);
nand U8342 (N_8342,N_7535,N_6201);
and U8343 (N_8343,N_6575,N_7412);
nand U8344 (N_8344,N_7206,N_6872);
nand U8345 (N_8345,N_7342,N_7354);
and U8346 (N_8346,N_6948,N_6533);
nand U8347 (N_8347,N_7590,N_6504);
nor U8348 (N_8348,N_6150,N_7882);
and U8349 (N_8349,N_7480,N_7712);
nand U8350 (N_8350,N_6938,N_7817);
and U8351 (N_8351,N_6800,N_6958);
nor U8352 (N_8352,N_6716,N_6687);
nor U8353 (N_8353,N_6739,N_7088);
nand U8354 (N_8354,N_6422,N_6635);
nor U8355 (N_8355,N_7425,N_6757);
or U8356 (N_8356,N_6374,N_7947);
or U8357 (N_8357,N_7290,N_6797);
xor U8358 (N_8358,N_7784,N_6879);
or U8359 (N_8359,N_6140,N_6842);
nor U8360 (N_8360,N_7497,N_6012);
nor U8361 (N_8361,N_6442,N_7370);
and U8362 (N_8362,N_6663,N_6768);
or U8363 (N_8363,N_7658,N_7077);
and U8364 (N_8364,N_6428,N_7487);
or U8365 (N_8365,N_7157,N_7111);
and U8366 (N_8366,N_7357,N_7744);
and U8367 (N_8367,N_6666,N_7563);
nor U8368 (N_8368,N_6844,N_6406);
and U8369 (N_8369,N_7214,N_7207);
nor U8370 (N_8370,N_7234,N_6452);
nor U8371 (N_8371,N_6252,N_7402);
or U8372 (N_8372,N_7238,N_7285);
nand U8373 (N_8373,N_6505,N_7451);
nor U8374 (N_8374,N_6741,N_7575);
nand U8375 (N_8375,N_6372,N_7204);
or U8376 (N_8376,N_7520,N_6322);
nand U8377 (N_8377,N_7746,N_7326);
or U8378 (N_8378,N_6899,N_6047);
or U8379 (N_8379,N_6217,N_6725);
or U8380 (N_8380,N_6531,N_7369);
nand U8381 (N_8381,N_6210,N_7009);
or U8382 (N_8382,N_7027,N_6485);
nor U8383 (N_8383,N_7036,N_6851);
and U8384 (N_8384,N_7722,N_7846);
nor U8385 (N_8385,N_7110,N_6593);
nand U8386 (N_8386,N_6934,N_6236);
or U8387 (N_8387,N_7097,N_6020);
or U8388 (N_8388,N_7643,N_7032);
nand U8389 (N_8389,N_6249,N_7037);
or U8390 (N_8390,N_7327,N_7826);
or U8391 (N_8391,N_7141,N_6703);
nor U8392 (N_8392,N_6142,N_6519);
or U8393 (N_8393,N_7641,N_6723);
nor U8394 (N_8394,N_6247,N_6711);
or U8395 (N_8395,N_7863,N_6021);
and U8396 (N_8396,N_7438,N_6486);
nor U8397 (N_8397,N_6919,N_7366);
or U8398 (N_8398,N_6562,N_7911);
or U8399 (N_8399,N_7988,N_7736);
nand U8400 (N_8400,N_6798,N_7682);
nand U8401 (N_8401,N_6601,N_6534);
nor U8402 (N_8402,N_6781,N_6694);
nand U8403 (N_8403,N_7875,N_6916);
and U8404 (N_8404,N_6516,N_6238);
or U8405 (N_8405,N_7221,N_6745);
nand U8406 (N_8406,N_6164,N_6633);
or U8407 (N_8407,N_7898,N_6364);
and U8408 (N_8408,N_6261,N_6891);
and U8409 (N_8409,N_6408,N_6493);
nand U8410 (N_8410,N_6545,N_7696);
and U8411 (N_8411,N_7571,N_6998);
nor U8412 (N_8412,N_7920,N_7070);
nand U8413 (N_8413,N_6821,N_7761);
and U8414 (N_8414,N_6270,N_7861);
or U8415 (N_8415,N_7719,N_7364);
nand U8416 (N_8416,N_7760,N_7567);
nand U8417 (N_8417,N_7545,N_6584);
or U8418 (N_8418,N_6145,N_7087);
or U8419 (N_8419,N_6255,N_6964);
and U8420 (N_8420,N_7183,N_6432);
nand U8421 (N_8421,N_7949,N_7638);
nand U8422 (N_8422,N_7691,N_7532);
nand U8423 (N_8423,N_7851,N_7134);
and U8424 (N_8424,N_7482,N_7673);
or U8425 (N_8425,N_6148,N_6527);
and U8426 (N_8426,N_6820,N_6212);
and U8427 (N_8427,N_6387,N_6587);
nor U8428 (N_8428,N_6132,N_7968);
and U8429 (N_8429,N_6483,N_7976);
and U8430 (N_8430,N_6860,N_6214);
and U8431 (N_8431,N_6287,N_6385);
nor U8432 (N_8432,N_7732,N_6224);
or U8433 (N_8433,N_7842,N_6620);
and U8434 (N_8434,N_6395,N_7549);
nand U8435 (N_8435,N_6194,N_7359);
nor U8436 (N_8436,N_6049,N_6412);
nand U8437 (N_8437,N_6867,N_6717);
nor U8438 (N_8438,N_7622,N_6528);
or U8439 (N_8439,N_7743,N_7980);
or U8440 (N_8440,N_7616,N_6931);
or U8441 (N_8441,N_6300,N_7050);
and U8442 (N_8442,N_7998,N_7569);
and U8443 (N_8443,N_6623,N_6576);
and U8444 (N_8444,N_6950,N_7795);
nor U8445 (N_8445,N_6925,N_6513);
or U8446 (N_8446,N_7387,N_7885);
or U8447 (N_8447,N_7449,N_7951);
nand U8448 (N_8448,N_7912,N_7178);
or U8449 (N_8449,N_6248,N_7265);
nand U8450 (N_8450,N_6076,N_7654);
nor U8451 (N_8451,N_7693,N_6543);
and U8452 (N_8452,N_7173,N_6004);
and U8453 (N_8453,N_7235,N_6392);
nor U8454 (N_8454,N_7220,N_6680);
and U8455 (N_8455,N_7106,N_6884);
and U8456 (N_8456,N_7508,N_6038);
nor U8457 (N_8457,N_7799,N_7833);
and U8458 (N_8458,N_7534,N_6975);
nor U8459 (N_8459,N_7635,N_7927);
nor U8460 (N_8460,N_7695,N_6921);
nor U8461 (N_8461,N_6952,N_7099);
and U8462 (N_8462,N_6358,N_6271);
nor U8463 (N_8463,N_7724,N_7598);
and U8464 (N_8464,N_7043,N_6579);
and U8465 (N_8465,N_7509,N_6608);
nand U8466 (N_8466,N_7666,N_6506);
and U8467 (N_8467,N_6634,N_7000);
or U8468 (N_8468,N_6034,N_7700);
xnor U8469 (N_8469,N_6402,N_6689);
or U8470 (N_8470,N_6092,N_6118);
nor U8471 (N_8471,N_6730,N_7940);
nand U8472 (N_8472,N_7789,N_7034);
and U8473 (N_8473,N_7513,N_6818);
and U8474 (N_8474,N_6002,N_6091);
nand U8475 (N_8475,N_7083,N_7227);
nor U8476 (N_8476,N_6161,N_6649);
or U8477 (N_8477,N_7125,N_6203);
and U8478 (N_8478,N_7627,N_6221);
or U8479 (N_8479,N_7767,N_7360);
nand U8480 (N_8480,N_7142,N_7517);
or U8481 (N_8481,N_7062,N_7512);
nand U8482 (N_8482,N_7171,N_7379);
nor U8483 (N_8483,N_6646,N_7908);
xor U8484 (N_8484,N_7044,N_7602);
or U8485 (N_8485,N_6658,N_6176);
and U8486 (N_8486,N_7889,N_6651);
nand U8487 (N_8487,N_6632,N_6081);
or U8488 (N_8488,N_6932,N_7507);
nor U8489 (N_8489,N_7630,N_6342);
nand U8490 (N_8490,N_6431,N_7372);
nor U8491 (N_8491,N_7786,N_6890);
nand U8492 (N_8492,N_6647,N_6051);
nor U8493 (N_8493,N_6953,N_6848);
nand U8494 (N_8494,N_7779,N_7936);
or U8495 (N_8495,N_6398,N_7406);
or U8496 (N_8496,N_7288,N_7283);
nor U8497 (N_8497,N_7910,N_7511);
nor U8498 (N_8498,N_6546,N_6957);
and U8499 (N_8499,N_7765,N_7256);
or U8500 (N_8500,N_6481,N_7624);
nand U8501 (N_8501,N_6105,N_6868);
nor U8502 (N_8502,N_6767,N_6956);
nand U8503 (N_8503,N_6594,N_7903);
and U8504 (N_8504,N_6572,N_6626);
nor U8505 (N_8505,N_7775,N_6404);
nand U8506 (N_8506,N_7371,N_6458);
and U8507 (N_8507,N_7403,N_6234);
and U8508 (N_8508,N_7414,N_6484);
and U8509 (N_8509,N_6379,N_7075);
nand U8510 (N_8510,N_6609,N_6197);
nand U8511 (N_8511,N_7014,N_7353);
nand U8512 (N_8512,N_7395,N_7704);
nor U8513 (N_8513,N_7072,N_6373);
and U8514 (N_8514,N_7432,N_6345);
or U8515 (N_8515,N_7252,N_7446);
nor U8516 (N_8516,N_7237,N_7670);
or U8517 (N_8517,N_6661,N_7592);
nor U8518 (N_8518,N_6999,N_7858);
nor U8519 (N_8519,N_7129,N_7867);
and U8520 (N_8520,N_6864,N_6169);
and U8521 (N_8521,N_7444,N_7287);
and U8522 (N_8522,N_6771,N_7679);
and U8523 (N_8523,N_6457,N_7282);
nor U8524 (N_8524,N_7362,N_6291);
and U8525 (N_8525,N_6571,N_7823);
and U8526 (N_8526,N_6008,N_7465);
and U8527 (N_8527,N_6959,N_7210);
or U8528 (N_8528,N_6944,N_7526);
nor U8529 (N_8529,N_6052,N_7909);
nand U8530 (N_8530,N_6541,N_7601);
or U8531 (N_8531,N_6473,N_6389);
nor U8532 (N_8532,N_6454,N_7595);
and U8533 (N_8533,N_6036,N_7033);
nand U8534 (N_8534,N_6410,N_7280);
nor U8535 (N_8535,N_6945,N_7711);
nand U8536 (N_8536,N_6419,N_6863);
nand U8537 (N_8537,N_7104,N_7853);
nand U8538 (N_8538,N_6928,N_7525);
or U8539 (N_8539,N_7281,N_6463);
and U8540 (N_8540,N_6941,N_7461);
nor U8541 (N_8541,N_7580,N_6028);
and U8542 (N_8542,N_7723,N_7742);
and U8543 (N_8543,N_6045,N_7478);
and U8544 (N_8544,N_6436,N_6637);
nand U8545 (N_8545,N_7381,N_6536);
nor U8546 (N_8546,N_6391,N_7161);
or U8547 (N_8547,N_7143,N_6377);
and U8548 (N_8548,N_6048,N_6459);
or U8549 (N_8549,N_6775,N_7329);
or U8550 (N_8550,N_6082,N_6735);
or U8551 (N_8551,N_6095,N_7703);
and U8552 (N_8552,N_6429,N_7818);
nand U8553 (N_8553,N_6942,N_7785);
nand U8554 (N_8554,N_7284,N_7012);
nor U8555 (N_8555,N_6870,N_7452);
or U8556 (N_8556,N_7836,N_6275);
and U8557 (N_8557,N_7538,N_6547);
nor U8558 (N_8558,N_7248,N_7123);
nor U8559 (N_8559,N_7209,N_7298);
nand U8560 (N_8560,N_6907,N_7768);
nor U8561 (N_8561,N_6846,N_6589);
xnor U8562 (N_8562,N_7100,N_7883);
nor U8563 (N_8563,N_6629,N_7992);
or U8564 (N_8564,N_7350,N_6136);
nand U8565 (N_8565,N_6370,N_6031);
nand U8566 (N_8566,N_7631,N_7310);
nor U8567 (N_8567,N_6721,N_7829);
nor U8568 (N_8568,N_7409,N_7576);
nand U8569 (N_8569,N_7510,N_7540);
and U8570 (N_8570,N_7612,N_6242);
nand U8571 (N_8571,N_7215,N_7303);
nand U8572 (N_8572,N_6494,N_7709);
nand U8573 (N_8573,N_6009,N_7328);
nand U8574 (N_8574,N_7445,N_6856);
and U8575 (N_8575,N_6222,N_7219);
or U8576 (N_8576,N_6993,N_6763);
and U8577 (N_8577,N_6067,N_6827);
nor U8578 (N_8578,N_6915,N_7239);
nand U8579 (N_8579,N_6691,N_6490);
or U8580 (N_8580,N_6102,N_7253);
or U8581 (N_8581,N_6978,N_7772);
xnor U8582 (N_8582,N_7436,N_7336);
and U8583 (N_8583,N_7163,N_7937);
nor U8584 (N_8584,N_6237,N_6243);
or U8585 (N_8585,N_6754,N_6695);
nor U8586 (N_8586,N_6756,N_6850);
or U8587 (N_8587,N_7959,N_7814);
and U8588 (N_8588,N_7705,N_7476);
and U8589 (N_8589,N_6075,N_7146);
nand U8590 (N_8590,N_6603,N_6886);
and U8591 (N_8591,N_7250,N_7637);
nand U8592 (N_8592,N_6384,N_7275);
and U8593 (N_8593,N_6556,N_6289);
nand U8594 (N_8594,N_6288,N_7984);
or U8595 (N_8595,N_6000,N_7080);
nor U8596 (N_8596,N_7128,N_7543);
nor U8597 (N_8597,N_7906,N_6298);
or U8598 (N_8598,N_6497,N_6645);
nand U8599 (N_8599,N_6196,N_6825);
nand U8600 (N_8600,N_7727,N_7933);
or U8601 (N_8601,N_6496,N_6582);
and U8602 (N_8602,N_7857,N_6151);
or U8603 (N_8603,N_7796,N_7190);
and U8604 (N_8604,N_6624,N_7721);
nand U8605 (N_8605,N_6901,N_7977);
or U8606 (N_8606,N_7931,N_7233);
and U8607 (N_8607,N_7783,N_7052);
nand U8608 (N_8608,N_6943,N_7230);
and U8609 (N_8609,N_6755,N_6225);
nand U8610 (N_8610,N_6641,N_7071);
nand U8611 (N_8611,N_6024,N_7808);
nor U8612 (N_8612,N_6097,N_6285);
nand U8613 (N_8613,N_7559,N_7341);
and U8614 (N_8614,N_7415,N_6281);
nand U8615 (N_8615,N_7021,N_7820);
xor U8616 (N_8616,N_6733,N_6697);
and U8617 (N_8617,N_7801,N_7264);
nand U8618 (N_8618,N_7243,N_6904);
or U8619 (N_8619,N_6617,N_6861);
nand U8620 (N_8620,N_6178,N_7730);
and U8621 (N_8621,N_6033,N_7355);
and U8622 (N_8622,N_7391,N_6479);
or U8623 (N_8623,N_6990,N_7089);
nor U8624 (N_8624,N_6276,N_6361);
or U8625 (N_8625,N_7558,N_7587);
or U8626 (N_8626,N_7453,N_6206);
nor U8627 (N_8627,N_7995,N_6682);
nor U8628 (N_8628,N_7892,N_6112);
nor U8629 (N_8629,N_6664,N_7493);
nand U8630 (N_8630,N_7193,N_6654);
nor U8631 (N_8631,N_7266,N_6269);
nand U8632 (N_8632,N_7437,N_7905);
and U8633 (N_8633,N_6414,N_6514);
nor U8634 (N_8634,N_6677,N_7945);
nor U8635 (N_8635,N_6518,N_6939);
nand U8636 (N_8636,N_7115,N_6318);
or U8637 (N_8637,N_6356,N_6453);
or U8638 (N_8638,N_6814,N_6124);
and U8639 (N_8639,N_6349,N_7468);
and U8640 (N_8640,N_7878,N_6790);
nand U8641 (N_8641,N_7388,N_7807);
or U8642 (N_8642,N_7119,N_7201);
or U8643 (N_8643,N_7278,N_7347);
or U8644 (N_8644,N_7439,N_7011);
and U8645 (N_8645,N_6489,N_6590);
nand U8646 (N_8646,N_6734,N_7573);
nor U8647 (N_8647,N_7039,N_6277);
nor U8648 (N_8648,N_6007,N_7456);
nor U8649 (N_8649,N_6253,N_6256);
or U8650 (N_8650,N_6761,N_6900);
nand U8651 (N_8651,N_6325,N_7610);
and U8652 (N_8652,N_6244,N_6153);
nand U8653 (N_8653,N_6444,N_6466);
xor U8654 (N_8654,N_6498,N_7997);
or U8655 (N_8655,N_6750,N_6202);
nand U8656 (N_8656,N_7322,N_7013);
nand U8657 (N_8657,N_6724,N_7473);
nand U8658 (N_8658,N_7952,N_6640);
and U8659 (N_8659,N_7149,N_6816);
or U8660 (N_8660,N_7815,N_6810);
and U8661 (N_8661,N_7291,N_7443);
and U8662 (N_8662,N_7699,N_6709);
nor U8663 (N_8663,N_7582,N_6525);
nand U8664 (N_8664,N_6588,N_6040);
or U8665 (N_8665,N_7954,N_7332);
nor U8666 (N_8666,N_7989,N_6437);
and U8667 (N_8667,N_6309,N_6061);
and U8668 (N_8668,N_7536,N_6050);
and U8669 (N_8669,N_6053,N_7297);
and U8670 (N_8670,N_6539,N_6859);
and U8671 (N_8671,N_6090,N_7561);
or U8672 (N_8672,N_6708,N_7320);
xnor U8673 (N_8673,N_7477,N_7527);
nand U8674 (N_8674,N_6568,N_6564);
nand U8675 (N_8675,N_6937,N_7975);
nor U8676 (N_8676,N_6168,N_7197);
nor U8677 (N_8677,N_7124,N_6336);
nor U8678 (N_8678,N_7553,N_7093);
nor U8679 (N_8679,N_6127,N_6170);
nor U8680 (N_8680,N_7113,N_6129);
nor U8681 (N_8681,N_7788,N_7716);
nor U8682 (N_8682,N_7167,N_7479);
nor U8683 (N_8683,N_7935,N_7891);
and U8684 (N_8684,N_7460,N_6520);
nand U8685 (N_8685,N_7121,N_6396);
and U8686 (N_8686,N_7212,N_7195);
nor U8687 (N_8687,N_7138,N_7868);
nand U8688 (N_8688,N_7978,N_7620);
or U8689 (N_8689,N_6982,N_7871);
or U8690 (N_8690,N_7745,N_7164);
nand U8691 (N_8691,N_6929,N_7963);
nand U8692 (N_8692,N_7135,N_6331);
and U8693 (N_8693,N_7983,N_6064);
or U8694 (N_8694,N_6405,N_7055);
nand U8695 (N_8695,N_7073,N_7066);
nor U8696 (N_8696,N_7114,N_7279);
or U8697 (N_8697,N_6376,N_7985);
or U8698 (N_8698,N_7579,N_7514);
nand U8699 (N_8699,N_6123,N_6877);
nand U8700 (N_8700,N_6971,N_7819);
nor U8701 (N_8701,N_7133,N_7356);
nand U8702 (N_8702,N_7269,N_7683);
xnor U8703 (N_8703,N_7057,N_7245);
or U8704 (N_8704,N_6911,N_7533);
or U8705 (N_8705,N_7764,N_6787);
nor U8706 (N_8706,N_7076,N_6918);
and U8707 (N_8707,N_6227,N_7918);
and U8708 (N_8708,N_6616,N_6100);
and U8709 (N_8709,N_6475,N_7023);
or U8710 (N_8710,N_6801,N_7351);
nor U8711 (N_8711,N_6366,N_7623);
nor U8712 (N_8712,N_6284,N_6445);
nand U8713 (N_8713,N_7780,N_7702);
or U8714 (N_8714,N_7411,N_7338);
nor U8715 (N_8715,N_7386,N_7471);
nand U8716 (N_8716,N_7755,N_6353);
and U8717 (N_8717,N_7651,N_6295);
and U8718 (N_8718,N_7960,N_6988);
nor U8719 (N_8719,N_6231,N_7045);
nand U8720 (N_8720,N_6424,N_6290);
nor U8721 (N_8721,N_7112,N_6973);
nor U8722 (N_8722,N_7675,N_6710);
and U8723 (N_8723,N_6335,N_6262);
nor U8724 (N_8724,N_7309,N_6940);
nor U8725 (N_8725,N_6354,N_7078);
nand U8726 (N_8726,N_7996,N_6726);
and U8727 (N_8727,N_7120,N_7018);
nand U8728 (N_8728,N_7873,N_6447);
nor U8729 (N_8729,N_7515,N_7669);
or U8730 (N_8730,N_7003,N_6773);
nor U8731 (N_8731,N_6439,N_6648);
nand U8732 (N_8732,N_7928,N_6855);
nand U8733 (N_8733,N_6685,N_6229);
or U8734 (N_8734,N_6344,N_6324);
or U8735 (N_8735,N_6314,N_7413);
nor U8736 (N_8736,N_7407,N_6776);
nand U8737 (N_8737,N_7668,N_6852);
and U8738 (N_8738,N_7435,N_6037);
nor U8739 (N_8739,N_6440,N_6809);
and U8740 (N_8740,N_6327,N_7943);
nor U8741 (N_8741,N_7729,N_6073);
and U8742 (N_8742,N_6304,N_7154);
nor U8743 (N_8743,N_7169,N_7649);
xor U8744 (N_8744,N_6228,N_7656);
and U8745 (N_8745,N_7152,N_7688);
or U8746 (N_8746,N_6367,N_6865);
nor U8747 (N_8747,N_6933,N_7019);
or U8748 (N_8748,N_7802,N_7661);
nor U8749 (N_8749,N_7484,N_7361);
nand U8750 (N_8750,N_6936,N_6819);
nand U8751 (N_8751,N_6357,N_6409);
or U8752 (N_8752,N_6910,N_7613);
xor U8753 (N_8753,N_6833,N_6215);
nand U8754 (N_8754,N_6070,N_7734);
and U8755 (N_8755,N_7464,N_7375);
or U8756 (N_8756,N_7228,N_6782);
nor U8757 (N_8757,N_6823,N_6246);
nand U8758 (N_8758,N_7657,N_7008);
nand U8759 (N_8759,N_6059,N_7644);
nor U8760 (N_8760,N_6282,N_7830);
and U8761 (N_8761,N_6837,N_7430);
nor U8762 (N_8762,N_7519,N_6598);
or U8763 (N_8763,N_7200,N_7855);
nor U8764 (N_8764,N_7915,N_6326);
nand U8765 (N_8765,N_7539,N_7429);
and U8766 (N_8766,N_6160,N_7029);
and U8767 (N_8767,N_6692,N_7961);
or U8768 (N_8768,N_6986,N_6949);
nor U8769 (N_8769,N_6382,N_6831);
and U8770 (N_8770,N_6511,N_7770);
and U8771 (N_8771,N_7969,N_7827);
and U8772 (N_8772,N_7463,N_7226);
and U8773 (N_8773,N_6114,N_7844);
and U8774 (N_8774,N_6989,N_6093);
nor U8775 (N_8775,N_6613,N_6542);
and U8776 (N_8776,N_7625,N_6961);
and U8777 (N_8777,N_7923,N_7085);
and U8778 (N_8778,N_7838,N_6488);
or U8779 (N_8779,N_6106,N_6824);
and U8780 (N_8780,N_7105,N_7606);
or U8781 (N_8781,N_7710,N_7006);
nand U8782 (N_8782,N_6139,N_7872);
nand U8783 (N_8783,N_6770,N_7901);
nand U8784 (N_8784,N_6394,N_6245);
nand U8785 (N_8785,N_6069,N_7401);
and U8786 (N_8786,N_6621,N_6469);
nor U8787 (N_8787,N_7841,N_7924);
or U8788 (N_8788,N_6553,N_7633);
nand U8789 (N_8789,N_6101,N_7258);
nor U8790 (N_8790,N_7876,N_7787);
nand U8791 (N_8791,N_7762,N_7216);
or U8792 (N_8792,N_7618,N_7805);
or U8793 (N_8793,N_6622,N_7544);
and U8794 (N_8794,N_7286,N_6438);
and U8795 (N_8795,N_6700,N_7339);
and U8796 (N_8796,N_6492,N_7301);
xor U8797 (N_8797,N_7941,N_7530);
nor U8798 (N_8798,N_6845,N_6555);
nor U8799 (N_8799,N_6251,N_7323);
nand U8800 (N_8800,N_7198,N_7939);
and U8801 (N_8801,N_6121,N_6172);
nor U8802 (N_8802,N_6896,N_6599);
nand U8803 (N_8803,N_6173,N_7864);
or U8804 (N_8804,N_7313,N_7680);
nand U8805 (N_8805,N_6866,N_6532);
nand U8806 (N_8806,N_7031,N_6972);
nand U8807 (N_8807,N_6362,N_6991);
and U8808 (N_8808,N_7272,N_6460);
or U8809 (N_8809,N_7632,N_6260);
and U8810 (N_8810,N_6175,N_7900);
nor U8811 (N_8811,N_6147,N_6704);
and U8812 (N_8812,N_6706,N_6969);
nor U8813 (N_8813,N_7241,N_7800);
nor U8814 (N_8814,N_6085,N_6015);
and U8815 (N_8815,N_6686,N_6098);
nand U8816 (N_8816,N_7589,N_6997);
nor U8817 (N_8817,N_7698,N_6657);
and U8818 (N_8818,N_6397,N_7318);
nand U8819 (N_8819,N_6163,N_7346);
nor U8820 (N_8820,N_7603,N_6115);
and U8821 (N_8821,N_7750,N_7181);
and U8822 (N_8822,N_7139,N_7153);
and U8823 (N_8823,N_6570,N_6137);
nor U8824 (N_8824,N_7340,N_7392);
and U8825 (N_8825,N_7170,N_6415);
nor U8826 (N_8826,N_6464,N_6472);
or U8827 (N_8827,N_6557,N_7542);
nand U8828 (N_8828,N_6141,N_6301);
nand U8829 (N_8829,N_7894,N_6560);
nand U8830 (N_8830,N_6401,N_6643);
or U8831 (N_8831,N_7179,N_6530);
nor U8832 (N_8832,N_7136,N_7617);
or U8833 (N_8833,N_7454,N_7343);
xnor U8834 (N_8834,N_6538,N_6585);
and U8835 (N_8835,N_6630,N_7879);
or U8836 (N_8836,N_6817,N_6727);
or U8837 (N_8837,N_7337,N_7907);
or U8838 (N_8838,N_6614,N_7503);
and U8839 (N_8839,N_7397,N_7733);
nand U8840 (N_8840,N_6889,N_7064);
or U8841 (N_8841,N_7316,N_7095);
or U8842 (N_8842,N_6566,N_6126);
and U8843 (N_8843,N_7222,N_6802);
or U8844 (N_8844,N_7648,N_7192);
and U8845 (N_8845,N_7474,N_6068);
nand U8846 (N_8846,N_6662,N_6056);
and U8847 (N_8847,N_6108,N_7946);
nor U8848 (N_8848,N_6135,N_6120);
or U8849 (N_8849,N_6549,N_6874);
nor U8850 (N_8850,N_7289,N_6672);
nor U8851 (N_8851,N_7852,N_7223);
and U8852 (N_8852,N_7058,N_7773);
and U8853 (N_8853,N_6563,N_7305);
nor U8854 (N_8854,N_7276,N_7839);
and U8855 (N_8855,N_7117,N_7020);
nor U8856 (N_8856,N_7565,N_6407);
nor U8857 (N_8857,N_7639,N_7394);
or U8858 (N_8858,N_6503,N_7458);
nand U8859 (N_8859,N_7747,N_6230);
and U8860 (N_8860,N_6390,N_6381);
nor U8861 (N_8861,N_6179,N_7735);
and U8862 (N_8862,N_6683,N_6834);
nand U8863 (N_8863,N_7348,N_7109);
and U8864 (N_8864,N_7255,N_7896);
or U8865 (N_8865,N_7790,N_6450);
nor U8866 (N_8866,N_6005,N_6805);
nand U8867 (N_8867,N_6055,N_6057);
and U8868 (N_8868,N_6156,N_7481);
nand U8869 (N_8869,N_6908,N_7840);
and U8870 (N_8870,N_6722,N_7177);
and U8871 (N_8871,N_7422,N_7701);
nor U8872 (N_8872,N_7191,N_6388);
nor U8873 (N_8873,N_6465,N_6551);
nor U8874 (N_8874,N_6660,N_6360);
and U8875 (N_8875,N_6857,N_6612);
and U8876 (N_8876,N_6766,N_6054);
and U8877 (N_8877,N_7674,N_7615);
nand U8878 (N_8878,N_6510,N_7038);
xor U8879 (N_8879,N_7131,N_6319);
or U8880 (N_8880,N_7993,N_7396);
or U8881 (N_8881,N_7782,N_6639);
and U8882 (N_8882,N_7528,N_7653);
nor U8883 (N_8883,N_6967,N_6947);
nand U8884 (N_8884,N_7921,N_6259);
and U8885 (N_8885,N_7300,N_7005);
or U8886 (N_8886,N_6411,N_6499);
nand U8887 (N_8887,N_6674,N_6240);
or U8888 (N_8888,N_7854,N_7974);
or U8889 (N_8889,N_6618,N_7421);
and U8890 (N_8890,N_6577,N_7754);
nor U8891 (N_8891,N_7257,N_6906);
and U8892 (N_8892,N_6583,N_6968);
and U8893 (N_8893,N_6329,N_7174);
nand U8894 (N_8894,N_7843,N_7470);
nand U8895 (N_8895,N_7490,N_6760);
nand U8896 (N_8896,N_6573,N_7431);
or U8897 (N_8897,N_6006,N_6780);
and U8898 (N_8898,N_7725,N_6752);
or U8899 (N_8899,N_7684,N_7090);
or U8900 (N_8900,N_7835,N_7804);
and U8901 (N_8901,N_6926,N_6294);
and U8902 (N_8902,N_7079,N_6981);
or U8903 (N_8903,N_7496,N_6675);
nand U8904 (N_8904,N_7363,N_6715);
nor U8905 (N_8905,N_7311,N_7913);
or U8906 (N_8906,N_7042,N_6207);
nor U8907 (N_8907,N_6333,N_6751);
and U8908 (N_8908,N_7389,N_6017);
xor U8909 (N_8909,N_6858,N_6574);
nand U8910 (N_8910,N_7739,N_6812);
and U8911 (N_8911,N_6280,N_7232);
nand U8912 (N_8912,N_6679,N_7130);
nand U8913 (N_8913,N_6337,N_6595);
nand U8914 (N_8914,N_6320,N_6569);
or U8915 (N_8915,N_7884,N_7888);
and U8916 (N_8916,N_6876,N_7483);
or U8917 (N_8917,N_7856,N_6707);
nand U8918 (N_8918,N_6258,N_6644);
and U8919 (N_8919,N_6746,N_7556);
nand U8920 (N_8920,N_7224,N_6903);
or U8921 (N_8921,N_7016,N_7263);
or U8922 (N_8922,N_6434,N_7405);
nor U8923 (N_8923,N_7792,N_6146);
nor U8924 (N_8924,N_7455,N_7715);
or U8925 (N_8925,N_7821,N_7098);
or U8926 (N_8926,N_7584,N_7365);
or U8927 (N_8927,N_6828,N_7344);
nand U8928 (N_8928,N_7267,N_7581);
or U8929 (N_8929,N_7010,N_7400);
or U8930 (N_8930,N_7678,N_7074);
and U8931 (N_8931,N_7591,N_6832);
or U8932 (N_8932,N_6188,N_6758);
and U8933 (N_8933,N_6266,N_6631);
or U8934 (N_8934,N_7236,N_6058);
and U8935 (N_8935,N_6226,N_7564);
or U8936 (N_8936,N_7865,N_7655);
nor U8937 (N_8937,N_6960,N_6165);
nor U8938 (N_8938,N_6264,N_6065);
and U8939 (N_8939,N_6074,N_7368);
nor U8940 (N_8940,N_7390,N_6080);
nand U8941 (N_8941,N_6792,N_6386);
xnor U8942 (N_8942,N_7424,N_7419);
or U8943 (N_8943,N_6893,N_6027);
nand U8944 (N_8944,N_7948,N_7557);
or U8945 (N_8945,N_7447,N_6219);
or U8946 (N_8946,N_6032,N_6987);
nor U8947 (N_8947,N_7717,N_6794);
and U8948 (N_8948,N_6299,N_6659);
nand U8949 (N_8949,N_6681,N_6853);
or U8950 (N_8950,N_7953,N_7893);
nor U8951 (N_8951,N_6155,N_6185);
nand U8952 (N_8952,N_6714,N_7600);
nor U8953 (N_8953,N_7626,N_6807);
or U8954 (N_8954,N_6198,N_7967);
and U8955 (N_8955,N_7502,N_6448);
nand U8956 (N_8956,N_7494,N_6062);
and U8957 (N_8957,N_7676,N_7586);
or U8958 (N_8958,N_6913,N_6883);
and U8959 (N_8959,N_6638,N_6671);
nor U8960 (N_8960,N_6213,N_7175);
and U8961 (N_8961,N_6471,N_7758);
and U8962 (N_8962,N_6888,N_6312);
nand U8963 (N_8963,N_7991,N_7427);
or U8964 (N_8964,N_7555,N_6789);
nand U8965 (N_8965,N_6184,N_7001);
or U8966 (N_8966,N_6125,N_7881);
and U8967 (N_8967,N_6892,N_6181);
and U8968 (N_8968,N_7247,N_7593);
nand U8969 (N_8969,N_6418,N_6749);
nand U8970 (N_8970,N_7810,N_7254);
nand U8971 (N_8971,N_6873,N_6338);
and U8972 (N_8972,N_7806,N_6786);
or U8973 (N_8973,N_6162,N_7367);
nand U8974 (N_8974,N_7162,N_7448);
nor U8975 (N_8975,N_7740,N_6495);
nand U8976 (N_8976,N_6927,N_7155);
nand U8977 (N_8977,N_7211,N_7082);
or U8978 (N_8978,N_6441,N_7261);
nand U8979 (N_8979,N_7500,N_6467);
nand U8980 (N_8980,N_7982,N_7277);
and U8981 (N_8981,N_6783,N_6535);
or U8982 (N_8982,N_7665,N_6205);
and U8983 (N_8983,N_7546,N_7423);
and U8984 (N_8984,N_6607,N_7659);
nand U8985 (N_8985,N_6887,N_7860);
nor U8986 (N_8986,N_7084,N_6283);
or U8987 (N_8987,N_6586,N_7469);
nor U8988 (N_8988,N_7385,N_6897);
nor U8989 (N_8989,N_6083,N_6232);
xor U8990 (N_8990,N_7585,N_7926);
nor U8991 (N_8991,N_7024,N_6811);
nand U8992 (N_8992,N_6808,N_7652);
or U8993 (N_8993,N_6186,N_6702);
nand U8994 (N_8994,N_6482,N_7462);
nor U8995 (N_8995,N_6191,N_7523);
nor U8996 (N_8996,N_6321,N_6462);
or U8997 (N_8997,N_7824,N_7116);
and U8998 (N_8998,N_6701,N_6869);
nor U8999 (N_8999,N_6393,N_7916);
nand U9000 (N_9000,N_7148,N_6536);
nand U9001 (N_9001,N_7953,N_6972);
nand U9002 (N_9002,N_6386,N_7077);
nand U9003 (N_9003,N_7207,N_7596);
nor U9004 (N_9004,N_6064,N_7049);
nand U9005 (N_9005,N_7255,N_7100);
nor U9006 (N_9006,N_6403,N_7336);
nand U9007 (N_9007,N_6334,N_6595);
nand U9008 (N_9008,N_7974,N_7696);
nor U9009 (N_9009,N_6373,N_6284);
and U9010 (N_9010,N_6473,N_7271);
nor U9011 (N_9011,N_7465,N_7530);
nand U9012 (N_9012,N_6424,N_7195);
xor U9013 (N_9013,N_6021,N_7105);
nor U9014 (N_9014,N_7043,N_6564);
nor U9015 (N_9015,N_6884,N_7085);
xnor U9016 (N_9016,N_7346,N_6942);
nor U9017 (N_9017,N_7056,N_6569);
xor U9018 (N_9018,N_6451,N_7442);
xor U9019 (N_9019,N_7127,N_6686);
and U9020 (N_9020,N_7396,N_7855);
or U9021 (N_9021,N_6669,N_6374);
nor U9022 (N_9022,N_6441,N_7036);
nand U9023 (N_9023,N_7736,N_6389);
or U9024 (N_9024,N_6154,N_7151);
nand U9025 (N_9025,N_6219,N_7282);
and U9026 (N_9026,N_7460,N_6247);
nand U9027 (N_9027,N_6121,N_7639);
nand U9028 (N_9028,N_7132,N_7435);
or U9029 (N_9029,N_7643,N_7468);
and U9030 (N_9030,N_7149,N_7898);
nor U9031 (N_9031,N_6383,N_6528);
nand U9032 (N_9032,N_6178,N_6052);
and U9033 (N_9033,N_7262,N_6752);
nor U9034 (N_9034,N_7152,N_6335);
and U9035 (N_9035,N_7187,N_6800);
or U9036 (N_9036,N_7531,N_6854);
nor U9037 (N_9037,N_6493,N_7649);
or U9038 (N_9038,N_7459,N_7983);
or U9039 (N_9039,N_6610,N_6544);
nor U9040 (N_9040,N_7674,N_6559);
and U9041 (N_9041,N_7768,N_6174);
nand U9042 (N_9042,N_7062,N_6308);
nand U9043 (N_9043,N_6195,N_6582);
and U9044 (N_9044,N_6314,N_7170);
and U9045 (N_9045,N_6371,N_6553);
or U9046 (N_9046,N_7056,N_6027);
and U9047 (N_9047,N_6548,N_6080);
nand U9048 (N_9048,N_6698,N_7369);
or U9049 (N_9049,N_6448,N_6269);
nor U9050 (N_9050,N_7159,N_6405);
and U9051 (N_9051,N_6396,N_7261);
or U9052 (N_9052,N_6827,N_7339);
or U9053 (N_9053,N_6625,N_7444);
nand U9054 (N_9054,N_6884,N_7637);
nand U9055 (N_9055,N_6725,N_6875);
nor U9056 (N_9056,N_6062,N_6136);
nand U9057 (N_9057,N_6406,N_6343);
xor U9058 (N_9058,N_6826,N_6523);
nand U9059 (N_9059,N_6664,N_6776);
xnor U9060 (N_9060,N_7374,N_6535);
and U9061 (N_9061,N_6407,N_7932);
nor U9062 (N_9062,N_6627,N_6809);
nand U9063 (N_9063,N_6178,N_7160);
and U9064 (N_9064,N_6244,N_6146);
nand U9065 (N_9065,N_6967,N_7559);
and U9066 (N_9066,N_6786,N_6916);
nor U9067 (N_9067,N_7338,N_7324);
nor U9068 (N_9068,N_6337,N_7506);
and U9069 (N_9069,N_7562,N_6789);
nor U9070 (N_9070,N_6250,N_6468);
nor U9071 (N_9071,N_6875,N_6343);
nor U9072 (N_9072,N_6823,N_7447);
or U9073 (N_9073,N_7448,N_6742);
nand U9074 (N_9074,N_7033,N_7122);
nor U9075 (N_9075,N_7246,N_7258);
or U9076 (N_9076,N_7005,N_7867);
or U9077 (N_9077,N_7579,N_6046);
nand U9078 (N_9078,N_7420,N_6099);
and U9079 (N_9079,N_7991,N_7964);
or U9080 (N_9080,N_7317,N_7746);
and U9081 (N_9081,N_7052,N_6794);
nor U9082 (N_9082,N_7930,N_6239);
nor U9083 (N_9083,N_7769,N_7727);
and U9084 (N_9084,N_6379,N_7453);
nor U9085 (N_9085,N_7353,N_6381);
and U9086 (N_9086,N_7279,N_7732);
and U9087 (N_9087,N_6726,N_7583);
or U9088 (N_9088,N_7709,N_6781);
nor U9089 (N_9089,N_7732,N_6174);
or U9090 (N_9090,N_6036,N_7920);
nor U9091 (N_9091,N_6489,N_7679);
nand U9092 (N_9092,N_6431,N_6589);
or U9093 (N_9093,N_7522,N_6895);
nor U9094 (N_9094,N_7773,N_7731);
nor U9095 (N_9095,N_6748,N_6308);
nand U9096 (N_9096,N_7188,N_7398);
or U9097 (N_9097,N_6090,N_6297);
xor U9098 (N_9098,N_7074,N_7484);
and U9099 (N_9099,N_6045,N_6774);
nor U9100 (N_9100,N_6046,N_7833);
nand U9101 (N_9101,N_6827,N_6720);
nor U9102 (N_9102,N_6794,N_7841);
and U9103 (N_9103,N_7580,N_6828);
or U9104 (N_9104,N_6416,N_6893);
nor U9105 (N_9105,N_6501,N_7316);
nor U9106 (N_9106,N_7411,N_6204);
or U9107 (N_9107,N_6308,N_6393);
nand U9108 (N_9108,N_6675,N_6301);
and U9109 (N_9109,N_7465,N_7975);
nand U9110 (N_9110,N_6771,N_7377);
and U9111 (N_9111,N_6528,N_6594);
xnor U9112 (N_9112,N_7851,N_7813);
nor U9113 (N_9113,N_6631,N_7232);
nor U9114 (N_9114,N_6869,N_7995);
nor U9115 (N_9115,N_7511,N_6380);
xnor U9116 (N_9116,N_7224,N_7835);
and U9117 (N_9117,N_7894,N_7708);
nand U9118 (N_9118,N_7293,N_6085);
nand U9119 (N_9119,N_7660,N_6601);
xnor U9120 (N_9120,N_6451,N_7906);
or U9121 (N_9121,N_7526,N_7671);
and U9122 (N_9122,N_7158,N_6465);
nor U9123 (N_9123,N_6306,N_7272);
and U9124 (N_9124,N_6551,N_6812);
nand U9125 (N_9125,N_6233,N_6848);
and U9126 (N_9126,N_7516,N_6636);
and U9127 (N_9127,N_7489,N_6819);
and U9128 (N_9128,N_7012,N_6038);
nand U9129 (N_9129,N_6702,N_7585);
and U9130 (N_9130,N_7933,N_6717);
and U9131 (N_9131,N_7365,N_7578);
nor U9132 (N_9132,N_6991,N_7601);
nand U9133 (N_9133,N_6285,N_6188);
and U9134 (N_9134,N_6979,N_7900);
nand U9135 (N_9135,N_6001,N_7572);
or U9136 (N_9136,N_7179,N_6755);
xnor U9137 (N_9137,N_6664,N_6369);
or U9138 (N_9138,N_7766,N_7454);
and U9139 (N_9139,N_7780,N_7400);
or U9140 (N_9140,N_7336,N_6492);
or U9141 (N_9141,N_6873,N_6904);
nor U9142 (N_9142,N_6355,N_6357);
and U9143 (N_9143,N_7725,N_6396);
and U9144 (N_9144,N_6664,N_6515);
or U9145 (N_9145,N_7896,N_7261);
nand U9146 (N_9146,N_6977,N_6517);
nor U9147 (N_9147,N_7075,N_6292);
and U9148 (N_9148,N_6452,N_7133);
or U9149 (N_9149,N_6553,N_6576);
and U9150 (N_9150,N_7940,N_6133);
nor U9151 (N_9151,N_7572,N_6716);
nand U9152 (N_9152,N_7133,N_7105);
or U9153 (N_9153,N_6086,N_7672);
and U9154 (N_9154,N_6442,N_7108);
and U9155 (N_9155,N_7839,N_6210);
nor U9156 (N_9156,N_7654,N_6428);
nor U9157 (N_9157,N_7420,N_6788);
or U9158 (N_9158,N_6854,N_7480);
or U9159 (N_9159,N_6038,N_6450);
xor U9160 (N_9160,N_7136,N_7089);
nor U9161 (N_9161,N_6178,N_6656);
nor U9162 (N_9162,N_6748,N_7206);
or U9163 (N_9163,N_7843,N_6121);
nor U9164 (N_9164,N_7136,N_7316);
or U9165 (N_9165,N_6256,N_6603);
nor U9166 (N_9166,N_7602,N_7139);
nor U9167 (N_9167,N_7225,N_7834);
or U9168 (N_9168,N_6474,N_6214);
and U9169 (N_9169,N_6455,N_7562);
nor U9170 (N_9170,N_6291,N_7297);
or U9171 (N_9171,N_6194,N_6674);
or U9172 (N_9172,N_6837,N_6016);
or U9173 (N_9173,N_7033,N_6081);
and U9174 (N_9174,N_7520,N_7518);
nand U9175 (N_9175,N_7396,N_6128);
xor U9176 (N_9176,N_6305,N_7811);
or U9177 (N_9177,N_6108,N_7615);
xnor U9178 (N_9178,N_6181,N_6089);
or U9179 (N_9179,N_6671,N_7925);
and U9180 (N_9180,N_7436,N_6383);
nor U9181 (N_9181,N_6551,N_7894);
nor U9182 (N_9182,N_6879,N_6722);
or U9183 (N_9183,N_6479,N_6020);
and U9184 (N_9184,N_7825,N_7780);
or U9185 (N_9185,N_7215,N_7016);
or U9186 (N_9186,N_6752,N_7440);
and U9187 (N_9187,N_6104,N_6816);
or U9188 (N_9188,N_6956,N_6530);
nor U9189 (N_9189,N_6593,N_6360);
or U9190 (N_9190,N_7191,N_7516);
and U9191 (N_9191,N_6617,N_7466);
xor U9192 (N_9192,N_7196,N_6989);
or U9193 (N_9193,N_6706,N_6712);
or U9194 (N_9194,N_7805,N_6447);
nand U9195 (N_9195,N_7119,N_7293);
and U9196 (N_9196,N_7237,N_6686);
nand U9197 (N_9197,N_7748,N_7577);
nor U9198 (N_9198,N_6926,N_6145);
and U9199 (N_9199,N_7008,N_6059);
nand U9200 (N_9200,N_7558,N_7951);
or U9201 (N_9201,N_7523,N_7836);
or U9202 (N_9202,N_6104,N_6196);
nor U9203 (N_9203,N_6954,N_7026);
and U9204 (N_9204,N_7987,N_6691);
and U9205 (N_9205,N_6085,N_7833);
or U9206 (N_9206,N_6326,N_6681);
and U9207 (N_9207,N_7127,N_7438);
or U9208 (N_9208,N_6986,N_7421);
nand U9209 (N_9209,N_7876,N_6552);
nor U9210 (N_9210,N_7491,N_6425);
nand U9211 (N_9211,N_6375,N_7332);
nor U9212 (N_9212,N_7173,N_6940);
and U9213 (N_9213,N_6138,N_7417);
and U9214 (N_9214,N_7750,N_6009);
nand U9215 (N_9215,N_7885,N_7543);
nor U9216 (N_9216,N_7337,N_6783);
or U9217 (N_9217,N_7412,N_6475);
nand U9218 (N_9218,N_6182,N_6767);
and U9219 (N_9219,N_7100,N_6411);
nand U9220 (N_9220,N_6061,N_7654);
nor U9221 (N_9221,N_7329,N_6050);
nor U9222 (N_9222,N_6037,N_6691);
nor U9223 (N_9223,N_7691,N_6367);
or U9224 (N_9224,N_7273,N_6596);
or U9225 (N_9225,N_7652,N_7137);
and U9226 (N_9226,N_6662,N_7991);
nor U9227 (N_9227,N_6285,N_7383);
or U9228 (N_9228,N_6471,N_6209);
and U9229 (N_9229,N_6199,N_6106);
nor U9230 (N_9230,N_7734,N_6139);
and U9231 (N_9231,N_6947,N_7784);
nor U9232 (N_9232,N_7919,N_6821);
nand U9233 (N_9233,N_7851,N_6651);
or U9234 (N_9234,N_7114,N_6896);
or U9235 (N_9235,N_7266,N_6140);
nand U9236 (N_9236,N_7345,N_7417);
nor U9237 (N_9237,N_7341,N_7053);
and U9238 (N_9238,N_6384,N_6358);
and U9239 (N_9239,N_6346,N_7067);
or U9240 (N_9240,N_6268,N_7557);
nand U9241 (N_9241,N_7001,N_6879);
nand U9242 (N_9242,N_6009,N_6230);
nand U9243 (N_9243,N_7830,N_7130);
or U9244 (N_9244,N_7370,N_7123);
nand U9245 (N_9245,N_6507,N_6681);
or U9246 (N_9246,N_6991,N_6019);
and U9247 (N_9247,N_7525,N_6211);
nor U9248 (N_9248,N_6121,N_6567);
and U9249 (N_9249,N_7701,N_6290);
or U9250 (N_9250,N_7925,N_7084);
nor U9251 (N_9251,N_6001,N_7296);
or U9252 (N_9252,N_7971,N_7395);
nor U9253 (N_9253,N_6965,N_7121);
nand U9254 (N_9254,N_6841,N_6976);
or U9255 (N_9255,N_7763,N_7630);
or U9256 (N_9256,N_6446,N_6897);
or U9257 (N_9257,N_6960,N_7092);
nor U9258 (N_9258,N_7479,N_7261);
or U9259 (N_9259,N_6020,N_6636);
xnor U9260 (N_9260,N_7911,N_6560);
or U9261 (N_9261,N_6611,N_6955);
and U9262 (N_9262,N_7373,N_7439);
and U9263 (N_9263,N_6690,N_7428);
or U9264 (N_9264,N_6470,N_7525);
nand U9265 (N_9265,N_7873,N_6409);
and U9266 (N_9266,N_7309,N_6523);
and U9267 (N_9267,N_7355,N_7272);
nand U9268 (N_9268,N_6309,N_7860);
nor U9269 (N_9269,N_7546,N_6853);
nand U9270 (N_9270,N_6226,N_6969);
and U9271 (N_9271,N_7422,N_6601);
nor U9272 (N_9272,N_6730,N_7312);
and U9273 (N_9273,N_7285,N_6774);
xnor U9274 (N_9274,N_6829,N_6526);
and U9275 (N_9275,N_7420,N_6050);
xor U9276 (N_9276,N_7307,N_6956);
nand U9277 (N_9277,N_7013,N_7045);
and U9278 (N_9278,N_6311,N_7552);
and U9279 (N_9279,N_6193,N_7609);
or U9280 (N_9280,N_7109,N_6876);
or U9281 (N_9281,N_7103,N_6840);
or U9282 (N_9282,N_7750,N_7569);
nand U9283 (N_9283,N_6103,N_7798);
and U9284 (N_9284,N_7974,N_7887);
nand U9285 (N_9285,N_6242,N_6799);
nand U9286 (N_9286,N_7479,N_7810);
nand U9287 (N_9287,N_7385,N_6794);
and U9288 (N_9288,N_6857,N_6217);
nand U9289 (N_9289,N_7913,N_7920);
or U9290 (N_9290,N_7806,N_7383);
or U9291 (N_9291,N_7702,N_6944);
or U9292 (N_9292,N_6264,N_7551);
or U9293 (N_9293,N_7504,N_6725);
and U9294 (N_9294,N_7391,N_7164);
nor U9295 (N_9295,N_7734,N_7373);
and U9296 (N_9296,N_7922,N_7735);
and U9297 (N_9297,N_6326,N_7270);
and U9298 (N_9298,N_7869,N_7279);
nor U9299 (N_9299,N_7006,N_6382);
nor U9300 (N_9300,N_7604,N_7892);
and U9301 (N_9301,N_6888,N_6392);
and U9302 (N_9302,N_6898,N_7326);
nor U9303 (N_9303,N_6262,N_7223);
and U9304 (N_9304,N_7166,N_6158);
xor U9305 (N_9305,N_6080,N_7958);
and U9306 (N_9306,N_7702,N_7056);
nor U9307 (N_9307,N_6469,N_6055);
nor U9308 (N_9308,N_7534,N_7061);
and U9309 (N_9309,N_7499,N_6735);
or U9310 (N_9310,N_7057,N_7076);
nor U9311 (N_9311,N_6377,N_6742);
and U9312 (N_9312,N_6972,N_6020);
or U9313 (N_9313,N_6102,N_6860);
nand U9314 (N_9314,N_6444,N_7217);
nor U9315 (N_9315,N_7245,N_6717);
nor U9316 (N_9316,N_7822,N_7245);
or U9317 (N_9317,N_6058,N_6702);
nand U9318 (N_9318,N_6142,N_7224);
nand U9319 (N_9319,N_6829,N_6930);
and U9320 (N_9320,N_7486,N_7369);
nor U9321 (N_9321,N_7689,N_6863);
or U9322 (N_9322,N_6784,N_6236);
nand U9323 (N_9323,N_7856,N_7236);
nand U9324 (N_9324,N_6118,N_7734);
or U9325 (N_9325,N_6903,N_7111);
or U9326 (N_9326,N_7784,N_7760);
nand U9327 (N_9327,N_7982,N_6963);
or U9328 (N_9328,N_7809,N_7838);
or U9329 (N_9329,N_7748,N_6737);
and U9330 (N_9330,N_6885,N_6081);
or U9331 (N_9331,N_7469,N_7163);
or U9332 (N_9332,N_7934,N_7200);
nor U9333 (N_9333,N_7610,N_7942);
nor U9334 (N_9334,N_7883,N_6650);
nand U9335 (N_9335,N_6065,N_6600);
and U9336 (N_9336,N_7614,N_7667);
or U9337 (N_9337,N_7710,N_7644);
and U9338 (N_9338,N_6826,N_6060);
nor U9339 (N_9339,N_7290,N_7645);
nand U9340 (N_9340,N_6782,N_6251);
and U9341 (N_9341,N_7060,N_6550);
nand U9342 (N_9342,N_6613,N_6171);
nand U9343 (N_9343,N_6681,N_7963);
nor U9344 (N_9344,N_6772,N_6987);
nor U9345 (N_9345,N_7237,N_7984);
and U9346 (N_9346,N_7446,N_6490);
or U9347 (N_9347,N_7605,N_7506);
nand U9348 (N_9348,N_7081,N_6572);
nor U9349 (N_9349,N_7038,N_7930);
nand U9350 (N_9350,N_7098,N_6015);
xnor U9351 (N_9351,N_6493,N_7667);
or U9352 (N_9352,N_6309,N_6962);
or U9353 (N_9353,N_7217,N_6091);
and U9354 (N_9354,N_6609,N_6855);
nand U9355 (N_9355,N_7775,N_6003);
nor U9356 (N_9356,N_6802,N_7491);
nor U9357 (N_9357,N_7753,N_7479);
or U9358 (N_9358,N_6524,N_6492);
and U9359 (N_9359,N_7429,N_6843);
or U9360 (N_9360,N_6727,N_7047);
nand U9361 (N_9361,N_7638,N_7120);
or U9362 (N_9362,N_7730,N_7728);
and U9363 (N_9363,N_7772,N_6952);
xor U9364 (N_9364,N_6301,N_7331);
nor U9365 (N_9365,N_7927,N_6008);
nor U9366 (N_9366,N_6670,N_7026);
nand U9367 (N_9367,N_6137,N_7447);
xnor U9368 (N_9368,N_7032,N_7875);
and U9369 (N_9369,N_6694,N_7011);
nor U9370 (N_9370,N_7577,N_7608);
nor U9371 (N_9371,N_6712,N_7731);
nand U9372 (N_9372,N_7635,N_7493);
or U9373 (N_9373,N_7593,N_7522);
nand U9374 (N_9374,N_7071,N_7548);
or U9375 (N_9375,N_6542,N_7208);
nand U9376 (N_9376,N_6408,N_7680);
and U9377 (N_9377,N_6734,N_7511);
nand U9378 (N_9378,N_7183,N_6772);
nor U9379 (N_9379,N_6885,N_6862);
nor U9380 (N_9380,N_6149,N_6607);
or U9381 (N_9381,N_6947,N_6906);
nand U9382 (N_9382,N_7254,N_7779);
nand U9383 (N_9383,N_6767,N_6642);
and U9384 (N_9384,N_7281,N_6744);
nand U9385 (N_9385,N_6076,N_7133);
and U9386 (N_9386,N_7518,N_7001);
and U9387 (N_9387,N_7052,N_7742);
nor U9388 (N_9388,N_6667,N_6697);
nor U9389 (N_9389,N_6095,N_6598);
nor U9390 (N_9390,N_7656,N_7151);
and U9391 (N_9391,N_6268,N_7033);
and U9392 (N_9392,N_6120,N_6306);
nand U9393 (N_9393,N_6960,N_7534);
or U9394 (N_9394,N_6729,N_6032);
or U9395 (N_9395,N_6474,N_6427);
and U9396 (N_9396,N_7462,N_6819);
nor U9397 (N_9397,N_6786,N_6731);
nand U9398 (N_9398,N_6677,N_6455);
or U9399 (N_9399,N_7614,N_6378);
nand U9400 (N_9400,N_7187,N_7170);
nand U9401 (N_9401,N_6821,N_6005);
or U9402 (N_9402,N_7882,N_7108);
or U9403 (N_9403,N_7076,N_7022);
and U9404 (N_9404,N_6278,N_7988);
or U9405 (N_9405,N_7187,N_7110);
xnor U9406 (N_9406,N_7046,N_6708);
nand U9407 (N_9407,N_7378,N_6178);
and U9408 (N_9408,N_6430,N_6702);
nand U9409 (N_9409,N_6740,N_7255);
nand U9410 (N_9410,N_7704,N_7259);
nor U9411 (N_9411,N_7047,N_7755);
nand U9412 (N_9412,N_7428,N_7412);
or U9413 (N_9413,N_7737,N_7272);
nand U9414 (N_9414,N_7685,N_7261);
nand U9415 (N_9415,N_7813,N_6814);
nand U9416 (N_9416,N_6583,N_7182);
and U9417 (N_9417,N_6300,N_6321);
and U9418 (N_9418,N_6129,N_7293);
nor U9419 (N_9419,N_6423,N_6182);
and U9420 (N_9420,N_7322,N_7696);
and U9421 (N_9421,N_6555,N_6166);
nand U9422 (N_9422,N_6135,N_7875);
or U9423 (N_9423,N_7774,N_6675);
or U9424 (N_9424,N_7100,N_6006);
and U9425 (N_9425,N_6088,N_7159);
or U9426 (N_9426,N_7536,N_7488);
nor U9427 (N_9427,N_7572,N_7503);
or U9428 (N_9428,N_6224,N_7654);
and U9429 (N_9429,N_7477,N_6377);
nor U9430 (N_9430,N_7455,N_7966);
nor U9431 (N_9431,N_6481,N_7178);
or U9432 (N_9432,N_6169,N_7677);
nand U9433 (N_9433,N_7280,N_6899);
and U9434 (N_9434,N_7116,N_7786);
nor U9435 (N_9435,N_7073,N_7337);
nand U9436 (N_9436,N_6259,N_6091);
nand U9437 (N_9437,N_6511,N_6352);
nand U9438 (N_9438,N_6232,N_7487);
nand U9439 (N_9439,N_6037,N_6449);
and U9440 (N_9440,N_6222,N_7472);
nand U9441 (N_9441,N_7615,N_6627);
nor U9442 (N_9442,N_7707,N_7942);
nor U9443 (N_9443,N_6613,N_7433);
or U9444 (N_9444,N_6846,N_6447);
and U9445 (N_9445,N_6051,N_6268);
nor U9446 (N_9446,N_6837,N_7608);
nor U9447 (N_9447,N_7727,N_6178);
and U9448 (N_9448,N_7733,N_6057);
nand U9449 (N_9449,N_7923,N_7043);
and U9450 (N_9450,N_7141,N_7155);
xnor U9451 (N_9451,N_7626,N_6410);
or U9452 (N_9452,N_7623,N_6745);
and U9453 (N_9453,N_6112,N_7046);
and U9454 (N_9454,N_6700,N_6070);
nor U9455 (N_9455,N_7373,N_6292);
nor U9456 (N_9456,N_7742,N_7571);
nand U9457 (N_9457,N_6614,N_6232);
nand U9458 (N_9458,N_7026,N_7942);
nand U9459 (N_9459,N_7329,N_7174);
nand U9460 (N_9460,N_6360,N_6613);
nand U9461 (N_9461,N_6959,N_6153);
nor U9462 (N_9462,N_7875,N_7468);
nor U9463 (N_9463,N_7345,N_6273);
nor U9464 (N_9464,N_6474,N_7246);
and U9465 (N_9465,N_6823,N_6969);
and U9466 (N_9466,N_6908,N_6805);
nand U9467 (N_9467,N_7490,N_6062);
nor U9468 (N_9468,N_7108,N_7154);
nor U9469 (N_9469,N_6625,N_7241);
and U9470 (N_9470,N_7351,N_6805);
or U9471 (N_9471,N_6675,N_6866);
nor U9472 (N_9472,N_6875,N_6947);
and U9473 (N_9473,N_6196,N_6907);
and U9474 (N_9474,N_7954,N_6118);
and U9475 (N_9475,N_7017,N_6626);
nand U9476 (N_9476,N_7638,N_7579);
nand U9477 (N_9477,N_7429,N_7311);
and U9478 (N_9478,N_6974,N_6708);
nor U9479 (N_9479,N_7453,N_6050);
nand U9480 (N_9480,N_6274,N_6262);
nor U9481 (N_9481,N_7484,N_6977);
or U9482 (N_9482,N_7031,N_6535);
nor U9483 (N_9483,N_7527,N_7478);
nor U9484 (N_9484,N_6811,N_6869);
and U9485 (N_9485,N_6931,N_7369);
or U9486 (N_9486,N_6303,N_6144);
nor U9487 (N_9487,N_7967,N_6928);
or U9488 (N_9488,N_6947,N_6418);
nor U9489 (N_9489,N_7156,N_7171);
and U9490 (N_9490,N_7150,N_6295);
or U9491 (N_9491,N_6536,N_7286);
or U9492 (N_9492,N_6262,N_6846);
nor U9493 (N_9493,N_6868,N_6756);
and U9494 (N_9494,N_6675,N_7909);
nor U9495 (N_9495,N_7288,N_7955);
nand U9496 (N_9496,N_7523,N_7619);
nand U9497 (N_9497,N_6322,N_6214);
nor U9498 (N_9498,N_6458,N_7379);
nor U9499 (N_9499,N_7270,N_7592);
and U9500 (N_9500,N_6019,N_7382);
and U9501 (N_9501,N_6851,N_6453);
nor U9502 (N_9502,N_6918,N_7564);
or U9503 (N_9503,N_7374,N_6293);
and U9504 (N_9504,N_6499,N_7256);
and U9505 (N_9505,N_7321,N_6084);
and U9506 (N_9506,N_7608,N_6445);
or U9507 (N_9507,N_6173,N_6573);
nand U9508 (N_9508,N_6699,N_7879);
and U9509 (N_9509,N_6541,N_6936);
xnor U9510 (N_9510,N_6721,N_7504);
and U9511 (N_9511,N_7612,N_6709);
nand U9512 (N_9512,N_7881,N_7946);
and U9513 (N_9513,N_6777,N_6975);
nor U9514 (N_9514,N_6199,N_7290);
nand U9515 (N_9515,N_6943,N_7555);
and U9516 (N_9516,N_6282,N_6127);
or U9517 (N_9517,N_7278,N_7591);
nor U9518 (N_9518,N_6984,N_6920);
or U9519 (N_9519,N_7363,N_7868);
and U9520 (N_9520,N_6501,N_7075);
nor U9521 (N_9521,N_6379,N_6255);
and U9522 (N_9522,N_7579,N_6837);
or U9523 (N_9523,N_6178,N_6571);
or U9524 (N_9524,N_7837,N_7179);
nand U9525 (N_9525,N_7760,N_7681);
or U9526 (N_9526,N_7651,N_7574);
or U9527 (N_9527,N_6305,N_7739);
nor U9528 (N_9528,N_6905,N_6508);
or U9529 (N_9529,N_6816,N_6589);
nand U9530 (N_9530,N_6506,N_6414);
nor U9531 (N_9531,N_6537,N_6291);
and U9532 (N_9532,N_7855,N_6637);
and U9533 (N_9533,N_7024,N_7901);
and U9534 (N_9534,N_6986,N_6351);
xnor U9535 (N_9535,N_6586,N_7727);
and U9536 (N_9536,N_6459,N_6861);
or U9537 (N_9537,N_6135,N_6207);
or U9538 (N_9538,N_7093,N_7506);
nand U9539 (N_9539,N_6565,N_7925);
or U9540 (N_9540,N_7268,N_6415);
and U9541 (N_9541,N_7006,N_7688);
nor U9542 (N_9542,N_7934,N_6142);
nand U9543 (N_9543,N_6225,N_6733);
nor U9544 (N_9544,N_6551,N_7816);
nand U9545 (N_9545,N_7782,N_7904);
or U9546 (N_9546,N_7124,N_7044);
nand U9547 (N_9547,N_6010,N_7496);
nand U9548 (N_9548,N_6080,N_7687);
or U9549 (N_9549,N_6750,N_7436);
and U9550 (N_9550,N_7695,N_7398);
nand U9551 (N_9551,N_6080,N_7930);
nand U9552 (N_9552,N_6828,N_7108);
nor U9553 (N_9553,N_7183,N_6194);
or U9554 (N_9554,N_7952,N_7130);
and U9555 (N_9555,N_6250,N_7321);
or U9556 (N_9556,N_7079,N_6033);
nand U9557 (N_9557,N_6175,N_6464);
nor U9558 (N_9558,N_6653,N_7214);
or U9559 (N_9559,N_6628,N_7375);
or U9560 (N_9560,N_7052,N_7619);
nor U9561 (N_9561,N_7110,N_7742);
nor U9562 (N_9562,N_6208,N_7349);
and U9563 (N_9563,N_7520,N_6153);
or U9564 (N_9564,N_7810,N_7389);
or U9565 (N_9565,N_6348,N_7786);
nand U9566 (N_9566,N_7193,N_6738);
xnor U9567 (N_9567,N_6142,N_7774);
or U9568 (N_9568,N_6946,N_7352);
nor U9569 (N_9569,N_7843,N_6041);
and U9570 (N_9570,N_7882,N_7883);
and U9571 (N_9571,N_6449,N_6658);
and U9572 (N_9572,N_7778,N_7973);
and U9573 (N_9573,N_6687,N_7558);
or U9574 (N_9574,N_6046,N_7773);
or U9575 (N_9575,N_7030,N_7782);
or U9576 (N_9576,N_7186,N_7158);
nand U9577 (N_9577,N_6220,N_6731);
or U9578 (N_9578,N_7900,N_7642);
or U9579 (N_9579,N_6265,N_6897);
xor U9580 (N_9580,N_6048,N_7382);
xnor U9581 (N_9581,N_6121,N_6761);
xnor U9582 (N_9582,N_7729,N_6643);
or U9583 (N_9583,N_6656,N_6519);
and U9584 (N_9584,N_7631,N_6101);
nand U9585 (N_9585,N_7263,N_6626);
nand U9586 (N_9586,N_7065,N_7133);
nor U9587 (N_9587,N_7164,N_7555);
and U9588 (N_9588,N_7671,N_6847);
nand U9589 (N_9589,N_7186,N_6898);
or U9590 (N_9590,N_7656,N_7185);
nor U9591 (N_9591,N_6096,N_7596);
nor U9592 (N_9592,N_6329,N_6604);
and U9593 (N_9593,N_6182,N_7419);
and U9594 (N_9594,N_6889,N_6203);
and U9595 (N_9595,N_6240,N_7446);
nor U9596 (N_9596,N_7888,N_7285);
and U9597 (N_9597,N_7348,N_7736);
nor U9598 (N_9598,N_6940,N_6484);
and U9599 (N_9599,N_6587,N_7034);
or U9600 (N_9600,N_7653,N_6239);
or U9601 (N_9601,N_7843,N_6045);
nor U9602 (N_9602,N_6406,N_6516);
and U9603 (N_9603,N_6381,N_6269);
and U9604 (N_9604,N_6386,N_6798);
or U9605 (N_9605,N_7421,N_6780);
and U9606 (N_9606,N_7477,N_7027);
nand U9607 (N_9607,N_6895,N_6225);
nand U9608 (N_9608,N_6365,N_6121);
or U9609 (N_9609,N_7719,N_6523);
and U9610 (N_9610,N_7866,N_7047);
nor U9611 (N_9611,N_6368,N_6892);
nand U9612 (N_9612,N_7227,N_6121);
nor U9613 (N_9613,N_7115,N_6300);
and U9614 (N_9614,N_6788,N_6883);
or U9615 (N_9615,N_7873,N_6270);
nor U9616 (N_9616,N_6696,N_7398);
nor U9617 (N_9617,N_6664,N_6519);
nand U9618 (N_9618,N_6083,N_7168);
nand U9619 (N_9619,N_6386,N_7019);
nor U9620 (N_9620,N_7160,N_7752);
nor U9621 (N_9621,N_7748,N_7805);
or U9622 (N_9622,N_7681,N_7185);
nand U9623 (N_9623,N_6162,N_7788);
nand U9624 (N_9624,N_6454,N_7995);
or U9625 (N_9625,N_6876,N_6435);
nor U9626 (N_9626,N_7265,N_6278);
nor U9627 (N_9627,N_6291,N_6189);
nand U9628 (N_9628,N_7984,N_6849);
nor U9629 (N_9629,N_6863,N_6653);
or U9630 (N_9630,N_7408,N_7474);
or U9631 (N_9631,N_6470,N_7152);
nor U9632 (N_9632,N_6869,N_7110);
nand U9633 (N_9633,N_7290,N_6616);
and U9634 (N_9634,N_7670,N_6119);
and U9635 (N_9635,N_6998,N_7840);
and U9636 (N_9636,N_6358,N_7109);
nand U9637 (N_9637,N_6062,N_7560);
or U9638 (N_9638,N_7193,N_6129);
or U9639 (N_9639,N_7506,N_7524);
and U9640 (N_9640,N_7293,N_7537);
and U9641 (N_9641,N_7886,N_7255);
and U9642 (N_9642,N_7937,N_7988);
and U9643 (N_9643,N_7050,N_6152);
or U9644 (N_9644,N_7155,N_6829);
nor U9645 (N_9645,N_7882,N_7776);
or U9646 (N_9646,N_6528,N_6431);
nor U9647 (N_9647,N_6529,N_6383);
nor U9648 (N_9648,N_7632,N_7070);
or U9649 (N_9649,N_7820,N_6113);
or U9650 (N_9650,N_6554,N_6566);
nand U9651 (N_9651,N_7334,N_6024);
or U9652 (N_9652,N_6152,N_7411);
or U9653 (N_9653,N_6883,N_6647);
nand U9654 (N_9654,N_6767,N_6936);
nor U9655 (N_9655,N_6964,N_7163);
or U9656 (N_9656,N_6411,N_6296);
nor U9657 (N_9657,N_6172,N_6665);
and U9658 (N_9658,N_6944,N_6841);
nand U9659 (N_9659,N_6904,N_7537);
nand U9660 (N_9660,N_6470,N_6380);
and U9661 (N_9661,N_6174,N_6859);
nand U9662 (N_9662,N_6015,N_7232);
or U9663 (N_9663,N_6417,N_6145);
or U9664 (N_9664,N_6502,N_7212);
nor U9665 (N_9665,N_7108,N_7092);
nor U9666 (N_9666,N_7494,N_7366);
and U9667 (N_9667,N_6704,N_6005);
and U9668 (N_9668,N_6990,N_6572);
and U9669 (N_9669,N_6451,N_6235);
nor U9670 (N_9670,N_7449,N_7921);
nor U9671 (N_9671,N_7133,N_7523);
and U9672 (N_9672,N_7729,N_7861);
nand U9673 (N_9673,N_7824,N_7396);
or U9674 (N_9674,N_7583,N_6794);
or U9675 (N_9675,N_6330,N_6195);
nor U9676 (N_9676,N_7045,N_6122);
nand U9677 (N_9677,N_6989,N_7139);
and U9678 (N_9678,N_6084,N_6651);
nor U9679 (N_9679,N_7114,N_6500);
nand U9680 (N_9680,N_6838,N_7894);
nor U9681 (N_9681,N_6237,N_7289);
and U9682 (N_9682,N_7668,N_7786);
or U9683 (N_9683,N_6007,N_7809);
nor U9684 (N_9684,N_7420,N_6878);
nand U9685 (N_9685,N_6195,N_7756);
or U9686 (N_9686,N_7923,N_6234);
nand U9687 (N_9687,N_7454,N_6006);
nor U9688 (N_9688,N_6254,N_6574);
nand U9689 (N_9689,N_7407,N_7999);
or U9690 (N_9690,N_7649,N_6726);
nor U9691 (N_9691,N_6998,N_6891);
xor U9692 (N_9692,N_6592,N_7392);
and U9693 (N_9693,N_6869,N_6845);
nor U9694 (N_9694,N_6233,N_7366);
or U9695 (N_9695,N_7377,N_7362);
nor U9696 (N_9696,N_6895,N_7484);
nor U9697 (N_9697,N_7398,N_6780);
nand U9698 (N_9698,N_6913,N_6472);
nand U9699 (N_9699,N_6641,N_7877);
nor U9700 (N_9700,N_6971,N_7628);
nor U9701 (N_9701,N_6736,N_7974);
and U9702 (N_9702,N_7937,N_6022);
and U9703 (N_9703,N_7514,N_6880);
or U9704 (N_9704,N_7860,N_6615);
xnor U9705 (N_9705,N_6516,N_6560);
nand U9706 (N_9706,N_6334,N_6056);
and U9707 (N_9707,N_6794,N_6199);
or U9708 (N_9708,N_6722,N_7589);
nor U9709 (N_9709,N_7832,N_7342);
and U9710 (N_9710,N_6833,N_6302);
nand U9711 (N_9711,N_7609,N_6445);
or U9712 (N_9712,N_7064,N_7730);
or U9713 (N_9713,N_6660,N_7004);
and U9714 (N_9714,N_7077,N_6838);
nor U9715 (N_9715,N_7419,N_6322);
nor U9716 (N_9716,N_7298,N_6343);
and U9717 (N_9717,N_6172,N_6965);
or U9718 (N_9718,N_6265,N_6955);
nand U9719 (N_9719,N_7490,N_7379);
or U9720 (N_9720,N_6348,N_7787);
nor U9721 (N_9721,N_6318,N_7128);
nand U9722 (N_9722,N_7805,N_6283);
nor U9723 (N_9723,N_7392,N_6517);
and U9724 (N_9724,N_6050,N_6002);
nor U9725 (N_9725,N_7018,N_6397);
nand U9726 (N_9726,N_7476,N_6602);
nand U9727 (N_9727,N_7901,N_6319);
nor U9728 (N_9728,N_7804,N_7024);
nand U9729 (N_9729,N_6946,N_6312);
or U9730 (N_9730,N_7277,N_6171);
and U9731 (N_9731,N_7195,N_7381);
nand U9732 (N_9732,N_7598,N_6155);
nand U9733 (N_9733,N_7417,N_6310);
and U9734 (N_9734,N_7458,N_6424);
and U9735 (N_9735,N_6736,N_6914);
nor U9736 (N_9736,N_6307,N_6414);
and U9737 (N_9737,N_7104,N_7818);
nand U9738 (N_9738,N_6169,N_6016);
nand U9739 (N_9739,N_7851,N_7159);
and U9740 (N_9740,N_7768,N_7702);
and U9741 (N_9741,N_7117,N_6073);
and U9742 (N_9742,N_7152,N_7471);
nor U9743 (N_9743,N_6735,N_6786);
nor U9744 (N_9744,N_6032,N_6691);
nand U9745 (N_9745,N_6539,N_7047);
nand U9746 (N_9746,N_6672,N_7181);
or U9747 (N_9747,N_6085,N_6003);
or U9748 (N_9748,N_7367,N_7777);
and U9749 (N_9749,N_7847,N_6237);
and U9750 (N_9750,N_6140,N_7190);
nand U9751 (N_9751,N_7891,N_7849);
or U9752 (N_9752,N_7098,N_7091);
nand U9753 (N_9753,N_6545,N_6373);
or U9754 (N_9754,N_7187,N_7515);
and U9755 (N_9755,N_7540,N_6298);
or U9756 (N_9756,N_7301,N_7426);
nor U9757 (N_9757,N_6014,N_6759);
and U9758 (N_9758,N_6670,N_7817);
and U9759 (N_9759,N_7376,N_7302);
and U9760 (N_9760,N_6093,N_7730);
nand U9761 (N_9761,N_7595,N_6950);
nor U9762 (N_9762,N_6465,N_6364);
or U9763 (N_9763,N_7676,N_7897);
and U9764 (N_9764,N_7360,N_7714);
nor U9765 (N_9765,N_6144,N_7876);
nor U9766 (N_9766,N_7886,N_7573);
and U9767 (N_9767,N_7645,N_6895);
or U9768 (N_9768,N_6497,N_7971);
and U9769 (N_9769,N_7122,N_7330);
or U9770 (N_9770,N_6732,N_6121);
or U9771 (N_9771,N_6551,N_7377);
or U9772 (N_9772,N_7259,N_6028);
or U9773 (N_9773,N_6432,N_7721);
nand U9774 (N_9774,N_7819,N_6857);
nor U9775 (N_9775,N_7181,N_6419);
nor U9776 (N_9776,N_6099,N_6103);
and U9777 (N_9777,N_6265,N_6184);
nor U9778 (N_9778,N_6533,N_6667);
and U9779 (N_9779,N_6298,N_7570);
nor U9780 (N_9780,N_6005,N_6494);
nor U9781 (N_9781,N_7598,N_7319);
or U9782 (N_9782,N_7916,N_6713);
nand U9783 (N_9783,N_6791,N_7028);
nand U9784 (N_9784,N_7896,N_7101);
or U9785 (N_9785,N_6325,N_6573);
nor U9786 (N_9786,N_7388,N_6827);
or U9787 (N_9787,N_7219,N_6387);
nand U9788 (N_9788,N_6840,N_6425);
and U9789 (N_9789,N_6539,N_6894);
and U9790 (N_9790,N_7326,N_7761);
nor U9791 (N_9791,N_6285,N_6937);
nor U9792 (N_9792,N_6630,N_7109);
and U9793 (N_9793,N_6205,N_7024);
and U9794 (N_9794,N_6381,N_7430);
nand U9795 (N_9795,N_6841,N_6597);
nor U9796 (N_9796,N_7686,N_7843);
or U9797 (N_9797,N_7889,N_7333);
or U9798 (N_9798,N_6301,N_6277);
xor U9799 (N_9799,N_7839,N_6591);
nand U9800 (N_9800,N_6358,N_7989);
nor U9801 (N_9801,N_6463,N_7973);
nand U9802 (N_9802,N_6813,N_6234);
and U9803 (N_9803,N_7440,N_7471);
nor U9804 (N_9804,N_7387,N_6961);
and U9805 (N_9805,N_6324,N_7525);
or U9806 (N_9806,N_6925,N_6075);
and U9807 (N_9807,N_7938,N_7597);
xnor U9808 (N_9808,N_6442,N_6676);
nor U9809 (N_9809,N_7944,N_7759);
nand U9810 (N_9810,N_6212,N_6401);
nand U9811 (N_9811,N_7573,N_7906);
and U9812 (N_9812,N_6486,N_7910);
and U9813 (N_9813,N_7069,N_6211);
or U9814 (N_9814,N_6063,N_7955);
and U9815 (N_9815,N_7095,N_7211);
or U9816 (N_9816,N_6034,N_6591);
nor U9817 (N_9817,N_7855,N_7257);
nor U9818 (N_9818,N_6957,N_6364);
and U9819 (N_9819,N_6925,N_6069);
nor U9820 (N_9820,N_7468,N_6220);
or U9821 (N_9821,N_6787,N_7771);
and U9822 (N_9822,N_6926,N_6987);
or U9823 (N_9823,N_7509,N_6435);
nor U9824 (N_9824,N_7931,N_7735);
or U9825 (N_9825,N_7638,N_6391);
or U9826 (N_9826,N_6073,N_6465);
nor U9827 (N_9827,N_7228,N_7413);
and U9828 (N_9828,N_7015,N_6560);
nor U9829 (N_9829,N_7443,N_7866);
nand U9830 (N_9830,N_7047,N_6154);
and U9831 (N_9831,N_7063,N_6108);
nor U9832 (N_9832,N_7609,N_6930);
and U9833 (N_9833,N_6013,N_7127);
or U9834 (N_9834,N_7160,N_6713);
or U9835 (N_9835,N_6036,N_7894);
nand U9836 (N_9836,N_7235,N_6092);
nor U9837 (N_9837,N_6849,N_7907);
and U9838 (N_9838,N_7159,N_6422);
or U9839 (N_9839,N_6710,N_6115);
nand U9840 (N_9840,N_6066,N_7391);
or U9841 (N_9841,N_7301,N_6487);
and U9842 (N_9842,N_6904,N_6901);
xnor U9843 (N_9843,N_7362,N_6741);
or U9844 (N_9844,N_6546,N_7838);
nor U9845 (N_9845,N_6135,N_7163);
nand U9846 (N_9846,N_7755,N_6111);
nand U9847 (N_9847,N_7648,N_6263);
nor U9848 (N_9848,N_6268,N_7597);
or U9849 (N_9849,N_7130,N_6294);
nand U9850 (N_9850,N_7471,N_6183);
nand U9851 (N_9851,N_7491,N_7806);
and U9852 (N_9852,N_6054,N_7765);
nor U9853 (N_9853,N_7315,N_7562);
or U9854 (N_9854,N_7159,N_6028);
and U9855 (N_9855,N_7016,N_6182);
and U9856 (N_9856,N_7710,N_7190);
or U9857 (N_9857,N_7464,N_7204);
and U9858 (N_9858,N_6379,N_7832);
nor U9859 (N_9859,N_6490,N_6915);
and U9860 (N_9860,N_6675,N_6287);
nand U9861 (N_9861,N_7974,N_6505);
nor U9862 (N_9862,N_6695,N_7301);
or U9863 (N_9863,N_6268,N_6269);
nor U9864 (N_9864,N_6870,N_6256);
xnor U9865 (N_9865,N_6187,N_6261);
or U9866 (N_9866,N_6183,N_6038);
nor U9867 (N_9867,N_6173,N_6667);
nand U9868 (N_9868,N_6975,N_7302);
or U9869 (N_9869,N_6953,N_6206);
nor U9870 (N_9870,N_7674,N_7150);
nand U9871 (N_9871,N_6785,N_7815);
nor U9872 (N_9872,N_7195,N_7475);
nor U9873 (N_9873,N_7217,N_6206);
and U9874 (N_9874,N_7515,N_7016);
nand U9875 (N_9875,N_6458,N_7884);
or U9876 (N_9876,N_7150,N_6064);
and U9877 (N_9877,N_7794,N_6785);
and U9878 (N_9878,N_7071,N_6882);
or U9879 (N_9879,N_6856,N_7661);
and U9880 (N_9880,N_6964,N_7974);
and U9881 (N_9881,N_7955,N_7853);
and U9882 (N_9882,N_7792,N_6751);
nor U9883 (N_9883,N_6427,N_7232);
nand U9884 (N_9884,N_6405,N_6141);
or U9885 (N_9885,N_7540,N_7810);
or U9886 (N_9886,N_7902,N_7600);
and U9887 (N_9887,N_6206,N_7276);
or U9888 (N_9888,N_7196,N_7437);
and U9889 (N_9889,N_6701,N_7539);
or U9890 (N_9890,N_6908,N_6902);
nor U9891 (N_9891,N_6336,N_7233);
and U9892 (N_9892,N_7188,N_6381);
nand U9893 (N_9893,N_6922,N_6998);
nand U9894 (N_9894,N_7778,N_7307);
and U9895 (N_9895,N_7479,N_7103);
or U9896 (N_9896,N_6819,N_6445);
nor U9897 (N_9897,N_6397,N_6827);
or U9898 (N_9898,N_7023,N_7091);
nand U9899 (N_9899,N_7429,N_6341);
nand U9900 (N_9900,N_6725,N_7198);
or U9901 (N_9901,N_6905,N_6197);
or U9902 (N_9902,N_6009,N_7202);
nand U9903 (N_9903,N_6448,N_7446);
and U9904 (N_9904,N_6653,N_6630);
and U9905 (N_9905,N_6721,N_7581);
nor U9906 (N_9906,N_6172,N_6277);
nand U9907 (N_9907,N_7508,N_6683);
and U9908 (N_9908,N_6536,N_6189);
nand U9909 (N_9909,N_6985,N_6461);
and U9910 (N_9910,N_6930,N_7921);
nand U9911 (N_9911,N_7227,N_7284);
and U9912 (N_9912,N_7214,N_6468);
and U9913 (N_9913,N_6228,N_7869);
and U9914 (N_9914,N_7542,N_6248);
and U9915 (N_9915,N_6484,N_6070);
or U9916 (N_9916,N_7748,N_6708);
or U9917 (N_9917,N_7933,N_7043);
and U9918 (N_9918,N_6075,N_6935);
nand U9919 (N_9919,N_7511,N_7921);
or U9920 (N_9920,N_6758,N_7126);
and U9921 (N_9921,N_7193,N_7699);
and U9922 (N_9922,N_7254,N_6306);
nor U9923 (N_9923,N_7907,N_6552);
nand U9924 (N_9924,N_6877,N_6085);
or U9925 (N_9925,N_6764,N_7740);
or U9926 (N_9926,N_6735,N_6051);
or U9927 (N_9927,N_6928,N_6628);
and U9928 (N_9928,N_6429,N_6304);
nor U9929 (N_9929,N_7916,N_6137);
nand U9930 (N_9930,N_7745,N_6341);
or U9931 (N_9931,N_7077,N_6346);
nand U9932 (N_9932,N_7658,N_6620);
or U9933 (N_9933,N_7335,N_7752);
nor U9934 (N_9934,N_6901,N_6004);
nor U9935 (N_9935,N_6381,N_6621);
xor U9936 (N_9936,N_6629,N_6942);
or U9937 (N_9937,N_7631,N_6106);
nand U9938 (N_9938,N_6936,N_7022);
or U9939 (N_9939,N_6098,N_7560);
nor U9940 (N_9940,N_7275,N_6912);
nor U9941 (N_9941,N_7153,N_7270);
and U9942 (N_9942,N_6244,N_6911);
nand U9943 (N_9943,N_7494,N_6622);
or U9944 (N_9944,N_6444,N_7486);
nand U9945 (N_9945,N_7148,N_6878);
nand U9946 (N_9946,N_6007,N_7795);
or U9947 (N_9947,N_6327,N_7542);
nor U9948 (N_9948,N_6587,N_6663);
and U9949 (N_9949,N_7940,N_6606);
xor U9950 (N_9950,N_7201,N_6448);
and U9951 (N_9951,N_7222,N_6921);
nor U9952 (N_9952,N_6572,N_7102);
nor U9953 (N_9953,N_7525,N_6617);
and U9954 (N_9954,N_6663,N_6751);
nor U9955 (N_9955,N_6376,N_6665);
and U9956 (N_9956,N_6516,N_7003);
or U9957 (N_9957,N_6421,N_6972);
or U9958 (N_9958,N_6470,N_6323);
nor U9959 (N_9959,N_6649,N_7333);
or U9960 (N_9960,N_7489,N_7147);
nor U9961 (N_9961,N_6876,N_7396);
nand U9962 (N_9962,N_7821,N_6238);
or U9963 (N_9963,N_7406,N_6796);
and U9964 (N_9964,N_7693,N_7148);
nand U9965 (N_9965,N_7319,N_7087);
nand U9966 (N_9966,N_7563,N_7056);
nand U9967 (N_9967,N_7138,N_6110);
or U9968 (N_9968,N_7877,N_7294);
or U9969 (N_9969,N_7940,N_7384);
or U9970 (N_9970,N_6146,N_7896);
and U9971 (N_9971,N_6275,N_7000);
nand U9972 (N_9972,N_6490,N_7961);
nor U9973 (N_9973,N_6273,N_6256);
and U9974 (N_9974,N_6897,N_7242);
xnor U9975 (N_9975,N_6803,N_6018);
or U9976 (N_9976,N_6216,N_6437);
and U9977 (N_9977,N_6998,N_6981);
or U9978 (N_9978,N_7630,N_7070);
and U9979 (N_9979,N_7101,N_6139);
nor U9980 (N_9980,N_7443,N_6727);
nand U9981 (N_9981,N_6235,N_6251);
or U9982 (N_9982,N_7584,N_7727);
or U9983 (N_9983,N_6262,N_6813);
and U9984 (N_9984,N_7780,N_7817);
or U9985 (N_9985,N_6493,N_7485);
and U9986 (N_9986,N_7647,N_7090);
nor U9987 (N_9987,N_7615,N_6964);
or U9988 (N_9988,N_6172,N_7216);
and U9989 (N_9989,N_7866,N_7533);
or U9990 (N_9990,N_6764,N_6605);
or U9991 (N_9991,N_6262,N_6958);
nor U9992 (N_9992,N_7175,N_7850);
or U9993 (N_9993,N_6824,N_7724);
xnor U9994 (N_9994,N_7192,N_6007);
or U9995 (N_9995,N_7740,N_7804);
or U9996 (N_9996,N_7564,N_6656);
and U9997 (N_9997,N_7089,N_7176);
and U9998 (N_9998,N_7494,N_7572);
or U9999 (N_9999,N_7599,N_6564);
nand UO_0 (O_0,N_8008,N_9565);
or UO_1 (O_1,N_8820,N_9779);
nand UO_2 (O_2,N_9879,N_9855);
nand UO_3 (O_3,N_9890,N_9290);
nand UO_4 (O_4,N_8207,N_8759);
and UO_5 (O_5,N_9989,N_8063);
and UO_6 (O_6,N_9852,N_9518);
or UO_7 (O_7,N_8683,N_8905);
and UO_8 (O_8,N_8706,N_8134);
nor UO_9 (O_9,N_9959,N_9607);
nand UO_10 (O_10,N_8684,N_9987);
and UO_11 (O_11,N_9939,N_8606);
nand UO_12 (O_12,N_8686,N_8525);
or UO_13 (O_13,N_9301,N_8888);
and UO_14 (O_14,N_9831,N_9485);
or UO_15 (O_15,N_9189,N_8476);
and UO_16 (O_16,N_8738,N_8286);
and UO_17 (O_17,N_8656,N_9960);
and UO_18 (O_18,N_8107,N_9193);
and UO_19 (O_19,N_9376,N_9042);
and UO_20 (O_20,N_9523,N_9913);
nand UO_21 (O_21,N_8547,N_9688);
nor UO_22 (O_22,N_9766,N_9126);
nand UO_23 (O_23,N_8210,N_8483);
and UO_24 (O_24,N_8687,N_8004);
nand UO_25 (O_25,N_8383,N_8522);
nand UO_26 (O_26,N_9866,N_9074);
nor UO_27 (O_27,N_9374,N_8195);
nand UO_28 (O_28,N_8647,N_8075);
nor UO_29 (O_29,N_9491,N_9787);
nor UO_30 (O_30,N_9436,N_8400);
or UO_31 (O_31,N_8612,N_9564);
nor UO_32 (O_32,N_8366,N_9156);
nor UO_33 (O_33,N_8358,N_9753);
or UO_34 (O_34,N_8623,N_8846);
or UO_35 (O_35,N_9459,N_9656);
and UO_36 (O_36,N_8182,N_9396);
nand UO_37 (O_37,N_8713,N_9957);
nand UO_38 (O_38,N_9245,N_8037);
or UO_39 (O_39,N_8450,N_8901);
nand UO_40 (O_40,N_9867,N_8564);
or UO_41 (O_41,N_9088,N_8590);
nand UO_42 (O_42,N_9676,N_8954);
nor UO_43 (O_43,N_8947,N_8094);
nand UO_44 (O_44,N_9673,N_8257);
nor UO_45 (O_45,N_8938,N_9535);
nor UO_46 (O_46,N_9743,N_8786);
nand UO_47 (O_47,N_8645,N_9257);
or UO_48 (O_48,N_8021,N_8263);
nand UO_49 (O_49,N_8598,N_9580);
and UO_50 (O_50,N_9319,N_8142);
and UO_51 (O_51,N_9697,N_9882);
nand UO_52 (O_52,N_9721,N_8085);
and UO_53 (O_53,N_9557,N_8951);
and UO_54 (O_54,N_9298,N_8272);
nor UO_55 (O_55,N_8720,N_9442);
or UO_56 (O_56,N_8513,N_8144);
nor UO_57 (O_57,N_8386,N_9754);
or UO_58 (O_58,N_9448,N_9487);
nand UO_59 (O_59,N_9776,N_9972);
nor UO_60 (O_60,N_9460,N_9799);
or UO_61 (O_61,N_8517,N_8099);
or UO_62 (O_62,N_8493,N_8068);
nand UO_63 (O_63,N_9716,N_8036);
nand UO_64 (O_64,N_8923,N_9143);
or UO_65 (O_65,N_9553,N_9043);
nand UO_66 (O_66,N_9503,N_8545);
and UO_67 (O_67,N_8092,N_9102);
and UO_68 (O_68,N_9624,N_8836);
and UO_69 (O_69,N_8763,N_8113);
nand UO_70 (O_70,N_9828,N_8666);
nor UO_71 (O_71,N_9424,N_9652);
and UO_72 (O_72,N_9416,N_8867);
or UO_73 (O_73,N_9420,N_8999);
or UO_74 (O_74,N_8540,N_8189);
nand UO_75 (O_75,N_8319,N_9609);
nor UO_76 (O_76,N_9663,N_8976);
or UO_77 (O_77,N_9452,N_8245);
or UO_78 (O_78,N_9014,N_9922);
nand UO_79 (O_79,N_9324,N_8172);
nor UO_80 (O_80,N_8697,N_9163);
xor UO_81 (O_81,N_8409,N_9060);
nand UO_82 (O_82,N_9525,N_8344);
nand UO_83 (O_83,N_9002,N_9215);
nand UO_84 (O_84,N_8180,N_8577);
nand UO_85 (O_85,N_8834,N_9870);
nand UO_86 (O_86,N_8163,N_8660);
nor UO_87 (O_87,N_8240,N_8445);
nor UO_88 (O_88,N_8485,N_8056);
and UO_89 (O_89,N_9615,N_9836);
or UO_90 (O_90,N_9197,N_9133);
nor UO_91 (O_91,N_8561,N_9194);
nor UO_92 (O_92,N_8716,N_9006);
xor UO_93 (O_93,N_9250,N_8979);
and UO_94 (O_94,N_8132,N_9978);
and UO_95 (O_95,N_8468,N_8842);
or UO_96 (O_96,N_9025,N_9207);
or UO_97 (O_97,N_8915,N_9864);
xnor UO_98 (O_98,N_8550,N_8223);
nand UO_99 (O_99,N_8749,N_9449);
nor UO_100 (O_100,N_8531,N_8760);
nand UO_101 (O_101,N_8397,N_8801);
nor UO_102 (O_102,N_8143,N_8331);
and UO_103 (O_103,N_8093,N_9367);
and UO_104 (O_104,N_9522,N_9405);
or UO_105 (O_105,N_9255,N_9486);
nor UO_106 (O_106,N_8110,N_9686);
and UO_107 (O_107,N_8605,N_9940);
or UO_108 (O_108,N_9954,N_8424);
nor UO_109 (O_109,N_8086,N_9480);
nand UO_110 (O_110,N_8548,N_8129);
and UO_111 (O_111,N_8352,N_9783);
nand UO_112 (O_112,N_8084,N_8309);
nand UO_113 (O_113,N_8768,N_8948);
and UO_114 (O_114,N_8511,N_9444);
or UO_115 (O_115,N_8524,N_9248);
and UO_116 (O_116,N_8261,N_8753);
nand UO_117 (O_117,N_8650,N_9413);
or UO_118 (O_118,N_8334,N_8364);
nor UO_119 (O_119,N_8233,N_9835);
nand UO_120 (O_120,N_9187,N_9506);
or UO_121 (O_121,N_9020,N_9058);
nand UO_122 (O_122,N_9033,N_8726);
and UO_123 (O_123,N_8600,N_9908);
nor UO_124 (O_124,N_9850,N_9203);
and UO_125 (O_125,N_9297,N_9756);
and UO_126 (O_126,N_9962,N_8042);
or UO_127 (O_127,N_9305,N_8480);
nor UO_128 (O_128,N_9176,N_9230);
and UO_129 (O_129,N_8870,N_9479);
nand UO_130 (O_130,N_9740,N_8961);
nor UO_131 (O_131,N_9802,N_8608);
nand UO_132 (O_132,N_8474,N_9899);
or UO_133 (O_133,N_8573,N_8487);
or UO_134 (O_134,N_8422,N_9131);
nor UO_135 (O_135,N_8494,N_8847);
or UO_136 (O_136,N_8964,N_9582);
or UO_137 (O_137,N_8446,N_8609);
nand UO_138 (O_138,N_9969,N_8554);
nor UO_139 (O_139,N_9572,N_8530);
nand UO_140 (O_140,N_8669,N_9004);
nor UO_141 (O_141,N_9808,N_9590);
and UO_142 (O_142,N_8664,N_9816);
and UO_143 (O_143,N_9272,N_8339);
nand UO_144 (O_144,N_8677,N_9847);
nand UO_145 (O_145,N_9161,N_9897);
and UO_146 (O_146,N_9046,N_9344);
or UO_147 (O_147,N_9340,N_8162);
nand UO_148 (O_148,N_8962,N_9251);
and UO_149 (O_149,N_8367,N_8398);
and UO_150 (O_150,N_8791,N_9650);
and UO_151 (O_151,N_8719,N_9429);
or UO_152 (O_152,N_9527,N_9169);
nor UO_153 (O_153,N_9072,N_8823);
nand UO_154 (O_154,N_9308,N_9118);
nor UO_155 (O_155,N_9596,N_8733);
nor UO_156 (O_156,N_9225,N_8774);
xnor UO_157 (O_157,N_9093,N_8102);
nor UO_158 (O_158,N_9139,N_8020);
nor UO_159 (O_159,N_8298,N_9682);
or UO_160 (O_160,N_9414,N_8735);
and UO_161 (O_161,N_9439,N_9037);
nand UO_162 (O_162,N_9270,N_8769);
nand UO_163 (O_163,N_9874,N_8009);
and UO_164 (O_164,N_8333,N_9415);
nand UO_165 (O_165,N_9375,N_8491);
nand UO_166 (O_166,N_8552,N_9877);
xnor UO_167 (O_167,N_8526,N_9310);
or UO_168 (O_168,N_8899,N_8795);
and UO_169 (O_169,N_9497,N_8244);
nor UO_170 (O_170,N_9819,N_9268);
nand UO_171 (O_171,N_8296,N_9026);
and UO_172 (O_172,N_9158,N_8676);
nand UO_173 (O_173,N_8855,N_9629);
nand UO_174 (O_174,N_9604,N_8934);
nand UO_175 (O_175,N_9979,N_8439);
nor UO_176 (O_176,N_8066,N_8698);
nand UO_177 (O_177,N_9066,N_9385);
nand UO_178 (O_178,N_9185,N_9354);
and UO_179 (O_179,N_9280,N_8630);
nand UO_180 (O_180,N_8978,N_9794);
and UO_181 (O_181,N_9705,N_8595);
nor UO_182 (O_182,N_8335,N_9791);
or UO_183 (O_183,N_9019,N_9181);
nand UO_184 (O_184,N_9910,N_8140);
and UO_185 (O_185,N_8740,N_9373);
nand UO_186 (O_186,N_9992,N_8931);
and UO_187 (O_187,N_9703,N_9923);
nand UO_188 (O_188,N_8765,N_9763);
or UO_189 (O_189,N_9392,N_8465);
nor UO_190 (O_190,N_9390,N_8024);
or UO_191 (O_191,N_9315,N_9346);
nor UO_192 (O_192,N_8844,N_8407);
or UO_193 (O_193,N_8481,N_8202);
or UO_194 (O_194,N_8062,N_8933);
or UO_195 (O_195,N_8861,N_9583);
nor UO_196 (O_196,N_9758,N_8019);
nand UO_197 (O_197,N_9638,N_9709);
and UO_198 (O_198,N_8370,N_8534);
nor UO_199 (O_199,N_9613,N_9691);
nand UO_200 (O_200,N_8939,N_8303);
or UO_201 (O_201,N_9653,N_8813);
nand UO_202 (O_202,N_9744,N_9332);
and UO_203 (O_203,N_8411,N_8808);
nor UO_204 (O_204,N_9115,N_8696);
nor UO_205 (O_205,N_8575,N_8067);
nor UO_206 (O_206,N_8260,N_9664);
and UO_207 (O_207,N_8940,N_9353);
or UO_208 (O_208,N_8586,N_9614);
and UO_209 (O_209,N_9745,N_9801);
nor UO_210 (O_210,N_8375,N_8796);
or UO_211 (O_211,N_8516,N_8389);
and UO_212 (O_212,N_9595,N_9488);
or UO_213 (O_213,N_8404,N_8259);
nor UO_214 (O_214,N_9274,N_8098);
nand UO_215 (O_215,N_8826,N_9575);
nor UO_216 (O_216,N_8845,N_8116);
or UO_217 (O_217,N_8248,N_8741);
and UO_218 (O_218,N_9199,N_9235);
or UO_219 (O_219,N_8184,N_9967);
nor UO_220 (O_220,N_9734,N_8185);
or UO_221 (O_221,N_9679,N_9868);
or UO_222 (O_222,N_9350,N_9528);
xnor UO_223 (O_223,N_8584,N_9127);
nand UO_224 (O_224,N_8044,N_8512);
nand UO_225 (O_225,N_9101,N_9496);
and UO_226 (O_226,N_9643,N_8641);
nor UO_227 (O_227,N_9533,N_9030);
or UO_228 (O_228,N_9063,N_9232);
nor UO_229 (O_229,N_9660,N_8253);
nor UO_230 (O_230,N_9265,N_8510);
nand UO_231 (O_231,N_9306,N_9473);
and UO_232 (O_232,N_8117,N_8015);
nor UO_233 (O_233,N_8835,N_9524);
and UO_234 (O_234,N_9012,N_9362);
nand UO_235 (O_235,N_8880,N_9100);
and UO_236 (O_236,N_8466,N_8072);
nand UO_237 (O_237,N_8262,N_9116);
and UO_238 (O_238,N_9944,N_9494);
or UO_239 (O_239,N_8755,N_8320);
and UO_240 (O_240,N_8998,N_9994);
nor UO_241 (O_241,N_8187,N_8077);
or UO_242 (O_242,N_9337,N_9851);
or UO_243 (O_243,N_9044,N_8891);
and UO_244 (O_244,N_8342,N_8239);
and UO_245 (O_245,N_8179,N_8960);
xnor UO_246 (O_246,N_8728,N_9206);
and UO_247 (O_247,N_9515,N_9051);
nor UO_248 (O_248,N_8448,N_9379);
or UO_249 (O_249,N_9343,N_9603);
nand UO_250 (O_250,N_9455,N_8599);
or UO_251 (O_251,N_8385,N_8781);
nand UO_252 (O_252,N_8498,N_9184);
nand UO_253 (O_253,N_9857,N_8509);
nand UO_254 (O_254,N_8237,N_8246);
nor UO_255 (O_255,N_9739,N_8393);
nand UO_256 (O_256,N_9351,N_9669);
nor UO_257 (O_257,N_9567,N_8887);
or UO_258 (O_258,N_8652,N_9084);
or UO_259 (O_259,N_9241,N_8913);
and UO_260 (O_260,N_8274,N_9099);
nor UO_261 (O_261,N_9382,N_8391);
nand UO_262 (O_262,N_9451,N_8292);
or UO_263 (O_263,N_8349,N_9065);
and UO_264 (O_264,N_9466,N_8046);
nor UO_265 (O_265,N_8316,N_8069);
and UO_266 (O_266,N_8152,N_9710);
nand UO_267 (O_267,N_9433,N_9138);
and UO_268 (O_268,N_9500,N_9469);
or UO_269 (O_269,N_9825,N_8369);
and UO_270 (O_270,N_8689,N_9408);
nor UO_271 (O_271,N_9894,N_8784);
or UO_272 (O_272,N_9948,N_9893);
nand UO_273 (O_273,N_8145,N_9177);
and UO_274 (O_274,N_9907,N_8432);
and UO_275 (O_275,N_8295,N_8321);
nand UO_276 (O_276,N_8308,N_8155);
nand UO_277 (O_277,N_9035,N_9589);
nand UO_278 (O_278,N_8161,N_8384);
xor UO_279 (O_279,N_9934,N_9339);
nor UO_280 (O_280,N_9117,N_8387);
nand UO_281 (O_281,N_9314,N_9841);
and UO_282 (O_282,N_8473,N_8247);
nor UO_283 (O_283,N_9210,N_8057);
nand UO_284 (O_284,N_9292,N_9123);
or UO_285 (O_285,N_8751,N_9722);
nor UO_286 (O_286,N_9789,N_8475);
nor UO_287 (O_287,N_9165,N_8770);
and UO_288 (O_288,N_8105,N_8382);
nand UO_289 (O_289,N_9316,N_8614);
nor UO_290 (O_290,N_8528,N_8154);
and UO_291 (O_291,N_9057,N_9964);
nor UO_292 (O_292,N_8275,N_8394);
nand UO_293 (O_293,N_8089,N_8956);
nand UO_294 (O_294,N_9038,N_8074);
nor UO_295 (O_295,N_8508,N_9563);
nand UO_296 (O_296,N_9208,N_9713);
nand UO_297 (O_297,N_8699,N_9718);
xnor UO_298 (O_298,N_8307,N_9036);
nor UO_299 (O_299,N_8455,N_9179);
nand UO_300 (O_300,N_8678,N_8563);
nand UO_301 (O_301,N_8114,N_9700);
nand UO_302 (O_302,N_8100,N_9174);
nand UO_303 (O_303,N_9406,N_9788);
nor UO_304 (O_304,N_9013,N_8279);
nand UO_305 (O_305,N_8843,N_8865);
and UO_306 (O_306,N_8277,N_9891);
nand UO_307 (O_307,N_8156,N_8425);
or UO_308 (O_308,N_9790,N_8365);
nand UO_309 (O_309,N_9837,N_8827);
xor UO_310 (O_310,N_9689,N_9103);
nand UO_311 (O_311,N_9201,N_9547);
nor UO_312 (O_312,N_8556,N_8220);
nor UO_313 (O_313,N_8983,N_9386);
and UO_314 (O_314,N_8695,N_9634);
nand UO_315 (O_315,N_8723,N_8249);
and UO_316 (O_316,N_8986,N_8111);
and UO_317 (O_317,N_9097,N_9467);
nor UO_318 (O_318,N_8871,N_8892);
nand UO_319 (O_319,N_9707,N_9956);
or UO_320 (O_320,N_9640,N_9380);
or UO_321 (O_321,N_9843,N_8588);
nand UO_322 (O_322,N_9782,N_8926);
nand UO_323 (O_323,N_9389,N_9434);
nand UO_324 (O_324,N_9630,N_9885);
nor UO_325 (O_325,N_8969,N_8766);
or UO_326 (O_326,N_9917,N_8756);
and UO_327 (O_327,N_8051,N_9735);
nand UO_328 (O_328,N_8872,N_8306);
and UO_329 (O_329,N_9261,N_9147);
xnor UO_330 (O_330,N_8081,N_8743);
nand UO_331 (O_331,N_8284,N_8718);
xor UO_332 (O_332,N_9173,N_8736);
and UO_333 (O_333,N_8591,N_8064);
and UO_334 (O_334,N_8711,N_9627);
nor UO_335 (O_335,N_9510,N_9973);
nor UO_336 (O_336,N_9062,N_9508);
and UO_337 (O_337,N_9205,N_8441);
nand UO_338 (O_338,N_9921,N_8967);
nor UO_339 (O_339,N_9202,N_9402);
or UO_340 (O_340,N_8615,N_8542);
or UO_341 (O_341,N_8514,N_9087);
and UO_342 (O_342,N_8930,N_8975);
and UO_343 (O_343,N_8109,N_8778);
and UO_344 (O_344,N_9661,N_9170);
and UO_345 (O_345,N_9136,N_9293);
nand UO_346 (O_346,N_9727,N_8443);
nand UO_347 (O_347,N_8235,N_8710);
or UO_348 (O_348,N_9311,N_8839);
nand UO_349 (O_349,N_9421,N_8750);
nor UO_350 (O_350,N_9931,N_9677);
and UO_351 (O_351,N_8038,N_8638);
and UO_352 (O_352,N_8170,N_9246);
nand UO_353 (O_353,N_8875,N_9073);
nand UO_354 (O_354,N_9279,N_8492);
nor UO_355 (O_355,N_9809,N_8764);
or UO_356 (O_356,N_8070,N_9276);
and UO_357 (O_357,N_8582,N_8538);
nand UO_358 (O_358,N_9585,N_8587);
or UO_359 (O_359,N_8372,N_9098);
xor UO_360 (O_360,N_8014,N_9914);
or UO_361 (O_361,N_9254,N_9334);
xor UO_362 (O_362,N_9342,N_9329);
and UO_363 (O_363,N_9372,N_8746);
nand UO_364 (O_364,N_9273,N_9492);
nand UO_365 (O_365,N_8000,N_9818);
and UO_366 (O_366,N_8862,N_9731);
xnor UO_367 (O_367,N_9426,N_9071);
nand UO_368 (O_368,N_9880,N_8819);
nand UO_369 (O_369,N_9681,N_8131);
or UO_370 (O_370,N_8635,N_9626);
nor UO_371 (O_371,N_9050,N_9095);
or UO_372 (O_372,N_9569,N_8535);
and UO_373 (O_373,N_8251,N_8456);
nand UO_374 (O_374,N_8022,N_8414);
nor UO_375 (O_375,N_8974,N_8644);
and UO_376 (O_376,N_9011,N_8779);
nor UO_377 (O_377,N_9995,N_8035);
nor UO_378 (O_378,N_8150,N_9404);
or UO_379 (O_379,N_9848,N_8374);
xnor UO_380 (O_380,N_8201,N_8027);
and UO_381 (O_381,N_8579,N_9238);
nor UO_382 (O_382,N_9154,N_9412);
nand UO_383 (O_383,N_8621,N_8204);
or UO_384 (O_384,N_8228,N_9243);
and UO_385 (O_385,N_9312,N_9089);
or UO_386 (O_386,N_9212,N_9277);
or UO_387 (O_387,N_9440,N_9619);
nor UO_388 (O_388,N_8482,N_9925);
or UO_389 (O_389,N_9064,N_8215);
nand UO_390 (O_390,N_9128,N_9015);
nand UO_391 (O_391,N_8671,N_9083);
and UO_392 (O_392,N_8953,N_8017);
nand UO_393 (O_393,N_9132,N_9916);
and UO_394 (O_394,N_9091,N_9129);
or UO_395 (O_395,N_8328,N_9384);
and UO_396 (O_396,N_8023,N_9383);
nor UO_397 (O_397,N_9331,N_9550);
or UO_398 (O_398,N_9952,N_8405);
nand UO_399 (O_399,N_8783,N_9330);
nor UO_400 (O_400,N_8620,N_8809);
and UO_401 (O_401,N_9516,N_9221);
nor UO_402 (O_402,N_9621,N_9023);
or UO_403 (O_403,N_9628,N_9474);
and UO_404 (O_404,N_8903,N_9168);
or UO_405 (O_405,N_9090,N_8060);
and UO_406 (O_406,N_9937,N_9949);
and UO_407 (O_407,N_9418,N_9253);
and UO_408 (O_408,N_9287,N_8618);
and UO_409 (O_409,N_8151,N_8636);
nand UO_410 (O_410,N_8838,N_9844);
and UO_411 (O_411,N_8196,N_8507);
nand UO_412 (O_412,N_9755,N_9104);
and UO_413 (O_413,N_8218,N_8885);
nand UO_414 (O_414,N_8558,N_8199);
nor UO_415 (O_415,N_8583,N_9796);
and UO_416 (O_416,N_9632,N_9566);
or UO_417 (O_417,N_8932,N_8176);
nand UO_418 (O_418,N_9605,N_8360);
xnor UO_419 (O_419,N_9081,N_9381);
nor UO_420 (O_420,N_9183,N_9399);
or UO_421 (O_421,N_9887,N_9764);
nand UO_422 (O_422,N_9548,N_8458);
nor UO_423 (O_423,N_8757,N_8704);
nor UO_424 (O_424,N_8104,N_8434);
nor UO_425 (O_425,N_9368,N_9435);
nand UO_426 (O_426,N_8688,N_9456);
nand UO_427 (O_427,N_8440,N_9120);
or UO_428 (O_428,N_9358,N_8078);
or UO_429 (O_429,N_9545,N_8700);
nand UO_430 (O_430,N_8868,N_8970);
nor UO_431 (O_431,N_8002,N_9651);
or UO_432 (O_432,N_9027,N_9996);
or UO_433 (O_433,N_8634,N_8079);
xnor UO_434 (O_434,N_9647,N_9574);
nor UO_435 (O_435,N_8153,N_8381);
or UO_436 (O_436,N_9049,N_8639);
and UO_437 (O_437,N_8811,N_8478);
nor UO_438 (O_438,N_8602,N_8546);
nor UO_439 (O_439,N_9539,N_9771);
nand UO_440 (O_440,N_8217,N_9370);
nand UO_441 (O_441,N_9839,N_8911);
or UO_442 (O_442,N_8996,N_9294);
and UO_443 (O_443,N_9291,N_9259);
nor UO_444 (O_444,N_9483,N_8410);
and UO_445 (O_445,N_8082,N_9834);
nand UO_446 (O_446,N_9611,N_8603);
nand UO_447 (O_447,N_9124,N_9662);
nor UO_448 (O_448,N_8581,N_8992);
and UO_449 (O_449,N_8841,N_9450);
nand UO_450 (O_450,N_8570,N_8812);
nand UO_451 (O_451,N_8830,N_9902);
xor UO_452 (O_452,N_8601,N_9388);
nor UO_453 (O_453,N_8506,N_8562);
or UO_454 (O_454,N_8649,N_9461);
and UO_455 (O_455,N_9854,N_8536);
and UO_456 (O_456,N_8869,N_9470);
nor UO_457 (O_457,N_8555,N_9729);
nand UO_458 (O_458,N_8447,N_8864);
or UO_459 (O_459,N_9130,N_9264);
nand UO_460 (O_460,N_8252,N_9878);
nand UO_461 (O_461,N_9657,N_8322);
nand UO_462 (O_462,N_8238,N_9457);
and UO_463 (O_463,N_9005,N_8617);
nor UO_464 (O_464,N_9976,N_9875);
xor UO_465 (O_465,N_8681,N_9558);
and UO_466 (O_466,N_9021,N_9706);
and UO_467 (O_467,N_8922,N_8884);
xor UO_468 (O_468,N_8423,N_8123);
or UO_469 (O_469,N_9410,N_8918);
nand UO_470 (O_470,N_9821,N_8628);
and UO_471 (O_471,N_9031,N_8462);
and UO_472 (O_472,N_8065,N_9338);
nand UO_473 (O_473,N_8258,N_8866);
or UO_474 (O_474,N_9182,N_9003);
nand UO_475 (O_475,N_8775,N_9366);
nand UO_476 (O_476,N_9053,N_8148);
or UO_477 (O_477,N_9529,N_9017);
nor UO_478 (O_478,N_9447,N_8003);
xnor UO_479 (O_479,N_9419,N_9371);
nand UO_480 (O_480,N_8090,N_8442);
nand UO_481 (O_481,N_9040,N_8661);
nand UO_482 (O_482,N_9556,N_9430);
nor UO_483 (O_483,N_9725,N_9690);
nor UO_484 (O_484,N_9471,N_8788);
and UO_485 (O_485,N_9534,N_9200);
nand UO_486 (O_486,N_8016,N_9930);
and UO_487 (O_487,N_8164,N_8594);
nand UO_488 (O_488,N_8988,N_8457);
and UO_489 (O_489,N_9610,N_8273);
or UO_490 (O_490,N_9059,N_9365);
nor UO_491 (O_491,N_9283,N_8031);
nor UO_492 (O_492,N_9458,N_9991);
nor UO_493 (O_493,N_9047,N_8327);
nand UO_494 (O_494,N_8255,N_9724);
nand UO_495 (O_495,N_9938,N_8361);
nor UO_496 (O_496,N_8011,N_9759);
nand UO_497 (O_497,N_8340,N_9812);
or UO_498 (O_498,N_9317,N_9299);
nand UO_499 (O_499,N_8730,N_8917);
or UO_500 (O_500,N_8054,N_9649);
nor UO_501 (O_501,N_8592,N_8006);
nand UO_502 (O_502,N_8290,N_9271);
nor UO_503 (O_503,N_9654,N_9094);
nor UO_504 (O_504,N_8236,N_9587);
nand UO_505 (O_505,N_8990,N_8902);
and UO_506 (O_506,N_9856,N_8504);
or UO_507 (O_507,N_9321,N_8205);
nor UO_508 (O_508,N_9432,N_8727);
nor UO_509 (O_509,N_9975,N_9428);
nor UO_510 (O_510,N_9501,N_8269);
xnor UO_511 (O_511,N_9927,N_8807);
nor UO_512 (O_512,N_9041,N_9813);
nor UO_513 (O_513,N_9263,N_8348);
or UO_514 (O_514,N_9167,N_8831);
and UO_515 (O_515,N_8413,N_8420);
or UO_516 (O_516,N_9318,N_9438);
or UO_517 (O_517,N_8544,N_9701);
nor UO_518 (O_518,N_9307,N_8373);
and UO_519 (O_519,N_9135,N_8080);
and UO_520 (O_520,N_8392,N_8668);
nor UO_521 (O_521,N_8095,N_9209);
and UO_522 (O_522,N_9400,N_9175);
and UO_523 (O_523,N_9820,N_8025);
nand UO_524 (O_524,N_8312,N_8833);
or UO_525 (O_525,N_8048,N_9905);
nor UO_526 (O_526,N_9260,N_8188);
or UO_527 (O_527,N_9863,N_8034);
nand UO_528 (O_528,N_8624,N_8174);
nand UO_529 (O_529,N_8908,N_8702);
nor UO_530 (O_530,N_8495,N_9068);
or UO_531 (O_531,N_8567,N_9219);
or UO_532 (O_532,N_9417,N_9303);
and UO_533 (O_533,N_8197,N_9119);
nor UO_534 (O_534,N_9929,N_9869);
nand UO_535 (O_535,N_8496,N_9082);
nor UO_536 (O_536,N_8276,N_9513);
nand UO_537 (O_537,N_8378,N_8910);
and UO_538 (O_538,N_9137,N_9559);
nand UO_539 (O_539,N_9797,N_9198);
or UO_540 (O_540,N_8679,N_9551);
nor UO_541 (O_541,N_9827,N_9981);
or UO_542 (O_542,N_8380,N_8428);
nand UO_543 (O_543,N_8136,N_9092);
nor UO_544 (O_544,N_9234,N_8800);
nand UO_545 (O_545,N_9378,N_8963);
or UO_546 (O_546,N_8744,N_8315);
nor UO_547 (O_547,N_9341,N_9160);
and UO_548 (O_548,N_9592,N_9267);
and UO_549 (O_549,N_9113,N_9369);
nor UO_550 (O_550,N_8229,N_9838);
nor UO_551 (O_551,N_8499,N_8026);
nand UO_552 (O_552,N_8173,N_8941);
nor UO_553 (O_553,N_9240,N_9577);
nor UO_554 (O_554,N_9145,N_9668);
and UO_555 (O_555,N_8565,N_8798);
nor UO_556 (O_556,N_9349,N_8005);
nand UO_557 (O_557,N_9275,N_9639);
nor UO_558 (O_558,N_8805,N_9737);
nand UO_559 (O_559,N_9685,N_8045);
and UO_560 (O_560,N_8777,N_8754);
or UO_561 (O_561,N_8216,N_9561);
nor UO_562 (O_562,N_8359,N_8851);
nand UO_563 (O_563,N_9159,N_9142);
nand UO_564 (O_564,N_8133,N_9853);
xnor UO_565 (O_565,N_9423,N_9886);
or UO_566 (O_566,N_8137,N_8505);
and UO_567 (O_567,N_8527,N_9001);
nor UO_568 (O_568,N_8814,N_8572);
nor UO_569 (O_569,N_8488,N_8463);
nand UO_570 (O_570,N_8231,N_9772);
and UO_571 (O_571,N_8821,N_9069);
and UO_572 (O_572,N_9859,N_8672);
or UO_573 (O_573,N_8049,N_8906);
and UO_574 (O_574,N_9984,N_9554);
nand UO_575 (O_575,N_8477,N_9482);
and UO_576 (O_576,N_8848,N_8178);
or UO_577 (O_577,N_9977,N_9295);
nor UO_578 (O_578,N_9757,N_9919);
nor UO_579 (O_579,N_8033,N_9993);
nand UO_580 (O_580,N_8318,N_9573);
and UO_581 (O_581,N_9407,N_8464);
nor UO_582 (O_582,N_9328,N_8659);
or UO_583 (O_583,N_9546,N_8341);
nand UO_584 (O_584,N_8467,N_9862);
or UO_585 (O_585,N_8460,N_9636);
nand UO_586 (O_586,N_8958,N_8472);
or UO_587 (O_587,N_8437,N_9281);
nor UO_588 (O_588,N_9356,N_9665);
or UO_589 (O_589,N_9171,N_9635);
nand UO_590 (O_590,N_8490,N_9107);
and UO_591 (O_591,N_8076,N_8816);
nand UO_592 (O_592,N_9571,N_8523);
nand UO_593 (O_593,N_9920,N_9552);
and UO_594 (O_594,N_8337,N_8141);
nand UO_595 (O_595,N_9327,N_9323);
xnor UO_596 (O_596,N_8832,N_8782);
nor UO_597 (O_597,N_9623,N_9586);
or UO_598 (O_598,N_9845,N_8310);
or UO_599 (O_599,N_8130,N_8789);
or UO_600 (O_600,N_8149,N_8715);
xnor UO_601 (O_601,N_8304,N_8521);
or UO_602 (O_602,N_9477,N_9108);
nor UO_603 (O_603,N_9218,N_8912);
and UO_604 (O_604,N_8430,N_8018);
and UO_605 (O_605,N_9347,N_9216);
nand UO_606 (O_606,N_8186,N_9646);
nand UO_607 (O_607,N_9749,N_8426);
nor UO_608 (O_608,N_8350,N_8850);
nor UO_609 (O_609,N_8376,N_8278);
nand UO_610 (O_610,N_8643,N_8052);
nor UO_611 (O_611,N_9164,N_9581);
and UO_612 (O_612,N_9555,N_8030);
nand UO_613 (O_613,N_9226,N_9588);
nor UO_614 (O_614,N_9067,N_8053);
nor UO_615 (O_615,N_8363,N_8806);
nand UO_616 (O_616,N_8585,N_8313);
nand UO_617 (O_617,N_9602,N_9075);
or UO_618 (O_618,N_8714,N_8662);
or UO_619 (O_619,N_8732,N_9191);
nand UO_620 (O_620,N_9437,N_8332);
nor UO_621 (O_621,N_9780,N_9824);
or UO_622 (O_622,N_8029,N_8646);
and UO_623 (O_623,N_9531,N_9599);
nor UO_624 (O_624,N_9741,N_9747);
and UO_625 (O_625,N_8725,N_9896);
and UO_626 (O_626,N_8532,N_9672);
and UO_627 (O_627,N_8752,N_9009);
nor UO_628 (O_628,N_8973,N_8627);
nor UO_629 (O_629,N_8890,N_8559);
nand UO_630 (O_630,N_8191,N_9536);
nand UO_631 (O_631,N_8435,N_8722);
xor UO_632 (O_632,N_8007,N_9865);
or UO_633 (O_633,N_8013,N_9965);
nand UO_634 (O_634,N_9288,N_9963);
xor UO_635 (O_635,N_8106,N_8803);
xnor UO_636 (O_636,N_8519,N_8707);
or UO_637 (O_637,N_9711,N_9262);
and UO_638 (O_638,N_8421,N_8950);
nor UO_639 (O_639,N_9830,N_8225);
and UO_640 (O_640,N_8914,N_8171);
nor UO_641 (O_641,N_8470,N_9222);
or UO_642 (O_642,N_8856,N_9730);
or UO_643 (O_643,N_9612,N_8626);
nand UO_644 (O_644,N_9096,N_9016);
nor UO_645 (O_645,N_9542,N_8989);
and UO_646 (O_646,N_9125,N_9178);
nor UO_647 (O_647,N_9022,N_8291);
nand UO_648 (O_648,N_8852,N_9898);
nor UO_649 (O_649,N_9765,N_8267);
or UO_650 (O_650,N_9633,N_8987);
and UO_651 (O_651,N_9909,N_9578);
nand UO_652 (O_652,N_8371,N_9224);
nand UO_653 (O_653,N_8345,N_9490);
nor UO_654 (O_654,N_9512,N_8772);
and UO_655 (O_655,N_9112,N_8972);
and UO_656 (O_656,N_8828,N_9761);
nand UO_657 (O_657,N_8165,N_9793);
and UO_658 (O_658,N_9078,N_8968);
and UO_659 (O_659,N_9947,N_8952);
nand UO_660 (O_660,N_8896,N_9008);
xnor UO_661 (O_661,N_9228,N_8761);
nor UO_662 (O_662,N_8282,N_8347);
nor UO_663 (O_663,N_8670,N_9625);
nor UO_664 (O_664,N_9325,N_9190);
and UO_665 (O_665,N_9694,N_8203);
or UO_666 (O_666,N_9769,N_9833);
nand UO_667 (O_667,N_9355,N_9670);
or UO_668 (O_668,N_8944,N_8166);
nand UO_669 (O_669,N_9666,N_9770);
or UO_670 (O_670,N_8119,N_9695);
nand UO_671 (O_671,N_9562,N_9425);
and UO_672 (O_672,N_9377,N_8857);
nor UO_673 (O_673,N_8955,N_9684);
or UO_674 (O_674,N_8898,N_8667);
and UO_675 (O_675,N_9266,N_9645);
or UO_676 (O_676,N_8604,N_8124);
or UO_677 (O_677,N_9530,N_9777);
nor UO_678 (O_678,N_8616,N_9109);
nand UO_679 (O_679,N_9901,N_8734);
or UO_680 (O_680,N_9683,N_9811);
nand UO_681 (O_681,N_8825,N_8329);
and UO_682 (O_682,N_8936,N_9239);
nand UO_683 (O_683,N_8444,N_9584);
nand UO_684 (O_684,N_8543,N_9803);
nor UO_685 (O_685,N_9805,N_9144);
nor UO_686 (O_686,N_9593,N_8459);
or UO_687 (O_687,N_9540,N_8091);
and UO_688 (O_688,N_8192,N_8121);
or UO_689 (O_689,N_9641,N_8338);
and UO_690 (O_690,N_9814,N_9895);
or UO_691 (O_691,N_8012,N_8860);
and UO_692 (O_692,N_9498,N_8703);
and UO_693 (O_693,N_8357,N_9918);
and UO_694 (O_694,N_9105,N_9153);
nand UO_695 (O_695,N_8146,N_8737);
nand UO_696 (O_696,N_9817,N_8904);
or UO_697 (O_697,N_9961,N_8576);
and UO_698 (O_698,N_8993,N_8351);
nand UO_699 (O_699,N_9720,N_9881);
or UO_700 (O_700,N_8942,N_8745);
and UO_701 (O_701,N_8658,N_8799);
or UO_702 (O_702,N_8680,N_8557);
or UO_703 (O_703,N_8965,N_9393);
nand UO_704 (O_704,N_9541,N_8767);
and UO_705 (O_705,N_8401,N_8227);
nand UO_706 (O_706,N_9950,N_9728);
and UO_707 (O_707,N_9000,N_9618);
nand UO_708 (O_708,N_9900,N_9717);
or UO_709 (O_709,N_8168,N_9284);
nor UO_710 (O_710,N_8484,N_8874);
or UO_711 (O_711,N_8043,N_8921);
or UO_712 (O_712,N_8709,N_8515);
nor UO_713 (O_713,N_8214,N_9086);
and UO_714 (O_714,N_8243,N_9708);
nand UO_715 (O_715,N_9526,N_8541);
nand UO_716 (O_716,N_9903,N_9247);
nor UO_717 (O_717,N_9752,N_8390);
nor UO_718 (O_718,N_9760,N_8115);
or UO_719 (O_719,N_9942,N_8073);
nor UO_720 (O_720,N_8882,N_8818);
nand UO_721 (O_721,N_9464,N_9394);
nor UO_722 (O_722,N_9990,N_8353);
nor UO_723 (O_723,N_9723,N_9778);
nand UO_724 (O_724,N_8580,N_9532);
nor UO_725 (O_725,N_9489,N_8537);
xnor UO_726 (O_726,N_9213,N_8840);
nand UO_727 (O_727,N_9807,N_9671);
or UO_728 (O_728,N_8981,N_8299);
nand UO_729 (O_729,N_8539,N_8047);
or UO_730 (O_730,N_9576,N_8101);
and UO_731 (O_731,N_8317,N_8705);
or UO_732 (O_732,N_9953,N_8731);
nor UO_733 (O_733,N_8927,N_9204);
xor UO_734 (O_734,N_8637,N_9968);
nand UO_735 (O_735,N_8461,N_9704);
or UO_736 (O_736,N_9945,N_8183);
nand UO_737 (O_737,N_8729,N_9076);
nor UO_738 (O_738,N_9823,N_8937);
or UO_739 (O_739,N_9244,N_9077);
xnor UO_740 (O_740,N_8787,N_9152);
and UO_741 (O_741,N_8673,N_9693);
xor UO_742 (O_742,N_8849,N_8001);
or UO_743 (O_743,N_8657,N_8997);
nand UO_744 (O_744,N_8957,N_9622);
or UO_745 (O_745,N_8311,N_8408);
or UO_746 (O_746,N_8226,N_8265);
and UO_747 (O_747,N_8945,N_9122);
and UO_748 (O_748,N_8254,N_8747);
or UO_749 (O_749,N_8395,N_8909);
nor UO_750 (O_750,N_8802,N_9443);
nand UO_751 (O_751,N_9282,N_9180);
or UO_752 (O_752,N_9986,N_8032);
nor UO_753 (O_753,N_9360,N_8596);
or UO_754 (O_754,N_8135,N_8502);
nor UO_755 (O_755,N_8566,N_9166);
or UO_756 (O_756,N_9499,N_9751);
and UO_757 (O_757,N_8041,N_8793);
nand UO_758 (O_758,N_9549,N_9935);
and UO_759 (O_759,N_8438,N_9698);
and UO_760 (O_760,N_8533,N_8881);
xnor UO_761 (O_761,N_8058,N_9514);
and UO_762 (O_762,N_8096,N_9220);
and UO_763 (O_763,N_9696,N_9980);
nand UO_764 (O_764,N_9217,N_8574);
and UO_765 (O_765,N_8578,N_9304);
or UO_766 (O_766,N_9932,N_8211);
nor UO_767 (O_767,N_9056,N_8433);
nor UO_768 (O_768,N_8631,N_9445);
nor UO_769 (O_769,N_8625,N_9223);
or UO_770 (O_770,N_8206,N_9591);
nor UO_771 (O_771,N_8356,N_8589);
or UO_772 (O_772,N_9883,N_8966);
nand UO_773 (O_773,N_9134,N_8055);
or UO_774 (O_774,N_9842,N_8497);
and UO_775 (O_775,N_9936,N_9229);
and UO_776 (O_776,N_8949,N_8549);
xor UO_777 (O_777,N_8792,N_9300);
or UO_778 (O_778,N_9674,N_9594);
nand UO_779 (O_779,N_9876,N_8610);
or UO_780 (O_780,N_9983,N_9278);
and UO_781 (O_781,N_9302,N_8859);
and UO_782 (O_782,N_8234,N_8242);
nor UO_783 (O_783,N_8607,N_9322);
and UO_784 (O_784,N_9079,N_8977);
nand UO_785 (O_785,N_9860,N_8929);
and UO_786 (O_786,N_8919,N_9560);
nor UO_787 (O_787,N_9320,N_9912);
or UO_788 (O_788,N_9463,N_8256);
nand UO_789 (O_789,N_8712,N_8412);
nor UO_790 (O_790,N_9884,N_9242);
and UO_791 (O_791,N_9151,N_8010);
nand UO_792 (O_792,N_9520,N_9462);
and UO_793 (O_793,N_9395,N_8167);
nand UO_794 (O_794,N_8059,N_9061);
and UO_795 (O_795,N_8264,N_8354);
nor UO_796 (O_796,N_8553,N_8685);
nand UO_797 (O_797,N_9422,N_9678);
and UO_798 (O_798,N_9141,N_8452);
nand UO_799 (O_799,N_9411,N_8103);
xnor UO_800 (O_800,N_8209,N_9052);
xor UO_801 (O_801,N_9988,N_9032);
and UO_802 (O_802,N_9773,N_9140);
nand UO_803 (O_803,N_9792,N_9692);
nor UO_804 (O_804,N_8346,N_9601);
nor UO_805 (O_805,N_9840,N_9804);
nand UO_806 (O_806,N_8108,N_9509);
nand UO_807 (O_807,N_9214,N_8655);
nor UO_808 (O_808,N_8980,N_8790);
or UO_809 (O_809,N_8417,N_8873);
nand UO_810 (O_810,N_9810,N_8889);
nor UO_811 (O_811,N_9832,N_8177);
nor UO_812 (O_812,N_8853,N_8717);
or UO_813 (O_813,N_8419,N_9849);
nor UO_814 (O_814,N_8924,N_8824);
nand UO_815 (O_815,N_8742,N_9924);
or UO_816 (O_816,N_9326,N_9762);
nor UO_817 (O_817,N_8281,N_9748);
nor UO_818 (O_818,N_9286,N_9502);
nand UO_819 (O_819,N_8040,N_8886);
and UO_820 (O_820,N_9114,N_9237);
nor UO_821 (O_821,N_9364,N_9733);
or UO_822 (O_822,N_9781,N_8593);
and UO_823 (O_823,N_8138,N_8039);
or UO_824 (O_824,N_8928,N_9946);
and UO_825 (O_825,N_9333,N_9999);
and UO_826 (O_826,N_9403,N_8406);
nor UO_827 (O_827,N_9504,N_9829);
and UO_828 (O_828,N_8230,N_9659);
nor UO_829 (O_829,N_8693,N_8280);
and UO_830 (O_830,N_9345,N_8648);
or UO_831 (O_831,N_8893,N_9507);
nand UO_832 (O_832,N_8479,N_9941);
nand UO_833 (O_833,N_8324,N_9401);
nor UO_834 (O_834,N_9029,N_9468);
nor UO_835 (O_835,N_9648,N_9409);
or UO_836 (O_836,N_8190,N_9775);
nor UO_837 (O_837,N_9675,N_9750);
and UO_838 (O_838,N_8355,N_9441);
and UO_839 (O_839,N_8415,N_8213);
xor UO_840 (O_840,N_9888,N_8569);
xor UO_841 (O_841,N_8431,N_9680);
nor UO_842 (O_842,N_8994,N_8436);
and UO_843 (O_843,N_9106,N_8748);
nor UO_844 (O_844,N_9822,N_8287);
xnor UO_845 (O_845,N_9667,N_9768);
and UO_846 (O_846,N_9475,N_8118);
nand UO_847 (O_847,N_8396,N_9786);
nand UO_848 (O_848,N_8837,N_9454);
and UO_849 (O_849,N_9699,N_8122);
nor UO_850 (O_850,N_8794,N_8785);
xor UO_851 (O_851,N_8453,N_9070);
nor UO_852 (O_852,N_8854,N_8403);
nor UO_853 (O_853,N_8503,N_9597);
and UO_854 (O_854,N_8560,N_9798);
and UO_855 (O_855,N_8829,N_9966);
or UO_856 (O_856,N_8200,N_8674);
or UO_857 (O_857,N_8762,N_9431);
or UO_858 (O_858,N_8489,N_8694);
or UO_859 (O_859,N_9958,N_8971);
xor UO_860 (O_860,N_8858,N_8721);
or UO_861 (O_861,N_8221,N_8427);
nand UO_862 (O_862,N_8863,N_8181);
nand UO_863 (O_863,N_8325,N_8271);
and UO_864 (O_864,N_8061,N_9495);
nor UO_865 (O_865,N_9568,N_8613);
or UO_866 (O_866,N_9195,N_9906);
nand UO_867 (O_867,N_9121,N_8330);
and UO_868 (O_868,N_9010,N_9543);
or UO_869 (O_869,N_8194,N_9858);
nand UO_870 (O_870,N_9915,N_8139);
nand UO_871 (O_871,N_8283,N_8399);
nor UO_872 (O_872,N_8501,N_9048);
and UO_873 (O_873,N_9517,N_9359);
and UO_874 (O_874,N_9719,N_9687);
nand UO_875 (O_875,N_8362,N_9034);
and UO_876 (O_876,N_8418,N_8551);
nor UO_877 (O_877,N_9055,N_8336);
nor UO_878 (O_878,N_9738,N_8301);
xor UO_879 (O_879,N_9655,N_9544);
and UO_880 (O_880,N_8175,N_8815);
or UO_881 (O_881,N_8916,N_8429);
and UO_882 (O_882,N_9774,N_9348);
and UO_883 (O_883,N_8897,N_8288);
nand UO_884 (O_884,N_9110,N_8198);
and UO_885 (O_885,N_8071,N_8159);
nand UO_886 (O_886,N_8402,N_9398);
or UO_887 (O_887,N_8879,N_9846);
nor UO_888 (O_888,N_9644,N_8083);
or UO_889 (O_889,N_8097,N_8776);
or UO_890 (O_890,N_9269,N_8241);
and UO_891 (O_891,N_8876,N_9926);
nand UO_892 (O_892,N_9800,N_9714);
nand UO_893 (O_893,N_8471,N_8571);
and UO_894 (O_894,N_8469,N_8654);
nand UO_895 (O_895,N_8653,N_9039);
nand UO_896 (O_896,N_9249,N_9974);
or UO_897 (O_897,N_9361,N_8293);
nand UO_898 (O_898,N_8804,N_9427);
nand UO_899 (O_899,N_8125,N_9742);
nand UO_900 (O_900,N_9608,N_8388);
or UO_901 (O_901,N_9537,N_8690);
and UO_902 (O_902,N_8294,N_8810);
nor UO_903 (O_903,N_8632,N_8127);
or UO_904 (O_904,N_9732,N_9080);
nand UO_905 (O_905,N_8894,N_9971);
xor UO_906 (O_906,N_8326,N_9872);
and UO_907 (O_907,N_9795,N_9149);
nand UO_908 (O_908,N_9943,N_8270);
nand UO_909 (O_909,N_8907,N_8112);
or UO_910 (O_910,N_8368,N_9712);
nand UO_911 (O_911,N_8232,N_9335);
or UO_912 (O_912,N_8991,N_8691);
nor UO_913 (O_913,N_9148,N_9889);
nor UO_914 (O_914,N_8266,N_9997);
and UO_915 (O_915,N_9702,N_9024);
nand UO_916 (O_916,N_9481,N_8629);
nor UO_917 (O_917,N_8300,N_9256);
and UO_918 (O_918,N_9472,N_8250);
nor UO_919 (O_919,N_9620,N_8486);
and UO_920 (O_920,N_9911,N_9054);
or UO_921 (O_921,N_8985,N_8701);
and UO_922 (O_922,N_9157,N_9642);
nor UO_923 (O_923,N_8771,N_9476);
and UO_924 (O_924,N_9186,N_8169);
nor UO_925 (O_925,N_8797,N_9465);
nor UO_926 (O_926,N_8050,N_8379);
and UO_927 (O_927,N_8451,N_8665);
nand UO_928 (O_928,N_8314,N_9085);
nor UO_929 (O_929,N_9028,N_9617);
nand UO_930 (O_930,N_8323,N_8633);
nand UO_931 (O_931,N_8959,N_8268);
nor UO_932 (O_932,N_8692,N_8212);
and UO_933 (O_933,N_8302,N_9387);
and UO_934 (O_934,N_9785,N_8682);
and UO_935 (O_935,N_9726,N_9658);
or UO_936 (O_936,N_9861,N_9970);
or UO_937 (O_937,N_9933,N_8285);
nand UO_938 (O_938,N_9928,N_9616);
nor UO_939 (O_939,N_8158,N_8758);
and UO_940 (O_940,N_9570,N_8449);
or UO_941 (O_941,N_9453,N_9637);
nor UO_942 (O_942,N_9252,N_9784);
nor UO_943 (O_943,N_9227,N_9211);
nor UO_944 (O_944,N_8611,N_8193);
or UO_945 (O_945,N_9007,N_9598);
nor UO_946 (O_946,N_8877,N_9231);
nand UO_947 (O_947,N_8895,N_9746);
nand UO_948 (O_948,N_9363,N_9631);
or UO_949 (O_949,N_8219,N_9478);
and UO_950 (O_950,N_8120,N_9045);
nand UO_951 (O_951,N_9309,N_9600);
or UO_952 (O_952,N_8147,N_9806);
or UO_953 (O_953,N_8640,N_8739);
or UO_954 (O_954,N_8619,N_9258);
or UO_955 (O_955,N_9767,N_8773);
and UO_956 (O_956,N_9951,N_8946);
or UO_957 (O_957,N_9826,N_8208);
nor UO_958 (O_958,N_9357,N_9397);
and UO_959 (O_959,N_9236,N_9296);
nor UO_960 (O_960,N_8297,N_9998);
nand UO_961 (O_961,N_9391,N_9736);
or UO_962 (O_962,N_8642,N_8126);
or UO_963 (O_963,N_9313,N_8982);
nand UO_964 (O_964,N_8900,N_9538);
nor UO_965 (O_965,N_8597,N_8663);
or UO_966 (O_966,N_9579,N_9505);
nor UO_967 (O_967,N_9352,N_8708);
nand UO_968 (O_968,N_8128,N_9155);
nor UO_969 (O_969,N_8878,N_9111);
nor UO_970 (O_970,N_8377,N_9196);
and UO_971 (O_971,N_8568,N_8622);
or UO_972 (O_972,N_9815,N_9484);
nor UO_973 (O_973,N_9892,N_9904);
or UO_974 (O_974,N_8529,N_8305);
or UO_975 (O_975,N_9873,N_9285);
and UO_976 (O_976,N_9955,N_9172);
nor UO_977 (O_977,N_8943,N_8160);
or UO_978 (O_978,N_8651,N_9493);
and UO_979 (O_979,N_8995,N_9192);
nand UO_980 (O_980,N_8724,N_8822);
or UO_981 (O_981,N_9233,N_8157);
nor UO_982 (O_982,N_9982,N_9985);
nand UO_983 (O_983,N_9446,N_9188);
nor UO_984 (O_984,N_9162,N_9289);
nor UO_985 (O_985,N_8500,N_8520);
nand UO_986 (O_986,N_8675,N_8343);
and UO_987 (O_987,N_9336,N_9018);
nor UO_988 (O_988,N_8222,N_9511);
nand UO_989 (O_989,N_8883,N_9715);
and UO_990 (O_990,N_8087,N_9519);
and UO_991 (O_991,N_9146,N_8984);
nand UO_992 (O_992,N_8454,N_8028);
nand UO_993 (O_993,N_8289,N_8780);
and UO_994 (O_994,N_8920,N_8088);
nor UO_995 (O_995,N_9871,N_9521);
nor UO_996 (O_996,N_8935,N_8224);
nand UO_997 (O_997,N_9606,N_8817);
nand UO_998 (O_998,N_8518,N_9150);
and UO_999 (O_999,N_8416,N_8925);
nor UO_1000 (O_1000,N_8559,N_8438);
xnor UO_1001 (O_1001,N_8903,N_9078);
or UO_1002 (O_1002,N_9630,N_8545);
nand UO_1003 (O_1003,N_9613,N_9615);
nand UO_1004 (O_1004,N_9062,N_9251);
nand UO_1005 (O_1005,N_8697,N_8135);
or UO_1006 (O_1006,N_9090,N_8722);
or UO_1007 (O_1007,N_8713,N_9883);
or UO_1008 (O_1008,N_8555,N_8301);
or UO_1009 (O_1009,N_8466,N_9535);
nor UO_1010 (O_1010,N_9905,N_9111);
or UO_1011 (O_1011,N_8693,N_9595);
or UO_1012 (O_1012,N_9148,N_9423);
or UO_1013 (O_1013,N_8615,N_9600);
or UO_1014 (O_1014,N_8403,N_9975);
nand UO_1015 (O_1015,N_9078,N_8536);
and UO_1016 (O_1016,N_8682,N_9232);
nor UO_1017 (O_1017,N_8712,N_8790);
or UO_1018 (O_1018,N_8013,N_8368);
and UO_1019 (O_1019,N_8742,N_9768);
nor UO_1020 (O_1020,N_9946,N_8429);
nor UO_1021 (O_1021,N_9144,N_9268);
nand UO_1022 (O_1022,N_8253,N_9269);
xor UO_1023 (O_1023,N_9730,N_8192);
and UO_1024 (O_1024,N_8138,N_9580);
nand UO_1025 (O_1025,N_8378,N_8524);
nand UO_1026 (O_1026,N_9173,N_9097);
or UO_1027 (O_1027,N_9460,N_8693);
and UO_1028 (O_1028,N_9723,N_8936);
nand UO_1029 (O_1029,N_9505,N_8835);
and UO_1030 (O_1030,N_9811,N_8174);
xnor UO_1031 (O_1031,N_8580,N_8681);
and UO_1032 (O_1032,N_8409,N_8054);
and UO_1033 (O_1033,N_9919,N_8270);
and UO_1034 (O_1034,N_9703,N_8661);
nand UO_1035 (O_1035,N_9688,N_9251);
nand UO_1036 (O_1036,N_8627,N_8665);
nand UO_1037 (O_1037,N_8044,N_8494);
nor UO_1038 (O_1038,N_9238,N_9679);
nand UO_1039 (O_1039,N_8534,N_9086);
and UO_1040 (O_1040,N_8306,N_8824);
and UO_1041 (O_1041,N_9235,N_8783);
nand UO_1042 (O_1042,N_8377,N_9984);
nor UO_1043 (O_1043,N_8411,N_9808);
xnor UO_1044 (O_1044,N_9714,N_9704);
nand UO_1045 (O_1045,N_8010,N_9382);
nand UO_1046 (O_1046,N_9382,N_8612);
xor UO_1047 (O_1047,N_9484,N_8958);
nand UO_1048 (O_1048,N_8679,N_8785);
or UO_1049 (O_1049,N_9384,N_8734);
nand UO_1050 (O_1050,N_8852,N_8221);
nand UO_1051 (O_1051,N_9751,N_8684);
nor UO_1052 (O_1052,N_9827,N_8159);
nor UO_1053 (O_1053,N_9102,N_8373);
nand UO_1054 (O_1054,N_9521,N_9356);
and UO_1055 (O_1055,N_9508,N_9585);
nor UO_1056 (O_1056,N_8605,N_9782);
or UO_1057 (O_1057,N_8142,N_9948);
nor UO_1058 (O_1058,N_8140,N_9564);
nor UO_1059 (O_1059,N_8163,N_8249);
nor UO_1060 (O_1060,N_9336,N_8964);
or UO_1061 (O_1061,N_8299,N_8101);
and UO_1062 (O_1062,N_8212,N_8532);
or UO_1063 (O_1063,N_9958,N_9800);
or UO_1064 (O_1064,N_8840,N_9910);
nor UO_1065 (O_1065,N_8537,N_9995);
and UO_1066 (O_1066,N_9285,N_8015);
or UO_1067 (O_1067,N_8315,N_9604);
and UO_1068 (O_1068,N_9962,N_9568);
nand UO_1069 (O_1069,N_9294,N_8535);
and UO_1070 (O_1070,N_9295,N_8610);
nand UO_1071 (O_1071,N_8347,N_9329);
or UO_1072 (O_1072,N_9593,N_8426);
and UO_1073 (O_1073,N_8598,N_8795);
or UO_1074 (O_1074,N_8696,N_9873);
or UO_1075 (O_1075,N_8968,N_9160);
or UO_1076 (O_1076,N_9328,N_9990);
nor UO_1077 (O_1077,N_9671,N_9759);
nand UO_1078 (O_1078,N_9019,N_8976);
or UO_1079 (O_1079,N_9187,N_8670);
nand UO_1080 (O_1080,N_8600,N_9306);
or UO_1081 (O_1081,N_9375,N_9782);
nor UO_1082 (O_1082,N_8655,N_8828);
and UO_1083 (O_1083,N_8777,N_8034);
and UO_1084 (O_1084,N_9117,N_9597);
nor UO_1085 (O_1085,N_8753,N_9894);
nor UO_1086 (O_1086,N_8406,N_9047);
and UO_1087 (O_1087,N_8007,N_9104);
nor UO_1088 (O_1088,N_9813,N_8148);
or UO_1089 (O_1089,N_9061,N_8896);
and UO_1090 (O_1090,N_8610,N_9983);
nor UO_1091 (O_1091,N_8474,N_9481);
nand UO_1092 (O_1092,N_8473,N_8209);
xor UO_1093 (O_1093,N_8282,N_9409);
nor UO_1094 (O_1094,N_8246,N_9184);
or UO_1095 (O_1095,N_9730,N_9048);
nor UO_1096 (O_1096,N_8914,N_9962);
nor UO_1097 (O_1097,N_8020,N_9686);
and UO_1098 (O_1098,N_9465,N_8490);
and UO_1099 (O_1099,N_8145,N_9937);
nand UO_1100 (O_1100,N_8558,N_9321);
xor UO_1101 (O_1101,N_8556,N_8994);
xnor UO_1102 (O_1102,N_8823,N_8865);
and UO_1103 (O_1103,N_9573,N_9919);
nand UO_1104 (O_1104,N_9521,N_9695);
nand UO_1105 (O_1105,N_9302,N_9247);
or UO_1106 (O_1106,N_9452,N_8827);
or UO_1107 (O_1107,N_8588,N_8561);
or UO_1108 (O_1108,N_9823,N_8235);
and UO_1109 (O_1109,N_8422,N_9783);
nor UO_1110 (O_1110,N_9653,N_9831);
and UO_1111 (O_1111,N_8949,N_9152);
nor UO_1112 (O_1112,N_9742,N_9645);
nand UO_1113 (O_1113,N_9762,N_9933);
and UO_1114 (O_1114,N_8100,N_9595);
nand UO_1115 (O_1115,N_9012,N_9863);
or UO_1116 (O_1116,N_9884,N_8710);
or UO_1117 (O_1117,N_9714,N_8166);
and UO_1118 (O_1118,N_9451,N_9768);
nor UO_1119 (O_1119,N_9602,N_8753);
nand UO_1120 (O_1120,N_8376,N_9092);
nor UO_1121 (O_1121,N_8498,N_8048);
nor UO_1122 (O_1122,N_8727,N_9008);
nand UO_1123 (O_1123,N_9001,N_9963);
nand UO_1124 (O_1124,N_9941,N_8801);
nor UO_1125 (O_1125,N_8598,N_9866);
nand UO_1126 (O_1126,N_9964,N_9401);
nand UO_1127 (O_1127,N_9194,N_8797);
xor UO_1128 (O_1128,N_8307,N_8225);
nor UO_1129 (O_1129,N_8841,N_9175);
nand UO_1130 (O_1130,N_8438,N_9637);
or UO_1131 (O_1131,N_8143,N_9191);
nor UO_1132 (O_1132,N_8500,N_9507);
and UO_1133 (O_1133,N_9467,N_9696);
and UO_1134 (O_1134,N_8857,N_9545);
and UO_1135 (O_1135,N_8527,N_9836);
nand UO_1136 (O_1136,N_8497,N_9701);
nand UO_1137 (O_1137,N_9426,N_9913);
and UO_1138 (O_1138,N_9811,N_8588);
nand UO_1139 (O_1139,N_8854,N_8277);
and UO_1140 (O_1140,N_8756,N_8645);
nor UO_1141 (O_1141,N_9210,N_9203);
nor UO_1142 (O_1142,N_9759,N_9933);
or UO_1143 (O_1143,N_9554,N_8820);
nor UO_1144 (O_1144,N_8415,N_9188);
and UO_1145 (O_1145,N_8110,N_9730);
or UO_1146 (O_1146,N_9629,N_8978);
nand UO_1147 (O_1147,N_9042,N_8800);
and UO_1148 (O_1148,N_9346,N_8261);
nand UO_1149 (O_1149,N_9471,N_9212);
and UO_1150 (O_1150,N_8952,N_8986);
nor UO_1151 (O_1151,N_8875,N_8970);
nand UO_1152 (O_1152,N_8139,N_8474);
or UO_1153 (O_1153,N_8437,N_9148);
and UO_1154 (O_1154,N_9909,N_8926);
or UO_1155 (O_1155,N_9092,N_8750);
or UO_1156 (O_1156,N_8371,N_8257);
or UO_1157 (O_1157,N_9753,N_9738);
nor UO_1158 (O_1158,N_9899,N_9986);
nand UO_1159 (O_1159,N_8290,N_9527);
and UO_1160 (O_1160,N_8670,N_8648);
or UO_1161 (O_1161,N_9625,N_9570);
and UO_1162 (O_1162,N_9276,N_8706);
and UO_1163 (O_1163,N_8434,N_8127);
and UO_1164 (O_1164,N_8225,N_9523);
nand UO_1165 (O_1165,N_9508,N_8389);
nor UO_1166 (O_1166,N_8705,N_8201);
and UO_1167 (O_1167,N_8303,N_8199);
nand UO_1168 (O_1168,N_8376,N_8365);
nor UO_1169 (O_1169,N_9449,N_8503);
or UO_1170 (O_1170,N_8143,N_9683);
and UO_1171 (O_1171,N_9343,N_8501);
nor UO_1172 (O_1172,N_9877,N_8665);
nand UO_1173 (O_1173,N_8715,N_8753);
nand UO_1174 (O_1174,N_8269,N_9591);
nor UO_1175 (O_1175,N_8853,N_8940);
nor UO_1176 (O_1176,N_9722,N_9661);
nor UO_1177 (O_1177,N_8274,N_8535);
or UO_1178 (O_1178,N_8877,N_8187);
nand UO_1179 (O_1179,N_8409,N_9670);
and UO_1180 (O_1180,N_9605,N_9542);
nand UO_1181 (O_1181,N_8963,N_9226);
or UO_1182 (O_1182,N_9276,N_8611);
nand UO_1183 (O_1183,N_9854,N_8735);
nor UO_1184 (O_1184,N_9653,N_9602);
nor UO_1185 (O_1185,N_8891,N_9457);
or UO_1186 (O_1186,N_8152,N_9107);
and UO_1187 (O_1187,N_9319,N_9697);
or UO_1188 (O_1188,N_8789,N_9548);
and UO_1189 (O_1189,N_8393,N_8870);
or UO_1190 (O_1190,N_8988,N_9253);
nor UO_1191 (O_1191,N_9272,N_8853);
and UO_1192 (O_1192,N_9723,N_9898);
or UO_1193 (O_1193,N_9148,N_8514);
nand UO_1194 (O_1194,N_9729,N_9273);
nor UO_1195 (O_1195,N_8278,N_9655);
and UO_1196 (O_1196,N_8801,N_8796);
nor UO_1197 (O_1197,N_9000,N_8221);
nor UO_1198 (O_1198,N_9717,N_8996);
or UO_1199 (O_1199,N_9044,N_9112);
or UO_1200 (O_1200,N_8692,N_8469);
nand UO_1201 (O_1201,N_8259,N_8992);
and UO_1202 (O_1202,N_9194,N_9502);
nand UO_1203 (O_1203,N_9162,N_9905);
nor UO_1204 (O_1204,N_8235,N_8929);
nor UO_1205 (O_1205,N_8884,N_9688);
nand UO_1206 (O_1206,N_9213,N_8537);
nand UO_1207 (O_1207,N_8388,N_8004);
and UO_1208 (O_1208,N_8348,N_8741);
nor UO_1209 (O_1209,N_8037,N_9051);
nor UO_1210 (O_1210,N_9058,N_9021);
nor UO_1211 (O_1211,N_9240,N_9158);
and UO_1212 (O_1212,N_8472,N_8034);
nand UO_1213 (O_1213,N_8737,N_9000);
and UO_1214 (O_1214,N_9844,N_9291);
or UO_1215 (O_1215,N_8269,N_8620);
and UO_1216 (O_1216,N_9333,N_8827);
and UO_1217 (O_1217,N_8732,N_8682);
nand UO_1218 (O_1218,N_9495,N_8438);
nand UO_1219 (O_1219,N_9531,N_9509);
or UO_1220 (O_1220,N_9343,N_8205);
nor UO_1221 (O_1221,N_9540,N_9836);
nor UO_1222 (O_1222,N_9562,N_8891);
nand UO_1223 (O_1223,N_9137,N_9238);
nor UO_1224 (O_1224,N_9064,N_8081);
nor UO_1225 (O_1225,N_8242,N_8505);
nand UO_1226 (O_1226,N_8894,N_9906);
nor UO_1227 (O_1227,N_8895,N_8216);
xnor UO_1228 (O_1228,N_9852,N_8690);
nor UO_1229 (O_1229,N_9573,N_8919);
nand UO_1230 (O_1230,N_9047,N_9835);
nand UO_1231 (O_1231,N_8336,N_9491);
or UO_1232 (O_1232,N_8545,N_9443);
nor UO_1233 (O_1233,N_9182,N_8122);
nor UO_1234 (O_1234,N_9241,N_9277);
nand UO_1235 (O_1235,N_9148,N_8177);
or UO_1236 (O_1236,N_8615,N_9175);
or UO_1237 (O_1237,N_8889,N_9650);
nand UO_1238 (O_1238,N_9589,N_8160);
nand UO_1239 (O_1239,N_9451,N_9037);
nand UO_1240 (O_1240,N_8227,N_8834);
or UO_1241 (O_1241,N_9629,N_9610);
and UO_1242 (O_1242,N_8392,N_9330);
and UO_1243 (O_1243,N_9169,N_9991);
xor UO_1244 (O_1244,N_9127,N_9702);
or UO_1245 (O_1245,N_9707,N_8677);
nand UO_1246 (O_1246,N_8229,N_9560);
nand UO_1247 (O_1247,N_9106,N_8723);
nand UO_1248 (O_1248,N_8072,N_9237);
nand UO_1249 (O_1249,N_9315,N_9872);
nor UO_1250 (O_1250,N_9378,N_9808);
nor UO_1251 (O_1251,N_8454,N_8019);
nand UO_1252 (O_1252,N_9014,N_8162);
nor UO_1253 (O_1253,N_8643,N_8542);
nor UO_1254 (O_1254,N_9588,N_9786);
or UO_1255 (O_1255,N_8015,N_9425);
nor UO_1256 (O_1256,N_9127,N_8026);
or UO_1257 (O_1257,N_9731,N_8818);
nor UO_1258 (O_1258,N_9240,N_9503);
or UO_1259 (O_1259,N_9306,N_8131);
or UO_1260 (O_1260,N_8938,N_8709);
nand UO_1261 (O_1261,N_8007,N_9063);
and UO_1262 (O_1262,N_9843,N_9982);
nor UO_1263 (O_1263,N_9509,N_8315);
and UO_1264 (O_1264,N_9494,N_9655);
or UO_1265 (O_1265,N_8972,N_8410);
nand UO_1266 (O_1266,N_8254,N_9438);
xnor UO_1267 (O_1267,N_8311,N_9153);
and UO_1268 (O_1268,N_8149,N_8342);
nand UO_1269 (O_1269,N_8487,N_8676);
nand UO_1270 (O_1270,N_9965,N_8966);
nor UO_1271 (O_1271,N_9653,N_9993);
or UO_1272 (O_1272,N_9871,N_8999);
nand UO_1273 (O_1273,N_9226,N_9620);
and UO_1274 (O_1274,N_9760,N_9433);
and UO_1275 (O_1275,N_9192,N_9788);
and UO_1276 (O_1276,N_8316,N_8756);
or UO_1277 (O_1277,N_9064,N_8651);
xnor UO_1278 (O_1278,N_9236,N_9733);
or UO_1279 (O_1279,N_9614,N_9792);
nor UO_1280 (O_1280,N_8982,N_9077);
or UO_1281 (O_1281,N_9066,N_9527);
nand UO_1282 (O_1282,N_9485,N_8611);
and UO_1283 (O_1283,N_9392,N_8878);
nor UO_1284 (O_1284,N_8114,N_8860);
nand UO_1285 (O_1285,N_8017,N_8097);
or UO_1286 (O_1286,N_8045,N_8334);
and UO_1287 (O_1287,N_8652,N_9961);
nor UO_1288 (O_1288,N_8398,N_9042);
or UO_1289 (O_1289,N_9374,N_9846);
and UO_1290 (O_1290,N_9292,N_9550);
nor UO_1291 (O_1291,N_8155,N_8971);
nand UO_1292 (O_1292,N_9896,N_8145);
and UO_1293 (O_1293,N_8851,N_8120);
nor UO_1294 (O_1294,N_9628,N_9292);
nor UO_1295 (O_1295,N_9601,N_9870);
nand UO_1296 (O_1296,N_8873,N_9639);
nand UO_1297 (O_1297,N_9026,N_8103);
or UO_1298 (O_1298,N_8646,N_9966);
nor UO_1299 (O_1299,N_8366,N_9382);
nor UO_1300 (O_1300,N_9205,N_9994);
nor UO_1301 (O_1301,N_8557,N_8660);
nand UO_1302 (O_1302,N_9224,N_9637);
nor UO_1303 (O_1303,N_9232,N_8740);
nand UO_1304 (O_1304,N_8354,N_9358);
nand UO_1305 (O_1305,N_8525,N_9445);
or UO_1306 (O_1306,N_8715,N_8231);
or UO_1307 (O_1307,N_8451,N_9011);
and UO_1308 (O_1308,N_8213,N_8289);
nor UO_1309 (O_1309,N_8235,N_9697);
and UO_1310 (O_1310,N_8921,N_8733);
nor UO_1311 (O_1311,N_9868,N_8532);
nor UO_1312 (O_1312,N_8017,N_9433);
nand UO_1313 (O_1313,N_8672,N_9770);
nor UO_1314 (O_1314,N_9363,N_8119);
nor UO_1315 (O_1315,N_9095,N_8146);
or UO_1316 (O_1316,N_8000,N_8360);
and UO_1317 (O_1317,N_8779,N_9187);
nand UO_1318 (O_1318,N_9210,N_8007);
nor UO_1319 (O_1319,N_9617,N_9571);
and UO_1320 (O_1320,N_8526,N_9234);
and UO_1321 (O_1321,N_8839,N_9981);
nor UO_1322 (O_1322,N_9174,N_8599);
nor UO_1323 (O_1323,N_9656,N_9890);
nand UO_1324 (O_1324,N_8801,N_9515);
nand UO_1325 (O_1325,N_8527,N_9401);
nand UO_1326 (O_1326,N_9578,N_8523);
and UO_1327 (O_1327,N_9059,N_8880);
nand UO_1328 (O_1328,N_8868,N_9776);
and UO_1329 (O_1329,N_9311,N_8152);
nor UO_1330 (O_1330,N_9357,N_9438);
and UO_1331 (O_1331,N_9859,N_9293);
nand UO_1332 (O_1332,N_9420,N_9231);
nor UO_1333 (O_1333,N_9389,N_8975);
nor UO_1334 (O_1334,N_8686,N_8335);
or UO_1335 (O_1335,N_8435,N_8919);
nor UO_1336 (O_1336,N_8168,N_9596);
or UO_1337 (O_1337,N_8627,N_9133);
or UO_1338 (O_1338,N_9273,N_8993);
nand UO_1339 (O_1339,N_9176,N_9096);
and UO_1340 (O_1340,N_8766,N_8880);
or UO_1341 (O_1341,N_8369,N_9081);
nor UO_1342 (O_1342,N_9096,N_8318);
or UO_1343 (O_1343,N_9269,N_8021);
and UO_1344 (O_1344,N_8070,N_8740);
and UO_1345 (O_1345,N_9452,N_8174);
or UO_1346 (O_1346,N_8352,N_8206);
and UO_1347 (O_1347,N_9500,N_9474);
nor UO_1348 (O_1348,N_9572,N_8543);
nor UO_1349 (O_1349,N_8774,N_8409);
nor UO_1350 (O_1350,N_8134,N_9094);
and UO_1351 (O_1351,N_8134,N_9039);
and UO_1352 (O_1352,N_8019,N_8477);
or UO_1353 (O_1353,N_8193,N_8201);
xor UO_1354 (O_1354,N_8123,N_9224);
or UO_1355 (O_1355,N_8771,N_8765);
nand UO_1356 (O_1356,N_8739,N_9743);
and UO_1357 (O_1357,N_8382,N_9526);
and UO_1358 (O_1358,N_9115,N_9660);
nand UO_1359 (O_1359,N_8777,N_8841);
nor UO_1360 (O_1360,N_9768,N_8866);
or UO_1361 (O_1361,N_8308,N_8598);
nand UO_1362 (O_1362,N_9053,N_8237);
and UO_1363 (O_1363,N_9535,N_9366);
nand UO_1364 (O_1364,N_8595,N_8027);
and UO_1365 (O_1365,N_9910,N_9510);
nor UO_1366 (O_1366,N_9571,N_9942);
nor UO_1367 (O_1367,N_8131,N_9647);
or UO_1368 (O_1368,N_8791,N_9944);
and UO_1369 (O_1369,N_8212,N_9112);
nor UO_1370 (O_1370,N_8286,N_8457);
nand UO_1371 (O_1371,N_8169,N_8418);
nor UO_1372 (O_1372,N_9115,N_8136);
nand UO_1373 (O_1373,N_8516,N_8750);
nand UO_1374 (O_1374,N_9482,N_8626);
and UO_1375 (O_1375,N_8520,N_9605);
or UO_1376 (O_1376,N_9570,N_9690);
and UO_1377 (O_1377,N_8319,N_8065);
or UO_1378 (O_1378,N_8646,N_8392);
or UO_1379 (O_1379,N_9415,N_8961);
and UO_1380 (O_1380,N_8067,N_9068);
nand UO_1381 (O_1381,N_8795,N_8010);
nor UO_1382 (O_1382,N_9639,N_8401);
or UO_1383 (O_1383,N_8547,N_8816);
and UO_1384 (O_1384,N_8742,N_9239);
or UO_1385 (O_1385,N_9684,N_9108);
or UO_1386 (O_1386,N_8506,N_9936);
nand UO_1387 (O_1387,N_9837,N_9318);
or UO_1388 (O_1388,N_8143,N_9216);
nand UO_1389 (O_1389,N_8469,N_9265);
and UO_1390 (O_1390,N_9937,N_9151);
nor UO_1391 (O_1391,N_8826,N_9446);
or UO_1392 (O_1392,N_9074,N_8501);
or UO_1393 (O_1393,N_8959,N_9949);
and UO_1394 (O_1394,N_9213,N_9508);
xor UO_1395 (O_1395,N_8381,N_9223);
nand UO_1396 (O_1396,N_8227,N_9346);
nor UO_1397 (O_1397,N_9952,N_9876);
or UO_1398 (O_1398,N_9458,N_8733);
nor UO_1399 (O_1399,N_8652,N_9987);
nor UO_1400 (O_1400,N_9037,N_9331);
nor UO_1401 (O_1401,N_8661,N_9986);
nand UO_1402 (O_1402,N_9719,N_9802);
and UO_1403 (O_1403,N_8721,N_8851);
and UO_1404 (O_1404,N_9526,N_9276);
nand UO_1405 (O_1405,N_8246,N_9291);
nand UO_1406 (O_1406,N_9570,N_9723);
xor UO_1407 (O_1407,N_9063,N_8192);
nand UO_1408 (O_1408,N_9611,N_9674);
and UO_1409 (O_1409,N_9623,N_9575);
nand UO_1410 (O_1410,N_8211,N_8539);
nor UO_1411 (O_1411,N_9456,N_8770);
and UO_1412 (O_1412,N_8706,N_8142);
nor UO_1413 (O_1413,N_9619,N_8955);
nand UO_1414 (O_1414,N_9127,N_9063);
xor UO_1415 (O_1415,N_9045,N_9542);
nor UO_1416 (O_1416,N_9927,N_8803);
nand UO_1417 (O_1417,N_8200,N_8150);
nor UO_1418 (O_1418,N_8989,N_9192);
xor UO_1419 (O_1419,N_8341,N_8312);
nor UO_1420 (O_1420,N_9541,N_8487);
and UO_1421 (O_1421,N_9931,N_8230);
or UO_1422 (O_1422,N_8875,N_9677);
xnor UO_1423 (O_1423,N_9585,N_9545);
or UO_1424 (O_1424,N_8998,N_8630);
or UO_1425 (O_1425,N_8792,N_8725);
or UO_1426 (O_1426,N_9979,N_9751);
nor UO_1427 (O_1427,N_9366,N_9259);
nand UO_1428 (O_1428,N_8132,N_9137);
nor UO_1429 (O_1429,N_9411,N_8951);
and UO_1430 (O_1430,N_8319,N_9755);
and UO_1431 (O_1431,N_8603,N_9184);
nand UO_1432 (O_1432,N_9518,N_8629);
and UO_1433 (O_1433,N_9980,N_8527);
nand UO_1434 (O_1434,N_8327,N_8334);
nor UO_1435 (O_1435,N_8585,N_8560);
or UO_1436 (O_1436,N_8179,N_9604);
and UO_1437 (O_1437,N_9992,N_8526);
nor UO_1438 (O_1438,N_9867,N_8974);
nand UO_1439 (O_1439,N_8882,N_8385);
and UO_1440 (O_1440,N_8161,N_8483);
or UO_1441 (O_1441,N_9001,N_9065);
or UO_1442 (O_1442,N_8853,N_8494);
nand UO_1443 (O_1443,N_8635,N_8338);
nand UO_1444 (O_1444,N_8203,N_9064);
or UO_1445 (O_1445,N_9539,N_8135);
and UO_1446 (O_1446,N_9736,N_8077);
and UO_1447 (O_1447,N_8543,N_9137);
and UO_1448 (O_1448,N_9615,N_9578);
and UO_1449 (O_1449,N_8755,N_8620);
or UO_1450 (O_1450,N_9120,N_8538);
and UO_1451 (O_1451,N_9054,N_9704);
nand UO_1452 (O_1452,N_9165,N_8613);
nand UO_1453 (O_1453,N_9612,N_9604);
nand UO_1454 (O_1454,N_8407,N_9238);
nor UO_1455 (O_1455,N_9447,N_9717);
or UO_1456 (O_1456,N_9517,N_9051);
nand UO_1457 (O_1457,N_8645,N_9944);
nand UO_1458 (O_1458,N_8200,N_8720);
or UO_1459 (O_1459,N_8248,N_9437);
and UO_1460 (O_1460,N_9788,N_8737);
nand UO_1461 (O_1461,N_8908,N_8879);
nor UO_1462 (O_1462,N_9410,N_8371);
nor UO_1463 (O_1463,N_8699,N_9593);
nor UO_1464 (O_1464,N_9837,N_8941);
and UO_1465 (O_1465,N_8053,N_9904);
or UO_1466 (O_1466,N_9620,N_9339);
xor UO_1467 (O_1467,N_9412,N_9695);
and UO_1468 (O_1468,N_9545,N_8629);
nand UO_1469 (O_1469,N_9770,N_8957);
nor UO_1470 (O_1470,N_8031,N_9390);
and UO_1471 (O_1471,N_9212,N_9088);
or UO_1472 (O_1472,N_8526,N_9410);
and UO_1473 (O_1473,N_8585,N_9103);
or UO_1474 (O_1474,N_8300,N_8247);
and UO_1475 (O_1475,N_9570,N_8697);
nor UO_1476 (O_1476,N_8098,N_8599);
or UO_1477 (O_1477,N_9353,N_9473);
nor UO_1478 (O_1478,N_9071,N_9719);
nor UO_1479 (O_1479,N_8394,N_8145);
nor UO_1480 (O_1480,N_8913,N_8978);
xnor UO_1481 (O_1481,N_8663,N_9232);
or UO_1482 (O_1482,N_8170,N_8021);
or UO_1483 (O_1483,N_9161,N_8955);
and UO_1484 (O_1484,N_9628,N_9853);
or UO_1485 (O_1485,N_9943,N_9216);
and UO_1486 (O_1486,N_9921,N_8274);
nor UO_1487 (O_1487,N_8441,N_9768);
and UO_1488 (O_1488,N_9820,N_9391);
nand UO_1489 (O_1489,N_8675,N_9633);
nand UO_1490 (O_1490,N_8581,N_8466);
or UO_1491 (O_1491,N_9174,N_9667);
or UO_1492 (O_1492,N_9298,N_8949);
and UO_1493 (O_1493,N_8734,N_8936);
or UO_1494 (O_1494,N_8324,N_8548);
xor UO_1495 (O_1495,N_9293,N_8316);
and UO_1496 (O_1496,N_9399,N_9190);
or UO_1497 (O_1497,N_8598,N_9385);
nand UO_1498 (O_1498,N_9747,N_9288);
nor UO_1499 (O_1499,N_9693,N_8239);
endmodule