module basic_1000_10000_1500_5_levels_2xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
and U0 (N_0,In_718,In_406);
nor U1 (N_1,In_631,In_429);
nor U2 (N_2,In_589,In_601);
or U3 (N_3,In_501,In_832);
nand U4 (N_4,In_155,In_934);
and U5 (N_5,In_957,In_489);
xor U6 (N_6,In_156,In_869);
and U7 (N_7,In_388,In_834);
and U8 (N_8,In_828,In_878);
xnor U9 (N_9,In_982,In_767);
or U10 (N_10,In_320,In_716);
and U11 (N_11,In_915,In_688);
and U12 (N_12,In_374,In_51);
and U13 (N_13,In_268,In_228);
nor U14 (N_14,In_562,In_160);
nor U15 (N_15,In_720,In_644);
nor U16 (N_16,In_573,In_71);
nor U17 (N_17,In_839,In_966);
and U18 (N_18,In_959,In_652);
nand U19 (N_19,In_564,In_849);
and U20 (N_20,In_124,In_276);
and U21 (N_21,In_393,In_129);
nand U22 (N_22,In_905,In_153);
and U23 (N_23,In_559,In_192);
nor U24 (N_24,In_838,In_497);
nor U25 (N_25,In_346,In_963);
nor U26 (N_26,In_74,In_978);
and U27 (N_27,In_146,In_8);
or U28 (N_28,In_969,In_35);
or U29 (N_29,In_45,In_523);
nand U30 (N_30,In_274,In_1);
and U31 (N_31,In_831,In_135);
nor U32 (N_32,In_163,In_603);
or U33 (N_33,In_18,In_223);
nand U34 (N_34,In_841,In_858);
or U35 (N_35,In_951,In_284);
nand U36 (N_36,In_974,In_270);
or U37 (N_37,In_505,In_184);
and U38 (N_38,In_425,In_151);
or U39 (N_39,In_702,In_64);
or U40 (N_40,In_239,In_109);
nand U41 (N_41,In_625,In_507);
or U42 (N_42,In_550,In_14);
and U43 (N_43,In_172,In_113);
and U44 (N_44,In_827,In_461);
nand U45 (N_45,In_5,In_948);
and U46 (N_46,In_924,In_332);
and U47 (N_47,In_793,In_66);
nand U48 (N_48,In_178,In_305);
nor U49 (N_49,In_862,In_536);
xor U50 (N_50,In_30,In_263);
nand U51 (N_51,In_758,In_571);
and U52 (N_52,In_221,In_235);
or U53 (N_53,In_954,In_903);
nor U54 (N_54,In_731,In_668);
nor U55 (N_55,In_300,In_280);
and U56 (N_56,In_619,In_233);
and U57 (N_57,In_732,In_605);
nand U58 (N_58,In_89,In_739);
or U59 (N_59,In_435,In_119);
nor U60 (N_60,In_719,In_889);
or U61 (N_61,In_190,In_80);
nand U62 (N_62,In_787,In_152);
and U63 (N_63,In_532,In_568);
or U64 (N_64,In_514,In_539);
nor U65 (N_65,In_939,In_994);
and U66 (N_66,In_945,In_604);
nor U67 (N_67,In_31,In_96);
or U68 (N_68,In_383,In_750);
or U69 (N_69,In_648,In_385);
or U70 (N_70,In_209,In_250);
xnor U71 (N_71,In_330,In_72);
nand U72 (N_72,In_896,In_317);
and U73 (N_73,In_993,In_456);
and U74 (N_74,In_701,In_174);
nor U75 (N_75,In_195,In_990);
nor U76 (N_76,In_961,In_682);
nor U77 (N_77,In_94,In_421);
nor U78 (N_78,In_240,In_213);
or U79 (N_79,In_43,In_823);
nand U80 (N_80,In_191,In_498);
xor U81 (N_81,In_0,In_721);
nor U82 (N_82,In_970,In_742);
and U83 (N_83,In_985,In_587);
nand U84 (N_84,In_337,In_848);
and U85 (N_85,In_588,In_748);
xnor U86 (N_86,In_917,In_774);
nor U87 (N_87,In_860,In_817);
nand U88 (N_88,In_729,In_251);
and U89 (N_89,In_806,In_710);
nand U90 (N_90,In_473,In_863);
nor U91 (N_91,In_303,In_665);
and U92 (N_92,In_438,In_125);
nand U93 (N_93,In_296,In_302);
nand U94 (N_94,In_369,In_890);
nor U95 (N_95,In_255,In_267);
and U96 (N_96,In_696,In_818);
nand U97 (N_97,In_496,In_667);
or U98 (N_98,In_671,In_411);
nor U99 (N_99,In_492,In_801);
and U100 (N_100,In_947,In_2);
nand U101 (N_101,In_215,In_304);
or U102 (N_102,In_902,In_36);
nor U103 (N_103,In_325,In_189);
nand U104 (N_104,In_976,In_457);
nor U105 (N_105,In_764,In_958);
nand U106 (N_106,In_484,In_164);
nor U107 (N_107,In_104,In_140);
and U108 (N_108,In_364,In_645);
or U109 (N_109,In_37,In_123);
nand U110 (N_110,In_469,In_854);
or U111 (N_111,In_387,In_145);
or U112 (N_112,In_139,In_509);
or U113 (N_113,In_508,In_458);
and U114 (N_114,In_620,In_628);
nor U115 (N_115,In_698,In_711);
and U116 (N_116,In_609,In_158);
nand U117 (N_117,In_499,In_674);
nand U118 (N_118,In_111,In_752);
nor U119 (N_119,In_446,In_621);
nand U120 (N_120,In_363,In_168);
nand U121 (N_121,In_180,In_786);
nand U122 (N_122,In_59,In_700);
nand U123 (N_123,In_776,In_289);
nand U124 (N_124,In_826,In_301);
or U125 (N_125,In_488,In_112);
or U126 (N_126,In_641,In_632);
and U127 (N_127,In_431,In_791);
nor U128 (N_128,In_813,In_697);
and U129 (N_129,In_259,In_326);
nand U130 (N_130,In_805,In_546);
nand U131 (N_131,In_535,In_840);
nand U132 (N_132,In_358,In_271);
and U133 (N_133,In_525,In_84);
and U134 (N_134,In_518,In_802);
nor U135 (N_135,In_12,In_264);
nor U136 (N_136,In_212,In_207);
and U137 (N_137,In_381,In_920);
and U138 (N_138,In_49,In_447);
and U139 (N_139,In_599,In_759);
and U140 (N_140,In_727,In_919);
or U141 (N_141,In_368,In_234);
and U142 (N_142,In_887,In_159);
and U143 (N_143,In_351,In_780);
or U144 (N_144,In_165,In_241);
or U145 (N_145,In_100,In_244);
nand U146 (N_146,In_590,In_20);
nor U147 (N_147,In_136,In_577);
or U148 (N_148,In_283,In_495);
nand U149 (N_149,In_127,In_441);
and U150 (N_150,In_871,In_946);
and U151 (N_151,In_968,In_232);
nand U152 (N_152,In_784,In_686);
nor U153 (N_153,In_114,In_888);
or U154 (N_154,In_713,In_809);
and U155 (N_155,In_730,In_455);
nor U156 (N_156,In_391,In_377);
nand U157 (N_157,In_837,In_524);
or U158 (N_158,In_88,In_214);
nand U159 (N_159,In_194,In_900);
or U160 (N_160,In_371,In_893);
and U161 (N_161,In_208,In_25);
or U162 (N_162,In_442,In_938);
nor U163 (N_163,In_647,In_6);
or U164 (N_164,In_563,In_687);
nor U165 (N_165,In_312,In_61);
nor U166 (N_166,In_650,In_877);
and U167 (N_167,In_996,In_299);
or U168 (N_168,In_973,In_188);
nand U169 (N_169,In_870,In_852);
and U170 (N_170,In_757,In_825);
or U171 (N_171,In_44,In_795);
and U172 (N_172,In_856,In_295);
nor U173 (N_173,In_790,In_851);
nand U174 (N_174,In_204,In_314);
nor U175 (N_175,In_844,In_81);
or U176 (N_176,In_176,In_389);
or U177 (N_177,In_777,In_487);
and U178 (N_178,In_380,In_4);
nand U179 (N_179,In_321,In_660);
nand U180 (N_180,In_740,In_897);
and U181 (N_181,In_278,In_908);
or U182 (N_182,In_79,In_50);
nand U183 (N_183,In_131,In_10);
or U184 (N_184,In_872,In_331);
nor U185 (N_185,In_717,In_964);
or U186 (N_186,In_308,In_940);
or U187 (N_187,In_310,In_15);
or U188 (N_188,In_38,In_699);
and U189 (N_189,In_673,In_803);
and U190 (N_190,In_983,In_999);
nor U191 (N_191,In_646,In_211);
nand U192 (N_192,In_462,In_556);
or U193 (N_193,In_493,In_785);
nand U194 (N_194,In_779,In_46);
or U195 (N_195,In_141,In_63);
and U196 (N_196,In_150,In_747);
or U197 (N_197,In_944,In_282);
nand U198 (N_198,In_980,In_467);
nor U199 (N_199,In_909,In_120);
nand U200 (N_200,In_681,In_770);
and U201 (N_201,In_340,In_744);
or U202 (N_202,In_422,In_899);
and U203 (N_203,In_936,In_875);
or U204 (N_204,In_333,In_677);
and U205 (N_205,In_766,In_728);
nand U206 (N_206,In_291,In_419);
nand U207 (N_207,In_929,In_692);
nand U208 (N_208,In_137,In_39);
nor U209 (N_209,In_988,In_572);
or U210 (N_210,In_933,In_471);
nor U211 (N_211,In_694,In_522);
or U212 (N_212,In_384,In_521);
nand U213 (N_213,In_935,In_110);
and U214 (N_214,In_42,In_685);
or U215 (N_215,In_734,In_943);
and U216 (N_216,In_676,In_480);
nand U217 (N_217,In_147,In_95);
nand U218 (N_218,In_847,In_78);
or U219 (N_219,In_477,In_819);
xor U220 (N_220,In_16,In_275);
nor U221 (N_221,In_29,In_403);
nand U222 (N_222,In_760,In_186);
nand U223 (N_223,In_771,In_753);
nand U224 (N_224,In_27,In_382);
nor U225 (N_225,In_132,In_751);
and U226 (N_226,In_997,In_737);
and U227 (N_227,In_205,In_815);
and U228 (N_228,In_584,In_77);
nor U229 (N_229,In_664,In_836);
nor U230 (N_230,In_3,In_121);
nand U231 (N_231,In_626,In_449);
nor U232 (N_232,In_183,In_638);
and U233 (N_233,In_773,In_754);
nand U234 (N_234,In_460,In_596);
nor U235 (N_235,In_723,In_93);
nand U236 (N_236,In_565,In_65);
nand U237 (N_237,In_470,In_395);
nand U238 (N_238,In_412,In_117);
or U239 (N_239,In_56,In_575);
nand U240 (N_240,In_576,In_262);
nor U241 (N_241,In_354,In_126);
and U242 (N_242,In_356,In_582);
nor U243 (N_243,In_611,In_666);
and U244 (N_244,In_143,In_62);
or U245 (N_245,In_528,In_541);
nand U246 (N_246,In_409,In_13);
and U247 (N_247,In_602,In_649);
and U248 (N_248,In_654,In_334);
or U249 (N_249,In_54,In_433);
and U250 (N_250,In_452,In_502);
and U251 (N_251,In_989,In_622);
nor U252 (N_252,In_83,In_594);
nand U253 (N_253,In_643,In_430);
or U254 (N_254,In_886,In_768);
and U255 (N_255,In_606,In_804);
nand U256 (N_256,In_226,In_87);
nand U257 (N_257,In_181,In_600);
and U258 (N_258,In_468,In_598);
nand U259 (N_259,In_635,In_689);
nand U260 (N_260,In_53,In_722);
or U261 (N_261,In_749,In_23);
and U262 (N_262,In_829,In_329);
and U263 (N_263,In_821,In_118);
nor U264 (N_264,In_311,In_554);
nand U265 (N_265,In_416,In_882);
nand U266 (N_266,In_952,In_70);
nand U267 (N_267,In_634,In_977);
nand U268 (N_268,In_246,In_593);
or U269 (N_269,In_218,In_396);
xor U270 (N_270,In_474,In_558);
xor U271 (N_271,In_7,In_675);
nor U272 (N_272,In_82,In_138);
xor U273 (N_273,In_257,In_971);
and U274 (N_274,In_891,In_914);
or U275 (N_275,In_134,In_128);
xor U276 (N_276,In_342,In_557);
and U277 (N_277,In_322,In_857);
nor U278 (N_278,In_219,In_448);
nor U279 (N_279,In_338,In_597);
nand U280 (N_280,In_916,In_824);
and U281 (N_281,In_617,In_355);
or U282 (N_282,In_911,In_103);
and U283 (N_283,In_451,In_781);
or U284 (N_284,In_91,In_906);
nor U285 (N_285,In_580,In_324);
nand U286 (N_286,In_285,In_515);
and U287 (N_287,In_309,In_569);
and U288 (N_288,In_531,In_177);
nand U289 (N_289,In_979,In_162);
nor U290 (N_290,In_220,In_570);
and U291 (N_291,In_352,In_534);
and U292 (N_292,In_424,In_185);
nor U293 (N_293,In_529,In_423);
or U294 (N_294,In_726,In_895);
and U295 (N_295,In_782,In_414);
or U296 (N_296,In_444,In_294);
and U297 (N_297,In_336,In_765);
nor U298 (N_298,In_868,In_490);
nor U299 (N_299,In_130,In_506);
nor U300 (N_300,In_975,In_17);
and U301 (N_301,In_171,In_341);
nand U302 (N_302,In_199,In_566);
or U303 (N_303,In_439,In_372);
and U304 (N_304,In_864,In_618);
nand U305 (N_305,In_392,In_820);
or U306 (N_306,In_743,In_797);
nand U307 (N_307,In_28,In_405);
nand U308 (N_308,In_273,In_706);
nand U309 (N_309,In_133,In_822);
nor U310 (N_310,In_76,In_453);
or U311 (N_311,In_527,In_608);
xnor U312 (N_312,In_833,In_814);
nand U313 (N_313,In_52,In_472);
nor U314 (N_314,In_479,In_703);
nand U315 (N_315,In_560,In_516);
nor U316 (N_316,In_500,In_401);
or U317 (N_317,In_200,In_735);
and U318 (N_318,In_148,In_835);
and U319 (N_319,In_142,In_553);
nand U320 (N_320,In_206,In_540);
and U321 (N_321,In_68,In_656);
and U322 (N_322,In_761,In_108);
and U323 (N_323,In_861,In_323);
and U324 (N_324,In_879,In_704);
nand U325 (N_325,In_481,In_986);
or U326 (N_326,In_48,In_542);
nand U327 (N_327,In_398,In_610);
and U328 (N_328,In_942,In_99);
nor U329 (N_329,In_658,In_581);
or U330 (N_330,In_261,In_253);
or U331 (N_331,In_607,In_443);
nor U332 (N_332,In_366,In_238);
and U333 (N_333,In_953,In_90);
nand U334 (N_334,In_578,In_695);
nand U335 (N_335,In_921,In_494);
nand U336 (N_336,In_885,In_167);
nand U337 (N_337,In_684,In_519);
nor U338 (N_338,In_436,In_705);
or U339 (N_339,In_427,In_454);
nor U340 (N_340,In_482,In_616);
nor U341 (N_341,In_67,In_633);
and U342 (N_342,In_991,In_231);
nand U343 (N_343,In_657,In_92);
or U344 (N_344,In_402,In_927);
and U345 (N_345,In_778,In_876);
nor U346 (N_346,In_122,In_98);
nor U347 (N_347,In_789,In_34);
or U348 (N_348,In_552,In_538);
or U349 (N_349,In_530,In_808);
and U350 (N_350,In_376,In_483);
or U351 (N_351,In_555,In_440);
nand U352 (N_352,In_286,In_437);
nor U353 (N_353,In_955,In_22);
nand U354 (N_354,In_663,In_816);
and U355 (N_355,In_811,In_995);
or U356 (N_356,In_69,In_865);
or U357 (N_357,In_707,In_335);
nor U358 (N_358,In_901,In_237);
or U359 (N_359,In_75,In_210);
nor U360 (N_360,In_157,In_343);
and U361 (N_361,In_510,In_397);
and U362 (N_362,In_866,In_745);
nor U363 (N_363,In_932,In_659);
nand U364 (N_364,In_894,In_624);
nor U365 (N_365,In_579,In_55);
nor U366 (N_366,In_873,In_24);
or U367 (N_367,In_595,In_170);
and U368 (N_368,In_339,In_923);
nor U369 (N_369,In_230,In_937);
nand U370 (N_370,In_420,In_661);
nor U371 (N_371,In_925,In_281);
or U372 (N_372,In_33,In_217);
nor U373 (N_373,In_222,In_949);
nand U374 (N_374,In_353,In_413);
nand U375 (N_375,In_533,In_842);
nor U376 (N_376,In_630,In_583);
nor U377 (N_377,In_591,In_367);
nand U378 (N_378,In_511,In_344);
nand U379 (N_379,In_883,In_792);
or U380 (N_380,In_623,In_418);
or U381 (N_381,In_960,In_288);
or U382 (N_382,In_105,In_272);
nand U383 (N_383,In_365,In_466);
nor U384 (N_384,In_922,In_57);
nand U385 (N_385,In_850,In_830);
or U386 (N_386,In_724,In_662);
nand U387 (N_387,In_485,In_173);
or U388 (N_388,In_672,In_637);
nand U389 (N_389,In_445,In_166);
nand U390 (N_390,In_491,In_375);
or U391 (N_391,In_812,In_892);
nor U392 (N_392,In_612,In_691);
nand U393 (N_393,In_783,In_898);
and U394 (N_394,In_874,In_772);
nor U395 (N_395,In_260,In_846);
or U396 (N_396,In_984,In_926);
nor U397 (N_397,In_361,In_972);
and U398 (N_398,In_690,In_102);
nor U399 (N_399,In_855,In_867);
and U400 (N_400,In_567,In_357);
nand U401 (N_401,In_520,In_243);
nand U402 (N_402,In_175,In_370);
and U403 (N_403,In_547,In_269);
or U404 (N_404,In_428,In_629);
or U405 (N_405,In_799,In_279);
and U406 (N_406,In_574,In_107);
nor U407 (N_407,In_265,In_586);
nand U408 (N_408,In_715,In_407);
nor U409 (N_409,In_26,In_47);
nand U410 (N_410,In_293,In_202);
or U411 (N_411,In_561,In_229);
and U412 (N_412,In_417,In_627);
nor U413 (N_413,In_544,In_328);
nand U414 (N_414,In_349,In_216);
and U415 (N_415,In_640,In_58);
or U416 (N_416,In_225,In_266);
or U417 (N_417,In_615,In_476);
or U418 (N_418,In_277,In_60);
and U419 (N_419,In_810,In_106);
nor U420 (N_420,In_585,In_306);
nand U421 (N_421,In_297,In_359);
nand U422 (N_422,In_478,In_307);
and U423 (N_423,In_680,In_670);
nor U424 (N_424,In_642,In_543);
or U425 (N_425,In_169,In_348);
and U426 (N_426,In_613,In_636);
nor U427 (N_427,In_517,In_154);
nand U428 (N_428,In_843,In_725);
or U429 (N_429,In_800,In_198);
and U430 (N_430,In_714,In_350);
nand U431 (N_431,In_503,In_224);
nor U432 (N_432,In_762,In_746);
and U433 (N_433,In_179,In_292);
and U434 (N_434,In_85,In_653);
nor U435 (N_435,In_904,In_981);
or U436 (N_436,In_807,In_709);
nor U437 (N_437,In_360,In_242);
xor U438 (N_438,In_32,In_639);
nor U439 (N_439,In_465,In_880);
nor U440 (N_440,In_651,In_537);
or U441 (N_441,In_287,In_551);
nor U442 (N_442,In_21,In_708);
xnor U443 (N_443,In_410,In_526);
or U444 (N_444,In_693,In_245);
nand U445 (N_445,In_40,In_733);
or U446 (N_446,In_434,In_11);
or U447 (N_447,In_415,In_373);
nor U448 (N_448,In_247,In_918);
nor U449 (N_449,In_19,In_512);
or U450 (N_450,In_378,In_97);
nor U451 (N_451,In_679,In_400);
or U452 (N_452,In_404,In_962);
and U453 (N_453,In_738,In_712);
or U454 (N_454,In_101,In_116);
and U455 (N_455,In_881,In_941);
and U456 (N_456,In_203,In_798);
nand U457 (N_457,In_201,In_227);
nor U458 (N_458,In_845,In_796);
xnor U459 (N_459,In_316,In_386);
nand U460 (N_460,In_592,In_930);
or U461 (N_461,In_187,In_678);
or U462 (N_462,In_290,In_9);
nand U463 (N_463,In_86,In_756);
or U464 (N_464,In_144,In_475);
nor U465 (N_465,In_459,In_504);
nand U466 (N_466,In_315,In_258);
nor U467 (N_467,In_965,In_956);
and U468 (N_468,In_998,In_362);
or U469 (N_469,In_193,In_859);
nand U470 (N_470,In_884,In_775);
nand U471 (N_471,In_853,In_683);
nor U472 (N_472,In_41,In_379);
or U473 (N_473,In_408,In_967);
or U474 (N_474,In_992,In_910);
nand U475 (N_475,In_345,In_73);
or U476 (N_476,In_788,In_347);
nand U477 (N_477,In_256,In_254);
and U478 (N_478,In_755,In_115);
or U479 (N_479,In_741,In_432);
and U480 (N_480,In_394,In_669);
and U481 (N_481,In_913,In_196);
nand U482 (N_482,In_236,In_464);
nor U483 (N_483,In_313,In_450);
xnor U484 (N_484,In_987,In_928);
and U485 (N_485,In_252,In_249);
or U486 (N_486,In_794,In_736);
nor U487 (N_487,In_426,In_545);
nand U488 (N_488,In_950,In_298);
nand U489 (N_489,In_318,In_549);
or U490 (N_490,In_614,In_763);
nor U491 (N_491,In_655,In_513);
or U492 (N_492,In_197,In_390);
and U493 (N_493,In_769,In_907);
xnor U494 (N_494,In_931,In_912);
and U495 (N_495,In_399,In_182);
and U496 (N_496,In_161,In_319);
nand U497 (N_497,In_248,In_463);
nor U498 (N_498,In_548,In_486);
or U499 (N_499,In_149,In_327);
or U500 (N_500,In_347,In_263);
nor U501 (N_501,In_612,In_744);
and U502 (N_502,In_0,In_876);
nand U503 (N_503,In_93,In_862);
nor U504 (N_504,In_900,In_368);
nor U505 (N_505,In_603,In_137);
nor U506 (N_506,In_52,In_497);
or U507 (N_507,In_979,In_182);
nand U508 (N_508,In_653,In_532);
nand U509 (N_509,In_558,In_950);
nand U510 (N_510,In_282,In_496);
nand U511 (N_511,In_746,In_13);
and U512 (N_512,In_296,In_478);
xnor U513 (N_513,In_487,In_328);
nand U514 (N_514,In_394,In_117);
and U515 (N_515,In_84,In_108);
or U516 (N_516,In_718,In_823);
or U517 (N_517,In_737,In_529);
nand U518 (N_518,In_591,In_82);
and U519 (N_519,In_489,In_708);
nand U520 (N_520,In_272,In_396);
nor U521 (N_521,In_736,In_399);
and U522 (N_522,In_229,In_143);
or U523 (N_523,In_88,In_142);
or U524 (N_524,In_420,In_807);
nand U525 (N_525,In_606,In_323);
xnor U526 (N_526,In_589,In_915);
or U527 (N_527,In_653,In_835);
nor U528 (N_528,In_750,In_684);
or U529 (N_529,In_882,In_846);
nand U530 (N_530,In_98,In_547);
nor U531 (N_531,In_893,In_706);
nand U532 (N_532,In_929,In_79);
nor U533 (N_533,In_894,In_816);
or U534 (N_534,In_775,In_337);
nand U535 (N_535,In_990,In_495);
nand U536 (N_536,In_933,In_706);
nor U537 (N_537,In_262,In_267);
or U538 (N_538,In_752,In_89);
or U539 (N_539,In_687,In_180);
and U540 (N_540,In_167,In_801);
and U541 (N_541,In_712,In_463);
nor U542 (N_542,In_396,In_582);
xnor U543 (N_543,In_366,In_890);
nand U544 (N_544,In_66,In_527);
nor U545 (N_545,In_451,In_502);
nor U546 (N_546,In_147,In_221);
nor U547 (N_547,In_890,In_213);
or U548 (N_548,In_376,In_364);
and U549 (N_549,In_365,In_661);
and U550 (N_550,In_789,In_932);
or U551 (N_551,In_25,In_577);
and U552 (N_552,In_848,In_500);
nand U553 (N_553,In_176,In_522);
or U554 (N_554,In_549,In_927);
nand U555 (N_555,In_317,In_262);
nor U556 (N_556,In_505,In_579);
nor U557 (N_557,In_339,In_366);
or U558 (N_558,In_331,In_678);
and U559 (N_559,In_794,In_481);
nand U560 (N_560,In_684,In_952);
nand U561 (N_561,In_967,In_456);
or U562 (N_562,In_167,In_75);
nand U563 (N_563,In_732,In_144);
or U564 (N_564,In_257,In_14);
or U565 (N_565,In_147,In_326);
or U566 (N_566,In_582,In_403);
or U567 (N_567,In_119,In_305);
and U568 (N_568,In_648,In_873);
or U569 (N_569,In_194,In_716);
nand U570 (N_570,In_88,In_489);
or U571 (N_571,In_147,In_850);
and U572 (N_572,In_264,In_645);
and U573 (N_573,In_656,In_102);
nor U574 (N_574,In_833,In_51);
nand U575 (N_575,In_354,In_608);
or U576 (N_576,In_79,In_349);
xor U577 (N_577,In_984,In_642);
and U578 (N_578,In_27,In_132);
or U579 (N_579,In_638,In_571);
and U580 (N_580,In_877,In_838);
and U581 (N_581,In_772,In_900);
nand U582 (N_582,In_950,In_925);
nor U583 (N_583,In_64,In_935);
nand U584 (N_584,In_958,In_835);
or U585 (N_585,In_945,In_650);
and U586 (N_586,In_553,In_385);
or U587 (N_587,In_462,In_460);
nand U588 (N_588,In_511,In_482);
or U589 (N_589,In_223,In_505);
and U590 (N_590,In_222,In_395);
nand U591 (N_591,In_735,In_577);
nand U592 (N_592,In_577,In_994);
nand U593 (N_593,In_867,In_826);
or U594 (N_594,In_447,In_255);
or U595 (N_595,In_567,In_70);
and U596 (N_596,In_496,In_234);
nor U597 (N_597,In_857,In_274);
nand U598 (N_598,In_258,In_205);
or U599 (N_599,In_833,In_655);
and U600 (N_600,In_623,In_852);
or U601 (N_601,In_912,In_343);
and U602 (N_602,In_726,In_900);
nor U603 (N_603,In_37,In_532);
and U604 (N_604,In_252,In_899);
nand U605 (N_605,In_762,In_77);
or U606 (N_606,In_460,In_606);
xnor U607 (N_607,In_768,In_568);
nand U608 (N_608,In_580,In_476);
nand U609 (N_609,In_13,In_385);
and U610 (N_610,In_759,In_330);
or U611 (N_611,In_542,In_184);
nand U612 (N_612,In_31,In_625);
or U613 (N_613,In_895,In_484);
and U614 (N_614,In_822,In_732);
or U615 (N_615,In_916,In_21);
and U616 (N_616,In_435,In_152);
nand U617 (N_617,In_67,In_915);
and U618 (N_618,In_49,In_194);
nand U619 (N_619,In_865,In_941);
nand U620 (N_620,In_307,In_614);
or U621 (N_621,In_570,In_392);
nor U622 (N_622,In_457,In_342);
nor U623 (N_623,In_767,In_180);
or U624 (N_624,In_33,In_748);
nor U625 (N_625,In_676,In_838);
nand U626 (N_626,In_585,In_530);
nor U627 (N_627,In_333,In_983);
nor U628 (N_628,In_219,In_570);
nor U629 (N_629,In_724,In_411);
or U630 (N_630,In_674,In_885);
or U631 (N_631,In_766,In_979);
or U632 (N_632,In_97,In_688);
nor U633 (N_633,In_624,In_626);
nand U634 (N_634,In_500,In_223);
and U635 (N_635,In_950,In_507);
or U636 (N_636,In_405,In_38);
nor U637 (N_637,In_204,In_535);
or U638 (N_638,In_203,In_106);
nand U639 (N_639,In_327,In_260);
and U640 (N_640,In_157,In_453);
nor U641 (N_641,In_445,In_982);
nor U642 (N_642,In_950,In_524);
nand U643 (N_643,In_353,In_827);
nor U644 (N_644,In_291,In_394);
nand U645 (N_645,In_680,In_26);
and U646 (N_646,In_823,In_635);
and U647 (N_647,In_333,In_15);
xor U648 (N_648,In_152,In_780);
nand U649 (N_649,In_136,In_696);
nand U650 (N_650,In_554,In_166);
nand U651 (N_651,In_700,In_242);
and U652 (N_652,In_688,In_875);
and U653 (N_653,In_984,In_204);
nor U654 (N_654,In_3,In_91);
and U655 (N_655,In_465,In_944);
nor U656 (N_656,In_938,In_374);
or U657 (N_657,In_768,In_552);
or U658 (N_658,In_615,In_998);
or U659 (N_659,In_161,In_365);
nand U660 (N_660,In_32,In_141);
and U661 (N_661,In_494,In_470);
or U662 (N_662,In_0,In_4);
nand U663 (N_663,In_728,In_773);
or U664 (N_664,In_102,In_777);
nor U665 (N_665,In_613,In_128);
and U666 (N_666,In_821,In_160);
and U667 (N_667,In_67,In_850);
or U668 (N_668,In_716,In_708);
and U669 (N_669,In_44,In_502);
or U670 (N_670,In_543,In_178);
and U671 (N_671,In_484,In_277);
nor U672 (N_672,In_803,In_576);
and U673 (N_673,In_694,In_259);
or U674 (N_674,In_627,In_890);
and U675 (N_675,In_421,In_296);
nand U676 (N_676,In_767,In_316);
or U677 (N_677,In_580,In_191);
nand U678 (N_678,In_603,In_631);
or U679 (N_679,In_725,In_830);
xnor U680 (N_680,In_560,In_95);
nand U681 (N_681,In_606,In_128);
nand U682 (N_682,In_37,In_624);
nor U683 (N_683,In_708,In_710);
nand U684 (N_684,In_863,In_409);
or U685 (N_685,In_958,In_137);
nor U686 (N_686,In_344,In_605);
or U687 (N_687,In_440,In_636);
and U688 (N_688,In_263,In_780);
and U689 (N_689,In_47,In_29);
or U690 (N_690,In_838,In_589);
or U691 (N_691,In_551,In_478);
nand U692 (N_692,In_731,In_765);
and U693 (N_693,In_357,In_765);
nor U694 (N_694,In_836,In_195);
xnor U695 (N_695,In_915,In_698);
nand U696 (N_696,In_656,In_720);
or U697 (N_697,In_61,In_250);
nand U698 (N_698,In_913,In_651);
nand U699 (N_699,In_658,In_105);
and U700 (N_700,In_986,In_762);
or U701 (N_701,In_258,In_128);
and U702 (N_702,In_639,In_669);
nand U703 (N_703,In_652,In_553);
and U704 (N_704,In_785,In_968);
or U705 (N_705,In_232,In_648);
or U706 (N_706,In_708,In_678);
nor U707 (N_707,In_280,In_682);
or U708 (N_708,In_126,In_831);
xnor U709 (N_709,In_48,In_989);
and U710 (N_710,In_195,In_919);
and U711 (N_711,In_168,In_186);
and U712 (N_712,In_336,In_460);
nand U713 (N_713,In_360,In_621);
or U714 (N_714,In_186,In_701);
and U715 (N_715,In_472,In_975);
or U716 (N_716,In_82,In_440);
nor U717 (N_717,In_876,In_435);
or U718 (N_718,In_382,In_3);
and U719 (N_719,In_874,In_771);
nand U720 (N_720,In_466,In_914);
and U721 (N_721,In_161,In_104);
and U722 (N_722,In_757,In_836);
nor U723 (N_723,In_380,In_412);
nor U724 (N_724,In_863,In_893);
nor U725 (N_725,In_888,In_167);
or U726 (N_726,In_388,In_612);
nor U727 (N_727,In_382,In_152);
xnor U728 (N_728,In_398,In_642);
nand U729 (N_729,In_908,In_443);
or U730 (N_730,In_95,In_256);
or U731 (N_731,In_980,In_833);
or U732 (N_732,In_938,In_724);
or U733 (N_733,In_123,In_866);
or U734 (N_734,In_36,In_222);
nand U735 (N_735,In_803,In_499);
or U736 (N_736,In_457,In_606);
and U737 (N_737,In_62,In_909);
nor U738 (N_738,In_195,In_570);
nand U739 (N_739,In_818,In_694);
or U740 (N_740,In_387,In_521);
nand U741 (N_741,In_367,In_424);
nor U742 (N_742,In_208,In_155);
or U743 (N_743,In_201,In_432);
and U744 (N_744,In_323,In_869);
or U745 (N_745,In_683,In_553);
nand U746 (N_746,In_313,In_264);
and U747 (N_747,In_61,In_684);
and U748 (N_748,In_718,In_190);
nor U749 (N_749,In_763,In_708);
or U750 (N_750,In_247,In_22);
and U751 (N_751,In_761,In_522);
nor U752 (N_752,In_77,In_151);
nor U753 (N_753,In_596,In_206);
or U754 (N_754,In_693,In_279);
nand U755 (N_755,In_385,In_484);
or U756 (N_756,In_697,In_12);
or U757 (N_757,In_300,In_441);
and U758 (N_758,In_759,In_960);
and U759 (N_759,In_237,In_999);
nor U760 (N_760,In_708,In_912);
nor U761 (N_761,In_416,In_202);
nand U762 (N_762,In_712,In_861);
nor U763 (N_763,In_45,In_662);
nor U764 (N_764,In_508,In_284);
or U765 (N_765,In_799,In_364);
nor U766 (N_766,In_133,In_640);
or U767 (N_767,In_162,In_471);
nor U768 (N_768,In_565,In_916);
nand U769 (N_769,In_276,In_193);
and U770 (N_770,In_603,In_933);
nand U771 (N_771,In_346,In_837);
nand U772 (N_772,In_74,In_240);
nand U773 (N_773,In_951,In_786);
nor U774 (N_774,In_284,In_272);
nand U775 (N_775,In_387,In_194);
nor U776 (N_776,In_159,In_39);
nor U777 (N_777,In_891,In_533);
or U778 (N_778,In_973,In_592);
nor U779 (N_779,In_750,In_324);
xor U780 (N_780,In_857,In_487);
nand U781 (N_781,In_617,In_652);
nor U782 (N_782,In_230,In_392);
or U783 (N_783,In_460,In_117);
nor U784 (N_784,In_291,In_335);
or U785 (N_785,In_815,In_436);
and U786 (N_786,In_281,In_234);
nor U787 (N_787,In_842,In_681);
nor U788 (N_788,In_631,In_497);
nor U789 (N_789,In_212,In_913);
nor U790 (N_790,In_277,In_564);
nor U791 (N_791,In_971,In_665);
or U792 (N_792,In_228,In_488);
nor U793 (N_793,In_738,In_521);
nand U794 (N_794,In_617,In_119);
or U795 (N_795,In_702,In_710);
or U796 (N_796,In_461,In_245);
and U797 (N_797,In_243,In_325);
nor U798 (N_798,In_153,In_275);
and U799 (N_799,In_94,In_555);
nand U800 (N_800,In_125,In_734);
nand U801 (N_801,In_320,In_621);
nor U802 (N_802,In_669,In_863);
or U803 (N_803,In_697,In_565);
or U804 (N_804,In_831,In_616);
nand U805 (N_805,In_105,In_241);
nand U806 (N_806,In_479,In_295);
nand U807 (N_807,In_557,In_895);
or U808 (N_808,In_566,In_912);
nor U809 (N_809,In_688,In_55);
or U810 (N_810,In_125,In_241);
nor U811 (N_811,In_868,In_471);
or U812 (N_812,In_601,In_738);
or U813 (N_813,In_656,In_85);
and U814 (N_814,In_534,In_773);
nand U815 (N_815,In_608,In_241);
nor U816 (N_816,In_997,In_230);
or U817 (N_817,In_948,In_789);
xnor U818 (N_818,In_373,In_739);
nand U819 (N_819,In_576,In_870);
and U820 (N_820,In_34,In_795);
nor U821 (N_821,In_889,In_863);
and U822 (N_822,In_733,In_667);
and U823 (N_823,In_294,In_875);
nor U824 (N_824,In_371,In_229);
nor U825 (N_825,In_69,In_933);
and U826 (N_826,In_861,In_910);
or U827 (N_827,In_920,In_603);
nand U828 (N_828,In_660,In_588);
or U829 (N_829,In_186,In_331);
or U830 (N_830,In_776,In_678);
and U831 (N_831,In_837,In_468);
nor U832 (N_832,In_303,In_166);
nor U833 (N_833,In_81,In_420);
nor U834 (N_834,In_160,In_778);
nor U835 (N_835,In_974,In_924);
and U836 (N_836,In_596,In_878);
or U837 (N_837,In_26,In_746);
and U838 (N_838,In_115,In_370);
or U839 (N_839,In_813,In_162);
and U840 (N_840,In_671,In_686);
nor U841 (N_841,In_822,In_83);
and U842 (N_842,In_751,In_180);
nand U843 (N_843,In_146,In_676);
or U844 (N_844,In_588,In_968);
or U845 (N_845,In_153,In_222);
or U846 (N_846,In_778,In_591);
or U847 (N_847,In_768,In_421);
nor U848 (N_848,In_387,In_662);
nand U849 (N_849,In_168,In_53);
nor U850 (N_850,In_329,In_765);
and U851 (N_851,In_357,In_71);
nand U852 (N_852,In_459,In_438);
nor U853 (N_853,In_484,In_252);
and U854 (N_854,In_161,In_456);
and U855 (N_855,In_518,In_741);
and U856 (N_856,In_811,In_649);
nor U857 (N_857,In_537,In_347);
xnor U858 (N_858,In_739,In_925);
and U859 (N_859,In_733,In_437);
nor U860 (N_860,In_791,In_998);
and U861 (N_861,In_336,In_67);
or U862 (N_862,In_494,In_68);
nor U863 (N_863,In_172,In_122);
or U864 (N_864,In_416,In_989);
nand U865 (N_865,In_916,In_696);
or U866 (N_866,In_796,In_26);
xor U867 (N_867,In_651,In_26);
or U868 (N_868,In_885,In_662);
nor U869 (N_869,In_722,In_367);
or U870 (N_870,In_501,In_18);
and U871 (N_871,In_129,In_478);
nor U872 (N_872,In_91,In_494);
or U873 (N_873,In_181,In_67);
or U874 (N_874,In_128,In_13);
or U875 (N_875,In_826,In_921);
nand U876 (N_876,In_273,In_557);
or U877 (N_877,In_374,In_334);
and U878 (N_878,In_791,In_13);
or U879 (N_879,In_798,In_576);
nand U880 (N_880,In_872,In_362);
or U881 (N_881,In_996,In_954);
nor U882 (N_882,In_188,In_980);
nor U883 (N_883,In_393,In_81);
nor U884 (N_884,In_280,In_618);
nand U885 (N_885,In_521,In_374);
nor U886 (N_886,In_161,In_11);
and U887 (N_887,In_606,In_126);
nand U888 (N_888,In_248,In_845);
nand U889 (N_889,In_100,In_260);
and U890 (N_890,In_133,In_13);
and U891 (N_891,In_833,In_82);
nand U892 (N_892,In_776,In_916);
and U893 (N_893,In_702,In_36);
nand U894 (N_894,In_893,In_622);
nor U895 (N_895,In_671,In_648);
and U896 (N_896,In_944,In_994);
nand U897 (N_897,In_609,In_98);
nor U898 (N_898,In_411,In_203);
nand U899 (N_899,In_136,In_331);
nor U900 (N_900,In_572,In_247);
nor U901 (N_901,In_893,In_542);
nand U902 (N_902,In_464,In_73);
and U903 (N_903,In_628,In_486);
and U904 (N_904,In_290,In_285);
or U905 (N_905,In_291,In_176);
nand U906 (N_906,In_778,In_25);
nor U907 (N_907,In_590,In_909);
nor U908 (N_908,In_764,In_331);
and U909 (N_909,In_729,In_875);
nor U910 (N_910,In_614,In_653);
nor U911 (N_911,In_941,In_393);
nor U912 (N_912,In_182,In_334);
nor U913 (N_913,In_427,In_351);
nand U914 (N_914,In_740,In_401);
nor U915 (N_915,In_355,In_498);
and U916 (N_916,In_380,In_372);
and U917 (N_917,In_355,In_545);
or U918 (N_918,In_982,In_552);
or U919 (N_919,In_365,In_504);
or U920 (N_920,In_276,In_540);
nor U921 (N_921,In_611,In_535);
or U922 (N_922,In_366,In_537);
nand U923 (N_923,In_573,In_612);
nor U924 (N_924,In_57,In_319);
nor U925 (N_925,In_699,In_563);
or U926 (N_926,In_659,In_100);
nor U927 (N_927,In_929,In_396);
and U928 (N_928,In_652,In_576);
nand U929 (N_929,In_540,In_513);
or U930 (N_930,In_415,In_887);
nand U931 (N_931,In_769,In_742);
or U932 (N_932,In_858,In_735);
or U933 (N_933,In_209,In_798);
or U934 (N_934,In_424,In_394);
nor U935 (N_935,In_899,In_869);
xor U936 (N_936,In_625,In_833);
or U937 (N_937,In_255,In_790);
or U938 (N_938,In_325,In_493);
nor U939 (N_939,In_467,In_750);
nor U940 (N_940,In_306,In_741);
or U941 (N_941,In_279,In_717);
nand U942 (N_942,In_831,In_667);
nor U943 (N_943,In_562,In_774);
or U944 (N_944,In_79,In_762);
nor U945 (N_945,In_398,In_439);
nor U946 (N_946,In_203,In_566);
and U947 (N_947,In_65,In_593);
and U948 (N_948,In_454,In_58);
and U949 (N_949,In_657,In_285);
nor U950 (N_950,In_821,In_341);
and U951 (N_951,In_928,In_786);
or U952 (N_952,In_335,In_149);
or U953 (N_953,In_775,In_640);
nand U954 (N_954,In_134,In_514);
nand U955 (N_955,In_112,In_983);
and U956 (N_956,In_125,In_692);
and U957 (N_957,In_675,In_691);
or U958 (N_958,In_841,In_512);
or U959 (N_959,In_95,In_393);
nor U960 (N_960,In_530,In_415);
or U961 (N_961,In_563,In_959);
and U962 (N_962,In_197,In_43);
nand U963 (N_963,In_79,In_846);
or U964 (N_964,In_924,In_748);
and U965 (N_965,In_172,In_559);
nand U966 (N_966,In_156,In_902);
and U967 (N_967,In_675,In_303);
nand U968 (N_968,In_584,In_180);
nand U969 (N_969,In_95,In_523);
and U970 (N_970,In_693,In_902);
nand U971 (N_971,In_974,In_641);
nand U972 (N_972,In_761,In_766);
nand U973 (N_973,In_205,In_576);
or U974 (N_974,In_369,In_485);
or U975 (N_975,In_316,In_650);
nand U976 (N_976,In_592,In_170);
nor U977 (N_977,In_508,In_391);
and U978 (N_978,In_646,In_486);
and U979 (N_979,In_534,In_658);
nor U980 (N_980,In_848,In_597);
or U981 (N_981,In_82,In_883);
nor U982 (N_982,In_176,In_444);
and U983 (N_983,In_913,In_51);
or U984 (N_984,In_573,In_874);
nand U985 (N_985,In_882,In_2);
and U986 (N_986,In_260,In_597);
nor U987 (N_987,In_407,In_616);
nor U988 (N_988,In_25,In_57);
and U989 (N_989,In_986,In_584);
or U990 (N_990,In_43,In_786);
nor U991 (N_991,In_929,In_981);
and U992 (N_992,In_628,In_789);
nand U993 (N_993,In_455,In_29);
nor U994 (N_994,In_501,In_901);
nand U995 (N_995,In_950,In_872);
nand U996 (N_996,In_910,In_518);
nand U997 (N_997,In_531,In_957);
nand U998 (N_998,In_82,In_139);
nor U999 (N_999,In_106,In_993);
nor U1000 (N_1000,In_320,In_189);
nand U1001 (N_1001,In_771,In_865);
and U1002 (N_1002,In_370,In_444);
nand U1003 (N_1003,In_174,In_548);
nand U1004 (N_1004,In_327,In_500);
and U1005 (N_1005,In_599,In_122);
nand U1006 (N_1006,In_535,In_455);
nor U1007 (N_1007,In_233,In_653);
nand U1008 (N_1008,In_640,In_980);
or U1009 (N_1009,In_692,In_724);
nand U1010 (N_1010,In_368,In_528);
and U1011 (N_1011,In_590,In_781);
nand U1012 (N_1012,In_82,In_121);
nand U1013 (N_1013,In_130,In_583);
and U1014 (N_1014,In_708,In_714);
nand U1015 (N_1015,In_139,In_126);
nand U1016 (N_1016,In_885,In_416);
nor U1017 (N_1017,In_590,In_886);
and U1018 (N_1018,In_970,In_889);
nor U1019 (N_1019,In_325,In_486);
nor U1020 (N_1020,In_676,In_406);
nor U1021 (N_1021,In_406,In_886);
and U1022 (N_1022,In_927,In_97);
nand U1023 (N_1023,In_252,In_758);
xnor U1024 (N_1024,In_813,In_272);
nand U1025 (N_1025,In_498,In_5);
or U1026 (N_1026,In_835,In_896);
and U1027 (N_1027,In_593,In_91);
nor U1028 (N_1028,In_80,In_532);
xnor U1029 (N_1029,In_837,In_428);
and U1030 (N_1030,In_991,In_962);
or U1031 (N_1031,In_602,In_860);
nand U1032 (N_1032,In_8,In_703);
nor U1033 (N_1033,In_135,In_397);
nor U1034 (N_1034,In_340,In_586);
or U1035 (N_1035,In_157,In_323);
nor U1036 (N_1036,In_331,In_394);
and U1037 (N_1037,In_996,In_900);
nand U1038 (N_1038,In_99,In_515);
nand U1039 (N_1039,In_103,In_206);
or U1040 (N_1040,In_794,In_926);
and U1041 (N_1041,In_717,In_14);
nand U1042 (N_1042,In_592,In_848);
nor U1043 (N_1043,In_183,In_285);
or U1044 (N_1044,In_676,In_304);
nor U1045 (N_1045,In_812,In_839);
and U1046 (N_1046,In_486,In_409);
nor U1047 (N_1047,In_562,In_868);
nor U1048 (N_1048,In_397,In_11);
or U1049 (N_1049,In_331,In_20);
nor U1050 (N_1050,In_359,In_747);
nand U1051 (N_1051,In_496,In_685);
nor U1052 (N_1052,In_88,In_715);
xnor U1053 (N_1053,In_1,In_136);
or U1054 (N_1054,In_872,In_429);
nand U1055 (N_1055,In_816,In_1);
nor U1056 (N_1056,In_231,In_204);
or U1057 (N_1057,In_82,In_799);
or U1058 (N_1058,In_793,In_246);
nand U1059 (N_1059,In_210,In_499);
or U1060 (N_1060,In_24,In_306);
nor U1061 (N_1061,In_650,In_337);
and U1062 (N_1062,In_792,In_706);
and U1063 (N_1063,In_361,In_793);
and U1064 (N_1064,In_292,In_339);
and U1065 (N_1065,In_977,In_34);
or U1066 (N_1066,In_43,In_769);
and U1067 (N_1067,In_990,In_666);
nand U1068 (N_1068,In_785,In_784);
or U1069 (N_1069,In_555,In_335);
and U1070 (N_1070,In_654,In_756);
or U1071 (N_1071,In_681,In_446);
nand U1072 (N_1072,In_922,In_600);
nand U1073 (N_1073,In_16,In_887);
xor U1074 (N_1074,In_66,In_284);
nand U1075 (N_1075,In_67,In_76);
and U1076 (N_1076,In_400,In_283);
or U1077 (N_1077,In_245,In_622);
or U1078 (N_1078,In_399,In_433);
xnor U1079 (N_1079,In_902,In_850);
nand U1080 (N_1080,In_78,In_687);
or U1081 (N_1081,In_586,In_814);
nor U1082 (N_1082,In_671,In_816);
or U1083 (N_1083,In_482,In_821);
xnor U1084 (N_1084,In_240,In_658);
or U1085 (N_1085,In_580,In_780);
or U1086 (N_1086,In_564,In_589);
nand U1087 (N_1087,In_480,In_226);
or U1088 (N_1088,In_265,In_651);
nor U1089 (N_1089,In_435,In_763);
nand U1090 (N_1090,In_286,In_891);
and U1091 (N_1091,In_589,In_922);
nand U1092 (N_1092,In_646,In_112);
or U1093 (N_1093,In_562,In_60);
or U1094 (N_1094,In_297,In_598);
or U1095 (N_1095,In_757,In_962);
nor U1096 (N_1096,In_207,In_649);
nor U1097 (N_1097,In_533,In_594);
and U1098 (N_1098,In_436,In_471);
or U1099 (N_1099,In_656,In_185);
or U1100 (N_1100,In_646,In_738);
nor U1101 (N_1101,In_89,In_5);
and U1102 (N_1102,In_131,In_99);
or U1103 (N_1103,In_632,In_574);
nor U1104 (N_1104,In_524,In_913);
nand U1105 (N_1105,In_926,In_194);
or U1106 (N_1106,In_518,In_885);
nand U1107 (N_1107,In_716,In_758);
and U1108 (N_1108,In_815,In_663);
or U1109 (N_1109,In_964,In_736);
and U1110 (N_1110,In_585,In_947);
or U1111 (N_1111,In_84,In_588);
nand U1112 (N_1112,In_3,In_751);
nor U1113 (N_1113,In_392,In_667);
nor U1114 (N_1114,In_833,In_911);
nand U1115 (N_1115,In_817,In_875);
nand U1116 (N_1116,In_477,In_971);
and U1117 (N_1117,In_5,In_651);
nand U1118 (N_1118,In_681,In_658);
and U1119 (N_1119,In_644,In_617);
or U1120 (N_1120,In_48,In_621);
or U1121 (N_1121,In_804,In_754);
and U1122 (N_1122,In_26,In_955);
nor U1123 (N_1123,In_658,In_325);
nand U1124 (N_1124,In_754,In_495);
or U1125 (N_1125,In_123,In_401);
and U1126 (N_1126,In_190,In_929);
or U1127 (N_1127,In_639,In_587);
and U1128 (N_1128,In_976,In_105);
nor U1129 (N_1129,In_705,In_519);
nor U1130 (N_1130,In_189,In_956);
or U1131 (N_1131,In_969,In_186);
and U1132 (N_1132,In_160,In_672);
or U1133 (N_1133,In_561,In_503);
nor U1134 (N_1134,In_885,In_833);
or U1135 (N_1135,In_288,In_9);
or U1136 (N_1136,In_769,In_570);
nand U1137 (N_1137,In_639,In_348);
nor U1138 (N_1138,In_142,In_699);
and U1139 (N_1139,In_796,In_799);
nand U1140 (N_1140,In_984,In_812);
nor U1141 (N_1141,In_876,In_546);
nor U1142 (N_1142,In_929,In_661);
and U1143 (N_1143,In_777,In_681);
nor U1144 (N_1144,In_493,In_646);
or U1145 (N_1145,In_335,In_282);
or U1146 (N_1146,In_162,In_108);
or U1147 (N_1147,In_589,In_673);
and U1148 (N_1148,In_481,In_982);
or U1149 (N_1149,In_703,In_609);
nand U1150 (N_1150,In_485,In_650);
nor U1151 (N_1151,In_970,In_276);
nand U1152 (N_1152,In_637,In_934);
nor U1153 (N_1153,In_707,In_581);
nor U1154 (N_1154,In_20,In_235);
or U1155 (N_1155,In_719,In_78);
and U1156 (N_1156,In_416,In_144);
nor U1157 (N_1157,In_442,In_317);
nor U1158 (N_1158,In_362,In_355);
and U1159 (N_1159,In_489,In_160);
or U1160 (N_1160,In_746,In_404);
nand U1161 (N_1161,In_229,In_699);
xnor U1162 (N_1162,In_267,In_963);
nand U1163 (N_1163,In_645,In_436);
nor U1164 (N_1164,In_446,In_5);
nor U1165 (N_1165,In_397,In_64);
xor U1166 (N_1166,In_47,In_318);
and U1167 (N_1167,In_450,In_387);
or U1168 (N_1168,In_403,In_543);
or U1169 (N_1169,In_620,In_982);
nand U1170 (N_1170,In_596,In_298);
or U1171 (N_1171,In_60,In_464);
nand U1172 (N_1172,In_803,In_807);
or U1173 (N_1173,In_233,In_325);
nor U1174 (N_1174,In_737,In_15);
nor U1175 (N_1175,In_175,In_252);
nor U1176 (N_1176,In_31,In_5);
or U1177 (N_1177,In_731,In_873);
nor U1178 (N_1178,In_36,In_143);
nor U1179 (N_1179,In_632,In_968);
nand U1180 (N_1180,In_970,In_228);
or U1181 (N_1181,In_140,In_837);
nand U1182 (N_1182,In_746,In_391);
nor U1183 (N_1183,In_509,In_807);
and U1184 (N_1184,In_123,In_61);
nor U1185 (N_1185,In_599,In_450);
nor U1186 (N_1186,In_229,In_350);
or U1187 (N_1187,In_81,In_957);
or U1188 (N_1188,In_92,In_118);
nand U1189 (N_1189,In_457,In_321);
and U1190 (N_1190,In_489,In_165);
or U1191 (N_1191,In_630,In_50);
and U1192 (N_1192,In_432,In_673);
nor U1193 (N_1193,In_394,In_450);
and U1194 (N_1194,In_258,In_642);
or U1195 (N_1195,In_508,In_699);
nand U1196 (N_1196,In_8,In_759);
and U1197 (N_1197,In_968,In_841);
nor U1198 (N_1198,In_310,In_787);
or U1199 (N_1199,In_348,In_645);
nor U1200 (N_1200,In_328,In_269);
or U1201 (N_1201,In_283,In_321);
nor U1202 (N_1202,In_994,In_146);
or U1203 (N_1203,In_381,In_377);
nor U1204 (N_1204,In_286,In_195);
or U1205 (N_1205,In_114,In_614);
nand U1206 (N_1206,In_495,In_685);
nand U1207 (N_1207,In_904,In_709);
and U1208 (N_1208,In_412,In_548);
and U1209 (N_1209,In_230,In_673);
xor U1210 (N_1210,In_189,In_220);
or U1211 (N_1211,In_761,In_360);
nor U1212 (N_1212,In_624,In_377);
nor U1213 (N_1213,In_106,In_854);
or U1214 (N_1214,In_650,In_866);
nand U1215 (N_1215,In_733,In_873);
or U1216 (N_1216,In_615,In_370);
nand U1217 (N_1217,In_887,In_47);
nand U1218 (N_1218,In_75,In_74);
xor U1219 (N_1219,In_161,In_462);
and U1220 (N_1220,In_873,In_764);
or U1221 (N_1221,In_644,In_562);
nand U1222 (N_1222,In_110,In_0);
nor U1223 (N_1223,In_225,In_104);
and U1224 (N_1224,In_788,In_794);
or U1225 (N_1225,In_787,In_209);
nor U1226 (N_1226,In_117,In_878);
and U1227 (N_1227,In_165,In_118);
nor U1228 (N_1228,In_359,In_912);
nor U1229 (N_1229,In_371,In_823);
and U1230 (N_1230,In_473,In_390);
nand U1231 (N_1231,In_945,In_619);
nor U1232 (N_1232,In_471,In_513);
nand U1233 (N_1233,In_968,In_746);
and U1234 (N_1234,In_774,In_951);
nand U1235 (N_1235,In_949,In_527);
nand U1236 (N_1236,In_572,In_648);
nor U1237 (N_1237,In_280,In_289);
or U1238 (N_1238,In_533,In_148);
nor U1239 (N_1239,In_770,In_808);
nand U1240 (N_1240,In_847,In_307);
xor U1241 (N_1241,In_203,In_357);
and U1242 (N_1242,In_821,In_462);
nand U1243 (N_1243,In_763,In_342);
nand U1244 (N_1244,In_340,In_99);
nor U1245 (N_1245,In_727,In_284);
nor U1246 (N_1246,In_462,In_268);
nor U1247 (N_1247,In_356,In_585);
or U1248 (N_1248,In_864,In_383);
or U1249 (N_1249,In_95,In_37);
nand U1250 (N_1250,In_337,In_397);
and U1251 (N_1251,In_23,In_773);
nand U1252 (N_1252,In_270,In_945);
xnor U1253 (N_1253,In_883,In_562);
nor U1254 (N_1254,In_948,In_366);
or U1255 (N_1255,In_340,In_13);
and U1256 (N_1256,In_316,In_476);
nand U1257 (N_1257,In_900,In_901);
nor U1258 (N_1258,In_341,In_164);
nand U1259 (N_1259,In_619,In_405);
and U1260 (N_1260,In_654,In_139);
or U1261 (N_1261,In_277,In_783);
nand U1262 (N_1262,In_376,In_565);
and U1263 (N_1263,In_707,In_430);
or U1264 (N_1264,In_116,In_58);
or U1265 (N_1265,In_136,In_945);
nand U1266 (N_1266,In_797,In_823);
or U1267 (N_1267,In_707,In_76);
nor U1268 (N_1268,In_361,In_133);
xor U1269 (N_1269,In_951,In_167);
nand U1270 (N_1270,In_432,In_582);
and U1271 (N_1271,In_350,In_396);
nand U1272 (N_1272,In_527,In_752);
nand U1273 (N_1273,In_795,In_260);
nor U1274 (N_1274,In_972,In_403);
or U1275 (N_1275,In_833,In_661);
nand U1276 (N_1276,In_738,In_165);
nand U1277 (N_1277,In_332,In_557);
or U1278 (N_1278,In_115,In_36);
and U1279 (N_1279,In_817,In_555);
and U1280 (N_1280,In_872,In_195);
nor U1281 (N_1281,In_165,In_907);
nor U1282 (N_1282,In_717,In_797);
and U1283 (N_1283,In_251,In_505);
nand U1284 (N_1284,In_976,In_733);
and U1285 (N_1285,In_318,In_79);
nand U1286 (N_1286,In_956,In_33);
xor U1287 (N_1287,In_997,In_690);
and U1288 (N_1288,In_297,In_133);
nor U1289 (N_1289,In_69,In_85);
nor U1290 (N_1290,In_427,In_623);
nand U1291 (N_1291,In_264,In_242);
or U1292 (N_1292,In_709,In_360);
and U1293 (N_1293,In_647,In_321);
and U1294 (N_1294,In_802,In_726);
nand U1295 (N_1295,In_731,In_982);
nor U1296 (N_1296,In_825,In_56);
or U1297 (N_1297,In_116,In_932);
nand U1298 (N_1298,In_959,In_591);
nor U1299 (N_1299,In_14,In_74);
or U1300 (N_1300,In_479,In_152);
nor U1301 (N_1301,In_632,In_906);
nor U1302 (N_1302,In_980,In_559);
nor U1303 (N_1303,In_334,In_669);
or U1304 (N_1304,In_391,In_729);
and U1305 (N_1305,In_622,In_228);
or U1306 (N_1306,In_291,In_240);
or U1307 (N_1307,In_284,In_169);
nor U1308 (N_1308,In_801,In_241);
nor U1309 (N_1309,In_652,In_746);
nand U1310 (N_1310,In_813,In_300);
and U1311 (N_1311,In_630,In_562);
and U1312 (N_1312,In_732,In_779);
nand U1313 (N_1313,In_812,In_503);
nand U1314 (N_1314,In_337,In_410);
or U1315 (N_1315,In_973,In_747);
nand U1316 (N_1316,In_855,In_111);
or U1317 (N_1317,In_375,In_349);
and U1318 (N_1318,In_739,In_643);
nand U1319 (N_1319,In_689,In_534);
and U1320 (N_1320,In_513,In_80);
nand U1321 (N_1321,In_766,In_488);
or U1322 (N_1322,In_685,In_728);
nand U1323 (N_1323,In_772,In_369);
nand U1324 (N_1324,In_487,In_162);
and U1325 (N_1325,In_760,In_762);
or U1326 (N_1326,In_743,In_921);
nand U1327 (N_1327,In_82,In_656);
nor U1328 (N_1328,In_162,In_824);
nor U1329 (N_1329,In_447,In_99);
nor U1330 (N_1330,In_168,In_566);
nor U1331 (N_1331,In_298,In_108);
and U1332 (N_1332,In_102,In_323);
and U1333 (N_1333,In_646,In_307);
nor U1334 (N_1334,In_989,In_258);
and U1335 (N_1335,In_840,In_294);
and U1336 (N_1336,In_292,In_465);
nor U1337 (N_1337,In_418,In_702);
xor U1338 (N_1338,In_630,In_152);
and U1339 (N_1339,In_66,In_677);
nor U1340 (N_1340,In_634,In_206);
nand U1341 (N_1341,In_918,In_802);
nor U1342 (N_1342,In_40,In_918);
or U1343 (N_1343,In_294,In_132);
and U1344 (N_1344,In_705,In_972);
or U1345 (N_1345,In_983,In_957);
nand U1346 (N_1346,In_739,In_270);
nand U1347 (N_1347,In_885,In_197);
nor U1348 (N_1348,In_97,In_15);
nand U1349 (N_1349,In_881,In_805);
nand U1350 (N_1350,In_699,In_854);
or U1351 (N_1351,In_260,In_502);
nand U1352 (N_1352,In_448,In_896);
and U1353 (N_1353,In_0,In_113);
or U1354 (N_1354,In_213,In_209);
nor U1355 (N_1355,In_628,In_363);
or U1356 (N_1356,In_587,In_495);
and U1357 (N_1357,In_615,In_915);
or U1358 (N_1358,In_489,In_553);
and U1359 (N_1359,In_640,In_125);
nand U1360 (N_1360,In_636,In_196);
nand U1361 (N_1361,In_259,In_619);
or U1362 (N_1362,In_9,In_996);
nor U1363 (N_1363,In_946,In_596);
nor U1364 (N_1364,In_607,In_123);
or U1365 (N_1365,In_190,In_271);
and U1366 (N_1366,In_280,In_693);
or U1367 (N_1367,In_41,In_716);
and U1368 (N_1368,In_507,In_431);
nor U1369 (N_1369,In_266,In_876);
or U1370 (N_1370,In_6,In_356);
nor U1371 (N_1371,In_105,In_343);
nand U1372 (N_1372,In_551,In_466);
nand U1373 (N_1373,In_987,In_410);
nor U1374 (N_1374,In_444,In_430);
and U1375 (N_1375,In_503,In_841);
and U1376 (N_1376,In_567,In_314);
nand U1377 (N_1377,In_98,In_719);
and U1378 (N_1378,In_123,In_705);
nand U1379 (N_1379,In_782,In_389);
or U1380 (N_1380,In_777,In_536);
and U1381 (N_1381,In_754,In_815);
and U1382 (N_1382,In_45,In_0);
nor U1383 (N_1383,In_750,In_798);
nand U1384 (N_1384,In_661,In_930);
nand U1385 (N_1385,In_86,In_488);
nand U1386 (N_1386,In_855,In_143);
nand U1387 (N_1387,In_810,In_466);
nor U1388 (N_1388,In_207,In_62);
nor U1389 (N_1389,In_567,In_736);
nand U1390 (N_1390,In_481,In_678);
nand U1391 (N_1391,In_768,In_627);
or U1392 (N_1392,In_667,In_754);
and U1393 (N_1393,In_463,In_963);
nand U1394 (N_1394,In_232,In_622);
or U1395 (N_1395,In_188,In_331);
nand U1396 (N_1396,In_597,In_204);
nand U1397 (N_1397,In_701,In_498);
or U1398 (N_1398,In_394,In_85);
and U1399 (N_1399,In_492,In_810);
nand U1400 (N_1400,In_580,In_408);
and U1401 (N_1401,In_788,In_53);
nand U1402 (N_1402,In_726,In_812);
nor U1403 (N_1403,In_996,In_774);
nor U1404 (N_1404,In_159,In_275);
nand U1405 (N_1405,In_146,In_699);
nor U1406 (N_1406,In_134,In_951);
or U1407 (N_1407,In_598,In_787);
nor U1408 (N_1408,In_799,In_764);
and U1409 (N_1409,In_567,In_422);
and U1410 (N_1410,In_615,In_86);
nand U1411 (N_1411,In_556,In_85);
and U1412 (N_1412,In_444,In_909);
or U1413 (N_1413,In_593,In_848);
or U1414 (N_1414,In_429,In_127);
nor U1415 (N_1415,In_958,In_286);
or U1416 (N_1416,In_159,In_366);
nor U1417 (N_1417,In_574,In_255);
nand U1418 (N_1418,In_994,In_594);
and U1419 (N_1419,In_188,In_130);
and U1420 (N_1420,In_980,In_736);
or U1421 (N_1421,In_38,In_673);
nand U1422 (N_1422,In_372,In_322);
nor U1423 (N_1423,In_383,In_120);
nand U1424 (N_1424,In_819,In_653);
or U1425 (N_1425,In_808,In_794);
nor U1426 (N_1426,In_823,In_567);
nor U1427 (N_1427,In_172,In_231);
nor U1428 (N_1428,In_523,In_990);
and U1429 (N_1429,In_855,In_456);
nand U1430 (N_1430,In_549,In_39);
and U1431 (N_1431,In_48,In_306);
or U1432 (N_1432,In_406,In_55);
nand U1433 (N_1433,In_803,In_333);
and U1434 (N_1434,In_772,In_333);
nor U1435 (N_1435,In_458,In_654);
nand U1436 (N_1436,In_701,In_998);
nand U1437 (N_1437,In_791,In_78);
and U1438 (N_1438,In_765,In_364);
nor U1439 (N_1439,In_953,In_581);
nand U1440 (N_1440,In_721,In_290);
nor U1441 (N_1441,In_953,In_327);
or U1442 (N_1442,In_720,In_807);
nand U1443 (N_1443,In_703,In_134);
and U1444 (N_1444,In_478,In_985);
nor U1445 (N_1445,In_951,In_333);
nor U1446 (N_1446,In_295,In_302);
nand U1447 (N_1447,In_513,In_480);
and U1448 (N_1448,In_740,In_355);
and U1449 (N_1449,In_339,In_902);
nor U1450 (N_1450,In_88,In_968);
nor U1451 (N_1451,In_513,In_687);
and U1452 (N_1452,In_279,In_85);
nor U1453 (N_1453,In_950,In_332);
nor U1454 (N_1454,In_80,In_10);
nand U1455 (N_1455,In_536,In_604);
nor U1456 (N_1456,In_300,In_591);
and U1457 (N_1457,In_505,In_934);
nor U1458 (N_1458,In_307,In_241);
or U1459 (N_1459,In_885,In_159);
or U1460 (N_1460,In_709,In_533);
or U1461 (N_1461,In_84,In_172);
or U1462 (N_1462,In_206,In_60);
nor U1463 (N_1463,In_335,In_199);
nor U1464 (N_1464,In_34,In_710);
nor U1465 (N_1465,In_7,In_20);
and U1466 (N_1466,In_330,In_681);
nand U1467 (N_1467,In_570,In_599);
nor U1468 (N_1468,In_198,In_200);
or U1469 (N_1469,In_24,In_592);
or U1470 (N_1470,In_818,In_161);
and U1471 (N_1471,In_66,In_864);
nand U1472 (N_1472,In_816,In_741);
nor U1473 (N_1473,In_266,In_521);
nand U1474 (N_1474,In_680,In_770);
nor U1475 (N_1475,In_677,In_75);
nor U1476 (N_1476,In_117,In_98);
nor U1477 (N_1477,In_819,In_727);
and U1478 (N_1478,In_834,In_792);
and U1479 (N_1479,In_90,In_189);
and U1480 (N_1480,In_445,In_425);
or U1481 (N_1481,In_340,In_890);
nor U1482 (N_1482,In_87,In_323);
nor U1483 (N_1483,In_448,In_376);
nor U1484 (N_1484,In_415,In_605);
or U1485 (N_1485,In_291,In_762);
or U1486 (N_1486,In_534,In_598);
or U1487 (N_1487,In_638,In_487);
nand U1488 (N_1488,In_146,In_94);
or U1489 (N_1489,In_906,In_102);
nand U1490 (N_1490,In_575,In_684);
xor U1491 (N_1491,In_678,In_863);
nor U1492 (N_1492,In_416,In_932);
or U1493 (N_1493,In_313,In_28);
or U1494 (N_1494,In_495,In_268);
or U1495 (N_1495,In_835,In_278);
nand U1496 (N_1496,In_346,In_293);
xor U1497 (N_1497,In_518,In_131);
and U1498 (N_1498,In_629,In_236);
nor U1499 (N_1499,In_212,In_862);
nor U1500 (N_1500,In_301,In_383);
and U1501 (N_1501,In_709,In_72);
nor U1502 (N_1502,In_514,In_179);
or U1503 (N_1503,In_473,In_911);
nand U1504 (N_1504,In_506,In_361);
and U1505 (N_1505,In_591,In_274);
or U1506 (N_1506,In_886,In_928);
or U1507 (N_1507,In_73,In_315);
nor U1508 (N_1508,In_953,In_738);
and U1509 (N_1509,In_1,In_425);
xor U1510 (N_1510,In_515,In_386);
nor U1511 (N_1511,In_4,In_671);
nor U1512 (N_1512,In_35,In_780);
or U1513 (N_1513,In_580,In_847);
and U1514 (N_1514,In_742,In_439);
nand U1515 (N_1515,In_421,In_961);
and U1516 (N_1516,In_976,In_297);
or U1517 (N_1517,In_283,In_366);
xor U1518 (N_1518,In_459,In_596);
or U1519 (N_1519,In_490,In_390);
nand U1520 (N_1520,In_442,In_258);
nor U1521 (N_1521,In_345,In_740);
and U1522 (N_1522,In_106,In_236);
and U1523 (N_1523,In_65,In_494);
nor U1524 (N_1524,In_79,In_542);
xnor U1525 (N_1525,In_9,In_410);
or U1526 (N_1526,In_804,In_57);
nor U1527 (N_1527,In_120,In_93);
or U1528 (N_1528,In_153,In_804);
and U1529 (N_1529,In_37,In_988);
or U1530 (N_1530,In_651,In_799);
xor U1531 (N_1531,In_947,In_744);
nand U1532 (N_1532,In_901,In_416);
nand U1533 (N_1533,In_212,In_605);
nor U1534 (N_1534,In_164,In_814);
and U1535 (N_1535,In_500,In_995);
and U1536 (N_1536,In_14,In_749);
nor U1537 (N_1537,In_135,In_607);
nor U1538 (N_1538,In_289,In_569);
nand U1539 (N_1539,In_677,In_350);
nor U1540 (N_1540,In_45,In_542);
nand U1541 (N_1541,In_122,In_483);
nor U1542 (N_1542,In_271,In_132);
nand U1543 (N_1543,In_663,In_208);
nand U1544 (N_1544,In_153,In_694);
nor U1545 (N_1545,In_740,In_215);
nand U1546 (N_1546,In_654,In_555);
or U1547 (N_1547,In_481,In_927);
or U1548 (N_1548,In_491,In_145);
or U1549 (N_1549,In_336,In_755);
nand U1550 (N_1550,In_515,In_369);
nor U1551 (N_1551,In_477,In_548);
xor U1552 (N_1552,In_167,In_642);
and U1553 (N_1553,In_850,In_544);
or U1554 (N_1554,In_109,In_296);
nand U1555 (N_1555,In_998,In_107);
nor U1556 (N_1556,In_817,In_282);
nand U1557 (N_1557,In_554,In_865);
or U1558 (N_1558,In_50,In_822);
and U1559 (N_1559,In_459,In_554);
and U1560 (N_1560,In_631,In_749);
nor U1561 (N_1561,In_968,In_338);
nand U1562 (N_1562,In_253,In_815);
or U1563 (N_1563,In_594,In_195);
or U1564 (N_1564,In_461,In_990);
or U1565 (N_1565,In_46,In_307);
or U1566 (N_1566,In_347,In_432);
nor U1567 (N_1567,In_71,In_489);
or U1568 (N_1568,In_851,In_503);
nand U1569 (N_1569,In_536,In_176);
nor U1570 (N_1570,In_92,In_55);
nand U1571 (N_1571,In_725,In_241);
and U1572 (N_1572,In_686,In_747);
or U1573 (N_1573,In_656,In_712);
or U1574 (N_1574,In_981,In_30);
nor U1575 (N_1575,In_438,In_476);
nor U1576 (N_1576,In_708,In_132);
and U1577 (N_1577,In_935,In_864);
nor U1578 (N_1578,In_301,In_755);
nor U1579 (N_1579,In_309,In_771);
nor U1580 (N_1580,In_213,In_612);
nand U1581 (N_1581,In_934,In_824);
nand U1582 (N_1582,In_91,In_640);
and U1583 (N_1583,In_713,In_479);
nand U1584 (N_1584,In_381,In_392);
or U1585 (N_1585,In_383,In_671);
and U1586 (N_1586,In_502,In_771);
or U1587 (N_1587,In_118,In_339);
or U1588 (N_1588,In_603,In_941);
or U1589 (N_1589,In_883,In_212);
or U1590 (N_1590,In_800,In_693);
or U1591 (N_1591,In_862,In_708);
and U1592 (N_1592,In_254,In_223);
and U1593 (N_1593,In_621,In_77);
or U1594 (N_1594,In_164,In_613);
and U1595 (N_1595,In_267,In_793);
or U1596 (N_1596,In_402,In_472);
nor U1597 (N_1597,In_870,In_499);
nand U1598 (N_1598,In_606,In_512);
and U1599 (N_1599,In_515,In_133);
and U1600 (N_1600,In_187,In_193);
or U1601 (N_1601,In_34,In_201);
nor U1602 (N_1602,In_97,In_2);
nand U1603 (N_1603,In_764,In_740);
or U1604 (N_1604,In_337,In_333);
nand U1605 (N_1605,In_62,In_969);
or U1606 (N_1606,In_766,In_392);
nor U1607 (N_1607,In_697,In_174);
nand U1608 (N_1608,In_403,In_490);
and U1609 (N_1609,In_765,In_465);
or U1610 (N_1610,In_711,In_652);
nand U1611 (N_1611,In_627,In_947);
nand U1612 (N_1612,In_829,In_306);
or U1613 (N_1613,In_319,In_820);
nand U1614 (N_1614,In_828,In_51);
and U1615 (N_1615,In_152,In_471);
or U1616 (N_1616,In_175,In_941);
xor U1617 (N_1617,In_685,In_263);
or U1618 (N_1618,In_591,In_670);
nor U1619 (N_1619,In_907,In_69);
nand U1620 (N_1620,In_833,In_44);
nor U1621 (N_1621,In_820,In_254);
nand U1622 (N_1622,In_794,In_224);
and U1623 (N_1623,In_712,In_21);
nand U1624 (N_1624,In_555,In_404);
nor U1625 (N_1625,In_591,In_482);
nor U1626 (N_1626,In_417,In_753);
nor U1627 (N_1627,In_40,In_568);
or U1628 (N_1628,In_946,In_205);
nand U1629 (N_1629,In_978,In_337);
nand U1630 (N_1630,In_359,In_293);
nor U1631 (N_1631,In_669,In_465);
and U1632 (N_1632,In_541,In_98);
or U1633 (N_1633,In_599,In_940);
and U1634 (N_1634,In_666,In_541);
or U1635 (N_1635,In_900,In_19);
and U1636 (N_1636,In_927,In_378);
and U1637 (N_1637,In_877,In_517);
nor U1638 (N_1638,In_446,In_511);
and U1639 (N_1639,In_887,In_321);
nand U1640 (N_1640,In_177,In_350);
or U1641 (N_1641,In_370,In_285);
nand U1642 (N_1642,In_511,In_970);
nand U1643 (N_1643,In_932,In_626);
nor U1644 (N_1644,In_94,In_397);
nor U1645 (N_1645,In_950,In_629);
and U1646 (N_1646,In_252,In_593);
or U1647 (N_1647,In_874,In_816);
and U1648 (N_1648,In_508,In_543);
nor U1649 (N_1649,In_355,In_169);
and U1650 (N_1650,In_495,In_704);
xnor U1651 (N_1651,In_512,In_358);
or U1652 (N_1652,In_909,In_663);
or U1653 (N_1653,In_912,In_245);
xnor U1654 (N_1654,In_960,In_981);
nand U1655 (N_1655,In_741,In_692);
or U1656 (N_1656,In_958,In_680);
nand U1657 (N_1657,In_545,In_4);
or U1658 (N_1658,In_506,In_925);
nor U1659 (N_1659,In_23,In_191);
or U1660 (N_1660,In_145,In_421);
nor U1661 (N_1661,In_631,In_191);
or U1662 (N_1662,In_247,In_131);
nor U1663 (N_1663,In_237,In_561);
nand U1664 (N_1664,In_32,In_236);
or U1665 (N_1665,In_619,In_340);
nor U1666 (N_1666,In_875,In_160);
or U1667 (N_1667,In_732,In_445);
or U1668 (N_1668,In_657,In_321);
xnor U1669 (N_1669,In_412,In_36);
nor U1670 (N_1670,In_408,In_311);
nor U1671 (N_1671,In_614,In_865);
or U1672 (N_1672,In_882,In_822);
and U1673 (N_1673,In_329,In_228);
nor U1674 (N_1674,In_463,In_544);
and U1675 (N_1675,In_730,In_569);
nor U1676 (N_1676,In_105,In_188);
nor U1677 (N_1677,In_994,In_716);
nor U1678 (N_1678,In_873,In_158);
nor U1679 (N_1679,In_341,In_304);
or U1680 (N_1680,In_38,In_843);
nor U1681 (N_1681,In_163,In_296);
or U1682 (N_1682,In_991,In_42);
nor U1683 (N_1683,In_484,In_779);
nor U1684 (N_1684,In_44,In_215);
nor U1685 (N_1685,In_773,In_504);
nor U1686 (N_1686,In_710,In_585);
or U1687 (N_1687,In_283,In_147);
xnor U1688 (N_1688,In_361,In_552);
or U1689 (N_1689,In_142,In_645);
nand U1690 (N_1690,In_757,In_729);
and U1691 (N_1691,In_742,In_762);
nand U1692 (N_1692,In_988,In_799);
and U1693 (N_1693,In_401,In_638);
and U1694 (N_1694,In_753,In_126);
and U1695 (N_1695,In_921,In_448);
nand U1696 (N_1696,In_757,In_61);
nand U1697 (N_1697,In_464,In_819);
nor U1698 (N_1698,In_662,In_169);
or U1699 (N_1699,In_201,In_156);
nor U1700 (N_1700,In_386,In_267);
and U1701 (N_1701,In_580,In_922);
and U1702 (N_1702,In_351,In_789);
nor U1703 (N_1703,In_184,In_122);
and U1704 (N_1704,In_722,In_339);
nor U1705 (N_1705,In_315,In_249);
or U1706 (N_1706,In_187,In_967);
nand U1707 (N_1707,In_510,In_412);
nor U1708 (N_1708,In_412,In_194);
nand U1709 (N_1709,In_990,In_408);
nor U1710 (N_1710,In_628,In_658);
nand U1711 (N_1711,In_530,In_742);
nand U1712 (N_1712,In_345,In_908);
or U1713 (N_1713,In_203,In_978);
or U1714 (N_1714,In_528,In_639);
nor U1715 (N_1715,In_315,In_161);
and U1716 (N_1716,In_139,In_197);
nand U1717 (N_1717,In_5,In_284);
and U1718 (N_1718,In_508,In_887);
and U1719 (N_1719,In_462,In_198);
nand U1720 (N_1720,In_920,In_460);
xnor U1721 (N_1721,In_12,In_367);
or U1722 (N_1722,In_358,In_981);
and U1723 (N_1723,In_242,In_846);
and U1724 (N_1724,In_356,In_392);
xor U1725 (N_1725,In_26,In_759);
nor U1726 (N_1726,In_736,In_959);
or U1727 (N_1727,In_881,In_291);
nand U1728 (N_1728,In_832,In_99);
nor U1729 (N_1729,In_0,In_811);
and U1730 (N_1730,In_77,In_682);
or U1731 (N_1731,In_103,In_994);
or U1732 (N_1732,In_249,In_907);
and U1733 (N_1733,In_686,In_239);
nor U1734 (N_1734,In_430,In_541);
nor U1735 (N_1735,In_668,In_204);
and U1736 (N_1736,In_407,In_718);
and U1737 (N_1737,In_491,In_582);
nor U1738 (N_1738,In_151,In_514);
or U1739 (N_1739,In_666,In_34);
nand U1740 (N_1740,In_194,In_819);
nor U1741 (N_1741,In_827,In_189);
and U1742 (N_1742,In_150,In_932);
and U1743 (N_1743,In_271,In_909);
xnor U1744 (N_1744,In_651,In_630);
nor U1745 (N_1745,In_976,In_993);
nand U1746 (N_1746,In_751,In_87);
nand U1747 (N_1747,In_988,In_672);
and U1748 (N_1748,In_947,In_505);
and U1749 (N_1749,In_376,In_91);
nor U1750 (N_1750,In_942,In_756);
xnor U1751 (N_1751,In_925,In_984);
or U1752 (N_1752,In_84,In_735);
nor U1753 (N_1753,In_859,In_512);
nor U1754 (N_1754,In_190,In_347);
or U1755 (N_1755,In_10,In_471);
xor U1756 (N_1756,In_522,In_426);
and U1757 (N_1757,In_277,In_488);
xor U1758 (N_1758,In_755,In_48);
and U1759 (N_1759,In_941,In_40);
or U1760 (N_1760,In_699,In_672);
and U1761 (N_1761,In_677,In_842);
and U1762 (N_1762,In_746,In_734);
and U1763 (N_1763,In_316,In_333);
and U1764 (N_1764,In_12,In_740);
and U1765 (N_1765,In_453,In_682);
or U1766 (N_1766,In_939,In_84);
or U1767 (N_1767,In_906,In_283);
or U1768 (N_1768,In_707,In_88);
nand U1769 (N_1769,In_111,In_482);
and U1770 (N_1770,In_854,In_921);
and U1771 (N_1771,In_693,In_492);
and U1772 (N_1772,In_741,In_119);
or U1773 (N_1773,In_374,In_20);
and U1774 (N_1774,In_427,In_343);
nand U1775 (N_1775,In_737,In_377);
nand U1776 (N_1776,In_49,In_488);
nor U1777 (N_1777,In_978,In_547);
nor U1778 (N_1778,In_598,In_378);
nor U1779 (N_1779,In_634,In_459);
and U1780 (N_1780,In_1,In_738);
or U1781 (N_1781,In_679,In_157);
or U1782 (N_1782,In_407,In_843);
and U1783 (N_1783,In_349,In_2);
nand U1784 (N_1784,In_460,In_370);
and U1785 (N_1785,In_665,In_727);
nand U1786 (N_1786,In_859,In_591);
or U1787 (N_1787,In_735,In_381);
and U1788 (N_1788,In_157,In_257);
and U1789 (N_1789,In_537,In_354);
nor U1790 (N_1790,In_761,In_410);
nor U1791 (N_1791,In_208,In_1);
or U1792 (N_1792,In_615,In_735);
nand U1793 (N_1793,In_747,In_718);
or U1794 (N_1794,In_669,In_696);
nor U1795 (N_1795,In_847,In_578);
nand U1796 (N_1796,In_275,In_681);
nor U1797 (N_1797,In_693,In_208);
and U1798 (N_1798,In_324,In_804);
nor U1799 (N_1799,In_150,In_914);
nor U1800 (N_1800,In_503,In_732);
and U1801 (N_1801,In_725,In_530);
and U1802 (N_1802,In_465,In_241);
nor U1803 (N_1803,In_295,In_351);
nand U1804 (N_1804,In_328,In_467);
nor U1805 (N_1805,In_348,In_521);
and U1806 (N_1806,In_953,In_424);
xor U1807 (N_1807,In_216,In_275);
nor U1808 (N_1808,In_944,In_742);
nand U1809 (N_1809,In_90,In_907);
and U1810 (N_1810,In_257,In_771);
and U1811 (N_1811,In_790,In_685);
nor U1812 (N_1812,In_707,In_538);
nor U1813 (N_1813,In_841,In_337);
nand U1814 (N_1814,In_345,In_895);
nor U1815 (N_1815,In_832,In_890);
and U1816 (N_1816,In_89,In_550);
or U1817 (N_1817,In_281,In_229);
xor U1818 (N_1818,In_741,In_930);
nand U1819 (N_1819,In_389,In_647);
nor U1820 (N_1820,In_926,In_534);
nor U1821 (N_1821,In_218,In_950);
and U1822 (N_1822,In_512,In_904);
nand U1823 (N_1823,In_653,In_300);
and U1824 (N_1824,In_324,In_784);
and U1825 (N_1825,In_552,In_135);
nand U1826 (N_1826,In_47,In_543);
and U1827 (N_1827,In_630,In_859);
or U1828 (N_1828,In_211,In_311);
xor U1829 (N_1829,In_895,In_13);
nor U1830 (N_1830,In_428,In_562);
or U1831 (N_1831,In_988,In_903);
and U1832 (N_1832,In_366,In_468);
nand U1833 (N_1833,In_788,In_777);
nand U1834 (N_1834,In_586,In_889);
or U1835 (N_1835,In_521,In_488);
nor U1836 (N_1836,In_536,In_877);
nor U1837 (N_1837,In_369,In_992);
and U1838 (N_1838,In_659,In_426);
nand U1839 (N_1839,In_368,In_820);
or U1840 (N_1840,In_554,In_800);
and U1841 (N_1841,In_522,In_417);
and U1842 (N_1842,In_614,In_471);
or U1843 (N_1843,In_963,In_931);
nor U1844 (N_1844,In_784,In_977);
and U1845 (N_1845,In_31,In_935);
or U1846 (N_1846,In_25,In_696);
nor U1847 (N_1847,In_967,In_740);
or U1848 (N_1848,In_318,In_219);
and U1849 (N_1849,In_465,In_801);
nor U1850 (N_1850,In_581,In_338);
nor U1851 (N_1851,In_438,In_561);
nor U1852 (N_1852,In_42,In_920);
nand U1853 (N_1853,In_973,In_649);
nand U1854 (N_1854,In_426,In_430);
nor U1855 (N_1855,In_990,In_559);
nand U1856 (N_1856,In_397,In_254);
nand U1857 (N_1857,In_593,In_686);
or U1858 (N_1858,In_895,In_258);
nand U1859 (N_1859,In_642,In_823);
nor U1860 (N_1860,In_34,In_11);
or U1861 (N_1861,In_436,In_3);
nand U1862 (N_1862,In_487,In_873);
nand U1863 (N_1863,In_619,In_15);
nor U1864 (N_1864,In_697,In_943);
or U1865 (N_1865,In_191,In_150);
and U1866 (N_1866,In_960,In_283);
and U1867 (N_1867,In_421,In_937);
and U1868 (N_1868,In_57,In_588);
or U1869 (N_1869,In_549,In_223);
and U1870 (N_1870,In_840,In_911);
or U1871 (N_1871,In_144,In_777);
or U1872 (N_1872,In_322,In_348);
and U1873 (N_1873,In_498,In_661);
xor U1874 (N_1874,In_320,In_427);
or U1875 (N_1875,In_222,In_574);
xor U1876 (N_1876,In_675,In_6);
or U1877 (N_1877,In_128,In_106);
nor U1878 (N_1878,In_932,In_389);
and U1879 (N_1879,In_34,In_207);
and U1880 (N_1880,In_627,In_314);
and U1881 (N_1881,In_391,In_461);
xor U1882 (N_1882,In_960,In_380);
xor U1883 (N_1883,In_597,In_240);
and U1884 (N_1884,In_884,In_639);
nor U1885 (N_1885,In_740,In_472);
nor U1886 (N_1886,In_605,In_535);
and U1887 (N_1887,In_627,In_216);
and U1888 (N_1888,In_597,In_253);
and U1889 (N_1889,In_804,In_524);
or U1890 (N_1890,In_227,In_113);
and U1891 (N_1891,In_773,In_181);
and U1892 (N_1892,In_511,In_351);
nand U1893 (N_1893,In_366,In_985);
or U1894 (N_1894,In_598,In_8);
nand U1895 (N_1895,In_908,In_900);
and U1896 (N_1896,In_481,In_770);
and U1897 (N_1897,In_675,In_541);
and U1898 (N_1898,In_181,In_613);
or U1899 (N_1899,In_334,In_259);
nor U1900 (N_1900,In_551,In_64);
or U1901 (N_1901,In_172,In_174);
nor U1902 (N_1902,In_96,In_494);
nor U1903 (N_1903,In_210,In_287);
and U1904 (N_1904,In_149,In_530);
nor U1905 (N_1905,In_279,In_778);
nand U1906 (N_1906,In_884,In_74);
or U1907 (N_1907,In_57,In_2);
nand U1908 (N_1908,In_672,In_78);
or U1909 (N_1909,In_885,In_377);
and U1910 (N_1910,In_489,In_362);
or U1911 (N_1911,In_929,In_234);
nand U1912 (N_1912,In_336,In_477);
and U1913 (N_1913,In_804,In_90);
nand U1914 (N_1914,In_190,In_278);
nor U1915 (N_1915,In_48,In_903);
nor U1916 (N_1916,In_701,In_681);
xnor U1917 (N_1917,In_957,In_675);
or U1918 (N_1918,In_105,In_27);
nand U1919 (N_1919,In_488,In_955);
and U1920 (N_1920,In_286,In_84);
and U1921 (N_1921,In_587,In_128);
nor U1922 (N_1922,In_413,In_790);
nor U1923 (N_1923,In_313,In_26);
or U1924 (N_1924,In_50,In_430);
and U1925 (N_1925,In_647,In_508);
nand U1926 (N_1926,In_709,In_71);
nor U1927 (N_1927,In_800,In_859);
nand U1928 (N_1928,In_570,In_699);
nand U1929 (N_1929,In_200,In_231);
nor U1930 (N_1930,In_614,In_535);
nor U1931 (N_1931,In_159,In_684);
nand U1932 (N_1932,In_843,In_369);
xnor U1933 (N_1933,In_24,In_735);
and U1934 (N_1934,In_897,In_713);
nor U1935 (N_1935,In_927,In_74);
or U1936 (N_1936,In_105,In_569);
nor U1937 (N_1937,In_421,In_956);
and U1938 (N_1938,In_399,In_472);
nand U1939 (N_1939,In_260,In_694);
or U1940 (N_1940,In_971,In_768);
nand U1941 (N_1941,In_897,In_63);
or U1942 (N_1942,In_309,In_404);
nand U1943 (N_1943,In_139,In_912);
xnor U1944 (N_1944,In_743,In_355);
nor U1945 (N_1945,In_2,In_761);
or U1946 (N_1946,In_876,In_717);
or U1947 (N_1947,In_683,In_224);
and U1948 (N_1948,In_690,In_696);
nor U1949 (N_1949,In_545,In_40);
nor U1950 (N_1950,In_72,In_408);
nand U1951 (N_1951,In_18,In_14);
nor U1952 (N_1952,In_721,In_925);
nor U1953 (N_1953,In_166,In_446);
or U1954 (N_1954,In_220,In_509);
nand U1955 (N_1955,In_961,In_890);
nand U1956 (N_1956,In_65,In_840);
and U1957 (N_1957,In_256,In_880);
nand U1958 (N_1958,In_999,In_435);
or U1959 (N_1959,In_173,In_794);
xnor U1960 (N_1960,In_670,In_312);
nor U1961 (N_1961,In_134,In_691);
nor U1962 (N_1962,In_486,In_971);
nand U1963 (N_1963,In_675,In_923);
nor U1964 (N_1964,In_6,In_716);
or U1965 (N_1965,In_33,In_51);
nor U1966 (N_1966,In_319,In_330);
and U1967 (N_1967,In_287,In_135);
xor U1968 (N_1968,In_491,In_305);
nand U1969 (N_1969,In_613,In_535);
and U1970 (N_1970,In_882,In_854);
xnor U1971 (N_1971,In_387,In_123);
or U1972 (N_1972,In_475,In_517);
or U1973 (N_1973,In_381,In_403);
nand U1974 (N_1974,In_596,In_269);
nand U1975 (N_1975,In_449,In_78);
and U1976 (N_1976,In_749,In_695);
nor U1977 (N_1977,In_261,In_302);
and U1978 (N_1978,In_659,In_446);
and U1979 (N_1979,In_225,In_708);
or U1980 (N_1980,In_331,In_637);
nor U1981 (N_1981,In_201,In_67);
and U1982 (N_1982,In_553,In_723);
nor U1983 (N_1983,In_50,In_327);
or U1984 (N_1984,In_288,In_217);
nor U1985 (N_1985,In_490,In_444);
xor U1986 (N_1986,In_20,In_648);
or U1987 (N_1987,In_381,In_723);
nor U1988 (N_1988,In_862,In_148);
and U1989 (N_1989,In_617,In_278);
nor U1990 (N_1990,In_29,In_968);
or U1991 (N_1991,In_559,In_387);
nor U1992 (N_1992,In_993,In_780);
and U1993 (N_1993,In_911,In_618);
nor U1994 (N_1994,In_948,In_512);
or U1995 (N_1995,In_336,In_648);
nand U1996 (N_1996,In_975,In_407);
or U1997 (N_1997,In_670,In_616);
nor U1998 (N_1998,In_142,In_748);
or U1999 (N_1999,In_76,In_228);
or U2000 (N_2000,N_1104,N_1526);
nand U2001 (N_2001,N_910,N_1254);
nand U2002 (N_2002,N_300,N_1281);
nand U2003 (N_2003,N_1961,N_768);
and U2004 (N_2004,N_1855,N_1935);
nand U2005 (N_2005,N_1103,N_1069);
or U2006 (N_2006,N_238,N_676);
or U2007 (N_2007,N_1385,N_1882);
or U2008 (N_2008,N_370,N_337);
nand U2009 (N_2009,N_786,N_787);
and U2010 (N_2010,N_1746,N_1464);
nor U2011 (N_2011,N_681,N_271);
xor U2012 (N_2012,N_1373,N_1943);
and U2013 (N_2013,N_1764,N_79);
and U2014 (N_2014,N_798,N_524);
nor U2015 (N_2015,N_1295,N_528);
or U2016 (N_2016,N_215,N_1874);
nor U2017 (N_2017,N_1335,N_1839);
or U2018 (N_2018,N_113,N_9);
and U2019 (N_2019,N_690,N_1794);
or U2020 (N_2020,N_1903,N_1890);
or U2021 (N_2021,N_1793,N_877);
nand U2022 (N_2022,N_1544,N_263);
or U2023 (N_2023,N_430,N_1534);
nor U2024 (N_2024,N_189,N_1367);
or U2025 (N_2025,N_584,N_821);
and U2026 (N_2026,N_921,N_398);
nor U2027 (N_2027,N_726,N_1609);
and U2028 (N_2028,N_851,N_1085);
and U2029 (N_2029,N_399,N_26);
nor U2030 (N_2030,N_423,N_1975);
nor U2031 (N_2031,N_1294,N_1226);
nor U2032 (N_2032,N_1770,N_1167);
or U2033 (N_2033,N_142,N_1590);
nand U2034 (N_2034,N_1704,N_1131);
nand U2035 (N_2035,N_1505,N_171);
nand U2036 (N_2036,N_1790,N_962);
nand U2037 (N_2037,N_606,N_201);
and U2038 (N_2038,N_1520,N_552);
nor U2039 (N_2039,N_465,N_598);
nand U2040 (N_2040,N_581,N_973);
or U2041 (N_2041,N_1743,N_1804);
or U2042 (N_2042,N_273,N_1679);
and U2043 (N_2043,N_1348,N_629);
nand U2044 (N_2044,N_751,N_82);
nor U2045 (N_2045,N_1431,N_1042);
nor U2046 (N_2046,N_449,N_439);
nand U2047 (N_2047,N_1419,N_299);
nor U2048 (N_2048,N_1267,N_344);
or U2049 (N_2049,N_1696,N_1875);
nand U2050 (N_2050,N_551,N_35);
or U2051 (N_2051,N_645,N_1511);
nor U2052 (N_2052,N_68,N_1988);
nand U2053 (N_2053,N_1989,N_1028);
nor U2054 (N_2054,N_794,N_545);
or U2055 (N_2055,N_1691,N_905);
nand U2056 (N_2056,N_863,N_646);
nor U2057 (N_2057,N_1977,N_148);
nor U2058 (N_2058,N_842,N_639);
or U2059 (N_2059,N_145,N_202);
or U2060 (N_2060,N_1249,N_1277);
and U2061 (N_2061,N_364,N_136);
or U2062 (N_2062,N_1260,N_683);
nand U2063 (N_2063,N_334,N_1016);
or U2064 (N_2064,N_1304,N_1135);
nand U2065 (N_2065,N_935,N_998);
and U2066 (N_2066,N_520,N_1991);
nand U2067 (N_2067,N_577,N_1391);
or U2068 (N_2068,N_290,N_812);
nor U2069 (N_2069,N_46,N_895);
nor U2070 (N_2070,N_72,N_941);
or U2071 (N_2071,N_746,N_414);
nor U2072 (N_2072,N_1917,N_924);
nand U2073 (N_2073,N_801,N_1381);
nor U2074 (N_2074,N_1153,N_727);
and U2075 (N_2075,N_1530,N_1633);
and U2076 (N_2076,N_1132,N_1193);
nor U2077 (N_2077,N_953,N_670);
nand U2078 (N_2078,N_1778,N_441);
nor U2079 (N_2079,N_760,N_1824);
nor U2080 (N_2080,N_1774,N_1569);
or U2081 (N_2081,N_1369,N_658);
or U2082 (N_2082,N_1773,N_1081);
nand U2083 (N_2083,N_694,N_1972);
and U2084 (N_2084,N_667,N_235);
and U2085 (N_2085,N_1741,N_1913);
nor U2086 (N_2086,N_731,N_1063);
or U2087 (N_2087,N_1666,N_1289);
or U2088 (N_2088,N_1263,N_1923);
nand U2089 (N_2089,N_892,N_1271);
nor U2090 (N_2090,N_425,N_722);
and U2091 (N_2091,N_1645,N_894);
or U2092 (N_2092,N_617,N_444);
or U2093 (N_2093,N_713,N_1995);
or U2094 (N_2094,N_1138,N_1198);
nand U2095 (N_2095,N_506,N_15);
and U2096 (N_2096,N_1756,N_1230);
and U2097 (N_2097,N_1521,N_1958);
nor U2098 (N_2098,N_567,N_599);
and U2099 (N_2099,N_1291,N_913);
nand U2100 (N_2100,N_226,N_1397);
nand U2101 (N_2101,N_138,N_554);
nor U2102 (N_2102,N_447,N_1967);
nor U2103 (N_2103,N_926,N_592);
and U2104 (N_2104,N_1683,N_338);
nand U2105 (N_2105,N_1358,N_523);
nand U2106 (N_2106,N_1911,N_1716);
nor U2107 (N_2107,N_216,N_1465);
nor U2108 (N_2108,N_395,N_806);
nand U2109 (N_2109,N_1605,N_1041);
nor U2110 (N_2110,N_1018,N_1133);
and U2111 (N_2111,N_254,N_1032);
nor U2112 (N_2112,N_203,N_1043);
or U2113 (N_2113,N_1997,N_67);
and U2114 (N_2114,N_1792,N_1428);
or U2115 (N_2115,N_677,N_1900);
nor U2116 (N_2116,N_418,N_1064);
nand U2117 (N_2117,N_297,N_1768);
nor U2118 (N_2118,N_340,N_1560);
nor U2119 (N_2119,N_1353,N_1719);
nand U2120 (N_2120,N_80,N_1417);
nor U2121 (N_2121,N_224,N_1757);
nor U2122 (N_2122,N_1784,N_600);
and U2123 (N_2123,N_912,N_1079);
nand U2124 (N_2124,N_1910,N_1282);
or U2125 (N_2125,N_361,N_390);
or U2126 (N_2126,N_1459,N_1318);
and U2127 (N_2127,N_1692,N_1467);
and U2128 (N_2128,N_362,N_1581);
and U2129 (N_2129,N_1026,N_1948);
or U2130 (N_2130,N_153,N_1729);
nand U2131 (N_2131,N_1306,N_453);
nor U2132 (N_2132,N_1448,N_73);
nand U2133 (N_2133,N_952,N_165);
nor U2134 (N_2134,N_1216,N_1818);
and U2135 (N_2135,N_633,N_988);
or U2136 (N_2136,N_1234,N_573);
nand U2137 (N_2137,N_1473,N_693);
and U2138 (N_2138,N_377,N_1058);
nor U2139 (N_2139,N_1504,N_967);
nand U2140 (N_2140,N_1585,N_1155);
or U2141 (N_2141,N_1287,N_1493);
nand U2142 (N_2142,N_743,N_1303);
nand U2143 (N_2143,N_999,N_576);
nor U2144 (N_2144,N_1182,N_1765);
or U2145 (N_2145,N_1430,N_1819);
nand U2146 (N_2146,N_473,N_994);
nor U2147 (N_2147,N_940,N_1675);
nand U2148 (N_2148,N_875,N_1019);
nand U2149 (N_2149,N_1107,N_227);
and U2150 (N_2150,N_596,N_682);
nor U2151 (N_2151,N_514,N_446);
and U2152 (N_2152,N_1331,N_69);
and U2153 (N_2153,N_91,N_881);
and U2154 (N_2154,N_1073,N_710);
nor U2155 (N_2155,N_656,N_1412);
nor U2156 (N_2156,N_163,N_415);
nand U2157 (N_2157,N_805,N_1034);
nand U2158 (N_2158,N_276,N_5);
and U2159 (N_2159,N_939,N_649);
or U2160 (N_2160,N_1293,N_1898);
or U2161 (N_2161,N_1405,N_1812);
nand U2162 (N_2162,N_1148,N_1408);
nand U2163 (N_2163,N_450,N_365);
and U2164 (N_2164,N_22,N_306);
and U2165 (N_2165,N_47,N_501);
nand U2166 (N_2166,N_257,N_348);
or U2167 (N_2167,N_1279,N_1524);
and U2168 (N_2168,N_1663,N_1258);
nor U2169 (N_2169,N_1203,N_1432);
or U2170 (N_2170,N_220,N_1747);
nor U2171 (N_2171,N_779,N_1469);
nand U2172 (N_2172,N_985,N_256);
nor U2173 (N_2173,N_661,N_1763);
and U2174 (N_2174,N_1139,N_1496);
or U2175 (N_2175,N_1264,N_25);
nor U2176 (N_2176,N_733,N_1788);
nand U2177 (N_2177,N_1508,N_118);
and U2178 (N_2178,N_979,N_1876);
nor U2179 (N_2179,N_1978,N_1549);
nand U2180 (N_2180,N_1572,N_237);
or U2181 (N_2181,N_1152,N_505);
or U2182 (N_2182,N_307,N_1648);
or U2183 (N_2183,N_652,N_1974);
nand U2184 (N_2184,N_1994,N_852);
and U2185 (N_2185,N_1754,N_1512);
nor U2186 (N_2186,N_129,N_1451);
and U2187 (N_2187,N_1596,N_745);
nand U2188 (N_2188,N_1119,N_1299);
and U2189 (N_2189,N_287,N_1556);
nand U2190 (N_2190,N_1246,N_126);
nand U2191 (N_2191,N_1668,N_1717);
or U2192 (N_2192,N_1895,N_1953);
and U2193 (N_2193,N_1838,N_1965);
and U2194 (N_2194,N_18,N_1191);
or U2195 (N_2195,N_1209,N_1113);
and U2196 (N_2196,N_484,N_1223);
or U2197 (N_2197,N_1364,N_1816);
nor U2198 (N_2198,N_572,N_247);
and U2199 (N_2199,N_927,N_1986);
and U2200 (N_2200,N_897,N_716);
or U2201 (N_2201,N_759,N_1212);
nor U2202 (N_2202,N_6,N_795);
nand U2203 (N_2203,N_1124,N_570);
or U2204 (N_2204,N_283,N_1425);
or U2205 (N_2205,N_380,N_997);
or U2206 (N_2206,N_412,N_1617);
or U2207 (N_2207,N_1087,N_1893);
nand U2208 (N_2208,N_756,N_655);
nand U2209 (N_2209,N_1372,N_566);
or U2210 (N_2210,N_62,N_75);
and U2211 (N_2211,N_359,N_267);
and U2212 (N_2212,N_1632,N_541);
or U2213 (N_2213,N_55,N_900);
and U2214 (N_2214,N_708,N_563);
or U2215 (N_2215,N_1561,N_834);
and U2216 (N_2216,N_1160,N_748);
nor U2217 (N_2217,N_1897,N_408);
nor U2218 (N_2218,N_986,N_1091);
nand U2219 (N_2219,N_1272,N_280);
and U2220 (N_2220,N_864,N_968);
and U2221 (N_2221,N_21,N_784);
nand U2222 (N_2222,N_714,N_1853);
and U2223 (N_2223,N_729,N_1035);
or U2224 (N_2224,N_1563,N_1003);
nand U2225 (N_2225,N_1108,N_1244);
nor U2226 (N_2226,N_146,N_636);
or U2227 (N_2227,N_1492,N_684);
nor U2228 (N_2228,N_144,N_1126);
nor U2229 (N_2229,N_29,N_1607);
or U2230 (N_2230,N_311,N_1421);
nand U2231 (N_2231,N_1460,N_938);
or U2232 (N_2232,N_1368,N_401);
or U2233 (N_2233,N_324,N_546);
nor U2234 (N_2234,N_1414,N_1224);
or U2235 (N_2235,N_1039,N_1462);
nand U2236 (N_2236,N_1439,N_1649);
xnor U2237 (N_2237,N_1865,N_1732);
nor U2238 (N_2238,N_1833,N_137);
nor U2239 (N_2239,N_500,N_54);
or U2240 (N_2240,N_1615,N_702);
nand U2241 (N_2241,N_76,N_312);
nor U2242 (N_2242,N_1049,N_1528);
nor U2243 (N_2243,N_454,N_1575);
and U2244 (N_2244,N_642,N_836);
and U2245 (N_2245,N_1976,N_1134);
or U2246 (N_2246,N_496,N_1030);
nand U2247 (N_2247,N_433,N_1858);
or U2248 (N_2248,N_1721,N_100);
nor U2249 (N_2249,N_1013,N_1905);
or U2250 (N_2250,N_1110,N_1093);
and U2251 (N_2251,N_1273,N_673);
nor U2252 (N_2252,N_835,N_1595);
or U2253 (N_2253,N_281,N_1981);
or U2254 (N_2254,N_1795,N_1005);
nor U2255 (N_2255,N_88,N_149);
and U2256 (N_2256,N_1519,N_815);
nand U2257 (N_2257,N_251,N_375);
nand U2258 (N_2258,N_173,N_250);
and U2259 (N_2259,N_1860,N_1342);
or U2260 (N_2260,N_1761,N_2);
or U2261 (N_2261,N_128,N_1944);
xnor U2262 (N_2262,N_1241,N_689);
and U2263 (N_2263,N_461,N_1695);
nand U2264 (N_2264,N_419,N_1947);
or U2265 (N_2265,N_1475,N_1536);
or U2266 (N_2266,N_1378,N_1352);
or U2267 (N_2267,N_1235,N_1316);
or U2268 (N_2268,N_1709,N_621);
or U2269 (N_2269,N_1051,N_167);
nor U2270 (N_2270,N_1513,N_1600);
nor U2271 (N_2271,N_143,N_1011);
or U2272 (N_2272,N_244,N_1877);
and U2273 (N_2273,N_557,N_1252);
or U2274 (N_2274,N_13,N_510);
and U2275 (N_2275,N_1597,N_252);
nor U2276 (N_2276,N_147,N_1120);
or U2277 (N_2277,N_1939,N_1515);
xnor U2278 (N_2278,N_1627,N_123);
nand U2279 (N_2279,N_363,N_948);
nor U2280 (N_2280,N_791,N_1688);
and U2281 (N_2281,N_1181,N_1338);
nand U2282 (N_2282,N_1843,N_1253);
and U2283 (N_2283,N_550,N_1621);
nor U2284 (N_2284,N_404,N_685);
or U2285 (N_2285,N_186,N_1476);
nand U2286 (N_2286,N_613,N_343);
or U2287 (N_2287,N_161,N_1037);
or U2288 (N_2288,N_824,N_105);
and U2289 (N_2289,N_638,N_177);
nor U2290 (N_2290,N_115,N_1629);
nor U2291 (N_2291,N_773,N_978);
or U2292 (N_2292,N_1737,N_1832);
nand U2293 (N_2293,N_230,N_49);
and U2294 (N_2294,N_1656,N_1546);
xnor U2295 (N_2295,N_777,N_588);
or U2296 (N_2296,N_1340,N_1548);
xor U2297 (N_2297,N_1749,N_1553);
nor U2298 (N_2298,N_918,N_1265);
and U2299 (N_2299,N_1712,N_1298);
nand U2300 (N_2300,N_909,N_1423);
or U2301 (N_2301,N_1933,N_1184);
or U2302 (N_2302,N_427,N_429);
and U2303 (N_2303,N_1047,N_853);
nand U2304 (N_2304,N_160,N_659);
nor U2305 (N_2305,N_28,N_1219);
and U2306 (N_2306,N_1227,N_1275);
nand U2307 (N_2307,N_492,N_886);
nand U2308 (N_2308,N_548,N_885);
and U2309 (N_2309,N_278,N_1742);
nor U2310 (N_2310,N_610,N_116);
or U2311 (N_2311,N_858,N_1361);
xor U2312 (N_2312,N_1570,N_1846);
or U2313 (N_2313,N_243,N_871);
nor U2314 (N_2314,N_1829,N_1738);
nand U2315 (N_2315,N_1969,N_332);
and U2316 (N_2316,N_982,N_992);
or U2317 (N_2317,N_1959,N_1847);
nor U2318 (N_2318,N_1859,N_1229);
nor U2319 (N_2319,N_1760,N_1029);
and U2320 (N_2320,N_1343,N_378);
nor U2321 (N_2321,N_960,N_1886);
nand U2322 (N_2322,N_48,N_603);
nor U2323 (N_2323,N_1157,N_1955);
nand U2324 (N_2324,N_95,N_564);
nor U2325 (N_2325,N_1884,N_1205);
or U2326 (N_2326,N_1831,N_1266);
nand U2327 (N_2327,N_1685,N_1963);
nand U2328 (N_2328,N_1333,N_286);
nand U2329 (N_2329,N_1887,N_1940);
and U2330 (N_2330,N_333,N_1813);
or U2331 (N_2331,N_1589,N_738);
or U2332 (N_2332,N_491,N_1936);
nand U2333 (N_2333,N_1677,N_1214);
nand U2334 (N_2334,N_1835,N_1602);
or U2335 (N_2335,N_1610,N_1236);
nand U2336 (N_2336,N_1731,N_1474);
and U2337 (N_2337,N_1114,N_264);
or U2338 (N_2338,N_1168,N_31);
nor U2339 (N_2339,N_1231,N_975);
nor U2340 (N_2340,N_808,N_1888);
nand U2341 (N_2341,N_458,N_1780);
nand U2342 (N_2342,N_1527,N_1931);
nor U2343 (N_2343,N_1486,N_1021);
and U2344 (N_2344,N_74,N_1066);
and U2345 (N_2345,N_1929,N_1769);
or U2346 (N_2346,N_1268,N_625);
nand U2347 (N_2347,N_555,N_700);
nand U2348 (N_2348,N_1097,N_1837);
and U2349 (N_2349,N_463,N_1753);
and U2350 (N_2350,N_644,N_1440);
or U2351 (N_2351,N_1671,N_1164);
xnor U2352 (N_2352,N_831,N_1517);
and U2353 (N_2353,N_1023,N_951);
nor U2354 (N_2354,N_1159,N_368);
and U2355 (N_2355,N_1388,N_99);
or U2356 (N_2356,N_1611,N_984);
nand U2357 (N_2357,N_1823,N_1466);
or U2358 (N_2358,N_1383,N_1449);
nand U2359 (N_2359,N_1187,N_1418);
nor U2360 (N_2360,N_562,N_1165);
or U2361 (N_2361,N_585,N_1643);
nor U2362 (N_2362,N_981,N_459);
and U2363 (N_2363,N_367,N_1389);
nor U2364 (N_2364,N_1543,N_929);
and U2365 (N_2365,N_1311,N_1797);
nand U2366 (N_2366,N_12,N_1673);
and U2367 (N_2367,N_204,N_819);
nand U2368 (N_2368,N_602,N_1409);
nand U2369 (N_2369,N_1872,N_175);
nand U2370 (N_2370,N_703,N_1601);
nor U2371 (N_2371,N_955,N_274);
nand U2372 (N_2372,N_780,N_1301);
nor U2373 (N_2373,N_1057,N_1463);
or U2374 (N_2374,N_891,N_1626);
nand U2375 (N_2375,N_1470,N_233);
or U2376 (N_2376,N_240,N_1541);
nor U2377 (N_2377,N_241,N_328);
nand U2378 (N_2378,N_972,N_1815);
and U2379 (N_2379,N_1163,N_1048);
and U2380 (N_2380,N_1158,N_1894);
nand U2381 (N_2381,N_1535,N_1270);
nand U2382 (N_2382,N_790,N_342);
nand U2383 (N_2383,N_521,N_1202);
and U2384 (N_2384,N_317,N_1111);
nand U2385 (N_2385,N_1022,N_925);
nand U2386 (N_2386,N_1127,N_1678);
or U2387 (N_2387,N_1118,N_1915);
nand U2388 (N_2388,N_1909,N_1162);
or U2389 (N_2389,N_37,N_931);
nor U2390 (N_2390,N_1879,N_832);
and U2391 (N_2391,N_1970,N_1927);
nor U2392 (N_2392,N_396,N_793);
and U2393 (N_2393,N_1485,N_919);
nand U2394 (N_2394,N_1919,N_1805);
nor U2395 (N_2395,N_1068,N_1151);
nor U2396 (N_2396,N_322,N_1783);
and U2397 (N_2397,N_1891,N_96);
or U2398 (N_2398,N_358,N_901);
nand U2399 (N_2399,N_1603,N_1772);
or U2400 (N_2400,N_862,N_111);
nand U2401 (N_2401,N_519,N_1307);
nand U2402 (N_2402,N_1916,N_1501);
and U2403 (N_2403,N_1146,N_640);
nor U2404 (N_2404,N_878,N_1055);
nor U2405 (N_2405,N_933,N_1889);
nand U2406 (N_2406,N_632,N_1161);
and U2407 (N_2407,N_1382,N_1004);
nor U2408 (N_2408,N_402,N_71);
or U2409 (N_2409,N_130,N_184);
and U2410 (N_2410,N_327,N_990);
and U2411 (N_2411,N_85,N_1053);
nand U2412 (N_2412,N_1437,N_1862);
nand U2413 (N_2413,N_1095,N_697);
nor U2414 (N_2414,N_1341,N_1061);
nor U2415 (N_2415,N_1359,N_33);
or U2416 (N_2416,N_489,N_351);
nand U2417 (N_2417,N_569,N_896);
nand U2418 (N_2418,N_477,N_219);
nor U2419 (N_2419,N_1122,N_1849);
xor U2420 (N_2420,N_42,N_284);
nand U2421 (N_2421,N_961,N_7);
and U2422 (N_2422,N_958,N_65);
and U2423 (N_2423,N_571,N_3);
and U2424 (N_2424,N_1950,N_345);
nand U2425 (N_2425,N_1370,N_275);
and U2426 (N_2426,N_1490,N_957);
nor U2427 (N_2427,N_19,N_1401);
xor U2428 (N_2428,N_1592,N_1210);
nand U2429 (N_2429,N_1908,N_1374);
xor U2430 (N_2430,N_1690,N_457);
nor U2431 (N_2431,N_903,N_906);
nand U2432 (N_2432,N_1559,N_4);
nor U2433 (N_2433,N_1142,N_493);
and U2434 (N_2434,N_1551,N_1274);
nand U2435 (N_2435,N_438,N_0);
nor U2436 (N_2436,N_674,N_182);
nor U2437 (N_2437,N_1098,N_1239);
or U2438 (N_2438,N_1481,N_1150);
and U2439 (N_2439,N_1123,N_316);
nor U2440 (N_2440,N_172,N_305);
and U2441 (N_2441,N_1208,N_498);
nand U2442 (N_2442,N_1290,N_388);
or U2443 (N_2443,N_480,N_1614);
nand U2444 (N_2444,N_1156,N_1101);
or U2445 (N_2445,N_669,N_150);
or U2446 (N_2446,N_908,N_213);
nor U2447 (N_2447,N_174,N_1982);
xor U2448 (N_2448,N_1902,N_108);
nor U2449 (N_2449,N_1925,N_1906);
and U2450 (N_2450,N_1325,N_730);
and U2451 (N_2451,N_758,N_1491);
nand U2452 (N_2452,N_1154,N_977);
and U2453 (N_2453,N_225,N_1577);
and U2454 (N_2454,N_568,N_928);
and U2455 (N_2455,N_1434,N_1722);
nor U2456 (N_2456,N_45,N_1863);
and U2457 (N_2457,N_591,N_1707);
and U2458 (N_2458,N_1094,N_1116);
nand U2459 (N_2459,N_1322,N_350);
and U2460 (N_2460,N_1999,N_579);
and U2461 (N_2461,N_662,N_1755);
nor U2462 (N_2462,N_792,N_1319);
and U2463 (N_2463,N_1129,N_1641);
or U2464 (N_2464,N_134,N_1427);
nand U2465 (N_2465,N_228,N_575);
nand U2466 (N_2466,N_1634,N_1078);
nor U2467 (N_2467,N_755,N_1868);
and U2468 (N_2468,N_1545,N_715);
nor U2469 (N_2469,N_1892,N_1321);
or U2470 (N_2470,N_64,N_52);
xnor U2471 (N_2471,N_1025,N_1062);
and U2472 (N_2472,N_814,N_1635);
and U2473 (N_2473,N_1809,N_1642);
nor U2474 (N_2474,N_1471,N_1308);
nor U2475 (N_2475,N_1144,N_1169);
nand U2476 (N_2476,N_1651,N_270);
or U2477 (N_2477,N_295,N_1215);
or U2478 (N_2478,N_1814,N_1720);
nand U2479 (N_2479,N_304,N_475);
or U2480 (N_2480,N_308,N_10);
and U2481 (N_2481,N_393,N_1736);
or U2482 (N_2482,N_612,N_1392);
nand U2483 (N_2483,N_883,N_1285);
nor U2484 (N_2484,N_1845,N_1752);
or U2485 (N_2485,N_1176,N_329);
and U2486 (N_2486,N_81,N_1881);
nor U2487 (N_2487,N_917,N_1776);
nand U2488 (N_2488,N_347,N_262);
nand U2489 (N_2489,N_1090,N_1194);
nand U2490 (N_2490,N_258,N_1330);
nand U2491 (N_2491,N_387,N_499);
nor U2492 (N_2492,N_1628,N_1584);
and U2493 (N_2493,N_1867,N_117);
nand U2494 (N_2494,N_587,N_1586);
nor U2495 (N_2495,N_1844,N_1362);
nor U2496 (N_2496,N_976,N_1937);
nand U2497 (N_2497,N_1002,N_1646);
xor U2498 (N_2498,N_1109,N_1658);
or U2499 (N_2499,N_1407,N_1604);
or U2500 (N_2500,N_911,N_1750);
and U2501 (N_2501,N_125,N_959);
nand U2502 (N_2502,N_30,N_718);
or U2503 (N_2503,N_1826,N_320);
nor U2504 (N_2504,N_255,N_1442);
or U2505 (N_2505,N_1024,N_1302);
and U2506 (N_2506,N_1350,N_1278);
or U2507 (N_2507,N_107,N_872);
and U2508 (N_2508,N_643,N_1177);
and U2509 (N_2509,N_1670,N_1949);
or U2510 (N_2510,N_1946,N_1957);
xnor U2511 (N_2511,N_428,N_721);
nand U2512 (N_2512,N_809,N_1197);
nor U2513 (N_2513,N_1326,N_1698);
and U2514 (N_2514,N_1713,N_1014);
and U2515 (N_2515,N_1723,N_242);
and U2516 (N_2516,N_970,N_761);
or U2517 (N_2517,N_339,N_511);
nor U2518 (N_2518,N_101,N_615);
nor U2519 (N_2519,N_531,N_512);
nor U2520 (N_2520,N_1482,N_386);
or U2521 (N_2521,N_1587,N_119);
or U2522 (N_2522,N_131,N_1775);
or U2523 (N_2523,N_1121,N_965);
and U2524 (N_2524,N_36,N_1983);
nand U2525 (N_2525,N_942,N_1516);
nor U2526 (N_2526,N_614,N_1071);
and U2527 (N_2527,N_272,N_628);
or U2528 (N_2528,N_293,N_1403);
nor U2529 (N_2529,N_1074,N_1125);
xnor U2530 (N_2530,N_1345,N_1740);
and U2531 (N_2531,N_354,N_1233);
and U2532 (N_2532,N_907,N_1446);
nand U2533 (N_2533,N_781,N_170);
nand U2534 (N_2534,N_650,N_1478);
nor U2535 (N_2535,N_678,N_1089);
nand U2536 (N_2536,N_497,N_717);
and U2537 (N_2537,N_1808,N_1638);
nor U2538 (N_2538,N_92,N_538);
xor U2539 (N_2539,N_1934,N_355);
and U2540 (N_2540,N_728,N_672);
or U2541 (N_2541,N_1687,N_604);
or U2542 (N_2542,N_486,N_695);
and U2543 (N_2543,N_782,N_1537);
nor U2544 (N_2544,N_503,N_1261);
nor U2545 (N_2545,N_874,N_178);
or U2546 (N_2546,N_1489,N_788);
nand U2547 (N_2547,N_1620,N_660);
or U2548 (N_2548,N_462,N_1455);
or U2549 (N_2549,N_1376,N_1075);
nor U2550 (N_2550,N_481,N_156);
and U2551 (N_2551,N_1714,N_1217);
and U2552 (N_2552,N_1284,N_485);
nand U2553 (N_2553,N_336,N_452);
nor U2554 (N_2554,N_106,N_58);
nand U2555 (N_2555,N_288,N_1598);
nor U2556 (N_2556,N_183,N_1568);
or U2557 (N_2557,N_1817,N_802);
nand U2558 (N_2558,N_1457,N_544);
nand U2559 (N_2559,N_389,N_1130);
nor U2560 (N_2560,N_1650,N_893);
nand U2561 (N_2561,N_1447,N_1371);
nor U2562 (N_2562,N_818,N_1309);
and U2563 (N_2563,N_89,N_86);
and U2564 (N_2564,N_1503,N_882);
nand U2565 (N_2565,N_822,N_772);
or U2566 (N_2566,N_223,N_1017);
nand U2567 (N_2567,N_90,N_1386);
and U2568 (N_2568,N_1510,N_487);
xnor U2569 (N_2569,N_622,N_1056);
or U2570 (N_2570,N_460,N_1242);
or U2571 (N_2571,N_826,N_1487);
and U2572 (N_2572,N_711,N_11);
and U2573 (N_2573,N_1394,N_1878);
and U2574 (N_2574,N_1065,N_950);
and U2575 (N_2575,N_1245,N_1213);
nor U2576 (N_2576,N_1238,N_837);
or U2577 (N_2577,N_374,N_1938);
and U2578 (N_2578,N_1077,N_854);
nand U2579 (N_2579,N_1998,N_1317);
or U2580 (N_2580,N_535,N_1038);
and U2581 (N_2581,N_155,N_1672);
or U2582 (N_2582,N_1869,N_1767);
xnor U2583 (N_2583,N_1705,N_200);
or U2584 (N_2584,N_1100,N_1008);
and U2585 (N_2585,N_1170,N_789);
or U2586 (N_2586,N_8,N_1237);
nand U2587 (N_2587,N_766,N_580);
nand U2588 (N_2588,N_1044,N_1701);
nor U2589 (N_2589,N_292,N_861);
or U2590 (N_2590,N_848,N_817);
nor U2591 (N_2591,N_382,N_740);
nand U2592 (N_2592,N_737,N_536);
nand U2593 (N_2593,N_23,N_1864);
nand U2594 (N_2594,N_843,N_739);
nor U2595 (N_2595,N_870,N_889);
or U2596 (N_2596,N_41,N_1010);
nor U2597 (N_2597,N_944,N_688);
or U2598 (N_2598,N_1012,N_1500);
or U2599 (N_2599,N_513,N_1357);
or U2600 (N_2600,N_1708,N_609);
and U2601 (N_2601,N_741,N_811);
or U2602 (N_2602,N_825,N_190);
and U2603 (N_2603,N_1006,N_314);
nor U2604 (N_2604,N_1762,N_1207);
nand U2605 (N_2605,N_561,N_627);
nor U2606 (N_2606,N_1533,N_1759);
nand U2607 (N_2607,N_221,N_1529);
and U2608 (N_2608,N_14,N_196);
nor U2609 (N_2609,N_1320,N_1676);
nor U2610 (N_2610,N_934,N_1802);
nand U2611 (N_2611,N_1576,N_1200);
or U2612 (N_2612,N_518,N_406);
or U2613 (N_2613,N_844,N_1637);
or U2614 (N_2614,N_206,N_282);
nand U2615 (N_2615,N_1914,N_1960);
or U2616 (N_2616,N_110,N_1147);
nand U2617 (N_2617,N_1099,N_679);
or U2618 (N_2618,N_1347,N_1420);
nor U2619 (N_2619,N_1964,N_1472);
and U2620 (N_2620,N_1667,N_816);
and U2621 (N_2621,N_799,N_1225);
nand U2622 (N_2622,N_764,N_914);
nand U2623 (N_2623,N_898,N_611);
and U2624 (N_2624,N_1178,N_1070);
and U2625 (N_2625,N_1599,N_1149);
nor U2626 (N_2626,N_260,N_124);
and U2627 (N_2627,N_1498,N_1112);
and U2628 (N_2628,N_1942,N_318);
xnor U2629 (N_2629,N_325,N_1117);
or U2630 (N_2630,N_185,N_1468);
or U2631 (N_2631,N_1854,N_904);
or U2632 (N_2632,N_1710,N_993);
nor U2633 (N_2633,N_607,N_1803);
nor U2634 (N_2634,N_771,N_734);
nor U2635 (N_2635,N_757,N_1866);
nand U2636 (N_2636,N_44,N_1700);
nand U2637 (N_2637,N_1088,N_1195);
or U2638 (N_2638,N_839,N_529);
and U2639 (N_2639,N_34,N_141);
nor U2640 (N_2640,N_51,N_1140);
and U2641 (N_2641,N_630,N_1941);
and U2642 (N_2642,N_704,N_279);
nand U2643 (N_2643,N_431,N_687);
nand U2644 (N_2644,N_647,N_849);
or U2645 (N_2645,N_93,N_869);
and U2646 (N_2646,N_1662,N_1532);
or U2647 (N_2647,N_1296,N_193);
nor U2648 (N_2648,N_1574,N_266);
and U2649 (N_2649,N_540,N_807);
or U2650 (N_2650,N_1166,N_833);
nor U2651 (N_2651,N_1429,N_234);
and U2652 (N_2652,N_315,N_943);
or U2653 (N_2653,N_1314,N_1619);
nor U2654 (N_2654,N_547,N_1415);
or U2655 (N_2655,N_1199,N_1962);
nand U2656 (N_2656,N_114,N_1329);
or U2657 (N_2657,N_464,N_43);
or U2658 (N_2658,N_1550,N_1618);
and U2659 (N_2659,N_188,N_855);
nand U2660 (N_2660,N_597,N_1665);
nand U2661 (N_2661,N_1228,N_346);
nor U2662 (N_2662,N_663,N_1661);
xnor U2663 (N_2663,N_665,N_1861);
or U2664 (N_2664,N_397,N_890);
nor U2665 (N_2665,N_1647,N_207);
or U2666 (N_2666,N_1789,N_168);
or U2667 (N_2667,N_1172,N_309);
and U2668 (N_2668,N_631,N_164);
nand U2669 (N_2669,N_456,N_634);
and U2670 (N_2670,N_1399,N_1912);
or U2671 (N_2671,N_1734,N_705);
nor U2672 (N_2672,N_1300,N_1435);
nor U2673 (N_2673,N_248,N_77);
or U2674 (N_2674,N_558,N_767);
nor U2675 (N_2675,N_1727,N_626);
nand U2676 (N_2676,N_549,N_1547);
or U2677 (N_2677,N_1377,N_783);
nor U2678 (N_2678,N_556,N_181);
and U2679 (N_2679,N_471,N_1232);
nand U2680 (N_2680,N_1880,N_360);
or U2681 (N_2681,N_1580,N_775);
or U2682 (N_2682,N_1188,N_1497);
or U2683 (N_2683,N_1840,N_653);
nand U2684 (N_2684,N_1128,N_920);
or U2685 (N_2685,N_1211,N_472);
nor U2686 (N_2686,N_620,N_1558);
or U2687 (N_2687,N_1416,N_50);
nand U2688 (N_2688,N_1718,N_1724);
nand U2689 (N_2689,N_470,N_1745);
and U2690 (N_2690,N_1625,N_974);
or U2691 (N_2691,N_1092,N_416);
nor U2692 (N_2692,N_723,N_850);
or U2693 (N_2693,N_1636,N_1286);
nor U2694 (N_2694,N_1883,N_157);
or U2695 (N_2695,N_1539,N_1297);
or U2696 (N_2696,N_1514,N_169);
or U2697 (N_2697,N_102,N_954);
or U2698 (N_2698,N_1441,N_1461);
nor U2699 (N_2699,N_902,N_1992);
nand U2700 (N_2700,N_289,N_437);
and U2701 (N_2701,N_1251,N_785);
nor U2702 (N_2702,N_671,N_1987);
nand U2703 (N_2703,N_1499,N_1644);
nor U2704 (N_2704,N_1332,N_1583);
nand U2705 (N_2705,N_1522,N_341);
nor U2706 (N_2706,N_302,N_1);
or U2707 (N_2707,N_525,N_754);
or U2708 (N_2708,N_1800,N_1821);
or U2709 (N_2709,N_20,N_1046);
and U2710 (N_2710,N_443,N_845);
or U2711 (N_2711,N_1591,N_1945);
nand U2712 (N_2712,N_385,N_1531);
nand U2713 (N_2713,N_371,N_1072);
nand U2714 (N_2714,N_1552,N_1175);
nor U2715 (N_2715,N_532,N_873);
nand U2716 (N_2716,N_1694,N_132);
nor U2717 (N_2717,N_331,N_543);
and U2718 (N_2718,N_515,N_83);
nand U2719 (N_2719,N_502,N_770);
or U2720 (N_2720,N_468,N_87);
or U2721 (N_2721,N_369,N_394);
and U2722 (N_2722,N_553,N_1920);
nor U2723 (N_2723,N_749,N_601);
nand U2724 (N_2724,N_152,N_989);
nand U2725 (N_2725,N_840,N_57);
or U2726 (N_2726,N_956,N_1654);
nor U2727 (N_2727,N_712,N_154);
nand U2728 (N_2728,N_1283,N_239);
nor U2729 (N_2729,N_1339,N_828);
and U2730 (N_2730,N_409,N_744);
and U2731 (N_2731,N_823,N_1806);
and U2732 (N_2732,N_1186,N_533);
nand U2733 (N_2733,N_1564,N_1822);
xor U2734 (N_2734,N_1836,N_1334);
nor U2735 (N_2735,N_373,N_1173);
and U2736 (N_2736,N_1400,N_84);
nand U2737 (N_2737,N_268,N_526);
nor U2738 (N_2738,N_616,N_245);
nor U2739 (N_2739,N_421,N_135);
xnor U2740 (N_2740,N_209,N_1096);
nor U2741 (N_2741,N_53,N_40);
nor U2742 (N_2742,N_542,N_1726);
and U2743 (N_2743,N_1810,N_210);
and U2744 (N_2744,N_949,N_1179);
nand U2745 (N_2745,N_1555,N_778);
or U2746 (N_2746,N_522,N_60);
nand U2747 (N_2747,N_1735,N_635);
and U2748 (N_2748,N_797,N_1766);
nor U2749 (N_2749,N_1183,N_753);
and U2750 (N_2750,N_1438,N_1366);
nor U2751 (N_2751,N_1932,N_559);
nand U2752 (N_2752,N_180,N_1424);
and U2753 (N_2753,N_1660,N_1956);
and U2754 (N_2754,N_1256,N_1608);
or U2755 (N_2755,N_494,N_1387);
nor U2756 (N_2756,N_432,N_208);
nor U2757 (N_2757,N_1777,N_194);
nor U2758 (N_2758,N_1711,N_1433);
nor U2759 (N_2759,N_1922,N_490);
nand U2760 (N_2760,N_158,N_735);
and U2761 (N_2761,N_736,N_205);
or U2762 (N_2762,N_720,N_1171);
nand U2763 (N_2763,N_1031,N_1973);
and U2764 (N_2764,N_236,N_127);
and U2765 (N_2765,N_199,N_1336);
and U2766 (N_2766,N_657,N_59);
or U2767 (N_2767,N_229,N_1578);
nand U2768 (N_2768,N_1483,N_488);
and U2769 (N_2769,N_442,N_1657);
nor U2770 (N_2770,N_403,N_1102);
nor U2771 (N_2771,N_1699,N_1080);
or U2772 (N_2772,N_1518,N_298);
or U2773 (N_2773,N_1054,N_1494);
nor U2774 (N_2774,N_1904,N_922);
nor U2775 (N_2775,N_1921,N_1851);
nor U2776 (N_2776,N_930,N_1422);
and U2777 (N_2777,N_1703,N_1684);
nand U2778 (N_2778,N_987,N_1060);
nor U2779 (N_2779,N_195,N_1848);
nand U2780 (N_2780,N_537,N_63);
and U2781 (N_2781,N_1827,N_1009);
nor U2782 (N_2782,N_1445,N_1706);
xor U2783 (N_2783,N_1189,N_1201);
nor U2784 (N_2784,N_574,N_1984);
xor U2785 (N_2785,N_1395,N_664);
nor U2786 (N_2786,N_517,N_1857);
nor U2787 (N_2787,N_1896,N_1811);
nand U2788 (N_2788,N_122,N_830);
or U2789 (N_2789,N_1739,N_1456);
nor U2790 (N_2790,N_560,N_530);
or U2791 (N_2791,N_269,N_1243);
or U2792 (N_2792,N_1830,N_1240);
nand U2793 (N_2793,N_1280,N_608);
nor U2794 (N_2794,N_451,N_1413);
nor U2795 (N_2795,N_407,N_1484);
nor U2796 (N_2796,N_1192,N_1033);
and U2797 (N_2797,N_1918,N_1758);
nor U2798 (N_2798,N_301,N_594);
nor U2799 (N_2799,N_1444,N_1174);
nand U2800 (N_2800,N_356,N_762);
nor U2801 (N_2801,N_1728,N_696);
and U2802 (N_2802,N_1801,N_1901);
nor U2803 (N_2803,N_218,N_319);
nor U2804 (N_2804,N_1681,N_411);
and U2805 (N_2805,N_641,N_747);
and U2806 (N_2806,N_750,N_1980);
nor U2807 (N_2807,N_353,N_868);
or U2808 (N_2808,N_1375,N_947);
nor U2809 (N_2809,N_1669,N_1796);
nand U2810 (N_2810,N_291,N_1507);
nor U2811 (N_2811,N_249,N_495);
or U2812 (N_2812,N_593,N_420);
nand U2813 (N_2813,N_605,N_1452);
and U2814 (N_2814,N_1479,N_1059);
nor U2815 (N_2815,N_191,N_1751);
xor U2816 (N_2816,N_372,N_277);
and U2817 (N_2817,N_1856,N_796);
nand U2818 (N_2818,N_1825,N_589);
nand U2819 (N_2819,N_1404,N_1027);
nor U2820 (N_2820,N_467,N_66);
or U2821 (N_2821,N_1979,N_915);
or U2822 (N_2822,N_1276,N_483);
and U2823 (N_2823,N_253,N_516);
or U2824 (N_2824,N_1040,N_1411);
xor U2825 (N_2825,N_383,N_1594);
or U2826 (N_2826,N_1871,N_1926);
nor U2827 (N_2827,N_1686,N_479);
and U2828 (N_2828,N_623,N_1488);
nor U2829 (N_2829,N_1453,N_61);
nor U2830 (N_2830,N_774,N_820);
or U2831 (N_2831,N_666,N_668);
nor U2832 (N_2832,N_381,N_648);
nand U2833 (N_2833,N_937,N_436);
or U2834 (N_2834,N_1624,N_1436);
nand U2835 (N_2835,N_804,N_1566);
or U2836 (N_2836,N_392,N_1384);
nand U2837 (N_2837,N_765,N_916);
nand U2838 (N_2838,N_1477,N_1573);
nand U2839 (N_2839,N_349,N_1398);
and U2840 (N_2840,N_565,N_527);
nand U2841 (N_2841,N_1565,N_829);
nor U2842 (N_2842,N_1365,N_38);
and U2843 (N_2843,N_1652,N_1020);
xor U2844 (N_2844,N_1250,N_991);
nand U2845 (N_2845,N_1664,N_1622);
or U2846 (N_2846,N_1593,N_56);
nand U2847 (N_2847,N_1682,N_112);
nand U2848 (N_2848,N_686,N_1410);
and U2849 (N_2849,N_1715,N_98);
nor U2850 (N_2850,N_867,N_159);
or U2851 (N_2851,N_1828,N_1106);
or U2852 (N_2852,N_120,N_1834);
or U2853 (N_2853,N_1402,N_321);
nor U2854 (N_2854,N_32,N_680);
nand U2855 (N_2855,N_448,N_724);
nand U2856 (N_2856,N_1952,N_800);
and U2857 (N_2857,N_222,N_330);
and U2858 (N_2858,N_1380,N_707);
and U2859 (N_2859,N_1786,N_214);
or U2860 (N_2860,N_326,N_1050);
nand U2861 (N_2861,N_1001,N_709);
nand U2862 (N_2862,N_1557,N_1015);
nor U2863 (N_2863,N_582,N_1655);
and U2864 (N_2864,N_880,N_534);
or U2865 (N_2865,N_422,N_78);
nor U2866 (N_2866,N_1495,N_1222);
nor U2867 (N_2867,N_691,N_1346);
or U2868 (N_2868,N_469,N_1288);
xnor U2869 (N_2869,N_1993,N_426);
nor U2870 (N_2870,N_1730,N_1180);
and U2871 (N_2871,N_376,N_846);
xor U2872 (N_2872,N_763,N_133);
nand U2873 (N_2873,N_1990,N_841);
or U2874 (N_2874,N_983,N_1907);
and U2875 (N_2875,N_70,N_742);
or U2876 (N_2876,N_879,N_838);
nor U2877 (N_2877,N_752,N_1145);
and U2878 (N_2878,N_1966,N_1328);
and U2879 (N_2879,N_1930,N_1137);
xor U2880 (N_2880,N_1702,N_259);
or U2881 (N_2881,N_859,N_424);
nand U2882 (N_2882,N_192,N_1725);
or U2883 (N_2883,N_109,N_1312);
or U2884 (N_2884,N_980,N_946);
and U2885 (N_2885,N_445,N_1337);
nor U2886 (N_2886,N_1538,N_1450);
and U2887 (N_2887,N_1779,N_1305);
nand U2888 (N_2888,N_590,N_1349);
nand U2889 (N_2889,N_675,N_701);
nor U2890 (N_2890,N_698,N_945);
or U2891 (N_2891,N_509,N_1351);
or U2892 (N_2892,N_539,N_1870);
nand U2893 (N_2893,N_1744,N_379);
or U2894 (N_2894,N_357,N_827);
or U2895 (N_2895,N_847,N_211);
nor U2896 (N_2896,N_1640,N_964);
nand U2897 (N_2897,N_769,N_1143);
nand U2898 (N_2898,N_654,N_504);
and U2899 (N_2899,N_923,N_583);
and U2900 (N_2900,N_776,N_618);
or U2901 (N_2901,N_1852,N_1680);
or U2902 (N_2902,N_860,N_1406);
and U2903 (N_2903,N_212,N_187);
or U2904 (N_2904,N_1313,N_866);
and U2905 (N_2905,N_198,N_1798);
or U2906 (N_2906,N_1659,N_578);
nand U2907 (N_2907,N_963,N_1220);
nor U2908 (N_2908,N_1689,N_1327);
nand U2909 (N_2909,N_162,N_508);
nand U2910 (N_2910,N_410,N_1363);
or U2911 (N_2911,N_231,N_651);
nor U2912 (N_2912,N_176,N_323);
nor U2913 (N_2913,N_1787,N_803);
nor U2914 (N_2914,N_1509,N_1697);
nor U2915 (N_2915,N_1968,N_476);
nand U2916 (N_2916,N_1396,N_857);
xor U2917 (N_2917,N_706,N_1542);
and U2918 (N_2918,N_1928,N_1355);
nand U2919 (N_2919,N_97,N_1248);
and U2920 (N_2920,N_1105,N_166);
nand U2921 (N_2921,N_1631,N_1579);
nor U2922 (N_2922,N_296,N_391);
nand U2923 (N_2923,N_1076,N_813);
nand U2924 (N_2924,N_966,N_1067);
nor U2925 (N_2925,N_1036,N_719);
nor U2926 (N_2926,N_17,N_996);
or U2927 (N_2927,N_1141,N_1782);
nor U2928 (N_2928,N_1393,N_121);
nand U2929 (N_2929,N_94,N_1443);
nand U2930 (N_2930,N_884,N_285);
nor U2931 (N_2931,N_261,N_1323);
nor U2932 (N_2932,N_1653,N_1842);
or U2933 (N_2933,N_1136,N_1257);
nor U2934 (N_2934,N_313,N_1996);
nand U2935 (N_2935,N_1185,N_1221);
or U2936 (N_2936,N_310,N_969);
nor U2937 (N_2937,N_27,N_624);
nor U2938 (N_2938,N_1315,N_995);
nand U2939 (N_2939,N_1115,N_366);
or U2940 (N_2940,N_1390,N_1255);
and U2941 (N_2941,N_1924,N_1899);
and U2942 (N_2942,N_232,N_434);
and U2943 (N_2943,N_384,N_1567);
nand U2944 (N_2944,N_294,N_1190);
or U2945 (N_2945,N_303,N_1310);
nand U2946 (N_2946,N_466,N_1007);
xnor U2947 (N_2947,N_1850,N_24);
or U2948 (N_2948,N_936,N_1083);
nor U2949 (N_2949,N_1354,N_1523);
nor U2950 (N_2950,N_1082,N_1791);
nor U2951 (N_2951,N_139,N_1454);
nor U2952 (N_2952,N_405,N_352);
and U2953 (N_2953,N_478,N_1084);
and U2954 (N_2954,N_440,N_619);
or U2955 (N_2955,N_1606,N_888);
or U2956 (N_2956,N_1506,N_1502);
or U2957 (N_2957,N_865,N_887);
and U2958 (N_2958,N_1360,N_1262);
nor U2959 (N_2959,N_1540,N_413);
or U2960 (N_2960,N_1324,N_1525);
or U2961 (N_2961,N_1218,N_151);
nor U2962 (N_2962,N_1426,N_1807);
or U2963 (N_2963,N_1693,N_692);
or U2964 (N_2964,N_1196,N_1480);
nor U2965 (N_2965,N_1582,N_179);
nand U2966 (N_2966,N_1841,N_1820);
or U2967 (N_2967,N_1292,N_435);
and U2968 (N_2968,N_1616,N_1951);
nand U2969 (N_2969,N_586,N_699);
or U2970 (N_2970,N_1571,N_1971);
nand U2971 (N_2971,N_335,N_1785);
nor U2972 (N_2972,N_1344,N_637);
nand U2973 (N_2973,N_1204,N_417);
and U2974 (N_2974,N_1873,N_876);
nor U2975 (N_2975,N_140,N_595);
nor U2976 (N_2976,N_1733,N_810);
xnor U2977 (N_2977,N_1458,N_1630);
xnor U2978 (N_2978,N_1045,N_1356);
nor U2979 (N_2979,N_1674,N_1562);
or U2980 (N_2980,N_1639,N_1269);
and U2981 (N_2981,N_1247,N_217);
and U2982 (N_2982,N_1000,N_16);
or U2983 (N_2983,N_265,N_1985);
nand U2984 (N_2984,N_932,N_455);
xnor U2985 (N_2985,N_103,N_507);
and U2986 (N_2986,N_474,N_1799);
nand U2987 (N_2987,N_732,N_856);
and U2988 (N_2988,N_104,N_1206);
and U2989 (N_2989,N_1259,N_1588);
nand U2990 (N_2990,N_1748,N_1781);
nand U2991 (N_2991,N_1613,N_725);
and U2992 (N_2992,N_246,N_899);
nand U2993 (N_2993,N_1379,N_971);
nor U2994 (N_2994,N_1612,N_1623);
xor U2995 (N_2995,N_197,N_1954);
or U2996 (N_2996,N_1771,N_1052);
or U2997 (N_2997,N_482,N_1554);
nor U2998 (N_2998,N_39,N_400);
or U2999 (N_2999,N_1086,N_1885);
and U3000 (N_3000,N_957,N_1037);
or U3001 (N_3001,N_316,N_555);
or U3002 (N_3002,N_1276,N_648);
or U3003 (N_3003,N_792,N_1049);
or U3004 (N_3004,N_1467,N_1818);
nand U3005 (N_3005,N_341,N_1093);
nor U3006 (N_3006,N_221,N_1902);
nand U3007 (N_3007,N_927,N_33);
and U3008 (N_3008,N_1331,N_263);
or U3009 (N_3009,N_694,N_323);
and U3010 (N_3010,N_1928,N_1834);
nor U3011 (N_3011,N_1650,N_1426);
and U3012 (N_3012,N_1710,N_975);
nor U3013 (N_3013,N_1271,N_727);
nor U3014 (N_3014,N_160,N_1252);
and U3015 (N_3015,N_798,N_758);
nand U3016 (N_3016,N_1822,N_1146);
or U3017 (N_3017,N_412,N_282);
nor U3018 (N_3018,N_404,N_97);
nor U3019 (N_3019,N_1492,N_849);
nor U3020 (N_3020,N_105,N_1666);
and U3021 (N_3021,N_1269,N_388);
or U3022 (N_3022,N_1728,N_1826);
nor U3023 (N_3023,N_1321,N_210);
nor U3024 (N_3024,N_697,N_936);
or U3025 (N_3025,N_808,N_1232);
and U3026 (N_3026,N_1970,N_604);
nand U3027 (N_3027,N_212,N_215);
nand U3028 (N_3028,N_859,N_262);
nor U3029 (N_3029,N_1262,N_1623);
nor U3030 (N_3030,N_3,N_1891);
or U3031 (N_3031,N_1796,N_978);
nand U3032 (N_3032,N_359,N_1601);
or U3033 (N_3033,N_985,N_1040);
xnor U3034 (N_3034,N_1142,N_175);
or U3035 (N_3035,N_1531,N_516);
and U3036 (N_3036,N_1947,N_484);
or U3037 (N_3037,N_1226,N_1586);
and U3038 (N_3038,N_702,N_493);
nor U3039 (N_3039,N_1405,N_1241);
nand U3040 (N_3040,N_1678,N_736);
or U3041 (N_3041,N_1344,N_424);
nand U3042 (N_3042,N_1649,N_1567);
nor U3043 (N_3043,N_983,N_1169);
nor U3044 (N_3044,N_1045,N_1347);
and U3045 (N_3045,N_145,N_1233);
nor U3046 (N_3046,N_741,N_1979);
or U3047 (N_3047,N_1971,N_750);
nand U3048 (N_3048,N_645,N_1641);
and U3049 (N_3049,N_874,N_113);
and U3050 (N_3050,N_1776,N_1967);
nor U3051 (N_3051,N_1923,N_1381);
or U3052 (N_3052,N_388,N_973);
or U3053 (N_3053,N_278,N_450);
or U3054 (N_3054,N_1161,N_310);
xnor U3055 (N_3055,N_808,N_72);
nor U3056 (N_3056,N_1400,N_795);
nand U3057 (N_3057,N_619,N_753);
nand U3058 (N_3058,N_1413,N_322);
nor U3059 (N_3059,N_937,N_924);
and U3060 (N_3060,N_1794,N_1096);
and U3061 (N_3061,N_809,N_762);
and U3062 (N_3062,N_1858,N_1775);
or U3063 (N_3063,N_1631,N_396);
or U3064 (N_3064,N_913,N_958);
nand U3065 (N_3065,N_1437,N_1616);
and U3066 (N_3066,N_80,N_1192);
nor U3067 (N_3067,N_1046,N_1913);
nand U3068 (N_3068,N_579,N_739);
and U3069 (N_3069,N_1199,N_1395);
or U3070 (N_3070,N_1302,N_654);
or U3071 (N_3071,N_442,N_1955);
or U3072 (N_3072,N_1276,N_1394);
nor U3073 (N_3073,N_702,N_1621);
or U3074 (N_3074,N_939,N_1130);
and U3075 (N_3075,N_604,N_55);
and U3076 (N_3076,N_1043,N_1201);
and U3077 (N_3077,N_1078,N_10);
and U3078 (N_3078,N_1909,N_1318);
or U3079 (N_3079,N_669,N_1445);
nor U3080 (N_3080,N_1272,N_939);
and U3081 (N_3081,N_1921,N_298);
and U3082 (N_3082,N_294,N_298);
nor U3083 (N_3083,N_812,N_958);
nor U3084 (N_3084,N_1423,N_906);
nand U3085 (N_3085,N_777,N_1603);
nor U3086 (N_3086,N_603,N_703);
xnor U3087 (N_3087,N_248,N_93);
or U3088 (N_3088,N_877,N_1315);
nor U3089 (N_3089,N_142,N_174);
nand U3090 (N_3090,N_1510,N_533);
nand U3091 (N_3091,N_32,N_1317);
and U3092 (N_3092,N_554,N_746);
or U3093 (N_3093,N_785,N_1341);
nor U3094 (N_3094,N_1514,N_495);
or U3095 (N_3095,N_1796,N_259);
and U3096 (N_3096,N_1806,N_69);
and U3097 (N_3097,N_984,N_56);
nand U3098 (N_3098,N_486,N_50);
nand U3099 (N_3099,N_146,N_21);
or U3100 (N_3100,N_1277,N_1737);
and U3101 (N_3101,N_506,N_358);
or U3102 (N_3102,N_292,N_1863);
or U3103 (N_3103,N_1146,N_189);
nor U3104 (N_3104,N_1599,N_55);
nor U3105 (N_3105,N_1678,N_224);
nor U3106 (N_3106,N_1224,N_1738);
nor U3107 (N_3107,N_1140,N_558);
nand U3108 (N_3108,N_1326,N_1412);
and U3109 (N_3109,N_708,N_1218);
nand U3110 (N_3110,N_440,N_379);
nor U3111 (N_3111,N_1289,N_768);
and U3112 (N_3112,N_813,N_341);
or U3113 (N_3113,N_1722,N_894);
or U3114 (N_3114,N_475,N_231);
nor U3115 (N_3115,N_479,N_194);
xor U3116 (N_3116,N_1814,N_1584);
nand U3117 (N_3117,N_741,N_627);
nor U3118 (N_3118,N_316,N_1986);
nor U3119 (N_3119,N_1644,N_1178);
and U3120 (N_3120,N_1179,N_1090);
nor U3121 (N_3121,N_161,N_1044);
nor U3122 (N_3122,N_1227,N_1536);
or U3123 (N_3123,N_492,N_1175);
or U3124 (N_3124,N_1054,N_990);
nor U3125 (N_3125,N_1226,N_1577);
nand U3126 (N_3126,N_893,N_955);
nand U3127 (N_3127,N_973,N_260);
or U3128 (N_3128,N_1148,N_1288);
nand U3129 (N_3129,N_615,N_333);
or U3130 (N_3130,N_1603,N_1233);
or U3131 (N_3131,N_1716,N_600);
and U3132 (N_3132,N_819,N_890);
nand U3133 (N_3133,N_1170,N_1539);
nand U3134 (N_3134,N_798,N_1540);
and U3135 (N_3135,N_1777,N_299);
or U3136 (N_3136,N_551,N_843);
nor U3137 (N_3137,N_1757,N_1291);
nor U3138 (N_3138,N_1175,N_1875);
or U3139 (N_3139,N_494,N_1452);
or U3140 (N_3140,N_360,N_387);
nand U3141 (N_3141,N_1927,N_719);
or U3142 (N_3142,N_113,N_524);
or U3143 (N_3143,N_1879,N_106);
or U3144 (N_3144,N_945,N_122);
and U3145 (N_3145,N_428,N_479);
nand U3146 (N_3146,N_343,N_1334);
and U3147 (N_3147,N_1262,N_1475);
and U3148 (N_3148,N_1287,N_1879);
nand U3149 (N_3149,N_1343,N_1120);
and U3150 (N_3150,N_102,N_1942);
nand U3151 (N_3151,N_285,N_870);
nor U3152 (N_3152,N_100,N_35);
nor U3153 (N_3153,N_248,N_216);
or U3154 (N_3154,N_16,N_1267);
nand U3155 (N_3155,N_900,N_787);
nand U3156 (N_3156,N_1344,N_1694);
nor U3157 (N_3157,N_1281,N_56);
or U3158 (N_3158,N_530,N_1538);
nand U3159 (N_3159,N_1060,N_1613);
nor U3160 (N_3160,N_328,N_975);
or U3161 (N_3161,N_502,N_1840);
nor U3162 (N_3162,N_1019,N_989);
nor U3163 (N_3163,N_1047,N_1448);
and U3164 (N_3164,N_237,N_818);
and U3165 (N_3165,N_1055,N_1504);
or U3166 (N_3166,N_1873,N_980);
or U3167 (N_3167,N_672,N_510);
and U3168 (N_3168,N_1914,N_410);
nand U3169 (N_3169,N_1665,N_1272);
or U3170 (N_3170,N_490,N_664);
and U3171 (N_3171,N_458,N_1753);
and U3172 (N_3172,N_330,N_1109);
and U3173 (N_3173,N_1421,N_1654);
xor U3174 (N_3174,N_1556,N_1902);
nand U3175 (N_3175,N_577,N_548);
or U3176 (N_3176,N_255,N_1644);
nor U3177 (N_3177,N_1379,N_1584);
or U3178 (N_3178,N_255,N_1208);
or U3179 (N_3179,N_527,N_37);
nor U3180 (N_3180,N_1940,N_528);
nand U3181 (N_3181,N_1071,N_1417);
or U3182 (N_3182,N_1217,N_1956);
and U3183 (N_3183,N_321,N_138);
xor U3184 (N_3184,N_1154,N_521);
or U3185 (N_3185,N_1358,N_1646);
nand U3186 (N_3186,N_244,N_54);
or U3187 (N_3187,N_1532,N_770);
nand U3188 (N_3188,N_477,N_1605);
nor U3189 (N_3189,N_1550,N_1161);
nor U3190 (N_3190,N_986,N_1893);
nor U3191 (N_3191,N_1819,N_858);
nand U3192 (N_3192,N_1313,N_585);
nand U3193 (N_3193,N_67,N_1498);
nand U3194 (N_3194,N_1620,N_942);
nand U3195 (N_3195,N_1744,N_1455);
nand U3196 (N_3196,N_1894,N_1133);
nor U3197 (N_3197,N_88,N_344);
or U3198 (N_3198,N_337,N_459);
nand U3199 (N_3199,N_1656,N_631);
nand U3200 (N_3200,N_632,N_1468);
or U3201 (N_3201,N_1851,N_858);
and U3202 (N_3202,N_909,N_554);
and U3203 (N_3203,N_244,N_912);
and U3204 (N_3204,N_616,N_1548);
nor U3205 (N_3205,N_527,N_447);
nor U3206 (N_3206,N_1905,N_1659);
and U3207 (N_3207,N_1093,N_108);
nand U3208 (N_3208,N_112,N_166);
or U3209 (N_3209,N_192,N_1597);
and U3210 (N_3210,N_307,N_514);
nor U3211 (N_3211,N_161,N_68);
nor U3212 (N_3212,N_484,N_130);
or U3213 (N_3213,N_522,N_1369);
xor U3214 (N_3214,N_926,N_1845);
and U3215 (N_3215,N_976,N_1916);
nor U3216 (N_3216,N_682,N_1443);
nor U3217 (N_3217,N_1310,N_213);
and U3218 (N_3218,N_1299,N_191);
or U3219 (N_3219,N_1832,N_1154);
nand U3220 (N_3220,N_234,N_157);
or U3221 (N_3221,N_1119,N_244);
or U3222 (N_3222,N_779,N_756);
nor U3223 (N_3223,N_1397,N_450);
and U3224 (N_3224,N_1047,N_376);
nand U3225 (N_3225,N_1708,N_1191);
nor U3226 (N_3226,N_1551,N_881);
nand U3227 (N_3227,N_346,N_220);
nor U3228 (N_3228,N_1154,N_706);
or U3229 (N_3229,N_1514,N_1240);
or U3230 (N_3230,N_1201,N_1666);
or U3231 (N_3231,N_1856,N_764);
or U3232 (N_3232,N_1172,N_1942);
or U3233 (N_3233,N_1727,N_599);
nand U3234 (N_3234,N_125,N_108);
or U3235 (N_3235,N_1204,N_797);
and U3236 (N_3236,N_501,N_1764);
and U3237 (N_3237,N_133,N_1993);
or U3238 (N_3238,N_1659,N_632);
nor U3239 (N_3239,N_1409,N_616);
nor U3240 (N_3240,N_807,N_423);
nand U3241 (N_3241,N_1224,N_336);
nand U3242 (N_3242,N_1686,N_306);
nor U3243 (N_3243,N_839,N_1843);
or U3244 (N_3244,N_1091,N_591);
nor U3245 (N_3245,N_1464,N_727);
or U3246 (N_3246,N_134,N_1109);
nand U3247 (N_3247,N_595,N_0);
or U3248 (N_3248,N_1233,N_178);
nand U3249 (N_3249,N_722,N_666);
and U3250 (N_3250,N_1025,N_375);
and U3251 (N_3251,N_1273,N_725);
nor U3252 (N_3252,N_463,N_1435);
nor U3253 (N_3253,N_1623,N_894);
or U3254 (N_3254,N_1261,N_196);
or U3255 (N_3255,N_669,N_434);
nor U3256 (N_3256,N_1608,N_1672);
and U3257 (N_3257,N_1136,N_1104);
nor U3258 (N_3258,N_603,N_792);
nor U3259 (N_3259,N_636,N_150);
nand U3260 (N_3260,N_242,N_79);
xnor U3261 (N_3261,N_1097,N_195);
nand U3262 (N_3262,N_1962,N_1926);
and U3263 (N_3263,N_27,N_42);
nand U3264 (N_3264,N_630,N_1796);
or U3265 (N_3265,N_1768,N_1722);
nand U3266 (N_3266,N_822,N_1677);
nor U3267 (N_3267,N_1285,N_1207);
and U3268 (N_3268,N_1718,N_1623);
and U3269 (N_3269,N_1890,N_944);
nand U3270 (N_3270,N_1351,N_1871);
xnor U3271 (N_3271,N_827,N_300);
nor U3272 (N_3272,N_806,N_925);
or U3273 (N_3273,N_748,N_1588);
and U3274 (N_3274,N_1831,N_902);
nor U3275 (N_3275,N_68,N_1755);
nor U3276 (N_3276,N_73,N_1653);
nor U3277 (N_3277,N_1504,N_1223);
or U3278 (N_3278,N_171,N_104);
and U3279 (N_3279,N_130,N_872);
nor U3280 (N_3280,N_323,N_1513);
and U3281 (N_3281,N_970,N_1007);
or U3282 (N_3282,N_1891,N_1416);
nand U3283 (N_3283,N_870,N_1305);
nand U3284 (N_3284,N_1306,N_1667);
nand U3285 (N_3285,N_1936,N_1515);
xnor U3286 (N_3286,N_967,N_76);
and U3287 (N_3287,N_187,N_1594);
nor U3288 (N_3288,N_211,N_1211);
nand U3289 (N_3289,N_881,N_308);
nand U3290 (N_3290,N_1506,N_1745);
nand U3291 (N_3291,N_606,N_110);
nand U3292 (N_3292,N_1415,N_89);
or U3293 (N_3293,N_1267,N_165);
and U3294 (N_3294,N_388,N_611);
nand U3295 (N_3295,N_1595,N_1736);
nand U3296 (N_3296,N_455,N_121);
nand U3297 (N_3297,N_881,N_1318);
nor U3298 (N_3298,N_186,N_1723);
nand U3299 (N_3299,N_992,N_1559);
or U3300 (N_3300,N_346,N_952);
nand U3301 (N_3301,N_662,N_1169);
or U3302 (N_3302,N_144,N_733);
xor U3303 (N_3303,N_563,N_660);
nor U3304 (N_3304,N_1488,N_58);
nand U3305 (N_3305,N_1699,N_743);
and U3306 (N_3306,N_548,N_1720);
nand U3307 (N_3307,N_999,N_1731);
nand U3308 (N_3308,N_1144,N_112);
nor U3309 (N_3309,N_247,N_1571);
or U3310 (N_3310,N_958,N_1336);
and U3311 (N_3311,N_733,N_1153);
or U3312 (N_3312,N_897,N_715);
nor U3313 (N_3313,N_755,N_812);
or U3314 (N_3314,N_1993,N_870);
nand U3315 (N_3315,N_714,N_1629);
nand U3316 (N_3316,N_77,N_118);
and U3317 (N_3317,N_1878,N_1588);
or U3318 (N_3318,N_720,N_150);
nand U3319 (N_3319,N_1010,N_87);
nor U3320 (N_3320,N_1567,N_443);
nand U3321 (N_3321,N_72,N_1270);
or U3322 (N_3322,N_1067,N_1044);
and U3323 (N_3323,N_563,N_1759);
nand U3324 (N_3324,N_1001,N_66);
nor U3325 (N_3325,N_1964,N_652);
and U3326 (N_3326,N_1573,N_640);
nand U3327 (N_3327,N_21,N_1037);
nand U3328 (N_3328,N_624,N_487);
and U3329 (N_3329,N_1655,N_1153);
nand U3330 (N_3330,N_1532,N_1079);
or U3331 (N_3331,N_1099,N_1935);
and U3332 (N_3332,N_1964,N_1452);
nor U3333 (N_3333,N_301,N_1598);
or U3334 (N_3334,N_1492,N_954);
nand U3335 (N_3335,N_720,N_555);
and U3336 (N_3336,N_1927,N_182);
and U3337 (N_3337,N_593,N_1410);
xor U3338 (N_3338,N_1904,N_1972);
or U3339 (N_3339,N_134,N_1094);
nand U3340 (N_3340,N_1959,N_1377);
nor U3341 (N_3341,N_1688,N_1570);
or U3342 (N_3342,N_1218,N_433);
and U3343 (N_3343,N_1898,N_1561);
and U3344 (N_3344,N_1144,N_169);
nand U3345 (N_3345,N_1696,N_1280);
or U3346 (N_3346,N_1636,N_794);
or U3347 (N_3347,N_258,N_1211);
and U3348 (N_3348,N_1639,N_774);
or U3349 (N_3349,N_401,N_1481);
or U3350 (N_3350,N_103,N_668);
and U3351 (N_3351,N_702,N_1830);
nor U3352 (N_3352,N_86,N_935);
nand U3353 (N_3353,N_993,N_1380);
and U3354 (N_3354,N_1396,N_1193);
or U3355 (N_3355,N_1605,N_42);
nor U3356 (N_3356,N_241,N_1949);
and U3357 (N_3357,N_228,N_818);
nor U3358 (N_3358,N_1104,N_437);
and U3359 (N_3359,N_392,N_1837);
and U3360 (N_3360,N_373,N_79);
or U3361 (N_3361,N_1463,N_1177);
and U3362 (N_3362,N_1579,N_1800);
nor U3363 (N_3363,N_315,N_1950);
or U3364 (N_3364,N_1786,N_1424);
nand U3365 (N_3365,N_1007,N_916);
or U3366 (N_3366,N_835,N_549);
nor U3367 (N_3367,N_984,N_650);
nand U3368 (N_3368,N_1873,N_1316);
or U3369 (N_3369,N_1932,N_80);
or U3370 (N_3370,N_411,N_559);
and U3371 (N_3371,N_1173,N_43);
or U3372 (N_3372,N_1645,N_1787);
nor U3373 (N_3373,N_967,N_1422);
or U3374 (N_3374,N_595,N_1306);
or U3375 (N_3375,N_1592,N_1136);
nor U3376 (N_3376,N_1637,N_1287);
xnor U3377 (N_3377,N_95,N_773);
and U3378 (N_3378,N_1601,N_1488);
or U3379 (N_3379,N_1077,N_923);
nand U3380 (N_3380,N_1821,N_1646);
nand U3381 (N_3381,N_1110,N_1238);
and U3382 (N_3382,N_1962,N_1908);
and U3383 (N_3383,N_1465,N_668);
nand U3384 (N_3384,N_1734,N_1771);
and U3385 (N_3385,N_1308,N_1743);
and U3386 (N_3386,N_636,N_1988);
or U3387 (N_3387,N_351,N_1935);
or U3388 (N_3388,N_1133,N_243);
or U3389 (N_3389,N_1619,N_805);
or U3390 (N_3390,N_358,N_466);
nor U3391 (N_3391,N_770,N_1063);
nand U3392 (N_3392,N_1658,N_1608);
nand U3393 (N_3393,N_1772,N_1999);
or U3394 (N_3394,N_102,N_731);
nand U3395 (N_3395,N_145,N_1982);
nor U3396 (N_3396,N_1732,N_1866);
or U3397 (N_3397,N_1518,N_506);
and U3398 (N_3398,N_1028,N_1090);
nand U3399 (N_3399,N_1554,N_1619);
nor U3400 (N_3400,N_734,N_762);
nor U3401 (N_3401,N_1238,N_300);
or U3402 (N_3402,N_1018,N_1973);
or U3403 (N_3403,N_159,N_1657);
and U3404 (N_3404,N_1316,N_1502);
and U3405 (N_3405,N_1686,N_187);
nor U3406 (N_3406,N_1327,N_1321);
nand U3407 (N_3407,N_568,N_1520);
nor U3408 (N_3408,N_1126,N_1529);
or U3409 (N_3409,N_1676,N_1808);
nand U3410 (N_3410,N_527,N_1040);
and U3411 (N_3411,N_191,N_136);
nand U3412 (N_3412,N_1459,N_1848);
or U3413 (N_3413,N_397,N_706);
nand U3414 (N_3414,N_61,N_423);
and U3415 (N_3415,N_1315,N_163);
or U3416 (N_3416,N_1053,N_815);
and U3417 (N_3417,N_970,N_1531);
nand U3418 (N_3418,N_1659,N_818);
and U3419 (N_3419,N_507,N_1878);
nand U3420 (N_3420,N_1272,N_406);
nand U3421 (N_3421,N_379,N_619);
nand U3422 (N_3422,N_1389,N_3);
or U3423 (N_3423,N_1168,N_1547);
nor U3424 (N_3424,N_1223,N_1368);
nor U3425 (N_3425,N_1440,N_1721);
and U3426 (N_3426,N_879,N_253);
and U3427 (N_3427,N_517,N_1253);
or U3428 (N_3428,N_946,N_1751);
nand U3429 (N_3429,N_1903,N_314);
nor U3430 (N_3430,N_1299,N_1072);
nor U3431 (N_3431,N_1528,N_1061);
nor U3432 (N_3432,N_984,N_1645);
and U3433 (N_3433,N_248,N_1105);
nor U3434 (N_3434,N_962,N_1307);
nand U3435 (N_3435,N_1239,N_1915);
nor U3436 (N_3436,N_1851,N_35);
nor U3437 (N_3437,N_504,N_1845);
nand U3438 (N_3438,N_1425,N_1601);
nor U3439 (N_3439,N_85,N_1552);
nor U3440 (N_3440,N_262,N_248);
nand U3441 (N_3441,N_1956,N_1122);
nand U3442 (N_3442,N_56,N_1790);
and U3443 (N_3443,N_1797,N_102);
nor U3444 (N_3444,N_830,N_209);
or U3445 (N_3445,N_863,N_25);
and U3446 (N_3446,N_469,N_1135);
or U3447 (N_3447,N_1500,N_30);
or U3448 (N_3448,N_315,N_555);
and U3449 (N_3449,N_25,N_1605);
nand U3450 (N_3450,N_1233,N_863);
or U3451 (N_3451,N_696,N_1993);
and U3452 (N_3452,N_312,N_692);
and U3453 (N_3453,N_1445,N_1178);
or U3454 (N_3454,N_159,N_1028);
or U3455 (N_3455,N_1246,N_1917);
xnor U3456 (N_3456,N_576,N_1268);
or U3457 (N_3457,N_1682,N_116);
nand U3458 (N_3458,N_536,N_210);
or U3459 (N_3459,N_148,N_1187);
or U3460 (N_3460,N_108,N_22);
nor U3461 (N_3461,N_1189,N_1115);
nand U3462 (N_3462,N_1125,N_431);
nor U3463 (N_3463,N_1837,N_1146);
nor U3464 (N_3464,N_1456,N_1467);
and U3465 (N_3465,N_1053,N_1102);
and U3466 (N_3466,N_1144,N_1738);
or U3467 (N_3467,N_1343,N_350);
nor U3468 (N_3468,N_433,N_576);
nor U3469 (N_3469,N_157,N_1941);
nor U3470 (N_3470,N_249,N_989);
nand U3471 (N_3471,N_1969,N_960);
or U3472 (N_3472,N_1007,N_1670);
and U3473 (N_3473,N_1171,N_1263);
or U3474 (N_3474,N_309,N_667);
nand U3475 (N_3475,N_1239,N_1952);
or U3476 (N_3476,N_183,N_824);
nand U3477 (N_3477,N_69,N_1266);
nand U3478 (N_3478,N_250,N_68);
or U3479 (N_3479,N_1348,N_1537);
and U3480 (N_3480,N_1108,N_452);
or U3481 (N_3481,N_742,N_197);
or U3482 (N_3482,N_1335,N_297);
and U3483 (N_3483,N_719,N_947);
or U3484 (N_3484,N_1935,N_1647);
nand U3485 (N_3485,N_1345,N_1755);
or U3486 (N_3486,N_965,N_1801);
nor U3487 (N_3487,N_356,N_1323);
nand U3488 (N_3488,N_1484,N_1668);
nand U3489 (N_3489,N_547,N_1012);
nor U3490 (N_3490,N_183,N_36);
and U3491 (N_3491,N_1205,N_272);
or U3492 (N_3492,N_937,N_522);
nand U3493 (N_3493,N_966,N_894);
nand U3494 (N_3494,N_190,N_1494);
nand U3495 (N_3495,N_319,N_873);
nand U3496 (N_3496,N_755,N_1088);
nand U3497 (N_3497,N_1205,N_304);
nand U3498 (N_3498,N_558,N_1603);
and U3499 (N_3499,N_540,N_1397);
nor U3500 (N_3500,N_1421,N_321);
or U3501 (N_3501,N_1706,N_1111);
xor U3502 (N_3502,N_240,N_1770);
and U3503 (N_3503,N_220,N_96);
nor U3504 (N_3504,N_1427,N_433);
or U3505 (N_3505,N_45,N_1236);
and U3506 (N_3506,N_75,N_912);
nor U3507 (N_3507,N_1207,N_1132);
nand U3508 (N_3508,N_1456,N_4);
nand U3509 (N_3509,N_1611,N_777);
and U3510 (N_3510,N_474,N_515);
or U3511 (N_3511,N_135,N_1079);
nor U3512 (N_3512,N_1880,N_830);
nand U3513 (N_3513,N_853,N_718);
nand U3514 (N_3514,N_1440,N_859);
and U3515 (N_3515,N_1351,N_1407);
nor U3516 (N_3516,N_296,N_643);
and U3517 (N_3517,N_863,N_1901);
nor U3518 (N_3518,N_126,N_100);
or U3519 (N_3519,N_156,N_1116);
nand U3520 (N_3520,N_1045,N_1558);
or U3521 (N_3521,N_603,N_264);
and U3522 (N_3522,N_1829,N_345);
nor U3523 (N_3523,N_1142,N_224);
nand U3524 (N_3524,N_8,N_476);
nand U3525 (N_3525,N_800,N_816);
nand U3526 (N_3526,N_1800,N_1781);
and U3527 (N_3527,N_1035,N_1485);
and U3528 (N_3528,N_1625,N_1864);
nand U3529 (N_3529,N_341,N_970);
nand U3530 (N_3530,N_1221,N_664);
nor U3531 (N_3531,N_1221,N_234);
nand U3532 (N_3532,N_3,N_354);
and U3533 (N_3533,N_1240,N_1519);
and U3534 (N_3534,N_1574,N_1124);
or U3535 (N_3535,N_361,N_228);
or U3536 (N_3536,N_1549,N_1218);
nor U3537 (N_3537,N_1774,N_1211);
and U3538 (N_3538,N_1350,N_125);
or U3539 (N_3539,N_52,N_626);
and U3540 (N_3540,N_1861,N_1340);
nor U3541 (N_3541,N_182,N_1183);
nor U3542 (N_3542,N_1325,N_333);
nor U3543 (N_3543,N_1,N_510);
nor U3544 (N_3544,N_1391,N_1395);
or U3545 (N_3545,N_244,N_1653);
nand U3546 (N_3546,N_1422,N_1218);
nor U3547 (N_3547,N_1354,N_251);
or U3548 (N_3548,N_729,N_66);
and U3549 (N_3549,N_389,N_103);
or U3550 (N_3550,N_932,N_462);
or U3551 (N_3551,N_360,N_1926);
or U3552 (N_3552,N_287,N_1254);
or U3553 (N_3553,N_1144,N_558);
or U3554 (N_3554,N_1298,N_1448);
and U3555 (N_3555,N_675,N_1837);
nand U3556 (N_3556,N_408,N_1274);
nor U3557 (N_3557,N_1952,N_368);
or U3558 (N_3558,N_1391,N_1456);
or U3559 (N_3559,N_1661,N_796);
nand U3560 (N_3560,N_878,N_1468);
or U3561 (N_3561,N_1477,N_1121);
nand U3562 (N_3562,N_1842,N_1029);
nor U3563 (N_3563,N_399,N_450);
or U3564 (N_3564,N_722,N_632);
nand U3565 (N_3565,N_659,N_29);
nand U3566 (N_3566,N_1003,N_621);
nand U3567 (N_3567,N_964,N_273);
or U3568 (N_3568,N_1412,N_1183);
nor U3569 (N_3569,N_1631,N_1850);
nor U3570 (N_3570,N_1310,N_1914);
nor U3571 (N_3571,N_685,N_521);
and U3572 (N_3572,N_297,N_160);
nand U3573 (N_3573,N_600,N_1698);
and U3574 (N_3574,N_493,N_1846);
and U3575 (N_3575,N_1634,N_833);
nor U3576 (N_3576,N_1280,N_1347);
nand U3577 (N_3577,N_1617,N_523);
nor U3578 (N_3578,N_518,N_1274);
or U3579 (N_3579,N_1234,N_900);
or U3580 (N_3580,N_296,N_268);
nand U3581 (N_3581,N_435,N_1178);
nor U3582 (N_3582,N_368,N_273);
and U3583 (N_3583,N_710,N_1695);
nand U3584 (N_3584,N_689,N_1394);
and U3585 (N_3585,N_215,N_501);
and U3586 (N_3586,N_496,N_956);
and U3587 (N_3587,N_1788,N_704);
or U3588 (N_3588,N_1176,N_171);
nor U3589 (N_3589,N_104,N_824);
nor U3590 (N_3590,N_616,N_1158);
and U3591 (N_3591,N_845,N_381);
and U3592 (N_3592,N_651,N_743);
or U3593 (N_3593,N_893,N_648);
nand U3594 (N_3594,N_70,N_159);
or U3595 (N_3595,N_1506,N_115);
nor U3596 (N_3596,N_1248,N_970);
nand U3597 (N_3597,N_1453,N_113);
or U3598 (N_3598,N_1395,N_1821);
nor U3599 (N_3599,N_1362,N_640);
or U3600 (N_3600,N_1464,N_1732);
nand U3601 (N_3601,N_1077,N_1187);
nand U3602 (N_3602,N_904,N_939);
nand U3603 (N_3603,N_93,N_1350);
or U3604 (N_3604,N_800,N_877);
or U3605 (N_3605,N_337,N_1978);
and U3606 (N_3606,N_655,N_502);
nor U3607 (N_3607,N_592,N_740);
or U3608 (N_3608,N_499,N_1181);
nor U3609 (N_3609,N_698,N_805);
and U3610 (N_3610,N_369,N_247);
nor U3611 (N_3611,N_1152,N_385);
nand U3612 (N_3612,N_945,N_899);
or U3613 (N_3613,N_1690,N_1662);
and U3614 (N_3614,N_1974,N_600);
or U3615 (N_3615,N_1792,N_1377);
nor U3616 (N_3616,N_527,N_1606);
and U3617 (N_3617,N_70,N_144);
and U3618 (N_3618,N_1600,N_871);
nor U3619 (N_3619,N_650,N_695);
or U3620 (N_3620,N_108,N_373);
or U3621 (N_3621,N_1004,N_151);
nand U3622 (N_3622,N_1480,N_1937);
nor U3623 (N_3623,N_40,N_1087);
nor U3624 (N_3624,N_1425,N_1370);
or U3625 (N_3625,N_648,N_1876);
or U3626 (N_3626,N_314,N_1508);
nand U3627 (N_3627,N_471,N_143);
nor U3628 (N_3628,N_1896,N_1189);
and U3629 (N_3629,N_1849,N_467);
nor U3630 (N_3630,N_1328,N_945);
nor U3631 (N_3631,N_1909,N_812);
nand U3632 (N_3632,N_1563,N_254);
and U3633 (N_3633,N_1797,N_1317);
nor U3634 (N_3634,N_1083,N_1780);
nand U3635 (N_3635,N_1774,N_1388);
nor U3636 (N_3636,N_1893,N_419);
nor U3637 (N_3637,N_1455,N_1740);
and U3638 (N_3638,N_88,N_483);
nor U3639 (N_3639,N_702,N_1574);
and U3640 (N_3640,N_952,N_1588);
nor U3641 (N_3641,N_285,N_865);
or U3642 (N_3642,N_120,N_1085);
or U3643 (N_3643,N_1984,N_681);
nand U3644 (N_3644,N_1344,N_854);
xor U3645 (N_3645,N_424,N_1578);
and U3646 (N_3646,N_1179,N_1490);
or U3647 (N_3647,N_1370,N_707);
or U3648 (N_3648,N_1938,N_869);
nor U3649 (N_3649,N_401,N_460);
nand U3650 (N_3650,N_1339,N_1179);
nor U3651 (N_3651,N_1073,N_1664);
and U3652 (N_3652,N_1530,N_1300);
nor U3653 (N_3653,N_1865,N_61);
nor U3654 (N_3654,N_190,N_1235);
nand U3655 (N_3655,N_1242,N_1234);
nand U3656 (N_3656,N_1588,N_729);
and U3657 (N_3657,N_246,N_365);
and U3658 (N_3658,N_1503,N_268);
or U3659 (N_3659,N_1848,N_7);
and U3660 (N_3660,N_646,N_148);
nand U3661 (N_3661,N_110,N_177);
nor U3662 (N_3662,N_1094,N_569);
nand U3663 (N_3663,N_1667,N_885);
nand U3664 (N_3664,N_1041,N_762);
nor U3665 (N_3665,N_918,N_722);
nand U3666 (N_3666,N_397,N_1934);
nor U3667 (N_3667,N_247,N_1695);
or U3668 (N_3668,N_887,N_241);
or U3669 (N_3669,N_331,N_601);
or U3670 (N_3670,N_1582,N_1168);
or U3671 (N_3671,N_65,N_1904);
and U3672 (N_3672,N_1786,N_901);
and U3673 (N_3673,N_1198,N_664);
nor U3674 (N_3674,N_548,N_1223);
nand U3675 (N_3675,N_1247,N_531);
nand U3676 (N_3676,N_1755,N_1381);
or U3677 (N_3677,N_1123,N_1453);
and U3678 (N_3678,N_1589,N_528);
nand U3679 (N_3679,N_995,N_1875);
nor U3680 (N_3680,N_863,N_1230);
nor U3681 (N_3681,N_97,N_347);
nor U3682 (N_3682,N_707,N_1580);
nor U3683 (N_3683,N_798,N_722);
nor U3684 (N_3684,N_235,N_475);
or U3685 (N_3685,N_1582,N_138);
or U3686 (N_3686,N_318,N_977);
and U3687 (N_3687,N_384,N_930);
or U3688 (N_3688,N_1648,N_1158);
or U3689 (N_3689,N_1645,N_1013);
and U3690 (N_3690,N_1223,N_805);
and U3691 (N_3691,N_749,N_1703);
xnor U3692 (N_3692,N_528,N_349);
or U3693 (N_3693,N_1646,N_1565);
nand U3694 (N_3694,N_1169,N_1522);
nand U3695 (N_3695,N_1126,N_1490);
nand U3696 (N_3696,N_617,N_317);
nand U3697 (N_3697,N_568,N_314);
nor U3698 (N_3698,N_1747,N_1434);
and U3699 (N_3699,N_824,N_714);
and U3700 (N_3700,N_1234,N_1346);
nor U3701 (N_3701,N_640,N_652);
and U3702 (N_3702,N_1280,N_1268);
nand U3703 (N_3703,N_1125,N_1149);
or U3704 (N_3704,N_152,N_553);
nand U3705 (N_3705,N_516,N_1783);
nor U3706 (N_3706,N_1287,N_1982);
nor U3707 (N_3707,N_1432,N_539);
and U3708 (N_3708,N_68,N_1169);
nor U3709 (N_3709,N_342,N_1623);
nor U3710 (N_3710,N_201,N_1670);
or U3711 (N_3711,N_799,N_251);
or U3712 (N_3712,N_1847,N_252);
or U3713 (N_3713,N_1200,N_1103);
and U3714 (N_3714,N_683,N_1881);
nor U3715 (N_3715,N_269,N_1981);
nand U3716 (N_3716,N_925,N_1437);
nand U3717 (N_3717,N_1967,N_664);
nand U3718 (N_3718,N_179,N_135);
and U3719 (N_3719,N_764,N_271);
and U3720 (N_3720,N_214,N_122);
nor U3721 (N_3721,N_1024,N_651);
nand U3722 (N_3722,N_1811,N_48);
nor U3723 (N_3723,N_1586,N_729);
nand U3724 (N_3724,N_1065,N_784);
nand U3725 (N_3725,N_1216,N_1170);
nand U3726 (N_3726,N_815,N_1261);
and U3727 (N_3727,N_457,N_360);
xor U3728 (N_3728,N_1442,N_1947);
nor U3729 (N_3729,N_792,N_1976);
and U3730 (N_3730,N_1104,N_677);
nand U3731 (N_3731,N_1932,N_1500);
and U3732 (N_3732,N_1051,N_261);
nor U3733 (N_3733,N_440,N_174);
and U3734 (N_3734,N_203,N_1443);
nand U3735 (N_3735,N_1614,N_808);
and U3736 (N_3736,N_1785,N_1450);
nor U3737 (N_3737,N_1657,N_341);
and U3738 (N_3738,N_75,N_1406);
or U3739 (N_3739,N_311,N_1075);
nand U3740 (N_3740,N_791,N_1960);
or U3741 (N_3741,N_1235,N_1332);
or U3742 (N_3742,N_754,N_336);
nand U3743 (N_3743,N_752,N_1880);
nand U3744 (N_3744,N_1384,N_241);
and U3745 (N_3745,N_1399,N_460);
nor U3746 (N_3746,N_466,N_763);
nor U3747 (N_3747,N_1756,N_967);
nand U3748 (N_3748,N_1842,N_306);
nand U3749 (N_3749,N_1879,N_1436);
and U3750 (N_3750,N_1962,N_1773);
nand U3751 (N_3751,N_1833,N_1334);
nand U3752 (N_3752,N_602,N_1907);
or U3753 (N_3753,N_1576,N_1457);
nand U3754 (N_3754,N_1879,N_194);
nor U3755 (N_3755,N_1045,N_64);
nor U3756 (N_3756,N_1179,N_1115);
nor U3757 (N_3757,N_1043,N_768);
nor U3758 (N_3758,N_276,N_1806);
nor U3759 (N_3759,N_379,N_635);
and U3760 (N_3760,N_536,N_1772);
or U3761 (N_3761,N_1225,N_268);
nor U3762 (N_3762,N_982,N_1402);
nor U3763 (N_3763,N_1000,N_1767);
or U3764 (N_3764,N_895,N_464);
and U3765 (N_3765,N_1509,N_958);
or U3766 (N_3766,N_856,N_843);
and U3767 (N_3767,N_399,N_172);
xor U3768 (N_3768,N_896,N_443);
and U3769 (N_3769,N_1701,N_168);
nor U3770 (N_3770,N_888,N_441);
nor U3771 (N_3771,N_739,N_1809);
nand U3772 (N_3772,N_485,N_71);
or U3773 (N_3773,N_1930,N_732);
nand U3774 (N_3774,N_1517,N_1709);
and U3775 (N_3775,N_1718,N_1796);
and U3776 (N_3776,N_350,N_979);
nor U3777 (N_3777,N_319,N_1450);
and U3778 (N_3778,N_1859,N_942);
nor U3779 (N_3779,N_1915,N_985);
nor U3780 (N_3780,N_1036,N_1214);
nor U3781 (N_3781,N_399,N_194);
and U3782 (N_3782,N_1007,N_737);
or U3783 (N_3783,N_1521,N_1577);
and U3784 (N_3784,N_1005,N_1916);
and U3785 (N_3785,N_1000,N_1802);
nand U3786 (N_3786,N_684,N_1988);
and U3787 (N_3787,N_994,N_1839);
or U3788 (N_3788,N_702,N_1609);
nor U3789 (N_3789,N_272,N_259);
and U3790 (N_3790,N_1628,N_1911);
and U3791 (N_3791,N_1690,N_849);
and U3792 (N_3792,N_1180,N_1457);
nor U3793 (N_3793,N_212,N_506);
xor U3794 (N_3794,N_412,N_673);
and U3795 (N_3795,N_1282,N_1696);
nor U3796 (N_3796,N_88,N_1034);
and U3797 (N_3797,N_714,N_1800);
and U3798 (N_3798,N_1349,N_1136);
nor U3799 (N_3799,N_23,N_1179);
nor U3800 (N_3800,N_1938,N_1641);
nor U3801 (N_3801,N_941,N_920);
nor U3802 (N_3802,N_1455,N_90);
or U3803 (N_3803,N_1053,N_374);
nand U3804 (N_3804,N_1484,N_1060);
nor U3805 (N_3805,N_1044,N_628);
nand U3806 (N_3806,N_1447,N_446);
or U3807 (N_3807,N_48,N_91);
and U3808 (N_3808,N_1964,N_1436);
or U3809 (N_3809,N_588,N_607);
nor U3810 (N_3810,N_1064,N_487);
nand U3811 (N_3811,N_999,N_969);
nor U3812 (N_3812,N_697,N_1685);
or U3813 (N_3813,N_1177,N_1107);
xor U3814 (N_3814,N_1223,N_881);
and U3815 (N_3815,N_43,N_1832);
nor U3816 (N_3816,N_239,N_329);
nor U3817 (N_3817,N_1418,N_903);
nand U3818 (N_3818,N_824,N_779);
nor U3819 (N_3819,N_246,N_1044);
and U3820 (N_3820,N_529,N_1473);
or U3821 (N_3821,N_180,N_422);
or U3822 (N_3822,N_1096,N_149);
nor U3823 (N_3823,N_1261,N_1553);
nand U3824 (N_3824,N_1337,N_56);
and U3825 (N_3825,N_929,N_324);
or U3826 (N_3826,N_1082,N_69);
nand U3827 (N_3827,N_836,N_1049);
and U3828 (N_3828,N_821,N_1861);
or U3829 (N_3829,N_690,N_227);
nor U3830 (N_3830,N_1772,N_1304);
nor U3831 (N_3831,N_1348,N_152);
nand U3832 (N_3832,N_1684,N_1790);
nor U3833 (N_3833,N_1350,N_1062);
nor U3834 (N_3834,N_1548,N_545);
nor U3835 (N_3835,N_1052,N_425);
nor U3836 (N_3836,N_1295,N_681);
and U3837 (N_3837,N_1220,N_1050);
nor U3838 (N_3838,N_1424,N_114);
nand U3839 (N_3839,N_433,N_1554);
nor U3840 (N_3840,N_159,N_804);
or U3841 (N_3841,N_938,N_998);
and U3842 (N_3842,N_1688,N_148);
nand U3843 (N_3843,N_118,N_366);
nor U3844 (N_3844,N_108,N_1601);
and U3845 (N_3845,N_122,N_808);
nor U3846 (N_3846,N_173,N_1156);
nand U3847 (N_3847,N_383,N_1279);
nor U3848 (N_3848,N_476,N_954);
nor U3849 (N_3849,N_851,N_1049);
or U3850 (N_3850,N_1373,N_606);
nor U3851 (N_3851,N_801,N_1073);
nor U3852 (N_3852,N_518,N_1727);
and U3853 (N_3853,N_1882,N_1479);
nor U3854 (N_3854,N_1166,N_370);
or U3855 (N_3855,N_918,N_1695);
and U3856 (N_3856,N_707,N_996);
xor U3857 (N_3857,N_708,N_1702);
or U3858 (N_3858,N_1720,N_1635);
nand U3859 (N_3859,N_669,N_766);
or U3860 (N_3860,N_1504,N_278);
nand U3861 (N_3861,N_1328,N_1943);
or U3862 (N_3862,N_1326,N_1643);
and U3863 (N_3863,N_850,N_947);
nor U3864 (N_3864,N_1457,N_1692);
and U3865 (N_3865,N_1421,N_859);
nand U3866 (N_3866,N_984,N_463);
and U3867 (N_3867,N_1837,N_864);
and U3868 (N_3868,N_758,N_842);
and U3869 (N_3869,N_1694,N_1301);
nor U3870 (N_3870,N_1455,N_1872);
nor U3871 (N_3871,N_38,N_986);
nor U3872 (N_3872,N_183,N_49);
and U3873 (N_3873,N_995,N_1798);
nor U3874 (N_3874,N_1972,N_37);
and U3875 (N_3875,N_820,N_1666);
nand U3876 (N_3876,N_1749,N_1913);
and U3877 (N_3877,N_141,N_529);
or U3878 (N_3878,N_839,N_989);
and U3879 (N_3879,N_1206,N_1663);
and U3880 (N_3880,N_150,N_509);
or U3881 (N_3881,N_720,N_207);
nand U3882 (N_3882,N_758,N_1804);
nand U3883 (N_3883,N_975,N_84);
nand U3884 (N_3884,N_1056,N_665);
nand U3885 (N_3885,N_1574,N_286);
and U3886 (N_3886,N_1593,N_58);
nor U3887 (N_3887,N_1764,N_1950);
or U3888 (N_3888,N_1991,N_404);
nor U3889 (N_3889,N_1593,N_302);
or U3890 (N_3890,N_1076,N_1077);
nor U3891 (N_3891,N_1806,N_1777);
nor U3892 (N_3892,N_1496,N_1195);
nand U3893 (N_3893,N_1718,N_1553);
or U3894 (N_3894,N_770,N_641);
nor U3895 (N_3895,N_460,N_616);
and U3896 (N_3896,N_393,N_611);
or U3897 (N_3897,N_754,N_438);
or U3898 (N_3898,N_1127,N_938);
nor U3899 (N_3899,N_916,N_1805);
nand U3900 (N_3900,N_1344,N_88);
and U3901 (N_3901,N_1290,N_1531);
nor U3902 (N_3902,N_1366,N_1675);
and U3903 (N_3903,N_365,N_452);
or U3904 (N_3904,N_1250,N_334);
and U3905 (N_3905,N_35,N_213);
or U3906 (N_3906,N_426,N_474);
nor U3907 (N_3907,N_119,N_163);
nand U3908 (N_3908,N_1005,N_9);
or U3909 (N_3909,N_1220,N_1639);
and U3910 (N_3910,N_1005,N_1597);
or U3911 (N_3911,N_1439,N_1496);
nor U3912 (N_3912,N_1699,N_521);
and U3913 (N_3913,N_1728,N_229);
and U3914 (N_3914,N_1505,N_572);
and U3915 (N_3915,N_1240,N_1189);
nor U3916 (N_3916,N_984,N_240);
nor U3917 (N_3917,N_1509,N_667);
or U3918 (N_3918,N_1425,N_125);
xor U3919 (N_3919,N_1496,N_1042);
nand U3920 (N_3920,N_223,N_138);
and U3921 (N_3921,N_437,N_700);
or U3922 (N_3922,N_1870,N_1838);
nor U3923 (N_3923,N_1003,N_546);
and U3924 (N_3924,N_587,N_347);
or U3925 (N_3925,N_1472,N_1774);
or U3926 (N_3926,N_677,N_595);
nand U3927 (N_3927,N_786,N_694);
and U3928 (N_3928,N_376,N_1991);
nor U3929 (N_3929,N_457,N_474);
nand U3930 (N_3930,N_230,N_678);
nand U3931 (N_3931,N_671,N_1208);
and U3932 (N_3932,N_285,N_375);
and U3933 (N_3933,N_1878,N_1216);
nand U3934 (N_3934,N_1883,N_86);
nor U3935 (N_3935,N_909,N_1757);
and U3936 (N_3936,N_1284,N_55);
xor U3937 (N_3937,N_1827,N_1446);
and U3938 (N_3938,N_578,N_1373);
or U3939 (N_3939,N_1217,N_258);
nor U3940 (N_3940,N_707,N_1932);
nand U3941 (N_3941,N_1687,N_1025);
and U3942 (N_3942,N_445,N_1665);
nor U3943 (N_3943,N_1601,N_320);
or U3944 (N_3944,N_1177,N_1607);
and U3945 (N_3945,N_1570,N_1043);
nor U3946 (N_3946,N_1234,N_1282);
nand U3947 (N_3947,N_1985,N_261);
nand U3948 (N_3948,N_1536,N_1558);
nand U3949 (N_3949,N_1036,N_485);
nor U3950 (N_3950,N_1653,N_1396);
nand U3951 (N_3951,N_298,N_1616);
nand U3952 (N_3952,N_1417,N_1869);
nor U3953 (N_3953,N_569,N_1079);
nor U3954 (N_3954,N_861,N_1895);
nand U3955 (N_3955,N_1825,N_655);
nor U3956 (N_3956,N_623,N_642);
xnor U3957 (N_3957,N_1068,N_305);
and U3958 (N_3958,N_802,N_1627);
nor U3959 (N_3959,N_987,N_885);
nand U3960 (N_3960,N_481,N_951);
nor U3961 (N_3961,N_1343,N_1113);
or U3962 (N_3962,N_1396,N_233);
nand U3963 (N_3963,N_215,N_1563);
and U3964 (N_3964,N_1487,N_1102);
nand U3965 (N_3965,N_1912,N_243);
nor U3966 (N_3966,N_1202,N_62);
or U3967 (N_3967,N_577,N_677);
nor U3968 (N_3968,N_1631,N_1609);
nor U3969 (N_3969,N_1526,N_120);
nand U3970 (N_3970,N_1057,N_1263);
and U3971 (N_3971,N_1875,N_743);
nand U3972 (N_3972,N_588,N_1982);
nor U3973 (N_3973,N_1174,N_223);
nor U3974 (N_3974,N_1513,N_416);
nand U3975 (N_3975,N_459,N_1125);
nand U3976 (N_3976,N_1542,N_1926);
or U3977 (N_3977,N_801,N_1474);
or U3978 (N_3978,N_1840,N_1991);
or U3979 (N_3979,N_901,N_935);
or U3980 (N_3980,N_779,N_1227);
and U3981 (N_3981,N_785,N_329);
or U3982 (N_3982,N_171,N_653);
or U3983 (N_3983,N_85,N_1678);
or U3984 (N_3984,N_632,N_587);
and U3985 (N_3985,N_1720,N_819);
nand U3986 (N_3986,N_451,N_1879);
and U3987 (N_3987,N_853,N_6);
nand U3988 (N_3988,N_888,N_1989);
or U3989 (N_3989,N_68,N_1724);
or U3990 (N_3990,N_1681,N_1797);
nand U3991 (N_3991,N_1048,N_1484);
or U3992 (N_3992,N_565,N_1613);
nor U3993 (N_3993,N_1464,N_274);
xor U3994 (N_3994,N_959,N_1982);
nor U3995 (N_3995,N_996,N_1034);
or U3996 (N_3996,N_1509,N_1118);
and U3997 (N_3997,N_1731,N_1215);
and U3998 (N_3998,N_908,N_1570);
or U3999 (N_3999,N_1535,N_1200);
nor U4000 (N_4000,N_3736,N_2189);
and U4001 (N_4001,N_2388,N_2790);
or U4002 (N_4002,N_3607,N_3130);
and U4003 (N_4003,N_2580,N_3680);
nand U4004 (N_4004,N_3242,N_2700);
and U4005 (N_4005,N_3351,N_2239);
and U4006 (N_4006,N_2227,N_2394);
nand U4007 (N_4007,N_3688,N_2714);
nor U4008 (N_4008,N_3784,N_3210);
and U4009 (N_4009,N_2565,N_3203);
or U4010 (N_4010,N_2750,N_3415);
nor U4011 (N_4011,N_3987,N_3327);
and U4012 (N_4012,N_3797,N_2999);
nand U4013 (N_4013,N_3893,N_2611);
and U4014 (N_4014,N_3950,N_2271);
or U4015 (N_4015,N_3246,N_2931);
nand U4016 (N_4016,N_2797,N_3709);
or U4017 (N_4017,N_2936,N_3883);
nor U4018 (N_4018,N_3886,N_2282);
or U4019 (N_4019,N_2658,N_3409);
or U4020 (N_4020,N_3953,N_3573);
and U4021 (N_4021,N_3978,N_2806);
or U4022 (N_4022,N_2799,N_3759);
nor U4023 (N_4023,N_3827,N_2769);
nor U4024 (N_4024,N_2829,N_2038);
or U4025 (N_4025,N_3534,N_3667);
nand U4026 (N_4026,N_3560,N_3606);
and U4027 (N_4027,N_2109,N_3374);
nand U4028 (N_4028,N_3931,N_2910);
nand U4029 (N_4029,N_2642,N_3404);
and U4030 (N_4030,N_2377,N_2311);
or U4031 (N_4031,N_2013,N_2967);
or U4032 (N_4032,N_3512,N_2672);
nor U4033 (N_4033,N_2869,N_3273);
nand U4034 (N_4034,N_3479,N_2043);
nand U4035 (N_4035,N_3822,N_2637);
and U4036 (N_4036,N_3553,N_3773);
and U4037 (N_4037,N_2175,N_3439);
and U4038 (N_4038,N_2649,N_2246);
nand U4039 (N_4039,N_2097,N_3287);
or U4040 (N_4040,N_2322,N_3256);
nor U4041 (N_4041,N_2346,N_3644);
nand U4042 (N_4042,N_3328,N_2119);
and U4043 (N_4043,N_3285,N_2005);
nor U4044 (N_4044,N_2582,N_3348);
and U4045 (N_4045,N_2634,N_2857);
nor U4046 (N_4046,N_3690,N_2655);
nor U4047 (N_4047,N_2809,N_2051);
nand U4048 (N_4048,N_2635,N_3569);
or U4049 (N_4049,N_3991,N_3433);
or U4050 (N_4050,N_3831,N_3320);
or U4051 (N_4051,N_3166,N_3755);
xor U4052 (N_4052,N_2904,N_2029);
and U4053 (N_4053,N_3032,N_2478);
and U4054 (N_4054,N_3686,N_2052);
nor U4055 (N_4055,N_2661,N_3758);
nor U4056 (N_4056,N_2357,N_3159);
nand U4057 (N_4057,N_2135,N_2512);
nand U4058 (N_4058,N_2289,N_2507);
nand U4059 (N_4059,N_2952,N_3856);
nor U4060 (N_4060,N_3395,N_3664);
or U4061 (N_4061,N_3340,N_3187);
nor U4062 (N_4062,N_2780,N_2674);
and U4063 (N_4063,N_2131,N_3948);
nand U4064 (N_4064,N_3006,N_2505);
and U4065 (N_4065,N_3448,N_2845);
nand U4066 (N_4066,N_2868,N_2430);
or U4067 (N_4067,N_3113,N_3005);
xor U4068 (N_4068,N_2179,N_2313);
nor U4069 (N_4069,N_2240,N_3862);
and U4070 (N_4070,N_2954,N_2222);
or U4071 (N_4071,N_3168,N_3460);
or U4072 (N_4072,N_3097,N_2354);
nor U4073 (N_4073,N_2698,N_3476);
or U4074 (N_4074,N_2784,N_2224);
nor U4075 (N_4075,N_3334,N_2735);
and U4076 (N_4076,N_3143,N_2673);
or U4077 (N_4077,N_3115,N_2390);
nand U4078 (N_4078,N_2939,N_3588);
or U4079 (N_4079,N_3417,N_2612);
and U4080 (N_4080,N_3945,N_2822);
nor U4081 (N_4081,N_3347,N_2881);
nor U4082 (N_4082,N_3385,N_2807);
nand U4083 (N_4083,N_2746,N_2641);
nor U4084 (N_4084,N_2073,N_2048);
or U4085 (N_4085,N_3807,N_3997);
nor U4086 (N_4086,N_2379,N_2712);
nand U4087 (N_4087,N_3453,N_2410);
or U4088 (N_4088,N_3576,N_2256);
and U4089 (N_4089,N_3592,N_2614);
nor U4090 (N_4090,N_3302,N_2166);
nor U4091 (N_4091,N_3048,N_3177);
nor U4092 (N_4092,N_2849,N_3154);
or U4093 (N_4093,N_2848,N_2552);
or U4094 (N_4094,N_3316,N_3330);
and U4095 (N_4095,N_3444,N_2278);
nand U4096 (N_4096,N_2703,N_3280);
or U4097 (N_4097,N_3610,N_3936);
and U4098 (N_4098,N_2428,N_2560);
and U4099 (N_4099,N_3603,N_3739);
nor U4100 (N_4100,N_2751,N_3258);
nand U4101 (N_4101,N_3493,N_3207);
or U4102 (N_4102,N_2104,N_2555);
or U4103 (N_4103,N_3894,N_2697);
nor U4104 (N_4104,N_2440,N_2009);
nor U4105 (N_4105,N_2820,N_2081);
or U4106 (N_4106,N_3707,N_2479);
or U4107 (N_4107,N_2449,N_3407);
nor U4108 (N_4108,N_3671,N_2362);
nor U4109 (N_4109,N_2206,N_3411);
or U4110 (N_4110,N_3632,N_3891);
nor U4111 (N_4111,N_3572,N_3400);
nand U4112 (N_4112,N_2453,N_2473);
nor U4113 (N_4113,N_3537,N_3823);
and U4114 (N_4114,N_3298,N_2685);
and U4115 (N_4115,N_2671,N_3440);
nor U4116 (N_4116,N_2554,N_3383);
nand U4117 (N_4117,N_3977,N_2546);
and U4118 (N_4118,N_2221,N_2125);
nand U4119 (N_4119,N_2965,N_3257);
nand U4120 (N_4120,N_3146,N_3757);
xor U4121 (N_4121,N_3546,N_3173);
or U4122 (N_4122,N_3416,N_2195);
and U4123 (N_4123,N_3854,N_2934);
or U4124 (N_4124,N_3148,N_3656);
or U4125 (N_4125,N_2046,N_2963);
and U4126 (N_4126,N_2991,N_3367);
nor U4127 (N_4127,N_3234,N_3182);
nor U4128 (N_4128,N_3729,N_2188);
or U4129 (N_4129,N_2485,N_3767);
and U4130 (N_4130,N_2108,N_3089);
and U4131 (N_4131,N_2676,N_2501);
nor U4132 (N_4132,N_2587,N_3092);
and U4133 (N_4133,N_3542,N_3410);
xor U4134 (N_4134,N_3034,N_2396);
and U4135 (N_4135,N_3908,N_3994);
nor U4136 (N_4136,N_2884,N_2747);
or U4137 (N_4137,N_2948,N_2475);
and U4138 (N_4138,N_3728,N_2645);
nor U4139 (N_4139,N_2850,N_3888);
nand U4140 (N_4140,N_2979,N_2129);
or U4141 (N_4141,N_3446,N_2815);
or U4142 (N_4142,N_3910,N_3284);
nand U4143 (N_4143,N_3892,N_2306);
xor U4144 (N_4144,N_2260,N_2011);
or U4145 (N_4145,N_2987,N_2941);
nor U4146 (N_4146,N_2412,N_2359);
or U4147 (N_4147,N_3749,N_2007);
and U4148 (N_4148,N_3804,N_3585);
and U4149 (N_4149,N_2481,N_3941);
and U4150 (N_4150,N_2981,N_3625);
nor U4151 (N_4151,N_3397,N_3300);
and U4152 (N_4152,N_3035,N_3150);
nand U4153 (N_4153,N_3106,N_3084);
nand U4154 (N_4154,N_2696,N_3488);
nor U4155 (N_4155,N_2464,N_2360);
or U4156 (N_4156,N_3080,N_3341);
and U4157 (N_4157,N_2927,N_2036);
or U4158 (N_4158,N_3007,N_3845);
or U4159 (N_4159,N_3108,N_2576);
nor U4160 (N_4160,N_2826,N_3740);
and U4161 (N_4161,N_3754,N_3838);
and U4162 (N_4162,N_3485,N_3060);
nand U4163 (N_4163,N_2732,N_3288);
nor U4164 (N_4164,N_2945,N_2436);
or U4165 (N_4165,N_3053,N_2032);
or U4166 (N_4166,N_2782,N_3903);
or U4167 (N_4167,N_3171,N_2235);
or U4168 (N_4168,N_2207,N_2586);
or U4169 (N_4169,N_3579,N_3121);
or U4170 (N_4170,N_2897,N_2093);
nand U4171 (N_4171,N_3536,N_3543);
or U4172 (N_4172,N_3186,N_2403);
or U4173 (N_4173,N_3408,N_2583);
nand U4174 (N_4174,N_2792,N_2037);
or U4175 (N_4175,N_2626,N_2717);
nand U4176 (N_4176,N_3642,N_3565);
nor U4177 (N_4177,N_3323,N_3215);
or U4178 (N_4178,N_2974,N_2124);
or U4179 (N_4179,N_2111,N_3355);
nor U4180 (N_4180,N_2681,N_3122);
nor U4181 (N_4181,N_3583,N_3024);
and U4182 (N_4182,N_2964,N_3547);
nand U4183 (N_4183,N_3081,N_3029);
nor U4184 (N_4184,N_3541,N_3277);
or U4185 (N_4185,N_3332,N_2662);
and U4186 (N_4186,N_3129,N_2808);
or U4187 (N_4187,N_3630,N_3079);
nor U4188 (N_4188,N_3466,N_2935);
and U4189 (N_4189,N_2392,N_2250);
or U4190 (N_4190,N_2123,N_3737);
and U4191 (N_4191,N_3524,N_3612);
or U4192 (N_4192,N_3529,N_2343);
or U4193 (N_4193,N_3343,N_3456);
or U4194 (N_4194,N_2255,N_3353);
or U4195 (N_4195,N_3509,N_3235);
nor U4196 (N_4196,N_3577,N_2245);
nor U4197 (N_4197,N_3438,N_3001);
nand U4198 (N_4198,N_2272,N_3363);
and U4199 (N_4199,N_2647,N_3361);
and U4200 (N_4200,N_2439,N_2352);
or U4201 (N_4201,N_2061,N_2744);
or U4202 (N_4202,N_2261,N_3458);
nand U4203 (N_4203,N_2937,N_3748);
and U4204 (N_4204,N_3684,N_2856);
nor U4205 (N_4205,N_3155,N_2940);
or U4206 (N_4206,N_3056,N_2349);
nand U4207 (N_4207,N_3939,N_3628);
nor U4208 (N_4208,N_3430,N_2543);
xor U4209 (N_4209,N_3745,N_2077);
or U4210 (N_4210,N_2985,N_3696);
or U4211 (N_4211,N_2545,N_2327);
and U4212 (N_4212,N_3490,N_2173);
nand U4213 (N_4213,N_2572,N_3682);
nand U4214 (N_4214,N_3641,N_3627);
and U4215 (N_4215,N_3314,N_3131);
or U4216 (N_4216,N_3788,N_2364);
nand U4217 (N_4217,N_3907,N_3000);
or U4218 (N_4218,N_2708,N_2702);
or U4219 (N_4219,N_3996,N_3850);
and U4220 (N_4220,N_2607,N_2372);
nand U4221 (N_4221,N_2281,N_2600);
and U4222 (N_4222,N_2140,N_2026);
and U4223 (N_4223,N_2774,N_2438);
nor U4224 (N_4224,N_3066,N_3836);
or U4225 (N_4225,N_3550,N_3508);
and U4226 (N_4226,N_2183,N_3959);
nand U4227 (N_4227,N_3801,N_3023);
nand U4228 (N_4228,N_2098,N_3137);
nor U4229 (N_4229,N_2068,N_3643);
nand U4230 (N_4230,N_3818,N_2793);
or U4231 (N_4231,N_3071,N_2315);
or U4232 (N_4232,N_3010,N_2157);
and U4233 (N_4233,N_3153,N_2594);
and U4234 (N_4234,N_3750,N_3431);
or U4235 (N_4235,N_3412,N_3070);
and U4236 (N_4236,N_3255,N_3114);
and U4237 (N_4237,N_2992,N_3392);
nor U4238 (N_4238,N_2960,N_3058);
or U4239 (N_4239,N_2204,N_3702);
and U4240 (N_4240,N_3999,N_3601);
nor U4241 (N_4241,N_3955,N_2251);
and U4242 (N_4242,N_2273,N_3318);
or U4243 (N_4243,N_2853,N_3321);
nand U4244 (N_4244,N_3160,N_2742);
or U4245 (N_4245,N_2729,N_3180);
nand U4246 (N_4246,N_3449,N_2921);
and U4247 (N_4247,N_2876,N_3076);
nand U4248 (N_4248,N_3350,N_3008);
and U4249 (N_4249,N_3175,N_2065);
and U4250 (N_4250,N_3502,N_3935);
or U4251 (N_4251,N_3083,N_3515);
or U4252 (N_4252,N_3816,N_3915);
nor U4253 (N_4253,N_2724,N_3631);
nand U4254 (N_4254,N_2942,N_2561);
nor U4255 (N_4255,N_3720,N_2603);
nor U4256 (N_4256,N_2928,N_3598);
or U4257 (N_4257,N_3857,N_2181);
nor U4258 (N_4258,N_2151,N_2519);
nand U4259 (N_4259,N_2898,N_3527);
and U4260 (N_4260,N_3518,N_3800);
nor U4261 (N_4261,N_2615,N_2092);
nor U4262 (N_4262,N_3659,N_3711);
nand U4263 (N_4263,N_2573,N_3937);
nor U4264 (N_4264,N_2492,N_3370);
and U4265 (N_4265,N_2923,N_2006);
or U4266 (N_4266,N_3026,N_3824);
nand U4267 (N_4267,N_3120,N_3971);
or U4268 (N_4268,N_2280,N_3510);
nand U4269 (N_4269,N_3764,N_2341);
nor U4270 (N_4270,N_3605,N_3934);
and U4271 (N_4271,N_2651,N_2844);
nor U4272 (N_4272,N_3184,N_3881);
and U4273 (N_4273,N_3099,N_2066);
nand U4274 (N_4274,N_2926,N_2514);
nor U4275 (N_4275,N_3609,N_2630);
and U4276 (N_4276,N_3983,N_3790);
nor U4277 (N_4277,N_2414,N_2145);
nor U4278 (N_4278,N_3296,N_2544);
and U4279 (N_4279,N_2989,N_2961);
nor U4280 (N_4280,N_3544,N_2162);
and U4281 (N_4281,N_2091,N_2667);
or U4282 (N_4282,N_3311,N_3140);
nand U4283 (N_4283,N_3507,N_3435);
nand U4284 (N_4284,N_2197,N_2000);
nor U4285 (N_4285,N_2798,N_2956);
and U4286 (N_4286,N_3900,N_2513);
or U4287 (N_4287,N_3687,N_3091);
and U4288 (N_4288,N_2663,N_2938);
and U4289 (N_4289,N_3722,N_2500);
or U4290 (N_4290,N_3861,N_3779);
nand U4291 (N_4291,N_2818,N_2616);
nand U4292 (N_4292,N_2033,N_3645);
and U4293 (N_4293,N_2382,N_3283);
nor U4294 (N_4294,N_3634,N_3497);
and U4295 (N_4295,N_3062,N_2053);
nor U4296 (N_4296,N_2613,N_2644);
nor U4297 (N_4297,N_2621,N_3357);
nand U4298 (N_4298,N_2292,N_2802);
and U4299 (N_4299,N_2027,N_2929);
nand U4300 (N_4300,N_3346,N_2319);
nand U4301 (N_4301,N_2393,N_2693);
xor U4302 (N_4302,N_3768,N_2760);
or U4303 (N_4303,N_3743,N_2977);
nor U4304 (N_4304,N_3443,N_3434);
nor U4305 (N_4305,N_2553,N_3128);
or U4306 (N_4306,N_2932,N_3895);
xnor U4307 (N_4307,N_2060,N_2020);
or U4308 (N_4308,N_3982,N_2435);
and U4309 (N_4309,N_2075,N_3653);
or U4310 (N_4310,N_2577,N_2851);
or U4311 (N_4311,N_3832,N_3679);
nor U4312 (N_4312,N_3303,N_2759);
nand U4313 (N_4313,N_3904,N_3414);
nor U4314 (N_4314,N_2623,N_2370);
or U4315 (N_4315,N_3020,N_3102);
nand U4316 (N_4316,N_2833,N_2827);
and U4317 (N_4317,N_3331,N_2527);
nand U4318 (N_4318,N_3317,N_2276);
nand U4319 (N_4319,N_2269,N_3078);
nor U4320 (N_4320,N_2537,N_2070);
or U4321 (N_4321,N_3014,N_2683);
nand U4322 (N_4322,N_2540,N_3563);
nor U4323 (N_4323,N_2950,N_3243);
nor U4324 (N_4324,N_2437,N_2959);
xnor U4325 (N_4325,N_2592,N_3013);
or U4326 (N_4326,N_3176,N_3803);
nor U4327 (N_4327,N_3551,N_2012);
or U4328 (N_4328,N_2886,N_2628);
and U4329 (N_4329,N_3594,N_2168);
and U4330 (N_4330,N_3947,N_3738);
nor U4331 (N_4331,N_2363,N_3238);
and U4332 (N_4332,N_3962,N_2010);
nor U4333 (N_4333,N_3360,N_2733);
or U4334 (N_4334,N_3698,N_2834);
or U4335 (N_4335,N_3517,N_2779);
nand U4336 (N_4336,N_2566,N_3830);
nor U4337 (N_4337,N_2726,N_3525);
and U4338 (N_4338,N_3972,N_2983);
nand U4339 (N_4339,N_3730,N_3792);
nand U4340 (N_4340,N_3295,N_3566);
or U4341 (N_4341,N_2116,N_3125);
nand U4342 (N_4342,N_2721,N_3199);
or U4343 (N_4343,N_3635,N_3090);
and U4344 (N_4344,N_2633,N_2190);
and U4345 (N_4345,N_2254,N_3202);
nand U4346 (N_4346,N_2230,N_2300);
nor U4347 (N_4347,N_3470,N_2223);
nor U4348 (N_4348,N_2218,N_3617);
nor U4349 (N_4349,N_3725,N_2409);
and U4350 (N_4350,N_2597,N_2174);
nand U4351 (N_4351,N_2090,N_3858);
nand U4352 (N_4352,N_2194,N_2045);
nor U4353 (N_4353,N_2099,N_3611);
or U4354 (N_4354,N_2214,N_3806);
or U4355 (N_4355,N_3855,N_3398);
nand U4356 (N_4356,N_2665,N_3269);
nor U4357 (N_4357,N_3956,N_3533);
xor U4358 (N_4358,N_2397,N_2244);
or U4359 (N_4359,N_3897,N_3652);
and U4360 (N_4360,N_2903,N_3123);
nor U4361 (N_4361,N_2212,N_2550);
nor U4362 (N_4362,N_2398,N_2297);
and U4363 (N_4363,N_3085,N_2973);
or U4364 (N_4364,N_3511,N_2533);
or U4365 (N_4365,N_2598,N_3194);
or U4366 (N_4366,N_2639,N_2529);
nor U4367 (N_4367,N_2406,N_3031);
nor U4368 (N_4368,N_2199,N_3335);
or U4369 (N_4369,N_3865,N_2944);
or U4370 (N_4370,N_2911,N_3169);
or U4371 (N_4371,N_2266,N_2459);
nand U4372 (N_4372,N_2494,N_3401);
and U4373 (N_4373,N_2812,N_2907);
nand U4374 (N_4374,N_3785,N_2407);
and U4375 (N_4375,N_3463,N_3494);
or U4376 (N_4376,N_2925,N_2765);
or U4377 (N_4377,N_3993,N_3217);
nand U4378 (N_4378,N_3821,N_3747);
or U4379 (N_4379,N_3437,N_2990);
nor U4380 (N_4380,N_2024,N_2542);
and U4381 (N_4381,N_3152,N_2395);
nor U4382 (N_4382,N_3228,N_2842);
or U4383 (N_4383,N_3798,N_2448);
nor U4384 (N_4384,N_2770,N_2581);
and U4385 (N_4385,N_2618,N_2520);
xor U4386 (N_4386,N_3778,N_2231);
or U4387 (N_4387,N_3386,N_3864);
or U4388 (N_4388,N_2404,N_2722);
and U4389 (N_4389,N_3232,N_2787);
nand U4390 (N_4390,N_2862,N_2314);
nor U4391 (N_4391,N_3593,N_2515);
nand U4392 (N_4392,N_2917,N_2740);
nor U4393 (N_4393,N_2356,N_2627);
and U4394 (N_4394,N_2495,N_3045);
nor U4395 (N_4395,N_2686,N_3112);
nor U4396 (N_4396,N_3751,N_2933);
and U4397 (N_4397,N_2426,N_3923);
nand U4398 (N_4398,N_2483,N_3849);
and U4399 (N_4399,N_2378,N_2203);
and U4400 (N_4400,N_2776,N_2585);
nand U4401 (N_4401,N_2386,N_2972);
nand U4402 (N_4402,N_3636,N_2433);
and U4403 (N_4403,N_2677,N_3828);
nand U4404 (N_4404,N_2772,N_3811);
nor U4405 (N_4405,N_2984,N_3796);
nand U4406 (N_4406,N_3265,N_2804);
and U4407 (N_4407,N_2795,N_3866);
and U4408 (N_4408,N_2215,N_3116);
nor U4409 (N_4409,N_3036,N_3561);
nand U4410 (N_4410,N_3842,N_2914);
nor U4411 (N_4411,N_3942,N_3837);
nand U4412 (N_4412,N_3629,N_3809);
nand U4413 (N_4413,N_3943,N_3963);
and U4414 (N_4414,N_2283,N_2087);
nor U4415 (N_4415,N_2988,N_2838);
or U4416 (N_4416,N_2518,N_2083);
nand U4417 (N_4417,N_3513,N_3608);
or U4418 (N_4418,N_2723,N_2718);
and U4419 (N_4419,N_2699,N_2267);
nor U4420 (N_4420,N_2472,N_2423);
or U4421 (N_4421,N_3322,N_2208);
nand U4422 (N_4422,N_2293,N_2536);
nor U4423 (N_4423,N_3793,N_3038);
or U4424 (N_4424,N_2568,N_3156);
nand U4425 (N_4425,N_2835,N_2526);
or U4426 (N_4426,N_2317,N_2457);
or U4427 (N_4427,N_2042,N_2657);
or U4428 (N_4428,N_2872,N_2730);
nand U4429 (N_4429,N_2896,N_2885);
and U4430 (N_4430,N_2801,N_2569);
nand U4431 (N_4431,N_2640,N_2069);
nor U4432 (N_4432,N_2427,N_3072);
and U4433 (N_4433,N_3851,N_2148);
nand U4434 (N_4434,N_2114,N_3003);
and U4435 (N_4435,N_3528,N_3491);
or U4436 (N_4436,N_3147,N_3464);
or U4437 (N_4437,N_3700,N_3174);
or U4438 (N_4438,N_2588,N_2172);
nand U4439 (N_4439,N_2447,N_2556);
nor U4440 (N_4440,N_3640,N_2517);
nand U4441 (N_4441,N_2996,N_2969);
nand U4442 (N_4442,N_2901,N_3069);
and U4443 (N_4443,N_3613,N_2285);
and U4444 (N_4444,N_3602,N_3872);
nand U4445 (N_4445,N_2737,N_3967);
nor U4446 (N_4446,N_2843,N_2480);
and U4447 (N_4447,N_2496,N_2811);
and U4448 (N_4448,N_3961,N_3789);
nand U4449 (N_4449,N_2079,N_2694);
nor U4450 (N_4450,N_3812,N_3587);
or U4451 (N_4451,N_3467,N_3393);
or U4452 (N_4452,N_3744,N_2134);
nor U4453 (N_4453,N_2847,N_2710);
xor U4454 (N_4454,N_3135,N_2023);
or U4455 (N_4455,N_2225,N_2351);
nand U4456 (N_4456,N_3964,N_3368);
and U4457 (N_4457,N_3372,N_2755);
and U4458 (N_4458,N_2490,N_3658);
and U4459 (N_4459,N_3521,N_2080);
nor U4460 (N_4460,N_3815,N_2211);
and U4461 (N_4461,N_3245,N_2022);
nand U4462 (N_4462,N_3701,N_2205);
or U4463 (N_4463,N_3204,N_2365);
and U4464 (N_4464,N_2373,N_3447);
and U4465 (N_4465,N_2191,N_3107);
nor U4466 (N_4466,N_2817,N_3377);
nand U4467 (N_4467,N_2946,N_2187);
nand U4468 (N_4468,N_3814,N_2014);
nand U4469 (N_4469,N_2487,N_3930);
nor U4470 (N_4470,N_3042,N_2017);
or U4471 (N_4471,N_2321,N_3500);
and U4472 (N_4472,N_3012,N_2691);
and U4473 (N_4473,N_2304,N_2652);
or U4474 (N_4474,N_3059,N_3519);
and U4475 (N_4475,N_2268,N_3380);
nor U4476 (N_4476,N_3158,N_2263);
or U4477 (N_4477,N_2711,N_2830);
or U4478 (N_4478,N_2736,N_2727);
and U4479 (N_4479,N_2656,N_2978);
and U4480 (N_4480,N_3041,N_2995);
or U4481 (N_4481,N_2380,N_2763);
xor U4482 (N_4482,N_2753,N_2400);
nor U4483 (N_4483,N_3132,N_3254);
nor U4484 (N_4484,N_2219,N_3639);
nor U4485 (N_4485,N_2170,N_2286);
or U4486 (N_4486,N_2059,N_2345);
or U4487 (N_4487,N_2078,N_3799);
nor U4488 (N_4488,N_3713,N_2589);
or U4489 (N_4489,N_2442,N_3867);
nor U4490 (N_4490,N_2361,N_3018);
nand U4491 (N_4491,N_3905,N_3044);
or U4492 (N_4492,N_3111,N_2624);
nand U4493 (N_4493,N_3365,N_2220);
or U4494 (N_4494,N_2270,N_2810);
xor U4495 (N_4495,N_2692,N_2559);
nor U4496 (N_4496,N_3802,N_3462);
nor U4497 (N_4497,N_3669,N_3819);
or U4498 (N_4498,N_3164,N_2713);
and U4499 (N_4499,N_2082,N_2035);
or U4500 (N_4500,N_3216,N_2466);
and U4501 (N_4501,N_3196,N_3649);
or U4502 (N_4502,N_3988,N_2295);
and U4503 (N_4503,N_2058,N_3535);
or U4504 (N_4504,N_3301,N_2031);
nor U4505 (N_4505,N_2084,N_2957);
and U4506 (N_4506,N_3279,N_2429);
nand U4507 (N_4507,N_2159,N_2424);
or U4508 (N_4508,N_3478,N_2675);
nand U4509 (N_4509,N_3957,N_3826);
or U4510 (N_4510,N_2154,N_2333);
and U4511 (N_4511,N_3271,N_2894);
nand U4512 (N_4512,N_2547,N_3002);
nand U4513 (N_4513,N_3661,N_2452);
or U4514 (N_4514,N_2121,N_3165);
and U4515 (N_4515,N_3324,N_3455);
nor U4516 (N_4516,N_2654,N_3557);
nor U4517 (N_4517,N_3817,N_2525);
nand U4518 (N_4518,N_3200,N_2855);
nor U4519 (N_4519,N_2874,N_3692);
or U4520 (N_4520,N_3637,N_3752);
nand U4521 (N_4521,N_2535,N_3151);
nor U4522 (N_4522,N_3902,N_2086);
and U4523 (N_4523,N_2030,N_2320);
nand U4524 (N_4524,N_2096,N_3025);
or U4525 (N_4525,N_2906,N_3161);
nor U4526 (N_4526,N_3672,N_3666);
nand U4527 (N_4527,N_2277,N_3336);
nor U4528 (N_4528,N_2136,N_3325);
nand U4529 (N_4529,N_2307,N_3782);
or U4530 (N_4530,N_2336,N_2101);
nor U4531 (N_4531,N_3213,N_3840);
and U4532 (N_4532,N_3975,N_2584);
xnor U4533 (N_4533,N_2137,N_3791);
or U4534 (N_4534,N_2670,N_3532);
nand U4535 (N_4535,N_2767,N_2242);
nor U4536 (N_4536,N_3540,N_2854);
and U4537 (N_4537,N_2326,N_2593);
and U4538 (N_4538,N_2126,N_3595);
and U4539 (N_4539,N_3844,N_3932);
or U4540 (N_4540,N_2132,N_3675);
nor U4541 (N_4541,N_3694,N_2381);
nand U4542 (N_4542,N_2421,N_3847);
nor U4543 (N_4543,N_2019,N_3017);
and U4544 (N_4544,N_3241,N_3871);
nand U4545 (N_4545,N_2103,N_2039);
nand U4546 (N_4546,N_3052,N_2625);
nand U4547 (N_4547,N_3226,N_3580);
nand U4548 (N_4548,N_2775,N_2766);
nand U4549 (N_4549,N_2332,N_2389);
nor U4550 (N_4550,N_3495,N_3712);
and U4551 (N_4551,N_3074,N_3960);
or U4552 (N_4552,N_2143,N_3061);
or U4553 (N_4553,N_2880,N_2570);
or U4554 (N_4554,N_3911,N_3364);
nand U4555 (N_4555,N_2419,N_2484);
or U4556 (N_4556,N_3506,N_3139);
xnor U4557 (N_4557,N_3291,N_2368);
nor U4558 (N_4558,N_2358,N_2888);
and U4559 (N_4559,N_2241,N_3138);
and U4560 (N_4560,N_2761,N_3781);
nand U4561 (N_4561,N_2653,N_3275);
or U4562 (N_4562,N_3413,N_3037);
nand U4563 (N_4563,N_2968,N_2041);
nand U4564 (N_4564,N_2557,N_2422);
nor U4565 (N_4565,N_2579,N_2434);
nor U4566 (N_4566,N_3646,N_2117);
or U4567 (N_4567,N_2416,N_2506);
or U4568 (N_4568,N_3589,N_3925);
or U4569 (N_4569,N_2476,N_3095);
or U4570 (N_4570,N_2110,N_3918);
or U4571 (N_4571,N_3538,N_3604);
and U4572 (N_4572,N_3501,N_3382);
nand U4573 (N_4573,N_3086,N_2279);
or U4574 (N_4574,N_3820,N_2474);
nor U4575 (N_4575,N_2163,N_3338);
or U4576 (N_4576,N_2201,N_2548);
nand U4577 (N_4577,N_3489,N_3616);
nand U4578 (N_4578,N_3869,N_3756);
or U4579 (N_4579,N_2344,N_3266);
nor U4580 (N_4580,N_3763,N_2161);
and U4581 (N_4581,N_3304,N_2768);
nand U4582 (N_4582,N_3727,N_3887);
or U4583 (N_4583,N_2509,N_3292);
nand U4584 (N_4584,N_2180,N_2376);
nand U4585 (N_4585,N_2617,N_3211);
nand U4586 (N_4586,N_2538,N_3685);
and U4587 (N_4587,N_3545,N_3775);
or U4588 (N_4588,N_3033,N_3568);
nor U4589 (N_4589,N_3333,N_2980);
nor U4590 (N_4590,N_2503,N_2156);
nand U4591 (N_4591,N_2113,N_3621);
nand U4592 (N_4592,N_2445,N_3101);
nor U4593 (N_4593,N_2497,N_3654);
nand U4594 (N_4594,N_3884,N_3890);
nor U4595 (N_4595,N_2040,N_2836);
nor U4596 (N_4596,N_3552,N_3668);
or U4597 (N_4597,N_3267,N_2420);
or U4598 (N_4598,N_2067,N_2706);
nand U4599 (N_4599,N_2057,N_3208);
nand U4600 (N_4600,N_3496,N_3620);
and U4601 (N_4601,N_3929,N_2047);
nor U4602 (N_4602,N_3825,N_2660);
and U4603 (N_4603,N_3795,N_2142);
nand U4604 (N_4604,N_2831,N_2678);
and U4605 (N_4605,N_3626,N_2725);
or U4606 (N_4606,N_3846,N_2824);
nor U4607 (N_4607,N_3976,N_3676);
nand U4608 (N_4608,N_3452,N_2028);
and U4609 (N_4609,N_3379,N_2102);
or U4610 (N_4610,N_3229,N_2467);
or U4611 (N_4611,N_3191,N_3833);
xor U4612 (N_4612,N_2741,N_2105);
xor U4613 (N_4613,N_3261,N_3420);
and U4614 (N_4614,N_3970,N_3721);
nand U4615 (N_4615,N_3969,N_3848);
nor U4616 (N_4616,N_3263,N_2088);
and U4617 (N_4617,N_2659,N_2469);
and U4618 (N_4618,N_3906,N_3530);
nand U4619 (N_4619,N_3181,N_3946);
or U4620 (N_4620,N_2858,N_2353);
nor U4621 (N_4621,N_2499,N_2127);
or U4622 (N_4622,N_3875,N_3293);
or U4623 (N_4623,N_3157,N_3623);
nand U4624 (N_4624,N_3657,N_3933);
nor U4625 (N_4625,N_3526,N_2604);
or U4626 (N_4626,N_2158,N_2294);
nor U4627 (N_4627,N_2924,N_3162);
or U4628 (N_4628,N_3928,N_3220);
or U4629 (N_4629,N_3040,N_3098);
nand U4630 (N_4630,N_3787,N_3233);
nand U4631 (N_4631,N_3468,N_2383);
or U4632 (N_4632,N_2828,N_2334);
nand U4633 (N_4633,N_3170,N_2669);
and U4634 (N_4634,N_2076,N_2541);
xor U4635 (N_4635,N_2912,N_3985);
or U4636 (N_4636,N_3896,N_3475);
nor U4637 (N_4637,N_2825,N_3968);
nor U4638 (N_4638,N_2595,N_3735);
or U4639 (N_4639,N_2122,N_3704);
nand U4640 (N_4640,N_2551,N_2044);
nor U4641 (N_4641,N_3877,N_3870);
or U4642 (N_4642,N_3600,N_3674);
or U4643 (N_4643,N_2636,N_2018);
and U4644 (N_4644,N_2909,N_2892);
and U4645 (N_4645,N_2549,N_2176);
nor U4646 (N_4646,N_3183,N_2491);
and U4647 (N_4647,N_2015,N_2387);
nand U4648 (N_4648,N_3222,N_2149);
nand U4649 (N_4649,N_2308,N_3581);
or U4650 (N_4650,N_2528,N_2994);
nand U4651 (N_4651,N_3651,N_3599);
nor U4652 (N_4652,N_3885,N_2680);
or U4653 (N_4653,N_2144,N_3922);
or U4654 (N_4654,N_2302,N_2578);
and U4655 (N_4655,N_2993,N_2878);
or U4656 (N_4656,N_2860,N_2200);
or U4657 (N_4657,N_2034,N_3761);
nand U4658 (N_4658,N_3426,N_3352);
and U4659 (N_4659,N_2182,N_3880);
xnor U4660 (N_4660,N_3909,N_3424);
or U4661 (N_4661,N_3919,N_3039);
nor U4662 (N_4662,N_2465,N_2210);
or U4663 (N_4663,N_2873,N_3133);
or U4664 (N_4664,N_3484,N_2922);
or U4665 (N_4665,N_2301,N_3231);
nand U4666 (N_4666,N_3859,N_3486);
and U4667 (N_4667,N_3559,N_3236);
nand U4668 (N_4668,N_2682,N_3944);
or U4669 (N_4669,N_3852,N_3376);
or U4670 (N_4670,N_3315,N_3305);
or U4671 (N_4671,N_2335,N_2839);
and U4672 (N_4672,N_3703,N_2488);
nand U4673 (N_4673,N_3899,N_2608);
or U4674 (N_4674,N_3055,N_2146);
nand U4675 (N_4675,N_2498,N_3973);
xor U4676 (N_4676,N_3144,N_2619);
nor U4677 (N_4677,N_3118,N_2508);
or U4678 (N_4678,N_3951,N_3454);
and U4679 (N_4679,N_3004,N_2728);
and U4680 (N_4680,N_3432,N_3021);
nor U4681 (N_4681,N_3843,N_3198);
nor U4682 (N_4682,N_2516,N_3381);
nand U4683 (N_4683,N_2716,N_3223);
and U4684 (N_4684,N_3655,N_3556);
or U4685 (N_4685,N_2169,N_3369);
or U4686 (N_4686,N_3927,N_3124);
or U4687 (N_4687,N_3399,N_2130);
nand U4688 (N_4688,N_3638,N_3860);
and U4689 (N_4689,N_3492,N_3185);
or U4690 (N_4690,N_3057,N_2754);
or U4691 (N_4691,N_2879,N_3665);
and U4692 (N_4692,N_3584,N_3068);
or U4693 (N_4693,N_2916,N_3878);
nor U4694 (N_4694,N_2415,N_3723);
and U4695 (N_4695,N_3765,N_3558);
and U4696 (N_4696,N_2021,N_3442);
nor U4697 (N_4697,N_2863,N_3681);
and U4698 (N_4698,N_2253,N_2316);
or U4699 (N_4699,N_2562,N_2895);
and U4700 (N_4700,N_2259,N_3221);
or U4701 (N_4701,N_2599,N_2919);
or U4702 (N_4702,N_3047,N_3248);
nand U4703 (N_4703,N_2369,N_3126);
and U4704 (N_4704,N_2511,N_2620);
nor U4705 (N_4705,N_3389,N_3774);
or U4706 (N_4706,N_2997,N_3349);
or U4707 (N_4707,N_2287,N_2323);
nand U4708 (N_4708,N_2745,N_2743);
or U4709 (N_4709,N_2638,N_2877);
nand U4710 (N_4710,N_3731,N_3974);
nand U4711 (N_4711,N_2152,N_3249);
and U4712 (N_4712,N_2739,N_3926);
or U4713 (N_4713,N_2213,N_2720);
nand U4714 (N_4714,N_2522,N_3306);
nor U4715 (N_4715,N_2609,N_2375);
nand U4716 (N_4716,N_2558,N_2049);
or U4717 (N_4717,N_3049,N_3345);
and U4718 (N_4718,N_2574,N_2451);
or U4719 (N_4719,N_3718,N_2056);
nor U4720 (N_4720,N_2785,N_3366);
and U4721 (N_4721,N_3618,N_3205);
nand U4722 (N_4722,N_3282,N_3436);
and U4723 (N_4723,N_3197,N_3054);
nand U4724 (N_4724,N_2258,N_2531);
or U4725 (N_4725,N_3046,N_3178);
nor U4726 (N_4726,N_3762,N_3050);
nand U4727 (N_4727,N_3274,N_2288);
or U4728 (N_4728,N_3808,N_2679);
or U4729 (N_4729,N_2003,N_2913);
nand U4730 (N_4730,N_2690,N_3251);
nand U4731 (N_4731,N_2477,N_2402);
or U4732 (N_4732,N_3660,N_3482);
and U4733 (N_4733,N_3247,N_2975);
nor U4734 (N_4734,N_2062,N_3384);
nor U4735 (N_4735,N_3766,N_3067);
and U4736 (N_4736,N_2186,N_3477);
or U4737 (N_4737,N_2871,N_3127);
nand U4738 (N_4738,N_2112,N_2217);
and U4739 (N_4739,N_3461,N_3917);
and U4740 (N_4740,N_3805,N_3777);
and U4741 (N_4741,N_3590,N_3418);
or U4742 (N_4742,N_2971,N_2882);
or U4743 (N_4743,N_2813,N_2237);
and U4744 (N_4744,N_2821,N_3691);
or U4745 (N_4745,N_3949,N_3104);
nand U4746 (N_4746,N_2337,N_2752);
xor U4747 (N_4747,N_3746,N_2339);
or U4748 (N_4748,N_2859,N_2366);
and U4749 (N_4749,N_3297,N_3405);
and U4750 (N_4750,N_3149,N_2107);
or U4751 (N_4751,N_3998,N_2050);
or U4752 (N_4752,N_2832,N_2530);
and U4753 (N_4753,N_2756,N_2106);
and U4754 (N_4754,N_3281,N_3624);
and U4755 (N_4755,N_2226,N_3406);
or U4756 (N_4756,N_2425,N_3504);
or U4757 (N_4757,N_3043,N_2631);
nor U4758 (N_4758,N_3662,N_2303);
nand U4759 (N_4759,N_2982,N_3834);
nor U4760 (N_4760,N_2800,N_2791);
or U4761 (N_4761,N_2184,N_3724);
nor U4762 (N_4762,N_2016,N_3480);
nor U4763 (N_4763,N_3531,N_3192);
and U4764 (N_4764,N_2115,N_2299);
xnor U4765 (N_4765,N_3073,N_2705);
or U4766 (N_4766,N_2100,N_3965);
nand U4767 (N_4767,N_3783,N_2918);
and U4768 (N_4768,N_2689,N_2601);
nor U4769 (N_4769,N_3853,N_2953);
and U4770 (N_4770,N_2296,N_3276);
and U4771 (N_4771,N_2072,N_2958);
nor U4772 (N_4772,N_3428,N_2202);
and U4773 (N_4773,N_2632,N_3310);
nand U4774 (N_4774,N_3342,N_2318);
nor U4775 (N_4775,N_2470,N_2865);
xor U4776 (N_4776,N_2391,N_2905);
and U4777 (N_4777,N_3879,N_3189);
and U4778 (N_4778,N_2325,N_3209);
and U4779 (N_4779,N_3075,N_3979);
or U4780 (N_4780,N_2861,N_2232);
or U4781 (N_4781,N_2902,N_2629);
or U4782 (N_4782,N_2709,N_3179);
or U4783 (N_4783,N_2605,N_2330);
nand U4784 (N_4784,N_2648,N_2171);
and U4785 (N_4785,N_2852,N_3571);
or U4786 (N_4786,N_3483,N_2610);
nand U4787 (N_4787,N_3394,N_3117);
or U4788 (N_4788,N_3319,N_2408);
or U4789 (N_4789,N_3574,N_2695);
and U4790 (N_4790,N_3813,N_2837);
nand U4791 (N_4791,N_3780,N_2177);
and U4792 (N_4792,N_2155,N_2883);
and U4793 (N_4793,N_3505,N_3995);
or U4794 (N_4794,N_3451,N_3921);
nor U4795 (N_4795,N_3190,N_3145);
or U4796 (N_4796,N_2731,N_3954);
nor U4797 (N_4797,N_2329,N_3278);
and U4798 (N_4798,N_3786,N_3992);
and U4799 (N_4799,N_3516,N_2970);
or U4800 (N_4800,N_2262,N_3699);
nor U4801 (N_4801,N_3633,N_2915);
nor U4802 (N_4802,N_2489,N_3354);
nand U4803 (N_4803,N_3422,N_3695);
nor U4804 (N_4804,N_3966,N_3219);
and U4805 (N_4805,N_2534,N_2216);
nor U4806 (N_4806,N_2778,N_3980);
nor U4807 (N_4807,N_3378,N_2371);
nor U4808 (N_4808,N_2650,N_3390);
and U4809 (N_4809,N_2738,N_2462);
nand U4810 (N_4810,N_2704,N_3810);
nand U4811 (N_4811,N_2247,N_2340);
or U4812 (N_4812,N_3403,N_2668);
nor U4813 (N_4813,N_3308,N_3465);
or U4814 (N_4814,N_2458,N_2120);
nor U4815 (N_4815,N_2265,N_2064);
nor U4816 (N_4816,N_2823,N_3253);
and U4817 (N_4817,N_3920,N_3615);
nand U4818 (N_4818,N_2900,N_2094);
nand U4819 (N_4819,N_2521,N_2955);
or U4820 (N_4820,N_2054,N_2748);
nor U4821 (N_4821,N_3421,N_3195);
and U4822 (N_4822,N_3371,N_2193);
nor U4823 (N_4823,N_2328,N_2417);
or U4824 (N_4824,N_3272,N_3100);
nor U4825 (N_4825,N_3110,N_3958);
and U4826 (N_4826,N_3741,N_3981);
and U4827 (N_4827,N_3423,N_3647);
nor U4828 (N_4828,N_3770,N_2455);
or U4829 (N_4829,N_2405,N_3224);
and U4830 (N_4830,N_3841,N_3710);
nand U4831 (N_4831,N_2486,N_3163);
and U4832 (N_4832,N_3717,N_3167);
or U4833 (N_4833,N_2870,N_3549);
and U4834 (N_4834,N_3670,N_3705);
or U4835 (N_4835,N_3225,N_2891);
nand U4836 (N_4836,N_2456,N_2875);
and U4837 (N_4837,N_2128,N_2074);
nand U4838 (N_4838,N_3916,N_2264);
nor U4839 (N_4839,N_3260,N_3359);
and U4840 (N_4840,N_3022,N_3650);
and U4841 (N_4841,N_3239,N_3912);
or U4842 (N_4842,N_2715,N_3402);
nand U4843 (N_4843,N_2866,N_2893);
and U4844 (N_4844,N_3459,N_3706);
and U4845 (N_4845,N_3760,N_3063);
nor U4846 (N_4846,N_2841,N_2147);
and U4847 (N_4847,N_3873,N_2342);
nor U4848 (N_4848,N_2133,N_3214);
nor U4849 (N_4849,N_2930,N_3141);
nor U4850 (N_4850,N_3889,N_3622);
and U4851 (N_4851,N_2643,N_2719);
or U4852 (N_4852,N_2291,N_3769);
nor U4853 (N_4853,N_3562,N_3868);
xnor U4854 (N_4854,N_3425,N_3259);
nand U4855 (N_4855,N_3450,N_2071);
or U4856 (N_4856,N_3733,N_2493);
nor U4857 (N_4857,N_3082,N_2867);
nor U4858 (N_4858,N_3678,N_2482);
nand U4859 (N_4859,N_2463,N_3498);
and U4860 (N_4860,N_2450,N_3742);
xnor U4861 (N_4861,N_3387,N_2348);
or U4862 (N_4862,N_2411,N_3874);
nand U4863 (N_4863,N_2840,N_2257);
nand U4864 (N_4864,N_2947,N_3719);
and U4865 (N_4865,N_3523,N_2539);
or U4866 (N_4866,N_3499,N_2966);
and U4867 (N_4867,N_3753,N_2602);
nand U4868 (N_4868,N_2532,N_3474);
or U4869 (N_4869,N_2846,N_3514);
nor U4870 (N_4870,N_2085,N_3570);
nand U4871 (N_4871,N_3520,N_3193);
nor U4872 (N_4872,N_2164,N_3294);
nand U4873 (N_4873,N_3309,N_2331);
or U4874 (N_4874,N_2819,N_3564);
and U4875 (N_4875,N_2228,N_3206);
and U4876 (N_4876,N_3109,N_2758);
and U4877 (N_4877,N_2347,N_3250);
or U4878 (N_4878,N_2471,N_3375);
nor U4879 (N_4879,N_3142,N_2814);
nor U4880 (N_4880,N_2803,N_3136);
or U4881 (N_4881,N_2773,N_2684);
nor U4882 (N_4882,N_3555,N_3028);
nand U4883 (N_4883,N_3901,N_3714);
nand U4884 (N_4884,N_3429,N_3481);
and U4885 (N_4885,N_3286,N_2749);
and U4886 (N_4886,N_3548,N_2305);
nand U4887 (N_4887,N_2764,N_2781);
and U4888 (N_4888,N_2777,N_3237);
or U4889 (N_4889,N_3105,N_2460);
nor U4890 (N_4890,N_3009,N_2002);
and U4891 (N_4891,N_2160,N_2095);
nand U4892 (N_4892,N_3794,N_2324);
nor U4893 (N_4893,N_3689,N_2510);
nand U4894 (N_4894,N_2198,N_2788);
nor U4895 (N_4895,N_2384,N_2504);
or U4896 (N_4896,N_3016,N_3619);
and U4897 (N_4897,N_3591,N_3356);
and U4898 (N_4898,N_2138,N_2350);
nor U4899 (N_4899,N_2233,N_3776);
nand U4900 (N_4900,N_2908,N_3270);
and U4901 (N_4901,N_2118,N_2355);
or U4902 (N_4902,N_2762,N_3172);
nand U4903 (N_4903,N_2274,N_3673);
and U4904 (N_4904,N_3472,N_2252);
and U4905 (N_4905,N_3596,N_3663);
nand U4906 (N_4906,N_3445,N_2943);
or U4907 (N_4907,N_3388,N_3575);
xor U4908 (N_4908,N_2986,N_2236);
and U4909 (N_4909,N_3441,N_2374);
or U4910 (N_4910,N_3715,N_3597);
or U4911 (N_4911,N_3227,N_3188);
or U4912 (N_4912,N_2796,N_3539);
or U4913 (N_4913,N_2243,N_3567);
or U4914 (N_4914,N_3391,N_3471);
nor U4915 (N_4915,N_2150,N_2590);
and U4916 (N_4916,N_3984,N_2783);
or U4917 (N_4917,N_3771,N_2004);
and U4918 (N_4918,N_2771,N_3093);
or U4919 (N_4919,N_2571,N_3027);
or U4920 (N_4920,N_2687,N_2290);
nor U4921 (N_4921,N_3487,N_2139);
nand U4922 (N_4922,N_3586,N_2298);
nor U4923 (N_4923,N_3924,N_2338);
nor U4924 (N_4924,N_3362,N_3262);
nor U4925 (N_4925,N_3011,N_3734);
or U4926 (N_4926,N_3307,N_2141);
or U4927 (N_4927,N_2887,N_2399);
or U4928 (N_4928,N_2431,N_3473);
nor U4929 (N_4929,N_2564,N_2454);
or U4930 (N_4930,N_2889,N_2310);
nand U4931 (N_4931,N_3863,N_2444);
nand U4932 (N_4932,N_3134,N_3289);
nor U4933 (N_4933,N_3503,N_2025);
and U4934 (N_4934,N_2523,N_3064);
or U4935 (N_4935,N_2786,N_2196);
nand U4936 (N_4936,N_2563,N_3290);
or U4937 (N_4937,N_2234,N_3952);
and U4938 (N_4938,N_3252,N_2502);
or U4939 (N_4939,N_2284,N_3337);
or U4940 (N_4940,N_2622,N_3065);
nor U4941 (N_4941,N_3582,N_2275);
nor U4942 (N_4942,N_2646,N_2167);
and U4943 (N_4943,N_3358,N_3457);
nor U4944 (N_4944,N_2432,N_3299);
or U4945 (N_4945,N_2249,N_2312);
nor U4946 (N_4946,N_2229,N_3940);
or U4947 (N_4947,N_3989,N_3077);
xnor U4948 (N_4948,N_3326,N_2591);
nand U4949 (N_4949,N_3419,N_2606);
nor U4950 (N_4950,N_3201,N_3051);
xnor U4951 (N_4951,N_3373,N_3264);
nor U4952 (N_4952,N_2248,N_3522);
nand U4953 (N_4953,N_3648,N_2920);
or U4954 (N_4954,N_2309,N_3268);
xnor U4955 (N_4955,N_2757,N_2178);
and U4956 (N_4956,N_3019,N_2575);
nand U4957 (N_4957,N_2089,N_2976);
or U4958 (N_4958,N_2998,N_2794);
xor U4959 (N_4959,N_3087,N_2192);
nor U4960 (N_4960,N_2899,N_3914);
nand U4961 (N_4961,N_3339,N_2001);
nand U4962 (N_4962,N_2524,N_2567);
and U4963 (N_4963,N_3835,N_2238);
or U4964 (N_4964,N_2816,N_2413);
and U4965 (N_4965,N_3772,N_3683);
or U4966 (N_4966,N_3839,N_3469);
or U4967 (N_4967,N_3578,N_2441);
nor U4968 (N_4968,N_3726,N_3030);
and U4969 (N_4969,N_3230,N_3829);
or U4970 (N_4970,N_3103,N_2367);
or U4971 (N_4971,N_2153,N_2185);
or U4972 (N_4972,N_3986,N_2864);
or U4973 (N_4973,N_3938,N_3015);
or U4974 (N_4974,N_3244,N_3882);
nand U4975 (N_4975,N_3913,N_3312);
and U4976 (N_4976,N_3732,N_2734);
and U4977 (N_4977,N_2701,N_3693);
nor U4978 (N_4978,N_2707,N_3708);
or U4979 (N_4979,N_3990,N_2789);
nor U4980 (N_4980,N_2209,N_2951);
xor U4981 (N_4981,N_3554,N_2165);
or U4982 (N_4982,N_2962,N_2055);
or U4983 (N_4983,N_3697,N_3313);
nor U4984 (N_4984,N_3218,N_3898);
nand U4985 (N_4985,N_2418,N_3344);
and U4986 (N_4986,N_3677,N_2805);
or U4987 (N_4987,N_2443,N_3329);
and U4988 (N_4988,N_2666,N_2063);
nor U4989 (N_4989,N_3119,N_2446);
and U4990 (N_4990,N_2385,N_3094);
or U4991 (N_4991,N_3716,N_2461);
xnor U4992 (N_4992,N_3096,N_2401);
nor U4993 (N_4993,N_3396,N_2890);
xor U4994 (N_4994,N_3240,N_3614);
and U4995 (N_4995,N_2468,N_2949);
and U4996 (N_4996,N_3212,N_2664);
nand U4997 (N_4997,N_3876,N_2596);
or U4998 (N_4998,N_3088,N_2688);
or U4999 (N_4999,N_3427,N_2008);
nor U5000 (N_5000,N_2220,N_2227);
nand U5001 (N_5001,N_3467,N_2820);
and U5002 (N_5002,N_3602,N_3269);
and U5003 (N_5003,N_3052,N_3876);
nor U5004 (N_5004,N_2540,N_3555);
nand U5005 (N_5005,N_2839,N_3295);
and U5006 (N_5006,N_3881,N_2352);
xnor U5007 (N_5007,N_2396,N_3728);
or U5008 (N_5008,N_2796,N_2936);
or U5009 (N_5009,N_2611,N_3106);
or U5010 (N_5010,N_2155,N_2544);
nor U5011 (N_5011,N_3310,N_2561);
nand U5012 (N_5012,N_2085,N_2781);
and U5013 (N_5013,N_3361,N_3789);
and U5014 (N_5014,N_2975,N_2664);
nand U5015 (N_5015,N_3941,N_2186);
or U5016 (N_5016,N_3145,N_3151);
nand U5017 (N_5017,N_3819,N_3289);
or U5018 (N_5018,N_2649,N_2461);
and U5019 (N_5019,N_3139,N_2752);
and U5020 (N_5020,N_2941,N_3334);
xor U5021 (N_5021,N_3174,N_3539);
nor U5022 (N_5022,N_2696,N_2643);
nor U5023 (N_5023,N_3188,N_3893);
nand U5024 (N_5024,N_3731,N_2362);
nand U5025 (N_5025,N_2339,N_3590);
nand U5026 (N_5026,N_3587,N_3323);
nor U5027 (N_5027,N_2220,N_2038);
nor U5028 (N_5028,N_3279,N_3407);
nor U5029 (N_5029,N_3073,N_2681);
or U5030 (N_5030,N_2682,N_2485);
or U5031 (N_5031,N_2117,N_3103);
or U5032 (N_5032,N_3632,N_3387);
nand U5033 (N_5033,N_3443,N_2636);
and U5034 (N_5034,N_2341,N_2021);
nor U5035 (N_5035,N_2236,N_3797);
and U5036 (N_5036,N_3578,N_3221);
or U5037 (N_5037,N_2541,N_3853);
or U5038 (N_5038,N_2605,N_3281);
or U5039 (N_5039,N_2556,N_3824);
nor U5040 (N_5040,N_2979,N_3393);
or U5041 (N_5041,N_3365,N_2483);
or U5042 (N_5042,N_3506,N_3145);
nor U5043 (N_5043,N_2322,N_2332);
and U5044 (N_5044,N_3194,N_3361);
or U5045 (N_5045,N_3861,N_2386);
or U5046 (N_5046,N_3412,N_3313);
nor U5047 (N_5047,N_2043,N_3237);
nor U5048 (N_5048,N_2790,N_2890);
and U5049 (N_5049,N_2784,N_3439);
nor U5050 (N_5050,N_2378,N_2416);
nand U5051 (N_5051,N_2061,N_2738);
or U5052 (N_5052,N_3741,N_3881);
and U5053 (N_5053,N_3307,N_2440);
and U5054 (N_5054,N_2657,N_2952);
or U5055 (N_5055,N_2876,N_3019);
nor U5056 (N_5056,N_2804,N_3038);
nand U5057 (N_5057,N_3686,N_3937);
nand U5058 (N_5058,N_2902,N_2586);
nor U5059 (N_5059,N_3100,N_3217);
and U5060 (N_5060,N_3180,N_3116);
nand U5061 (N_5061,N_3451,N_3855);
or U5062 (N_5062,N_3909,N_2864);
nand U5063 (N_5063,N_2973,N_2845);
or U5064 (N_5064,N_2002,N_3577);
and U5065 (N_5065,N_2950,N_2444);
or U5066 (N_5066,N_3267,N_3570);
and U5067 (N_5067,N_2377,N_3396);
nand U5068 (N_5068,N_2775,N_2691);
or U5069 (N_5069,N_2425,N_2181);
and U5070 (N_5070,N_3715,N_3104);
or U5071 (N_5071,N_2647,N_2611);
nand U5072 (N_5072,N_3882,N_3066);
nor U5073 (N_5073,N_3953,N_3778);
nor U5074 (N_5074,N_3908,N_3006);
or U5075 (N_5075,N_3695,N_3770);
nand U5076 (N_5076,N_3915,N_2265);
and U5077 (N_5077,N_3556,N_2161);
or U5078 (N_5078,N_3575,N_3026);
nor U5079 (N_5079,N_2257,N_2850);
nor U5080 (N_5080,N_2145,N_2085);
nor U5081 (N_5081,N_3411,N_2854);
and U5082 (N_5082,N_2325,N_3989);
nor U5083 (N_5083,N_3628,N_2801);
or U5084 (N_5084,N_3109,N_3504);
or U5085 (N_5085,N_2631,N_3508);
nand U5086 (N_5086,N_3424,N_2826);
and U5087 (N_5087,N_3606,N_2453);
nand U5088 (N_5088,N_3484,N_2397);
and U5089 (N_5089,N_2316,N_2464);
and U5090 (N_5090,N_3819,N_3848);
or U5091 (N_5091,N_3856,N_2433);
and U5092 (N_5092,N_2024,N_3096);
nand U5093 (N_5093,N_2621,N_3209);
xor U5094 (N_5094,N_3023,N_3124);
nand U5095 (N_5095,N_2870,N_3579);
and U5096 (N_5096,N_2905,N_2535);
or U5097 (N_5097,N_3811,N_2649);
and U5098 (N_5098,N_3240,N_2890);
nand U5099 (N_5099,N_2708,N_2798);
xnor U5100 (N_5100,N_3990,N_2483);
nand U5101 (N_5101,N_2278,N_3359);
and U5102 (N_5102,N_3110,N_3947);
nand U5103 (N_5103,N_2424,N_3081);
and U5104 (N_5104,N_2042,N_2260);
nand U5105 (N_5105,N_2613,N_2318);
xor U5106 (N_5106,N_2296,N_2369);
nor U5107 (N_5107,N_2172,N_2161);
nand U5108 (N_5108,N_3213,N_2636);
and U5109 (N_5109,N_3212,N_2224);
and U5110 (N_5110,N_3151,N_3081);
or U5111 (N_5111,N_2628,N_2212);
or U5112 (N_5112,N_3973,N_3004);
xor U5113 (N_5113,N_3202,N_2170);
nand U5114 (N_5114,N_3372,N_2236);
nand U5115 (N_5115,N_3479,N_2251);
or U5116 (N_5116,N_3267,N_2641);
and U5117 (N_5117,N_3091,N_2399);
and U5118 (N_5118,N_3406,N_3747);
nand U5119 (N_5119,N_2139,N_2360);
nand U5120 (N_5120,N_2591,N_3460);
nor U5121 (N_5121,N_2568,N_3947);
nand U5122 (N_5122,N_3298,N_3798);
or U5123 (N_5123,N_3219,N_3639);
or U5124 (N_5124,N_3790,N_3565);
nor U5125 (N_5125,N_2071,N_3007);
nand U5126 (N_5126,N_2637,N_3734);
xnor U5127 (N_5127,N_3470,N_3481);
or U5128 (N_5128,N_3955,N_3289);
and U5129 (N_5129,N_2266,N_3753);
or U5130 (N_5130,N_2477,N_2879);
and U5131 (N_5131,N_2598,N_3354);
xor U5132 (N_5132,N_2389,N_2384);
or U5133 (N_5133,N_3005,N_2140);
or U5134 (N_5134,N_3634,N_3486);
nor U5135 (N_5135,N_3235,N_2039);
and U5136 (N_5136,N_2213,N_3355);
or U5137 (N_5137,N_3122,N_2170);
nand U5138 (N_5138,N_3205,N_3727);
nand U5139 (N_5139,N_2869,N_3910);
nand U5140 (N_5140,N_3810,N_2156);
or U5141 (N_5141,N_2009,N_3144);
and U5142 (N_5142,N_2281,N_2194);
and U5143 (N_5143,N_3084,N_3053);
nand U5144 (N_5144,N_3427,N_2223);
or U5145 (N_5145,N_2273,N_3947);
nor U5146 (N_5146,N_2053,N_2979);
nor U5147 (N_5147,N_3376,N_3079);
or U5148 (N_5148,N_2992,N_3186);
and U5149 (N_5149,N_3973,N_2373);
nand U5150 (N_5150,N_2673,N_2097);
and U5151 (N_5151,N_2644,N_2970);
and U5152 (N_5152,N_2816,N_2612);
nor U5153 (N_5153,N_2747,N_2328);
nand U5154 (N_5154,N_3719,N_2228);
nand U5155 (N_5155,N_3750,N_2467);
nand U5156 (N_5156,N_3229,N_2767);
or U5157 (N_5157,N_2158,N_3515);
xnor U5158 (N_5158,N_3148,N_3655);
nand U5159 (N_5159,N_3381,N_2264);
nor U5160 (N_5160,N_3669,N_2444);
and U5161 (N_5161,N_2057,N_3179);
xor U5162 (N_5162,N_2570,N_3417);
and U5163 (N_5163,N_3472,N_3614);
xnor U5164 (N_5164,N_2731,N_3421);
and U5165 (N_5165,N_2970,N_3573);
or U5166 (N_5166,N_3019,N_3580);
nand U5167 (N_5167,N_3155,N_2768);
nand U5168 (N_5168,N_2042,N_3258);
nor U5169 (N_5169,N_3507,N_3132);
or U5170 (N_5170,N_3296,N_2335);
or U5171 (N_5171,N_2854,N_3634);
and U5172 (N_5172,N_2266,N_2457);
or U5173 (N_5173,N_3273,N_2021);
and U5174 (N_5174,N_2996,N_3926);
and U5175 (N_5175,N_2681,N_2214);
nand U5176 (N_5176,N_2318,N_3604);
nor U5177 (N_5177,N_2166,N_2479);
nand U5178 (N_5178,N_3741,N_3036);
or U5179 (N_5179,N_2933,N_2299);
and U5180 (N_5180,N_2801,N_2808);
or U5181 (N_5181,N_2475,N_2404);
nand U5182 (N_5182,N_2180,N_2657);
or U5183 (N_5183,N_2373,N_3153);
nand U5184 (N_5184,N_2654,N_2591);
or U5185 (N_5185,N_3089,N_2452);
and U5186 (N_5186,N_2429,N_3049);
nand U5187 (N_5187,N_2640,N_2565);
nor U5188 (N_5188,N_2700,N_2519);
nand U5189 (N_5189,N_2019,N_3572);
and U5190 (N_5190,N_3267,N_2785);
or U5191 (N_5191,N_3584,N_3771);
or U5192 (N_5192,N_2754,N_3625);
nor U5193 (N_5193,N_2849,N_2868);
or U5194 (N_5194,N_2861,N_3785);
nand U5195 (N_5195,N_3624,N_3342);
nor U5196 (N_5196,N_3548,N_3857);
nor U5197 (N_5197,N_3224,N_3411);
and U5198 (N_5198,N_2286,N_2178);
nand U5199 (N_5199,N_2273,N_2920);
nand U5200 (N_5200,N_3584,N_2552);
nand U5201 (N_5201,N_3459,N_3022);
nor U5202 (N_5202,N_2683,N_3922);
and U5203 (N_5203,N_2439,N_3233);
nor U5204 (N_5204,N_3757,N_2395);
and U5205 (N_5205,N_2995,N_3316);
or U5206 (N_5206,N_2152,N_3287);
nand U5207 (N_5207,N_2148,N_3874);
and U5208 (N_5208,N_3903,N_3598);
nand U5209 (N_5209,N_2245,N_2523);
nor U5210 (N_5210,N_2433,N_3433);
and U5211 (N_5211,N_3544,N_2441);
and U5212 (N_5212,N_2113,N_3035);
or U5213 (N_5213,N_2563,N_2119);
or U5214 (N_5214,N_2924,N_2815);
nand U5215 (N_5215,N_3236,N_3729);
nand U5216 (N_5216,N_3773,N_3939);
nand U5217 (N_5217,N_3629,N_2842);
or U5218 (N_5218,N_3965,N_3407);
and U5219 (N_5219,N_2347,N_2208);
nand U5220 (N_5220,N_3262,N_3492);
and U5221 (N_5221,N_2928,N_2423);
or U5222 (N_5222,N_2117,N_2915);
xor U5223 (N_5223,N_3613,N_2799);
nor U5224 (N_5224,N_3918,N_2258);
and U5225 (N_5225,N_3525,N_3462);
and U5226 (N_5226,N_2065,N_2853);
nand U5227 (N_5227,N_2904,N_3377);
nor U5228 (N_5228,N_3029,N_2271);
nor U5229 (N_5229,N_2988,N_2362);
or U5230 (N_5230,N_3526,N_2925);
nand U5231 (N_5231,N_2678,N_3740);
nand U5232 (N_5232,N_3645,N_3836);
nand U5233 (N_5233,N_3490,N_2784);
nand U5234 (N_5234,N_2185,N_2172);
or U5235 (N_5235,N_3837,N_3367);
and U5236 (N_5236,N_3536,N_3333);
nor U5237 (N_5237,N_3976,N_2864);
and U5238 (N_5238,N_3640,N_2630);
nand U5239 (N_5239,N_2042,N_2611);
nand U5240 (N_5240,N_3747,N_2421);
nand U5241 (N_5241,N_3934,N_3751);
nor U5242 (N_5242,N_3391,N_3957);
nand U5243 (N_5243,N_2775,N_3048);
nor U5244 (N_5244,N_2886,N_3836);
and U5245 (N_5245,N_3262,N_2623);
nand U5246 (N_5246,N_2969,N_3893);
xnor U5247 (N_5247,N_2531,N_2650);
nand U5248 (N_5248,N_3710,N_3651);
nand U5249 (N_5249,N_2231,N_2016);
nand U5250 (N_5250,N_2622,N_3861);
nand U5251 (N_5251,N_3655,N_3177);
or U5252 (N_5252,N_2390,N_3943);
nand U5253 (N_5253,N_3048,N_3624);
nor U5254 (N_5254,N_3624,N_3446);
nand U5255 (N_5255,N_3097,N_2940);
or U5256 (N_5256,N_3345,N_3659);
nor U5257 (N_5257,N_3364,N_2098);
or U5258 (N_5258,N_2163,N_2237);
and U5259 (N_5259,N_3654,N_2783);
nor U5260 (N_5260,N_3077,N_3885);
nor U5261 (N_5261,N_3746,N_3483);
nor U5262 (N_5262,N_3816,N_3579);
nand U5263 (N_5263,N_3513,N_3941);
xor U5264 (N_5264,N_3951,N_2061);
nor U5265 (N_5265,N_3430,N_3426);
nand U5266 (N_5266,N_2883,N_2190);
and U5267 (N_5267,N_3240,N_3497);
or U5268 (N_5268,N_3332,N_3092);
nand U5269 (N_5269,N_3399,N_2167);
and U5270 (N_5270,N_3995,N_2658);
and U5271 (N_5271,N_3057,N_3132);
nor U5272 (N_5272,N_3686,N_2427);
or U5273 (N_5273,N_3239,N_2502);
nor U5274 (N_5274,N_3053,N_2100);
xor U5275 (N_5275,N_2700,N_3617);
nand U5276 (N_5276,N_2993,N_2986);
or U5277 (N_5277,N_2329,N_3954);
nand U5278 (N_5278,N_2797,N_3436);
nand U5279 (N_5279,N_3923,N_2621);
nand U5280 (N_5280,N_3389,N_3692);
or U5281 (N_5281,N_3737,N_2244);
and U5282 (N_5282,N_2024,N_3007);
nor U5283 (N_5283,N_3958,N_2605);
nor U5284 (N_5284,N_3201,N_2658);
or U5285 (N_5285,N_3905,N_3652);
and U5286 (N_5286,N_2454,N_3643);
and U5287 (N_5287,N_2005,N_2322);
xor U5288 (N_5288,N_3894,N_2871);
or U5289 (N_5289,N_2328,N_3134);
or U5290 (N_5290,N_2900,N_3234);
nor U5291 (N_5291,N_3857,N_3492);
and U5292 (N_5292,N_2196,N_3574);
nand U5293 (N_5293,N_3028,N_3416);
nand U5294 (N_5294,N_3397,N_2008);
nor U5295 (N_5295,N_2200,N_3726);
and U5296 (N_5296,N_3586,N_2654);
nand U5297 (N_5297,N_2048,N_3301);
nand U5298 (N_5298,N_3554,N_2916);
xnor U5299 (N_5299,N_3289,N_3455);
nand U5300 (N_5300,N_3948,N_2807);
or U5301 (N_5301,N_3952,N_3645);
nand U5302 (N_5302,N_2224,N_2536);
or U5303 (N_5303,N_2799,N_3128);
nand U5304 (N_5304,N_3687,N_2179);
and U5305 (N_5305,N_3382,N_3591);
nand U5306 (N_5306,N_3841,N_3329);
and U5307 (N_5307,N_2182,N_3976);
nor U5308 (N_5308,N_3071,N_2438);
or U5309 (N_5309,N_2170,N_3571);
or U5310 (N_5310,N_3043,N_2954);
nand U5311 (N_5311,N_2086,N_2703);
nand U5312 (N_5312,N_2333,N_2955);
and U5313 (N_5313,N_3387,N_3312);
nor U5314 (N_5314,N_3235,N_2187);
nand U5315 (N_5315,N_3740,N_3963);
nor U5316 (N_5316,N_3310,N_3468);
nor U5317 (N_5317,N_2672,N_3029);
or U5318 (N_5318,N_3410,N_2490);
and U5319 (N_5319,N_3416,N_2171);
nor U5320 (N_5320,N_3694,N_2099);
nor U5321 (N_5321,N_3077,N_3440);
nor U5322 (N_5322,N_2594,N_2290);
and U5323 (N_5323,N_3704,N_2556);
nand U5324 (N_5324,N_2636,N_2779);
and U5325 (N_5325,N_2396,N_3799);
or U5326 (N_5326,N_3336,N_2684);
or U5327 (N_5327,N_3017,N_2031);
or U5328 (N_5328,N_2159,N_3627);
nand U5329 (N_5329,N_2315,N_2404);
nor U5330 (N_5330,N_2548,N_2949);
and U5331 (N_5331,N_2945,N_3366);
and U5332 (N_5332,N_3341,N_2238);
xnor U5333 (N_5333,N_2786,N_3430);
nor U5334 (N_5334,N_3479,N_2520);
and U5335 (N_5335,N_2788,N_3352);
or U5336 (N_5336,N_3282,N_3474);
and U5337 (N_5337,N_2242,N_2541);
or U5338 (N_5338,N_3713,N_2174);
nand U5339 (N_5339,N_3851,N_3442);
or U5340 (N_5340,N_2793,N_2037);
nand U5341 (N_5341,N_2667,N_3042);
nand U5342 (N_5342,N_3182,N_3924);
nand U5343 (N_5343,N_2682,N_3953);
and U5344 (N_5344,N_2915,N_3728);
xnor U5345 (N_5345,N_2416,N_3649);
nor U5346 (N_5346,N_2600,N_2493);
and U5347 (N_5347,N_3637,N_3917);
or U5348 (N_5348,N_2278,N_3150);
or U5349 (N_5349,N_3303,N_3683);
nand U5350 (N_5350,N_2285,N_3482);
or U5351 (N_5351,N_3704,N_3401);
or U5352 (N_5352,N_2715,N_2485);
and U5353 (N_5353,N_2390,N_3778);
nor U5354 (N_5354,N_2138,N_3004);
nor U5355 (N_5355,N_3230,N_3890);
nor U5356 (N_5356,N_3987,N_3925);
nor U5357 (N_5357,N_2914,N_3578);
and U5358 (N_5358,N_3692,N_2133);
nor U5359 (N_5359,N_3083,N_3796);
nand U5360 (N_5360,N_3998,N_3231);
nor U5361 (N_5361,N_2902,N_3629);
or U5362 (N_5362,N_3083,N_3107);
xor U5363 (N_5363,N_2835,N_2944);
and U5364 (N_5364,N_2930,N_3889);
nor U5365 (N_5365,N_2379,N_3140);
nor U5366 (N_5366,N_2629,N_2260);
nor U5367 (N_5367,N_2439,N_3004);
nand U5368 (N_5368,N_2604,N_2025);
and U5369 (N_5369,N_3059,N_3419);
and U5370 (N_5370,N_2520,N_3922);
nand U5371 (N_5371,N_2551,N_2761);
and U5372 (N_5372,N_3500,N_2039);
nor U5373 (N_5373,N_3307,N_3292);
nand U5374 (N_5374,N_3021,N_2993);
or U5375 (N_5375,N_2995,N_3476);
nor U5376 (N_5376,N_2463,N_3047);
or U5377 (N_5377,N_2510,N_3607);
or U5378 (N_5378,N_3906,N_3990);
and U5379 (N_5379,N_3011,N_2635);
nand U5380 (N_5380,N_3397,N_2098);
or U5381 (N_5381,N_3667,N_3817);
nor U5382 (N_5382,N_3219,N_3029);
or U5383 (N_5383,N_2247,N_3382);
or U5384 (N_5384,N_3602,N_2276);
nor U5385 (N_5385,N_2689,N_3076);
or U5386 (N_5386,N_2001,N_2931);
and U5387 (N_5387,N_3867,N_2750);
nor U5388 (N_5388,N_2385,N_2792);
and U5389 (N_5389,N_2043,N_2530);
nand U5390 (N_5390,N_3302,N_3127);
nand U5391 (N_5391,N_2077,N_2420);
and U5392 (N_5392,N_2964,N_3538);
nor U5393 (N_5393,N_2758,N_2436);
nand U5394 (N_5394,N_2504,N_2661);
nand U5395 (N_5395,N_2302,N_2604);
or U5396 (N_5396,N_3219,N_3937);
xor U5397 (N_5397,N_2952,N_2438);
or U5398 (N_5398,N_3962,N_3108);
or U5399 (N_5399,N_3692,N_2302);
nand U5400 (N_5400,N_2719,N_2867);
nor U5401 (N_5401,N_3536,N_3292);
and U5402 (N_5402,N_2788,N_2696);
nand U5403 (N_5403,N_2923,N_2061);
nand U5404 (N_5404,N_3248,N_3111);
or U5405 (N_5405,N_3858,N_2720);
or U5406 (N_5406,N_3738,N_2430);
and U5407 (N_5407,N_3354,N_2916);
nand U5408 (N_5408,N_2666,N_3997);
nor U5409 (N_5409,N_2945,N_3931);
or U5410 (N_5410,N_3677,N_2239);
nand U5411 (N_5411,N_2924,N_2209);
and U5412 (N_5412,N_3914,N_2974);
and U5413 (N_5413,N_3373,N_3003);
and U5414 (N_5414,N_2507,N_3645);
nand U5415 (N_5415,N_3719,N_2992);
nor U5416 (N_5416,N_2818,N_3234);
nand U5417 (N_5417,N_3340,N_3118);
nor U5418 (N_5418,N_3416,N_3079);
and U5419 (N_5419,N_2224,N_3769);
or U5420 (N_5420,N_2394,N_3172);
nand U5421 (N_5421,N_2961,N_2122);
or U5422 (N_5422,N_3940,N_2720);
and U5423 (N_5423,N_3616,N_3820);
xor U5424 (N_5424,N_2595,N_3266);
nor U5425 (N_5425,N_2208,N_2519);
or U5426 (N_5426,N_3541,N_3569);
and U5427 (N_5427,N_3789,N_2824);
and U5428 (N_5428,N_2490,N_2996);
nor U5429 (N_5429,N_3081,N_2051);
or U5430 (N_5430,N_3444,N_3774);
or U5431 (N_5431,N_2255,N_2008);
nand U5432 (N_5432,N_3107,N_3986);
and U5433 (N_5433,N_3394,N_2549);
or U5434 (N_5434,N_2171,N_3340);
and U5435 (N_5435,N_2748,N_2727);
or U5436 (N_5436,N_2250,N_2104);
and U5437 (N_5437,N_2503,N_2377);
nor U5438 (N_5438,N_2759,N_2043);
nand U5439 (N_5439,N_2738,N_2978);
nand U5440 (N_5440,N_3683,N_2840);
nand U5441 (N_5441,N_2914,N_2071);
xnor U5442 (N_5442,N_2388,N_3600);
nor U5443 (N_5443,N_3164,N_3908);
and U5444 (N_5444,N_3393,N_3885);
nand U5445 (N_5445,N_2150,N_3303);
and U5446 (N_5446,N_3467,N_2166);
and U5447 (N_5447,N_2189,N_2370);
or U5448 (N_5448,N_3312,N_3637);
or U5449 (N_5449,N_2703,N_3573);
or U5450 (N_5450,N_3694,N_3722);
or U5451 (N_5451,N_2622,N_2032);
and U5452 (N_5452,N_3207,N_3469);
or U5453 (N_5453,N_2346,N_2432);
nor U5454 (N_5454,N_2973,N_2399);
nand U5455 (N_5455,N_2653,N_3970);
and U5456 (N_5456,N_2255,N_2970);
or U5457 (N_5457,N_3841,N_2449);
and U5458 (N_5458,N_2001,N_2045);
and U5459 (N_5459,N_2553,N_3001);
nor U5460 (N_5460,N_3934,N_2398);
and U5461 (N_5461,N_2965,N_2464);
or U5462 (N_5462,N_2660,N_2280);
nand U5463 (N_5463,N_2305,N_3586);
nor U5464 (N_5464,N_2557,N_2975);
nand U5465 (N_5465,N_2051,N_3766);
nor U5466 (N_5466,N_3146,N_2246);
and U5467 (N_5467,N_3226,N_3400);
and U5468 (N_5468,N_2241,N_3895);
nand U5469 (N_5469,N_2455,N_3111);
or U5470 (N_5470,N_2776,N_3054);
nand U5471 (N_5471,N_3985,N_3814);
and U5472 (N_5472,N_3609,N_2205);
and U5473 (N_5473,N_2985,N_2637);
or U5474 (N_5474,N_3818,N_3607);
nand U5475 (N_5475,N_2847,N_2216);
nor U5476 (N_5476,N_2167,N_2511);
nand U5477 (N_5477,N_3050,N_3115);
nand U5478 (N_5478,N_2664,N_3809);
nor U5479 (N_5479,N_2752,N_2602);
nand U5480 (N_5480,N_2714,N_2128);
nor U5481 (N_5481,N_3300,N_2109);
nor U5482 (N_5482,N_3543,N_3746);
and U5483 (N_5483,N_3052,N_3709);
and U5484 (N_5484,N_2649,N_3315);
or U5485 (N_5485,N_3046,N_2392);
nor U5486 (N_5486,N_3658,N_3777);
and U5487 (N_5487,N_3873,N_2302);
nor U5488 (N_5488,N_2711,N_3248);
nor U5489 (N_5489,N_2110,N_3128);
or U5490 (N_5490,N_3508,N_2915);
nor U5491 (N_5491,N_2643,N_2428);
and U5492 (N_5492,N_3867,N_3657);
nor U5493 (N_5493,N_3354,N_2792);
or U5494 (N_5494,N_2856,N_2693);
or U5495 (N_5495,N_3035,N_2268);
nor U5496 (N_5496,N_3992,N_3230);
or U5497 (N_5497,N_2068,N_2125);
and U5498 (N_5498,N_3509,N_3403);
and U5499 (N_5499,N_2665,N_3873);
nand U5500 (N_5500,N_2567,N_3926);
nand U5501 (N_5501,N_3644,N_2056);
and U5502 (N_5502,N_3609,N_2833);
and U5503 (N_5503,N_2609,N_3027);
nor U5504 (N_5504,N_3109,N_3880);
or U5505 (N_5505,N_3233,N_2993);
nand U5506 (N_5506,N_2580,N_3006);
or U5507 (N_5507,N_2402,N_3679);
nor U5508 (N_5508,N_3186,N_2819);
and U5509 (N_5509,N_2424,N_2828);
nand U5510 (N_5510,N_3566,N_2034);
nand U5511 (N_5511,N_3914,N_2992);
or U5512 (N_5512,N_2258,N_3219);
and U5513 (N_5513,N_3959,N_3975);
or U5514 (N_5514,N_3760,N_3432);
xnor U5515 (N_5515,N_3659,N_3978);
and U5516 (N_5516,N_3477,N_3456);
nor U5517 (N_5517,N_2822,N_3683);
nand U5518 (N_5518,N_3881,N_3797);
nand U5519 (N_5519,N_3168,N_2673);
or U5520 (N_5520,N_2315,N_2221);
nor U5521 (N_5521,N_2728,N_3369);
nor U5522 (N_5522,N_3365,N_2198);
nor U5523 (N_5523,N_2849,N_3829);
or U5524 (N_5524,N_3035,N_3263);
or U5525 (N_5525,N_2392,N_2726);
nor U5526 (N_5526,N_3036,N_2068);
nand U5527 (N_5527,N_3547,N_3825);
nor U5528 (N_5528,N_2299,N_3080);
and U5529 (N_5529,N_2204,N_3403);
or U5530 (N_5530,N_3436,N_3169);
nor U5531 (N_5531,N_3646,N_2674);
and U5532 (N_5532,N_3712,N_2605);
nand U5533 (N_5533,N_2713,N_2361);
or U5534 (N_5534,N_3426,N_2333);
and U5535 (N_5535,N_3466,N_2778);
or U5536 (N_5536,N_2498,N_3139);
or U5537 (N_5537,N_3278,N_2067);
and U5538 (N_5538,N_3657,N_2667);
nor U5539 (N_5539,N_2232,N_3384);
and U5540 (N_5540,N_3050,N_3634);
and U5541 (N_5541,N_3548,N_2507);
or U5542 (N_5542,N_2996,N_3846);
nand U5543 (N_5543,N_3651,N_2167);
nand U5544 (N_5544,N_3714,N_3324);
xor U5545 (N_5545,N_2670,N_3786);
and U5546 (N_5546,N_3620,N_2846);
nand U5547 (N_5547,N_3421,N_3356);
and U5548 (N_5548,N_3217,N_2873);
nor U5549 (N_5549,N_2841,N_3757);
or U5550 (N_5550,N_3599,N_2638);
or U5551 (N_5551,N_2252,N_3338);
nand U5552 (N_5552,N_2453,N_2166);
nor U5553 (N_5553,N_3861,N_3919);
nor U5554 (N_5554,N_2234,N_3516);
nor U5555 (N_5555,N_3175,N_2486);
or U5556 (N_5556,N_2641,N_3601);
xnor U5557 (N_5557,N_2129,N_2279);
or U5558 (N_5558,N_2568,N_3929);
or U5559 (N_5559,N_2776,N_2056);
nor U5560 (N_5560,N_3908,N_3974);
or U5561 (N_5561,N_3867,N_2902);
nand U5562 (N_5562,N_3745,N_2519);
nor U5563 (N_5563,N_2410,N_2124);
and U5564 (N_5564,N_3653,N_2259);
nand U5565 (N_5565,N_2220,N_3635);
or U5566 (N_5566,N_3696,N_2348);
nor U5567 (N_5567,N_3248,N_3571);
or U5568 (N_5568,N_2326,N_2407);
nand U5569 (N_5569,N_2765,N_2041);
nand U5570 (N_5570,N_2765,N_3759);
and U5571 (N_5571,N_2216,N_2879);
and U5572 (N_5572,N_2793,N_3103);
and U5573 (N_5573,N_2930,N_2447);
nand U5574 (N_5574,N_3896,N_2632);
or U5575 (N_5575,N_2414,N_3335);
xor U5576 (N_5576,N_2085,N_2770);
nand U5577 (N_5577,N_2486,N_2335);
or U5578 (N_5578,N_2131,N_3199);
nand U5579 (N_5579,N_2550,N_2953);
or U5580 (N_5580,N_2443,N_3792);
or U5581 (N_5581,N_2460,N_3899);
nand U5582 (N_5582,N_2226,N_3714);
nor U5583 (N_5583,N_3892,N_2654);
or U5584 (N_5584,N_3062,N_3094);
and U5585 (N_5585,N_3200,N_2613);
or U5586 (N_5586,N_2357,N_2728);
or U5587 (N_5587,N_2111,N_3400);
nand U5588 (N_5588,N_2403,N_2939);
or U5589 (N_5589,N_2292,N_3090);
nand U5590 (N_5590,N_3182,N_3859);
nor U5591 (N_5591,N_2148,N_3660);
nand U5592 (N_5592,N_2910,N_3511);
nand U5593 (N_5593,N_3615,N_3955);
and U5594 (N_5594,N_2696,N_2251);
nor U5595 (N_5595,N_2405,N_3348);
nand U5596 (N_5596,N_2109,N_3108);
or U5597 (N_5597,N_3381,N_3236);
and U5598 (N_5598,N_3519,N_3066);
and U5599 (N_5599,N_2559,N_3716);
nand U5600 (N_5600,N_3527,N_3694);
nor U5601 (N_5601,N_3674,N_2710);
and U5602 (N_5602,N_3871,N_3536);
nor U5603 (N_5603,N_3065,N_2019);
and U5604 (N_5604,N_3800,N_2318);
nand U5605 (N_5605,N_2923,N_2752);
nand U5606 (N_5606,N_3998,N_3971);
or U5607 (N_5607,N_2579,N_3834);
nand U5608 (N_5608,N_3825,N_3441);
nor U5609 (N_5609,N_2246,N_2382);
nor U5610 (N_5610,N_2066,N_3978);
and U5611 (N_5611,N_2372,N_2436);
or U5612 (N_5612,N_3227,N_3071);
or U5613 (N_5613,N_3749,N_3800);
or U5614 (N_5614,N_3577,N_3015);
and U5615 (N_5615,N_3010,N_3360);
nor U5616 (N_5616,N_3658,N_3026);
and U5617 (N_5617,N_3885,N_2327);
nand U5618 (N_5618,N_2131,N_2431);
nand U5619 (N_5619,N_3305,N_3556);
nand U5620 (N_5620,N_2503,N_2362);
or U5621 (N_5621,N_3057,N_2037);
or U5622 (N_5622,N_3865,N_3909);
nand U5623 (N_5623,N_2566,N_2173);
and U5624 (N_5624,N_3860,N_2682);
nor U5625 (N_5625,N_3936,N_3580);
or U5626 (N_5626,N_3285,N_3893);
nor U5627 (N_5627,N_3221,N_2143);
nand U5628 (N_5628,N_2217,N_3000);
and U5629 (N_5629,N_2508,N_2923);
nand U5630 (N_5630,N_2950,N_3167);
nand U5631 (N_5631,N_2652,N_3274);
nor U5632 (N_5632,N_3924,N_2981);
nand U5633 (N_5633,N_2539,N_3745);
nor U5634 (N_5634,N_3030,N_3655);
nor U5635 (N_5635,N_2442,N_2638);
or U5636 (N_5636,N_2753,N_2877);
and U5637 (N_5637,N_2603,N_3816);
and U5638 (N_5638,N_2781,N_3954);
nand U5639 (N_5639,N_3710,N_2230);
nand U5640 (N_5640,N_3075,N_2770);
or U5641 (N_5641,N_3174,N_2739);
nand U5642 (N_5642,N_3398,N_2673);
and U5643 (N_5643,N_2077,N_2625);
or U5644 (N_5644,N_2036,N_3615);
nand U5645 (N_5645,N_3288,N_3284);
nand U5646 (N_5646,N_3277,N_3243);
and U5647 (N_5647,N_3683,N_3765);
nor U5648 (N_5648,N_3527,N_2078);
nor U5649 (N_5649,N_3609,N_2703);
or U5650 (N_5650,N_3652,N_3202);
nor U5651 (N_5651,N_3522,N_3791);
nand U5652 (N_5652,N_2579,N_3467);
nand U5653 (N_5653,N_2559,N_2553);
and U5654 (N_5654,N_2612,N_2632);
or U5655 (N_5655,N_3343,N_2511);
or U5656 (N_5656,N_2337,N_3486);
nor U5657 (N_5657,N_3758,N_3223);
nor U5658 (N_5658,N_2853,N_2657);
or U5659 (N_5659,N_2092,N_3563);
nor U5660 (N_5660,N_2726,N_3822);
and U5661 (N_5661,N_3695,N_2667);
nor U5662 (N_5662,N_3098,N_3480);
or U5663 (N_5663,N_2442,N_3455);
nand U5664 (N_5664,N_2830,N_2668);
nor U5665 (N_5665,N_3626,N_3330);
nand U5666 (N_5666,N_2056,N_2462);
xor U5667 (N_5667,N_2535,N_3596);
and U5668 (N_5668,N_2006,N_2079);
nand U5669 (N_5669,N_2417,N_3066);
and U5670 (N_5670,N_2219,N_3553);
nand U5671 (N_5671,N_2922,N_2920);
or U5672 (N_5672,N_3476,N_3595);
or U5673 (N_5673,N_3450,N_3934);
nor U5674 (N_5674,N_2256,N_2722);
nor U5675 (N_5675,N_2118,N_2890);
nor U5676 (N_5676,N_3474,N_3226);
or U5677 (N_5677,N_2542,N_2413);
or U5678 (N_5678,N_3745,N_2763);
or U5679 (N_5679,N_2882,N_3600);
nand U5680 (N_5680,N_2566,N_2185);
nand U5681 (N_5681,N_3928,N_2809);
or U5682 (N_5682,N_3771,N_3039);
nand U5683 (N_5683,N_3705,N_2166);
xor U5684 (N_5684,N_2365,N_2915);
and U5685 (N_5685,N_3432,N_2170);
or U5686 (N_5686,N_2987,N_3598);
nand U5687 (N_5687,N_2445,N_3723);
nand U5688 (N_5688,N_3427,N_3965);
nand U5689 (N_5689,N_3180,N_2670);
nor U5690 (N_5690,N_3475,N_3580);
nor U5691 (N_5691,N_3462,N_3701);
or U5692 (N_5692,N_2410,N_3804);
and U5693 (N_5693,N_2378,N_3905);
nor U5694 (N_5694,N_3512,N_2461);
nor U5695 (N_5695,N_2410,N_3729);
and U5696 (N_5696,N_2855,N_2626);
and U5697 (N_5697,N_2631,N_3255);
and U5698 (N_5698,N_3666,N_3636);
nor U5699 (N_5699,N_3615,N_3797);
nand U5700 (N_5700,N_3059,N_2613);
and U5701 (N_5701,N_3788,N_3689);
xnor U5702 (N_5702,N_3006,N_2286);
nand U5703 (N_5703,N_3103,N_3623);
nor U5704 (N_5704,N_2227,N_2051);
nand U5705 (N_5705,N_3139,N_2032);
nand U5706 (N_5706,N_3295,N_3920);
nor U5707 (N_5707,N_3041,N_3061);
nor U5708 (N_5708,N_3455,N_3355);
or U5709 (N_5709,N_2102,N_3197);
nor U5710 (N_5710,N_2592,N_2171);
nand U5711 (N_5711,N_3327,N_2876);
nand U5712 (N_5712,N_3993,N_3272);
nor U5713 (N_5713,N_3464,N_3060);
or U5714 (N_5714,N_3858,N_3723);
nor U5715 (N_5715,N_2272,N_2013);
nor U5716 (N_5716,N_3923,N_3541);
nor U5717 (N_5717,N_2663,N_2433);
nor U5718 (N_5718,N_3558,N_2008);
or U5719 (N_5719,N_2020,N_2985);
and U5720 (N_5720,N_2309,N_2472);
and U5721 (N_5721,N_3112,N_3272);
or U5722 (N_5722,N_2620,N_2144);
nand U5723 (N_5723,N_2764,N_2268);
or U5724 (N_5724,N_2474,N_3520);
nor U5725 (N_5725,N_2099,N_2653);
and U5726 (N_5726,N_2465,N_3068);
or U5727 (N_5727,N_2941,N_3210);
nor U5728 (N_5728,N_2018,N_2424);
or U5729 (N_5729,N_2909,N_2964);
nor U5730 (N_5730,N_3062,N_2120);
or U5731 (N_5731,N_3545,N_3897);
or U5732 (N_5732,N_3617,N_2869);
xnor U5733 (N_5733,N_2734,N_2936);
nor U5734 (N_5734,N_3951,N_3496);
or U5735 (N_5735,N_2186,N_2004);
nor U5736 (N_5736,N_2801,N_3623);
or U5737 (N_5737,N_2422,N_3370);
nand U5738 (N_5738,N_2509,N_2423);
or U5739 (N_5739,N_3215,N_3153);
nor U5740 (N_5740,N_3375,N_3366);
nor U5741 (N_5741,N_3529,N_2682);
and U5742 (N_5742,N_3270,N_3454);
nor U5743 (N_5743,N_2412,N_3293);
xnor U5744 (N_5744,N_2242,N_3841);
or U5745 (N_5745,N_2906,N_2692);
and U5746 (N_5746,N_3917,N_3565);
nand U5747 (N_5747,N_3027,N_3290);
or U5748 (N_5748,N_2049,N_3492);
or U5749 (N_5749,N_2160,N_3690);
nand U5750 (N_5750,N_3554,N_2086);
and U5751 (N_5751,N_2550,N_2727);
and U5752 (N_5752,N_3330,N_2938);
nor U5753 (N_5753,N_2503,N_3099);
or U5754 (N_5754,N_3387,N_3294);
nor U5755 (N_5755,N_2181,N_3242);
nor U5756 (N_5756,N_3619,N_2405);
or U5757 (N_5757,N_3808,N_3910);
nand U5758 (N_5758,N_3727,N_2979);
nand U5759 (N_5759,N_3481,N_3946);
or U5760 (N_5760,N_3055,N_2300);
and U5761 (N_5761,N_2513,N_2479);
and U5762 (N_5762,N_3378,N_2185);
nor U5763 (N_5763,N_3622,N_2554);
or U5764 (N_5764,N_2373,N_3556);
or U5765 (N_5765,N_2888,N_2678);
nand U5766 (N_5766,N_3698,N_3189);
nand U5767 (N_5767,N_2154,N_2400);
nor U5768 (N_5768,N_2921,N_3909);
nand U5769 (N_5769,N_2117,N_3206);
nand U5770 (N_5770,N_3585,N_2513);
or U5771 (N_5771,N_3976,N_2927);
nand U5772 (N_5772,N_2031,N_2295);
nor U5773 (N_5773,N_2452,N_3268);
or U5774 (N_5774,N_3051,N_2366);
nand U5775 (N_5775,N_2921,N_2878);
nand U5776 (N_5776,N_3755,N_3246);
or U5777 (N_5777,N_3344,N_3314);
and U5778 (N_5778,N_2785,N_3383);
nor U5779 (N_5779,N_3418,N_3780);
or U5780 (N_5780,N_3200,N_3073);
nor U5781 (N_5781,N_2963,N_3741);
nor U5782 (N_5782,N_3012,N_3969);
nand U5783 (N_5783,N_2036,N_2032);
or U5784 (N_5784,N_2321,N_3382);
nor U5785 (N_5785,N_2264,N_2702);
and U5786 (N_5786,N_2611,N_2433);
nand U5787 (N_5787,N_3863,N_2761);
nand U5788 (N_5788,N_2415,N_3794);
nand U5789 (N_5789,N_2380,N_3876);
nor U5790 (N_5790,N_2954,N_3749);
nor U5791 (N_5791,N_2531,N_2658);
nand U5792 (N_5792,N_2531,N_3162);
nor U5793 (N_5793,N_2053,N_2957);
or U5794 (N_5794,N_3351,N_3290);
nor U5795 (N_5795,N_3385,N_2021);
and U5796 (N_5796,N_2815,N_3863);
nand U5797 (N_5797,N_2101,N_2058);
and U5798 (N_5798,N_2696,N_2634);
nand U5799 (N_5799,N_2554,N_3922);
nand U5800 (N_5800,N_2284,N_2888);
or U5801 (N_5801,N_3225,N_2860);
or U5802 (N_5802,N_2022,N_3500);
or U5803 (N_5803,N_3019,N_3392);
nand U5804 (N_5804,N_2544,N_3424);
or U5805 (N_5805,N_2768,N_3657);
and U5806 (N_5806,N_3430,N_2011);
nand U5807 (N_5807,N_3544,N_3550);
nand U5808 (N_5808,N_3743,N_2707);
and U5809 (N_5809,N_3160,N_2616);
or U5810 (N_5810,N_3670,N_2756);
and U5811 (N_5811,N_3908,N_2624);
nand U5812 (N_5812,N_3701,N_2098);
and U5813 (N_5813,N_2042,N_2144);
or U5814 (N_5814,N_3291,N_2099);
nand U5815 (N_5815,N_3281,N_3841);
nor U5816 (N_5816,N_3122,N_2492);
nand U5817 (N_5817,N_2186,N_2985);
nor U5818 (N_5818,N_3872,N_3010);
nand U5819 (N_5819,N_2851,N_3802);
nor U5820 (N_5820,N_3916,N_2344);
nor U5821 (N_5821,N_2007,N_3552);
nor U5822 (N_5822,N_3788,N_2308);
nor U5823 (N_5823,N_2233,N_3977);
nand U5824 (N_5824,N_3945,N_3482);
nor U5825 (N_5825,N_3921,N_2902);
nand U5826 (N_5826,N_3044,N_2826);
xnor U5827 (N_5827,N_3300,N_3789);
nand U5828 (N_5828,N_3841,N_2186);
nand U5829 (N_5829,N_3112,N_3707);
nand U5830 (N_5830,N_3936,N_3856);
nor U5831 (N_5831,N_3187,N_3864);
nor U5832 (N_5832,N_3873,N_2437);
nand U5833 (N_5833,N_3706,N_2332);
and U5834 (N_5834,N_2784,N_3720);
nand U5835 (N_5835,N_2483,N_2594);
xor U5836 (N_5836,N_3724,N_2965);
or U5837 (N_5837,N_2216,N_3919);
and U5838 (N_5838,N_2459,N_3277);
nor U5839 (N_5839,N_3747,N_2788);
nor U5840 (N_5840,N_2691,N_2187);
nand U5841 (N_5841,N_2454,N_2249);
and U5842 (N_5842,N_3282,N_3010);
and U5843 (N_5843,N_3397,N_2058);
nand U5844 (N_5844,N_3532,N_3462);
and U5845 (N_5845,N_2106,N_2412);
nand U5846 (N_5846,N_2640,N_3087);
and U5847 (N_5847,N_2138,N_2167);
xor U5848 (N_5848,N_3619,N_2095);
nor U5849 (N_5849,N_3466,N_3158);
nand U5850 (N_5850,N_3679,N_2586);
or U5851 (N_5851,N_3934,N_2618);
and U5852 (N_5852,N_2367,N_2626);
nand U5853 (N_5853,N_3122,N_2485);
nand U5854 (N_5854,N_3510,N_2591);
nand U5855 (N_5855,N_2027,N_2810);
and U5856 (N_5856,N_3925,N_3942);
nor U5857 (N_5857,N_2246,N_3311);
nor U5858 (N_5858,N_3897,N_2385);
nor U5859 (N_5859,N_3260,N_2726);
nand U5860 (N_5860,N_2572,N_3337);
nor U5861 (N_5861,N_2066,N_2032);
nand U5862 (N_5862,N_3144,N_2949);
and U5863 (N_5863,N_2473,N_2819);
nand U5864 (N_5864,N_3636,N_2417);
nand U5865 (N_5865,N_3796,N_3978);
nor U5866 (N_5866,N_3084,N_3121);
nor U5867 (N_5867,N_2707,N_3456);
and U5868 (N_5868,N_3390,N_2568);
nor U5869 (N_5869,N_2264,N_2445);
or U5870 (N_5870,N_3272,N_2485);
or U5871 (N_5871,N_2289,N_2745);
and U5872 (N_5872,N_3634,N_3043);
or U5873 (N_5873,N_3844,N_2372);
nand U5874 (N_5874,N_2512,N_2902);
and U5875 (N_5875,N_3634,N_3535);
xor U5876 (N_5876,N_2542,N_2321);
and U5877 (N_5877,N_2418,N_2435);
or U5878 (N_5878,N_3434,N_3893);
nand U5879 (N_5879,N_2053,N_2475);
nor U5880 (N_5880,N_3187,N_2537);
and U5881 (N_5881,N_3374,N_2966);
nand U5882 (N_5882,N_3357,N_2394);
nor U5883 (N_5883,N_3615,N_3972);
and U5884 (N_5884,N_2985,N_3717);
or U5885 (N_5885,N_2131,N_2906);
and U5886 (N_5886,N_2338,N_2688);
nand U5887 (N_5887,N_3387,N_3985);
nor U5888 (N_5888,N_2614,N_3704);
and U5889 (N_5889,N_2351,N_2003);
nand U5890 (N_5890,N_2436,N_3251);
nand U5891 (N_5891,N_2003,N_2258);
nand U5892 (N_5892,N_2837,N_2107);
or U5893 (N_5893,N_2698,N_2511);
or U5894 (N_5894,N_3148,N_3368);
or U5895 (N_5895,N_3205,N_3969);
nand U5896 (N_5896,N_3161,N_3675);
nand U5897 (N_5897,N_2305,N_3665);
nor U5898 (N_5898,N_2256,N_2100);
nand U5899 (N_5899,N_2929,N_3515);
or U5900 (N_5900,N_3941,N_3705);
nand U5901 (N_5901,N_3834,N_2211);
or U5902 (N_5902,N_3631,N_3676);
and U5903 (N_5903,N_2228,N_2313);
and U5904 (N_5904,N_2454,N_2866);
xor U5905 (N_5905,N_2861,N_2342);
nor U5906 (N_5906,N_2426,N_2555);
or U5907 (N_5907,N_3424,N_3268);
nor U5908 (N_5908,N_3076,N_3350);
and U5909 (N_5909,N_2278,N_2549);
nand U5910 (N_5910,N_2467,N_3453);
and U5911 (N_5911,N_3605,N_3023);
nand U5912 (N_5912,N_2774,N_2692);
and U5913 (N_5913,N_3951,N_3288);
or U5914 (N_5914,N_3207,N_3927);
and U5915 (N_5915,N_2979,N_3489);
nand U5916 (N_5916,N_3762,N_2346);
nor U5917 (N_5917,N_3514,N_3731);
and U5918 (N_5918,N_3005,N_3066);
and U5919 (N_5919,N_2265,N_3406);
nand U5920 (N_5920,N_3346,N_2898);
or U5921 (N_5921,N_2196,N_3178);
and U5922 (N_5922,N_2364,N_3570);
and U5923 (N_5923,N_3478,N_2655);
nor U5924 (N_5924,N_2754,N_3320);
nor U5925 (N_5925,N_3645,N_3446);
nand U5926 (N_5926,N_3048,N_3213);
nand U5927 (N_5927,N_2986,N_3719);
and U5928 (N_5928,N_3999,N_2330);
nand U5929 (N_5929,N_2805,N_3190);
nor U5930 (N_5930,N_3535,N_3362);
or U5931 (N_5931,N_2692,N_2388);
nor U5932 (N_5932,N_3632,N_2610);
nand U5933 (N_5933,N_2682,N_3281);
nand U5934 (N_5934,N_3786,N_2038);
or U5935 (N_5935,N_2217,N_3450);
and U5936 (N_5936,N_2596,N_2123);
or U5937 (N_5937,N_2003,N_3580);
and U5938 (N_5938,N_2200,N_2497);
nor U5939 (N_5939,N_2378,N_2201);
or U5940 (N_5940,N_3745,N_2602);
nor U5941 (N_5941,N_2545,N_3232);
nor U5942 (N_5942,N_3841,N_3555);
and U5943 (N_5943,N_3677,N_2777);
nand U5944 (N_5944,N_3133,N_3768);
and U5945 (N_5945,N_2565,N_3790);
nor U5946 (N_5946,N_2108,N_3561);
and U5947 (N_5947,N_2042,N_2790);
nand U5948 (N_5948,N_3473,N_2634);
xnor U5949 (N_5949,N_2265,N_2849);
or U5950 (N_5950,N_3533,N_2892);
and U5951 (N_5951,N_3602,N_3976);
nand U5952 (N_5952,N_2489,N_3843);
nand U5953 (N_5953,N_2072,N_3633);
and U5954 (N_5954,N_3224,N_3739);
and U5955 (N_5955,N_3042,N_2501);
nor U5956 (N_5956,N_3627,N_2037);
or U5957 (N_5957,N_3354,N_3603);
nand U5958 (N_5958,N_3134,N_3336);
nor U5959 (N_5959,N_2007,N_3476);
nor U5960 (N_5960,N_2737,N_2267);
nand U5961 (N_5961,N_2897,N_2249);
and U5962 (N_5962,N_3241,N_2119);
nor U5963 (N_5963,N_3415,N_2086);
nor U5964 (N_5964,N_3351,N_3180);
or U5965 (N_5965,N_3604,N_2186);
nor U5966 (N_5966,N_3887,N_3627);
xnor U5967 (N_5967,N_2146,N_3515);
nand U5968 (N_5968,N_3355,N_3058);
nor U5969 (N_5969,N_3095,N_3982);
or U5970 (N_5970,N_2919,N_3121);
nand U5971 (N_5971,N_2007,N_2988);
and U5972 (N_5972,N_3191,N_3782);
nand U5973 (N_5973,N_3211,N_2019);
nor U5974 (N_5974,N_3923,N_3506);
nor U5975 (N_5975,N_3844,N_3101);
nand U5976 (N_5976,N_3452,N_3549);
and U5977 (N_5977,N_2525,N_3453);
nand U5978 (N_5978,N_2788,N_2624);
and U5979 (N_5979,N_3964,N_2147);
and U5980 (N_5980,N_2043,N_2161);
nand U5981 (N_5981,N_2299,N_3381);
nand U5982 (N_5982,N_3957,N_3332);
nor U5983 (N_5983,N_2445,N_3861);
or U5984 (N_5984,N_2256,N_2429);
and U5985 (N_5985,N_3733,N_2593);
or U5986 (N_5986,N_3113,N_2469);
nor U5987 (N_5987,N_3479,N_2797);
nor U5988 (N_5988,N_3005,N_2712);
nor U5989 (N_5989,N_3767,N_3563);
or U5990 (N_5990,N_2706,N_2206);
nor U5991 (N_5991,N_3640,N_3382);
nor U5992 (N_5992,N_3352,N_3776);
nand U5993 (N_5993,N_2058,N_2506);
nor U5994 (N_5994,N_3416,N_3742);
nor U5995 (N_5995,N_3907,N_3605);
or U5996 (N_5996,N_3772,N_2459);
nand U5997 (N_5997,N_2067,N_3057);
nand U5998 (N_5998,N_3592,N_3789);
and U5999 (N_5999,N_3482,N_3931);
nor U6000 (N_6000,N_5196,N_4225);
nand U6001 (N_6001,N_5063,N_4209);
or U6002 (N_6002,N_5481,N_4931);
nand U6003 (N_6003,N_5230,N_4747);
nor U6004 (N_6004,N_4401,N_5467);
nor U6005 (N_6005,N_5014,N_4379);
nand U6006 (N_6006,N_4929,N_5113);
nand U6007 (N_6007,N_4997,N_5816);
nor U6008 (N_6008,N_4575,N_4163);
nor U6009 (N_6009,N_5912,N_5074);
nand U6010 (N_6010,N_5359,N_5708);
nand U6011 (N_6011,N_4740,N_5147);
and U6012 (N_6012,N_5652,N_4979);
and U6013 (N_6013,N_5123,N_4887);
and U6014 (N_6014,N_4812,N_5983);
and U6015 (N_6015,N_5465,N_4171);
and U6016 (N_6016,N_5223,N_4573);
or U6017 (N_6017,N_5535,N_4462);
and U6018 (N_6018,N_4988,N_4722);
nand U6019 (N_6019,N_4344,N_5870);
or U6020 (N_6020,N_5096,N_4598);
and U6021 (N_6021,N_4756,N_5441);
nor U6022 (N_6022,N_5410,N_4113);
nor U6023 (N_6023,N_5597,N_5140);
and U6024 (N_6024,N_4958,N_4565);
and U6025 (N_6025,N_4198,N_4847);
and U6026 (N_6026,N_4184,N_5706);
nor U6027 (N_6027,N_5973,N_4024);
nand U6028 (N_6028,N_5571,N_4153);
nor U6029 (N_6029,N_5177,N_4146);
and U6030 (N_6030,N_5087,N_4915);
nand U6031 (N_6031,N_4674,N_4214);
or U6032 (N_6032,N_4129,N_4571);
and U6033 (N_6033,N_4597,N_5601);
or U6034 (N_6034,N_5056,N_5026);
and U6035 (N_6035,N_5061,N_5784);
nand U6036 (N_6036,N_5842,N_5115);
nor U6037 (N_6037,N_5009,N_4823);
and U6038 (N_6038,N_4547,N_4307);
nor U6039 (N_6039,N_4730,N_4581);
nor U6040 (N_6040,N_5516,N_4249);
nor U6041 (N_6041,N_4215,N_5126);
and U6042 (N_6042,N_4441,N_4291);
and U6043 (N_6043,N_5015,N_5653);
or U6044 (N_6044,N_4874,N_4033);
nor U6045 (N_6045,N_5422,N_4155);
nand U6046 (N_6046,N_4270,N_4704);
and U6047 (N_6047,N_5710,N_5363);
nand U6048 (N_6048,N_5683,N_4533);
and U6049 (N_6049,N_4443,N_5709);
nor U6050 (N_6050,N_5689,N_4772);
nand U6051 (N_6051,N_4158,N_5540);
nand U6052 (N_6052,N_4051,N_4869);
nand U6053 (N_6053,N_4494,N_5360);
nand U6054 (N_6054,N_4309,N_5233);
nor U6055 (N_6055,N_4138,N_5867);
and U6056 (N_6056,N_5275,N_5331);
nand U6057 (N_6057,N_5081,N_4658);
xnor U6058 (N_6058,N_5023,N_5594);
or U6059 (N_6059,N_4172,N_4067);
or U6060 (N_6060,N_4147,N_5750);
nor U6061 (N_6061,N_4070,N_4527);
or U6062 (N_6062,N_5592,N_5137);
and U6063 (N_6063,N_5962,N_4851);
nand U6064 (N_6064,N_5338,N_5656);
nor U6065 (N_6065,N_4310,N_4422);
or U6066 (N_6066,N_4473,N_5333);
or U6067 (N_6067,N_5823,N_4805);
or U6068 (N_6068,N_4752,N_5863);
nor U6069 (N_6069,N_5805,N_5278);
nand U6070 (N_6070,N_5725,N_4457);
and U6071 (N_6071,N_5478,N_4058);
nand U6072 (N_6072,N_5088,N_5949);
or U6073 (N_6073,N_4993,N_5555);
or U6074 (N_6074,N_5578,N_4135);
nand U6075 (N_6075,N_4074,N_4435);
and U6076 (N_6076,N_4778,N_4061);
nand U6077 (N_6077,N_4817,N_4328);
and U6078 (N_6078,N_4056,N_4157);
nor U6079 (N_6079,N_4875,N_4286);
xnor U6080 (N_6080,N_5937,N_5513);
and U6081 (N_6081,N_5313,N_5854);
nand U6082 (N_6082,N_4140,N_4479);
nand U6083 (N_6083,N_4345,N_5099);
nand U6084 (N_6084,N_4322,N_4032);
nor U6085 (N_6085,N_4945,N_4230);
or U6086 (N_6086,N_5212,N_4671);
and U6087 (N_6087,N_4319,N_4925);
nand U6088 (N_6088,N_4118,N_5511);
nand U6089 (N_6089,N_5872,N_5766);
nand U6090 (N_6090,N_4275,N_4323);
or U6091 (N_6091,N_5118,N_4264);
nor U6092 (N_6092,N_5617,N_5092);
nor U6093 (N_6093,N_4470,N_4811);
nor U6094 (N_6094,N_4040,N_5728);
and U6095 (N_6095,N_4705,N_4072);
and U6096 (N_6096,N_5141,N_5925);
and U6097 (N_6097,N_4902,N_4006);
nor U6098 (N_6098,N_4743,N_5844);
nor U6099 (N_6099,N_5828,N_4097);
and U6100 (N_6100,N_4446,N_5544);
xnor U6101 (N_6101,N_4712,N_4354);
nand U6102 (N_6102,N_4130,N_5714);
or U6103 (N_6103,N_4487,N_5255);
and U6104 (N_6104,N_4739,N_5988);
nand U6105 (N_6105,N_4391,N_5538);
and U6106 (N_6106,N_4947,N_5616);
and U6107 (N_6107,N_4903,N_4976);
or U6108 (N_6108,N_5120,N_4090);
nor U6109 (N_6109,N_5839,N_4134);
and U6110 (N_6110,N_4458,N_5899);
nor U6111 (N_6111,N_5454,N_5902);
and U6112 (N_6112,N_5877,N_4289);
or U6113 (N_6113,N_4549,N_5146);
nor U6114 (N_6114,N_5724,N_5488);
nor U6115 (N_6115,N_5969,N_4834);
or U6116 (N_6116,N_4290,N_5200);
nand U6117 (N_6117,N_4604,N_4795);
nor U6118 (N_6118,N_5035,N_5394);
nand U6119 (N_6119,N_5694,N_5778);
nand U6120 (N_6120,N_5835,N_5453);
and U6121 (N_6121,N_5191,N_5636);
or U6122 (N_6122,N_4126,N_5105);
or U6123 (N_6123,N_4055,N_4418);
or U6124 (N_6124,N_5631,N_5320);
or U6125 (N_6125,N_5504,N_4689);
nand U6126 (N_6126,N_5443,N_5432);
and U6127 (N_6127,N_5249,N_5271);
nand U6128 (N_6128,N_5067,N_4848);
xor U6129 (N_6129,N_5852,N_5878);
nor U6130 (N_6130,N_5319,N_4934);
or U6131 (N_6131,N_4666,N_4992);
and U6132 (N_6132,N_5183,N_5507);
and U6133 (N_6133,N_4169,N_4905);
nor U6134 (N_6134,N_4116,N_5545);
and U6135 (N_6135,N_5554,N_5368);
nor U6136 (N_6136,N_5590,N_4259);
or U6137 (N_6137,N_5431,N_4092);
nor U6138 (N_6138,N_4687,N_4237);
nor U6139 (N_6139,N_5859,N_4193);
and U6140 (N_6140,N_5938,N_5259);
or U6141 (N_6141,N_4480,N_4601);
nor U6142 (N_6142,N_4477,N_4166);
nor U6143 (N_6143,N_5756,N_4577);
nor U6144 (N_6144,N_4205,N_4330);
and U6145 (N_6145,N_5471,N_4190);
and U6146 (N_6146,N_5101,N_4818);
nor U6147 (N_6147,N_4626,N_4912);
or U6148 (N_6148,N_4326,N_5225);
nor U6149 (N_6149,N_5711,N_4497);
nor U6150 (N_6150,N_4724,N_5868);
and U6151 (N_6151,N_4766,N_5794);
or U6152 (N_6152,N_4893,N_4211);
nor U6153 (N_6153,N_4396,N_5598);
or U6154 (N_6154,N_4510,N_5384);
and U6155 (N_6155,N_4895,N_4797);
nand U6156 (N_6156,N_4474,N_4349);
or U6157 (N_6157,N_4484,N_5595);
or U6158 (N_6158,N_5845,N_5989);
nor U6159 (N_6159,N_4989,N_4132);
or U6160 (N_6160,N_4159,N_5559);
nor U6161 (N_6161,N_5059,N_5857);
and U6162 (N_6162,N_4376,N_5898);
or U6163 (N_6163,N_5730,N_5678);
nor U6164 (N_6164,N_4420,N_4566);
nand U6165 (N_6165,N_5326,N_5029);
and U6166 (N_6166,N_4896,N_4331);
nor U6167 (N_6167,N_5186,N_4068);
and U6168 (N_6168,N_4620,N_4570);
and U6169 (N_6169,N_5517,N_4599);
nor U6170 (N_6170,N_5502,N_5715);
and U6171 (N_6171,N_5165,N_4721);
or U6172 (N_6172,N_4372,N_4605);
or U6173 (N_6173,N_4417,N_4252);
or U6174 (N_6174,N_5787,N_5232);
and U6175 (N_6175,N_4936,N_4187);
nor U6176 (N_6176,N_5312,N_4651);
xor U6177 (N_6177,N_4383,N_5619);
and U6178 (N_6178,N_4488,N_4318);
and U6179 (N_6179,N_5943,N_5676);
xor U6180 (N_6180,N_5090,N_4608);
or U6181 (N_6181,N_5344,N_5643);
nor U6182 (N_6182,N_5028,N_5748);
xnor U6183 (N_6183,N_4585,N_4445);
nor U6184 (N_6184,N_4016,N_5495);
nor U6185 (N_6185,N_5414,N_4516);
and U6186 (N_6186,N_4280,N_4406);
nor U6187 (N_6187,N_4862,N_5455);
and U6188 (N_6188,N_5966,N_5397);
nor U6189 (N_6189,N_4334,N_5365);
nand U6190 (N_6190,N_5248,N_4346);
nor U6191 (N_6191,N_5022,N_4112);
or U6192 (N_6192,N_5767,N_5956);
nand U6193 (N_6193,N_4253,N_4625);
and U6194 (N_6194,N_4386,N_4867);
nor U6195 (N_6195,N_4078,N_4174);
and U6196 (N_6196,N_5875,N_5716);
or U6197 (N_6197,N_4481,N_4048);
or U6198 (N_6198,N_5833,N_4063);
and U6199 (N_6199,N_5896,N_4492);
and U6200 (N_6200,N_5037,N_4922);
nor U6201 (N_6201,N_4195,N_4521);
and U6202 (N_6202,N_5679,N_5758);
nor U6203 (N_6203,N_5698,N_5489);
nor U6204 (N_6204,N_5985,N_5121);
nand U6205 (N_6205,N_5175,N_4222);
nor U6206 (N_6206,N_5144,N_4640);
and U6207 (N_6207,N_5219,N_4537);
nand U6208 (N_6208,N_5251,N_4871);
nor U6209 (N_6209,N_4419,N_5670);
and U6210 (N_6210,N_4025,N_5884);
and U6211 (N_6211,N_4127,N_5523);
and U6212 (N_6212,N_4935,N_5855);
or U6213 (N_6213,N_4557,N_5550);
nor U6214 (N_6214,N_5646,N_5905);
nand U6215 (N_6215,N_4831,N_5849);
and U6216 (N_6216,N_5494,N_4731);
or U6217 (N_6217,N_5935,N_5277);
nand U6218 (N_6218,N_5654,N_5135);
nand U6219 (N_6219,N_4273,N_4444);
and U6220 (N_6220,N_4432,N_5524);
or U6221 (N_6221,N_4489,N_4607);
or U6222 (N_6222,N_5776,N_4107);
and U6223 (N_6223,N_4927,N_5952);
nand U6224 (N_6224,N_5407,N_4125);
or U6225 (N_6225,N_4115,N_5560);
or U6226 (N_6226,N_5586,N_5040);
and U6227 (N_6227,N_5429,N_4631);
and U6228 (N_6228,N_5768,N_5366);
or U6229 (N_6229,N_5690,N_5939);
and U6230 (N_6230,N_5085,N_4426);
nand U6231 (N_6231,N_4296,N_4483);
nor U6232 (N_6232,N_5658,N_5600);
or U6233 (N_6233,N_4007,N_5972);
or U6234 (N_6234,N_5428,N_5328);
and U6235 (N_6235,N_4353,N_5389);
and U6236 (N_6236,N_4873,N_5562);
nand U6237 (N_6237,N_4734,N_4294);
or U6238 (N_6238,N_5286,N_4629);
or U6239 (N_6239,N_4676,N_5720);
and U6240 (N_6240,N_5083,N_4365);
nand U6241 (N_6241,N_4828,N_4799);
nor U6242 (N_6242,N_4921,N_4117);
and U6243 (N_6243,N_5945,N_5841);
nor U6244 (N_6244,N_5336,N_5874);
or U6245 (N_6245,N_4121,N_4042);
nand U6246 (N_6246,N_5624,N_5139);
nand U6247 (N_6247,N_4644,N_4940);
nand U6248 (N_6248,N_5542,N_5546);
and U6249 (N_6249,N_5179,N_4486);
and U6250 (N_6250,N_4911,N_5886);
and U6251 (N_6251,N_5158,N_4358);
nand U6252 (N_6252,N_5473,N_4202);
nand U6253 (N_6253,N_5587,N_5738);
or U6254 (N_6254,N_5496,N_5589);
nand U6255 (N_6255,N_5114,N_5370);
and U6256 (N_6256,N_4216,N_4083);
or U6257 (N_6257,N_4578,N_4909);
nor U6258 (N_6258,N_5532,N_4244);
nand U6259 (N_6259,N_5804,N_5942);
and U6260 (N_6260,N_4540,N_4005);
nand U6261 (N_6261,N_4775,N_5457);
nor U6262 (N_6262,N_4881,N_4161);
nand U6263 (N_6263,N_5439,N_5379);
or U6264 (N_6264,N_4711,N_5462);
nand U6265 (N_6265,N_4335,N_5563);
nand U6266 (N_6266,N_4239,N_4295);
nand U6267 (N_6267,N_4325,N_4939);
or U6268 (N_6268,N_4256,N_5591);
nand U6269 (N_6269,N_5607,N_5673);
nor U6270 (N_6270,N_4863,N_4539);
or U6271 (N_6271,N_5736,N_4877);
or U6272 (N_6272,N_5712,N_4229);
nor U6273 (N_6273,N_5045,N_4960);
or U6274 (N_6274,N_5469,N_4329);
nor U6275 (N_6275,N_4550,N_5041);
or U6276 (N_6276,N_4251,N_4675);
nand U6277 (N_6277,N_5387,N_5001);
and U6278 (N_6278,N_4170,N_5075);
and U6279 (N_6279,N_5926,N_4890);
nor U6280 (N_6280,N_5947,N_5528);
or U6281 (N_6281,N_5411,N_5953);
and U6282 (N_6282,N_4589,N_4762);
or U6283 (N_6283,N_4231,N_5227);
and U6284 (N_6284,N_4023,N_5871);
nor U6285 (N_6285,N_5779,N_4771);
or U6286 (N_6286,N_5188,N_5071);
nand U6287 (N_6287,N_4899,N_5820);
nand U6288 (N_6288,N_5285,N_4248);
and U6289 (N_6289,N_5306,N_5948);
nand U6290 (N_6290,N_4891,N_4637);
xor U6291 (N_6291,N_4368,N_5050);
and U6292 (N_6292,N_4703,N_5311);
and U6293 (N_6293,N_5463,N_4199);
nor U6294 (N_6294,N_5330,N_4652);
and U6295 (N_6295,N_5065,N_5780);
nand U6296 (N_6296,N_4995,N_4080);
or U6297 (N_6297,N_4846,N_4971);
nor U6298 (N_6298,N_4816,N_5548);
nor U6299 (N_6299,N_5644,N_5556);
nor U6300 (N_6300,N_4459,N_4627);
nand U6301 (N_6301,N_4260,N_4039);
nor U6302 (N_6302,N_5451,N_5686);
or U6303 (N_6303,N_4036,N_4094);
and U6304 (N_6304,N_4543,N_5681);
and U6305 (N_6305,N_4034,N_5440);
and U6306 (N_6306,N_5765,N_4966);
and U6307 (N_6307,N_4523,N_5752);
and U6308 (N_6308,N_5322,N_5396);
or U6309 (N_6309,N_4969,N_4279);
and U6310 (N_6310,N_5826,N_5593);
or U6311 (N_6311,N_4564,N_5491);
nor U6312 (N_6312,N_5731,N_4498);
and U6313 (N_6313,N_5873,N_4183);
nand U6314 (N_6314,N_5419,N_5246);
nand U6315 (N_6315,N_4888,N_5222);
nor U6316 (N_6316,N_4892,N_4104);
or U6317 (N_6317,N_4228,N_4619);
nor U6318 (N_6318,N_5773,N_4210);
nand U6319 (N_6319,N_5066,N_4490);
or U6320 (N_6320,N_5124,N_5485);
nand U6321 (N_6321,N_5672,N_5922);
and U6322 (N_6322,N_4613,N_5723);
nor U6323 (N_6323,N_5732,N_5830);
xor U6324 (N_6324,N_4574,N_5660);
nor U6325 (N_6325,N_4408,N_5514);
nor U6326 (N_6326,N_5498,N_5913);
nand U6327 (N_6327,N_5142,N_4388);
nor U6328 (N_6328,N_4649,N_4587);
xor U6329 (N_6329,N_5818,N_4719);
nor U6330 (N_6330,N_4269,N_4041);
and U6331 (N_6331,N_4173,N_4341);
or U6332 (N_6332,N_5650,N_5053);
or U6333 (N_6333,N_4824,N_4563);
nor U6334 (N_6334,N_4636,N_4086);
or U6335 (N_6335,N_5763,N_5298);
nand U6336 (N_6336,N_5499,N_4833);
and U6337 (N_6337,N_5819,N_4615);
or U6338 (N_6338,N_5573,N_4994);
and U6339 (N_6339,N_5645,N_4491);
nand U6340 (N_6340,N_5889,N_5642);
or U6341 (N_6341,N_5080,N_5282);
nand U6342 (N_6342,N_4999,N_5011);
and U6343 (N_6343,N_4733,N_5194);
nor U6344 (N_6344,N_5615,N_4363);
nand U6345 (N_6345,N_5641,N_4332);
nor U6346 (N_6346,N_5385,N_4845);
and U6347 (N_6347,N_5981,N_4413);
and U6348 (N_6348,N_5490,N_5699);
xor U6349 (N_6349,N_4713,N_4367);
and U6350 (N_6350,N_5401,N_5418);
nor U6351 (N_6351,N_5149,N_4245);
xor U6352 (N_6352,N_4254,N_5004);
xnor U6353 (N_6353,N_4064,N_4438);
nor U6354 (N_6354,N_4904,N_5769);
or U6355 (N_6355,N_5605,N_5167);
nand U6356 (N_6356,N_5604,N_4044);
or U6357 (N_6357,N_4433,N_4013);
nand U6358 (N_6358,N_4440,N_4562);
or U6359 (N_6359,N_5549,N_4001);
nand U6360 (N_6360,N_4050,N_4065);
nand U6361 (N_6361,N_5622,N_5057);
nand U6362 (N_6362,N_4777,N_4937);
nor U6363 (N_6363,N_4351,N_4327);
nor U6364 (N_6364,N_5008,N_4456);
nor U6365 (N_6365,N_5713,N_5792);
nand U6366 (N_6366,N_4784,N_4263);
or U6367 (N_6367,N_4425,N_4633);
and U6368 (N_6368,N_5042,N_5971);
nor U6369 (N_6369,N_5695,N_5184);
nor U6370 (N_6370,N_5603,N_4352);
nand U6371 (N_6371,N_5892,N_4829);
and U6372 (N_6372,N_5376,N_5880);
nor U6373 (N_6373,N_5999,N_4077);
and U6374 (N_6374,N_5416,N_4535);
nand U6375 (N_6375,N_4678,N_4900);
or U6376 (N_6376,N_5089,N_4151);
nor U6377 (N_6377,N_4801,N_4439);
and U6378 (N_6378,N_5734,N_4381);
nand U6379 (N_6379,N_5903,N_5588);
and U6380 (N_6380,N_5793,N_5790);
and U6381 (N_6381,N_4879,N_5772);
and U6382 (N_6382,N_4946,N_5210);
or U6383 (N_6383,N_5975,N_4924);
and U6384 (N_6384,N_5343,N_5424);
nand U6385 (N_6385,N_5244,N_4528);
and U6386 (N_6386,N_5984,N_5521);
or U6387 (N_6387,N_4665,N_4953);
or U6388 (N_6388,N_5202,N_4447);
nor U6389 (N_6389,N_5822,N_5209);
and U6390 (N_6390,N_5228,N_5073);
and U6391 (N_6391,N_5257,N_4390);
nand U6392 (N_6392,N_4482,N_5515);
and U6393 (N_6393,N_5881,N_5677);
or U6394 (N_6394,N_4588,N_4788);
or U6395 (N_6395,N_5408,N_5858);
nand U6396 (N_6396,N_4505,N_4854);
nor U6397 (N_6397,N_5335,N_5657);
or U6398 (N_6398,N_5661,N_4819);
and U6399 (N_6399,N_5375,N_4669);
nor U6400 (N_6400,N_5479,N_5580);
xnor U6401 (N_6401,N_5309,N_5203);
and U6402 (N_6402,N_4360,N_5316);
nand U6403 (N_6403,N_4317,N_5904);
nand U6404 (N_6404,N_4430,N_4506);
nand U6405 (N_6405,N_5751,N_4201);
and U6406 (N_6406,N_5374,N_4460);
nor U6407 (N_6407,N_5812,N_5486);
and U6408 (N_6408,N_4003,N_5132);
nor U6409 (N_6409,N_5430,N_5036);
and U6410 (N_6410,N_4536,N_4612);
or U6411 (N_6411,N_5032,N_4411);
nor U6412 (N_6412,N_4266,N_4100);
or U6413 (N_6413,N_5051,N_4144);
or U6414 (N_6414,N_4688,N_4677);
nor U6415 (N_6415,N_5238,N_4503);
or U6416 (N_6416,N_5630,N_4624);
and U6417 (N_6417,N_5978,N_5434);
nor U6418 (N_6418,N_5287,N_5910);
nor U6419 (N_6419,N_5951,N_4943);
or U6420 (N_6420,N_5526,N_4808);
and U6421 (N_6421,N_5464,N_4876);
or U6422 (N_6422,N_4427,N_5688);
nand U6423 (N_6423,N_4405,N_4672);
and U6424 (N_6424,N_5152,N_4791);
or U6425 (N_6425,N_5628,N_4394);
nor U6426 (N_6426,N_4765,N_5433);
nand U6427 (N_6427,N_4787,N_4271);
nand U6428 (N_6428,N_5332,N_5252);
nor U6429 (N_6429,N_4384,N_5740);
and U6430 (N_6430,N_4038,N_4982);
and U6431 (N_6431,N_4313,N_5572);
nand U6432 (N_6432,N_5106,N_4333);
nor U6433 (N_6433,N_5475,N_4800);
nand U6434 (N_6434,N_5729,N_5638);
and U6435 (N_6435,N_5914,N_5078);
nand U6436 (N_6436,N_5258,N_5979);
nand U6437 (N_6437,N_5476,N_5378);
nand U6438 (N_6438,N_5019,N_4737);
nand U6439 (N_6439,N_4793,N_4815);
and U6440 (N_6440,N_5721,N_5371);
and U6441 (N_6441,N_5104,N_4224);
nor U6442 (N_6442,N_4218,N_5131);
and U6443 (N_6443,N_4047,N_5110);
or U6444 (N_6444,N_4683,N_5762);
or U6445 (N_6445,N_5837,N_5425);
nand U6446 (N_6446,N_4957,N_4268);
nand U6447 (N_6447,N_5302,N_5272);
nor U6448 (N_6448,N_5856,N_5500);
nor U6449 (N_6449,N_5193,N_4293);
nor U6450 (N_6450,N_5299,N_5497);
and U6451 (N_6451,N_5924,N_5757);
or U6452 (N_6452,N_4773,N_5204);
and U6453 (N_6453,N_5577,N_5530);
or U6454 (N_6454,N_5421,N_5130);
or U6455 (N_6455,N_5831,N_4814);
or U6456 (N_6456,N_5417,N_5569);
nor U6457 (N_6457,N_4403,N_5692);
nand U6458 (N_6458,N_4987,N_4544);
nor U6459 (N_6459,N_4062,N_4162);
or U6460 (N_6460,N_4998,N_5651);
xnor U6461 (N_6461,N_4022,N_4015);
nand U6462 (N_6462,N_4866,N_5799);
nand U6463 (N_6463,N_4395,N_4021);
nor U6464 (N_6464,N_5908,N_4694);
nor U6465 (N_6465,N_5602,N_5509);
or U6466 (N_6466,N_4926,N_4792);
and U6467 (N_6467,N_4339,N_4389);
nand U6468 (N_6468,N_5317,N_4301);
nand U6469 (N_6469,N_5484,N_4894);
and U6470 (N_6470,N_5348,N_5821);
or U6471 (N_6471,N_5290,N_5518);
xnor U6472 (N_6472,N_5405,N_4701);
or U6473 (N_6473,N_4910,N_4298);
nor U6474 (N_6474,N_5682,N_4579);
and U6475 (N_6475,N_4504,N_5525);
or U6476 (N_6476,N_4710,N_5005);
or U6477 (N_6477,N_4542,N_4247);
nor U6478 (N_6478,N_4541,N_4517);
or U6479 (N_6479,N_4639,N_5997);
nand U6480 (N_6480,N_5707,N_5575);
nor U6481 (N_6481,N_5024,N_5006);
nand U6482 (N_6482,N_4750,N_4567);
nand U6483 (N_6483,N_5649,N_5119);
nand U6484 (N_6484,N_4622,N_5279);
and U6485 (N_6485,N_4179,N_5543);
nand U6486 (N_6486,N_4099,N_4402);
xor U6487 (N_6487,N_5231,N_5460);
nor U6488 (N_6488,N_4507,N_4968);
xor U6489 (N_6489,N_4803,N_4308);
nand U6490 (N_6490,N_5129,N_5351);
nand U6491 (N_6491,N_5260,N_4780);
nand U6492 (N_6492,N_5668,N_5062);
nor U6493 (N_6493,N_4534,N_5280);
and U6494 (N_6494,N_4594,N_4820);
nand U6495 (N_6495,N_4188,N_5192);
nand U6496 (N_6496,N_5959,N_4697);
and U6497 (N_6497,N_4556,N_5472);
nand U6498 (N_6498,N_5125,N_4180);
nor U6499 (N_6499,N_4670,N_4970);
and U6500 (N_6500,N_4371,N_4250);
nor U6501 (N_6501,N_5111,N_5585);
or U6502 (N_6502,N_4096,N_4206);
or U6503 (N_6503,N_5452,N_5100);
and U6504 (N_6504,N_5388,N_5522);
or U6505 (N_6505,N_4399,N_4614);
or U6506 (N_6506,N_5741,N_4150);
or U6507 (N_6507,N_4685,N_4840);
or U6508 (N_6508,N_5304,N_4602);
nand U6509 (N_6509,N_4606,N_5380);
or U6510 (N_6510,N_4826,N_5329);
xor U6511 (N_6511,N_4977,N_4208);
nor U6512 (N_6512,N_4628,N_5323);
nor U6513 (N_6513,N_4884,N_5927);
and U6514 (N_6514,N_5836,N_4284);
nor U6515 (N_6515,N_5308,N_4786);
or U6516 (N_6516,N_4303,N_4682);
nor U6517 (N_6517,N_4880,N_5195);
nand U6518 (N_6518,N_5300,N_4176);
and U6519 (N_6519,N_4142,N_4240);
nand U6520 (N_6520,N_4967,N_4356);
or U6521 (N_6521,N_5996,N_4508);
nand U6522 (N_6522,N_4493,N_4223);
nor U6523 (N_6523,N_4496,N_5531);
nand U6524 (N_6524,N_5847,N_4431);
and U6525 (N_6525,N_4843,N_5865);
nor U6526 (N_6526,N_4751,N_4246);
and U6527 (N_6527,N_4119,N_5666);
nand U6528 (N_6528,N_5861,N_4568);
nor U6529 (N_6529,N_5611,N_5296);
or U6530 (N_6530,N_5869,N_5632);
nand U6531 (N_6531,N_5923,N_5404);
and U6532 (N_6532,N_4415,N_4769);
nand U6533 (N_6533,N_5684,N_4133);
nand U6534 (N_6534,N_5020,N_5327);
or U6535 (N_6535,N_4524,N_5138);
and U6536 (N_6536,N_4378,N_5944);
or U6537 (N_6537,N_4714,N_5506);
and U6538 (N_6538,N_5318,N_5353);
and U6539 (N_6539,N_4321,N_5955);
nor U6540 (N_6540,N_4538,N_5701);
and U6541 (N_6541,N_4928,N_4105);
nand U6542 (N_6542,N_5093,N_5153);
and U6543 (N_6543,N_4810,N_4079);
nand U6544 (N_6544,N_4583,N_4287);
or U6545 (N_6545,N_4128,N_5685);
nand U6546 (N_6546,N_5253,N_5064);
and U6547 (N_6547,N_4956,N_5002);
xnor U6548 (N_6548,N_4227,N_4436);
or U6549 (N_6549,N_4359,N_5533);
nor U6550 (N_6550,N_4108,N_4576);
nor U6551 (N_6551,N_5536,N_5276);
nor U6552 (N_6552,N_4745,N_5726);
or U6553 (N_6553,N_4110,N_4707);
and U6554 (N_6554,N_5640,N_5618);
nor U6555 (N_6555,N_5274,N_4716);
or U6556 (N_6556,N_5742,N_4634);
and U6557 (N_6557,N_5840,N_5609);
or U6558 (N_6558,N_4990,N_4783);
or U6559 (N_6559,N_5663,N_5033);
and U6560 (N_6560,N_4850,N_4409);
nor U6561 (N_6561,N_5807,N_5164);
xor U6562 (N_6562,N_5931,N_5626);
nand U6563 (N_6563,N_5704,N_4580);
nor U6564 (N_6564,N_5116,N_5176);
nand U6565 (N_6565,N_4680,N_5055);
and U6566 (N_6566,N_4996,N_5608);
nor U6567 (N_6567,N_4661,N_4111);
nand U6568 (N_6568,N_4770,N_4392);
nor U6569 (N_6569,N_5627,N_4272);
nor U6570 (N_6570,N_5901,N_5315);
nor U6571 (N_6571,N_4642,N_4343);
nand U6572 (N_6572,N_4790,N_4681);
and U6573 (N_6573,N_5749,N_4156);
and U6574 (N_6574,N_4098,N_5288);
nor U6575 (N_6575,N_5743,N_5367);
nand U6576 (N_6576,N_5218,N_4261);
or U6577 (N_6577,N_5885,N_5637);
nor U6578 (N_6578,N_4495,N_5437);
or U6579 (N_6579,N_5553,N_4026);
xor U6580 (N_6580,N_5091,N_4555);
and U6581 (N_6581,N_5505,N_4122);
and U6582 (N_6582,N_5534,N_4917);
or U6583 (N_6583,N_5474,N_5862);
nor U6584 (N_6584,N_4844,N_4525);
or U6585 (N_6585,N_5084,N_4720);
or U6586 (N_6586,N_5929,N_5224);
or U6587 (N_6587,N_5510,N_5697);
nand U6588 (N_6588,N_5117,N_4469);
nor U6589 (N_6589,N_5614,N_4760);
or U6590 (N_6590,N_5154,N_4693);
nand U6591 (N_6591,N_5963,N_5566);
and U6592 (N_6592,N_5393,N_5703);
xnor U6593 (N_6593,N_5825,N_5781);
or U6594 (N_6594,N_5007,N_5635);
nand U6595 (N_6595,N_4914,N_4569);
and U6596 (N_6596,N_4212,N_4088);
nand U6597 (N_6597,N_5127,N_4630);
nor U6598 (N_6598,N_5570,N_4638);
nor U6599 (N_6599,N_5163,N_5148);
and U6600 (N_6600,N_4238,N_5447);
or U6601 (N_6601,N_4145,N_5814);
and U6602 (N_6602,N_5941,N_5161);
or U6603 (N_6603,N_5797,N_5492);
nor U6604 (N_6604,N_4868,N_4428);
nor U6605 (N_6605,N_4164,N_4668);
nand U6606 (N_6606,N_4030,N_4748);
nand U6607 (N_6607,N_4476,N_4611);
nand U6608 (N_6608,N_4472,N_5890);
nand U6609 (N_6609,N_4220,N_4434);
nand U6610 (N_6610,N_4882,N_5894);
or U6611 (N_6611,N_4856,N_5806);
or U6612 (N_6612,N_5568,N_4715);
nor U6613 (N_6613,N_5800,N_4449);
or U6614 (N_6614,N_5970,N_4382);
or U6615 (N_6615,N_4203,N_5879);
or U6616 (N_6616,N_4609,N_5582);
xor U6617 (N_6617,N_5347,N_4553);
or U6618 (N_6618,N_5995,N_4725);
nor U6619 (N_6619,N_5000,N_4961);
and U6620 (N_6620,N_4742,N_4551);
nor U6621 (N_6621,N_5383,N_4466);
nor U6622 (N_6622,N_5391,N_5342);
nand U6623 (N_6623,N_4370,N_4653);
and U6624 (N_6624,N_4154,N_4191);
nand U6625 (N_6625,N_4759,N_5345);
nor U6626 (N_6626,N_5242,N_4763);
nand U6627 (N_6627,N_4101,N_5174);
nor U6628 (N_6628,N_4276,N_5846);
or U6629 (N_6629,N_5190,N_4031);
nand U6630 (N_6630,N_4861,N_4974);
and U6631 (N_6631,N_4610,N_5373);
nor U6632 (N_6632,N_5940,N_5283);
nand U6633 (N_6633,N_5851,N_5199);
nor U6634 (N_6634,N_5564,N_5221);
and U6635 (N_6635,N_4813,N_4908);
and U6636 (N_6636,N_4410,N_4362);
or U6637 (N_6637,N_5620,N_5159);
and U6638 (N_6638,N_5086,N_5128);
and U6639 (N_6639,N_5082,N_4374);
nand U6640 (N_6640,N_5567,N_4586);
and U6641 (N_6641,N_4336,N_5558);
and U6642 (N_6642,N_5965,N_4387);
and U6643 (N_6643,N_5964,N_4338);
and U6644 (N_6644,N_4776,N_5581);
nor U6645 (N_6645,N_5579,N_4949);
nand U6646 (N_6646,N_5334,N_4071);
or U6647 (N_6647,N_4702,N_4471);
nand U6648 (N_6648,N_4018,N_4149);
nand U6649 (N_6649,N_5900,N_5435);
and U6650 (N_6650,N_4274,N_5705);
nor U6651 (N_6651,N_5409,N_5906);
or U6652 (N_6652,N_5888,N_5017);
or U6653 (N_6653,N_4727,N_4085);
or U6654 (N_6654,N_4082,N_5596);
nand U6655 (N_6655,N_5266,N_5046);
or U6656 (N_6656,N_5395,N_5891);
and U6657 (N_6657,N_5702,N_5234);
and U6658 (N_6658,N_4849,N_5216);
or U6659 (N_6659,N_4746,N_5982);
nor U6660 (N_6660,N_4009,N_4029);
nor U6661 (N_6661,N_5012,N_5958);
and U6662 (N_6662,N_4398,N_5477);
and U6663 (N_6663,N_4963,N_5245);
or U6664 (N_6664,N_5264,N_5827);
nand U6665 (N_6665,N_4515,N_4554);
or U6666 (N_6666,N_4621,N_5480);
nand U6667 (N_6667,N_4204,N_5832);
nor U6668 (N_6668,N_5217,N_4311);
nand U6669 (N_6669,N_4511,N_4236);
and U6670 (N_6670,N_4832,N_4185);
or U6671 (N_6671,N_5034,N_5003);
or U6672 (N_6672,N_4706,N_4114);
nor U6673 (N_6673,N_5990,N_5883);
nor U6674 (N_6674,N_4020,N_4177);
nand U6675 (N_6675,N_4753,N_4708);
nand U6676 (N_6676,N_5362,N_5446);
and U6677 (N_6677,N_4821,N_5031);
and U6678 (N_6678,N_4278,N_4522);
or U6679 (N_6679,N_5449,N_5289);
and U6680 (N_6680,N_5427,N_4738);
and U6681 (N_6681,N_5519,N_5357);
and U6682 (N_6682,N_4729,N_4423);
or U6683 (N_6683,N_5102,N_5537);
and U6684 (N_6684,N_4450,N_5612);
nor U6685 (N_6685,N_4004,N_5917);
or U6686 (N_6686,N_5717,N_5811);
nor U6687 (N_6687,N_4809,N_5256);
and U6688 (N_6688,N_5267,N_4393);
and U6689 (N_6689,N_5508,N_4530);
or U6690 (N_6690,N_4768,N_5181);
nor U6691 (N_6691,N_4841,N_4350);
nand U6692 (N_6692,N_4827,N_4304);
or U6693 (N_6693,N_4648,N_5760);
nand U6694 (N_6694,N_5412,N_4948);
nor U6695 (N_6695,N_4475,N_4027);
or U6696 (N_6696,N_5789,N_5254);
and U6697 (N_6697,N_5044,N_5205);
or U6698 (N_6698,N_5932,N_5450);
and U6699 (N_6699,N_4641,N_4053);
nand U6700 (N_6700,N_4103,N_4897);
nand U6701 (N_6701,N_5423,N_4728);
or U6702 (N_6702,N_4448,N_5895);
nor U6703 (N_6703,N_4437,N_4454);
and U6704 (N_6704,N_4442,N_5722);
and U6705 (N_6705,N_4500,N_5468);
or U6706 (N_6706,N_4774,N_4019);
or U6707 (N_6707,N_5994,N_5786);
nand U6708 (N_6708,N_5070,N_4842);
nor U6709 (N_6709,N_5442,N_5314);
nor U6710 (N_6710,N_5829,N_5747);
nand U6711 (N_6711,N_4913,N_4830);
or U6712 (N_6712,N_4855,N_4741);
nor U6713 (N_6713,N_5539,N_4052);
and U6714 (N_6714,N_4340,N_5226);
nand U6715 (N_6715,N_5934,N_5341);
nand U6716 (N_6716,N_5662,N_4950);
or U6717 (N_6717,N_5108,N_5415);
nor U6718 (N_6718,N_4189,N_4690);
nand U6719 (N_6719,N_4299,N_5783);
nand U6720 (N_6720,N_5122,N_5897);
xor U6721 (N_6721,N_4717,N_4324);
nor U6722 (N_6722,N_4593,N_5356);
and U6723 (N_6723,N_5606,N_5301);
or U6724 (N_6724,N_5170,N_5187);
nand U6725 (N_6725,N_5961,N_5458);
nand U6726 (N_6726,N_5240,N_5459);
nand U6727 (N_6727,N_4046,N_4964);
nand U6728 (N_6728,N_4181,N_5236);
nand U6729 (N_6729,N_4478,N_4292);
nand U6730 (N_6730,N_4532,N_5785);
and U6731 (N_6731,N_4141,N_5503);
or U6732 (N_6732,N_4089,N_5625);
or U6733 (N_6733,N_5584,N_4075);
nor U6734 (N_6734,N_4785,N_5261);
nor U6735 (N_6735,N_4235,N_5361);
and U6736 (N_6736,N_5220,N_5921);
xnor U6737 (N_6737,N_5198,N_4518);
or U6738 (N_6738,N_4035,N_5399);
nand U6739 (N_6739,N_5853,N_4519);
or U6740 (N_6740,N_5700,N_4400);
nand U6741 (N_6741,N_4698,N_4858);
or U6742 (N_6742,N_4603,N_5243);
and U6743 (N_6743,N_5933,N_4463);
or U6744 (N_6744,N_5864,N_4552);
or U6745 (N_6745,N_4749,N_4499);
or U6746 (N_6746,N_4942,N_5991);
nand U6747 (N_6747,N_5305,N_5048);
and U6748 (N_6748,N_4014,N_5381);
or U6749 (N_6749,N_4980,N_4011);
or U6750 (N_6750,N_5954,N_4646);
or U6751 (N_6751,N_5173,N_5583);
or U6752 (N_6752,N_4316,N_5977);
nand U6753 (N_6753,N_4485,N_5946);
and U6754 (N_6754,N_5887,N_4520);
and U6755 (N_6755,N_5107,N_4468);
and U6756 (N_6756,N_4194,N_5143);
nand U6757 (N_6757,N_5882,N_5438);
or U6758 (N_6758,N_5671,N_5664);
nand U6759 (N_6759,N_5398,N_5824);
or U6760 (N_6760,N_4596,N_5273);
or U6761 (N_6761,N_5512,N_5103);
nor U6762 (N_6762,N_4196,N_5976);
or U6763 (N_6763,N_4081,N_4165);
nor U6764 (N_6764,N_5777,N_5160);
nand U6765 (N_6765,N_4959,N_5669);
or U6766 (N_6766,N_5696,N_4373);
or U6767 (N_6767,N_5796,N_4872);
nor U6768 (N_6768,N_4561,N_5456);
and U6769 (N_6769,N_4757,N_4087);
nand U6770 (N_6770,N_4424,N_5269);
nand U6771 (N_6771,N_5667,N_4377);
nor U6772 (N_6772,N_5876,N_4213);
or U6773 (N_6773,N_4796,N_5998);
or U6774 (N_6774,N_4735,N_5155);
nand U6775 (N_6775,N_4012,N_5094);
and U6776 (N_6776,N_5501,N_4955);
or U6777 (N_6777,N_5719,N_4559);
xnor U6778 (N_6778,N_5403,N_5809);
nor U6779 (N_6779,N_4870,N_5850);
nand U6780 (N_6780,N_4686,N_4919);
and U6781 (N_6781,N_4380,N_4654);
nand U6782 (N_6782,N_4962,N_5529);
nor U6783 (N_6783,N_5295,N_5813);
nand U6784 (N_6784,N_4804,N_5737);
and U6785 (N_6785,N_4091,N_4200);
nor U6786 (N_6786,N_5727,N_4277);
nand U6787 (N_6787,N_4513,N_4656);
nor U6788 (N_6788,N_5974,N_5150);
nor U6789 (N_6789,N_5038,N_4412);
or U6790 (N_6790,N_5551,N_5915);
or U6791 (N_6791,N_5054,N_5097);
and U6792 (N_6792,N_5613,N_5674);
nand U6793 (N_6793,N_5576,N_4529);
and U6794 (N_6794,N_5386,N_4838);
nand U6795 (N_6795,N_4825,N_5426);
and U6796 (N_6796,N_5206,N_4017);
and U6797 (N_6797,N_5303,N_5801);
nor U6798 (N_6798,N_4347,N_4985);
xor U6799 (N_6799,N_4660,N_4560);
and U6800 (N_6800,N_4952,N_5262);
nand U6801 (N_6801,N_5920,N_5733);
or U6802 (N_6802,N_5400,N_5021);
nand U6803 (N_6803,N_5659,N_5265);
or U6804 (N_6804,N_5178,N_5687);
nand U6805 (N_6805,N_4452,N_4167);
and U6806 (N_6806,N_4531,N_4857);
nor U6807 (N_6807,N_5634,N_4679);
and U6808 (N_6808,N_4696,N_4002);
nand U6809 (N_6809,N_4764,N_4084);
or U6810 (N_6810,N_4000,N_5647);
and U6811 (N_6811,N_4692,N_5860);
or U6812 (N_6812,N_5077,N_5281);
or U6813 (N_6813,N_5109,N_4718);
nand U6814 (N_6814,N_5466,N_5992);
and U6815 (N_6815,N_4501,N_4673);
and U6816 (N_6816,N_4691,N_4779);
and U6817 (N_6817,N_4152,N_5151);
nand U6818 (N_6818,N_4281,N_5098);
and U6819 (N_6819,N_5241,N_4465);
nor U6820 (N_6820,N_4933,N_4421);
nand U6821 (N_6821,N_4767,N_4972);
nand U6822 (N_6822,N_4057,N_5655);
nand U6823 (N_6823,N_5541,N_4923);
and U6824 (N_6824,N_4907,N_5382);
xor U6825 (N_6825,N_5207,N_5967);
or U6826 (N_6826,N_4109,N_5795);
and U6827 (N_6827,N_4918,N_4657);
nor U6828 (N_6828,N_5755,N_4986);
xnor U6829 (N_6829,N_4582,N_4514);
nor U6830 (N_6830,N_5621,N_5291);
nand U6831 (N_6831,N_4455,N_4357);
and U6832 (N_6832,N_4978,N_4590);
nand U6833 (N_6833,N_5049,N_4054);
and U6834 (N_6834,N_4645,N_4732);
and U6835 (N_6835,N_4558,N_5390);
nand U6836 (N_6836,N_4136,N_5774);
xor U6837 (N_6837,N_5770,N_4755);
nand U6838 (N_6838,N_4632,N_4226);
nor U6839 (N_6839,N_5043,N_5076);
or U6840 (N_6840,N_4878,N_4073);
and U6841 (N_6841,N_5134,N_4617);
nand U6842 (N_6842,N_5761,N_4010);
and U6843 (N_6843,N_5986,N_4736);
nor U6844 (N_6844,N_4207,N_5445);
nand U6845 (N_6845,N_4726,N_4429);
nand U6846 (N_6846,N_4837,N_5133);
xor U6847 (N_6847,N_4397,N_4106);
nand U6848 (N_6848,N_4182,N_4916);
nand U6849 (N_6849,N_5349,N_5325);
or U6850 (N_6850,N_4526,N_4973);
nor U6851 (N_6851,N_5547,N_4901);
and U6852 (N_6852,N_5145,N_5557);
xnor U6853 (N_6853,N_5182,N_5239);
and U6854 (N_6854,N_4600,N_4288);
or U6855 (N_6855,N_5675,N_4257);
and U6856 (N_6856,N_4616,N_5753);
nand U6857 (N_6857,N_4069,N_4148);
nor U6858 (N_6858,N_5718,N_4572);
and U6859 (N_6859,N_5247,N_4283);
or U6860 (N_6860,N_5648,N_4744);
or U6861 (N_6861,N_5810,N_4802);
nor U6862 (N_6862,N_5633,N_5928);
nor U6863 (N_6863,N_4635,N_4342);
nand U6864 (N_6864,N_4407,N_5292);
nor U6865 (N_6865,N_4684,N_4664);
nand U6866 (N_6866,N_5815,N_4983);
nand U6867 (N_6867,N_4839,N_5211);
and U6868 (N_6868,N_5957,N_4700);
or U6869 (N_6869,N_4124,N_5911);
xnor U6870 (N_6870,N_4852,N_5866);
nand U6871 (N_6871,N_5214,N_5775);
or U6872 (N_6872,N_5782,N_4306);
nand U6873 (N_6873,N_4659,N_5746);
or U6874 (N_6874,N_4219,N_4512);
or U6875 (N_6875,N_4548,N_4794);
and U6876 (N_6876,N_5095,N_4889);
nand U6877 (N_6877,N_5482,N_4965);
nand U6878 (N_6878,N_4502,N_5069);
nand U6879 (N_6879,N_4836,N_5838);
or U6880 (N_6880,N_5739,N_4028);
nand U6881 (N_6881,N_4059,N_4467);
nand U6882 (N_6882,N_5893,N_4139);
nor U6883 (N_6883,N_5561,N_5907);
nor U6884 (N_6884,N_5337,N_5030);
nor U6885 (N_6885,N_5834,N_5039);
or U6886 (N_6886,N_4093,N_4618);
nor U6887 (N_6887,N_4464,N_4300);
and U6888 (N_6888,N_4584,N_5321);
nand U6889 (N_6889,N_4414,N_5307);
nor U6890 (N_6890,N_5461,N_4835);
and U6891 (N_6891,N_4885,N_4375);
and U6892 (N_6892,N_5171,N_4461);
and U6893 (N_6893,N_5639,N_5010);
nand U6894 (N_6894,N_4242,N_4758);
xor U6895 (N_6895,N_5918,N_5754);
and U6896 (N_6896,N_4781,N_4258);
or U6897 (N_6897,N_5487,N_5552);
nand U6898 (N_6898,N_5162,N_4951);
and U6899 (N_6899,N_5665,N_5354);
and U6900 (N_6900,N_5993,N_4348);
or U6901 (N_6901,N_5293,N_5339);
or U6902 (N_6902,N_4695,N_4320);
or U6903 (N_6903,N_5027,N_5372);
and U6904 (N_6904,N_4102,N_4243);
nand U6905 (N_6905,N_5980,N_5803);
or U6906 (N_6906,N_4197,N_4545);
and U6907 (N_6907,N_4941,N_4509);
nand U6908 (N_6908,N_5680,N_5169);
and U6909 (N_6909,N_4623,N_5058);
or U6910 (N_6910,N_4416,N_5340);
or U6911 (N_6911,N_5250,N_4860);
or U6912 (N_6912,N_5358,N_4232);
or U6913 (N_6913,N_4045,N_4761);
nor U6914 (N_6914,N_4807,N_5987);
and U6915 (N_6915,N_4667,N_5294);
xnor U6916 (N_6916,N_4369,N_4364);
nor U6917 (N_6917,N_5157,N_5527);
nor U6918 (N_6918,N_5936,N_4255);
or U6919 (N_6919,N_5691,N_4662);
and U6920 (N_6920,N_4699,N_4008);
nand U6921 (N_6921,N_5420,N_4168);
and U6922 (N_6922,N_5791,N_4991);
and U6923 (N_6923,N_4981,N_5599);
or U6924 (N_6924,N_4297,N_5208);
nand U6925 (N_6925,N_5848,N_4650);
nor U6926 (N_6926,N_5745,N_4938);
nand U6927 (N_6927,N_5802,N_4806);
nand U6928 (N_6928,N_4647,N_5172);
and U6929 (N_6929,N_5201,N_5268);
nor U6930 (N_6930,N_4120,N_5215);
and U6931 (N_6931,N_4267,N_5156);
nand U6932 (N_6932,N_4192,N_4859);
nand U6933 (N_6933,N_4385,N_5930);
nand U6934 (N_6934,N_4186,N_5392);
nor U6935 (N_6935,N_5413,N_5310);
nor U6936 (N_6936,N_4709,N_4234);
or U6937 (N_6937,N_4944,N_4305);
or U6938 (N_6938,N_4886,N_4366);
and U6939 (N_6939,N_5610,N_5018);
or U6940 (N_6940,N_5950,N_5436);
and U6941 (N_6941,N_4984,N_4822);
and U6942 (N_6942,N_4451,N_5185);
or U6943 (N_6943,N_5355,N_4043);
nor U6944 (N_6944,N_5350,N_4798);
nor U6945 (N_6945,N_5079,N_5735);
nor U6946 (N_6946,N_5968,N_5297);
and U6947 (N_6947,N_4789,N_4723);
and U6948 (N_6948,N_4595,N_5808);
nor U6949 (N_6949,N_4175,N_5047);
nand U6950 (N_6950,N_5013,N_5352);
and U6951 (N_6951,N_5916,N_4643);
nand U6952 (N_6952,N_4591,N_5324);
and U6953 (N_6953,N_5817,N_5377);
and U6954 (N_6954,N_5168,N_4453);
nand U6955 (N_6955,N_4314,N_5284);
and U6956 (N_6956,N_4930,N_4663);
nor U6957 (N_6957,N_5060,N_4853);
or U6958 (N_6958,N_4143,N_5112);
nor U6959 (N_6959,N_4060,N_5909);
nand U6960 (N_6960,N_5213,N_5068);
or U6961 (N_6961,N_4546,N_4932);
nor U6962 (N_6962,N_4312,N_5180);
nand U6963 (N_6963,N_4864,N_5764);
and U6964 (N_6964,N_5843,N_5166);
or U6965 (N_6965,N_5237,N_5520);
and U6966 (N_6966,N_4592,N_4920);
nor U6967 (N_6967,N_4782,N_5759);
or U6968 (N_6968,N_4123,N_4131);
nor U6969 (N_6969,N_4898,N_4404);
or U6970 (N_6970,N_4337,N_4233);
nand U6971 (N_6971,N_4066,N_5369);
nor U6972 (N_6972,N_4265,N_4355);
or U6973 (N_6973,N_5565,N_4160);
xor U6974 (N_6974,N_5364,N_4221);
and U6975 (N_6975,N_5229,N_5623);
and U6976 (N_6976,N_5025,N_5493);
nand U6977 (N_6977,N_4217,N_5693);
or U6978 (N_6978,N_4095,N_5788);
xnor U6979 (N_6979,N_5263,N_5771);
and U6980 (N_6980,N_4137,N_4954);
and U6981 (N_6981,N_4178,N_4655);
nor U6982 (N_6982,N_5470,N_4906);
nor U6983 (N_6983,N_4865,N_5346);
or U6984 (N_6984,N_5960,N_5744);
nor U6985 (N_6985,N_4754,N_4285);
or U6986 (N_6986,N_5235,N_4076);
nor U6987 (N_6987,N_5136,N_4883);
and U6988 (N_6988,N_5483,N_5406);
or U6989 (N_6989,N_5919,N_5574);
nor U6990 (N_6990,N_5444,N_4361);
and U6991 (N_6991,N_5189,N_4049);
nor U6992 (N_6992,N_4282,N_4262);
and U6993 (N_6993,N_5197,N_4037);
and U6994 (N_6994,N_5072,N_4975);
or U6995 (N_6995,N_5798,N_4315);
nand U6996 (N_6996,N_5052,N_5016);
nor U6997 (N_6997,N_5270,N_5448);
or U6998 (N_6998,N_4302,N_4241);
or U6999 (N_6999,N_5629,N_5402);
nor U7000 (N_7000,N_4768,N_5886);
nor U7001 (N_7001,N_4244,N_4729);
nor U7002 (N_7002,N_4909,N_4124);
nor U7003 (N_7003,N_5643,N_4495);
nand U7004 (N_7004,N_5175,N_5664);
and U7005 (N_7005,N_4973,N_4851);
or U7006 (N_7006,N_4659,N_5877);
and U7007 (N_7007,N_4581,N_5679);
nand U7008 (N_7008,N_4501,N_5277);
nor U7009 (N_7009,N_5043,N_4303);
or U7010 (N_7010,N_5474,N_4874);
or U7011 (N_7011,N_5557,N_4339);
or U7012 (N_7012,N_4460,N_4659);
nand U7013 (N_7013,N_4327,N_5332);
nand U7014 (N_7014,N_4202,N_5031);
nand U7015 (N_7015,N_4035,N_4236);
or U7016 (N_7016,N_4272,N_5483);
and U7017 (N_7017,N_4030,N_5781);
nand U7018 (N_7018,N_5941,N_5354);
or U7019 (N_7019,N_5135,N_5263);
nor U7020 (N_7020,N_4133,N_4472);
or U7021 (N_7021,N_4730,N_5869);
nand U7022 (N_7022,N_5582,N_5557);
nor U7023 (N_7023,N_5224,N_4748);
nand U7024 (N_7024,N_4430,N_4327);
and U7025 (N_7025,N_5466,N_4457);
nor U7026 (N_7026,N_4873,N_5027);
and U7027 (N_7027,N_4610,N_4871);
xnor U7028 (N_7028,N_4301,N_4035);
nor U7029 (N_7029,N_4541,N_5543);
or U7030 (N_7030,N_5842,N_4096);
and U7031 (N_7031,N_4945,N_5048);
nand U7032 (N_7032,N_4114,N_4260);
xor U7033 (N_7033,N_5362,N_5104);
or U7034 (N_7034,N_4937,N_4216);
or U7035 (N_7035,N_5750,N_4864);
nor U7036 (N_7036,N_5586,N_4878);
nand U7037 (N_7037,N_5747,N_5590);
and U7038 (N_7038,N_5927,N_4581);
or U7039 (N_7039,N_5604,N_5207);
or U7040 (N_7040,N_5323,N_5816);
nand U7041 (N_7041,N_4582,N_5131);
nand U7042 (N_7042,N_5213,N_4472);
and U7043 (N_7043,N_4030,N_4665);
or U7044 (N_7044,N_5115,N_5505);
nor U7045 (N_7045,N_4347,N_5490);
or U7046 (N_7046,N_5827,N_5586);
or U7047 (N_7047,N_4314,N_5409);
nand U7048 (N_7048,N_4738,N_5228);
and U7049 (N_7049,N_4454,N_4023);
nor U7050 (N_7050,N_4693,N_4788);
nand U7051 (N_7051,N_4500,N_4052);
nand U7052 (N_7052,N_5382,N_4892);
nand U7053 (N_7053,N_4482,N_5206);
nand U7054 (N_7054,N_5281,N_5935);
and U7055 (N_7055,N_5732,N_4223);
or U7056 (N_7056,N_4906,N_4938);
nor U7057 (N_7057,N_5333,N_5612);
nand U7058 (N_7058,N_4503,N_4398);
nand U7059 (N_7059,N_5574,N_5323);
and U7060 (N_7060,N_4362,N_5992);
or U7061 (N_7061,N_4795,N_4739);
nor U7062 (N_7062,N_5840,N_5242);
nand U7063 (N_7063,N_5358,N_5348);
and U7064 (N_7064,N_5666,N_5889);
nor U7065 (N_7065,N_5131,N_4363);
nand U7066 (N_7066,N_5267,N_4804);
and U7067 (N_7067,N_4701,N_4939);
or U7068 (N_7068,N_5416,N_5517);
or U7069 (N_7069,N_4917,N_5836);
and U7070 (N_7070,N_4449,N_5187);
nor U7071 (N_7071,N_4677,N_5633);
and U7072 (N_7072,N_5561,N_4362);
nand U7073 (N_7073,N_5584,N_5856);
and U7074 (N_7074,N_4771,N_5925);
or U7075 (N_7075,N_4588,N_4784);
and U7076 (N_7076,N_5791,N_4228);
nand U7077 (N_7077,N_5387,N_5076);
or U7078 (N_7078,N_5262,N_5118);
and U7079 (N_7079,N_5488,N_5451);
nand U7080 (N_7080,N_5301,N_4010);
or U7081 (N_7081,N_4504,N_5179);
nand U7082 (N_7082,N_5331,N_4827);
and U7083 (N_7083,N_4533,N_4377);
or U7084 (N_7084,N_4747,N_4158);
xnor U7085 (N_7085,N_5024,N_4331);
nand U7086 (N_7086,N_4461,N_4814);
nor U7087 (N_7087,N_4345,N_5632);
and U7088 (N_7088,N_4047,N_5039);
nor U7089 (N_7089,N_4757,N_4596);
and U7090 (N_7090,N_4994,N_5913);
or U7091 (N_7091,N_4977,N_4305);
nand U7092 (N_7092,N_5117,N_4586);
nand U7093 (N_7093,N_5845,N_5660);
nand U7094 (N_7094,N_4031,N_4379);
nor U7095 (N_7095,N_4795,N_4120);
xnor U7096 (N_7096,N_4354,N_5702);
nand U7097 (N_7097,N_5195,N_4773);
and U7098 (N_7098,N_5091,N_4325);
or U7099 (N_7099,N_4341,N_4466);
nor U7100 (N_7100,N_4845,N_4850);
nand U7101 (N_7101,N_5039,N_4852);
and U7102 (N_7102,N_5455,N_4689);
or U7103 (N_7103,N_4954,N_5151);
nor U7104 (N_7104,N_4085,N_4016);
nor U7105 (N_7105,N_5259,N_4846);
nor U7106 (N_7106,N_5108,N_5034);
nand U7107 (N_7107,N_5814,N_5641);
and U7108 (N_7108,N_4047,N_5086);
or U7109 (N_7109,N_5322,N_4275);
and U7110 (N_7110,N_5690,N_5072);
and U7111 (N_7111,N_4887,N_4682);
or U7112 (N_7112,N_4842,N_4292);
nand U7113 (N_7113,N_4936,N_5610);
xnor U7114 (N_7114,N_4247,N_5894);
nor U7115 (N_7115,N_5614,N_4699);
nor U7116 (N_7116,N_5248,N_5643);
and U7117 (N_7117,N_5622,N_5424);
and U7118 (N_7118,N_4506,N_4234);
and U7119 (N_7119,N_5497,N_5584);
or U7120 (N_7120,N_5588,N_4959);
nor U7121 (N_7121,N_5632,N_4129);
or U7122 (N_7122,N_5019,N_5205);
xor U7123 (N_7123,N_4837,N_4057);
nand U7124 (N_7124,N_4608,N_5859);
or U7125 (N_7125,N_5836,N_4301);
xnor U7126 (N_7126,N_4665,N_5755);
nor U7127 (N_7127,N_4990,N_5200);
nand U7128 (N_7128,N_4625,N_5205);
and U7129 (N_7129,N_5252,N_4628);
and U7130 (N_7130,N_4605,N_4434);
nand U7131 (N_7131,N_5997,N_4748);
and U7132 (N_7132,N_5645,N_5658);
and U7133 (N_7133,N_4994,N_5940);
nor U7134 (N_7134,N_4020,N_5229);
and U7135 (N_7135,N_4228,N_5740);
and U7136 (N_7136,N_5911,N_5585);
nor U7137 (N_7137,N_5190,N_4783);
nor U7138 (N_7138,N_5926,N_5108);
nor U7139 (N_7139,N_5274,N_4044);
nand U7140 (N_7140,N_4929,N_4278);
nand U7141 (N_7141,N_5201,N_4108);
nand U7142 (N_7142,N_5205,N_5095);
nand U7143 (N_7143,N_4169,N_4664);
nand U7144 (N_7144,N_5281,N_5030);
xor U7145 (N_7145,N_5214,N_4947);
and U7146 (N_7146,N_5547,N_5203);
and U7147 (N_7147,N_4318,N_4734);
and U7148 (N_7148,N_4279,N_5314);
nand U7149 (N_7149,N_5026,N_5401);
and U7150 (N_7150,N_4048,N_5033);
and U7151 (N_7151,N_4492,N_5139);
xor U7152 (N_7152,N_4537,N_5759);
and U7153 (N_7153,N_4327,N_4061);
or U7154 (N_7154,N_5205,N_5553);
nor U7155 (N_7155,N_4633,N_5467);
nor U7156 (N_7156,N_5553,N_4546);
and U7157 (N_7157,N_5570,N_4917);
nor U7158 (N_7158,N_4361,N_4965);
xnor U7159 (N_7159,N_5192,N_4878);
nand U7160 (N_7160,N_5337,N_5144);
and U7161 (N_7161,N_4491,N_4801);
nor U7162 (N_7162,N_5197,N_5702);
nand U7163 (N_7163,N_5706,N_4176);
or U7164 (N_7164,N_5438,N_5683);
and U7165 (N_7165,N_4511,N_5305);
xor U7166 (N_7166,N_5130,N_5792);
and U7167 (N_7167,N_4095,N_4554);
nand U7168 (N_7168,N_5308,N_4635);
nor U7169 (N_7169,N_4764,N_5388);
or U7170 (N_7170,N_5930,N_5724);
or U7171 (N_7171,N_4742,N_5471);
nand U7172 (N_7172,N_5001,N_4721);
nand U7173 (N_7173,N_5353,N_5543);
nand U7174 (N_7174,N_4936,N_5115);
or U7175 (N_7175,N_4868,N_4141);
nor U7176 (N_7176,N_5036,N_4841);
or U7177 (N_7177,N_4304,N_5964);
or U7178 (N_7178,N_4718,N_5133);
and U7179 (N_7179,N_4234,N_5036);
nand U7180 (N_7180,N_5558,N_4486);
and U7181 (N_7181,N_4553,N_4456);
xnor U7182 (N_7182,N_4917,N_5954);
nand U7183 (N_7183,N_4358,N_4691);
nor U7184 (N_7184,N_5811,N_5682);
nor U7185 (N_7185,N_4972,N_4913);
and U7186 (N_7186,N_5250,N_5374);
or U7187 (N_7187,N_5724,N_4104);
nand U7188 (N_7188,N_4722,N_4204);
nor U7189 (N_7189,N_5633,N_5784);
nor U7190 (N_7190,N_4229,N_5060);
and U7191 (N_7191,N_4348,N_5002);
nor U7192 (N_7192,N_4518,N_5102);
nor U7193 (N_7193,N_5653,N_4917);
nand U7194 (N_7194,N_5864,N_4124);
and U7195 (N_7195,N_4041,N_4573);
nor U7196 (N_7196,N_4512,N_5757);
or U7197 (N_7197,N_4859,N_5288);
nand U7198 (N_7198,N_5361,N_5166);
nand U7199 (N_7199,N_5204,N_5286);
or U7200 (N_7200,N_5928,N_5520);
or U7201 (N_7201,N_4564,N_5115);
and U7202 (N_7202,N_4498,N_4634);
nor U7203 (N_7203,N_5981,N_5842);
and U7204 (N_7204,N_5826,N_5869);
or U7205 (N_7205,N_5656,N_4944);
nor U7206 (N_7206,N_4383,N_5943);
nor U7207 (N_7207,N_4615,N_4710);
or U7208 (N_7208,N_4255,N_4715);
and U7209 (N_7209,N_4527,N_4561);
nor U7210 (N_7210,N_4987,N_5080);
nand U7211 (N_7211,N_4519,N_4427);
and U7212 (N_7212,N_5613,N_5070);
nand U7213 (N_7213,N_4522,N_4105);
nand U7214 (N_7214,N_5699,N_4899);
and U7215 (N_7215,N_5738,N_5807);
or U7216 (N_7216,N_4927,N_4745);
nand U7217 (N_7217,N_5485,N_4653);
or U7218 (N_7218,N_4125,N_4130);
nand U7219 (N_7219,N_4347,N_4988);
nand U7220 (N_7220,N_5580,N_5009);
and U7221 (N_7221,N_5742,N_4874);
nand U7222 (N_7222,N_4801,N_4233);
and U7223 (N_7223,N_5219,N_5927);
and U7224 (N_7224,N_4452,N_4832);
nor U7225 (N_7225,N_5230,N_4622);
or U7226 (N_7226,N_4248,N_4387);
nor U7227 (N_7227,N_5026,N_4256);
nor U7228 (N_7228,N_4236,N_5962);
nand U7229 (N_7229,N_5473,N_4766);
xnor U7230 (N_7230,N_4008,N_5972);
or U7231 (N_7231,N_5738,N_5098);
or U7232 (N_7232,N_5316,N_4311);
or U7233 (N_7233,N_5371,N_4155);
and U7234 (N_7234,N_5332,N_5492);
or U7235 (N_7235,N_5056,N_4581);
nor U7236 (N_7236,N_5818,N_5982);
or U7237 (N_7237,N_4247,N_4194);
or U7238 (N_7238,N_4039,N_4634);
nor U7239 (N_7239,N_4169,N_4958);
or U7240 (N_7240,N_5381,N_5651);
or U7241 (N_7241,N_4603,N_4340);
nor U7242 (N_7242,N_4180,N_4647);
nand U7243 (N_7243,N_5975,N_5512);
or U7244 (N_7244,N_4474,N_5424);
xnor U7245 (N_7245,N_5158,N_5739);
xnor U7246 (N_7246,N_5681,N_5095);
nand U7247 (N_7247,N_4371,N_4165);
nor U7248 (N_7248,N_5136,N_5241);
and U7249 (N_7249,N_4136,N_4350);
or U7250 (N_7250,N_4473,N_5640);
nor U7251 (N_7251,N_4620,N_4062);
xnor U7252 (N_7252,N_4139,N_4196);
nand U7253 (N_7253,N_5592,N_5515);
or U7254 (N_7254,N_5983,N_5324);
nand U7255 (N_7255,N_5837,N_4711);
nand U7256 (N_7256,N_5663,N_4850);
nand U7257 (N_7257,N_4896,N_4211);
and U7258 (N_7258,N_4318,N_5045);
nor U7259 (N_7259,N_4067,N_5421);
nand U7260 (N_7260,N_4952,N_5608);
or U7261 (N_7261,N_4546,N_5845);
and U7262 (N_7262,N_4362,N_4535);
or U7263 (N_7263,N_4144,N_5321);
nor U7264 (N_7264,N_4914,N_5159);
nor U7265 (N_7265,N_5291,N_4951);
nor U7266 (N_7266,N_4513,N_4774);
nor U7267 (N_7267,N_4439,N_5884);
nand U7268 (N_7268,N_4740,N_4486);
or U7269 (N_7269,N_4034,N_4437);
or U7270 (N_7270,N_5512,N_4024);
nand U7271 (N_7271,N_4237,N_4515);
and U7272 (N_7272,N_5514,N_4971);
and U7273 (N_7273,N_4928,N_4106);
or U7274 (N_7274,N_4750,N_4124);
nor U7275 (N_7275,N_4223,N_5907);
nor U7276 (N_7276,N_5235,N_5779);
and U7277 (N_7277,N_5497,N_4803);
and U7278 (N_7278,N_4779,N_4096);
nor U7279 (N_7279,N_5545,N_4931);
or U7280 (N_7280,N_4647,N_4161);
nand U7281 (N_7281,N_4292,N_4486);
nand U7282 (N_7282,N_4547,N_5987);
and U7283 (N_7283,N_5186,N_5754);
nand U7284 (N_7284,N_5146,N_5070);
nor U7285 (N_7285,N_4486,N_5857);
and U7286 (N_7286,N_5135,N_5847);
or U7287 (N_7287,N_4839,N_5698);
and U7288 (N_7288,N_5509,N_5935);
nor U7289 (N_7289,N_4499,N_4011);
or U7290 (N_7290,N_4447,N_5605);
nand U7291 (N_7291,N_4406,N_5710);
or U7292 (N_7292,N_4654,N_5191);
and U7293 (N_7293,N_4306,N_5644);
or U7294 (N_7294,N_5651,N_4675);
and U7295 (N_7295,N_4807,N_4069);
or U7296 (N_7296,N_4906,N_4398);
nor U7297 (N_7297,N_5998,N_4846);
nor U7298 (N_7298,N_5189,N_5455);
and U7299 (N_7299,N_5830,N_4079);
nand U7300 (N_7300,N_5415,N_5330);
or U7301 (N_7301,N_4034,N_5722);
nand U7302 (N_7302,N_5780,N_4434);
and U7303 (N_7303,N_4296,N_4649);
or U7304 (N_7304,N_4128,N_5640);
or U7305 (N_7305,N_5520,N_4212);
xnor U7306 (N_7306,N_5599,N_5372);
or U7307 (N_7307,N_5459,N_4276);
nor U7308 (N_7308,N_5280,N_4880);
nor U7309 (N_7309,N_4523,N_4941);
or U7310 (N_7310,N_4239,N_4629);
or U7311 (N_7311,N_5219,N_5672);
nand U7312 (N_7312,N_4649,N_5607);
or U7313 (N_7313,N_5010,N_5187);
nand U7314 (N_7314,N_4628,N_4995);
and U7315 (N_7315,N_4211,N_4875);
xnor U7316 (N_7316,N_4857,N_4234);
or U7317 (N_7317,N_4010,N_4100);
nand U7318 (N_7318,N_4623,N_5712);
or U7319 (N_7319,N_5311,N_4216);
or U7320 (N_7320,N_4158,N_4778);
nor U7321 (N_7321,N_4060,N_5823);
nand U7322 (N_7322,N_4825,N_5409);
nand U7323 (N_7323,N_5494,N_5197);
or U7324 (N_7324,N_5650,N_4670);
or U7325 (N_7325,N_4575,N_4934);
nand U7326 (N_7326,N_5658,N_4676);
or U7327 (N_7327,N_5457,N_5835);
and U7328 (N_7328,N_5128,N_5454);
and U7329 (N_7329,N_5881,N_5784);
nand U7330 (N_7330,N_5666,N_5493);
nor U7331 (N_7331,N_5937,N_4352);
nor U7332 (N_7332,N_4481,N_4147);
and U7333 (N_7333,N_5952,N_4644);
nor U7334 (N_7334,N_5271,N_5330);
and U7335 (N_7335,N_5145,N_4443);
nor U7336 (N_7336,N_4112,N_5179);
or U7337 (N_7337,N_4571,N_5551);
or U7338 (N_7338,N_4034,N_5139);
or U7339 (N_7339,N_5319,N_5332);
and U7340 (N_7340,N_4140,N_4130);
or U7341 (N_7341,N_4014,N_4900);
nand U7342 (N_7342,N_5193,N_4972);
nor U7343 (N_7343,N_4474,N_5078);
nand U7344 (N_7344,N_4340,N_5294);
nand U7345 (N_7345,N_5917,N_4371);
or U7346 (N_7346,N_5225,N_5160);
or U7347 (N_7347,N_4278,N_4991);
and U7348 (N_7348,N_5011,N_5047);
nor U7349 (N_7349,N_5093,N_4469);
nor U7350 (N_7350,N_4081,N_4026);
nand U7351 (N_7351,N_4511,N_5367);
or U7352 (N_7352,N_5961,N_5244);
and U7353 (N_7353,N_5120,N_5267);
and U7354 (N_7354,N_5290,N_4067);
or U7355 (N_7355,N_5337,N_5958);
or U7356 (N_7356,N_5380,N_5323);
or U7357 (N_7357,N_5026,N_4988);
or U7358 (N_7358,N_4186,N_5457);
nor U7359 (N_7359,N_4196,N_5566);
or U7360 (N_7360,N_5500,N_5825);
nand U7361 (N_7361,N_5191,N_4963);
nand U7362 (N_7362,N_5991,N_4824);
nor U7363 (N_7363,N_5502,N_5951);
nor U7364 (N_7364,N_4530,N_5338);
nand U7365 (N_7365,N_4951,N_5903);
nand U7366 (N_7366,N_4847,N_5642);
nand U7367 (N_7367,N_4186,N_5900);
nor U7368 (N_7368,N_4107,N_5698);
nor U7369 (N_7369,N_4976,N_5063);
nand U7370 (N_7370,N_5343,N_4872);
and U7371 (N_7371,N_5727,N_5494);
xor U7372 (N_7372,N_5881,N_4975);
and U7373 (N_7373,N_4287,N_5615);
or U7374 (N_7374,N_4834,N_5126);
nand U7375 (N_7375,N_5528,N_4525);
nor U7376 (N_7376,N_5905,N_5090);
and U7377 (N_7377,N_4333,N_4398);
and U7378 (N_7378,N_5048,N_5999);
nand U7379 (N_7379,N_4756,N_4915);
or U7380 (N_7380,N_4276,N_5856);
nor U7381 (N_7381,N_4417,N_4904);
and U7382 (N_7382,N_5643,N_5713);
or U7383 (N_7383,N_5807,N_4881);
and U7384 (N_7384,N_4696,N_4165);
nand U7385 (N_7385,N_4660,N_4675);
or U7386 (N_7386,N_4164,N_4268);
nand U7387 (N_7387,N_4184,N_4862);
or U7388 (N_7388,N_5350,N_5990);
or U7389 (N_7389,N_5912,N_5503);
nor U7390 (N_7390,N_5994,N_4600);
nor U7391 (N_7391,N_4298,N_4457);
nor U7392 (N_7392,N_4018,N_4522);
and U7393 (N_7393,N_4571,N_4079);
and U7394 (N_7394,N_4119,N_5205);
and U7395 (N_7395,N_5355,N_5406);
nand U7396 (N_7396,N_4169,N_5918);
nor U7397 (N_7397,N_4738,N_4545);
nor U7398 (N_7398,N_4197,N_4216);
and U7399 (N_7399,N_4381,N_4685);
nand U7400 (N_7400,N_4089,N_4194);
and U7401 (N_7401,N_5514,N_4225);
or U7402 (N_7402,N_4030,N_5139);
nor U7403 (N_7403,N_4561,N_5970);
nand U7404 (N_7404,N_4921,N_4853);
and U7405 (N_7405,N_5272,N_5589);
and U7406 (N_7406,N_5438,N_5131);
and U7407 (N_7407,N_5409,N_5872);
nor U7408 (N_7408,N_5670,N_5143);
and U7409 (N_7409,N_5177,N_4101);
and U7410 (N_7410,N_5333,N_4319);
nand U7411 (N_7411,N_4790,N_4391);
and U7412 (N_7412,N_4126,N_4524);
or U7413 (N_7413,N_5393,N_4726);
or U7414 (N_7414,N_4339,N_5335);
nor U7415 (N_7415,N_4808,N_5305);
nand U7416 (N_7416,N_4749,N_4147);
or U7417 (N_7417,N_5441,N_4870);
xnor U7418 (N_7418,N_4377,N_4126);
and U7419 (N_7419,N_5636,N_5084);
xnor U7420 (N_7420,N_4695,N_4223);
and U7421 (N_7421,N_4730,N_4336);
nand U7422 (N_7422,N_5047,N_4210);
and U7423 (N_7423,N_5451,N_4609);
nor U7424 (N_7424,N_4365,N_5911);
and U7425 (N_7425,N_5034,N_4233);
nand U7426 (N_7426,N_5295,N_5094);
and U7427 (N_7427,N_5333,N_4920);
nand U7428 (N_7428,N_4921,N_4109);
nand U7429 (N_7429,N_4347,N_5546);
nand U7430 (N_7430,N_5914,N_4848);
xor U7431 (N_7431,N_5321,N_4120);
and U7432 (N_7432,N_4394,N_4064);
nand U7433 (N_7433,N_4656,N_5409);
or U7434 (N_7434,N_4645,N_5080);
nor U7435 (N_7435,N_4881,N_4528);
nand U7436 (N_7436,N_5934,N_4881);
nor U7437 (N_7437,N_5128,N_5134);
nand U7438 (N_7438,N_4936,N_4287);
nand U7439 (N_7439,N_4378,N_4522);
or U7440 (N_7440,N_4512,N_4348);
nand U7441 (N_7441,N_4813,N_4392);
nor U7442 (N_7442,N_5057,N_5749);
nor U7443 (N_7443,N_4773,N_5332);
nor U7444 (N_7444,N_4155,N_4032);
or U7445 (N_7445,N_5860,N_5836);
nor U7446 (N_7446,N_5738,N_5737);
or U7447 (N_7447,N_5969,N_5448);
nand U7448 (N_7448,N_5201,N_4760);
or U7449 (N_7449,N_4932,N_4198);
and U7450 (N_7450,N_4625,N_5117);
nor U7451 (N_7451,N_4646,N_4435);
nand U7452 (N_7452,N_5578,N_5111);
or U7453 (N_7453,N_4124,N_5508);
or U7454 (N_7454,N_4221,N_4665);
nor U7455 (N_7455,N_5493,N_5264);
nand U7456 (N_7456,N_4280,N_5521);
nand U7457 (N_7457,N_5729,N_4741);
xor U7458 (N_7458,N_4814,N_5504);
and U7459 (N_7459,N_5340,N_4805);
and U7460 (N_7460,N_5026,N_5587);
or U7461 (N_7461,N_5414,N_5295);
or U7462 (N_7462,N_4936,N_5405);
and U7463 (N_7463,N_4392,N_5893);
nor U7464 (N_7464,N_4031,N_5509);
xnor U7465 (N_7465,N_5074,N_4686);
or U7466 (N_7466,N_4949,N_4767);
nand U7467 (N_7467,N_5669,N_5716);
nor U7468 (N_7468,N_5449,N_5567);
nor U7469 (N_7469,N_5167,N_4275);
nor U7470 (N_7470,N_4889,N_4215);
or U7471 (N_7471,N_5019,N_4525);
or U7472 (N_7472,N_4298,N_5402);
xor U7473 (N_7473,N_5004,N_4550);
nand U7474 (N_7474,N_5640,N_4454);
nand U7475 (N_7475,N_4593,N_5100);
and U7476 (N_7476,N_4131,N_5315);
nand U7477 (N_7477,N_4963,N_5170);
nor U7478 (N_7478,N_5905,N_5351);
or U7479 (N_7479,N_5631,N_4774);
and U7480 (N_7480,N_5973,N_4980);
nand U7481 (N_7481,N_5354,N_4598);
nor U7482 (N_7482,N_5552,N_4848);
nor U7483 (N_7483,N_5312,N_4926);
or U7484 (N_7484,N_4498,N_4660);
nor U7485 (N_7485,N_5448,N_4802);
xor U7486 (N_7486,N_5870,N_5344);
nor U7487 (N_7487,N_4193,N_4247);
and U7488 (N_7488,N_4975,N_4751);
nand U7489 (N_7489,N_5131,N_4839);
nand U7490 (N_7490,N_4685,N_4256);
or U7491 (N_7491,N_4861,N_5575);
or U7492 (N_7492,N_5441,N_4936);
or U7493 (N_7493,N_5667,N_4323);
nand U7494 (N_7494,N_5070,N_4253);
or U7495 (N_7495,N_5510,N_4326);
or U7496 (N_7496,N_4464,N_4293);
nand U7497 (N_7497,N_5833,N_4700);
nor U7498 (N_7498,N_4951,N_5348);
nand U7499 (N_7499,N_4271,N_4202);
nor U7500 (N_7500,N_4876,N_4572);
and U7501 (N_7501,N_4129,N_5745);
and U7502 (N_7502,N_5233,N_4229);
or U7503 (N_7503,N_5034,N_5561);
nand U7504 (N_7504,N_4755,N_5538);
or U7505 (N_7505,N_5421,N_4455);
nand U7506 (N_7506,N_4815,N_4652);
and U7507 (N_7507,N_4133,N_4474);
nor U7508 (N_7508,N_4454,N_5330);
or U7509 (N_7509,N_4663,N_5939);
nand U7510 (N_7510,N_4413,N_5118);
nor U7511 (N_7511,N_4249,N_4991);
nand U7512 (N_7512,N_4292,N_4163);
and U7513 (N_7513,N_4717,N_5555);
nand U7514 (N_7514,N_5395,N_5544);
and U7515 (N_7515,N_4700,N_5027);
or U7516 (N_7516,N_5745,N_4822);
or U7517 (N_7517,N_5579,N_4738);
and U7518 (N_7518,N_4717,N_5069);
and U7519 (N_7519,N_5459,N_5827);
nand U7520 (N_7520,N_4262,N_5588);
and U7521 (N_7521,N_5606,N_5299);
nor U7522 (N_7522,N_5947,N_4246);
nor U7523 (N_7523,N_4869,N_5328);
or U7524 (N_7524,N_4468,N_5219);
and U7525 (N_7525,N_5671,N_4501);
nor U7526 (N_7526,N_5848,N_5857);
nand U7527 (N_7527,N_5195,N_4537);
nor U7528 (N_7528,N_5290,N_4214);
nand U7529 (N_7529,N_5906,N_5768);
nor U7530 (N_7530,N_4747,N_5269);
and U7531 (N_7531,N_4469,N_5858);
nor U7532 (N_7532,N_4883,N_4286);
nor U7533 (N_7533,N_5516,N_4620);
nor U7534 (N_7534,N_4209,N_4306);
nand U7535 (N_7535,N_5858,N_4086);
and U7536 (N_7536,N_4506,N_4038);
or U7537 (N_7537,N_4590,N_4356);
and U7538 (N_7538,N_5622,N_4280);
or U7539 (N_7539,N_5573,N_5287);
nor U7540 (N_7540,N_5067,N_4317);
xor U7541 (N_7541,N_5437,N_4206);
and U7542 (N_7542,N_5271,N_4671);
nor U7543 (N_7543,N_5010,N_5510);
or U7544 (N_7544,N_5818,N_5249);
and U7545 (N_7545,N_4632,N_5524);
nand U7546 (N_7546,N_4827,N_4667);
nor U7547 (N_7547,N_4195,N_5216);
or U7548 (N_7548,N_4678,N_4086);
or U7549 (N_7549,N_4948,N_5630);
nand U7550 (N_7550,N_4138,N_4538);
or U7551 (N_7551,N_5719,N_5812);
nor U7552 (N_7552,N_4432,N_4586);
xnor U7553 (N_7553,N_5291,N_5795);
nor U7554 (N_7554,N_4986,N_5437);
nand U7555 (N_7555,N_4908,N_4513);
and U7556 (N_7556,N_5611,N_5488);
or U7557 (N_7557,N_4829,N_5143);
nand U7558 (N_7558,N_4256,N_5465);
nor U7559 (N_7559,N_5365,N_4232);
nor U7560 (N_7560,N_4323,N_5356);
nand U7561 (N_7561,N_5895,N_5215);
or U7562 (N_7562,N_4321,N_4989);
nand U7563 (N_7563,N_5172,N_4164);
nor U7564 (N_7564,N_5538,N_5906);
and U7565 (N_7565,N_5094,N_5291);
and U7566 (N_7566,N_4808,N_4127);
nor U7567 (N_7567,N_5275,N_5660);
nand U7568 (N_7568,N_5094,N_5622);
and U7569 (N_7569,N_5582,N_4952);
and U7570 (N_7570,N_4086,N_4603);
nor U7571 (N_7571,N_5172,N_4348);
or U7572 (N_7572,N_4570,N_4407);
nor U7573 (N_7573,N_4532,N_5390);
and U7574 (N_7574,N_5072,N_5357);
and U7575 (N_7575,N_4174,N_5049);
or U7576 (N_7576,N_4644,N_5526);
nor U7577 (N_7577,N_5792,N_5979);
nor U7578 (N_7578,N_4293,N_4251);
or U7579 (N_7579,N_4195,N_5369);
or U7580 (N_7580,N_4527,N_5802);
nand U7581 (N_7581,N_5849,N_5597);
and U7582 (N_7582,N_5546,N_4960);
nand U7583 (N_7583,N_5692,N_5295);
or U7584 (N_7584,N_5203,N_5349);
nor U7585 (N_7585,N_4250,N_5045);
or U7586 (N_7586,N_5661,N_4420);
and U7587 (N_7587,N_5779,N_5675);
nand U7588 (N_7588,N_4388,N_5741);
nor U7589 (N_7589,N_4106,N_4952);
nand U7590 (N_7590,N_4834,N_5719);
nand U7591 (N_7591,N_4082,N_4122);
nor U7592 (N_7592,N_4211,N_4645);
nand U7593 (N_7593,N_4281,N_5584);
nor U7594 (N_7594,N_5203,N_4109);
nand U7595 (N_7595,N_5353,N_5799);
nor U7596 (N_7596,N_4636,N_5814);
and U7597 (N_7597,N_4755,N_4627);
nor U7598 (N_7598,N_4914,N_4617);
nor U7599 (N_7599,N_4689,N_5707);
and U7600 (N_7600,N_4331,N_5813);
nand U7601 (N_7601,N_4366,N_4590);
and U7602 (N_7602,N_5654,N_4560);
nor U7603 (N_7603,N_5500,N_4195);
nand U7604 (N_7604,N_5461,N_4062);
xnor U7605 (N_7605,N_4822,N_4028);
nand U7606 (N_7606,N_5258,N_5334);
nor U7607 (N_7607,N_4793,N_5695);
or U7608 (N_7608,N_4082,N_5581);
and U7609 (N_7609,N_5831,N_5017);
nor U7610 (N_7610,N_5988,N_4716);
or U7611 (N_7611,N_4336,N_5965);
or U7612 (N_7612,N_4052,N_5252);
and U7613 (N_7613,N_4083,N_4702);
nor U7614 (N_7614,N_4375,N_5424);
or U7615 (N_7615,N_4164,N_4235);
and U7616 (N_7616,N_4255,N_5446);
nor U7617 (N_7617,N_4760,N_4132);
or U7618 (N_7618,N_5602,N_5088);
nand U7619 (N_7619,N_5301,N_5625);
or U7620 (N_7620,N_5329,N_4825);
and U7621 (N_7621,N_5896,N_5182);
nor U7622 (N_7622,N_5216,N_4426);
nand U7623 (N_7623,N_5368,N_5622);
and U7624 (N_7624,N_5933,N_5209);
nor U7625 (N_7625,N_4209,N_5637);
xor U7626 (N_7626,N_5166,N_4548);
or U7627 (N_7627,N_4871,N_5902);
nand U7628 (N_7628,N_4554,N_4882);
or U7629 (N_7629,N_5998,N_4366);
and U7630 (N_7630,N_4217,N_4922);
or U7631 (N_7631,N_5816,N_4785);
nor U7632 (N_7632,N_5111,N_5222);
nand U7633 (N_7633,N_5359,N_4051);
nand U7634 (N_7634,N_4085,N_5641);
and U7635 (N_7635,N_4803,N_4967);
and U7636 (N_7636,N_5895,N_5317);
nor U7637 (N_7637,N_5954,N_4885);
or U7638 (N_7638,N_5660,N_5322);
or U7639 (N_7639,N_5708,N_5322);
and U7640 (N_7640,N_4092,N_5817);
nand U7641 (N_7641,N_4865,N_5689);
nor U7642 (N_7642,N_5545,N_4371);
and U7643 (N_7643,N_4892,N_5350);
nor U7644 (N_7644,N_5964,N_5948);
or U7645 (N_7645,N_4059,N_5591);
nand U7646 (N_7646,N_4611,N_5917);
nand U7647 (N_7647,N_5477,N_4331);
xor U7648 (N_7648,N_5490,N_4633);
or U7649 (N_7649,N_5317,N_4773);
and U7650 (N_7650,N_5149,N_5303);
or U7651 (N_7651,N_5297,N_4942);
nor U7652 (N_7652,N_4357,N_4801);
nand U7653 (N_7653,N_5808,N_4513);
nor U7654 (N_7654,N_5398,N_4309);
nor U7655 (N_7655,N_4033,N_5836);
nor U7656 (N_7656,N_5395,N_5429);
nand U7657 (N_7657,N_5403,N_5598);
nand U7658 (N_7658,N_4080,N_5270);
xor U7659 (N_7659,N_5808,N_4746);
and U7660 (N_7660,N_5885,N_5932);
nand U7661 (N_7661,N_5067,N_5674);
or U7662 (N_7662,N_5214,N_4959);
and U7663 (N_7663,N_4219,N_5065);
nand U7664 (N_7664,N_4089,N_5568);
nand U7665 (N_7665,N_5050,N_4656);
or U7666 (N_7666,N_4721,N_5117);
nand U7667 (N_7667,N_5583,N_4313);
or U7668 (N_7668,N_5310,N_4818);
nor U7669 (N_7669,N_5050,N_4302);
nor U7670 (N_7670,N_4431,N_4366);
nand U7671 (N_7671,N_5506,N_5824);
or U7672 (N_7672,N_5056,N_4206);
nor U7673 (N_7673,N_5216,N_4906);
nand U7674 (N_7674,N_5396,N_4284);
nor U7675 (N_7675,N_4340,N_5769);
and U7676 (N_7676,N_5576,N_4056);
nor U7677 (N_7677,N_5553,N_5282);
or U7678 (N_7678,N_5931,N_5764);
nor U7679 (N_7679,N_4920,N_4575);
or U7680 (N_7680,N_4967,N_4771);
or U7681 (N_7681,N_4035,N_5967);
nor U7682 (N_7682,N_5824,N_4601);
nand U7683 (N_7683,N_5246,N_4108);
nand U7684 (N_7684,N_4334,N_5407);
nand U7685 (N_7685,N_5739,N_5883);
nand U7686 (N_7686,N_4318,N_4612);
and U7687 (N_7687,N_5158,N_5897);
and U7688 (N_7688,N_4145,N_5700);
nor U7689 (N_7689,N_4394,N_5604);
and U7690 (N_7690,N_5929,N_4859);
and U7691 (N_7691,N_5582,N_5564);
nand U7692 (N_7692,N_4668,N_4787);
nand U7693 (N_7693,N_5966,N_4457);
or U7694 (N_7694,N_5667,N_4061);
nor U7695 (N_7695,N_4533,N_5214);
and U7696 (N_7696,N_4912,N_5690);
nor U7697 (N_7697,N_4620,N_5087);
or U7698 (N_7698,N_5588,N_5561);
or U7699 (N_7699,N_4934,N_5131);
nand U7700 (N_7700,N_4157,N_4319);
nand U7701 (N_7701,N_4934,N_5204);
nor U7702 (N_7702,N_5309,N_5685);
or U7703 (N_7703,N_5878,N_5648);
and U7704 (N_7704,N_5794,N_4340);
and U7705 (N_7705,N_5869,N_4754);
or U7706 (N_7706,N_4302,N_4018);
nand U7707 (N_7707,N_5497,N_5317);
nor U7708 (N_7708,N_4765,N_5506);
nand U7709 (N_7709,N_5198,N_4655);
nor U7710 (N_7710,N_5612,N_4231);
and U7711 (N_7711,N_4033,N_4615);
nand U7712 (N_7712,N_5509,N_4729);
nor U7713 (N_7713,N_4834,N_5593);
or U7714 (N_7714,N_4319,N_5503);
or U7715 (N_7715,N_5923,N_4323);
and U7716 (N_7716,N_4523,N_5974);
or U7717 (N_7717,N_5059,N_5426);
and U7718 (N_7718,N_5439,N_4984);
nand U7719 (N_7719,N_4491,N_4020);
or U7720 (N_7720,N_4204,N_5565);
nor U7721 (N_7721,N_4886,N_5247);
nor U7722 (N_7722,N_4625,N_4109);
and U7723 (N_7723,N_5739,N_5275);
nor U7724 (N_7724,N_4827,N_5578);
nand U7725 (N_7725,N_5398,N_4214);
or U7726 (N_7726,N_4922,N_5103);
nand U7727 (N_7727,N_4225,N_4489);
xnor U7728 (N_7728,N_4871,N_4953);
nor U7729 (N_7729,N_4660,N_5172);
or U7730 (N_7730,N_4958,N_5368);
and U7731 (N_7731,N_5639,N_5093);
and U7732 (N_7732,N_5094,N_5332);
nand U7733 (N_7733,N_4151,N_4260);
and U7734 (N_7734,N_5004,N_5193);
nand U7735 (N_7735,N_4466,N_4146);
and U7736 (N_7736,N_4163,N_5767);
nand U7737 (N_7737,N_4669,N_4201);
xor U7738 (N_7738,N_4930,N_4104);
and U7739 (N_7739,N_5008,N_4183);
and U7740 (N_7740,N_5547,N_5992);
nand U7741 (N_7741,N_5868,N_4828);
and U7742 (N_7742,N_4585,N_5980);
and U7743 (N_7743,N_5621,N_5184);
nor U7744 (N_7744,N_4442,N_5783);
or U7745 (N_7745,N_4177,N_4363);
or U7746 (N_7746,N_4388,N_4726);
and U7747 (N_7747,N_4727,N_4609);
or U7748 (N_7748,N_5781,N_4628);
or U7749 (N_7749,N_5901,N_4894);
nand U7750 (N_7750,N_4543,N_4306);
and U7751 (N_7751,N_4671,N_4215);
nor U7752 (N_7752,N_4960,N_5349);
or U7753 (N_7753,N_4383,N_4029);
or U7754 (N_7754,N_5602,N_5679);
nand U7755 (N_7755,N_5812,N_5283);
or U7756 (N_7756,N_5422,N_5327);
and U7757 (N_7757,N_4033,N_4047);
xor U7758 (N_7758,N_4486,N_5349);
nor U7759 (N_7759,N_5701,N_4966);
and U7760 (N_7760,N_5887,N_5663);
nor U7761 (N_7761,N_4209,N_4166);
nand U7762 (N_7762,N_4151,N_4017);
and U7763 (N_7763,N_4957,N_4504);
or U7764 (N_7764,N_4178,N_4321);
nor U7765 (N_7765,N_5622,N_4637);
or U7766 (N_7766,N_4749,N_4630);
or U7767 (N_7767,N_4325,N_4683);
or U7768 (N_7768,N_5772,N_4646);
and U7769 (N_7769,N_5697,N_4726);
and U7770 (N_7770,N_5120,N_4123);
and U7771 (N_7771,N_5011,N_5521);
or U7772 (N_7772,N_5071,N_5545);
or U7773 (N_7773,N_5731,N_4426);
and U7774 (N_7774,N_5734,N_5507);
and U7775 (N_7775,N_5919,N_5992);
or U7776 (N_7776,N_4949,N_5633);
or U7777 (N_7777,N_4264,N_5628);
nand U7778 (N_7778,N_5544,N_4348);
nand U7779 (N_7779,N_5541,N_5464);
nand U7780 (N_7780,N_5400,N_5848);
nor U7781 (N_7781,N_5988,N_4866);
or U7782 (N_7782,N_4708,N_4040);
or U7783 (N_7783,N_4857,N_5692);
and U7784 (N_7784,N_4645,N_5178);
nor U7785 (N_7785,N_5864,N_5764);
nand U7786 (N_7786,N_4757,N_4853);
nand U7787 (N_7787,N_5697,N_4383);
nand U7788 (N_7788,N_5706,N_5413);
nor U7789 (N_7789,N_4369,N_4271);
or U7790 (N_7790,N_4665,N_5895);
nor U7791 (N_7791,N_4897,N_5631);
nor U7792 (N_7792,N_5228,N_4593);
xnor U7793 (N_7793,N_5245,N_4692);
or U7794 (N_7794,N_5644,N_4715);
and U7795 (N_7795,N_4717,N_4977);
nor U7796 (N_7796,N_5617,N_5718);
nand U7797 (N_7797,N_5125,N_4066);
and U7798 (N_7798,N_5788,N_4208);
nand U7799 (N_7799,N_5310,N_5994);
nor U7800 (N_7800,N_5274,N_4010);
and U7801 (N_7801,N_5129,N_5553);
nor U7802 (N_7802,N_5992,N_4456);
nor U7803 (N_7803,N_5276,N_4577);
nand U7804 (N_7804,N_5969,N_4241);
and U7805 (N_7805,N_4196,N_4363);
or U7806 (N_7806,N_4691,N_5728);
nor U7807 (N_7807,N_5765,N_5527);
nand U7808 (N_7808,N_4227,N_5847);
or U7809 (N_7809,N_5955,N_4458);
nand U7810 (N_7810,N_4138,N_4703);
nor U7811 (N_7811,N_4877,N_5462);
or U7812 (N_7812,N_5253,N_5058);
nor U7813 (N_7813,N_4247,N_4869);
nand U7814 (N_7814,N_5083,N_4024);
or U7815 (N_7815,N_4168,N_5500);
or U7816 (N_7816,N_5272,N_5361);
nor U7817 (N_7817,N_5155,N_4131);
and U7818 (N_7818,N_5881,N_5100);
and U7819 (N_7819,N_4521,N_4736);
and U7820 (N_7820,N_4096,N_5473);
or U7821 (N_7821,N_4202,N_4404);
nand U7822 (N_7822,N_4222,N_5542);
or U7823 (N_7823,N_5960,N_4456);
nor U7824 (N_7824,N_5282,N_4399);
and U7825 (N_7825,N_5656,N_4747);
and U7826 (N_7826,N_4394,N_4293);
nand U7827 (N_7827,N_4093,N_4144);
or U7828 (N_7828,N_4975,N_5701);
nor U7829 (N_7829,N_5864,N_4275);
or U7830 (N_7830,N_5262,N_5475);
and U7831 (N_7831,N_4025,N_4026);
and U7832 (N_7832,N_4907,N_4750);
nor U7833 (N_7833,N_5771,N_5032);
nor U7834 (N_7834,N_4917,N_5816);
and U7835 (N_7835,N_5915,N_5682);
or U7836 (N_7836,N_4675,N_5674);
nand U7837 (N_7837,N_5195,N_5724);
nor U7838 (N_7838,N_4152,N_5389);
or U7839 (N_7839,N_4458,N_5619);
nand U7840 (N_7840,N_5608,N_4512);
nand U7841 (N_7841,N_4301,N_4146);
nand U7842 (N_7842,N_5680,N_4984);
or U7843 (N_7843,N_4770,N_4473);
and U7844 (N_7844,N_4972,N_4595);
or U7845 (N_7845,N_5708,N_5300);
nor U7846 (N_7846,N_4348,N_5879);
or U7847 (N_7847,N_4078,N_5805);
and U7848 (N_7848,N_5786,N_5083);
nor U7849 (N_7849,N_4253,N_5384);
or U7850 (N_7850,N_5455,N_4141);
or U7851 (N_7851,N_4987,N_4479);
or U7852 (N_7852,N_5095,N_5908);
xor U7853 (N_7853,N_4753,N_4108);
nor U7854 (N_7854,N_5520,N_4080);
or U7855 (N_7855,N_5281,N_4888);
and U7856 (N_7856,N_5051,N_5793);
or U7857 (N_7857,N_4065,N_4430);
nand U7858 (N_7858,N_4989,N_4693);
nand U7859 (N_7859,N_5424,N_4063);
nand U7860 (N_7860,N_4342,N_4092);
or U7861 (N_7861,N_4720,N_5517);
xor U7862 (N_7862,N_4117,N_5777);
nand U7863 (N_7863,N_4802,N_5901);
or U7864 (N_7864,N_5985,N_5746);
and U7865 (N_7865,N_4027,N_4993);
nand U7866 (N_7866,N_5917,N_4470);
or U7867 (N_7867,N_4570,N_5386);
or U7868 (N_7868,N_4462,N_5652);
nand U7869 (N_7869,N_5825,N_4019);
nor U7870 (N_7870,N_5372,N_5490);
and U7871 (N_7871,N_4903,N_4006);
nand U7872 (N_7872,N_4308,N_4822);
nand U7873 (N_7873,N_5812,N_4192);
and U7874 (N_7874,N_5479,N_5836);
nand U7875 (N_7875,N_5954,N_4413);
or U7876 (N_7876,N_5397,N_4206);
nor U7877 (N_7877,N_5675,N_5041);
nand U7878 (N_7878,N_4324,N_4456);
and U7879 (N_7879,N_5550,N_5343);
xor U7880 (N_7880,N_4776,N_5295);
nor U7881 (N_7881,N_5376,N_4711);
nand U7882 (N_7882,N_5199,N_4035);
nand U7883 (N_7883,N_5067,N_4684);
nor U7884 (N_7884,N_5502,N_4658);
nand U7885 (N_7885,N_4387,N_4817);
nand U7886 (N_7886,N_5418,N_5498);
nand U7887 (N_7887,N_4689,N_5918);
or U7888 (N_7888,N_5221,N_5271);
and U7889 (N_7889,N_4464,N_5574);
and U7890 (N_7890,N_5324,N_4784);
or U7891 (N_7891,N_5015,N_5483);
or U7892 (N_7892,N_4772,N_5957);
and U7893 (N_7893,N_5925,N_4660);
and U7894 (N_7894,N_5629,N_4160);
nor U7895 (N_7895,N_4947,N_4498);
xor U7896 (N_7896,N_5760,N_5398);
and U7897 (N_7897,N_4260,N_4965);
or U7898 (N_7898,N_5181,N_4873);
or U7899 (N_7899,N_5823,N_4916);
nor U7900 (N_7900,N_5256,N_4536);
or U7901 (N_7901,N_4434,N_4302);
nor U7902 (N_7902,N_5950,N_5444);
nor U7903 (N_7903,N_5829,N_5248);
and U7904 (N_7904,N_4369,N_4759);
nor U7905 (N_7905,N_4487,N_5567);
or U7906 (N_7906,N_5885,N_5515);
nand U7907 (N_7907,N_4846,N_4943);
and U7908 (N_7908,N_4620,N_5656);
nand U7909 (N_7909,N_4051,N_4228);
or U7910 (N_7910,N_4933,N_5285);
nand U7911 (N_7911,N_5128,N_5274);
or U7912 (N_7912,N_5568,N_4731);
nor U7913 (N_7913,N_5527,N_5141);
or U7914 (N_7914,N_4164,N_5435);
or U7915 (N_7915,N_5668,N_4884);
or U7916 (N_7916,N_5564,N_4410);
nor U7917 (N_7917,N_5541,N_4099);
nor U7918 (N_7918,N_5799,N_4320);
nor U7919 (N_7919,N_5975,N_5547);
or U7920 (N_7920,N_4932,N_4539);
nand U7921 (N_7921,N_4168,N_4371);
or U7922 (N_7922,N_5440,N_5921);
and U7923 (N_7923,N_5795,N_4579);
or U7924 (N_7924,N_4809,N_5637);
or U7925 (N_7925,N_4136,N_4273);
nor U7926 (N_7926,N_4298,N_5856);
and U7927 (N_7927,N_4237,N_4598);
nand U7928 (N_7928,N_5562,N_4215);
or U7929 (N_7929,N_4614,N_5861);
or U7930 (N_7930,N_4692,N_5019);
or U7931 (N_7931,N_5230,N_5786);
and U7932 (N_7932,N_4898,N_4250);
or U7933 (N_7933,N_5707,N_5813);
and U7934 (N_7934,N_4191,N_4169);
and U7935 (N_7935,N_4810,N_4242);
nor U7936 (N_7936,N_4985,N_4254);
nor U7937 (N_7937,N_4577,N_4976);
or U7938 (N_7938,N_5499,N_5525);
nor U7939 (N_7939,N_4547,N_4707);
nor U7940 (N_7940,N_4546,N_4023);
and U7941 (N_7941,N_5818,N_4776);
nor U7942 (N_7942,N_5619,N_4463);
nor U7943 (N_7943,N_4242,N_4267);
or U7944 (N_7944,N_5890,N_5088);
and U7945 (N_7945,N_4087,N_5959);
nand U7946 (N_7946,N_4715,N_4880);
nand U7947 (N_7947,N_4274,N_4278);
and U7948 (N_7948,N_4083,N_4005);
nor U7949 (N_7949,N_4221,N_4883);
and U7950 (N_7950,N_4747,N_4441);
or U7951 (N_7951,N_5309,N_5742);
or U7952 (N_7952,N_5906,N_4306);
nand U7953 (N_7953,N_4262,N_4952);
or U7954 (N_7954,N_5173,N_5299);
nand U7955 (N_7955,N_5323,N_5365);
nor U7956 (N_7956,N_5032,N_4582);
nor U7957 (N_7957,N_4170,N_4788);
and U7958 (N_7958,N_4046,N_4966);
and U7959 (N_7959,N_4774,N_5728);
or U7960 (N_7960,N_5934,N_5422);
or U7961 (N_7961,N_4122,N_4546);
nand U7962 (N_7962,N_4568,N_5378);
and U7963 (N_7963,N_5601,N_4816);
or U7964 (N_7964,N_5161,N_4672);
nand U7965 (N_7965,N_4455,N_4511);
or U7966 (N_7966,N_4124,N_4282);
nor U7967 (N_7967,N_4275,N_5647);
or U7968 (N_7968,N_5763,N_4464);
nor U7969 (N_7969,N_5390,N_4765);
and U7970 (N_7970,N_4036,N_4869);
or U7971 (N_7971,N_5858,N_5019);
nand U7972 (N_7972,N_5271,N_5427);
and U7973 (N_7973,N_5544,N_4713);
nor U7974 (N_7974,N_4448,N_4071);
and U7975 (N_7975,N_4674,N_5217);
nand U7976 (N_7976,N_4313,N_5931);
nand U7977 (N_7977,N_4095,N_4546);
or U7978 (N_7978,N_5913,N_5940);
or U7979 (N_7979,N_5530,N_5111);
or U7980 (N_7980,N_5397,N_4028);
or U7981 (N_7981,N_5578,N_5783);
or U7982 (N_7982,N_5084,N_5956);
and U7983 (N_7983,N_5184,N_4710);
nor U7984 (N_7984,N_5930,N_4647);
nand U7985 (N_7985,N_4280,N_4779);
nor U7986 (N_7986,N_5447,N_5769);
nor U7987 (N_7987,N_5848,N_5414);
nor U7988 (N_7988,N_5841,N_5055);
and U7989 (N_7989,N_4135,N_4657);
and U7990 (N_7990,N_5609,N_5794);
nand U7991 (N_7991,N_4416,N_4622);
or U7992 (N_7992,N_4102,N_4012);
nor U7993 (N_7993,N_5415,N_5891);
nand U7994 (N_7994,N_5024,N_4976);
or U7995 (N_7995,N_4099,N_4375);
or U7996 (N_7996,N_5036,N_5188);
or U7997 (N_7997,N_5978,N_4322);
and U7998 (N_7998,N_4244,N_5184);
nor U7999 (N_7999,N_5247,N_4834);
nor U8000 (N_8000,N_6493,N_6274);
nand U8001 (N_8001,N_7300,N_6218);
nor U8002 (N_8002,N_6385,N_6133);
nand U8003 (N_8003,N_6322,N_7455);
and U8004 (N_8004,N_6230,N_6446);
nand U8005 (N_8005,N_7856,N_6096);
or U8006 (N_8006,N_7371,N_6032);
nor U8007 (N_8007,N_6361,N_7574);
or U8008 (N_8008,N_6691,N_6292);
and U8009 (N_8009,N_6772,N_6089);
nand U8010 (N_8010,N_7241,N_7427);
or U8011 (N_8011,N_6502,N_6549);
and U8012 (N_8012,N_6741,N_7362);
nor U8013 (N_8013,N_7720,N_7740);
and U8014 (N_8014,N_7925,N_6428);
nor U8015 (N_8015,N_6994,N_7335);
nor U8016 (N_8016,N_7726,N_6011);
or U8017 (N_8017,N_6153,N_7761);
and U8018 (N_8018,N_7178,N_6368);
nand U8019 (N_8019,N_7200,N_6574);
nor U8020 (N_8020,N_6263,N_7941);
or U8021 (N_8021,N_6855,N_7638);
nand U8022 (N_8022,N_7542,N_6588);
nand U8023 (N_8023,N_6087,N_7714);
and U8024 (N_8024,N_7217,N_6255);
or U8025 (N_8025,N_7258,N_7474);
or U8026 (N_8026,N_6989,N_6929);
and U8027 (N_8027,N_7063,N_6395);
nand U8028 (N_8028,N_6550,N_7346);
or U8029 (N_8029,N_6145,N_6935);
or U8030 (N_8030,N_7195,N_6443);
or U8031 (N_8031,N_6578,N_7845);
or U8032 (N_8032,N_7735,N_7751);
and U8033 (N_8033,N_7464,N_6885);
nand U8034 (N_8034,N_7776,N_6942);
or U8035 (N_8035,N_6670,N_6807);
nor U8036 (N_8036,N_6100,N_7489);
or U8037 (N_8037,N_7290,N_6513);
or U8038 (N_8038,N_6496,N_6727);
nand U8039 (N_8039,N_7727,N_7216);
xor U8040 (N_8040,N_7855,N_7811);
and U8041 (N_8041,N_7254,N_7480);
or U8042 (N_8042,N_6005,N_6362);
nand U8043 (N_8043,N_6162,N_6234);
or U8044 (N_8044,N_7301,N_7255);
or U8045 (N_8045,N_6532,N_7633);
nor U8046 (N_8046,N_7327,N_6376);
or U8047 (N_8047,N_7968,N_6390);
nand U8048 (N_8048,N_7957,N_7481);
nor U8049 (N_8049,N_7503,N_7533);
nand U8050 (N_8050,N_7004,N_6375);
nand U8051 (N_8051,N_7662,N_6637);
and U8052 (N_8052,N_6258,N_7450);
xor U8053 (N_8053,N_7332,N_6102);
nand U8054 (N_8054,N_6280,N_7853);
nand U8055 (N_8055,N_6504,N_7611);
nor U8056 (N_8056,N_7494,N_6478);
or U8057 (N_8057,N_6115,N_7958);
or U8058 (N_8058,N_6497,N_7094);
nor U8059 (N_8059,N_6667,N_6468);
and U8060 (N_8060,N_6004,N_7598);
nor U8061 (N_8061,N_7786,N_7848);
nor U8062 (N_8062,N_6127,N_7657);
and U8063 (N_8063,N_7066,N_7885);
nand U8064 (N_8064,N_6290,N_6778);
nor U8065 (N_8065,N_6046,N_6774);
or U8066 (N_8066,N_7838,N_7270);
or U8067 (N_8067,N_6628,N_6914);
and U8068 (N_8068,N_6076,N_6633);
or U8069 (N_8069,N_6895,N_7172);
or U8070 (N_8070,N_7682,N_6034);
and U8071 (N_8071,N_6505,N_7296);
nand U8072 (N_8072,N_7459,N_6624);
xor U8073 (N_8073,N_7160,N_6590);
and U8074 (N_8074,N_6186,N_6283);
nand U8075 (N_8075,N_7753,N_6328);
or U8076 (N_8076,N_7488,N_7147);
nand U8077 (N_8077,N_6192,N_7084);
nand U8078 (N_8078,N_7402,N_7443);
or U8079 (N_8079,N_6179,N_6349);
nand U8080 (N_8080,N_6853,N_6970);
and U8081 (N_8081,N_6854,N_7846);
or U8082 (N_8082,N_6101,N_7940);
nor U8083 (N_8083,N_6306,N_7515);
and U8084 (N_8084,N_7413,N_6320);
nor U8085 (N_8085,N_7275,N_6698);
and U8086 (N_8086,N_6587,N_7458);
or U8087 (N_8087,N_7634,N_6503);
and U8088 (N_8088,N_7830,N_7596);
or U8089 (N_8089,N_7658,N_7113);
nand U8090 (N_8090,N_7866,N_7582);
nand U8091 (N_8091,N_7131,N_7651);
and U8092 (N_8092,N_7681,N_7642);
and U8093 (N_8093,N_7243,N_6238);
or U8094 (N_8094,N_7857,N_6081);
and U8095 (N_8095,N_6334,N_6090);
or U8096 (N_8096,N_7414,N_6938);
nand U8097 (N_8097,N_6526,N_7679);
nand U8098 (N_8098,N_6545,N_6605);
nor U8099 (N_8099,N_7279,N_7356);
and U8100 (N_8100,N_7504,N_6780);
and U8101 (N_8101,N_7024,N_6596);
nand U8102 (N_8102,N_7422,N_6615);
nand U8103 (N_8103,N_6232,N_7567);
or U8104 (N_8104,N_6770,N_6050);
nand U8105 (N_8105,N_6971,N_6891);
nand U8106 (N_8106,N_7894,N_6785);
or U8107 (N_8107,N_6058,N_6437);
nand U8108 (N_8108,N_7755,N_6174);
nand U8109 (N_8109,N_6211,N_6309);
and U8110 (N_8110,N_7036,N_7931);
and U8111 (N_8111,N_7905,N_6117);
nor U8112 (N_8112,N_6052,N_6538);
and U8113 (N_8113,N_6939,N_7017);
or U8114 (N_8114,N_7706,N_7222);
or U8115 (N_8115,N_6351,N_7881);
nor U8116 (N_8116,N_7475,N_6178);
and U8117 (N_8117,N_7707,N_7153);
xnor U8118 (N_8118,N_7057,N_6374);
nand U8119 (N_8119,N_6165,N_6015);
nor U8120 (N_8120,N_6905,N_7010);
nor U8121 (N_8121,N_7096,N_6111);
nor U8122 (N_8122,N_6459,N_6874);
or U8123 (N_8123,N_6422,N_7588);
xnor U8124 (N_8124,N_7308,N_7793);
or U8125 (N_8125,N_6248,N_7770);
nor U8126 (N_8126,N_6472,N_6867);
and U8127 (N_8127,N_6715,N_6683);
nor U8128 (N_8128,N_7961,N_7944);
nand U8129 (N_8129,N_7325,N_7892);
nor U8130 (N_8130,N_7593,N_6489);
or U8131 (N_8131,N_7112,N_6959);
and U8132 (N_8132,N_6722,N_6723);
and U8133 (N_8133,N_7954,N_6851);
nor U8134 (N_8134,N_7659,N_7268);
nor U8135 (N_8135,N_6591,N_7164);
nand U8136 (N_8136,N_6233,N_6729);
nand U8137 (N_8137,N_7146,N_6427);
nand U8138 (N_8138,N_6105,N_7077);
and U8139 (N_8139,N_7765,N_7778);
and U8140 (N_8140,N_6817,N_7635);
or U8141 (N_8141,N_6932,N_6924);
and U8142 (N_8142,N_7877,N_6771);
or U8143 (N_8143,N_6528,N_7874);
or U8144 (N_8144,N_7052,N_7445);
and U8145 (N_8145,N_6169,N_6287);
or U8146 (N_8146,N_7276,N_6242);
nor U8147 (N_8147,N_7266,N_6217);
or U8148 (N_8148,N_6200,N_6921);
and U8149 (N_8149,N_7257,N_7293);
or U8150 (N_8150,N_6837,N_6572);
and U8151 (N_8151,N_6739,N_7784);
xor U8152 (N_8152,N_6980,N_7232);
or U8153 (N_8153,N_7585,N_7058);
and U8154 (N_8154,N_7444,N_6531);
nand U8155 (N_8155,N_7530,N_6933);
and U8156 (N_8156,N_7460,N_7380);
nand U8157 (N_8157,N_6412,N_7525);
nand U8158 (N_8158,N_6630,N_6696);
xnor U8159 (N_8159,N_7123,N_7591);
nor U8160 (N_8160,N_6110,N_6709);
nor U8161 (N_8161,N_7338,N_6802);
and U8162 (N_8162,N_7230,N_7182);
or U8163 (N_8163,N_6663,N_7151);
nor U8164 (N_8164,N_7190,N_7538);
nand U8165 (N_8165,N_6647,N_7867);
nor U8166 (N_8166,N_6887,N_6231);
nor U8167 (N_8167,N_6847,N_7655);
and U8168 (N_8168,N_7355,N_6239);
nor U8169 (N_8169,N_6080,N_6061);
and U8170 (N_8170,N_7436,N_6952);
nand U8171 (N_8171,N_6960,N_7605);
nor U8172 (N_8172,N_6273,N_7660);
or U8173 (N_8173,N_7779,N_7732);
and U8174 (N_8174,N_6718,N_7395);
nor U8175 (N_8175,N_6797,N_7875);
nand U8176 (N_8176,N_7724,N_7183);
or U8177 (N_8177,N_6347,N_7368);
nor U8178 (N_8178,N_6296,N_7067);
nor U8179 (N_8179,N_6552,N_7245);
or U8180 (N_8180,N_7742,N_7630);
or U8181 (N_8181,N_6660,N_6638);
and U8182 (N_8182,N_6713,N_6808);
nor U8183 (N_8183,N_6191,N_7055);
or U8184 (N_8184,N_7448,N_7080);
nand U8185 (N_8185,N_6652,N_7713);
and U8186 (N_8186,N_6302,N_6492);
nor U8187 (N_8187,N_7558,N_6579);
or U8188 (N_8188,N_6400,N_6640);
nor U8189 (N_8189,N_6702,N_7981);
and U8190 (N_8190,N_6359,N_6403);
xor U8191 (N_8191,N_6609,N_6398);
nor U8192 (N_8192,N_7637,N_6405);
nand U8193 (N_8193,N_6346,N_7526);
or U8194 (N_8194,N_7683,N_6927);
or U8195 (N_8195,N_6235,N_6171);
nand U8196 (N_8196,N_6956,N_7076);
nor U8197 (N_8197,N_6453,N_6031);
nor U8198 (N_8198,N_6986,N_6278);
or U8199 (N_8199,N_7697,N_7691);
or U8200 (N_8200,N_7795,N_6372);
nor U8201 (N_8201,N_6471,N_6196);
nand U8202 (N_8202,N_7367,N_6991);
and U8203 (N_8203,N_7271,N_6800);
and U8204 (N_8204,N_7365,N_6114);
and U8205 (N_8205,N_6122,N_6546);
or U8206 (N_8206,N_7331,N_6355);
or U8207 (N_8207,N_7433,N_7420);
or U8208 (N_8208,N_7393,N_7832);
or U8209 (N_8209,N_6634,N_7214);
or U8210 (N_8210,N_6260,N_6285);
nor U8211 (N_8211,N_6069,N_6955);
and U8212 (N_8212,N_6295,N_7208);
nand U8213 (N_8213,N_6898,N_7044);
and U8214 (N_8214,N_6023,N_6918);
and U8215 (N_8215,N_7127,N_6075);
nand U8216 (N_8216,N_6210,N_7302);
nand U8217 (N_8217,N_7099,N_6612);
nand U8218 (N_8218,N_7839,N_7749);
nor U8219 (N_8219,N_7221,N_6088);
and U8220 (N_8220,N_7689,N_7942);
and U8221 (N_8221,N_7895,N_6181);
and U8222 (N_8222,N_7834,N_6144);
or U8223 (N_8223,N_7640,N_7813);
and U8224 (N_8224,N_7267,N_7675);
and U8225 (N_8225,N_7921,N_6301);
nand U8226 (N_8226,N_6139,N_7240);
nor U8227 (N_8227,N_6595,N_6893);
nand U8228 (N_8228,N_6404,N_6903);
nand U8229 (N_8229,N_6170,N_6305);
or U8230 (N_8230,N_6430,N_6650);
and U8231 (N_8231,N_6265,N_7913);
nand U8232 (N_8232,N_7403,N_7476);
nand U8233 (N_8233,N_7979,N_6944);
or U8234 (N_8234,N_7361,N_6877);
and U8235 (N_8235,N_6768,N_7406);
or U8236 (N_8236,N_7535,N_7752);
nand U8237 (N_8237,N_7298,N_6469);
or U8238 (N_8238,N_7023,N_6821);
nor U8239 (N_8239,N_7141,N_7704);
nor U8240 (N_8240,N_7390,N_7934);
or U8241 (N_8241,N_6414,N_6070);
nand U8242 (N_8242,N_7359,N_6910);
or U8243 (N_8243,N_6465,N_6336);
and U8244 (N_8244,N_6190,N_7159);
xnor U8245 (N_8245,N_7677,N_6098);
and U8246 (N_8246,N_6920,N_6432);
nor U8247 (N_8247,N_7625,N_6544);
nand U8248 (N_8248,N_6262,N_6187);
nand U8249 (N_8249,N_7976,N_6694);
and U8250 (N_8250,N_7008,N_6752);
or U8251 (N_8251,N_6244,N_7757);
nor U8252 (N_8252,N_7815,N_6714);
nand U8253 (N_8253,N_6480,N_7246);
or U8254 (N_8254,N_7982,N_7452);
nand U8255 (N_8255,N_6142,N_6749);
xnor U8256 (N_8256,N_6279,N_7614);
nor U8257 (N_8257,N_6473,N_6731);
or U8258 (N_8258,N_7386,N_6182);
nor U8259 (N_8259,N_7577,N_7064);
nand U8260 (N_8260,N_7528,N_6216);
nor U8261 (N_8261,N_6677,N_7927);
nor U8262 (N_8262,N_6726,N_7360);
or U8263 (N_8263,N_6530,N_6123);
xor U8264 (N_8264,N_6733,N_6108);
nor U8265 (N_8265,N_7788,N_7138);
or U8266 (N_8266,N_6711,N_7817);
or U8267 (N_8267,N_7973,N_7062);
nor U8268 (N_8268,N_6379,N_6879);
or U8269 (N_8269,N_7003,N_6413);
nand U8270 (N_8270,N_7608,N_6215);
nor U8271 (N_8271,N_6458,N_7952);
nand U8272 (N_8272,N_7495,N_6205);
nor U8273 (N_8273,N_7553,N_7345);
nor U8274 (N_8274,N_7666,N_6394);
and U8275 (N_8275,N_7703,N_6167);
nand U8276 (N_8276,N_6317,N_7589);
and U8277 (N_8277,N_7334,N_7569);
nor U8278 (N_8278,N_7859,N_6845);
nor U8279 (N_8279,N_6534,N_7862);
nand U8280 (N_8280,N_6150,N_7167);
nor U8281 (N_8281,N_6417,N_6904);
or U8282 (N_8282,N_7518,N_7060);
or U8283 (N_8283,N_7728,N_7226);
nand U8284 (N_8284,N_6212,N_6401);
and U8285 (N_8285,N_6483,N_6685);
nor U8286 (N_8286,N_6318,N_6018);
nand U8287 (N_8287,N_7858,N_6063);
and U8288 (N_8288,N_7841,N_7229);
or U8289 (N_8289,N_7373,N_6455);
nor U8290 (N_8290,N_6119,N_7224);
or U8291 (N_8291,N_7854,N_6022);
nand U8292 (N_8292,N_7928,N_6676);
nand U8293 (N_8293,N_6491,N_7133);
nand U8294 (N_8294,N_7235,N_7708);
nand U8295 (N_8295,N_6999,N_6341);
nand U8296 (N_8296,N_7483,N_7110);
nand U8297 (N_8297,N_6352,N_6849);
or U8298 (N_8298,N_7871,N_7026);
nand U8299 (N_8299,N_6149,N_6024);
nand U8300 (N_8300,N_6957,N_6277);
and U8301 (N_8301,N_7321,N_7328);
and U8302 (N_8302,N_6449,N_6565);
and U8303 (N_8303,N_7185,N_7378);
nand U8304 (N_8304,N_6071,N_7397);
and U8305 (N_8305,N_6020,N_6717);
nand U8306 (N_8306,N_7725,N_6928);
and U8307 (N_8307,N_6477,N_6901);
xor U8308 (N_8308,N_6902,N_7644);
nand U8309 (N_8309,N_7478,N_7011);
nor U8310 (N_8310,N_6500,N_7676);
nand U8311 (N_8311,N_7180,N_6906);
or U8312 (N_8312,N_6668,N_7006);
and U8313 (N_8313,N_7796,N_7033);
nor U8314 (N_8314,N_6976,N_7576);
and U8315 (N_8315,N_7654,N_7620);
nand U8316 (N_8316,N_6930,N_6725);
nor U8317 (N_8317,N_7915,N_6747);
and U8318 (N_8318,N_7808,N_7668);
and U8319 (N_8319,N_6391,N_6256);
nand U8320 (N_8320,N_6784,N_7031);
and U8321 (N_8321,N_6570,N_7069);
nand U8322 (N_8322,N_7259,N_7363);
and U8323 (N_8323,N_7912,N_7392);
nand U8324 (N_8324,N_6060,N_6326);
and U8325 (N_8325,N_7583,N_7398);
or U8326 (N_8326,N_6342,N_7597);
nand U8327 (N_8327,N_7696,N_7029);
nor U8328 (N_8328,N_6183,N_7065);
or U8329 (N_8329,N_7194,N_6822);
and U8330 (N_8330,N_7449,N_7790);
and U8331 (N_8331,N_6766,N_7804);
and U8332 (N_8332,N_7656,N_7040);
or U8333 (N_8333,N_7169,N_7517);
nand U8334 (N_8334,N_6353,N_7670);
and U8335 (N_8335,N_7016,N_7090);
nand U8336 (N_8336,N_7442,N_6213);
and U8337 (N_8337,N_7264,N_6969);
nor U8338 (N_8338,N_7309,N_7107);
nand U8339 (N_8339,N_6019,N_6626);
and U8340 (N_8340,N_6160,N_6763);
nor U8341 (N_8341,N_7119,N_7693);
and U8342 (N_8342,N_7391,N_6864);
and U8343 (N_8343,N_6601,N_6863);
or U8344 (N_8344,N_7739,N_7946);
or U8345 (N_8345,N_7079,N_6053);
and U8346 (N_8346,N_6720,N_7074);
nand U8347 (N_8347,N_6486,N_6961);
or U8348 (N_8348,N_6298,N_6567);
nor U8349 (N_8349,N_7695,N_7157);
or U8350 (N_8350,N_7537,N_7295);
or U8351 (N_8351,N_6745,N_6629);
and U8352 (N_8352,N_7179,N_6831);
and U8353 (N_8353,N_7181,N_6762);
or U8354 (N_8354,N_7204,N_7672);
and U8355 (N_8355,N_6383,N_7326);
nor U8356 (N_8356,N_7082,N_6356);
nor U8357 (N_8357,N_7315,N_6131);
nor U8358 (N_8358,N_7203,N_7700);
nand U8359 (N_8359,N_6225,N_7985);
nor U8360 (N_8360,N_7409,N_7125);
nor U8361 (N_8361,N_7501,N_6045);
nor U8362 (N_8362,N_6981,N_7350);
or U8363 (N_8363,N_6293,N_7998);
or U8364 (N_8364,N_7103,N_7565);
and U8365 (N_8365,N_6646,N_6421);
or U8366 (N_8366,N_7917,N_6716);
nor U8367 (N_8367,N_6365,N_6852);
and U8368 (N_8368,N_7626,N_7771);
or U8369 (N_8369,N_6476,N_7711);
nand U8370 (N_8370,N_7206,N_7836);
nor U8371 (N_8371,N_7247,N_7333);
or U8372 (N_8372,N_7760,N_6997);
nor U8373 (N_8373,N_7799,N_6386);
nand U8374 (N_8374,N_7073,N_7539);
and U8375 (N_8375,N_7712,N_7888);
nor U8376 (N_8376,N_7508,N_6724);
and U8377 (N_8377,N_6641,N_6943);
or U8378 (N_8378,N_7143,N_7890);
nor U8379 (N_8379,N_7234,N_6913);
and U8380 (N_8380,N_7903,N_7384);
nand U8381 (N_8381,N_7860,N_7089);
nor U8382 (N_8382,N_6543,N_6016);
and U8383 (N_8383,N_7613,N_6012);
nor U8384 (N_8384,N_6884,N_7375);
and U8385 (N_8385,N_7186,N_7631);
or U8386 (N_8386,N_7212,N_6790);
nor U8387 (N_8387,N_6585,N_6072);
or U8388 (N_8388,N_7897,N_6840);
nand U8389 (N_8389,N_7906,N_7320);
and U8390 (N_8390,N_6878,N_7828);
or U8391 (N_8391,N_6589,N_7000);
nor U8392 (N_8392,N_7935,N_6614);
nor U8393 (N_8393,N_7566,N_6744);
nor U8394 (N_8394,N_7075,N_6697);
nor U8395 (N_8395,N_7868,N_7262);
nand U8396 (N_8396,N_7665,N_6039);
or U8397 (N_8397,N_6158,N_7319);
nor U8398 (N_8398,N_6484,N_6059);
nor U8399 (N_8399,N_6339,N_6533);
nand U8400 (N_8400,N_7163,N_7046);
nand U8401 (N_8401,N_6692,N_7081);
or U8402 (N_8402,N_6041,N_6632);
and U8403 (N_8403,N_6452,N_6673);
and U8404 (N_8404,N_7498,N_6340);
and U8405 (N_8405,N_7898,N_6580);
nor U8406 (N_8406,N_6161,N_7819);
nand U8407 (N_8407,N_7312,N_6104);
nand U8408 (N_8408,N_7009,N_7516);
nand U8409 (N_8409,N_6796,N_7963);
and U8410 (N_8410,N_6291,N_6987);
nand U8411 (N_8411,N_7030,N_6838);
or U8412 (N_8412,N_7643,N_7166);
or U8413 (N_8413,N_6425,N_7507);
or U8414 (N_8414,N_6824,N_7490);
and U8415 (N_8415,N_7314,N_6621);
nor U8416 (N_8416,N_6049,N_7568);
or U8417 (N_8417,N_6220,N_7156);
and U8418 (N_8418,N_7197,N_7387);
nand U8419 (N_8419,N_6582,N_6982);
or U8420 (N_8420,N_6661,N_6345);
or U8421 (N_8421,N_6511,N_6776);
nor U8422 (N_8422,N_6799,N_7358);
nand U8423 (N_8423,N_7184,N_7242);
nor U8424 (N_8424,N_6889,N_7344);
and U8425 (N_8425,N_7015,N_7134);
and U8426 (N_8426,N_7685,N_6962);
or U8427 (N_8427,N_7109,N_6508);
nor U8428 (N_8428,N_7733,N_6861);
nand U8429 (N_8429,N_7272,N_7557);
nor U8430 (N_8430,N_6839,N_7383);
and U8431 (N_8431,N_6332,N_7410);
or U8432 (N_8432,N_6788,N_6463);
or U8433 (N_8433,N_6586,N_7926);
nand U8434 (N_8434,N_7136,N_6806);
or U8435 (N_8435,N_7872,N_6042);
or U8436 (N_8436,N_6276,N_6958);
nor U8437 (N_8437,N_6311,N_7698);
and U8438 (N_8438,N_7806,N_6708);
nand U8439 (N_8439,N_6393,N_7850);
and U8440 (N_8440,N_6789,N_7105);
nand U8441 (N_8441,N_6056,N_6501);
or U8442 (N_8442,N_6740,N_6557);
nand U8443 (N_8443,N_7852,N_6227);
nor U8444 (N_8444,N_6040,N_7924);
nor U8445 (N_8445,N_6793,N_7715);
nand U8446 (N_8446,N_7821,N_7457);
nand U8447 (N_8447,N_6219,N_6786);
or U8448 (N_8448,N_6541,N_7541);
nand U8449 (N_8449,N_7191,N_6872);
and U8450 (N_8450,N_6564,N_7174);
nand U8451 (N_8451,N_6810,N_6602);
and U8452 (N_8452,N_7369,N_6257);
nor U8453 (N_8453,N_7260,N_7606);
and U8454 (N_8454,N_7282,N_6253);
nand U8455 (N_8455,N_7994,N_7018);
and U8456 (N_8456,N_6517,N_6389);
and U8457 (N_8457,N_6300,N_7536);
nand U8458 (N_8458,N_6998,N_6573);
nand U8459 (N_8459,N_6571,N_6876);
or U8460 (N_8460,N_6767,N_7607);
nor U8461 (N_8461,N_6499,N_7288);
nor U8462 (N_8462,N_7299,N_7984);
nor U8463 (N_8463,N_7964,N_6655);
nand U8464 (N_8464,N_7822,N_6972);
and U8465 (N_8465,N_6429,N_7650);
and U8466 (N_8466,N_7645,N_6335);
and U8467 (N_8467,N_6424,N_6523);
or U8468 (N_8468,N_7218,N_7198);
nor U8469 (N_8469,N_7324,N_7559);
nor U8470 (N_8470,N_7610,N_7261);
or U8471 (N_8471,N_7896,N_7794);
xor U8472 (N_8472,N_6803,N_6035);
or U8473 (N_8473,N_6835,N_6267);
nand U8474 (N_8474,N_7418,N_7002);
nor U8475 (N_8475,N_7472,N_7734);
nor U8476 (N_8476,N_6409,N_7990);
nor U8477 (N_8477,N_7624,N_7124);
and U8478 (N_8478,N_7086,N_6689);
xnor U8479 (N_8479,N_6323,N_6859);
nor U8480 (N_8480,N_6204,N_6710);
nand U8481 (N_8481,N_7937,N_7401);
nor U8482 (N_8482,N_7661,N_6606);
and U8483 (N_8483,N_6965,N_6966);
nand U8484 (N_8484,N_6487,N_7746);
nand U8485 (N_8485,N_6520,N_6608);
nand U8486 (N_8486,N_7987,N_7933);
and U8487 (N_8487,N_7021,N_6915);
or U8488 (N_8488,N_6164,N_7783);
or U8489 (N_8489,N_6703,N_6013);
nor U8490 (N_8490,N_6156,N_7285);
nand U8491 (N_8491,N_6091,N_6354);
or U8492 (N_8492,N_7148,N_7548);
nor U8493 (N_8493,N_7253,N_6241);
nor U8494 (N_8494,N_6568,N_7762);
nand U8495 (N_8495,N_6199,N_6438);
nor U8496 (N_8496,N_6313,N_7014);
and U8497 (N_8497,N_6542,N_6448);
and U8498 (N_8498,N_6540,N_7722);
nand U8499 (N_8499,N_6791,N_6209);
or U8500 (N_8500,N_6054,N_7883);
nor U8501 (N_8501,N_7612,N_6275);
or U8502 (N_8502,N_7114,N_7428);
nand U8503 (N_8503,N_6555,N_7438);
nand U8504 (N_8504,N_6314,N_6636);
or U8505 (N_8505,N_6514,N_6085);
or U8506 (N_8506,N_6125,N_7189);
or U8507 (N_8507,N_7265,N_7231);
nor U8508 (N_8508,N_6581,N_7965);
and U8509 (N_8509,N_6719,N_6193);
nand U8510 (N_8510,N_6524,N_6147);
and U8511 (N_8511,N_7774,N_7962);
and U8512 (N_8512,N_6721,N_6264);
nand U8513 (N_8513,N_6176,N_6594);
nor U8514 (N_8514,N_7664,N_6858);
and U8515 (N_8515,N_6925,N_6936);
and U8516 (N_8516,N_6307,N_6880);
nor U8517 (N_8517,N_7307,N_6820);
nor U8518 (N_8518,N_7087,N_7150);
nor U8519 (N_8519,N_6135,N_6946);
nand U8520 (N_8520,N_6569,N_7223);
nor U8521 (N_8521,N_7723,N_7818);
nand U8522 (N_8522,N_6418,N_7863);
nor U8523 (N_8523,N_6559,N_6221);
and U8524 (N_8524,N_6095,N_6554);
nand U8525 (N_8525,N_6420,N_6862);
and U8526 (N_8526,N_6475,N_6129);
and U8527 (N_8527,N_7341,N_7463);
or U8528 (N_8528,N_6750,N_6436);
nor U8529 (N_8529,N_6795,N_7955);
or U8530 (N_8530,N_7812,N_6494);
nand U8531 (N_8531,N_7977,N_7085);
or U8532 (N_8532,N_6856,N_6627);
nor U8533 (N_8533,N_7602,N_7256);
nand U8534 (N_8534,N_6860,N_6047);
nor U8535 (N_8535,N_7599,N_7527);
nor U8536 (N_8536,N_6882,N_6194);
nor U8537 (N_8537,N_7330,N_7461);
nand U8538 (N_8538,N_6699,N_6945);
or U8539 (N_8539,N_7947,N_7152);
nor U8540 (N_8540,N_6639,N_7844);
and U8541 (N_8541,N_6266,N_6402);
and U8542 (N_8542,N_6208,N_6188);
or U8543 (N_8543,N_6021,N_7477);
nor U8544 (N_8544,N_6426,N_7056);
nand U8545 (N_8545,N_7120,N_6746);
nor U8546 (N_8546,N_7616,N_6246);
and U8547 (N_8547,N_6575,N_6804);
nor U8548 (N_8548,N_6649,N_6963);
or U8549 (N_8549,N_7649,N_7487);
or U8550 (N_8550,N_6657,N_6134);
and U8551 (N_8551,N_7505,N_7663);
or U8552 (N_8552,N_7465,N_7907);
and U8553 (N_8553,N_7587,N_7512);
nor U8554 (N_8554,N_6635,N_6488);
nand U8555 (N_8555,N_6152,N_7560);
nand U8556 (N_8556,N_7193,N_7317);
and U8557 (N_8557,N_7211,N_7580);
or U8558 (N_8558,N_7205,N_7078);
nor U8559 (N_8559,N_7807,N_7540);
nand U8560 (N_8560,N_6734,N_6259);
xor U8561 (N_8561,N_6038,N_6392);
and U8562 (N_8562,N_6457,N_7594);
nand U8563 (N_8563,N_7429,N_7423);
or U8564 (N_8564,N_6990,N_6704);
and U8565 (N_8565,N_7621,N_6521);
nand U8566 (N_8566,N_6367,N_6758);
and U8567 (N_8567,N_7286,N_6084);
or U8568 (N_8568,N_6850,N_7646);
nor U8569 (N_8569,N_7581,N_6408);
or U8570 (N_8570,N_6159,N_7311);
nand U8571 (N_8571,N_7609,N_6360);
and U8572 (N_8572,N_6551,N_6754);
or U8573 (N_8573,N_7432,N_7430);
and U8574 (N_8574,N_7730,N_6593);
and U8575 (N_8575,N_6556,N_6558);
and U8576 (N_8576,N_6113,N_7400);
nor U8577 (N_8577,N_6842,N_7564);
or U8578 (N_8578,N_7043,N_6143);
or U8579 (N_8579,N_6826,N_7377);
or U8580 (N_8580,N_6396,N_6203);
nand U8581 (N_8581,N_6120,N_6330);
and U8582 (N_8582,N_6783,N_7709);
nand U8583 (N_8583,N_6979,N_6166);
and U8584 (N_8584,N_7759,N_7995);
and U8585 (N_8585,N_6712,N_6512);
and U8586 (N_8586,N_6207,N_7546);
and U8587 (N_8587,N_6434,N_7101);
nand U8588 (N_8588,N_6055,N_7949);
and U8589 (N_8589,N_6684,N_6949);
and U8590 (N_8590,N_7108,N_6737);
and U8591 (N_8591,N_7738,N_6440);
nor U8592 (N_8592,N_7446,N_7978);
or U8593 (N_8593,N_6563,N_6656);
nor U8594 (N_8594,N_7284,N_7870);
nand U8595 (N_8595,N_6760,N_7632);
or U8596 (N_8596,N_6319,N_7176);
nor U8597 (N_8597,N_6481,N_6387);
and U8598 (N_8598,N_6679,N_6083);
and U8599 (N_8599,N_7415,N_7139);
nor U8600 (N_8600,N_6671,N_6482);
or U8601 (N_8601,N_7054,N_7847);
nor U8602 (N_8602,N_7684,N_7128);
and U8603 (N_8603,N_7622,N_7831);
nor U8604 (N_8604,N_7554,N_6813);
and U8605 (N_8605,N_6525,N_7399);
and U8606 (N_8606,N_6106,N_7027);
nand U8607 (N_8607,N_7469,N_6299);
and U8608 (N_8608,N_7227,N_6964);
nor U8609 (N_8609,N_6562,N_6001);
nand U8610 (N_8610,N_6645,N_6948);
nand U8611 (N_8611,N_7766,N_6583);
or U8612 (N_8612,N_7374,N_6027);
xnor U8613 (N_8613,N_7922,N_7337);
nor U8614 (N_8614,N_6818,N_6917);
nand U8615 (N_8615,N_7833,N_6777);
and U8616 (N_8616,N_7969,N_7088);
and U8617 (N_8617,N_6338,N_7532);
nor U8618 (N_8618,N_7513,N_6331);
and U8619 (N_8619,N_7353,N_6841);
and U8620 (N_8620,N_7207,N_7149);
and U8621 (N_8621,N_6653,N_7142);
or U8622 (N_8622,N_7878,N_7322);
nand U8623 (N_8623,N_7485,N_7690);
nor U8624 (N_8624,N_7950,N_6406);
nor U8625 (N_8625,N_7028,N_7175);
nor U8626 (N_8626,N_7165,N_7425);
nor U8627 (N_8627,N_6003,N_6553);
nor U8628 (N_8628,N_6705,N_7801);
nand U8629 (N_8629,N_7604,N_7652);
or U8630 (N_8630,N_6576,N_7986);
and U8631 (N_8631,N_7687,N_7641);
nor U8632 (N_8632,N_7747,N_6598);
xor U8633 (N_8633,N_6140,N_6873);
and U8634 (N_8634,N_7861,N_6329);
and U8635 (N_8635,N_7556,N_7617);
nand U8636 (N_8636,N_6658,N_6812);
nand U8637 (N_8637,N_6082,N_7287);
and U8638 (N_8638,N_6675,N_6097);
nor U8639 (N_8639,N_7750,N_6600);
and U8640 (N_8640,N_6155,N_7627);
or U8641 (N_8641,N_7201,N_7745);
nor U8642 (N_8642,N_6967,N_7692);
nand U8643 (N_8643,N_7435,N_7013);
and U8644 (N_8644,N_7603,N_6431);
or U8645 (N_8645,N_6214,N_7283);
and U8646 (N_8646,N_6222,N_7772);
nor U8647 (N_8647,N_7154,N_7405);
and U8648 (N_8648,N_7876,N_7869);
nand U8649 (N_8649,N_6008,N_6922);
and U8650 (N_8650,N_7579,N_7382);
nor U8651 (N_8651,N_7615,N_6358);
or U8652 (N_8652,N_6377,N_6756);
nor U8653 (N_8653,N_7803,N_6919);
and U8654 (N_8654,N_7484,N_7177);
nand U8655 (N_8655,N_6566,N_7336);
nand U8656 (N_8656,N_7918,N_7236);
nor U8657 (N_8657,N_6173,N_7923);
nor U8658 (N_8658,N_6268,N_6669);
xor U8659 (N_8659,N_7005,N_7520);
or U8660 (N_8660,N_6537,N_6324);
or U8661 (N_8661,N_6730,N_7274);
or U8662 (N_8662,N_7550,N_7741);
or U8663 (N_8663,N_7424,N_7252);
and U8664 (N_8664,N_7511,N_7767);
or U8665 (N_8665,N_6033,N_6761);
or U8666 (N_8666,N_7104,N_7547);
or U8667 (N_8667,N_6249,N_7434);
nand U8668 (N_8668,N_7161,N_7938);
nor U8669 (N_8669,N_7744,N_7843);
nand U8670 (N_8670,N_6951,N_7389);
nor U8671 (N_8671,N_6495,N_6700);
xnor U8672 (N_8672,N_7805,N_7768);
or U8673 (N_8673,N_6177,N_7468);
and U8674 (N_8674,N_7210,N_6801);
nand U8675 (N_8675,N_6674,N_6094);
nor U8676 (N_8676,N_6371,N_6798);
or U8677 (N_8677,N_7372,N_7170);
and U8678 (N_8678,N_6009,N_7278);
nand U8679 (N_8679,N_7041,N_7993);
nand U8680 (N_8680,N_7305,N_6975);
nand U8681 (N_8681,N_6197,N_6198);
or U8682 (N_8682,N_7780,N_6282);
and U8683 (N_8683,N_6732,N_6315);
or U8684 (N_8684,N_6782,N_6077);
or U8685 (N_8685,N_7441,N_7310);
nand U8686 (N_8686,N_6787,N_7269);
and U8687 (N_8687,N_6896,N_6926);
and U8688 (N_8688,N_6043,N_7019);
nand U8689 (N_8689,N_6954,N_6823);
xnor U8690 (N_8690,N_7972,N_6738);
xor U8691 (N_8691,N_7352,N_7048);
and U8692 (N_8692,N_6461,N_7549);
nand U8693 (N_8693,N_7510,N_6435);
xor U8694 (N_8694,N_6619,N_6126);
and U8695 (N_8695,N_7462,N_7717);
nand U8696 (N_8696,N_6868,N_7792);
xnor U8697 (N_8697,N_7718,N_7440);
nand U8698 (N_8698,N_6378,N_7721);
nand U8699 (N_8699,N_6451,N_6736);
nor U8700 (N_8700,N_7479,N_7244);
or U8701 (N_8701,N_7902,N_7966);
or U8702 (N_8702,N_6103,N_6237);
xor U8703 (N_8703,N_7304,N_6857);
or U8704 (N_8704,N_6539,N_7787);
or U8705 (N_8705,N_7118,N_6974);
and U8706 (N_8706,N_6229,N_6261);
and U8707 (N_8707,N_6366,N_6223);
and U8708 (N_8708,N_7238,N_6000);
nand U8709 (N_8709,N_6832,N_6289);
and U8710 (N_8710,N_6779,N_7904);
and U8711 (N_8711,N_7342,N_6441);
or U8712 (N_8712,N_6875,N_6067);
or U8713 (N_8713,N_7158,N_7835);
and U8714 (N_8714,N_7702,N_6506);
and U8715 (N_8715,N_6892,N_6611);
or U8716 (N_8716,N_6931,N_7509);
nand U8717 (N_8717,N_7887,N_6834);
nor U8718 (N_8718,N_6825,N_7671);
and U8719 (N_8719,N_7220,N_6308);
or U8720 (N_8720,N_6916,N_7820);
and U8721 (N_8721,N_7093,N_6687);
nor U8722 (N_8722,N_6093,N_7743);
or U8723 (N_8723,N_6757,N_6245);
and U8724 (N_8724,N_6680,N_7578);
and U8725 (N_8725,N_7225,N_7144);
nor U8726 (N_8726,N_6755,N_6454);
nand U8727 (N_8727,N_7249,N_7523);
nor U8728 (N_8728,N_7097,N_6664);
nor U8729 (N_8729,N_7126,N_7705);
nor U8730 (N_8730,N_7168,N_7500);
nor U8731 (N_8731,N_6527,N_7826);
nand U8732 (N_8732,N_6651,N_7900);
nand U8733 (N_8733,N_6662,N_6252);
and U8734 (N_8734,N_6597,N_7758);
and U8735 (N_8735,N_6466,N_6599);
nand U8736 (N_8736,N_7072,N_7098);
nand U8737 (N_8737,N_6014,N_6029);
and U8738 (N_8738,N_6765,N_6247);
nand U8739 (N_8739,N_6444,N_7970);
nor U8740 (N_8740,N_7421,N_7899);
nor U8741 (N_8741,N_6201,N_6068);
nand U8742 (N_8742,N_7800,N_7719);
and U8743 (N_8743,N_7281,N_7534);
nor U8744 (N_8744,N_7466,N_7070);
nand U8745 (N_8745,N_6843,N_6333);
nand U8746 (N_8746,N_6397,N_6509);
or U8747 (N_8747,N_6348,N_6381);
and U8748 (N_8748,N_7851,N_7388);
or U8749 (N_8749,N_6607,N_6682);
nand U8750 (N_8750,N_7882,N_6086);
and U8751 (N_8751,N_6659,N_7411);
nor U8752 (N_8752,N_7601,N_7376);
xnor U8753 (N_8753,N_7797,N_6666);
nor U8754 (N_8754,N_6529,N_6686);
nor U8755 (N_8755,N_7092,N_7187);
nand U8756 (N_8756,N_7381,N_6672);
nor U8757 (N_8757,N_7102,N_6118);
nor U8758 (N_8758,N_7280,N_6984);
nand U8759 (N_8759,N_6547,N_7053);
nand U8760 (N_8760,N_7291,N_6030);
and U8761 (N_8761,N_7042,N_7636);
nor U8762 (N_8762,N_6467,N_7891);
or U8763 (N_8763,N_7145,N_6099);
nor U8764 (N_8764,N_6648,N_6226);
and U8765 (N_8765,N_6130,N_7571);
or U8766 (N_8766,N_7499,N_7531);
nor U8767 (N_8767,N_7482,N_7453);
or U8768 (N_8768,N_6168,N_6848);
or U8769 (N_8769,N_7116,N_7034);
xnor U8770 (N_8770,N_7357,N_6109);
or U8771 (N_8771,N_6995,N_7667);
or U8772 (N_8772,N_6415,N_7496);
nor U8773 (N_8773,N_7038,N_7678);
and U8774 (N_8774,N_6992,N_6151);
nor U8775 (N_8775,N_6978,N_6894);
nand U8776 (N_8776,N_7901,N_6092);
nand U8777 (N_8777,N_6792,N_6827);
nor U8778 (N_8778,N_6107,N_7842);
nor U8779 (N_8779,N_6002,N_6370);
nor U8780 (N_8780,N_6138,N_6037);
or U8781 (N_8781,N_7417,N_7932);
or U8782 (N_8782,N_7454,N_7997);
or U8783 (N_8783,N_7318,N_7773);
nand U8784 (N_8784,N_6419,N_7920);
and U8785 (N_8785,N_7343,N_7996);
or U8786 (N_8786,N_6357,N_7840);
and U8787 (N_8787,N_6871,N_7584);
xor U8788 (N_8788,N_6272,N_7959);
nand U8789 (N_8789,N_6310,N_7292);
nor U8790 (N_8790,N_7929,N_6644);
nor U8791 (N_8791,N_7673,N_6604);
nand U8792 (N_8792,N_7729,N_6206);
and U8793 (N_8793,N_6157,N_7313);
or U8794 (N_8794,N_7590,N_6116);
nor U8795 (N_8795,N_7756,N_6678);
nor U8796 (N_8796,N_6316,N_7192);
nor U8797 (N_8797,N_7629,N_6620);
nor U8798 (N_8798,N_7623,N_6490);
and U8799 (N_8799,N_7595,N_7639);
nand U8800 (N_8800,N_6180,N_6006);
nand U8801 (N_8801,N_6516,N_6507);
nor U8802 (N_8802,N_6814,N_6136);
nand U8803 (N_8803,N_7199,N_6026);
nand U8804 (N_8804,N_7802,N_6616);
and U8805 (N_8805,N_7791,N_7020);
and U8806 (N_8806,N_7140,N_6294);
and U8807 (N_8807,N_6498,N_7716);
and U8808 (N_8808,N_7297,N_6781);
nor U8809 (N_8809,N_6707,N_6977);
and U8810 (N_8810,N_7880,N_7910);
nand U8811 (N_8811,N_6128,N_7879);
nor U8812 (N_8812,N_6343,N_7991);
and U8813 (N_8813,N_7137,N_6240);
or U8814 (N_8814,N_6074,N_7370);
nand U8815 (N_8815,N_7306,N_7135);
and U8816 (N_8816,N_7980,N_7763);
and U8817 (N_8817,N_7956,N_7456);
and U8818 (N_8818,N_7519,N_7111);
or U8819 (N_8819,N_6172,N_7347);
nand U8820 (N_8820,N_7555,N_6665);
or U8821 (N_8821,N_6830,N_7239);
and U8822 (N_8822,N_7404,N_6141);
and U8823 (N_8823,N_7543,N_6610);
and U8824 (N_8824,N_6941,N_6010);
nor U8825 (N_8825,N_6753,N_6470);
nor U8826 (N_8826,N_6121,N_6828);
nand U8827 (N_8827,N_7524,N_7506);
nor U8828 (N_8828,N_7971,N_7619);
nor U8829 (N_8829,N_6866,N_6881);
or U8830 (N_8830,N_7379,N_6078);
nand U8831 (N_8831,N_7045,N_6809);
or U8832 (N_8832,N_7967,N_7939);
nand U8833 (N_8833,N_6456,N_7059);
and U8834 (N_8834,N_7575,N_6057);
and U8835 (N_8835,N_6695,N_6816);
and U8836 (N_8836,N_7573,N_6869);
nand U8837 (N_8837,N_6846,N_6983);
nor U8838 (N_8838,N_6759,N_6643);
and U8839 (N_8839,N_6735,N_7893);
and U8840 (N_8840,N_7930,N_6380);
and U8841 (N_8841,N_7426,N_7025);
or U8842 (N_8842,N_7447,N_7809);
nor U8843 (N_8843,N_7731,N_6728);
nand U8844 (N_8844,N_6897,N_7001);
and U8845 (N_8845,N_6439,N_6617);
or U8846 (N_8846,N_7688,N_7233);
and U8847 (N_8847,N_6815,N_6474);
and U8848 (N_8848,N_7789,N_6561);
nand U8849 (N_8849,N_7354,N_7316);
and U8850 (N_8850,N_6048,N_7394);
nand U8851 (N_8851,N_6416,N_6202);
nor U8852 (N_8852,N_6228,N_7303);
or U8853 (N_8853,N_6518,N_6751);
nor U8854 (N_8854,N_7674,N_7699);
nor U8855 (N_8855,N_7936,N_6254);
nand U8856 (N_8856,N_7407,N_7451);
nor U8857 (N_8857,N_7486,N_7095);
nand U8858 (N_8858,N_6950,N_6373);
nand U8859 (N_8859,N_6065,N_7497);
nor U8860 (N_8860,N_7439,N_6993);
or U8861 (N_8861,N_6618,N_7348);
nand U8862 (N_8862,N_6773,N_6775);
nor U8863 (N_8863,N_6577,N_6062);
and U8864 (N_8864,N_7769,N_7694);
and U8865 (N_8865,N_7736,N_6243);
nor U8866 (N_8866,N_7351,N_7289);
or U8867 (N_8867,N_7908,N_6947);
and U8868 (N_8868,N_6560,N_6462);
nand U8869 (N_8869,N_6883,N_7785);
and U8870 (N_8870,N_7237,N_7162);
or U8871 (N_8871,N_6028,N_6250);
and U8872 (N_8872,N_7999,N_7686);
nor U8873 (N_8873,N_7117,N_6433);
nor U8874 (N_8874,N_7364,N_6706);
nor U8875 (N_8875,N_7251,N_6584);
and U8876 (N_8876,N_7471,N_7521);
nand U8877 (N_8877,N_7983,N_6693);
or U8878 (N_8878,N_6519,N_6051);
nor U8879 (N_8879,N_6908,N_7943);
or U8880 (N_8880,N_6690,N_7068);
and U8881 (N_8881,N_6146,N_6485);
nor U8882 (N_8882,N_6742,N_6912);
and U8883 (N_8883,N_7492,N_7188);
nand U8884 (N_8884,N_6423,N_6764);
or U8885 (N_8885,N_6805,N_7814);
nor U8886 (N_8886,N_7816,N_7561);
nand U8887 (N_8887,N_7889,N_7544);
or U8888 (N_8888,N_6642,N_7992);
nand U8889 (N_8889,N_7171,N_6923);
or U8890 (N_8890,N_6536,N_6369);
and U8891 (N_8891,N_7798,N_7215);
or U8892 (N_8892,N_6284,N_7051);
nor U8893 (N_8893,N_7039,N_6124);
or U8894 (N_8894,N_7106,N_7975);
and U8895 (N_8895,N_6269,N_6535);
nor U8896 (N_8896,N_6407,N_6154);
nand U8897 (N_8897,N_7837,N_7173);
nand U8898 (N_8898,N_6688,N_6464);
nor U8899 (N_8899,N_6271,N_6286);
nand U8900 (N_8900,N_6836,N_7551);
or U8901 (N_8901,N_6044,N_6907);
and U8902 (N_8902,N_7628,N_6603);
or U8903 (N_8903,N_6794,N_7764);
nand U8904 (N_8904,N_6411,N_7748);
nand U8905 (N_8905,N_6363,N_7514);
and U8906 (N_8906,N_6953,N_7100);
and U8907 (N_8907,N_7873,N_6515);
and U8908 (N_8908,N_6934,N_7007);
nand U8909 (N_8909,N_7960,N_6327);
nor U8910 (N_8910,N_7349,N_7829);
nand U8911 (N_8911,N_6985,N_6937);
and U8912 (N_8912,N_7083,N_6701);
nor U8913 (N_8913,N_7754,N_7155);
and U8914 (N_8914,N_7653,N_7974);
and U8915 (N_8915,N_7470,N_7737);
or U8916 (N_8916,N_7071,N_7115);
and U8917 (N_8917,N_7049,N_7781);
and U8918 (N_8918,N_7948,N_6007);
nor U8919 (N_8919,N_7864,N_6940);
nor U8920 (N_8920,N_7522,N_7277);
and U8921 (N_8921,N_6163,N_7129);
xnor U8922 (N_8922,N_7037,N_6622);
or U8923 (N_8923,N_6175,N_7592);
or U8924 (N_8924,N_7849,N_6184);
or U8925 (N_8925,N_6270,N_7777);
and U8926 (N_8926,N_7775,N_6479);
or U8927 (N_8927,N_7570,N_7916);
or U8928 (N_8928,N_7196,N_6968);
or U8929 (N_8929,N_6900,N_7782);
nor U8930 (N_8930,N_7600,N_6321);
nand U8931 (N_8931,N_6522,N_6410);
nand U8932 (N_8932,N_7416,N_7669);
nor U8933 (N_8933,N_6073,N_7122);
nand U8934 (N_8934,N_7473,N_6304);
xor U8935 (N_8935,N_6988,N_7132);
nor U8936 (N_8936,N_7914,N_6450);
or U8937 (N_8937,N_6442,N_6460);
nand U8938 (N_8938,N_7273,N_7825);
nor U8939 (N_8939,N_7951,N_7012);
nand U8940 (N_8940,N_6350,N_6388);
and U8941 (N_8941,N_7491,N_7545);
nor U8942 (N_8942,N_6066,N_7988);
and U8943 (N_8943,N_7586,N_6819);
or U8944 (N_8944,N_6654,N_7909);
nor U8945 (N_8945,N_6036,N_7437);
and U8946 (N_8946,N_6748,N_7562);
or U8947 (N_8947,N_7431,N_6185);
nand U8948 (N_8948,N_7886,N_7823);
or U8949 (N_8949,N_7294,N_6132);
nor U8950 (N_8950,N_6899,N_6973);
nand U8951 (N_8951,N_6017,N_7047);
and U8952 (N_8952,N_6909,N_7339);
nand U8953 (N_8953,N_7563,N_7493);
and U8954 (N_8954,N_6079,N_6844);
or U8955 (N_8955,N_6445,N_6064);
and U8956 (N_8956,N_6337,N_6148);
nand U8957 (N_8957,N_7467,N_7647);
nand U8958 (N_8958,N_7219,N_7502);
and U8959 (N_8959,N_7618,N_6888);
and U8960 (N_8960,N_6025,N_6743);
and U8961 (N_8961,N_6829,N_7340);
nor U8962 (N_8962,N_6112,N_6281);
nor U8963 (N_8963,N_7323,N_6870);
nor U8964 (N_8964,N_7366,N_6224);
nand U8965 (N_8965,N_6344,N_7035);
nand U8966 (N_8966,N_7552,N_7827);
or U8967 (N_8967,N_7022,N_7050);
and U8968 (N_8968,N_6236,N_7919);
nor U8969 (N_8969,N_7989,N_6303);
and U8970 (N_8970,N_7824,N_6382);
and U8971 (N_8971,N_7329,N_6288);
and U8972 (N_8972,N_7213,N_7202);
nand U8973 (N_8973,N_6195,N_7648);
and U8974 (N_8974,N_6833,N_6399);
or U8975 (N_8975,N_6631,N_6681);
or U8976 (N_8976,N_6297,N_7412);
and U8977 (N_8977,N_6548,N_6189);
xnor U8978 (N_8978,N_7250,N_7061);
nor U8979 (N_8979,N_6865,N_7945);
nand U8980 (N_8980,N_6886,N_6623);
or U8981 (N_8981,N_6911,N_7408);
nor U8982 (N_8982,N_7865,N_6364);
nor U8983 (N_8983,N_6592,N_7529);
and U8984 (N_8984,N_7810,N_7032);
xnor U8985 (N_8985,N_7385,N_7884);
or U8986 (N_8986,N_7209,N_7419);
and U8987 (N_8987,N_6312,N_7263);
or U8988 (N_8988,N_6510,N_6625);
or U8989 (N_8989,N_7121,N_7091);
and U8990 (N_8990,N_6384,N_7396);
and U8991 (N_8991,N_6996,N_6251);
and U8992 (N_8992,N_7710,N_7911);
and U8993 (N_8993,N_6447,N_6325);
and U8994 (N_8994,N_7953,N_7248);
or U8995 (N_8995,N_7701,N_6769);
or U8996 (N_8996,N_7130,N_6137);
or U8997 (N_8997,N_7680,N_6890);
nor U8998 (N_8998,N_6811,N_6613);
nand U8999 (N_8999,N_7228,N_7572);
or U9000 (N_9000,N_7330,N_7386);
nor U9001 (N_9001,N_7490,N_7597);
and U9002 (N_9002,N_6790,N_6538);
nand U9003 (N_9003,N_7401,N_6616);
or U9004 (N_9004,N_6323,N_7174);
and U9005 (N_9005,N_7677,N_7669);
or U9006 (N_9006,N_6749,N_6973);
and U9007 (N_9007,N_7480,N_6957);
or U9008 (N_9008,N_6218,N_7745);
nand U9009 (N_9009,N_6305,N_6361);
and U9010 (N_9010,N_6470,N_7163);
nor U9011 (N_9011,N_7008,N_7756);
or U9012 (N_9012,N_7468,N_7625);
nand U9013 (N_9013,N_7671,N_6191);
or U9014 (N_9014,N_6517,N_6446);
or U9015 (N_9015,N_6074,N_6222);
nand U9016 (N_9016,N_6447,N_7290);
nand U9017 (N_9017,N_6943,N_7381);
and U9018 (N_9018,N_6142,N_6325);
nand U9019 (N_9019,N_7770,N_7551);
nand U9020 (N_9020,N_6564,N_6037);
nor U9021 (N_9021,N_7674,N_7332);
and U9022 (N_9022,N_7066,N_7765);
nor U9023 (N_9023,N_7341,N_7261);
nor U9024 (N_9024,N_7082,N_6935);
nor U9025 (N_9025,N_7350,N_7183);
nor U9026 (N_9026,N_6976,N_7345);
and U9027 (N_9027,N_7629,N_6725);
nor U9028 (N_9028,N_6470,N_6850);
and U9029 (N_9029,N_6499,N_7826);
nor U9030 (N_9030,N_6676,N_7086);
nand U9031 (N_9031,N_7631,N_6458);
or U9032 (N_9032,N_7447,N_6330);
nor U9033 (N_9033,N_7715,N_7483);
and U9034 (N_9034,N_6211,N_7785);
and U9035 (N_9035,N_6062,N_6230);
nand U9036 (N_9036,N_6016,N_7444);
nand U9037 (N_9037,N_7585,N_7493);
nor U9038 (N_9038,N_6750,N_7984);
and U9039 (N_9039,N_7356,N_7476);
and U9040 (N_9040,N_7734,N_6448);
and U9041 (N_9041,N_7224,N_7474);
nor U9042 (N_9042,N_6207,N_6264);
and U9043 (N_9043,N_6646,N_6933);
nor U9044 (N_9044,N_7661,N_7465);
and U9045 (N_9045,N_6774,N_7160);
nand U9046 (N_9046,N_7434,N_7099);
nand U9047 (N_9047,N_6403,N_6617);
nor U9048 (N_9048,N_6879,N_7347);
and U9049 (N_9049,N_6918,N_6977);
nand U9050 (N_9050,N_6380,N_6161);
or U9051 (N_9051,N_7182,N_7437);
nor U9052 (N_9052,N_7193,N_6208);
nor U9053 (N_9053,N_7024,N_6483);
nand U9054 (N_9054,N_7999,N_7989);
or U9055 (N_9055,N_6582,N_6132);
and U9056 (N_9056,N_6328,N_6874);
nor U9057 (N_9057,N_7215,N_6694);
nor U9058 (N_9058,N_6833,N_7773);
nand U9059 (N_9059,N_7710,N_6854);
or U9060 (N_9060,N_6476,N_7671);
nor U9061 (N_9061,N_7820,N_7424);
xor U9062 (N_9062,N_6688,N_7508);
nand U9063 (N_9063,N_7521,N_7187);
nand U9064 (N_9064,N_7343,N_7279);
nor U9065 (N_9065,N_6530,N_7494);
nand U9066 (N_9066,N_6444,N_7022);
or U9067 (N_9067,N_7377,N_6954);
xnor U9068 (N_9068,N_6282,N_6742);
and U9069 (N_9069,N_6330,N_6392);
nor U9070 (N_9070,N_7815,N_6535);
or U9071 (N_9071,N_6792,N_7164);
nor U9072 (N_9072,N_6923,N_6045);
nor U9073 (N_9073,N_7834,N_6103);
or U9074 (N_9074,N_7464,N_6695);
nand U9075 (N_9075,N_7229,N_7965);
nor U9076 (N_9076,N_6778,N_7649);
or U9077 (N_9077,N_6739,N_6237);
and U9078 (N_9078,N_6015,N_6848);
nand U9079 (N_9079,N_7428,N_7044);
nor U9080 (N_9080,N_6337,N_6703);
or U9081 (N_9081,N_7883,N_6926);
and U9082 (N_9082,N_7992,N_7566);
or U9083 (N_9083,N_7063,N_7630);
and U9084 (N_9084,N_7477,N_7099);
and U9085 (N_9085,N_6943,N_6985);
nor U9086 (N_9086,N_6110,N_6509);
and U9087 (N_9087,N_6963,N_7534);
nand U9088 (N_9088,N_7640,N_7134);
nand U9089 (N_9089,N_7685,N_7887);
nand U9090 (N_9090,N_7200,N_7252);
or U9091 (N_9091,N_7405,N_7792);
xor U9092 (N_9092,N_7820,N_6229);
nor U9093 (N_9093,N_6306,N_6289);
nor U9094 (N_9094,N_6824,N_6040);
and U9095 (N_9095,N_7418,N_6302);
and U9096 (N_9096,N_7251,N_6052);
or U9097 (N_9097,N_7682,N_7385);
nand U9098 (N_9098,N_7694,N_6561);
or U9099 (N_9099,N_6652,N_6617);
or U9100 (N_9100,N_7721,N_6434);
or U9101 (N_9101,N_7000,N_6104);
nand U9102 (N_9102,N_7839,N_7265);
or U9103 (N_9103,N_6261,N_6052);
or U9104 (N_9104,N_7420,N_7266);
nand U9105 (N_9105,N_7208,N_7186);
and U9106 (N_9106,N_7397,N_6569);
nor U9107 (N_9107,N_6978,N_7694);
or U9108 (N_9108,N_7329,N_6025);
and U9109 (N_9109,N_6509,N_6452);
xor U9110 (N_9110,N_6513,N_6067);
or U9111 (N_9111,N_7926,N_6587);
nor U9112 (N_9112,N_6610,N_7527);
nand U9113 (N_9113,N_7091,N_7967);
nand U9114 (N_9114,N_6989,N_7988);
or U9115 (N_9115,N_7859,N_7200);
or U9116 (N_9116,N_6862,N_6508);
nor U9117 (N_9117,N_7003,N_6419);
or U9118 (N_9118,N_6612,N_7090);
nand U9119 (N_9119,N_6273,N_7837);
nor U9120 (N_9120,N_7126,N_7019);
or U9121 (N_9121,N_7488,N_6503);
and U9122 (N_9122,N_7939,N_6351);
nor U9123 (N_9123,N_7735,N_7378);
nor U9124 (N_9124,N_6394,N_6929);
or U9125 (N_9125,N_6555,N_6915);
nand U9126 (N_9126,N_7548,N_6434);
nand U9127 (N_9127,N_7680,N_7541);
or U9128 (N_9128,N_6221,N_6751);
and U9129 (N_9129,N_7617,N_7130);
nand U9130 (N_9130,N_6555,N_6762);
or U9131 (N_9131,N_7725,N_6782);
nor U9132 (N_9132,N_7273,N_7247);
xnor U9133 (N_9133,N_7688,N_7235);
or U9134 (N_9134,N_7215,N_7713);
nor U9135 (N_9135,N_6834,N_7901);
and U9136 (N_9136,N_6164,N_7542);
nand U9137 (N_9137,N_6105,N_6937);
nand U9138 (N_9138,N_7300,N_6059);
nand U9139 (N_9139,N_6320,N_6351);
nand U9140 (N_9140,N_7857,N_7152);
or U9141 (N_9141,N_7981,N_7965);
nand U9142 (N_9142,N_6162,N_6394);
nand U9143 (N_9143,N_6263,N_6881);
and U9144 (N_9144,N_7259,N_7436);
nand U9145 (N_9145,N_7870,N_6520);
or U9146 (N_9146,N_6188,N_7506);
and U9147 (N_9147,N_6501,N_7250);
or U9148 (N_9148,N_6823,N_6614);
xor U9149 (N_9149,N_6494,N_6192);
nand U9150 (N_9150,N_7906,N_6380);
nand U9151 (N_9151,N_7618,N_7492);
and U9152 (N_9152,N_6769,N_7895);
nor U9153 (N_9153,N_7222,N_7896);
and U9154 (N_9154,N_7365,N_6607);
or U9155 (N_9155,N_6448,N_6252);
or U9156 (N_9156,N_7388,N_7546);
or U9157 (N_9157,N_6227,N_7340);
nand U9158 (N_9158,N_7777,N_7377);
nor U9159 (N_9159,N_7509,N_7920);
or U9160 (N_9160,N_7564,N_6100);
nand U9161 (N_9161,N_7295,N_7442);
nor U9162 (N_9162,N_7621,N_7151);
nor U9163 (N_9163,N_6153,N_6981);
nor U9164 (N_9164,N_6266,N_7359);
nand U9165 (N_9165,N_7560,N_7567);
nand U9166 (N_9166,N_6713,N_7578);
and U9167 (N_9167,N_7875,N_7175);
and U9168 (N_9168,N_6388,N_7319);
nand U9169 (N_9169,N_6460,N_7776);
nand U9170 (N_9170,N_6455,N_7975);
and U9171 (N_9171,N_6380,N_6033);
nand U9172 (N_9172,N_7019,N_7091);
nor U9173 (N_9173,N_6556,N_6594);
or U9174 (N_9174,N_7109,N_6935);
nand U9175 (N_9175,N_7278,N_7522);
and U9176 (N_9176,N_6098,N_6115);
nor U9177 (N_9177,N_7865,N_6367);
and U9178 (N_9178,N_7563,N_7360);
nand U9179 (N_9179,N_7958,N_7287);
nand U9180 (N_9180,N_7381,N_7361);
or U9181 (N_9181,N_7856,N_6655);
nor U9182 (N_9182,N_7107,N_6739);
nand U9183 (N_9183,N_7301,N_7011);
nand U9184 (N_9184,N_6395,N_7960);
or U9185 (N_9185,N_7984,N_6833);
and U9186 (N_9186,N_7348,N_7371);
and U9187 (N_9187,N_7785,N_6401);
nand U9188 (N_9188,N_7474,N_7908);
or U9189 (N_9189,N_6838,N_7192);
or U9190 (N_9190,N_7283,N_6363);
and U9191 (N_9191,N_6456,N_7653);
or U9192 (N_9192,N_6675,N_7513);
nand U9193 (N_9193,N_6964,N_6088);
or U9194 (N_9194,N_6317,N_7709);
nor U9195 (N_9195,N_6089,N_7623);
nand U9196 (N_9196,N_6030,N_7327);
nor U9197 (N_9197,N_6240,N_7383);
nand U9198 (N_9198,N_6784,N_7557);
or U9199 (N_9199,N_6647,N_6203);
nand U9200 (N_9200,N_6250,N_7323);
nor U9201 (N_9201,N_7340,N_7317);
nand U9202 (N_9202,N_7677,N_7232);
nor U9203 (N_9203,N_7482,N_6846);
and U9204 (N_9204,N_6758,N_7889);
and U9205 (N_9205,N_7919,N_7986);
or U9206 (N_9206,N_6929,N_7784);
nand U9207 (N_9207,N_7566,N_7656);
or U9208 (N_9208,N_7462,N_6812);
and U9209 (N_9209,N_7108,N_6230);
nor U9210 (N_9210,N_6170,N_6371);
and U9211 (N_9211,N_6250,N_6439);
or U9212 (N_9212,N_7918,N_6270);
or U9213 (N_9213,N_7606,N_7087);
nor U9214 (N_9214,N_6920,N_7004);
or U9215 (N_9215,N_7340,N_7036);
and U9216 (N_9216,N_7945,N_7578);
or U9217 (N_9217,N_7139,N_7333);
nor U9218 (N_9218,N_7984,N_6036);
nor U9219 (N_9219,N_6752,N_7219);
nand U9220 (N_9220,N_6754,N_7870);
nand U9221 (N_9221,N_7540,N_7382);
and U9222 (N_9222,N_7195,N_6905);
nor U9223 (N_9223,N_7627,N_7168);
or U9224 (N_9224,N_7539,N_7331);
and U9225 (N_9225,N_6252,N_7039);
nand U9226 (N_9226,N_7223,N_7889);
or U9227 (N_9227,N_7974,N_7030);
and U9228 (N_9228,N_7886,N_6317);
and U9229 (N_9229,N_6362,N_7280);
nor U9230 (N_9230,N_7821,N_6408);
nand U9231 (N_9231,N_7552,N_7910);
nand U9232 (N_9232,N_7006,N_6423);
nor U9233 (N_9233,N_7084,N_6988);
and U9234 (N_9234,N_7927,N_6667);
nand U9235 (N_9235,N_7553,N_6530);
nor U9236 (N_9236,N_6312,N_7841);
or U9237 (N_9237,N_7035,N_6569);
nor U9238 (N_9238,N_6559,N_7900);
and U9239 (N_9239,N_7285,N_7253);
nor U9240 (N_9240,N_6550,N_7812);
or U9241 (N_9241,N_6587,N_6727);
nor U9242 (N_9242,N_6415,N_7050);
or U9243 (N_9243,N_6076,N_7640);
nor U9244 (N_9244,N_6340,N_7638);
and U9245 (N_9245,N_7893,N_7809);
xnor U9246 (N_9246,N_7454,N_6353);
and U9247 (N_9247,N_6350,N_6522);
and U9248 (N_9248,N_7316,N_6251);
nor U9249 (N_9249,N_7210,N_6672);
and U9250 (N_9250,N_6793,N_7615);
or U9251 (N_9251,N_7364,N_7008);
nand U9252 (N_9252,N_6453,N_6170);
or U9253 (N_9253,N_6267,N_7503);
and U9254 (N_9254,N_6896,N_7475);
nand U9255 (N_9255,N_6611,N_7891);
nand U9256 (N_9256,N_7701,N_6846);
nand U9257 (N_9257,N_7869,N_7861);
nor U9258 (N_9258,N_7302,N_7386);
and U9259 (N_9259,N_6705,N_7330);
nand U9260 (N_9260,N_6690,N_6743);
nand U9261 (N_9261,N_6282,N_7887);
and U9262 (N_9262,N_6000,N_6676);
or U9263 (N_9263,N_6993,N_6393);
and U9264 (N_9264,N_6324,N_7074);
nand U9265 (N_9265,N_7710,N_6593);
or U9266 (N_9266,N_7891,N_6753);
or U9267 (N_9267,N_7878,N_7797);
and U9268 (N_9268,N_6305,N_7979);
and U9269 (N_9269,N_7066,N_6763);
or U9270 (N_9270,N_6475,N_7290);
and U9271 (N_9271,N_6014,N_6780);
xor U9272 (N_9272,N_7324,N_6475);
or U9273 (N_9273,N_6661,N_6804);
and U9274 (N_9274,N_7517,N_7987);
and U9275 (N_9275,N_6405,N_6558);
nor U9276 (N_9276,N_6876,N_7535);
and U9277 (N_9277,N_6227,N_7280);
nand U9278 (N_9278,N_6693,N_6102);
or U9279 (N_9279,N_7602,N_7133);
nand U9280 (N_9280,N_6960,N_6774);
nor U9281 (N_9281,N_6326,N_6591);
nand U9282 (N_9282,N_6160,N_7084);
nor U9283 (N_9283,N_7613,N_7538);
and U9284 (N_9284,N_6952,N_7649);
and U9285 (N_9285,N_7487,N_7313);
or U9286 (N_9286,N_7406,N_6920);
or U9287 (N_9287,N_6649,N_7293);
and U9288 (N_9288,N_7879,N_6738);
or U9289 (N_9289,N_6868,N_6597);
nor U9290 (N_9290,N_7186,N_6015);
nor U9291 (N_9291,N_7414,N_6979);
and U9292 (N_9292,N_7327,N_6467);
and U9293 (N_9293,N_6196,N_7528);
xor U9294 (N_9294,N_6423,N_6499);
and U9295 (N_9295,N_7916,N_6095);
nor U9296 (N_9296,N_7660,N_6096);
nor U9297 (N_9297,N_7900,N_6079);
nor U9298 (N_9298,N_7374,N_6199);
nor U9299 (N_9299,N_7902,N_7264);
nand U9300 (N_9300,N_6308,N_7358);
and U9301 (N_9301,N_7262,N_6849);
nor U9302 (N_9302,N_7395,N_7535);
nand U9303 (N_9303,N_6293,N_7044);
nand U9304 (N_9304,N_7967,N_7339);
or U9305 (N_9305,N_6975,N_6015);
nand U9306 (N_9306,N_7978,N_6765);
nor U9307 (N_9307,N_7855,N_6306);
or U9308 (N_9308,N_6226,N_7444);
nor U9309 (N_9309,N_6901,N_6518);
or U9310 (N_9310,N_6023,N_6479);
nor U9311 (N_9311,N_7371,N_7965);
nand U9312 (N_9312,N_7181,N_6515);
nor U9313 (N_9313,N_7327,N_6526);
or U9314 (N_9314,N_6085,N_6191);
or U9315 (N_9315,N_7233,N_7208);
and U9316 (N_9316,N_6795,N_6898);
and U9317 (N_9317,N_6730,N_6915);
nor U9318 (N_9318,N_6688,N_7056);
or U9319 (N_9319,N_6004,N_7855);
nand U9320 (N_9320,N_6516,N_7987);
nand U9321 (N_9321,N_6502,N_7438);
nand U9322 (N_9322,N_6003,N_7278);
nand U9323 (N_9323,N_6714,N_6354);
nor U9324 (N_9324,N_6903,N_6495);
nand U9325 (N_9325,N_6012,N_7642);
nand U9326 (N_9326,N_7626,N_6250);
nor U9327 (N_9327,N_6416,N_6938);
or U9328 (N_9328,N_6798,N_7055);
or U9329 (N_9329,N_6610,N_6355);
nand U9330 (N_9330,N_6759,N_6745);
and U9331 (N_9331,N_7198,N_6454);
nand U9332 (N_9332,N_6481,N_6574);
nor U9333 (N_9333,N_7339,N_7315);
nand U9334 (N_9334,N_7854,N_6228);
or U9335 (N_9335,N_7691,N_7746);
nor U9336 (N_9336,N_6346,N_7282);
or U9337 (N_9337,N_7445,N_6555);
nand U9338 (N_9338,N_6472,N_7131);
nor U9339 (N_9339,N_6092,N_6934);
nand U9340 (N_9340,N_7393,N_7540);
and U9341 (N_9341,N_6908,N_7660);
nand U9342 (N_9342,N_6555,N_6276);
and U9343 (N_9343,N_7723,N_6777);
nand U9344 (N_9344,N_6225,N_7126);
nor U9345 (N_9345,N_6963,N_7250);
xor U9346 (N_9346,N_7430,N_6488);
and U9347 (N_9347,N_7750,N_7887);
nor U9348 (N_9348,N_6375,N_7849);
or U9349 (N_9349,N_6478,N_7089);
nor U9350 (N_9350,N_6119,N_6934);
nand U9351 (N_9351,N_7972,N_7273);
and U9352 (N_9352,N_6334,N_7890);
nand U9353 (N_9353,N_6574,N_6181);
and U9354 (N_9354,N_7814,N_6357);
nor U9355 (N_9355,N_6849,N_6987);
xnor U9356 (N_9356,N_6130,N_6082);
or U9357 (N_9357,N_6712,N_7300);
or U9358 (N_9358,N_7855,N_6747);
nor U9359 (N_9359,N_7890,N_6207);
nand U9360 (N_9360,N_7183,N_6755);
or U9361 (N_9361,N_6193,N_7525);
and U9362 (N_9362,N_6384,N_7575);
nor U9363 (N_9363,N_6900,N_6074);
or U9364 (N_9364,N_7842,N_7150);
or U9365 (N_9365,N_7656,N_7827);
or U9366 (N_9366,N_6290,N_6493);
nand U9367 (N_9367,N_7136,N_7441);
nand U9368 (N_9368,N_6844,N_7210);
nor U9369 (N_9369,N_7099,N_6081);
nand U9370 (N_9370,N_6716,N_7597);
and U9371 (N_9371,N_7363,N_7828);
nor U9372 (N_9372,N_7724,N_7646);
or U9373 (N_9373,N_7560,N_7918);
nor U9374 (N_9374,N_6002,N_6937);
nor U9375 (N_9375,N_6502,N_6366);
and U9376 (N_9376,N_6051,N_7639);
nand U9377 (N_9377,N_6997,N_7886);
nor U9378 (N_9378,N_6746,N_6977);
or U9379 (N_9379,N_6875,N_7541);
nand U9380 (N_9380,N_6315,N_7012);
nor U9381 (N_9381,N_7292,N_7059);
nand U9382 (N_9382,N_6635,N_6050);
or U9383 (N_9383,N_6598,N_6190);
and U9384 (N_9384,N_6390,N_7533);
or U9385 (N_9385,N_7515,N_7280);
nand U9386 (N_9386,N_6869,N_6318);
nor U9387 (N_9387,N_7884,N_7597);
or U9388 (N_9388,N_6479,N_6755);
and U9389 (N_9389,N_7394,N_6006);
and U9390 (N_9390,N_7937,N_7727);
or U9391 (N_9391,N_7435,N_6302);
or U9392 (N_9392,N_6334,N_6788);
or U9393 (N_9393,N_7807,N_7072);
nand U9394 (N_9394,N_6918,N_7686);
and U9395 (N_9395,N_7346,N_7735);
or U9396 (N_9396,N_6704,N_7795);
or U9397 (N_9397,N_7356,N_6497);
and U9398 (N_9398,N_7618,N_6238);
nor U9399 (N_9399,N_6183,N_6785);
and U9400 (N_9400,N_6573,N_7251);
nor U9401 (N_9401,N_6232,N_7541);
and U9402 (N_9402,N_7251,N_6361);
and U9403 (N_9403,N_6255,N_7608);
or U9404 (N_9404,N_7850,N_7913);
and U9405 (N_9405,N_6651,N_7493);
and U9406 (N_9406,N_7918,N_6947);
or U9407 (N_9407,N_6783,N_7988);
and U9408 (N_9408,N_6783,N_7457);
nor U9409 (N_9409,N_6709,N_6813);
nor U9410 (N_9410,N_6052,N_6057);
xnor U9411 (N_9411,N_6230,N_6575);
or U9412 (N_9412,N_7355,N_7755);
and U9413 (N_9413,N_6937,N_7753);
and U9414 (N_9414,N_6505,N_6745);
nor U9415 (N_9415,N_6719,N_7323);
or U9416 (N_9416,N_6903,N_6875);
or U9417 (N_9417,N_6426,N_7233);
and U9418 (N_9418,N_6618,N_6640);
and U9419 (N_9419,N_7367,N_6024);
and U9420 (N_9420,N_6420,N_6306);
nor U9421 (N_9421,N_7138,N_6440);
nor U9422 (N_9422,N_6871,N_7225);
nand U9423 (N_9423,N_6056,N_7468);
nand U9424 (N_9424,N_7019,N_6740);
nor U9425 (N_9425,N_7419,N_6998);
nand U9426 (N_9426,N_7154,N_6635);
or U9427 (N_9427,N_7140,N_7735);
or U9428 (N_9428,N_6857,N_7830);
nor U9429 (N_9429,N_6035,N_6579);
xnor U9430 (N_9430,N_7745,N_7702);
or U9431 (N_9431,N_6955,N_6397);
nor U9432 (N_9432,N_6455,N_7766);
nor U9433 (N_9433,N_7157,N_6415);
or U9434 (N_9434,N_6230,N_7637);
or U9435 (N_9435,N_6978,N_7888);
and U9436 (N_9436,N_6275,N_7115);
and U9437 (N_9437,N_6249,N_7138);
nor U9438 (N_9438,N_7434,N_6062);
or U9439 (N_9439,N_6400,N_7410);
or U9440 (N_9440,N_6104,N_6253);
nor U9441 (N_9441,N_7672,N_7563);
or U9442 (N_9442,N_6865,N_6936);
and U9443 (N_9443,N_6708,N_7538);
and U9444 (N_9444,N_7613,N_7448);
nor U9445 (N_9445,N_6866,N_7417);
or U9446 (N_9446,N_6894,N_7260);
nor U9447 (N_9447,N_6066,N_7991);
or U9448 (N_9448,N_6556,N_7538);
nor U9449 (N_9449,N_7401,N_6304);
nor U9450 (N_9450,N_7547,N_6336);
nor U9451 (N_9451,N_6475,N_6962);
or U9452 (N_9452,N_7345,N_7103);
and U9453 (N_9453,N_7357,N_6265);
and U9454 (N_9454,N_6020,N_7546);
nand U9455 (N_9455,N_6054,N_7947);
nand U9456 (N_9456,N_6465,N_6286);
nand U9457 (N_9457,N_6844,N_7357);
nor U9458 (N_9458,N_6514,N_6355);
or U9459 (N_9459,N_7520,N_7460);
and U9460 (N_9460,N_6496,N_6468);
and U9461 (N_9461,N_6959,N_6966);
or U9462 (N_9462,N_6137,N_6696);
or U9463 (N_9463,N_6905,N_6691);
nand U9464 (N_9464,N_6169,N_6525);
or U9465 (N_9465,N_7309,N_7042);
and U9466 (N_9466,N_7935,N_7925);
or U9467 (N_9467,N_6398,N_6519);
and U9468 (N_9468,N_6248,N_6903);
nor U9469 (N_9469,N_6843,N_7625);
and U9470 (N_9470,N_7338,N_6155);
and U9471 (N_9471,N_6740,N_6217);
and U9472 (N_9472,N_7140,N_6675);
nor U9473 (N_9473,N_7485,N_7580);
and U9474 (N_9474,N_6261,N_7805);
nand U9475 (N_9475,N_7968,N_6089);
and U9476 (N_9476,N_6386,N_6365);
nor U9477 (N_9477,N_7095,N_6157);
and U9478 (N_9478,N_6863,N_7684);
nand U9479 (N_9479,N_6497,N_7525);
or U9480 (N_9480,N_6201,N_6521);
xor U9481 (N_9481,N_6305,N_7091);
nand U9482 (N_9482,N_7311,N_6415);
nand U9483 (N_9483,N_7833,N_7815);
nor U9484 (N_9484,N_7578,N_7094);
nand U9485 (N_9485,N_7708,N_7244);
nand U9486 (N_9486,N_7525,N_7855);
nor U9487 (N_9487,N_7209,N_7429);
or U9488 (N_9488,N_6037,N_6000);
or U9489 (N_9489,N_7306,N_7987);
nor U9490 (N_9490,N_7339,N_7900);
nor U9491 (N_9491,N_6259,N_7234);
and U9492 (N_9492,N_7968,N_6315);
or U9493 (N_9493,N_6411,N_7656);
nand U9494 (N_9494,N_6827,N_7578);
or U9495 (N_9495,N_6289,N_7331);
and U9496 (N_9496,N_7965,N_6065);
and U9497 (N_9497,N_7903,N_6940);
and U9498 (N_9498,N_6951,N_6545);
nor U9499 (N_9499,N_7821,N_7458);
nor U9500 (N_9500,N_6522,N_6891);
or U9501 (N_9501,N_6101,N_7968);
and U9502 (N_9502,N_7442,N_7068);
and U9503 (N_9503,N_6686,N_6555);
and U9504 (N_9504,N_7213,N_7435);
nand U9505 (N_9505,N_6538,N_7112);
nand U9506 (N_9506,N_6872,N_6205);
xor U9507 (N_9507,N_7153,N_6381);
and U9508 (N_9508,N_6626,N_6703);
nor U9509 (N_9509,N_6566,N_7610);
or U9510 (N_9510,N_7480,N_6248);
nor U9511 (N_9511,N_7030,N_6416);
or U9512 (N_9512,N_6554,N_7253);
nor U9513 (N_9513,N_7432,N_6317);
nor U9514 (N_9514,N_6220,N_6018);
or U9515 (N_9515,N_7318,N_7576);
nand U9516 (N_9516,N_7827,N_6914);
or U9517 (N_9517,N_7074,N_6063);
nor U9518 (N_9518,N_7097,N_7183);
or U9519 (N_9519,N_6887,N_6121);
xnor U9520 (N_9520,N_6736,N_7696);
xor U9521 (N_9521,N_6571,N_6034);
nand U9522 (N_9522,N_6977,N_7432);
nand U9523 (N_9523,N_7489,N_7921);
or U9524 (N_9524,N_7237,N_6144);
or U9525 (N_9525,N_6051,N_7729);
or U9526 (N_9526,N_7837,N_7015);
and U9527 (N_9527,N_7451,N_6387);
nand U9528 (N_9528,N_6144,N_6979);
nand U9529 (N_9529,N_7391,N_6170);
nand U9530 (N_9530,N_7576,N_6671);
or U9531 (N_9531,N_7704,N_7785);
or U9532 (N_9532,N_7279,N_7941);
nand U9533 (N_9533,N_7920,N_6703);
nand U9534 (N_9534,N_7029,N_7203);
and U9535 (N_9535,N_6388,N_7966);
nand U9536 (N_9536,N_7603,N_7394);
nand U9537 (N_9537,N_6705,N_6621);
and U9538 (N_9538,N_7438,N_7226);
nand U9539 (N_9539,N_6782,N_6686);
or U9540 (N_9540,N_7996,N_7697);
or U9541 (N_9541,N_7330,N_7655);
nand U9542 (N_9542,N_6402,N_7339);
nand U9543 (N_9543,N_6067,N_6607);
and U9544 (N_9544,N_6296,N_7820);
or U9545 (N_9545,N_7960,N_6247);
xnor U9546 (N_9546,N_6507,N_6595);
nand U9547 (N_9547,N_6057,N_6034);
nor U9548 (N_9548,N_7729,N_7596);
and U9549 (N_9549,N_6679,N_6786);
nor U9550 (N_9550,N_6299,N_7722);
and U9551 (N_9551,N_7286,N_7407);
or U9552 (N_9552,N_6487,N_6824);
nand U9553 (N_9553,N_6992,N_7463);
or U9554 (N_9554,N_6128,N_6047);
nand U9555 (N_9555,N_7424,N_6471);
or U9556 (N_9556,N_7997,N_6453);
nor U9557 (N_9557,N_6569,N_6060);
and U9558 (N_9558,N_6280,N_6722);
or U9559 (N_9559,N_7662,N_7215);
nand U9560 (N_9560,N_6240,N_6268);
nand U9561 (N_9561,N_7166,N_7191);
or U9562 (N_9562,N_7431,N_7259);
or U9563 (N_9563,N_7246,N_7090);
and U9564 (N_9564,N_7446,N_6913);
or U9565 (N_9565,N_6239,N_7490);
nand U9566 (N_9566,N_7359,N_7855);
and U9567 (N_9567,N_7353,N_7659);
and U9568 (N_9568,N_7954,N_6903);
or U9569 (N_9569,N_6613,N_7808);
nor U9570 (N_9570,N_7906,N_7092);
nor U9571 (N_9571,N_7606,N_7502);
or U9572 (N_9572,N_6176,N_7028);
nor U9573 (N_9573,N_7905,N_7383);
or U9574 (N_9574,N_6466,N_6088);
nor U9575 (N_9575,N_7896,N_6202);
or U9576 (N_9576,N_6463,N_7049);
nor U9577 (N_9577,N_6569,N_6140);
nor U9578 (N_9578,N_6101,N_7771);
and U9579 (N_9579,N_7330,N_6723);
or U9580 (N_9580,N_7154,N_6451);
nand U9581 (N_9581,N_7880,N_7365);
or U9582 (N_9582,N_6751,N_6873);
nand U9583 (N_9583,N_7237,N_6836);
nand U9584 (N_9584,N_6833,N_7211);
or U9585 (N_9585,N_7984,N_6636);
and U9586 (N_9586,N_7808,N_7262);
or U9587 (N_9587,N_6474,N_6275);
nor U9588 (N_9588,N_7298,N_6548);
and U9589 (N_9589,N_6261,N_6293);
nor U9590 (N_9590,N_7652,N_6622);
nor U9591 (N_9591,N_6689,N_7500);
and U9592 (N_9592,N_7284,N_6292);
nand U9593 (N_9593,N_7499,N_7725);
or U9594 (N_9594,N_6111,N_7309);
nor U9595 (N_9595,N_6266,N_7435);
and U9596 (N_9596,N_6584,N_6943);
and U9597 (N_9597,N_7264,N_7722);
or U9598 (N_9598,N_6748,N_7618);
and U9599 (N_9599,N_7449,N_6961);
nand U9600 (N_9600,N_6148,N_7455);
or U9601 (N_9601,N_6240,N_7588);
or U9602 (N_9602,N_6007,N_7914);
or U9603 (N_9603,N_7923,N_6067);
or U9604 (N_9604,N_7640,N_6727);
or U9605 (N_9605,N_7634,N_6997);
nor U9606 (N_9606,N_6951,N_6193);
or U9607 (N_9607,N_6744,N_6398);
or U9608 (N_9608,N_7254,N_6222);
nand U9609 (N_9609,N_6754,N_7254);
xnor U9610 (N_9610,N_6444,N_7540);
xnor U9611 (N_9611,N_6356,N_6832);
nor U9612 (N_9612,N_6350,N_6281);
xnor U9613 (N_9613,N_6180,N_6633);
and U9614 (N_9614,N_7295,N_6311);
or U9615 (N_9615,N_7045,N_7572);
and U9616 (N_9616,N_6164,N_7744);
or U9617 (N_9617,N_6350,N_7572);
or U9618 (N_9618,N_7836,N_6977);
or U9619 (N_9619,N_6543,N_7531);
and U9620 (N_9620,N_6969,N_6954);
xor U9621 (N_9621,N_7886,N_6542);
nor U9622 (N_9622,N_6603,N_6400);
or U9623 (N_9623,N_6322,N_7907);
or U9624 (N_9624,N_6561,N_6085);
nand U9625 (N_9625,N_7290,N_6795);
or U9626 (N_9626,N_6281,N_7603);
nand U9627 (N_9627,N_7905,N_6054);
nor U9628 (N_9628,N_7671,N_6752);
and U9629 (N_9629,N_7595,N_6206);
or U9630 (N_9630,N_6138,N_7485);
nand U9631 (N_9631,N_7495,N_6268);
and U9632 (N_9632,N_7992,N_7915);
nand U9633 (N_9633,N_7687,N_6401);
nor U9634 (N_9634,N_7661,N_6100);
or U9635 (N_9635,N_7682,N_7469);
and U9636 (N_9636,N_6442,N_7342);
and U9637 (N_9637,N_6465,N_7590);
nor U9638 (N_9638,N_6637,N_6887);
or U9639 (N_9639,N_6146,N_6420);
or U9640 (N_9640,N_7183,N_6519);
xnor U9641 (N_9641,N_6344,N_7042);
nor U9642 (N_9642,N_6905,N_7350);
nand U9643 (N_9643,N_7401,N_7155);
or U9644 (N_9644,N_6665,N_7609);
nor U9645 (N_9645,N_7265,N_6338);
nand U9646 (N_9646,N_6030,N_7226);
nand U9647 (N_9647,N_6456,N_6728);
nand U9648 (N_9648,N_7050,N_7456);
and U9649 (N_9649,N_6532,N_6943);
nand U9650 (N_9650,N_6762,N_6342);
nand U9651 (N_9651,N_7396,N_6473);
nand U9652 (N_9652,N_7941,N_6011);
nand U9653 (N_9653,N_6458,N_6046);
nor U9654 (N_9654,N_7900,N_7228);
or U9655 (N_9655,N_7456,N_6557);
or U9656 (N_9656,N_7804,N_6749);
or U9657 (N_9657,N_6700,N_6697);
and U9658 (N_9658,N_6258,N_6976);
and U9659 (N_9659,N_7296,N_7868);
nor U9660 (N_9660,N_7718,N_6321);
and U9661 (N_9661,N_7833,N_6635);
nand U9662 (N_9662,N_6505,N_7727);
nor U9663 (N_9663,N_7797,N_7752);
nand U9664 (N_9664,N_7579,N_7115);
nand U9665 (N_9665,N_6727,N_6615);
nand U9666 (N_9666,N_7436,N_6268);
nor U9667 (N_9667,N_7849,N_6182);
nor U9668 (N_9668,N_6107,N_6880);
nor U9669 (N_9669,N_7336,N_7849);
nand U9670 (N_9670,N_7000,N_6187);
and U9671 (N_9671,N_6809,N_7369);
or U9672 (N_9672,N_7773,N_6997);
nor U9673 (N_9673,N_6947,N_7978);
nand U9674 (N_9674,N_7730,N_6950);
nand U9675 (N_9675,N_7294,N_6548);
nor U9676 (N_9676,N_6377,N_7151);
nand U9677 (N_9677,N_6884,N_7684);
nand U9678 (N_9678,N_6638,N_6281);
and U9679 (N_9679,N_7333,N_6341);
or U9680 (N_9680,N_6473,N_6359);
nand U9681 (N_9681,N_6592,N_6114);
or U9682 (N_9682,N_6731,N_7941);
or U9683 (N_9683,N_6366,N_7570);
or U9684 (N_9684,N_7098,N_7923);
xor U9685 (N_9685,N_6202,N_6449);
nand U9686 (N_9686,N_7357,N_6022);
nand U9687 (N_9687,N_7405,N_6538);
and U9688 (N_9688,N_6169,N_6067);
and U9689 (N_9689,N_6473,N_7355);
and U9690 (N_9690,N_7798,N_6730);
xor U9691 (N_9691,N_6460,N_7788);
and U9692 (N_9692,N_6968,N_7771);
and U9693 (N_9693,N_6679,N_7655);
and U9694 (N_9694,N_7798,N_7461);
nand U9695 (N_9695,N_7072,N_6304);
nor U9696 (N_9696,N_7859,N_7013);
or U9697 (N_9697,N_6372,N_7331);
and U9698 (N_9698,N_6543,N_7342);
or U9699 (N_9699,N_7277,N_7695);
and U9700 (N_9700,N_7954,N_6790);
nand U9701 (N_9701,N_6353,N_6920);
xor U9702 (N_9702,N_7427,N_7608);
nand U9703 (N_9703,N_7711,N_6977);
and U9704 (N_9704,N_6384,N_6631);
or U9705 (N_9705,N_6977,N_6874);
xnor U9706 (N_9706,N_7082,N_6792);
nor U9707 (N_9707,N_7782,N_6790);
and U9708 (N_9708,N_7440,N_6774);
nand U9709 (N_9709,N_7443,N_7801);
and U9710 (N_9710,N_6229,N_6358);
and U9711 (N_9711,N_6976,N_7073);
and U9712 (N_9712,N_6703,N_7501);
and U9713 (N_9713,N_6790,N_7931);
nand U9714 (N_9714,N_6558,N_6518);
nor U9715 (N_9715,N_7559,N_6843);
nor U9716 (N_9716,N_6075,N_7228);
nor U9717 (N_9717,N_6151,N_6460);
nand U9718 (N_9718,N_6976,N_6483);
and U9719 (N_9719,N_6212,N_6728);
nand U9720 (N_9720,N_6603,N_7827);
and U9721 (N_9721,N_7884,N_7715);
nor U9722 (N_9722,N_7409,N_6684);
nand U9723 (N_9723,N_6147,N_7407);
or U9724 (N_9724,N_7537,N_6735);
nor U9725 (N_9725,N_6038,N_7030);
and U9726 (N_9726,N_7965,N_7830);
nor U9727 (N_9727,N_7013,N_6364);
nor U9728 (N_9728,N_7662,N_7306);
nor U9729 (N_9729,N_7518,N_7209);
nor U9730 (N_9730,N_6041,N_7523);
and U9731 (N_9731,N_6980,N_7696);
and U9732 (N_9732,N_6370,N_7075);
and U9733 (N_9733,N_6361,N_7302);
and U9734 (N_9734,N_7804,N_6351);
nor U9735 (N_9735,N_7876,N_6189);
nand U9736 (N_9736,N_6306,N_6913);
or U9737 (N_9737,N_7434,N_7598);
nor U9738 (N_9738,N_6160,N_6412);
nand U9739 (N_9739,N_7514,N_7699);
nor U9740 (N_9740,N_6470,N_7697);
or U9741 (N_9741,N_6417,N_6544);
nand U9742 (N_9742,N_6653,N_7945);
or U9743 (N_9743,N_7076,N_6596);
nor U9744 (N_9744,N_6687,N_7685);
and U9745 (N_9745,N_7939,N_7769);
nand U9746 (N_9746,N_7774,N_7393);
and U9747 (N_9747,N_6152,N_6826);
nand U9748 (N_9748,N_6181,N_6779);
and U9749 (N_9749,N_6673,N_6996);
or U9750 (N_9750,N_6120,N_6020);
and U9751 (N_9751,N_6800,N_7213);
nand U9752 (N_9752,N_7223,N_7356);
or U9753 (N_9753,N_7096,N_6395);
nand U9754 (N_9754,N_7382,N_7454);
nand U9755 (N_9755,N_6560,N_7746);
or U9756 (N_9756,N_6565,N_6378);
nor U9757 (N_9757,N_7067,N_7723);
nand U9758 (N_9758,N_6197,N_6341);
nand U9759 (N_9759,N_7432,N_7752);
nand U9760 (N_9760,N_7383,N_7898);
and U9761 (N_9761,N_7370,N_7777);
nand U9762 (N_9762,N_6848,N_7043);
and U9763 (N_9763,N_6712,N_6033);
nand U9764 (N_9764,N_7758,N_6134);
nor U9765 (N_9765,N_7391,N_7770);
xor U9766 (N_9766,N_7520,N_7011);
nor U9767 (N_9767,N_6388,N_6242);
or U9768 (N_9768,N_7454,N_6140);
nand U9769 (N_9769,N_6526,N_7105);
and U9770 (N_9770,N_6498,N_7155);
nand U9771 (N_9771,N_7418,N_7039);
or U9772 (N_9772,N_7146,N_6664);
and U9773 (N_9773,N_6174,N_6184);
nor U9774 (N_9774,N_7490,N_7272);
or U9775 (N_9775,N_7187,N_6601);
nand U9776 (N_9776,N_7305,N_7883);
and U9777 (N_9777,N_7835,N_7555);
nand U9778 (N_9778,N_7239,N_6149);
nor U9779 (N_9779,N_7673,N_7707);
nor U9780 (N_9780,N_6449,N_6812);
and U9781 (N_9781,N_7591,N_6062);
or U9782 (N_9782,N_6711,N_6919);
nand U9783 (N_9783,N_7901,N_6582);
nand U9784 (N_9784,N_6901,N_7912);
nor U9785 (N_9785,N_7554,N_7448);
or U9786 (N_9786,N_7680,N_6699);
and U9787 (N_9787,N_6481,N_6735);
nand U9788 (N_9788,N_6743,N_7789);
and U9789 (N_9789,N_7407,N_6037);
and U9790 (N_9790,N_7267,N_6323);
nand U9791 (N_9791,N_7469,N_6397);
nand U9792 (N_9792,N_6324,N_7176);
nor U9793 (N_9793,N_6144,N_7483);
xnor U9794 (N_9794,N_6658,N_7401);
and U9795 (N_9795,N_6257,N_6046);
nor U9796 (N_9796,N_6085,N_7638);
nand U9797 (N_9797,N_6147,N_7092);
or U9798 (N_9798,N_6104,N_6022);
and U9799 (N_9799,N_6657,N_6645);
nand U9800 (N_9800,N_6948,N_6583);
nor U9801 (N_9801,N_7331,N_7605);
and U9802 (N_9802,N_6997,N_7504);
nand U9803 (N_9803,N_6445,N_7676);
and U9804 (N_9804,N_7613,N_7061);
or U9805 (N_9805,N_6066,N_7427);
or U9806 (N_9806,N_6486,N_7847);
and U9807 (N_9807,N_6635,N_7579);
or U9808 (N_9808,N_6805,N_7321);
nand U9809 (N_9809,N_7581,N_7689);
and U9810 (N_9810,N_6580,N_6057);
or U9811 (N_9811,N_6544,N_6269);
xor U9812 (N_9812,N_6881,N_7378);
xor U9813 (N_9813,N_6627,N_6078);
xnor U9814 (N_9814,N_7256,N_6017);
or U9815 (N_9815,N_6125,N_7972);
xor U9816 (N_9816,N_7559,N_7555);
or U9817 (N_9817,N_7720,N_7106);
nand U9818 (N_9818,N_7131,N_7037);
nand U9819 (N_9819,N_7630,N_7199);
and U9820 (N_9820,N_6963,N_7883);
nor U9821 (N_9821,N_7447,N_6237);
nor U9822 (N_9822,N_6416,N_6002);
nand U9823 (N_9823,N_6074,N_7905);
xor U9824 (N_9824,N_6256,N_7659);
nor U9825 (N_9825,N_6810,N_6904);
nor U9826 (N_9826,N_6659,N_7793);
and U9827 (N_9827,N_7933,N_6958);
nand U9828 (N_9828,N_6010,N_7958);
and U9829 (N_9829,N_7906,N_7603);
nor U9830 (N_9830,N_7743,N_7558);
nand U9831 (N_9831,N_6399,N_7109);
nand U9832 (N_9832,N_7792,N_7761);
or U9833 (N_9833,N_6080,N_6477);
or U9834 (N_9834,N_7551,N_6535);
nor U9835 (N_9835,N_6601,N_6908);
and U9836 (N_9836,N_6548,N_6874);
nand U9837 (N_9837,N_6572,N_6205);
nand U9838 (N_9838,N_6420,N_7068);
nor U9839 (N_9839,N_7675,N_6196);
and U9840 (N_9840,N_6891,N_6949);
nand U9841 (N_9841,N_7787,N_7650);
or U9842 (N_9842,N_6754,N_7861);
nor U9843 (N_9843,N_7494,N_6411);
and U9844 (N_9844,N_7727,N_7955);
nand U9845 (N_9845,N_6847,N_7432);
nand U9846 (N_9846,N_6373,N_7891);
nand U9847 (N_9847,N_7550,N_7782);
and U9848 (N_9848,N_6343,N_6750);
nor U9849 (N_9849,N_7850,N_7763);
and U9850 (N_9850,N_6576,N_6019);
or U9851 (N_9851,N_6170,N_7946);
and U9852 (N_9852,N_7140,N_7618);
nand U9853 (N_9853,N_6446,N_7495);
nor U9854 (N_9854,N_7321,N_6916);
and U9855 (N_9855,N_7555,N_7240);
nor U9856 (N_9856,N_7052,N_6083);
xor U9857 (N_9857,N_6351,N_7417);
nor U9858 (N_9858,N_6339,N_7030);
nor U9859 (N_9859,N_6944,N_6428);
nand U9860 (N_9860,N_6559,N_6606);
or U9861 (N_9861,N_6517,N_6514);
or U9862 (N_9862,N_7670,N_7032);
and U9863 (N_9863,N_6266,N_6095);
xor U9864 (N_9864,N_7600,N_6449);
nand U9865 (N_9865,N_6746,N_6455);
nor U9866 (N_9866,N_7626,N_6054);
xnor U9867 (N_9867,N_7051,N_7377);
or U9868 (N_9868,N_6317,N_6494);
or U9869 (N_9869,N_6303,N_7051);
or U9870 (N_9870,N_6856,N_6401);
nor U9871 (N_9871,N_6152,N_6099);
nor U9872 (N_9872,N_6722,N_6728);
or U9873 (N_9873,N_7585,N_6838);
nand U9874 (N_9874,N_6251,N_6818);
nor U9875 (N_9875,N_6699,N_6661);
nor U9876 (N_9876,N_6834,N_7929);
nor U9877 (N_9877,N_6831,N_7936);
and U9878 (N_9878,N_7682,N_7252);
and U9879 (N_9879,N_6055,N_6955);
or U9880 (N_9880,N_6605,N_6655);
or U9881 (N_9881,N_7875,N_7832);
nand U9882 (N_9882,N_7706,N_7243);
nor U9883 (N_9883,N_6092,N_7569);
or U9884 (N_9884,N_7413,N_7644);
xor U9885 (N_9885,N_6932,N_6291);
or U9886 (N_9886,N_6843,N_7772);
nor U9887 (N_9887,N_7825,N_7996);
nand U9888 (N_9888,N_6180,N_6927);
nand U9889 (N_9889,N_6183,N_7913);
and U9890 (N_9890,N_6033,N_6594);
or U9891 (N_9891,N_7567,N_7195);
and U9892 (N_9892,N_7319,N_6685);
or U9893 (N_9893,N_7382,N_6918);
and U9894 (N_9894,N_7956,N_6150);
nand U9895 (N_9895,N_6605,N_6632);
nand U9896 (N_9896,N_7094,N_7600);
and U9897 (N_9897,N_6087,N_6587);
nand U9898 (N_9898,N_6021,N_6274);
nand U9899 (N_9899,N_7865,N_7999);
nor U9900 (N_9900,N_7497,N_6192);
or U9901 (N_9901,N_7188,N_7028);
and U9902 (N_9902,N_6161,N_6261);
nor U9903 (N_9903,N_7588,N_6637);
nor U9904 (N_9904,N_7506,N_6509);
nand U9905 (N_9905,N_7590,N_6487);
or U9906 (N_9906,N_7802,N_6121);
and U9907 (N_9907,N_7257,N_7089);
nor U9908 (N_9908,N_7206,N_6144);
nor U9909 (N_9909,N_7428,N_6494);
nand U9910 (N_9910,N_7002,N_7723);
nand U9911 (N_9911,N_7571,N_6219);
or U9912 (N_9912,N_6882,N_7968);
nor U9913 (N_9913,N_7372,N_6486);
nand U9914 (N_9914,N_6485,N_7415);
and U9915 (N_9915,N_7736,N_6975);
and U9916 (N_9916,N_6148,N_6608);
nor U9917 (N_9917,N_6311,N_6148);
or U9918 (N_9918,N_7390,N_6288);
or U9919 (N_9919,N_7597,N_6704);
or U9920 (N_9920,N_6852,N_7260);
or U9921 (N_9921,N_6288,N_6971);
nand U9922 (N_9922,N_6024,N_7268);
or U9923 (N_9923,N_7246,N_6838);
nor U9924 (N_9924,N_7286,N_6129);
and U9925 (N_9925,N_7168,N_7591);
nand U9926 (N_9926,N_6335,N_7182);
nand U9927 (N_9927,N_7738,N_7356);
and U9928 (N_9928,N_6283,N_7457);
nor U9929 (N_9929,N_7261,N_6342);
nor U9930 (N_9930,N_7292,N_6475);
nand U9931 (N_9931,N_7656,N_7081);
nand U9932 (N_9932,N_6858,N_6146);
or U9933 (N_9933,N_7519,N_6493);
xor U9934 (N_9934,N_7382,N_6584);
and U9935 (N_9935,N_6610,N_7619);
and U9936 (N_9936,N_7304,N_7500);
or U9937 (N_9937,N_6996,N_6159);
or U9938 (N_9938,N_6996,N_7964);
or U9939 (N_9939,N_6817,N_6730);
xnor U9940 (N_9940,N_7708,N_7512);
nor U9941 (N_9941,N_6074,N_7349);
and U9942 (N_9942,N_7858,N_7738);
or U9943 (N_9943,N_7649,N_6681);
nor U9944 (N_9944,N_7847,N_7855);
nand U9945 (N_9945,N_6181,N_6904);
and U9946 (N_9946,N_6437,N_6499);
or U9947 (N_9947,N_6372,N_6609);
nor U9948 (N_9948,N_6226,N_6478);
and U9949 (N_9949,N_6754,N_6847);
and U9950 (N_9950,N_7916,N_7368);
xor U9951 (N_9951,N_6112,N_7837);
or U9952 (N_9952,N_6715,N_6255);
xor U9953 (N_9953,N_7688,N_7018);
nand U9954 (N_9954,N_7866,N_7906);
nor U9955 (N_9955,N_6707,N_7802);
and U9956 (N_9956,N_6874,N_6829);
or U9957 (N_9957,N_7010,N_7778);
or U9958 (N_9958,N_6593,N_7459);
nor U9959 (N_9959,N_7878,N_7401);
nand U9960 (N_9960,N_6034,N_7349);
nand U9961 (N_9961,N_7369,N_6019);
nor U9962 (N_9962,N_6067,N_6511);
nand U9963 (N_9963,N_7018,N_7032);
or U9964 (N_9964,N_6670,N_6335);
nand U9965 (N_9965,N_6780,N_6592);
nor U9966 (N_9966,N_7095,N_6046);
and U9967 (N_9967,N_6647,N_6631);
nor U9968 (N_9968,N_7064,N_7657);
and U9969 (N_9969,N_6045,N_6422);
nand U9970 (N_9970,N_6400,N_7266);
or U9971 (N_9971,N_7901,N_6400);
nor U9972 (N_9972,N_6270,N_6440);
and U9973 (N_9973,N_7781,N_7350);
or U9974 (N_9974,N_7008,N_6431);
and U9975 (N_9975,N_7254,N_6558);
nand U9976 (N_9976,N_6340,N_7840);
nand U9977 (N_9977,N_7562,N_7917);
and U9978 (N_9978,N_6023,N_7189);
and U9979 (N_9979,N_6152,N_6811);
and U9980 (N_9980,N_6621,N_7973);
nand U9981 (N_9981,N_6331,N_6747);
nor U9982 (N_9982,N_6321,N_6699);
nand U9983 (N_9983,N_7058,N_6172);
nor U9984 (N_9984,N_6181,N_6913);
nand U9985 (N_9985,N_6802,N_7634);
nand U9986 (N_9986,N_7467,N_6779);
nand U9987 (N_9987,N_6701,N_6214);
or U9988 (N_9988,N_6938,N_6747);
nand U9989 (N_9989,N_7807,N_7019);
nor U9990 (N_9990,N_6093,N_6510);
nor U9991 (N_9991,N_7102,N_7715);
xnor U9992 (N_9992,N_7007,N_7295);
and U9993 (N_9993,N_6430,N_7382);
and U9994 (N_9994,N_6516,N_7992);
nand U9995 (N_9995,N_6040,N_7136);
or U9996 (N_9996,N_6727,N_7686);
nor U9997 (N_9997,N_7241,N_7621);
xor U9998 (N_9998,N_6112,N_6367);
nand U9999 (N_9999,N_7737,N_7027);
and UO_0 (O_0,N_9934,N_9727);
nand UO_1 (O_1,N_9075,N_9797);
or UO_2 (O_2,N_8161,N_8719);
nor UO_3 (O_3,N_9429,N_8412);
or UO_4 (O_4,N_8417,N_9752);
nand UO_5 (O_5,N_9605,N_8835);
and UO_6 (O_6,N_9718,N_8225);
nand UO_7 (O_7,N_9629,N_9792);
nand UO_8 (O_8,N_8216,N_8771);
nand UO_9 (O_9,N_8142,N_9400);
nor UO_10 (O_10,N_9973,N_9354);
or UO_11 (O_11,N_9307,N_9452);
or UO_12 (O_12,N_8507,N_9288);
nor UO_13 (O_13,N_8777,N_8050);
nand UO_14 (O_14,N_8644,N_8188);
xnor UO_15 (O_15,N_9543,N_9790);
and UO_16 (O_16,N_8569,N_8911);
and UO_17 (O_17,N_9302,N_8479);
and UO_18 (O_18,N_9321,N_9559);
nor UO_19 (O_19,N_9977,N_8187);
nor UO_20 (O_20,N_9177,N_9289);
or UO_21 (O_21,N_8388,N_9395);
nand UO_22 (O_22,N_9172,N_9178);
and UO_23 (O_23,N_9526,N_9217);
and UO_24 (O_24,N_9905,N_9606);
and UO_25 (O_25,N_8859,N_9392);
and UO_26 (O_26,N_8914,N_8334);
or UO_27 (O_27,N_8692,N_9087);
nand UO_28 (O_28,N_8755,N_9781);
nand UO_29 (O_29,N_8100,N_9733);
or UO_30 (O_30,N_9138,N_9428);
nand UO_31 (O_31,N_9917,N_8491);
nor UO_32 (O_32,N_9532,N_8520);
nand UO_33 (O_33,N_8839,N_9823);
nand UO_34 (O_34,N_9184,N_9711);
xnor UO_35 (O_35,N_8582,N_8384);
nor UO_36 (O_36,N_9545,N_8567);
nor UO_37 (O_37,N_8028,N_8634);
nor UO_38 (O_38,N_9084,N_8333);
nor UO_39 (O_39,N_8979,N_9802);
xor UO_40 (O_40,N_9616,N_8966);
xor UO_41 (O_41,N_9788,N_9997);
and UO_42 (O_42,N_8592,N_8872);
nand UO_43 (O_43,N_8353,N_8375);
and UO_44 (O_44,N_8555,N_9607);
nor UO_45 (O_45,N_8217,N_9574);
or UO_46 (O_46,N_8999,N_9534);
xnor UO_47 (O_47,N_9859,N_8181);
nand UO_48 (O_48,N_9393,N_8305);
and UO_49 (O_49,N_9194,N_9709);
nand UO_50 (O_50,N_8513,N_9538);
or UO_51 (O_51,N_8814,N_9215);
nor UO_52 (O_52,N_9432,N_8741);
and UO_53 (O_53,N_8822,N_8763);
nor UO_54 (O_54,N_9502,N_9407);
and UO_55 (O_55,N_8072,N_9698);
and UO_56 (O_56,N_9266,N_9234);
nor UO_57 (O_57,N_9004,N_9482);
xnor UO_58 (O_58,N_9547,N_8599);
nor UO_59 (O_59,N_9907,N_8572);
and UO_60 (O_60,N_8543,N_9332);
nand UO_61 (O_61,N_9098,N_8036);
nand UO_62 (O_62,N_9967,N_9783);
and UO_63 (O_63,N_9147,N_9258);
nand UO_64 (O_64,N_8938,N_9331);
or UO_65 (O_65,N_8199,N_9920);
or UO_66 (O_66,N_9751,N_8259);
nor UO_67 (O_67,N_9628,N_8930);
nor UO_68 (O_68,N_8092,N_9657);
nor UO_69 (O_69,N_9436,N_9986);
nand UO_70 (O_70,N_8194,N_8237);
or UO_71 (O_71,N_9238,N_9621);
or UO_72 (O_72,N_8389,N_8150);
or UO_73 (O_73,N_8166,N_8815);
nor UO_74 (O_74,N_9149,N_8064);
or UO_75 (O_75,N_8271,N_9459);
and UO_76 (O_76,N_9180,N_9068);
or UO_77 (O_77,N_9773,N_9069);
nor UO_78 (O_78,N_9350,N_8667);
nor UO_79 (O_79,N_8831,N_8099);
or UO_80 (O_80,N_9873,N_9142);
nor UO_81 (O_81,N_9578,N_9342);
and UO_82 (O_82,N_8845,N_8364);
nor UO_83 (O_83,N_9897,N_9760);
and UO_84 (O_84,N_8936,N_9155);
and UO_85 (O_85,N_8866,N_8368);
or UO_86 (O_86,N_8971,N_8970);
nor UO_87 (O_87,N_9328,N_8214);
or UO_88 (O_88,N_8029,N_8343);
nor UO_89 (O_89,N_9885,N_9219);
or UO_90 (O_90,N_8516,N_9654);
nand UO_91 (O_91,N_8801,N_9642);
nor UO_92 (O_92,N_9093,N_9467);
nor UO_93 (O_93,N_8697,N_8629);
nor UO_94 (O_94,N_8729,N_8898);
and UO_95 (O_95,N_8608,N_9473);
nor UO_96 (O_96,N_9228,N_8648);
nor UO_97 (O_97,N_8503,N_9937);
and UO_98 (O_98,N_8292,N_9670);
nand UO_99 (O_99,N_9542,N_8945);
and UO_100 (O_100,N_9434,N_8481);
nor UO_101 (O_101,N_9814,N_9813);
nor UO_102 (O_102,N_8880,N_9148);
nor UO_103 (O_103,N_8601,N_8861);
nor UO_104 (O_104,N_9314,N_9213);
and UO_105 (O_105,N_9041,N_8242);
and UO_106 (O_106,N_8458,N_8082);
and UO_107 (O_107,N_9222,N_8110);
and UO_108 (O_108,N_8957,N_8309);
nand UO_109 (O_109,N_8710,N_9015);
nand UO_110 (O_110,N_8427,N_8813);
and UO_111 (O_111,N_8650,N_9281);
nor UO_112 (O_112,N_8612,N_8034);
or UO_113 (O_113,N_9819,N_9540);
or UO_114 (O_114,N_8984,N_8933);
nor UO_115 (O_115,N_9017,N_8120);
nor UO_116 (O_116,N_9655,N_8376);
nor UO_117 (O_117,N_8631,N_8649);
and UO_118 (O_118,N_9283,N_9457);
nand UO_119 (O_119,N_9193,N_8824);
and UO_120 (O_120,N_9984,N_9020);
nand UO_121 (O_121,N_8665,N_9141);
or UO_122 (O_122,N_8836,N_9168);
nand UO_123 (O_123,N_9623,N_9380);
xor UO_124 (O_124,N_8251,N_8734);
or UO_125 (O_125,N_8189,N_9130);
nor UO_126 (O_126,N_9656,N_9679);
nand UO_127 (O_127,N_8020,N_8978);
xor UO_128 (O_128,N_9770,N_8234);
nand UO_129 (O_129,N_9704,N_8675);
nand UO_130 (O_130,N_9622,N_9179);
and UO_131 (O_131,N_9517,N_8672);
xor UO_132 (O_132,N_8043,N_9170);
nand UO_133 (O_133,N_9516,N_9728);
nor UO_134 (O_134,N_8809,N_8439);
nand UO_135 (O_135,N_8553,N_8291);
or UO_136 (O_136,N_9027,N_8358);
nand UO_137 (O_137,N_9563,N_9318);
or UO_138 (O_138,N_8399,N_8992);
nor UO_139 (O_139,N_8195,N_9626);
nand UO_140 (O_140,N_8917,N_8511);
nand UO_141 (O_141,N_8793,N_8867);
or UO_142 (O_142,N_8619,N_8956);
or UO_143 (O_143,N_8006,N_9351);
nor UO_144 (O_144,N_9748,N_9528);
xnor UO_145 (O_145,N_8404,N_8838);
and UO_146 (O_146,N_9593,N_9188);
or UO_147 (O_147,N_8097,N_9385);
nand UO_148 (O_148,N_9793,N_9203);
nor UO_149 (O_149,N_8063,N_8828);
or UO_150 (O_150,N_8937,N_9114);
nor UO_151 (O_151,N_8910,N_8282);
or UO_152 (O_152,N_9465,N_9608);
nand UO_153 (O_153,N_9880,N_9868);
nand UO_154 (O_154,N_8246,N_8972);
nand UO_155 (O_155,N_9946,N_8126);
and UO_156 (O_156,N_9135,N_8136);
nor UO_157 (O_157,N_9049,N_8000);
and UO_158 (O_158,N_9794,N_9836);
or UO_159 (O_159,N_9272,N_8202);
nor UO_160 (O_160,N_9828,N_8762);
and UO_161 (O_161,N_9335,N_9086);
nor UO_162 (O_162,N_9022,N_9001);
and UO_163 (O_163,N_9384,N_9000);
or UO_164 (O_164,N_8642,N_9954);
nand UO_165 (O_165,N_9014,N_9163);
nand UO_166 (O_166,N_8902,N_9466);
and UO_167 (O_167,N_9613,N_8725);
nand UO_168 (O_168,N_8862,N_9031);
nand UO_169 (O_169,N_8780,N_9922);
nand UO_170 (O_170,N_8953,N_9682);
nor UO_171 (O_171,N_9056,N_8379);
and UO_172 (O_172,N_8726,N_9570);
nor UO_173 (O_173,N_8119,N_8366);
or UO_174 (O_174,N_9507,N_8611);
nand UO_175 (O_175,N_9745,N_8244);
nand UO_176 (O_176,N_9693,N_8805);
or UO_177 (O_177,N_9401,N_9769);
nor UO_178 (O_178,N_8269,N_8227);
or UO_179 (O_179,N_8253,N_9415);
nor UO_180 (O_180,N_9514,N_8863);
nand UO_181 (O_181,N_8764,N_9550);
nand UO_182 (O_182,N_8800,N_9107);
nand UO_183 (O_183,N_9681,N_8756);
or UO_184 (O_184,N_9486,N_9129);
and UO_185 (O_185,N_9830,N_9494);
nor UO_186 (O_186,N_8974,N_9064);
or UO_187 (O_187,N_8736,N_8906);
and UO_188 (O_188,N_8329,N_9694);
nor UO_189 (O_189,N_9487,N_9744);
nand UO_190 (O_190,N_8350,N_9377);
nand UO_191 (O_191,N_8791,N_8620);
nand UO_192 (O_192,N_9050,N_9039);
and UO_193 (O_193,N_8745,N_9592);
nand UO_194 (O_194,N_9341,N_8101);
nand UO_195 (O_195,N_9264,N_8913);
or UO_196 (O_196,N_9060,N_9275);
and UO_197 (O_197,N_9619,N_9376);
nand UO_198 (O_198,N_8009,N_9110);
or UO_199 (O_199,N_8703,N_8127);
and UO_200 (O_200,N_8066,N_9749);
nand UO_201 (O_201,N_9750,N_8302);
or UO_202 (O_202,N_8407,N_8812);
nor UO_203 (O_203,N_8206,N_9826);
or UO_204 (O_204,N_9011,N_8735);
or UO_205 (O_205,N_8664,N_8348);
nand UO_206 (O_206,N_8738,N_8335);
and UO_207 (O_207,N_8431,N_9105);
or UO_208 (O_208,N_9667,N_8157);
or UO_209 (O_209,N_9865,N_8449);
and UO_210 (O_210,N_9715,N_8109);
and UO_211 (O_211,N_8873,N_9097);
nor UO_212 (O_212,N_8044,N_8443);
xor UO_213 (O_213,N_9462,N_8095);
or UO_214 (O_214,N_9333,N_9892);
nor UO_215 (O_215,N_8156,N_8495);
or UO_216 (O_216,N_8709,N_9697);
nand UO_217 (O_217,N_9556,N_9730);
or UO_218 (O_218,N_9689,N_8517);
or UO_219 (O_219,N_9779,N_8639);
and UO_220 (O_220,N_8073,N_9356);
nor UO_221 (O_221,N_9208,N_9504);
nand UO_222 (O_222,N_8032,N_9383);
nand UO_223 (O_223,N_9630,N_8848);
nand UO_224 (O_224,N_8480,N_9856);
nor UO_225 (O_225,N_8975,N_9471);
nand UO_226 (O_226,N_8580,N_9403);
xnor UO_227 (O_227,N_9840,N_8689);
nor UO_228 (O_228,N_8576,N_8461);
or UO_229 (O_229,N_8472,N_8182);
and UO_230 (O_230,N_9460,N_9546);
nand UO_231 (O_231,N_8145,N_9051);
nor UO_232 (O_232,N_9363,N_9386);
nor UO_233 (O_233,N_8258,N_8625);
nand UO_234 (O_234,N_9025,N_8395);
and UO_235 (O_235,N_9210,N_9349);
or UO_236 (O_236,N_8342,N_9690);
nand UO_237 (O_237,N_8964,N_8071);
nand UO_238 (O_238,N_8121,N_8519);
nor UO_239 (O_239,N_9080,N_8566);
nor UO_240 (O_240,N_9006,N_9162);
or UO_241 (O_241,N_8765,N_9270);
or UO_242 (O_242,N_9531,N_9405);
or UO_243 (O_243,N_8323,N_8113);
xor UO_244 (O_244,N_8135,N_9417);
xnor UO_245 (O_245,N_8578,N_8536);
nor UO_246 (O_246,N_8018,N_8179);
or UO_247 (O_247,N_9544,N_8514);
or UO_248 (O_248,N_8371,N_9777);
and UO_249 (O_249,N_8792,N_8786);
or UO_250 (O_250,N_9820,N_9942);
or UO_251 (O_251,N_9662,N_9348);
and UO_252 (O_252,N_8160,N_8465);
or UO_253 (O_253,N_8941,N_8604);
nand UO_254 (O_254,N_8463,N_8767);
nor UO_255 (O_255,N_8737,N_8635);
nand UO_256 (O_256,N_9186,N_8818);
nor UO_257 (O_257,N_9933,N_9477);
or UO_258 (O_258,N_9449,N_9646);
nand UO_259 (O_259,N_8939,N_9975);
nor UO_260 (O_260,N_9833,N_9644);
or UO_261 (O_261,N_8124,N_8833);
or UO_262 (O_262,N_8727,N_8823);
and UO_263 (O_263,N_9480,N_8233);
and UO_264 (O_264,N_9995,N_8946);
or UO_265 (O_265,N_9716,N_9190);
or UO_266 (O_266,N_9604,N_9311);
and UO_267 (O_267,N_8056,N_9438);
and UO_268 (O_268,N_8162,N_8143);
nor UO_269 (O_269,N_9719,N_8285);
and UO_270 (O_270,N_9095,N_8279);
nor UO_271 (O_271,N_9879,N_8674);
xor UO_272 (O_272,N_8477,N_9557);
or UO_273 (O_273,N_9869,N_8958);
and UO_274 (O_274,N_8130,N_8210);
nand UO_275 (O_275,N_9468,N_8355);
and UO_276 (O_276,N_8215,N_8441);
and UO_277 (O_277,N_8406,N_8455);
or UO_278 (O_278,N_8111,N_9941);
or UO_279 (O_279,N_8435,N_8026);
and UO_280 (O_280,N_9059,N_9675);
nor UO_281 (O_281,N_8988,N_8893);
or UO_282 (O_282,N_8122,N_9280);
nor UO_283 (O_283,N_9003,N_9916);
and UO_284 (O_284,N_9308,N_9082);
nor UO_285 (O_285,N_9855,N_8666);
and UO_286 (O_286,N_8001,N_9888);
and UO_287 (O_287,N_8462,N_9843);
and UO_288 (O_288,N_8386,N_9365);
and UO_289 (O_289,N_8784,N_9512);
and UO_290 (O_290,N_9085,N_9309);
or UO_291 (O_291,N_9611,N_9652);
nor UO_292 (O_292,N_8591,N_8451);
xnor UO_293 (O_293,N_9033,N_9548);
or UO_294 (O_294,N_8897,N_8192);
and UO_295 (O_295,N_9767,N_8915);
nor UO_296 (O_296,N_8139,N_8277);
nand UO_297 (O_297,N_9490,N_8087);
and UO_298 (O_298,N_9418,N_9419);
nor UO_299 (O_299,N_8250,N_8345);
and UO_300 (O_300,N_8023,N_8947);
nand UO_301 (O_301,N_8422,N_8991);
xnor UO_302 (O_302,N_9404,N_9045);
nor UO_303 (O_303,N_8304,N_9965);
and UO_304 (O_304,N_9424,N_9566);
or UO_305 (O_305,N_8594,N_9343);
nand UO_306 (O_306,N_9982,N_8661);
nand UO_307 (O_307,N_8381,N_8058);
or UO_308 (O_308,N_8403,N_8884);
or UO_309 (O_309,N_9765,N_8372);
and UO_310 (O_310,N_9591,N_8038);
nand UO_311 (O_311,N_8331,N_9878);
and UO_312 (O_312,N_9273,N_8270);
and UO_313 (O_313,N_8545,N_8228);
nor UO_314 (O_314,N_8724,N_8096);
and UO_315 (O_315,N_8560,N_8008);
nand UO_316 (O_316,N_9699,N_8769);
nand UO_317 (O_317,N_9073,N_9245);
and UO_318 (O_318,N_8327,N_9124);
or UO_319 (O_319,N_9653,N_9599);
and UO_320 (O_320,N_9988,N_9672);
or UO_321 (O_321,N_8021,N_8452);
nor UO_322 (O_322,N_8506,N_9587);
and UO_323 (O_323,N_8132,N_8577);
and UO_324 (O_324,N_9316,N_9235);
or UO_325 (O_325,N_8821,N_9506);
nor UO_326 (O_326,N_8478,N_9702);
nor UO_327 (O_327,N_8600,N_9346);
nor UO_328 (O_328,N_8040,N_8858);
nand UO_329 (O_329,N_9464,N_8949);
or UO_330 (O_330,N_8437,N_8289);
or UO_331 (O_331,N_9996,N_8610);
or UO_332 (O_332,N_9650,N_9347);
nor UO_333 (O_333,N_8400,N_8523);
and UO_334 (O_334,N_9918,N_9530);
and UO_335 (O_335,N_8052,N_8987);
and UO_336 (O_336,N_9382,N_8349);
or UO_337 (O_337,N_9005,N_8829);
or UO_338 (O_338,N_8450,N_9929);
and UO_339 (O_339,N_8854,N_9212);
xor UO_340 (O_340,N_8810,N_8249);
nand UO_341 (O_341,N_9772,N_8537);
and UO_342 (O_342,N_9796,N_9478);
and UO_343 (O_343,N_9101,N_8453);
and UO_344 (O_344,N_8899,N_8985);
or UO_345 (O_345,N_8061,N_8380);
or UO_346 (O_346,N_9241,N_9860);
nand UO_347 (O_347,N_8834,N_8267);
or UO_348 (O_348,N_9047,N_9396);
or UO_349 (O_349,N_8301,N_9666);
nand UO_350 (O_350,N_9362,N_8943);
or UO_351 (O_351,N_9372,N_8447);
and UO_352 (O_352,N_8876,N_9572);
nor UO_353 (O_353,N_9055,N_8474);
or UO_354 (O_354,N_8901,N_8434);
nor UO_355 (O_355,N_9755,N_8394);
and UO_356 (O_356,N_9100,N_8844);
or UO_357 (O_357,N_9236,N_8895);
nor UO_358 (O_358,N_9040,N_8993);
and UO_359 (O_359,N_8330,N_8896);
or UO_360 (O_360,N_9771,N_9071);
nor UO_361 (O_361,N_8847,N_8405);
or UO_362 (O_362,N_8654,N_8257);
nand UO_363 (O_363,N_9024,N_9503);
or UO_364 (O_364,N_9867,N_9758);
nand UO_365 (O_365,N_8245,N_8207);
nor UO_366 (O_366,N_8299,N_8921);
nand UO_367 (O_367,N_8235,N_8656);
and UO_368 (O_368,N_9639,N_8616);
xnor UO_369 (O_369,N_8418,N_8676);
and UO_370 (O_370,N_8796,N_8870);
nor UO_371 (O_371,N_8841,N_8278);
and UO_372 (O_372,N_8565,N_8391);
nand UO_373 (O_373,N_8721,N_9881);
and UO_374 (O_374,N_9090,N_9782);
and UO_375 (O_375,N_8759,N_9551);
nand UO_376 (O_376,N_8193,N_9565);
nor UO_377 (O_377,N_8500,N_9156);
xnor UO_378 (O_378,N_8761,N_8432);
nand UO_379 (O_379,N_8347,N_9176);
or UO_380 (O_380,N_8067,N_9315);
nand UO_381 (O_381,N_9994,N_8722);
or UO_382 (O_382,N_9999,N_8626);
and UO_383 (O_383,N_8996,N_9932);
nor UO_384 (O_384,N_8169,N_8003);
or UO_385 (O_385,N_9450,N_9609);
nand UO_386 (O_386,N_9858,N_9617);
xnor UO_387 (O_387,N_8842,N_9541);
and UO_388 (O_388,N_9576,N_8211);
nor UO_389 (O_389,N_9577,N_9019);
nor UO_390 (O_390,N_8630,N_9474);
nor UO_391 (O_391,N_8534,N_9943);
nor UO_392 (O_392,N_8178,N_8923);
nor UO_393 (O_393,N_8027,N_9271);
or UO_394 (O_394,N_9077,N_8012);
nor UO_395 (O_395,N_9352,N_8484);
and UO_396 (O_396,N_9221,N_8025);
and UO_397 (O_397,N_9255,N_9846);
nor UO_398 (O_398,N_8397,N_9035);
nand UO_399 (O_399,N_8374,N_9936);
nor UO_400 (O_400,N_9002,N_8387);
nand UO_401 (O_401,N_8326,N_8098);
and UO_402 (O_402,N_9322,N_9935);
nand UO_403 (O_403,N_9589,N_8473);
nand UO_404 (O_404,N_9807,N_9475);
nor UO_405 (O_405,N_9276,N_9567);
or UO_406 (O_406,N_9371,N_9723);
nor UO_407 (O_407,N_8321,N_9201);
nand UO_408 (O_408,N_8995,N_9286);
or UO_409 (O_409,N_9731,N_9710);
nand UO_410 (O_410,N_9537,N_9625);
nand UO_411 (O_411,N_8310,N_9809);
xnor UO_412 (O_412,N_9079,N_9323);
or UO_413 (O_413,N_8502,N_8529);
or UO_414 (O_414,N_8541,N_9787);
nor UO_415 (O_415,N_9143,N_8524);
nand UO_416 (O_416,N_8637,N_9575);
and UO_417 (O_417,N_8693,N_8205);
nor UO_418 (O_418,N_8579,N_9924);
or UO_419 (O_419,N_8934,N_8927);
nor UO_420 (O_420,N_9960,N_9296);
and UO_421 (O_421,N_9013,N_9146);
nor UO_422 (O_422,N_8615,N_9944);
nand UO_423 (O_423,N_8392,N_9725);
nor UO_424 (O_424,N_8652,N_9306);
nand UO_425 (O_425,N_9360,N_9956);
nand UO_426 (O_426,N_9303,N_8521);
nor UO_427 (O_427,N_8284,N_8039);
or UO_428 (O_428,N_8222,N_8681);
nand UO_429 (O_429,N_8487,N_9324);
nand UO_430 (O_430,N_9757,N_9612);
nand UO_431 (O_431,N_8877,N_8468);
or UO_432 (O_432,N_9866,N_9786);
or UO_433 (O_433,N_9601,N_8772);
nand UO_434 (O_434,N_8622,N_9265);
xnor UO_435 (O_435,N_8236,N_8307);
nor UO_436 (O_436,N_8527,N_9010);
nor UO_437 (O_437,N_9983,N_8445);
and UO_438 (O_438,N_9552,N_8886);
nor UO_439 (O_439,N_9908,N_8885);
or UO_440 (O_440,N_8114,N_8636);
and UO_441 (O_441,N_9214,N_8268);
or UO_442 (O_442,N_9870,N_9927);
nor UO_443 (O_443,N_8010,N_9992);
or UO_444 (O_444,N_8981,N_9596);
nor UO_445 (O_445,N_8808,N_9078);
nor UO_446 (O_446,N_9738,N_8717);
xnor UO_447 (O_447,N_8940,N_8874);
nor UO_448 (O_448,N_9046,N_8501);
and UO_449 (O_449,N_8294,N_8146);
and UO_450 (O_450,N_8557,N_9980);
and UO_451 (O_451,N_8887,N_8951);
nand UO_452 (O_452,N_8846,N_9513);
or UO_453 (O_453,N_9412,N_9906);
or UO_454 (O_454,N_8782,N_8151);
nor UO_455 (O_455,N_8853,N_9966);
nor UO_456 (O_456,N_9640,N_9445);
nand UO_457 (O_457,N_9741,N_9268);
and UO_458 (O_458,N_8425,N_9799);
nand UO_459 (O_459,N_8632,N_9237);
nor UO_460 (O_460,N_8508,N_8617);
and UO_461 (O_461,N_8558,N_9030);
or UO_462 (O_462,N_9220,N_8730);
nand UO_463 (O_463,N_8024,N_9803);
and UO_464 (O_464,N_9126,N_8746);
or UO_465 (O_465,N_9028,N_9632);
and UO_466 (O_466,N_8252,N_8276);
and UO_467 (O_467,N_8633,N_9614);
or UO_468 (O_468,N_9753,N_8223);
nand UO_469 (O_469,N_9312,N_9903);
and UO_470 (O_470,N_8679,N_9940);
nor UO_471 (O_471,N_9397,N_8483);
nor UO_472 (O_472,N_9740,N_9125);
nand UO_473 (O_473,N_8699,N_9915);
nor UO_474 (O_474,N_8533,N_9167);
nand UO_475 (O_475,N_9416,N_8286);
and UO_476 (O_476,N_8022,N_9427);
or UO_477 (O_477,N_9610,N_9962);
and UO_478 (O_478,N_8104,N_9092);
and UO_479 (O_479,N_8288,N_8783);
nor UO_480 (O_480,N_8457,N_8315);
nand UO_481 (O_481,N_8948,N_8275);
and UO_482 (O_482,N_8147,N_9884);
nand UO_483 (O_483,N_8125,N_8655);
and UO_484 (O_484,N_9326,N_9109);
nor UO_485 (O_485,N_8590,N_9195);
nand UO_486 (O_486,N_9132,N_9206);
nor UO_487 (O_487,N_9676,N_9847);
nand UO_488 (O_488,N_8776,N_9463);
or UO_489 (O_489,N_9810,N_8817);
and UO_490 (O_490,N_9827,N_8377);
and UO_491 (O_491,N_9595,N_9677);
or UO_492 (O_492,N_8538,N_9585);
or UO_493 (O_493,N_8997,N_9103);
and UO_494 (O_494,N_8811,N_8747);
and UO_495 (O_495,N_9579,N_8239);
xor UO_496 (O_496,N_8266,N_8200);
or UO_497 (O_497,N_9390,N_9104);
nand UO_498 (O_498,N_8748,N_9600);
or UO_499 (O_499,N_9964,N_9998);
or UO_500 (O_500,N_9345,N_8401);
and UO_501 (O_501,N_9862,N_9317);
nand UO_502 (O_502,N_8751,N_8370);
nor UO_503 (O_503,N_9497,N_9701);
nor UO_504 (O_504,N_9991,N_8002);
nor UO_505 (O_505,N_9204,N_9052);
nand UO_506 (O_506,N_8303,N_8967);
nand UO_507 (O_507,N_8882,N_9951);
or UO_508 (O_508,N_8197,N_8928);
nand UO_509 (O_509,N_9008,N_9774);
nor UO_510 (O_510,N_8879,N_9375);
and UO_511 (O_511,N_8894,N_9558);
or UO_512 (O_512,N_8059,N_8712);
and UO_513 (O_513,N_8528,N_9737);
or UO_514 (O_514,N_8108,N_8961);
or UO_515 (O_515,N_8154,N_8701);
and UO_516 (O_516,N_9889,N_8019);
and UO_517 (O_517,N_8409,N_9455);
nand UO_518 (O_518,N_9373,N_9123);
nor UO_519 (O_519,N_9958,N_9634);
or UO_520 (O_520,N_8778,N_9131);
and UO_521 (O_521,N_9108,N_9357);
nor UO_522 (O_522,N_8281,N_9152);
and UO_523 (O_523,N_9259,N_8141);
xnor UO_524 (O_524,N_9358,N_8180);
or UO_525 (O_525,N_8184,N_9066);
nand UO_526 (O_526,N_9310,N_9928);
or UO_527 (O_527,N_9925,N_9597);
nand UO_528 (O_528,N_9638,N_9230);
nor UO_529 (O_529,N_9726,N_8696);
or UO_530 (O_530,N_9454,N_9290);
nor UO_531 (O_531,N_8924,N_9279);
nand UO_532 (O_532,N_8094,N_9300);
nor UO_533 (O_533,N_8708,N_9674);
nand UO_534 (O_534,N_9153,N_8360);
and UO_535 (O_535,N_9239,N_9853);
or UO_536 (O_536,N_8265,N_9325);
and UO_537 (O_537,N_8865,N_9705);
nand UO_538 (O_538,N_9624,N_9972);
nand UO_539 (O_539,N_9067,N_8905);
or UO_540 (O_540,N_9501,N_8891);
nand UO_541 (O_541,N_9057,N_9987);
or UO_542 (O_542,N_9872,N_8243);
nor UO_543 (O_543,N_8153,N_8504);
nor UO_544 (O_544,N_9007,N_8486);
xor UO_545 (O_545,N_8005,N_9479);
and UO_546 (O_546,N_8883,N_8651);
or UO_547 (O_547,N_8830,N_8732);
nor UO_548 (O_548,N_8089,N_9065);
nand UO_549 (O_549,N_8317,N_9089);
or UO_550 (O_550,N_8552,N_9437);
nor UO_551 (O_551,N_9446,N_9631);
and UO_552 (O_552,N_9949,N_9660);
and UO_553 (O_553,N_9329,N_9742);
nor UO_554 (O_554,N_8584,N_8356);
nand UO_555 (O_555,N_8641,N_8410);
nor UO_556 (O_556,N_9811,N_8671);
nor UO_557 (O_557,N_9298,N_8718);
and UO_558 (O_558,N_9253,N_9293);
xor UO_559 (O_559,N_8081,N_9535);
and UO_560 (O_560,N_8843,N_9931);
nor UO_561 (O_561,N_8624,N_8138);
nor UO_562 (O_562,N_9144,N_8720);
nor UO_563 (O_563,N_9026,N_8918);
or UO_564 (O_564,N_9036,N_8573);
nand UO_565 (O_565,N_8702,N_8170);
xnor UO_566 (O_566,N_9732,N_9252);
nor UO_567 (O_567,N_8658,N_9590);
nor UO_568 (O_568,N_9784,N_8361);
nor UO_569 (O_569,N_8176,N_9914);
and UO_570 (O_570,N_8442,N_9527);
nand UO_571 (O_571,N_8920,N_8768);
and UO_572 (O_572,N_8952,N_9118);
and UO_573 (O_573,N_9893,N_8855);
nor UO_574 (O_574,N_9883,N_8128);
xnor UO_575 (O_575,N_8396,N_8295);
nand UO_576 (O_576,N_9500,N_9083);
or UO_577 (O_577,N_8165,N_8976);
nand UO_578 (O_578,N_9173,N_8739);
nand UO_579 (O_579,N_9284,N_9489);
nor UO_580 (O_580,N_8428,N_8436);
or UO_581 (O_581,N_9425,N_9854);
and UO_582 (O_582,N_9508,N_8173);
and UO_583 (O_583,N_9175,N_8522);
or UO_584 (O_584,N_8300,N_9336);
or UO_585 (O_585,N_9254,N_8587);
or UO_586 (O_586,N_8378,N_8998);
nand UO_587 (O_587,N_8959,N_9824);
nor UO_588 (O_588,N_9313,N_9091);
and UO_589 (O_589,N_8030,N_9399);
nand UO_590 (O_590,N_8123,N_9549);
or UO_591 (O_591,N_9044,N_8969);
nand UO_592 (O_592,N_8469,N_9244);
and UO_593 (O_593,N_8414,N_9402);
or UO_594 (O_594,N_9260,N_8088);
or UO_595 (O_595,N_9721,N_9422);
nor UO_596 (O_596,N_9297,N_9829);
or UO_597 (O_597,N_8682,N_9451);
or UO_598 (O_598,N_8670,N_9301);
and UO_599 (O_599,N_8657,N_9122);
nand UO_600 (O_600,N_9665,N_9910);
nand UO_601 (O_601,N_8586,N_8174);
or UO_602 (O_602,N_8628,N_9554);
and UO_603 (O_603,N_9678,N_9900);
nor UO_604 (O_604,N_9911,N_9106);
and UO_605 (O_605,N_8583,N_8488);
or UO_606 (O_606,N_9661,N_8677);
and UO_607 (O_607,N_8512,N_9871);
or UO_608 (O_608,N_8103,N_9361);
nor UO_609 (O_609,N_9816,N_9778);
nand UO_610 (O_610,N_8663,N_9158);
nand UO_611 (O_611,N_8685,N_8416);
nor UO_612 (O_612,N_8875,N_8048);
nor UO_613 (O_613,N_9240,N_9978);
and UO_614 (O_614,N_8925,N_9334);
nand UO_615 (O_615,N_9834,N_9320);
nand UO_616 (O_616,N_8163,N_8322);
and UO_617 (O_617,N_8041,N_8175);
nand UO_618 (O_618,N_9561,N_9447);
and UO_619 (O_619,N_9248,N_8224);
nand UO_620 (O_620,N_8869,N_8888);
nand UO_621 (O_621,N_8332,N_8904);
nor UO_622 (O_622,N_8646,N_8264);
or UO_623 (O_623,N_9722,N_9115);
nand UO_624 (O_624,N_8691,N_8788);
or UO_625 (O_625,N_8298,N_8444);
nor UO_626 (O_626,N_8602,N_8492);
xnor UO_627 (O_627,N_8185,N_9707);
and UO_628 (O_628,N_8944,N_9564);
nand UO_629 (O_629,N_9406,N_9112);
nor UO_630 (O_630,N_9229,N_8464);
and UO_631 (O_631,N_9430,N_8398);
nor UO_632 (O_632,N_8466,N_9651);
nor UO_633 (O_633,N_8743,N_8070);
or UO_634 (O_634,N_8562,N_8482);
or UO_635 (O_635,N_9948,N_9505);
nand UO_636 (O_636,N_8962,N_8563);
nand UO_637 (O_637,N_8903,N_9861);
or UO_638 (O_638,N_9562,N_9246);
or UO_639 (O_639,N_9495,N_8868);
and UO_640 (O_640,N_9825,N_8989);
and UO_641 (O_641,N_8352,N_9038);
and UO_642 (O_642,N_9603,N_8864);
and UO_643 (O_643,N_9615,N_8973);
or UO_644 (O_644,N_9898,N_9775);
and UO_645 (O_645,N_8881,N_8475);
or UO_646 (O_646,N_8744,N_8561);
nand UO_647 (O_647,N_8158,N_9410);
nand UO_648 (O_648,N_8660,N_9818);
or UO_649 (O_649,N_8208,N_9043);
and UO_650 (O_650,N_9340,N_8339);
and UO_651 (O_651,N_8546,N_8890);
and UO_652 (O_652,N_8686,N_8787);
nand UO_653 (O_653,N_8826,N_8051);
nand UO_654 (O_654,N_8490,N_9521);
or UO_655 (O_655,N_8262,N_8004);
or UO_656 (O_656,N_8499,N_9062);
and UO_657 (O_657,N_9832,N_9481);
and UO_658 (O_658,N_8438,N_8550);
or UO_659 (O_659,N_8338,N_8505);
nor UO_660 (O_660,N_8714,N_9048);
nor UO_661 (O_661,N_9461,N_8336);
and UO_662 (O_662,N_8232,N_8367);
nand UO_663 (O_663,N_8860,N_8673);
or UO_664 (O_664,N_8155,N_9863);
nand UO_665 (O_665,N_9939,N_9021);
nor UO_666 (O_666,N_8700,N_8668);
nor UO_667 (O_667,N_8935,N_9319);
or UO_668 (O_668,N_9768,N_8609);
xnor UO_669 (O_669,N_8454,N_8554);
nand UO_670 (O_670,N_8017,N_9938);
nand UO_671 (O_671,N_9469,N_8926);
and UO_672 (O_672,N_8293,N_8083);
or UO_673 (O_673,N_8530,N_9837);
and UO_674 (O_674,N_9113,N_9166);
and UO_675 (O_675,N_9411,N_9806);
or UO_676 (O_676,N_8698,N_9766);
nand UO_677 (O_677,N_8013,N_9519);
nand UO_678 (O_678,N_8856,N_9160);
nand UO_679 (O_679,N_9979,N_9216);
nor UO_680 (O_680,N_9374,N_8102);
or UO_681 (O_681,N_9523,N_9930);
and UO_682 (O_682,N_9974,N_9174);
or UO_683 (O_683,N_9720,N_8694);
or UO_684 (O_684,N_9029,N_9842);
nand UO_685 (O_685,N_9525,N_8383);
nand UO_686 (O_686,N_8990,N_9472);
nand UO_687 (O_687,N_8871,N_8711);
or UO_688 (O_688,N_9121,N_9838);
and UO_689 (O_689,N_8105,N_9736);
xnor UO_690 (O_690,N_8852,N_8752);
or UO_691 (O_691,N_9181,N_9339);
or UO_692 (O_692,N_8758,N_9586);
nor UO_693 (O_693,N_9952,N_8750);
or UO_694 (O_694,N_9522,N_8645);
and UO_695 (O_695,N_9685,N_8042);
and UO_696 (O_696,N_8713,N_8016);
nand UO_697 (O_697,N_9762,N_9553);
nand UO_698 (O_698,N_8426,N_8593);
and UO_699 (O_699,N_8797,N_9588);
or UO_700 (O_700,N_9636,N_8518);
nand UO_701 (O_701,N_8749,N_9243);
nand UO_702 (O_702,N_9493,N_9439);
nand UO_703 (O_703,N_9267,N_9696);
and UO_704 (O_704,N_8683,N_9224);
xor UO_705 (O_705,N_9759,N_9673);
and UO_706 (O_706,N_9691,N_8263);
nand UO_707 (O_707,N_8074,N_9583);
and UO_708 (O_708,N_8055,N_9128);
or UO_709 (O_709,N_8117,N_9582);
nand UO_710 (O_710,N_9695,N_9291);
nand UO_711 (O_711,N_8621,N_8240);
nor UO_712 (O_712,N_8084,N_8695);
and UO_713 (O_713,N_8733,N_8798);
and UO_714 (O_714,N_9161,N_8900);
and UO_715 (O_715,N_9692,N_8757);
nand UO_716 (O_716,N_9886,N_8148);
or UO_717 (O_717,N_9641,N_8290);
and UO_718 (O_718,N_8647,N_8241);
or UO_719 (O_719,N_8093,N_9687);
nor UO_720 (O_720,N_8680,N_8247);
nand UO_721 (O_721,N_8539,N_8402);
nand UO_722 (O_722,N_8047,N_8011);
nor UO_723 (O_723,N_8053,N_8045);
or UO_724 (O_724,N_9637,N_9812);
xor UO_725 (O_725,N_8955,N_9111);
or UO_726 (O_726,N_8606,N_8167);
and UO_727 (O_727,N_9839,N_8287);
nor UO_728 (O_728,N_8152,N_9841);
nor UO_729 (O_729,N_9042,N_9849);
or UO_730 (O_730,N_9227,N_8614);
and UO_731 (O_731,N_9199,N_9072);
nand UO_732 (O_732,N_9815,N_9169);
nor UO_733 (O_733,N_9441,N_8218);
nand UO_734 (O_734,N_9198,N_8035);
nor UO_735 (O_735,N_8819,N_8889);
nand UO_736 (O_736,N_9269,N_9278);
nand UO_737 (O_737,N_9485,N_9891);
nand UO_738 (O_738,N_9684,N_9945);
or UO_739 (O_739,N_9164,N_8433);
or UO_740 (O_740,N_8684,N_9539);
or UO_741 (O_741,N_9102,N_8408);
nand UO_742 (O_742,N_9223,N_9119);
nand UO_743 (O_743,N_8986,N_9518);
nand UO_744 (O_744,N_9458,N_8548);
nor UO_745 (O_745,N_9780,N_9985);
and UO_746 (O_746,N_8470,N_8046);
or UO_747 (O_747,N_8781,N_8107);
or UO_748 (O_748,N_8688,N_8607);
or UO_749 (O_749,N_8931,N_8742);
and UO_750 (O_750,N_9285,N_9294);
nor UO_751 (O_751,N_9568,N_8133);
or UO_752 (O_752,N_8049,N_9099);
or UO_753 (O_753,N_8807,N_8618);
nor UO_754 (O_754,N_9848,N_9963);
nand UO_755 (O_755,N_9492,N_8707);
nand UO_756 (O_756,N_8706,N_8705);
nor UO_757 (O_757,N_9569,N_9327);
and UO_758 (O_758,N_9421,N_8213);
and UO_759 (O_759,N_8344,N_9524);
or UO_760 (O_760,N_9499,N_9909);
and UO_761 (O_761,N_8570,N_9231);
nor UO_762 (O_762,N_9754,N_9391);
and UO_763 (O_763,N_9249,N_9904);
nand UO_764 (O_764,N_8851,N_8559);
nand UO_765 (O_765,N_9763,N_9151);
nand UO_766 (O_766,N_9488,N_9094);
nor UO_767 (O_767,N_8785,N_9032);
and UO_768 (O_768,N_9686,N_8510);
or UO_769 (O_769,N_8892,N_8489);
and UO_770 (O_770,N_9185,N_8597);
nor UO_771 (O_771,N_9145,N_8254);
or UO_772 (O_772,N_8581,N_9137);
nand UO_773 (O_773,N_9511,N_9895);
and UO_774 (O_774,N_9808,N_9061);
and UO_775 (O_775,N_9584,N_9453);
and UO_776 (O_776,N_8308,N_9875);
and UO_777 (O_777,N_8341,N_9706);
nand UO_778 (O_778,N_9232,N_8068);
and UO_779 (O_779,N_9668,N_8078);
and UO_780 (O_780,N_9633,N_9157);
xnor UO_781 (O_781,N_8283,N_8850);
and UO_782 (O_782,N_8037,N_9703);
or UO_783 (O_783,N_8916,N_8728);
xor UO_784 (O_784,N_8613,N_9159);
and UO_785 (O_785,N_8415,N_9664);
nand UO_786 (O_786,N_9627,N_8354);
nor UO_787 (O_787,N_8090,N_8789);
nand UO_788 (O_788,N_9287,N_9444);
xnor UO_789 (O_789,N_9096,N_8932);
nand UO_790 (O_790,N_9054,N_8226);
or UO_791 (O_791,N_9009,N_8968);
or UO_792 (O_792,N_9913,N_8775);
nand UO_793 (O_793,N_8159,N_9483);
nor UO_794 (O_794,N_9533,N_8598);
nand UO_795 (O_795,N_9620,N_9926);
or UO_796 (O_796,N_8365,N_8238);
nor UO_797 (O_797,N_8219,N_8754);
or UO_798 (O_798,N_9209,N_9389);
nand UO_799 (O_799,N_9366,N_8779);
nor UO_800 (O_800,N_8575,N_8908);
and UO_801 (O_801,N_9990,N_8069);
nand UO_802 (O_802,N_9355,N_8203);
nor UO_803 (O_803,N_8351,N_9700);
nor UO_804 (O_804,N_8509,N_8640);
or UO_805 (O_805,N_9894,N_8313);
and UO_806 (O_806,N_9344,N_8273);
and UO_807 (O_807,N_8085,N_8007);
nand UO_808 (O_808,N_9127,N_9016);
nor UO_809 (O_809,N_8542,N_8060);
nor UO_810 (O_810,N_8363,N_8115);
nor UO_811 (O_811,N_9225,N_8186);
nor UO_812 (O_812,N_9955,N_9023);
nor UO_813 (O_813,N_9801,N_9256);
nand UO_814 (O_814,N_9414,N_8296);
nor UO_815 (O_815,N_8773,N_9764);
nand UO_816 (O_816,N_9182,N_8086);
and UO_817 (O_817,N_9845,N_9969);
or UO_818 (O_818,N_9018,N_9262);
and UO_819 (O_819,N_8311,N_9852);
or UO_820 (O_820,N_9981,N_8596);
and UO_821 (O_821,N_8171,N_8909);
or UO_822 (O_822,N_9817,N_9735);
and UO_823 (O_823,N_8802,N_9165);
and UO_824 (O_824,N_9408,N_9902);
and UO_825 (O_825,N_8716,N_8079);
and UO_826 (O_826,N_9140,N_8603);
or UO_827 (O_827,N_8362,N_8907);
or UO_828 (O_828,N_8816,N_8460);
nor UO_829 (O_829,N_8054,N_8731);
nor UO_830 (O_830,N_8390,N_8129);
nand UO_831 (O_831,N_8033,N_9671);
and UO_832 (O_832,N_9805,N_8140);
nand UO_833 (O_833,N_9598,N_9420);
nor UO_834 (O_834,N_8994,N_9795);
and UO_835 (O_835,N_9835,N_8977);
nor UO_836 (O_836,N_8574,N_8498);
nand UO_837 (O_837,N_9034,N_8168);
nand UO_838 (O_838,N_9789,N_9251);
xnor UO_839 (O_839,N_8525,N_9635);
or UO_840 (O_840,N_8929,N_8799);
and UO_841 (O_841,N_9058,N_9257);
nand UO_842 (O_842,N_9299,N_8261);
and UO_843 (O_843,N_8827,N_8316);
and UO_844 (O_844,N_8723,N_9717);
and UO_845 (O_845,N_8320,N_9890);
nand UO_846 (O_846,N_8448,N_9196);
nand UO_847 (O_847,N_9435,N_8515);
nand UO_848 (O_848,N_8965,N_8031);
nand UO_849 (O_849,N_8467,N_8653);
nor UO_850 (O_850,N_9989,N_8420);
or UO_851 (O_851,N_8172,N_8134);
and UO_852 (O_852,N_8221,N_8411);
or UO_853 (O_853,N_9761,N_8878);
nand UO_854 (O_854,N_8456,N_9171);
and UO_855 (O_855,N_9498,N_8091);
and UO_856 (O_856,N_8669,N_8678);
and UO_857 (O_857,N_8106,N_9187);
nand UO_858 (O_858,N_8198,N_9571);
or UO_859 (O_859,N_8190,N_8191);
and UO_860 (O_860,N_9116,N_9857);
nor UO_861 (O_861,N_8919,N_9851);
nand UO_862 (O_862,N_8740,N_9456);
or UO_863 (O_863,N_8328,N_8623);
nor UO_864 (O_864,N_9442,N_9822);
nand UO_865 (O_865,N_8766,N_8212);
nand UO_866 (O_866,N_8280,N_9282);
nand UO_867 (O_867,N_8346,N_8704);
nor UO_868 (O_868,N_9440,N_9304);
nor UO_869 (O_869,N_8963,N_9821);
and UO_870 (O_870,N_8413,N_8485);
and UO_871 (O_871,N_8248,N_9971);
nand UO_872 (O_872,N_8532,N_9581);
nor UO_873 (O_873,N_8564,N_9560);
nor UO_874 (O_874,N_9226,N_8589);
nand UO_875 (O_875,N_8832,N_8643);
nor UO_876 (O_876,N_8446,N_9743);
or UO_877 (O_877,N_9183,N_8983);
or UO_878 (O_878,N_8220,N_9150);
nand UO_879 (O_879,N_8715,N_9555);
nor UO_880 (O_880,N_8382,N_9877);
nand UO_881 (O_881,N_9864,N_9887);
or UO_882 (O_882,N_8075,N_8531);
nor UO_883 (O_883,N_9359,N_8183);
nand UO_884 (O_884,N_9139,N_9683);
and UO_885 (O_885,N_8149,N_9529);
or UO_886 (O_886,N_8137,N_9423);
nand UO_887 (O_887,N_9976,N_9120);
nor UO_888 (O_888,N_8980,N_8209);
nor UO_889 (O_889,N_9154,N_9443);
nor UO_890 (O_890,N_9713,N_9053);
and UO_891 (O_891,N_9580,N_8144);
nor UO_892 (O_892,N_8325,N_9263);
or UO_893 (O_893,N_8256,N_8585);
or UO_894 (O_894,N_8638,N_8540);
nor UO_895 (O_895,N_8795,N_8496);
nor UO_896 (O_896,N_9896,N_8393);
xnor UO_897 (O_897,N_8076,N_8357);
nor UO_898 (O_898,N_9876,N_9850);
xnor UO_899 (O_899,N_8337,N_8820);
nor UO_900 (O_900,N_9433,N_9669);
nor UO_901 (O_901,N_9714,N_9277);
nor UO_902 (O_902,N_9520,N_9133);
nand UO_903 (O_903,N_8065,N_8837);
nand UO_904 (O_904,N_9515,N_9993);
and UO_905 (O_905,N_8430,N_8204);
and UO_906 (O_906,N_9961,N_9200);
nor UO_907 (O_907,N_8359,N_9250);
or UO_908 (O_908,N_9746,N_9968);
nand UO_909 (O_909,N_9643,N_8790);
or UO_910 (O_910,N_9136,N_9658);
or UO_911 (O_911,N_9536,N_8177);
or UO_912 (O_912,N_8164,N_8571);
or UO_913 (O_913,N_9394,N_8306);
and UO_914 (O_914,N_8230,N_8687);
and UO_915 (O_915,N_8429,N_8062);
and UO_916 (O_916,N_9509,N_8423);
nor UO_917 (O_917,N_8471,N_8774);
nor UO_918 (O_918,N_9923,N_9649);
and UO_919 (O_919,N_8912,N_8274);
nand UO_920 (O_920,N_9409,N_9804);
nand UO_921 (O_921,N_9659,N_8659);
nand UO_922 (O_922,N_9680,N_9950);
nor UO_923 (O_923,N_9618,N_8369);
and UO_924 (O_924,N_8494,N_9970);
and UO_925 (O_925,N_9688,N_9947);
or UO_926 (O_926,N_9901,N_9337);
or UO_927 (O_927,N_8535,N_8922);
nand UO_928 (O_928,N_9292,N_8551);
or UO_929 (O_929,N_9957,N_9088);
and UO_930 (O_930,N_8760,N_9189);
nand UO_931 (O_931,N_9353,N_9387);
nand UO_932 (O_932,N_8255,N_9381);
and UO_933 (O_933,N_9261,N_8340);
or UO_934 (O_934,N_9431,N_9037);
nor UO_935 (O_935,N_9081,N_9074);
and UO_936 (O_936,N_8319,N_9496);
and UO_937 (O_937,N_9338,N_8950);
and UO_938 (O_938,N_9724,N_8196);
nand UO_939 (O_939,N_9785,N_9242);
nand UO_940 (O_940,N_9197,N_9191);
or UO_941 (O_941,N_9734,N_8440);
nor UO_942 (O_942,N_8588,N_8015);
or UO_943 (O_943,N_9426,N_8942);
or UO_944 (O_944,N_9117,N_9953);
nor UO_945 (O_945,N_9364,N_8803);
nand UO_946 (O_946,N_9134,N_8605);
or UO_947 (O_947,N_8318,N_9076);
nor UO_948 (O_948,N_9063,N_9874);
nand UO_949 (O_949,N_8116,N_8131);
nor UO_950 (O_950,N_9247,N_8229);
or UO_951 (O_951,N_9379,N_8421);
and UO_952 (O_952,N_8806,N_8419);
and UO_953 (O_953,N_9899,N_8112);
nand UO_954 (O_954,N_9645,N_8954);
or UO_955 (O_955,N_9756,N_8385);
nand UO_956 (O_956,N_8794,N_9448);
nor UO_957 (O_957,N_9919,N_8547);
or UO_958 (O_958,N_9470,N_8459);
or UO_959 (O_959,N_8544,N_9573);
nand UO_960 (O_960,N_9070,N_9378);
nand UO_961 (O_961,N_8840,N_9844);
or UO_962 (O_962,N_9491,N_9739);
or UO_963 (O_963,N_9798,N_9211);
and UO_964 (O_964,N_8493,N_8804);
or UO_965 (O_965,N_8549,N_8960);
or UO_966 (O_966,N_8526,N_8314);
nor UO_967 (O_967,N_8201,N_9729);
and UO_968 (O_968,N_9370,N_8849);
or UO_969 (O_969,N_9398,N_9274);
nand UO_970 (O_970,N_8324,N_9776);
nand UO_971 (O_971,N_8424,N_9368);
nand UO_972 (O_972,N_9369,N_8373);
and UO_973 (O_973,N_9202,N_9207);
nand UO_974 (O_974,N_9747,N_8662);
and UO_975 (O_975,N_8118,N_9602);
and UO_976 (O_976,N_9413,N_9800);
and UO_977 (O_977,N_9192,N_8595);
nand UO_978 (O_978,N_8753,N_8312);
nand UO_979 (O_979,N_8690,N_8568);
nor UO_980 (O_980,N_8077,N_8556);
or UO_981 (O_981,N_8497,N_9663);
nand UO_982 (O_982,N_9484,N_9218);
nand UO_983 (O_983,N_9791,N_9647);
nor UO_984 (O_984,N_9959,N_8057);
or UO_985 (O_985,N_9330,N_8297);
and UO_986 (O_986,N_9831,N_8260);
nor UO_987 (O_987,N_9921,N_8770);
nand UO_988 (O_988,N_9648,N_9712);
nand UO_989 (O_989,N_9510,N_9295);
nand UO_990 (O_990,N_8272,N_9594);
nand UO_991 (O_991,N_9367,N_8080);
nor UO_992 (O_992,N_8627,N_9233);
and UO_993 (O_993,N_9012,N_9305);
and UO_994 (O_994,N_9476,N_8825);
and UO_995 (O_995,N_9388,N_8231);
nor UO_996 (O_996,N_9205,N_8476);
nor UO_997 (O_997,N_8014,N_8857);
and UO_998 (O_998,N_9912,N_8982);
and UO_999 (O_999,N_9882,N_9708);
and UO_1000 (O_1000,N_9270,N_8769);
or UO_1001 (O_1001,N_9626,N_9581);
and UO_1002 (O_1002,N_9821,N_8288);
or UO_1003 (O_1003,N_9251,N_9905);
or UO_1004 (O_1004,N_9701,N_8905);
and UO_1005 (O_1005,N_9189,N_9989);
and UO_1006 (O_1006,N_9470,N_9338);
nand UO_1007 (O_1007,N_8963,N_9116);
or UO_1008 (O_1008,N_8401,N_8468);
and UO_1009 (O_1009,N_8725,N_8090);
or UO_1010 (O_1010,N_8286,N_9017);
nor UO_1011 (O_1011,N_9543,N_9800);
nor UO_1012 (O_1012,N_8438,N_8071);
or UO_1013 (O_1013,N_8301,N_9076);
nand UO_1014 (O_1014,N_9111,N_9522);
nand UO_1015 (O_1015,N_8313,N_8942);
or UO_1016 (O_1016,N_9971,N_8544);
nand UO_1017 (O_1017,N_9200,N_9195);
nand UO_1018 (O_1018,N_9877,N_9569);
xnor UO_1019 (O_1019,N_8259,N_9598);
or UO_1020 (O_1020,N_9874,N_8579);
or UO_1021 (O_1021,N_9474,N_9663);
and UO_1022 (O_1022,N_9641,N_9628);
or UO_1023 (O_1023,N_9921,N_8379);
nor UO_1024 (O_1024,N_8385,N_9596);
nor UO_1025 (O_1025,N_8503,N_9735);
or UO_1026 (O_1026,N_8951,N_8307);
nand UO_1027 (O_1027,N_9895,N_9465);
and UO_1028 (O_1028,N_8690,N_8041);
or UO_1029 (O_1029,N_9078,N_8202);
nand UO_1030 (O_1030,N_8616,N_9610);
or UO_1031 (O_1031,N_8930,N_9007);
nand UO_1032 (O_1032,N_9483,N_8818);
and UO_1033 (O_1033,N_8645,N_8890);
nand UO_1034 (O_1034,N_8132,N_9370);
or UO_1035 (O_1035,N_9704,N_8204);
nor UO_1036 (O_1036,N_8817,N_8194);
nand UO_1037 (O_1037,N_8761,N_8465);
and UO_1038 (O_1038,N_9594,N_9055);
nand UO_1039 (O_1039,N_9392,N_8693);
or UO_1040 (O_1040,N_8198,N_8296);
xor UO_1041 (O_1041,N_9807,N_8066);
or UO_1042 (O_1042,N_9278,N_9381);
or UO_1043 (O_1043,N_8298,N_8520);
nor UO_1044 (O_1044,N_8622,N_8198);
and UO_1045 (O_1045,N_9425,N_9620);
nor UO_1046 (O_1046,N_9417,N_8171);
nand UO_1047 (O_1047,N_8415,N_8681);
or UO_1048 (O_1048,N_9295,N_9613);
and UO_1049 (O_1049,N_9774,N_8515);
nor UO_1050 (O_1050,N_8563,N_8794);
nand UO_1051 (O_1051,N_8185,N_8855);
nand UO_1052 (O_1052,N_8430,N_8012);
or UO_1053 (O_1053,N_9928,N_8793);
nor UO_1054 (O_1054,N_9513,N_9501);
nor UO_1055 (O_1055,N_8337,N_8513);
and UO_1056 (O_1056,N_8440,N_8685);
or UO_1057 (O_1057,N_8775,N_9509);
nor UO_1058 (O_1058,N_8371,N_9450);
nor UO_1059 (O_1059,N_9774,N_8956);
nor UO_1060 (O_1060,N_9821,N_8735);
nand UO_1061 (O_1061,N_9519,N_9071);
and UO_1062 (O_1062,N_9915,N_8953);
or UO_1063 (O_1063,N_8466,N_8668);
nor UO_1064 (O_1064,N_8816,N_8404);
nand UO_1065 (O_1065,N_9768,N_9443);
nor UO_1066 (O_1066,N_9363,N_8067);
nor UO_1067 (O_1067,N_8255,N_9029);
and UO_1068 (O_1068,N_8610,N_9991);
and UO_1069 (O_1069,N_8634,N_9282);
or UO_1070 (O_1070,N_9109,N_9169);
xnor UO_1071 (O_1071,N_9243,N_8733);
and UO_1072 (O_1072,N_8310,N_9148);
nand UO_1073 (O_1073,N_9314,N_9794);
nand UO_1074 (O_1074,N_9826,N_9081);
and UO_1075 (O_1075,N_9430,N_9881);
and UO_1076 (O_1076,N_8877,N_9267);
nand UO_1077 (O_1077,N_9669,N_9036);
nor UO_1078 (O_1078,N_9865,N_8865);
or UO_1079 (O_1079,N_8984,N_8488);
nor UO_1080 (O_1080,N_9271,N_9545);
or UO_1081 (O_1081,N_8050,N_8356);
nand UO_1082 (O_1082,N_9579,N_8738);
nor UO_1083 (O_1083,N_8392,N_8438);
xor UO_1084 (O_1084,N_9573,N_8341);
or UO_1085 (O_1085,N_8950,N_8893);
nor UO_1086 (O_1086,N_9337,N_9292);
or UO_1087 (O_1087,N_9400,N_8684);
or UO_1088 (O_1088,N_8111,N_8324);
or UO_1089 (O_1089,N_8813,N_8387);
nand UO_1090 (O_1090,N_9126,N_9221);
and UO_1091 (O_1091,N_8336,N_8219);
and UO_1092 (O_1092,N_9911,N_8311);
nor UO_1093 (O_1093,N_8394,N_8160);
and UO_1094 (O_1094,N_9400,N_9761);
nand UO_1095 (O_1095,N_9801,N_9369);
or UO_1096 (O_1096,N_9021,N_8953);
nand UO_1097 (O_1097,N_9011,N_8167);
nand UO_1098 (O_1098,N_9605,N_8498);
nand UO_1099 (O_1099,N_9907,N_8377);
nor UO_1100 (O_1100,N_9056,N_9237);
nor UO_1101 (O_1101,N_8703,N_8439);
nand UO_1102 (O_1102,N_8827,N_9396);
or UO_1103 (O_1103,N_8233,N_8683);
nand UO_1104 (O_1104,N_8035,N_8187);
nand UO_1105 (O_1105,N_9359,N_9847);
and UO_1106 (O_1106,N_8499,N_9161);
and UO_1107 (O_1107,N_8910,N_8140);
nor UO_1108 (O_1108,N_9983,N_8995);
nand UO_1109 (O_1109,N_8670,N_9647);
xor UO_1110 (O_1110,N_8578,N_8991);
and UO_1111 (O_1111,N_9810,N_9284);
and UO_1112 (O_1112,N_9493,N_9769);
nand UO_1113 (O_1113,N_8483,N_8458);
or UO_1114 (O_1114,N_8099,N_9147);
and UO_1115 (O_1115,N_9883,N_8145);
nor UO_1116 (O_1116,N_8239,N_9276);
or UO_1117 (O_1117,N_8742,N_8140);
and UO_1118 (O_1118,N_9090,N_9407);
nor UO_1119 (O_1119,N_8897,N_8974);
nand UO_1120 (O_1120,N_8253,N_8523);
or UO_1121 (O_1121,N_9154,N_8334);
nand UO_1122 (O_1122,N_9531,N_8562);
nand UO_1123 (O_1123,N_8980,N_9854);
nand UO_1124 (O_1124,N_8570,N_8200);
nand UO_1125 (O_1125,N_9869,N_9614);
or UO_1126 (O_1126,N_9571,N_8032);
and UO_1127 (O_1127,N_8053,N_8751);
nor UO_1128 (O_1128,N_8813,N_8765);
and UO_1129 (O_1129,N_8255,N_8170);
nor UO_1130 (O_1130,N_8261,N_9234);
nand UO_1131 (O_1131,N_8662,N_8846);
nor UO_1132 (O_1132,N_8855,N_8440);
or UO_1133 (O_1133,N_8303,N_9598);
nand UO_1134 (O_1134,N_8205,N_9310);
nor UO_1135 (O_1135,N_8044,N_9223);
nor UO_1136 (O_1136,N_9406,N_8478);
and UO_1137 (O_1137,N_8223,N_9777);
nor UO_1138 (O_1138,N_9294,N_9373);
or UO_1139 (O_1139,N_9389,N_8758);
nand UO_1140 (O_1140,N_8698,N_8280);
or UO_1141 (O_1141,N_9829,N_8481);
and UO_1142 (O_1142,N_9913,N_9890);
nand UO_1143 (O_1143,N_9053,N_9022);
or UO_1144 (O_1144,N_9174,N_8294);
or UO_1145 (O_1145,N_8146,N_8599);
nor UO_1146 (O_1146,N_8879,N_8282);
nor UO_1147 (O_1147,N_9313,N_9789);
nor UO_1148 (O_1148,N_8371,N_9955);
nor UO_1149 (O_1149,N_9716,N_9070);
and UO_1150 (O_1150,N_8319,N_9114);
nor UO_1151 (O_1151,N_9648,N_9089);
nand UO_1152 (O_1152,N_8421,N_8025);
nand UO_1153 (O_1153,N_8033,N_9738);
nand UO_1154 (O_1154,N_9820,N_9160);
nor UO_1155 (O_1155,N_8578,N_8350);
or UO_1156 (O_1156,N_8495,N_9906);
and UO_1157 (O_1157,N_8732,N_8666);
nor UO_1158 (O_1158,N_9496,N_9993);
and UO_1159 (O_1159,N_8767,N_8330);
nor UO_1160 (O_1160,N_8331,N_9940);
and UO_1161 (O_1161,N_8809,N_8515);
or UO_1162 (O_1162,N_9083,N_8037);
nor UO_1163 (O_1163,N_9940,N_8171);
nand UO_1164 (O_1164,N_9487,N_9806);
nor UO_1165 (O_1165,N_8150,N_8009);
nand UO_1166 (O_1166,N_8210,N_8614);
and UO_1167 (O_1167,N_8234,N_8068);
and UO_1168 (O_1168,N_9130,N_9372);
nand UO_1169 (O_1169,N_8277,N_8243);
and UO_1170 (O_1170,N_9311,N_9512);
nand UO_1171 (O_1171,N_8437,N_8156);
and UO_1172 (O_1172,N_9633,N_9276);
nor UO_1173 (O_1173,N_8643,N_8793);
and UO_1174 (O_1174,N_9843,N_9654);
nand UO_1175 (O_1175,N_9497,N_9484);
or UO_1176 (O_1176,N_9863,N_8506);
and UO_1177 (O_1177,N_8947,N_9001);
or UO_1178 (O_1178,N_9353,N_8574);
and UO_1179 (O_1179,N_9086,N_8833);
nor UO_1180 (O_1180,N_8738,N_9948);
nor UO_1181 (O_1181,N_8452,N_9204);
nand UO_1182 (O_1182,N_8565,N_9913);
nand UO_1183 (O_1183,N_9878,N_8538);
and UO_1184 (O_1184,N_8890,N_8863);
nor UO_1185 (O_1185,N_9504,N_9164);
or UO_1186 (O_1186,N_8276,N_9286);
and UO_1187 (O_1187,N_9673,N_8833);
and UO_1188 (O_1188,N_9539,N_8815);
or UO_1189 (O_1189,N_9633,N_8935);
nor UO_1190 (O_1190,N_9383,N_8527);
or UO_1191 (O_1191,N_8814,N_8213);
xor UO_1192 (O_1192,N_8855,N_8218);
or UO_1193 (O_1193,N_8062,N_8756);
nand UO_1194 (O_1194,N_9711,N_8114);
or UO_1195 (O_1195,N_9659,N_9129);
and UO_1196 (O_1196,N_8339,N_8836);
nand UO_1197 (O_1197,N_8633,N_8567);
and UO_1198 (O_1198,N_9098,N_9321);
or UO_1199 (O_1199,N_9228,N_8423);
nand UO_1200 (O_1200,N_9605,N_8387);
or UO_1201 (O_1201,N_8547,N_8100);
nand UO_1202 (O_1202,N_9803,N_8827);
nand UO_1203 (O_1203,N_9169,N_8768);
and UO_1204 (O_1204,N_8019,N_8016);
or UO_1205 (O_1205,N_9836,N_8830);
nor UO_1206 (O_1206,N_9707,N_9956);
nand UO_1207 (O_1207,N_9567,N_9542);
nor UO_1208 (O_1208,N_8422,N_9238);
or UO_1209 (O_1209,N_8321,N_8208);
nor UO_1210 (O_1210,N_9669,N_8690);
nand UO_1211 (O_1211,N_8343,N_8865);
or UO_1212 (O_1212,N_9859,N_9407);
nand UO_1213 (O_1213,N_9535,N_8505);
xnor UO_1214 (O_1214,N_8750,N_8345);
or UO_1215 (O_1215,N_8827,N_8276);
nand UO_1216 (O_1216,N_9787,N_9572);
nand UO_1217 (O_1217,N_9242,N_8159);
nand UO_1218 (O_1218,N_8131,N_8234);
nor UO_1219 (O_1219,N_9805,N_8394);
nor UO_1220 (O_1220,N_8512,N_9094);
or UO_1221 (O_1221,N_9027,N_8647);
and UO_1222 (O_1222,N_8562,N_8854);
xor UO_1223 (O_1223,N_8036,N_8688);
nand UO_1224 (O_1224,N_9567,N_9279);
or UO_1225 (O_1225,N_8090,N_9895);
and UO_1226 (O_1226,N_9954,N_9511);
nor UO_1227 (O_1227,N_9888,N_9942);
nor UO_1228 (O_1228,N_8796,N_8232);
nand UO_1229 (O_1229,N_8293,N_8922);
nand UO_1230 (O_1230,N_8374,N_9331);
and UO_1231 (O_1231,N_9092,N_8013);
nor UO_1232 (O_1232,N_9434,N_9535);
or UO_1233 (O_1233,N_8185,N_9423);
nor UO_1234 (O_1234,N_9462,N_9063);
nor UO_1235 (O_1235,N_9073,N_8057);
and UO_1236 (O_1236,N_8733,N_9442);
nand UO_1237 (O_1237,N_9927,N_9622);
or UO_1238 (O_1238,N_8311,N_9473);
nand UO_1239 (O_1239,N_9901,N_8044);
and UO_1240 (O_1240,N_8416,N_8932);
nor UO_1241 (O_1241,N_9195,N_9359);
nand UO_1242 (O_1242,N_9392,N_8503);
nor UO_1243 (O_1243,N_8621,N_9497);
nand UO_1244 (O_1244,N_9060,N_8956);
or UO_1245 (O_1245,N_8100,N_9173);
or UO_1246 (O_1246,N_8963,N_9454);
nor UO_1247 (O_1247,N_9772,N_8509);
or UO_1248 (O_1248,N_9400,N_9404);
or UO_1249 (O_1249,N_8553,N_9354);
nor UO_1250 (O_1250,N_9070,N_8023);
xor UO_1251 (O_1251,N_8550,N_9698);
nor UO_1252 (O_1252,N_8411,N_8654);
and UO_1253 (O_1253,N_8928,N_8358);
or UO_1254 (O_1254,N_8099,N_9486);
and UO_1255 (O_1255,N_8414,N_9445);
nor UO_1256 (O_1256,N_8159,N_8025);
or UO_1257 (O_1257,N_8425,N_9357);
nand UO_1258 (O_1258,N_8976,N_9964);
and UO_1259 (O_1259,N_9501,N_8791);
or UO_1260 (O_1260,N_9961,N_9678);
nor UO_1261 (O_1261,N_8875,N_8234);
nor UO_1262 (O_1262,N_8619,N_9168);
and UO_1263 (O_1263,N_9152,N_8722);
nor UO_1264 (O_1264,N_9349,N_9700);
and UO_1265 (O_1265,N_8457,N_9619);
nand UO_1266 (O_1266,N_9587,N_9254);
nor UO_1267 (O_1267,N_9673,N_9276);
and UO_1268 (O_1268,N_8464,N_9455);
nand UO_1269 (O_1269,N_9361,N_9444);
and UO_1270 (O_1270,N_9438,N_9014);
or UO_1271 (O_1271,N_8799,N_8800);
or UO_1272 (O_1272,N_9068,N_9376);
nand UO_1273 (O_1273,N_8277,N_9415);
nor UO_1274 (O_1274,N_8835,N_9966);
nand UO_1275 (O_1275,N_8629,N_9971);
xnor UO_1276 (O_1276,N_8326,N_9765);
nor UO_1277 (O_1277,N_8535,N_8090);
or UO_1278 (O_1278,N_8818,N_9273);
nand UO_1279 (O_1279,N_8729,N_8442);
nor UO_1280 (O_1280,N_8311,N_8919);
and UO_1281 (O_1281,N_9256,N_9860);
nor UO_1282 (O_1282,N_9457,N_8441);
and UO_1283 (O_1283,N_9703,N_9437);
nand UO_1284 (O_1284,N_8477,N_8909);
and UO_1285 (O_1285,N_9437,N_9109);
and UO_1286 (O_1286,N_9945,N_9230);
and UO_1287 (O_1287,N_9898,N_9216);
nand UO_1288 (O_1288,N_8307,N_8616);
nand UO_1289 (O_1289,N_9681,N_9473);
nor UO_1290 (O_1290,N_8681,N_9276);
or UO_1291 (O_1291,N_8439,N_9347);
or UO_1292 (O_1292,N_9861,N_9338);
xnor UO_1293 (O_1293,N_8215,N_9610);
nand UO_1294 (O_1294,N_8273,N_9777);
nor UO_1295 (O_1295,N_9299,N_8697);
and UO_1296 (O_1296,N_9268,N_9445);
or UO_1297 (O_1297,N_8859,N_9686);
or UO_1298 (O_1298,N_9635,N_9221);
and UO_1299 (O_1299,N_9647,N_8648);
nor UO_1300 (O_1300,N_9442,N_8550);
or UO_1301 (O_1301,N_9596,N_8585);
nand UO_1302 (O_1302,N_8094,N_9676);
or UO_1303 (O_1303,N_8196,N_9257);
xor UO_1304 (O_1304,N_8484,N_8466);
nand UO_1305 (O_1305,N_9906,N_8597);
nand UO_1306 (O_1306,N_8659,N_9057);
xnor UO_1307 (O_1307,N_8282,N_8215);
or UO_1308 (O_1308,N_9714,N_8548);
nor UO_1309 (O_1309,N_8807,N_9275);
and UO_1310 (O_1310,N_8710,N_8016);
nand UO_1311 (O_1311,N_9318,N_8847);
nand UO_1312 (O_1312,N_9650,N_9331);
and UO_1313 (O_1313,N_9230,N_9377);
nor UO_1314 (O_1314,N_9474,N_9874);
nand UO_1315 (O_1315,N_9089,N_8224);
nand UO_1316 (O_1316,N_9106,N_9879);
nand UO_1317 (O_1317,N_8000,N_8373);
and UO_1318 (O_1318,N_8383,N_9047);
or UO_1319 (O_1319,N_9173,N_8367);
or UO_1320 (O_1320,N_9107,N_9615);
nor UO_1321 (O_1321,N_8821,N_8033);
nand UO_1322 (O_1322,N_8695,N_8744);
or UO_1323 (O_1323,N_8954,N_9622);
nand UO_1324 (O_1324,N_9813,N_9805);
nand UO_1325 (O_1325,N_8396,N_9679);
or UO_1326 (O_1326,N_9468,N_9345);
nand UO_1327 (O_1327,N_9751,N_9842);
or UO_1328 (O_1328,N_8531,N_8446);
nor UO_1329 (O_1329,N_8297,N_9214);
and UO_1330 (O_1330,N_8921,N_8574);
xnor UO_1331 (O_1331,N_9155,N_9842);
nor UO_1332 (O_1332,N_8756,N_9237);
nor UO_1333 (O_1333,N_9112,N_8430);
or UO_1334 (O_1334,N_8067,N_8752);
nor UO_1335 (O_1335,N_9547,N_8023);
or UO_1336 (O_1336,N_9077,N_9784);
or UO_1337 (O_1337,N_8381,N_8388);
nor UO_1338 (O_1338,N_8582,N_9377);
nand UO_1339 (O_1339,N_8362,N_8848);
nor UO_1340 (O_1340,N_8512,N_8557);
nand UO_1341 (O_1341,N_9755,N_8749);
and UO_1342 (O_1342,N_8591,N_8793);
or UO_1343 (O_1343,N_8929,N_8238);
nand UO_1344 (O_1344,N_9436,N_9481);
nor UO_1345 (O_1345,N_9479,N_9209);
nor UO_1346 (O_1346,N_8624,N_8758);
nand UO_1347 (O_1347,N_8272,N_8336);
or UO_1348 (O_1348,N_9778,N_9435);
nor UO_1349 (O_1349,N_9840,N_9398);
nor UO_1350 (O_1350,N_9610,N_9863);
or UO_1351 (O_1351,N_9500,N_8860);
xnor UO_1352 (O_1352,N_8587,N_8131);
and UO_1353 (O_1353,N_9673,N_8862);
and UO_1354 (O_1354,N_8074,N_9998);
or UO_1355 (O_1355,N_8388,N_9089);
and UO_1356 (O_1356,N_9066,N_9560);
nor UO_1357 (O_1357,N_8857,N_8670);
and UO_1358 (O_1358,N_8116,N_8090);
nor UO_1359 (O_1359,N_9470,N_9231);
nor UO_1360 (O_1360,N_8805,N_9761);
nand UO_1361 (O_1361,N_8285,N_8808);
and UO_1362 (O_1362,N_8890,N_9289);
or UO_1363 (O_1363,N_8672,N_9687);
or UO_1364 (O_1364,N_9984,N_9670);
or UO_1365 (O_1365,N_9962,N_8727);
nor UO_1366 (O_1366,N_9966,N_8121);
or UO_1367 (O_1367,N_8427,N_8171);
nor UO_1368 (O_1368,N_9882,N_8830);
nor UO_1369 (O_1369,N_9017,N_9979);
and UO_1370 (O_1370,N_9403,N_8370);
or UO_1371 (O_1371,N_8703,N_9524);
xor UO_1372 (O_1372,N_8624,N_9447);
nand UO_1373 (O_1373,N_9336,N_8500);
nor UO_1374 (O_1374,N_9921,N_8864);
nand UO_1375 (O_1375,N_9984,N_8714);
and UO_1376 (O_1376,N_9000,N_9576);
nor UO_1377 (O_1377,N_9037,N_8498);
nand UO_1378 (O_1378,N_8747,N_8639);
or UO_1379 (O_1379,N_9366,N_9405);
nand UO_1380 (O_1380,N_9289,N_8759);
nand UO_1381 (O_1381,N_9047,N_9036);
and UO_1382 (O_1382,N_8331,N_9930);
nand UO_1383 (O_1383,N_8220,N_8612);
xnor UO_1384 (O_1384,N_8204,N_8796);
or UO_1385 (O_1385,N_9533,N_9811);
nand UO_1386 (O_1386,N_8597,N_8321);
nor UO_1387 (O_1387,N_8703,N_8580);
or UO_1388 (O_1388,N_8579,N_9519);
nand UO_1389 (O_1389,N_8185,N_8188);
or UO_1390 (O_1390,N_9200,N_8584);
nand UO_1391 (O_1391,N_9478,N_8423);
and UO_1392 (O_1392,N_8088,N_8275);
nor UO_1393 (O_1393,N_8755,N_8319);
nand UO_1394 (O_1394,N_9269,N_9874);
or UO_1395 (O_1395,N_9932,N_8739);
and UO_1396 (O_1396,N_8336,N_9649);
and UO_1397 (O_1397,N_9991,N_8326);
or UO_1398 (O_1398,N_8764,N_9598);
nor UO_1399 (O_1399,N_8845,N_9890);
nor UO_1400 (O_1400,N_9001,N_8043);
nand UO_1401 (O_1401,N_9961,N_8557);
nor UO_1402 (O_1402,N_8856,N_9626);
xor UO_1403 (O_1403,N_9814,N_8108);
or UO_1404 (O_1404,N_8208,N_8859);
nand UO_1405 (O_1405,N_9735,N_9638);
and UO_1406 (O_1406,N_8433,N_8176);
nor UO_1407 (O_1407,N_9225,N_8113);
or UO_1408 (O_1408,N_8448,N_8061);
and UO_1409 (O_1409,N_8731,N_9620);
and UO_1410 (O_1410,N_9167,N_8917);
nand UO_1411 (O_1411,N_8912,N_9046);
or UO_1412 (O_1412,N_9062,N_9835);
or UO_1413 (O_1413,N_8671,N_9253);
and UO_1414 (O_1414,N_9157,N_8448);
or UO_1415 (O_1415,N_9555,N_9190);
and UO_1416 (O_1416,N_9990,N_8672);
and UO_1417 (O_1417,N_8305,N_9837);
and UO_1418 (O_1418,N_9169,N_8181);
and UO_1419 (O_1419,N_8087,N_8561);
nor UO_1420 (O_1420,N_8606,N_9499);
and UO_1421 (O_1421,N_9639,N_9599);
nand UO_1422 (O_1422,N_8795,N_9877);
nor UO_1423 (O_1423,N_9028,N_9291);
or UO_1424 (O_1424,N_9592,N_9649);
or UO_1425 (O_1425,N_8405,N_9118);
or UO_1426 (O_1426,N_8604,N_9101);
and UO_1427 (O_1427,N_8325,N_8401);
or UO_1428 (O_1428,N_9386,N_8577);
and UO_1429 (O_1429,N_9380,N_8496);
nor UO_1430 (O_1430,N_9950,N_9526);
nor UO_1431 (O_1431,N_9267,N_9329);
nor UO_1432 (O_1432,N_9159,N_9478);
and UO_1433 (O_1433,N_9439,N_9680);
nand UO_1434 (O_1434,N_8892,N_8714);
and UO_1435 (O_1435,N_9128,N_8711);
and UO_1436 (O_1436,N_9744,N_9686);
and UO_1437 (O_1437,N_8192,N_9507);
and UO_1438 (O_1438,N_8939,N_8736);
nor UO_1439 (O_1439,N_9082,N_9840);
nand UO_1440 (O_1440,N_8102,N_8492);
and UO_1441 (O_1441,N_9350,N_8471);
nor UO_1442 (O_1442,N_8945,N_9954);
and UO_1443 (O_1443,N_8570,N_8855);
nor UO_1444 (O_1444,N_8674,N_9600);
nand UO_1445 (O_1445,N_9384,N_9452);
and UO_1446 (O_1446,N_8523,N_9522);
or UO_1447 (O_1447,N_9184,N_8854);
nor UO_1448 (O_1448,N_8063,N_9294);
or UO_1449 (O_1449,N_8357,N_9013);
and UO_1450 (O_1450,N_8114,N_8170);
or UO_1451 (O_1451,N_8713,N_8888);
nand UO_1452 (O_1452,N_9227,N_8344);
nor UO_1453 (O_1453,N_9433,N_8563);
nor UO_1454 (O_1454,N_8986,N_9295);
xor UO_1455 (O_1455,N_8904,N_9238);
or UO_1456 (O_1456,N_8897,N_8411);
or UO_1457 (O_1457,N_9192,N_9033);
nand UO_1458 (O_1458,N_9369,N_9786);
nand UO_1459 (O_1459,N_9502,N_9075);
or UO_1460 (O_1460,N_9625,N_8811);
nand UO_1461 (O_1461,N_8926,N_8479);
nor UO_1462 (O_1462,N_8650,N_9773);
and UO_1463 (O_1463,N_8421,N_9948);
and UO_1464 (O_1464,N_8486,N_8851);
and UO_1465 (O_1465,N_9243,N_9458);
and UO_1466 (O_1466,N_9536,N_8885);
nand UO_1467 (O_1467,N_8371,N_8568);
nor UO_1468 (O_1468,N_8488,N_8724);
or UO_1469 (O_1469,N_8242,N_9146);
and UO_1470 (O_1470,N_8148,N_9362);
nand UO_1471 (O_1471,N_8881,N_8620);
nor UO_1472 (O_1472,N_8010,N_8448);
or UO_1473 (O_1473,N_8910,N_8310);
nand UO_1474 (O_1474,N_9801,N_9859);
and UO_1475 (O_1475,N_9285,N_8254);
nand UO_1476 (O_1476,N_8235,N_9088);
and UO_1477 (O_1477,N_8781,N_9812);
nor UO_1478 (O_1478,N_9811,N_9735);
nand UO_1479 (O_1479,N_9991,N_9895);
and UO_1480 (O_1480,N_9692,N_9700);
or UO_1481 (O_1481,N_9039,N_8595);
nand UO_1482 (O_1482,N_8687,N_9717);
nand UO_1483 (O_1483,N_8066,N_8928);
nand UO_1484 (O_1484,N_8918,N_9615);
nor UO_1485 (O_1485,N_9897,N_9687);
nand UO_1486 (O_1486,N_9923,N_9412);
nor UO_1487 (O_1487,N_8842,N_8361);
nand UO_1488 (O_1488,N_8947,N_9176);
nand UO_1489 (O_1489,N_9020,N_8978);
and UO_1490 (O_1490,N_8182,N_9139);
nor UO_1491 (O_1491,N_9559,N_9291);
and UO_1492 (O_1492,N_9526,N_9171);
nor UO_1493 (O_1493,N_9994,N_8974);
and UO_1494 (O_1494,N_9667,N_9615);
or UO_1495 (O_1495,N_8864,N_8140);
and UO_1496 (O_1496,N_8761,N_8082);
nand UO_1497 (O_1497,N_9381,N_8043);
or UO_1498 (O_1498,N_9209,N_8910);
or UO_1499 (O_1499,N_9005,N_9828);
endmodule