module basic_2000_20000_2500_4_levels_1xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
and U0 (N_0,In_46,In_1507);
or U1 (N_1,In_547,In_599);
and U2 (N_2,In_1376,In_658);
or U3 (N_3,In_575,In_886);
nand U4 (N_4,In_398,In_1010);
nand U5 (N_5,In_168,In_1736);
nor U6 (N_6,In_96,In_1346);
or U7 (N_7,In_1598,In_1636);
nor U8 (N_8,In_432,In_955);
nor U9 (N_9,In_188,In_1066);
nand U10 (N_10,In_1142,In_277);
nor U11 (N_11,In_1664,In_1472);
nor U12 (N_12,In_1498,In_238);
and U13 (N_13,In_267,In_996);
or U14 (N_14,In_1063,In_1169);
or U15 (N_15,In_1809,In_1709);
nor U16 (N_16,In_1785,In_889);
nor U17 (N_17,In_1547,In_1108);
xnor U18 (N_18,In_1612,In_607);
and U19 (N_19,In_1482,In_1445);
nand U20 (N_20,In_1077,In_1470);
nand U21 (N_21,In_287,In_1473);
nor U22 (N_22,In_1048,In_1533);
or U23 (N_23,In_483,In_486);
or U24 (N_24,In_278,In_581);
nand U25 (N_25,In_1509,In_985);
nor U26 (N_26,In_1041,In_1002);
xnor U27 (N_27,In_951,In_691);
or U28 (N_28,In_1278,In_1946);
or U29 (N_29,In_733,In_121);
nor U30 (N_30,In_1984,In_1361);
nor U31 (N_31,In_674,In_1592);
and U32 (N_32,In_353,In_1569);
nand U33 (N_33,In_846,In_364);
nand U34 (N_34,In_373,In_1495);
and U35 (N_35,In_1799,In_103);
nor U36 (N_36,In_781,In_1735);
nor U37 (N_37,In_1618,In_1317);
nand U38 (N_38,In_617,In_98);
nand U39 (N_39,In_1730,In_1577);
nor U40 (N_40,In_1893,In_1170);
or U41 (N_41,In_1897,In_427);
nor U42 (N_42,In_1739,In_895);
nand U43 (N_43,In_945,In_331);
and U44 (N_44,In_196,In_653);
nor U45 (N_45,In_295,In_1012);
nand U46 (N_46,In_828,In_1844);
or U47 (N_47,In_150,In_19);
and U48 (N_48,In_700,In_1476);
nor U49 (N_49,In_181,In_642);
nor U50 (N_50,In_975,In_988);
nand U51 (N_51,In_1798,In_1653);
nand U52 (N_52,In_1028,In_167);
nor U53 (N_53,In_1816,In_28);
and U54 (N_54,In_134,In_1997);
or U55 (N_55,In_1995,In_294);
nand U56 (N_56,In_803,In_860);
nand U57 (N_57,In_527,In_1761);
or U58 (N_58,In_237,In_419);
and U59 (N_59,In_1585,In_913);
or U60 (N_60,In_990,In_980);
and U61 (N_61,In_1033,In_1682);
and U62 (N_62,In_1345,In_810);
and U63 (N_63,In_1936,In_1680);
nor U64 (N_64,In_564,In_900);
nand U65 (N_65,In_1326,In_887);
nand U66 (N_66,In_548,In_436);
nand U67 (N_67,In_644,In_256);
and U68 (N_68,In_1237,In_54);
or U69 (N_69,In_1433,In_613);
nor U70 (N_70,In_1186,In_1518);
nand U71 (N_71,In_1210,In_589);
or U72 (N_72,In_1502,In_943);
and U73 (N_73,In_762,In_1665);
nand U74 (N_74,In_553,In_709);
nand U75 (N_75,In_624,In_313);
nor U76 (N_76,In_1155,In_1778);
and U77 (N_77,In_588,In_1536);
nor U78 (N_78,In_1973,In_715);
nor U79 (N_79,In_1375,In_1490);
nor U80 (N_80,In_723,In_285);
or U81 (N_81,In_1937,In_1295);
or U82 (N_82,In_1537,In_207);
nand U83 (N_83,In_1694,In_42);
or U84 (N_84,In_494,In_560);
nor U85 (N_85,In_1684,In_1539);
and U86 (N_86,In_471,In_602);
and U87 (N_87,In_1444,In_1707);
or U88 (N_88,In_41,In_1659);
or U89 (N_89,In_571,In_234);
or U90 (N_90,In_920,In_1261);
and U91 (N_91,In_1886,In_119);
nand U92 (N_92,In_1710,In_837);
nor U93 (N_93,In_1681,In_74);
nand U94 (N_94,In_1872,In_378);
or U95 (N_95,In_739,In_123);
nor U96 (N_96,In_515,In_1203);
nor U97 (N_97,In_253,In_429);
and U98 (N_98,In_1934,In_239);
nand U99 (N_99,In_1944,In_9);
and U100 (N_100,In_1296,In_995);
nand U101 (N_101,In_1045,In_898);
and U102 (N_102,In_396,In_355);
and U103 (N_103,In_1905,In_1145);
and U104 (N_104,In_1,In_1439);
or U105 (N_105,In_1561,In_72);
and U106 (N_106,In_1961,In_1136);
and U107 (N_107,In_344,In_879);
or U108 (N_108,In_1581,In_909);
nor U109 (N_109,In_1418,In_1725);
and U110 (N_110,In_1945,In_1738);
nand U111 (N_111,In_540,In_169);
nor U112 (N_112,In_764,In_1545);
nand U113 (N_113,In_844,In_1953);
nand U114 (N_114,In_286,In_482);
nor U115 (N_115,In_790,In_908);
nor U116 (N_116,In_408,In_131);
nor U117 (N_117,In_50,In_941);
and U118 (N_118,In_1718,In_88);
and U119 (N_119,In_1670,In_90);
nand U120 (N_120,In_447,In_1562);
and U121 (N_121,In_1667,In_415);
or U122 (N_122,In_829,In_1020);
or U123 (N_123,In_817,In_437);
or U124 (N_124,In_881,In_276);
nand U125 (N_125,In_1929,In_792);
nand U126 (N_126,In_1051,In_712);
xor U127 (N_127,In_1016,In_1907);
or U128 (N_128,In_274,In_272);
and U129 (N_129,In_1234,In_1001);
nand U130 (N_130,In_1368,In_418);
nor U131 (N_131,In_1546,In_1397);
nor U132 (N_132,In_798,In_1312);
and U133 (N_133,In_978,In_565);
or U134 (N_134,In_1031,In_389);
and U135 (N_135,In_1180,In_1340);
nand U136 (N_136,In_1188,In_680);
or U137 (N_137,In_1752,In_921);
nor U138 (N_138,In_1315,In_580);
nor U139 (N_139,In_485,In_1348);
nand U140 (N_140,In_768,In_620);
or U141 (N_141,In_374,In_750);
nor U142 (N_142,In_209,In_1405);
xnor U143 (N_143,In_1624,In_760);
or U144 (N_144,In_1631,In_965);
and U145 (N_145,In_173,In_1156);
and U146 (N_146,In_1434,In_628);
nor U147 (N_147,In_1733,In_539);
nor U148 (N_148,In_1658,In_1425);
or U149 (N_149,In_651,In_1438);
and U150 (N_150,In_1862,In_962);
nor U151 (N_151,In_214,In_1268);
and U152 (N_152,In_481,In_614);
and U153 (N_153,In_1111,In_1891);
nand U154 (N_154,In_1018,In_967);
and U155 (N_155,In_1780,In_1269);
nand U156 (N_156,In_627,In_1369);
and U157 (N_157,In_81,In_306);
and U158 (N_158,In_1690,In_194);
or U159 (N_159,In_976,In_146);
nand U160 (N_160,In_422,In_1745);
and U161 (N_161,In_1060,In_843);
and U162 (N_162,In_1205,In_1924);
and U163 (N_163,In_915,In_1426);
or U164 (N_164,In_1072,In_155);
nor U165 (N_165,In_280,In_159);
or U166 (N_166,In_1208,In_1055);
or U167 (N_167,In_707,In_635);
nand U168 (N_168,In_1367,In_1892);
and U169 (N_169,In_1480,In_1489);
or U170 (N_170,In_861,In_596);
nand U171 (N_171,In_1305,In_94);
nand U172 (N_172,In_1641,In_337);
nand U173 (N_173,In_732,In_228);
nand U174 (N_174,In_1272,In_1544);
or U175 (N_175,In_1309,In_882);
and U176 (N_176,In_1115,In_1040);
and U177 (N_177,In_672,In_518);
nand U178 (N_178,In_1616,In_690);
and U179 (N_179,In_1906,In_77);
xor U180 (N_180,In_1164,In_724);
nand U181 (N_181,In_25,In_1882);
nand U182 (N_182,In_1042,In_770);
nor U183 (N_183,In_1625,In_1783);
and U184 (N_184,In_1078,In_1231);
nand U185 (N_185,In_1697,In_1527);
and U186 (N_186,In_578,In_821);
and U187 (N_187,In_590,In_1899);
and U188 (N_188,In_749,In_345);
or U189 (N_189,In_1009,In_149);
nor U190 (N_190,In_125,In_1409);
or U191 (N_191,In_1609,In_536);
and U192 (N_192,In_1337,In_328);
nand U193 (N_193,In_323,In_1974);
or U194 (N_194,In_1408,In_1629);
and U195 (N_195,In_1039,In_1091);
and U196 (N_196,In_1611,In_1904);
or U197 (N_197,In_1784,In_1976);
and U198 (N_198,In_1228,In_938);
and U199 (N_199,In_1746,In_1824);
nor U200 (N_200,In_1335,In_761);
xnor U201 (N_201,In_47,In_1271);
nand U202 (N_202,In_1313,In_1558);
nand U203 (N_203,In_1441,In_1004);
nand U204 (N_204,In_603,In_30);
and U205 (N_205,In_44,In_79);
nand U206 (N_206,In_307,In_1727);
and U207 (N_207,In_1298,In_1466);
nand U208 (N_208,In_1711,In_950);
nor U209 (N_209,In_1877,In_1801);
and U210 (N_210,In_314,In_1006);
and U211 (N_211,In_655,In_1255);
or U212 (N_212,In_917,In_457);
nor U213 (N_213,In_891,In_1384);
nor U214 (N_214,In_1525,In_1756);
or U215 (N_215,In_16,In_964);
nor U216 (N_216,In_1771,In_1566);
nor U217 (N_217,In_201,In_1501);
nor U218 (N_218,In_1747,In_1407);
nor U219 (N_219,In_316,In_1233);
nand U220 (N_220,In_394,In_1484);
nand U221 (N_221,In_1206,In_1217);
nor U222 (N_222,In_1097,In_634);
and U223 (N_223,In_302,In_1574);
nand U224 (N_224,In_1822,In_210);
nand U225 (N_225,In_1938,In_431);
nor U226 (N_226,In_1640,In_1879);
and U227 (N_227,In_754,In_893);
nand U228 (N_228,In_1989,In_1182);
nand U229 (N_229,In_1005,In_1549);
or U230 (N_230,In_1227,In_379);
xnor U231 (N_231,In_1493,In_1378);
nand U232 (N_232,In_142,In_1578);
or U233 (N_233,In_960,In_1504);
nand U234 (N_234,In_751,In_1925);
nand U235 (N_235,In_866,In_1957);
or U236 (N_236,In_1845,In_1671);
or U237 (N_237,In_771,In_3);
nor U238 (N_238,In_216,In_1267);
nand U239 (N_239,In_623,In_0);
nand U240 (N_240,In_1417,In_979);
nand U241 (N_241,In_193,In_1692);
nand U242 (N_242,In_1503,In_554);
nand U243 (N_243,In_1095,In_722);
nor U244 (N_244,In_626,In_1543);
and U245 (N_245,In_1793,In_1532);
nand U246 (N_246,In_55,In_877);
and U247 (N_247,In_385,In_442);
nor U248 (N_248,In_959,In_192);
or U249 (N_249,In_1792,In_372);
nor U250 (N_250,In_1068,In_1540);
or U251 (N_251,In_91,In_890);
nor U252 (N_252,In_298,In_1099);
nor U253 (N_253,In_1225,In_139);
and U254 (N_254,In_458,In_641);
nor U255 (N_255,In_530,In_1252);
nor U256 (N_256,In_1332,In_638);
or U257 (N_257,In_75,In_968);
and U258 (N_258,In_80,In_1909);
nor U259 (N_259,In_101,In_692);
and U260 (N_260,In_1633,In_734);
nor U261 (N_261,In_1442,In_1849);
nor U262 (N_262,In_769,In_1555);
and U263 (N_263,In_1486,In_1635);
or U264 (N_264,In_1959,In_1021);
and U265 (N_265,In_1978,In_1122);
and U266 (N_266,In_686,In_1413);
nor U267 (N_267,In_1322,In_1386);
nor U268 (N_268,In_117,In_1732);
or U269 (N_269,In_1400,In_694);
and U270 (N_270,In_1754,In_1123);
nand U271 (N_271,In_594,In_550);
nand U272 (N_272,In_1173,In_296);
and U273 (N_273,In_1406,In_1103);
nand U274 (N_274,In_1679,In_1686);
or U275 (N_275,In_1570,In_802);
and U276 (N_276,In_204,In_1294);
and U277 (N_277,In_217,In_1067);
or U278 (N_278,In_2,In_1150);
nand U279 (N_279,In_1149,In_148);
or U280 (N_280,In_1087,In_1812);
nand U281 (N_281,In_122,In_93);
nand U282 (N_282,In_1782,In_1024);
xnor U283 (N_283,In_1870,In_1120);
xnor U284 (N_284,In_433,In_1204);
or U285 (N_285,In_1435,In_435);
or U286 (N_286,In_1716,In_1483);
nand U287 (N_287,In_868,In_698);
and U288 (N_288,In_794,In_544);
nand U289 (N_289,In_914,In_197);
or U290 (N_290,In_375,In_926);
and U291 (N_291,In_929,In_585);
or U292 (N_292,In_991,In_880);
nor U293 (N_293,In_1791,In_1279);
nor U294 (N_294,In_1963,In_677);
or U295 (N_295,In_450,In_1284);
nand U296 (N_296,In_704,In_649);
nand U297 (N_297,In_1590,In_1837);
nand U298 (N_298,In_1250,In_1669);
or U299 (N_299,In_392,In_1402);
nand U300 (N_300,In_1513,In_521);
nor U301 (N_301,In_1648,In_488);
or U302 (N_302,In_259,In_1875);
nand U303 (N_303,In_555,In_1130);
nand U304 (N_304,In_1049,In_289);
or U305 (N_305,In_1319,In_1253);
nor U306 (N_306,In_789,In_993);
nor U307 (N_307,In_765,In_687);
nor U308 (N_308,In_1787,In_934);
and U309 (N_309,In_832,In_1573);
or U310 (N_310,In_1646,In_947);
or U311 (N_311,In_346,In_386);
and U312 (N_312,In_1596,In_1788);
or U313 (N_313,In_1769,In_543);
and U314 (N_314,In_784,In_775);
nand U315 (N_315,In_693,In_1617);
and U316 (N_316,In_158,In_1919);
and U317 (N_317,In_84,In_1955);
nand U318 (N_318,In_412,In_176);
nor U319 (N_319,In_983,In_1069);
and U320 (N_320,In_291,In_1642);
and U321 (N_321,In_673,In_787);
nand U322 (N_322,In_1510,In_744);
and U323 (N_323,In_1215,In_1750);
nand U324 (N_324,In_1448,In_906);
nor U325 (N_325,In_558,In_1722);
nor U326 (N_326,In_160,In_816);
nor U327 (N_327,In_356,In_1815);
or U328 (N_328,In_939,In_845);
or U329 (N_329,In_1894,In_352);
nor U330 (N_330,In_128,In_1249);
nand U331 (N_331,In_338,In_1548);
and U332 (N_332,In_17,In_714);
nor U333 (N_333,In_927,In_1551);
nor U334 (N_334,In_1918,In_606);
or U335 (N_335,In_533,In_141);
or U336 (N_336,In_1415,In_1007);
and U337 (N_337,In_1129,In_73);
or U338 (N_338,In_466,In_1118);
nor U339 (N_339,In_1096,In_1167);
or U340 (N_340,In_1354,In_166);
nand U341 (N_341,In_1290,In_636);
xor U342 (N_342,In_1459,In_360);
and U343 (N_343,In_29,In_855);
nor U344 (N_344,In_1954,In_1841);
nor U345 (N_345,In_1890,In_742);
and U346 (N_346,In_317,In_1230);
and U347 (N_347,In_1981,In_1179);
or U348 (N_348,In_721,In_421);
nor U349 (N_349,In_1572,In_1796);
nor U350 (N_350,In_414,In_156);
or U351 (N_351,In_671,In_664);
or U352 (N_352,In_933,In_682);
nor U353 (N_353,In_1958,In_703);
or U354 (N_354,In_1113,In_248);
nor U355 (N_355,In_1135,In_1913);
xor U356 (N_356,In_1393,In_1776);
nand U357 (N_357,In_227,In_556);
nand U358 (N_358,In_1382,In_1373);
or U359 (N_359,In_263,In_660);
nor U360 (N_360,In_1274,In_611);
nand U361 (N_361,In_391,In_1770);
nor U362 (N_362,In_251,In_1263);
nor U363 (N_363,In_902,In_710);
nor U364 (N_364,In_332,In_1583);
or U365 (N_365,In_1744,In_369);
nor U366 (N_366,In_930,In_1000);
and U367 (N_367,In_1133,In_1853);
and U368 (N_368,In_1092,In_1620);
nor U369 (N_369,In_83,In_676);
nor U370 (N_370,In_650,In_215);
or U371 (N_371,In_1314,In_1356);
nor U372 (N_372,In_873,In_1508);
and U373 (N_373,In_1582,In_258);
or U374 (N_374,In_785,In_1474);
nand U375 (N_375,In_647,In_202);
nand U376 (N_376,In_1813,In_1107);
or U377 (N_377,In_1994,In_697);
and U378 (N_378,In_1286,In_70);
and U379 (N_379,In_247,In_186);
nor U380 (N_380,In_1467,In_1440);
nand U381 (N_381,In_819,In_870);
nor U382 (N_382,In_1488,In_923);
nor U383 (N_383,In_667,In_455);
or U384 (N_384,In_1324,In_240);
or U385 (N_385,In_399,In_395);
or U386 (N_386,In_1044,In_497);
nor U387 (N_387,In_1338,In_778);
nor U388 (N_388,In_1093,In_1226);
nand U389 (N_389,In_1117,In_484);
and U390 (N_390,In_224,In_205);
nand U391 (N_391,In_1085,In_476);
nand U392 (N_392,In_164,In_1717);
or U393 (N_393,In_163,In_718);
nand U394 (N_394,In_478,In_111);
or U395 (N_395,In_309,In_577);
or U396 (N_396,In_969,In_779);
nand U397 (N_397,In_67,In_1755);
and U398 (N_398,In_1985,In_393);
or U399 (N_399,In_281,In_1749);
or U400 (N_400,In_579,In_897);
and U401 (N_401,In_1471,In_190);
nor U402 (N_402,In_1606,In_706);
and U403 (N_403,In_1158,In_1726);
nor U404 (N_404,In_1172,In_1980);
nand U405 (N_405,In_1915,In_1969);
and U406 (N_406,In_557,In_806);
or U407 (N_407,In_1621,In_1610);
and U408 (N_408,In_1956,In_684);
nand U409 (N_409,In_1410,In_1302);
or U410 (N_410,In_1644,In_640);
and U411 (N_411,In_1810,In_397);
nand U412 (N_412,In_212,In_68);
or U413 (N_413,In_509,In_1280);
nand U414 (N_414,In_454,In_1251);
and U415 (N_415,In_1479,In_1678);
nor U416 (N_416,In_1602,In_1057);
xnor U417 (N_417,In_417,In_1901);
nand U418 (N_418,In_1839,In_270);
or U419 (N_419,In_1851,In_1177);
nand U420 (N_420,In_1162,In_1637);
or U421 (N_421,In_1399,In_467);
nand U422 (N_422,In_1370,In_566);
or U423 (N_423,In_563,In_717);
nor U424 (N_424,In_878,In_1289);
nor U425 (N_425,In_1181,In_1881);
nor U426 (N_426,In_469,In_865);
nand U427 (N_427,In_305,In_1157);
nand U428 (N_428,In_242,In_1589);
nand U429 (N_429,In_725,In_1232);
and U430 (N_430,In_430,In_1242);
or U431 (N_431,In_97,In_1935);
nor U432 (N_432,In_958,In_525);
or U433 (N_433,In_24,In_1270);
nand U434 (N_434,In_1383,In_490);
nor U435 (N_435,In_1902,In_404);
nand U436 (N_436,In_859,In_1529);
nor U437 (N_437,In_1437,In_974);
and U438 (N_438,In_1677,In_221);
nand U439 (N_439,In_480,In_1866);
nand U440 (N_440,In_1328,In_942);
nand U441 (N_441,In_1422,In_468);
and U442 (N_442,In_1660,In_984);
nand U443 (N_443,In_1454,In_919);
and U444 (N_444,In_1306,In_1923);
nand U445 (N_445,In_1468,In_14);
and U446 (N_446,In_1987,In_463);
nand U447 (N_447,In_508,In_32);
or U448 (N_448,In_1240,In_922);
or U449 (N_449,In_1143,In_1395);
or U450 (N_450,In_1174,In_910);
or U451 (N_451,In_1349,In_705);
nor U452 (N_452,In_459,In_1411);
nor U453 (N_453,In_140,In_1404);
or U454 (N_454,In_1163,In_1112);
and U455 (N_455,In_446,In_1990);
and U456 (N_456,In_33,In_1663);
and U457 (N_457,In_1623,In_1342);
or U458 (N_458,In_1283,In_1241);
or U459 (N_459,In_1880,In_1083);
and U460 (N_460,In_66,In_1576);
or U461 (N_461,In_1421,In_255);
nor U462 (N_462,In_688,In_474);
nand U463 (N_463,In_1595,In_918);
or U464 (N_464,In_1947,In_1248);
nand U465 (N_465,In_211,In_905);
and U466 (N_466,In_1926,In_1807);
or U467 (N_467,In_473,In_948);
and U468 (N_468,In_405,In_598);
or U469 (N_469,In_1975,In_699);
or U470 (N_470,In_932,In_833);
xnor U471 (N_471,In_1282,In_1605);
nand U472 (N_472,In_1355,In_1523);
and U473 (N_473,In_1706,In_154);
nand U474 (N_474,In_1821,In_1685);
nand U475 (N_475,In_998,In_487);
and U476 (N_476,In_179,In_505);
nor U477 (N_477,In_60,In_341);
and U478 (N_478,In_1497,In_402);
nor U479 (N_479,In_319,In_1676);
and U480 (N_480,In_1615,In_1514);
or U481 (N_481,In_1672,In_1571);
nand U482 (N_482,In_137,In_516);
nor U483 (N_483,In_273,In_752);
nand U484 (N_484,In_406,In_1127);
nor U485 (N_485,In_290,In_1260);
nor U486 (N_486,In_1693,In_127);
or U487 (N_487,In_1931,In_1275);
nor U488 (N_488,In_973,In_208);
nor U489 (N_489,In_1737,In_1800);
nand U490 (N_490,In_1264,In_1797);
or U491 (N_491,In_971,In_981);
and U492 (N_492,In_1634,In_89);
or U493 (N_493,In_65,In_1374);
nor U494 (N_494,In_1119,In_340);
nor U495 (N_495,In_147,In_180);
or U496 (N_496,In_342,In_716);
or U497 (N_497,In_534,In_1524);
nor U498 (N_498,In_746,In_439);
nand U499 (N_499,In_994,In_321);
or U500 (N_500,In_189,In_776);
nor U501 (N_501,In_1481,In_1458);
nand U502 (N_502,In_549,In_92);
nand U503 (N_503,In_452,In_851);
nand U504 (N_504,In_1757,In_1952);
or U505 (N_505,In_591,In_87);
nor U506 (N_506,In_368,In_1825);
or U507 (N_507,In_875,In_1239);
or U508 (N_508,In_1147,In_1160);
or U509 (N_509,In_1889,In_308);
and U510 (N_510,In_1427,In_1601);
nand U511 (N_511,In_1491,In_1950);
nor U512 (N_512,In_1238,In_362);
nand U513 (N_513,In_380,In_576);
nand U514 (N_514,In_145,In_57);
or U515 (N_515,In_1013,In_1064);
nand U516 (N_516,In_1432,In_1917);
nor U517 (N_517,In_1651,In_1416);
nand U518 (N_518,In_76,In_763);
and U519 (N_519,In_184,In_1789);
nand U520 (N_520,In_1061,In_1124);
nand U521 (N_521,In_1728,In_569);
or U522 (N_522,In_1146,In_1485);
nand U523 (N_523,In_1358,In_1948);
and U524 (N_524,In_37,In_1833);
and U525 (N_525,In_223,In_261);
or U526 (N_526,In_820,In_1325);
nand U527 (N_527,In_681,In_1032);
nand U528 (N_528,In_997,In_1689);
or U529 (N_529,In_1786,In_1456);
and U530 (N_530,In_479,In_612);
and U531 (N_531,In_1398,In_567);
and U532 (N_532,In_663,In_170);
nor U533 (N_533,In_1713,In_738);
and U534 (N_534,In_823,In_325);
and U535 (N_535,In_165,In_796);
and U536 (N_536,In_1297,In_318);
nor U537 (N_537,In_772,In_440);
nand U538 (N_538,In_63,In_1878);
nor U539 (N_539,In_1806,In_1098);
nor U540 (N_540,In_783,In_1622);
nand U541 (N_541,In_1630,In_500);
or U542 (N_542,In_726,In_532);
nand U543 (N_543,In_999,In_100);
and U544 (N_544,In_219,In_284);
and U545 (N_545,In_504,In_434);
nand U546 (N_546,In_595,In_1766);
nand U547 (N_547,In_1236,In_1287);
nor U548 (N_548,In_1109,In_523);
or U549 (N_549,In_1436,In_1996);
and U550 (N_550,In_683,In_659);
or U551 (N_551,In_1259,In_1350);
nor U552 (N_552,In_226,In_1702);
nand U553 (N_553,In_1939,In_115);
or U554 (N_554,In_126,In_648);
or U555 (N_555,In_416,In_735);
or U556 (N_556,In_793,In_1385);
nor U557 (N_557,In_1229,In_1563);
nor U558 (N_558,In_916,In_574);
and U559 (N_559,In_1911,In_1246);
or U560 (N_560,In_1829,In_957);
or U561 (N_561,In_759,In_1675);
nor U562 (N_562,In_327,In_1074);
nor U563 (N_563,In_1308,In_1559);
and U564 (N_564,In_1628,In_1964);
nor U565 (N_565,In_1698,In_1365);
and U566 (N_566,In_1394,In_529);
nor U567 (N_567,In_1614,In_1568);
and U568 (N_568,In_848,In_1025);
and U569 (N_569,In_443,In_1245);
and U570 (N_570,In_110,In_11);
nor U571 (N_571,In_1867,In_1584);
and U572 (N_572,In_1360,In_5);
nor U573 (N_573,In_1301,In_609);
and U574 (N_574,In_62,In_1126);
nor U575 (N_575,In_570,In_743);
or U576 (N_576,In_737,In_911);
nand U577 (N_577,In_304,In_1650);
nor U578 (N_578,In_1362,In_1310);
and U579 (N_579,In_1632,In_1811);
or U580 (N_580,In_453,In_243);
and U581 (N_581,In_1656,In_646);
nor U582 (N_582,In_1243,In_266);
or U583 (N_583,In_657,In_625);
and U584 (N_584,In_330,In_1075);
nor U585 (N_585,In_1080,In_637);
and U586 (N_586,In_1714,In_376);
and U587 (N_587,In_472,In_1277);
and U588 (N_588,In_252,In_59);
and U589 (N_589,In_757,In_936);
nor U590 (N_590,In_275,In_1854);
and U591 (N_591,In_1565,In_36);
and U592 (N_592,In_1940,In_800);
nor U593 (N_593,In_1626,In_1960);
or U594 (N_594,In_1094,In_824);
nor U595 (N_595,In_1101,In_894);
and U596 (N_596,In_1553,In_1125);
nor U597 (N_597,In_357,In_986);
nor U598 (N_598,In_1873,In_27);
nand U599 (N_599,In_1392,In_441);
nand U600 (N_600,In_526,In_538);
and U601 (N_601,In_1219,In_4);
and U602 (N_602,In_185,In_448);
nor U603 (N_603,In_1803,In_86);
or U604 (N_604,In_311,In_853);
or U605 (N_605,In_1772,In_1207);
and U606 (N_606,In_124,In_1201);
nand U607 (N_607,In_961,In_1139);
and U608 (N_608,In_989,In_1887);
and U609 (N_609,In_177,In_1148);
nand U610 (N_610,In_1723,In_1357);
nor U611 (N_611,In_654,In_834);
or U612 (N_612,In_1494,In_840);
nor U613 (N_613,In_233,In_174);
nor U614 (N_614,In_827,In_1412);
nor U615 (N_615,In_812,In_600);
nor U616 (N_616,In_982,In_756);
nand U617 (N_617,In_852,In_883);
and U618 (N_618,In_678,In_1183);
or U619 (N_619,In_183,In_1666);
nand U620 (N_620,In_1414,In_424);
or U621 (N_621,In_583,In_363);
or U622 (N_622,In_949,In_780);
nor U623 (N_623,In_511,In_1379);
and U624 (N_624,In_1916,In_254);
nor U625 (N_625,In_109,In_728);
nor U626 (N_626,In_1216,In_679);
nand U627 (N_627,In_52,In_615);
or U628 (N_628,In_551,In_1218);
and U629 (N_629,In_1564,In_1982);
nand U630 (N_630,In_114,In_1446);
nand U631 (N_631,In_1176,In_1767);
or U632 (N_632,In_1820,In_708);
or U633 (N_633,In_175,In_847);
nor U634 (N_634,In_195,In_1774);
or U635 (N_635,In_1654,In_888);
and U636 (N_636,In_1594,In_857);
and U637 (N_637,In_970,In_801);
and U638 (N_638,In_1447,In_1034);
and U639 (N_639,In_21,In_78);
or U640 (N_640,In_1535,In_952);
or U641 (N_641,In_1779,In_1639);
nor U642 (N_642,In_354,In_1088);
or U643 (N_643,In_731,In_130);
and U644 (N_644,In_1521,In_1760);
nor U645 (N_645,In_1700,In_622);
nand U646 (N_646,In_18,In_1455);
nand U647 (N_647,In_552,In_1200);
or U648 (N_648,In_22,In_1835);
nor U649 (N_649,In_1366,In_1986);
nor U650 (N_650,In_135,In_1850);
nand U651 (N_651,In_1165,In_428);
nand U652 (N_652,In_1460,In_1499);
and U653 (N_653,In_112,In_1884);
nor U654 (N_654,In_884,In_206);
nand U655 (N_655,In_1554,In_1993);
and U656 (N_656,In_1258,In_1505);
and U657 (N_657,In_489,In_1865);
nand U658 (N_658,In_172,In_43);
and U659 (N_659,In_1257,In_444);
and U660 (N_660,In_1705,In_1102);
or U661 (N_661,In_1552,In_282);
or U662 (N_662,In_966,In_907);
or U663 (N_663,In_506,In_1304);
or U664 (N_664,In_1247,In_102);
nor U665 (N_665,In_26,In_1450);
nand U666 (N_666,In_1190,In_519);
or U667 (N_667,In_669,In_1453);
nand U668 (N_668,In_461,In_1153);
nor U669 (N_669,In_1967,In_387);
or U670 (N_670,In_1344,In_528);
nand U671 (N_671,In_1808,In_1871);
or U672 (N_672,In_213,In_407);
or U673 (N_673,In_629,In_1992);
nor U674 (N_674,In_661,In_1557);
and U675 (N_675,In_940,In_814);
or U676 (N_676,In_1244,In_359);
or U677 (N_677,In_531,In_1015);
nand U678 (N_678,In_713,In_849);
or U679 (N_679,In_410,In_161);
or U680 (N_680,In_1983,In_1613);
or U681 (N_681,In_1390,In_1619);
and U682 (N_682,In_665,In_1429);
nand U683 (N_683,In_1895,In_987);
nor U684 (N_684,In_279,In_587);
or U685 (N_685,In_773,In_236);
nor U686 (N_686,In_1965,In_178);
nor U687 (N_687,In_1364,In_1979);
or U688 (N_688,In_711,In_411);
or U689 (N_689,In_401,In_831);
nor U690 (N_690,In_413,In_1330);
nor U691 (N_691,In_1604,In_1168);
or U692 (N_692,In_69,In_1910);
nand U693 (N_693,In_871,In_292);
and U694 (N_694,In_618,In_1864);
or U695 (N_695,In_1802,In_822);
or U696 (N_696,In_1817,In_899);
nand U697 (N_697,In_171,In_39);
nor U698 (N_698,In_1826,In_1443);
or U699 (N_699,In_510,In_1198);
nor U700 (N_700,In_885,In_856);
or U701 (N_701,In_1273,In_1311);
or U702 (N_702,In_249,In_56);
nand U703 (N_703,In_268,In_1086);
nand U704 (N_704,In_1863,In_1528);
and U705 (N_705,In_95,In_1475);
nand U706 (N_706,In_61,In_1281);
nor U707 (N_707,In_1159,In_462);
nand U708 (N_708,In_1140,In_1645);
or U709 (N_709,In_1520,In_815);
nand U710 (N_710,In_1464,In_106);
or U711 (N_711,In_892,In_1154);
and U712 (N_712,In_1542,In_1017);
nand U713 (N_713,In_597,In_1898);
nor U714 (N_714,In_1235,In_231);
and U715 (N_715,In_333,In_1588);
nand U716 (N_716,In_1703,In_1587);
nor U717 (N_717,In_1860,In_388);
nor U718 (N_718,In_1209,In_928);
or U719 (N_719,In_1171,In_1674);
or U720 (N_720,In_501,In_1457);
and U721 (N_721,In_426,In_670);
nor U722 (N_722,In_1189,In_774);
nand U723 (N_723,In_1266,In_1134);
nor U724 (N_724,In_1089,In_1962);
nor U725 (N_725,In_198,In_1035);
or U726 (N_726,In_1043,In_324);
nor U727 (N_727,In_1823,In_1599);
nor U728 (N_728,In_1729,In_1781);
nand U729 (N_729,In_445,In_1191);
nand U730 (N_730,In_6,In_40);
nor U731 (N_731,In_753,In_795);
or U732 (N_732,In_524,In_334);
nor U733 (N_733,In_685,In_791);
nor U734 (N_734,In_1423,In_537);
and U735 (N_735,In_605,In_1742);
nor U736 (N_736,In_390,In_1285);
nand U737 (N_737,In_1541,In_203);
nor U738 (N_738,In_1343,In_666);
or U739 (N_739,In_1868,In_1765);
nand U740 (N_740,In_1818,In_944);
nor U741 (N_741,In_199,In_545);
nand U742 (N_742,In_568,In_1175);
or U743 (N_743,In_1105,In_1144);
or U744 (N_744,In_12,In_1515);
nor U745 (N_745,In_1420,In_804);
nor U746 (N_746,In_876,In_118);
nor U747 (N_747,In_633,In_1731);
or U748 (N_748,In_593,In_1538);
or U749 (N_749,In_935,In_1687);
nor U750 (N_750,In_143,In_1321);
and U751 (N_751,In_1401,In_1327);
or U752 (N_752,In_1657,In_358);
or U753 (N_753,In_1708,In_1469);
nor U754 (N_754,In_187,In_361);
and U755 (N_755,In_1668,In_1734);
nand U756 (N_756,In_1419,In_499);
nand U757 (N_757,In_872,In_1424);
nor U758 (N_758,In_491,In_1452);
or U759 (N_759,In_1777,In_105);
and U760 (N_760,In_1359,In_15);
and U761 (N_761,In_517,In_1451);
nand U762 (N_762,In_1831,In_1347);
or U763 (N_763,In_370,In_869);
nor U764 (N_764,In_1449,In_1517);
nor U765 (N_765,In_1082,In_559);
or U766 (N_766,In_1673,In_610);
and U767 (N_767,In_1988,In_1333);
or U768 (N_768,In_1371,In_1152);
and U769 (N_769,In_786,In_1323);
nand U770 (N_770,In_1196,In_748);
or U771 (N_771,In_1597,In_297);
nand U772 (N_772,In_1223,In_1116);
or U773 (N_773,In_365,In_782);
and U774 (N_774,In_1719,In_225);
or U775 (N_775,In_1516,In_107);
nand U776 (N_776,In_1874,In_245);
nor U777 (N_777,In_1859,In_1531);
and U778 (N_778,In_322,In_1790);
nand U779 (N_779,In_1762,In_1966);
and U780 (N_780,In_1027,In_1608);
or U781 (N_781,In_420,In_864);
or U782 (N_782,In_1699,In_423);
or U783 (N_783,In_818,In_1023);
and U784 (N_784,In_874,In_1114);
or U785 (N_785,In_1843,In_310);
nand U786 (N_786,In_1998,In_854);
or U787 (N_787,In_586,In_1288);
nand U788 (N_788,In_1556,In_1836);
nor U789 (N_789,In_108,In_835);
and U790 (N_790,In_797,In_38);
and U791 (N_791,In_235,In_116);
or U792 (N_792,In_1828,In_1951);
or U793 (N_793,In_502,In_1003);
xor U794 (N_794,In_799,In_513);
nand U795 (N_795,In_1912,In_246);
and U796 (N_796,In_903,In_303);
and U797 (N_797,In_931,In_1840);
or U798 (N_798,In_1256,In_1930);
nand U799 (N_799,In_619,In_260);
nand U800 (N_800,In_632,In_736);
and U801 (N_801,In_1580,In_1794);
or U802 (N_802,In_230,In_956);
and U803 (N_803,In_1184,In_1104);
nor U804 (N_804,In_1971,In_1059);
or U805 (N_805,In_45,In_1896);
nand U806 (N_806,In_1942,In_1759);
nor U807 (N_807,In_1071,In_23);
nand U808 (N_808,In_120,In_1941);
and U809 (N_809,In_1462,In_1030);
and U810 (N_810,In_573,In_1026);
nor U811 (N_811,In_572,In_946);
nand U812 (N_812,In_1773,In_1084);
and U813 (N_813,In_1593,In_562);
or U814 (N_814,In_1512,In_643);
and U815 (N_815,In_1047,In_1943);
and U816 (N_816,In_8,In_229);
nor U817 (N_817,In_1291,In_1053);
nand U818 (N_818,In_85,In_1352);
nor U819 (N_819,In_264,In_343);
or U820 (N_820,In_465,In_1652);
nand U821 (N_821,In_777,In_315);
nor U822 (N_822,In_244,In_162);
nand U823 (N_823,In_113,In_977);
or U824 (N_824,In_1293,In_218);
and U825 (N_825,In_1151,In_542);
or U826 (N_826,In_477,In_13);
nor U827 (N_827,In_1991,In_507);
nor U828 (N_828,In_862,In_755);
nand U829 (N_829,In_924,In_727);
xnor U830 (N_830,In_1764,In_1661);
nor U831 (N_831,In_1496,In_1932);
nor U832 (N_832,In_53,In_767);
or U833 (N_833,In_809,In_157);
nand U834 (N_834,In_152,In_830);
or U835 (N_835,In_604,In_1724);
and U836 (N_836,In_367,In_645);
or U837 (N_837,In_1202,In_1492);
or U838 (N_838,In_1999,In_1712);
nand U839 (N_839,In_621,In_1076);
or U840 (N_840,In_1848,In_1056);
nand U841 (N_841,In_350,In_129);
or U842 (N_842,In_841,In_1511);
and U843 (N_843,In_896,In_1178);
and U844 (N_844,In_729,In_1968);
and U845 (N_845,In_1607,In_1396);
nand U846 (N_846,In_1688,In_1876);
or U847 (N_847,In_937,In_1842);
nand U848 (N_848,In_300,In_1187);
or U849 (N_849,In_720,In_826);
and U850 (N_850,In_496,In_1329);
and U851 (N_851,In_1185,In_1334);
nor U852 (N_852,In_339,In_582);
and U853 (N_853,In_1741,In_301);
nand U854 (N_854,In_449,In_1062);
nor U855 (N_855,In_1970,In_668);
nand U856 (N_856,In_1194,In_348);
nor U857 (N_857,In_808,In_1627);
and U858 (N_858,In_512,In_972);
nand U859 (N_859,In_329,In_1011);
nor U860 (N_860,In_153,In_1022);
or U861 (N_861,In_1197,In_912);
and U862 (N_862,In_1381,In_925);
nor U863 (N_863,In_1768,In_1430);
or U864 (N_864,In_1908,In_470);
nand U865 (N_865,In_788,In_1751);
nor U866 (N_866,In_696,In_1534);
or U867 (N_867,In_1805,In_1166);
or U868 (N_868,In_745,In_601);
and U869 (N_869,In_1500,In_1477);
nor U870 (N_870,In_1221,In_1740);
and U871 (N_871,In_1363,In_535);
nand U872 (N_872,In_1389,In_82);
nand U873 (N_873,In_1847,In_1530);
and U874 (N_874,In_1292,In_1254);
nor U875 (N_875,In_7,In_1046);
nor U876 (N_876,In_1037,In_1106);
nand U877 (N_877,In_1900,In_1341);
nand U878 (N_878,In_1691,In_1795);
or U879 (N_879,In_1428,In_132);
nor U880 (N_880,In_1603,In_1100);
nor U881 (N_881,In_460,In_1195);
nand U882 (N_882,In_1019,In_1299);
nor U883 (N_883,In_1058,In_1199);
nand U884 (N_884,In_349,In_241);
or U885 (N_885,In_1914,In_1856);
or U886 (N_886,In_1193,In_425);
nand U887 (N_887,In_1567,In_1307);
and U888 (N_888,In_1550,In_1073);
and U889 (N_889,In_1036,In_1560);
and U890 (N_890,In_584,In_377);
or U891 (N_891,In_1161,In_151);
nor U892 (N_892,In_1351,In_409);
or U893 (N_893,In_1353,In_1522);
nor U894 (N_894,In_51,In_1403);
nand U895 (N_895,In_366,In_1132);
nor U896 (N_896,In_35,In_1649);
or U897 (N_897,In_1224,In_825);
nand U898 (N_898,In_514,In_31);
nor U899 (N_899,In_702,In_730);
nor U900 (N_900,In_451,In_1721);
nor U901 (N_901,In_1377,In_138);
and U902 (N_902,In_1331,In_766);
and U903 (N_903,In_144,In_904);
and U904 (N_904,In_1380,In_963);
xnor U905 (N_905,In_1487,In_1883);
or U906 (N_906,In_1461,In_1519);
and U907 (N_907,In_561,In_1029);
nor U908 (N_908,In_608,In_1701);
or U909 (N_909,In_250,In_1830);
and U910 (N_910,In_741,In_1339);
nand U911 (N_911,In_1855,In_689);
and U912 (N_912,In_1922,In_1885);
and U913 (N_913,In_283,In_1038);
nand U914 (N_914,In_1526,In_269);
xor U915 (N_915,In_1695,In_1478);
nor U916 (N_916,In_1138,In_954);
or U917 (N_917,In_498,In_1110);
nor U918 (N_918,In_1387,In_1775);
nand U919 (N_919,In_522,In_1303);
nand U920 (N_920,In_1591,In_492);
or U921 (N_921,In_520,In_456);
nor U922 (N_922,In_630,In_133);
or U923 (N_923,In_836,In_842);
nand U924 (N_924,In_1050,In_867);
nand U925 (N_925,In_1131,In_1933);
or U926 (N_926,In_1065,In_740);
nor U927 (N_927,In_1949,In_1336);
nand U928 (N_928,In_719,In_1720);
nor U929 (N_929,In_1819,In_384);
nor U930 (N_930,In_1014,In_1222);
nor U931 (N_931,In_1834,In_1391);
nor U932 (N_932,In_1300,In_1318);
or U933 (N_933,In_1586,In_675);
and U934 (N_934,In_1869,In_695);
or U935 (N_935,In_1903,In_1079);
nand U936 (N_936,In_662,In_381);
or U937 (N_937,In_701,In_71);
nor U938 (N_938,In_953,In_1638);
nor U939 (N_939,In_1827,In_901);
and U940 (N_940,In_288,In_64);
nand U941 (N_941,In_858,In_616);
or U942 (N_942,In_850,In_1070);
nor U943 (N_943,In_541,In_1220);
or U944 (N_944,In_495,In_1128);
and U945 (N_945,In_1372,In_1643);
nor U946 (N_946,In_863,In_1748);
and U947 (N_947,In_1212,In_1388);
xnor U948 (N_948,In_371,In_1575);
and U949 (N_949,In_807,In_320);
nand U950 (N_950,In_1265,In_1431);
and U951 (N_951,In_652,In_838);
and U952 (N_952,In_1137,In_1008);
and U953 (N_953,In_1141,In_1753);
nor U954 (N_954,In_335,In_232);
and U955 (N_955,In_1211,In_758);
and U956 (N_956,In_592,In_438);
nor U957 (N_957,In_639,In_805);
nor U958 (N_958,In_1081,In_383);
nand U959 (N_959,In_464,In_403);
xnor U960 (N_960,In_10,In_34);
or U961 (N_961,In_811,In_351);
xnor U962 (N_962,In_257,In_1743);
and U963 (N_963,In_1052,In_1888);
nor U964 (N_964,In_1090,In_656);
or U965 (N_965,In_191,In_1977);
and U966 (N_966,In_1763,In_631);
nor U967 (N_967,In_382,In_1320);
and U968 (N_968,In_1316,In_299);
or U969 (N_969,In_1861,In_293);
nor U970 (N_970,In_992,In_1758);
nor U971 (N_971,In_1832,In_1715);
nor U972 (N_972,In_1814,In_49);
and U973 (N_973,In_493,In_1972);
nand U974 (N_974,In_1276,In_1262);
nand U975 (N_975,In_1921,In_1852);
or U976 (N_976,In_813,In_1600);
or U977 (N_977,In_182,In_48);
or U978 (N_978,In_1655,In_347);
nand U979 (N_979,In_336,In_1846);
and U980 (N_980,In_747,In_503);
or U981 (N_981,In_1662,In_839);
nand U982 (N_982,In_1213,In_1927);
and U983 (N_983,In_1683,In_104);
and U984 (N_984,In_20,In_475);
and U985 (N_985,In_99,In_1192);
nor U986 (N_986,In_136,In_1054);
and U987 (N_987,In_220,In_1506);
and U988 (N_988,In_1214,In_1647);
nor U989 (N_989,In_1804,In_200);
nor U990 (N_990,In_1857,In_1463);
or U991 (N_991,In_1579,In_1704);
nand U992 (N_992,In_1858,In_546);
or U993 (N_993,In_400,In_1838);
or U994 (N_994,In_1920,In_222);
and U995 (N_995,In_1121,In_58);
nor U996 (N_996,In_1465,In_326);
or U997 (N_997,In_262,In_271);
or U998 (N_998,In_265,In_1928);
nor U999 (N_999,In_1696,In_312);
and U1000 (N_1000,In_193,In_1339);
nor U1001 (N_1001,In_59,In_912);
and U1002 (N_1002,In_1932,In_1533);
or U1003 (N_1003,In_1061,In_1506);
nand U1004 (N_1004,In_1572,In_1732);
nor U1005 (N_1005,In_1659,In_1987);
nand U1006 (N_1006,In_290,In_1670);
and U1007 (N_1007,In_989,In_622);
or U1008 (N_1008,In_4,In_1056);
and U1009 (N_1009,In_393,In_325);
nor U1010 (N_1010,In_572,In_363);
nor U1011 (N_1011,In_1845,In_726);
nand U1012 (N_1012,In_1424,In_214);
or U1013 (N_1013,In_348,In_1859);
nor U1014 (N_1014,In_419,In_1972);
nand U1015 (N_1015,In_1570,In_1610);
nor U1016 (N_1016,In_1311,In_799);
nand U1017 (N_1017,In_1601,In_525);
or U1018 (N_1018,In_375,In_793);
and U1019 (N_1019,In_391,In_1512);
nand U1020 (N_1020,In_1744,In_1948);
and U1021 (N_1021,In_712,In_1257);
nand U1022 (N_1022,In_1505,In_408);
and U1023 (N_1023,In_1567,In_3);
nor U1024 (N_1024,In_128,In_355);
nand U1025 (N_1025,In_1540,In_677);
nor U1026 (N_1026,In_526,In_572);
nor U1027 (N_1027,In_1813,In_1160);
nand U1028 (N_1028,In_552,In_1460);
nor U1029 (N_1029,In_1385,In_1639);
nor U1030 (N_1030,In_457,In_1610);
and U1031 (N_1031,In_648,In_1556);
nor U1032 (N_1032,In_571,In_1780);
and U1033 (N_1033,In_467,In_1258);
and U1034 (N_1034,In_1679,In_875);
and U1035 (N_1035,In_650,In_1075);
or U1036 (N_1036,In_1971,In_283);
or U1037 (N_1037,In_1597,In_1405);
nand U1038 (N_1038,In_1928,In_1399);
and U1039 (N_1039,In_515,In_721);
nand U1040 (N_1040,In_1406,In_1463);
or U1041 (N_1041,In_616,In_129);
nor U1042 (N_1042,In_65,In_319);
and U1043 (N_1043,In_465,In_1499);
nor U1044 (N_1044,In_1319,In_1616);
xor U1045 (N_1045,In_268,In_1747);
nand U1046 (N_1046,In_1078,In_1156);
or U1047 (N_1047,In_1057,In_706);
and U1048 (N_1048,In_1436,In_43);
nand U1049 (N_1049,In_1202,In_1087);
nand U1050 (N_1050,In_1194,In_1187);
nor U1051 (N_1051,In_885,In_729);
nand U1052 (N_1052,In_481,In_687);
and U1053 (N_1053,In_1651,In_997);
nor U1054 (N_1054,In_638,In_926);
or U1055 (N_1055,In_763,In_1164);
or U1056 (N_1056,In_1193,In_32);
or U1057 (N_1057,In_737,In_141);
nor U1058 (N_1058,In_316,In_1185);
xnor U1059 (N_1059,In_1649,In_1719);
or U1060 (N_1060,In_1113,In_354);
nand U1061 (N_1061,In_809,In_873);
nor U1062 (N_1062,In_1988,In_1759);
nor U1063 (N_1063,In_924,In_1518);
and U1064 (N_1064,In_538,In_1858);
and U1065 (N_1065,In_253,In_1187);
nand U1066 (N_1066,In_1982,In_526);
or U1067 (N_1067,In_1086,In_1063);
nand U1068 (N_1068,In_414,In_453);
or U1069 (N_1069,In_137,In_885);
nor U1070 (N_1070,In_1288,In_706);
nand U1071 (N_1071,In_266,In_1596);
and U1072 (N_1072,In_733,In_1062);
and U1073 (N_1073,In_143,In_1031);
or U1074 (N_1074,In_284,In_199);
and U1075 (N_1075,In_1178,In_1480);
or U1076 (N_1076,In_1063,In_1000);
nand U1077 (N_1077,In_561,In_1838);
nor U1078 (N_1078,In_74,In_376);
nor U1079 (N_1079,In_658,In_1370);
and U1080 (N_1080,In_1897,In_762);
nor U1081 (N_1081,In_1709,In_697);
and U1082 (N_1082,In_1952,In_494);
or U1083 (N_1083,In_1728,In_1989);
nand U1084 (N_1084,In_1521,In_873);
nor U1085 (N_1085,In_149,In_1458);
or U1086 (N_1086,In_1763,In_1856);
nor U1087 (N_1087,In_1193,In_1727);
or U1088 (N_1088,In_1587,In_405);
nor U1089 (N_1089,In_1840,In_1334);
nor U1090 (N_1090,In_218,In_369);
nor U1091 (N_1091,In_1406,In_205);
nor U1092 (N_1092,In_1575,In_1492);
or U1093 (N_1093,In_1282,In_882);
and U1094 (N_1094,In_111,In_1810);
nand U1095 (N_1095,In_661,In_1041);
nor U1096 (N_1096,In_1395,In_1190);
or U1097 (N_1097,In_1428,In_225);
and U1098 (N_1098,In_1932,In_1554);
nor U1099 (N_1099,In_1205,In_379);
nand U1100 (N_1100,In_1101,In_533);
and U1101 (N_1101,In_1004,In_312);
or U1102 (N_1102,In_1206,In_384);
nand U1103 (N_1103,In_1162,In_557);
nand U1104 (N_1104,In_771,In_1778);
or U1105 (N_1105,In_505,In_209);
and U1106 (N_1106,In_1126,In_1124);
xnor U1107 (N_1107,In_1733,In_1952);
nand U1108 (N_1108,In_975,In_1475);
nor U1109 (N_1109,In_1495,In_1890);
nand U1110 (N_1110,In_1168,In_262);
nor U1111 (N_1111,In_753,In_1241);
nor U1112 (N_1112,In_1644,In_40);
nand U1113 (N_1113,In_489,In_1028);
or U1114 (N_1114,In_1748,In_1425);
nand U1115 (N_1115,In_39,In_634);
or U1116 (N_1116,In_927,In_762);
nor U1117 (N_1117,In_815,In_914);
xnor U1118 (N_1118,In_1915,In_1125);
nor U1119 (N_1119,In_1138,In_307);
or U1120 (N_1120,In_159,In_1431);
nor U1121 (N_1121,In_518,In_1696);
nor U1122 (N_1122,In_1671,In_669);
nor U1123 (N_1123,In_103,In_920);
nand U1124 (N_1124,In_1987,In_858);
nor U1125 (N_1125,In_842,In_749);
nand U1126 (N_1126,In_420,In_1242);
nor U1127 (N_1127,In_1535,In_350);
nand U1128 (N_1128,In_445,In_748);
nand U1129 (N_1129,In_920,In_518);
nor U1130 (N_1130,In_1588,In_709);
and U1131 (N_1131,In_1404,In_327);
nor U1132 (N_1132,In_1841,In_1980);
and U1133 (N_1133,In_61,In_1711);
nor U1134 (N_1134,In_1395,In_1459);
or U1135 (N_1135,In_1367,In_706);
nor U1136 (N_1136,In_46,In_1135);
nand U1137 (N_1137,In_869,In_576);
nand U1138 (N_1138,In_189,In_1562);
or U1139 (N_1139,In_1634,In_1826);
and U1140 (N_1140,In_999,In_1663);
and U1141 (N_1141,In_1940,In_942);
nor U1142 (N_1142,In_370,In_1983);
nand U1143 (N_1143,In_1542,In_969);
nand U1144 (N_1144,In_562,In_1328);
or U1145 (N_1145,In_1250,In_1158);
nor U1146 (N_1146,In_1636,In_903);
and U1147 (N_1147,In_69,In_411);
nand U1148 (N_1148,In_1641,In_1245);
and U1149 (N_1149,In_1070,In_825);
nand U1150 (N_1150,In_432,In_1890);
nand U1151 (N_1151,In_189,In_921);
and U1152 (N_1152,In_311,In_1207);
nor U1153 (N_1153,In_769,In_1900);
or U1154 (N_1154,In_1373,In_384);
or U1155 (N_1155,In_131,In_549);
nand U1156 (N_1156,In_1953,In_1711);
or U1157 (N_1157,In_1453,In_837);
nor U1158 (N_1158,In_739,In_1631);
or U1159 (N_1159,In_672,In_1234);
and U1160 (N_1160,In_878,In_393);
nand U1161 (N_1161,In_1230,In_19);
or U1162 (N_1162,In_1728,In_620);
nor U1163 (N_1163,In_570,In_1704);
nand U1164 (N_1164,In_1343,In_330);
nor U1165 (N_1165,In_534,In_191);
xor U1166 (N_1166,In_794,In_1443);
nand U1167 (N_1167,In_1030,In_1958);
nand U1168 (N_1168,In_767,In_400);
nand U1169 (N_1169,In_1770,In_1768);
nor U1170 (N_1170,In_888,In_1897);
nand U1171 (N_1171,In_1895,In_1702);
and U1172 (N_1172,In_998,In_1609);
nor U1173 (N_1173,In_298,In_1984);
nand U1174 (N_1174,In_1984,In_997);
nand U1175 (N_1175,In_770,In_188);
nand U1176 (N_1176,In_269,In_584);
and U1177 (N_1177,In_593,In_1614);
or U1178 (N_1178,In_765,In_1753);
nor U1179 (N_1179,In_1903,In_67);
and U1180 (N_1180,In_491,In_1744);
nor U1181 (N_1181,In_1510,In_849);
and U1182 (N_1182,In_618,In_136);
nand U1183 (N_1183,In_662,In_403);
nand U1184 (N_1184,In_1366,In_45);
or U1185 (N_1185,In_1705,In_1396);
and U1186 (N_1186,In_145,In_1494);
or U1187 (N_1187,In_939,In_1341);
or U1188 (N_1188,In_1038,In_1476);
and U1189 (N_1189,In_218,In_1809);
and U1190 (N_1190,In_1426,In_1765);
nand U1191 (N_1191,In_1756,In_644);
and U1192 (N_1192,In_1982,In_452);
nor U1193 (N_1193,In_1677,In_1580);
and U1194 (N_1194,In_852,In_1136);
or U1195 (N_1195,In_1542,In_963);
nor U1196 (N_1196,In_1592,In_1663);
or U1197 (N_1197,In_1061,In_1089);
and U1198 (N_1198,In_189,In_1783);
xnor U1199 (N_1199,In_181,In_1121);
or U1200 (N_1200,In_1803,In_1615);
or U1201 (N_1201,In_710,In_742);
and U1202 (N_1202,In_581,In_1678);
and U1203 (N_1203,In_949,In_1189);
nand U1204 (N_1204,In_77,In_1249);
nor U1205 (N_1205,In_1220,In_219);
nand U1206 (N_1206,In_1361,In_628);
and U1207 (N_1207,In_1420,In_1133);
nor U1208 (N_1208,In_538,In_1247);
or U1209 (N_1209,In_1611,In_1627);
and U1210 (N_1210,In_636,In_827);
and U1211 (N_1211,In_1795,In_1675);
nand U1212 (N_1212,In_584,In_149);
or U1213 (N_1213,In_1488,In_1880);
nand U1214 (N_1214,In_871,In_1845);
nand U1215 (N_1215,In_830,In_1803);
or U1216 (N_1216,In_1648,In_1904);
nor U1217 (N_1217,In_941,In_1290);
or U1218 (N_1218,In_467,In_1133);
nor U1219 (N_1219,In_1853,In_1062);
or U1220 (N_1220,In_73,In_60);
or U1221 (N_1221,In_1199,In_488);
nor U1222 (N_1222,In_1662,In_911);
and U1223 (N_1223,In_1617,In_12);
nand U1224 (N_1224,In_950,In_1281);
nor U1225 (N_1225,In_272,In_154);
nor U1226 (N_1226,In_760,In_90);
nor U1227 (N_1227,In_1865,In_1963);
nor U1228 (N_1228,In_131,In_1647);
or U1229 (N_1229,In_103,In_944);
nor U1230 (N_1230,In_434,In_1674);
nand U1231 (N_1231,In_1977,In_833);
and U1232 (N_1232,In_592,In_1461);
nor U1233 (N_1233,In_1818,In_1274);
nand U1234 (N_1234,In_742,In_546);
nor U1235 (N_1235,In_1417,In_1248);
nor U1236 (N_1236,In_136,In_1731);
or U1237 (N_1237,In_1731,In_665);
nor U1238 (N_1238,In_733,In_1822);
nand U1239 (N_1239,In_339,In_1846);
nor U1240 (N_1240,In_464,In_153);
or U1241 (N_1241,In_871,In_986);
or U1242 (N_1242,In_1469,In_1400);
xnor U1243 (N_1243,In_371,In_117);
nand U1244 (N_1244,In_536,In_1875);
nand U1245 (N_1245,In_305,In_411);
nand U1246 (N_1246,In_615,In_966);
nand U1247 (N_1247,In_125,In_177);
nor U1248 (N_1248,In_109,In_1323);
nand U1249 (N_1249,In_38,In_553);
or U1250 (N_1250,In_311,In_851);
or U1251 (N_1251,In_153,In_162);
or U1252 (N_1252,In_718,In_236);
and U1253 (N_1253,In_330,In_1065);
nand U1254 (N_1254,In_1062,In_336);
and U1255 (N_1255,In_1936,In_1807);
nor U1256 (N_1256,In_1718,In_1701);
nor U1257 (N_1257,In_532,In_381);
nor U1258 (N_1258,In_72,In_846);
and U1259 (N_1259,In_930,In_477);
nand U1260 (N_1260,In_327,In_1449);
or U1261 (N_1261,In_1200,In_1583);
nand U1262 (N_1262,In_958,In_670);
nor U1263 (N_1263,In_12,In_1454);
nor U1264 (N_1264,In_876,In_742);
or U1265 (N_1265,In_250,In_843);
nor U1266 (N_1266,In_1083,In_1259);
nor U1267 (N_1267,In_549,In_343);
nor U1268 (N_1268,In_1137,In_1282);
nor U1269 (N_1269,In_525,In_834);
nor U1270 (N_1270,In_1934,In_469);
nand U1271 (N_1271,In_249,In_1698);
and U1272 (N_1272,In_799,In_234);
or U1273 (N_1273,In_444,In_642);
nor U1274 (N_1274,In_698,In_561);
and U1275 (N_1275,In_895,In_1462);
or U1276 (N_1276,In_408,In_803);
nor U1277 (N_1277,In_1493,In_368);
xnor U1278 (N_1278,In_1090,In_1915);
nand U1279 (N_1279,In_101,In_325);
or U1280 (N_1280,In_393,In_1937);
or U1281 (N_1281,In_59,In_1281);
or U1282 (N_1282,In_1333,In_96);
nand U1283 (N_1283,In_1010,In_1660);
nand U1284 (N_1284,In_865,In_165);
and U1285 (N_1285,In_1084,In_853);
and U1286 (N_1286,In_1157,In_1842);
nor U1287 (N_1287,In_1215,In_1071);
nor U1288 (N_1288,In_410,In_63);
or U1289 (N_1289,In_670,In_1528);
and U1290 (N_1290,In_1856,In_693);
or U1291 (N_1291,In_1356,In_1395);
nand U1292 (N_1292,In_1608,In_1156);
nor U1293 (N_1293,In_400,In_615);
nand U1294 (N_1294,In_512,In_1722);
and U1295 (N_1295,In_1670,In_740);
nor U1296 (N_1296,In_1014,In_435);
nor U1297 (N_1297,In_348,In_1962);
nand U1298 (N_1298,In_301,In_1830);
or U1299 (N_1299,In_1205,In_1843);
or U1300 (N_1300,In_1669,In_662);
or U1301 (N_1301,In_178,In_1568);
or U1302 (N_1302,In_1005,In_1057);
nor U1303 (N_1303,In_918,In_630);
or U1304 (N_1304,In_357,In_1279);
and U1305 (N_1305,In_1436,In_1054);
nor U1306 (N_1306,In_116,In_1330);
and U1307 (N_1307,In_1590,In_1536);
nor U1308 (N_1308,In_357,In_1775);
and U1309 (N_1309,In_1719,In_1690);
and U1310 (N_1310,In_1051,In_1185);
nor U1311 (N_1311,In_1222,In_1497);
nand U1312 (N_1312,In_1768,In_262);
and U1313 (N_1313,In_1047,In_256);
nor U1314 (N_1314,In_427,In_108);
nor U1315 (N_1315,In_1696,In_1811);
or U1316 (N_1316,In_1810,In_991);
or U1317 (N_1317,In_101,In_267);
or U1318 (N_1318,In_1850,In_11);
nor U1319 (N_1319,In_1374,In_1617);
nor U1320 (N_1320,In_752,In_915);
nor U1321 (N_1321,In_1079,In_229);
and U1322 (N_1322,In_190,In_443);
nor U1323 (N_1323,In_252,In_615);
and U1324 (N_1324,In_1621,In_1177);
nand U1325 (N_1325,In_514,In_114);
nand U1326 (N_1326,In_476,In_717);
and U1327 (N_1327,In_486,In_745);
nor U1328 (N_1328,In_1506,In_1873);
and U1329 (N_1329,In_1013,In_1119);
nor U1330 (N_1330,In_1023,In_1625);
nand U1331 (N_1331,In_586,In_1387);
or U1332 (N_1332,In_1249,In_189);
or U1333 (N_1333,In_1844,In_49);
nand U1334 (N_1334,In_1458,In_54);
nand U1335 (N_1335,In_1995,In_887);
or U1336 (N_1336,In_30,In_184);
nand U1337 (N_1337,In_59,In_1795);
nor U1338 (N_1338,In_1588,In_977);
nand U1339 (N_1339,In_341,In_1315);
or U1340 (N_1340,In_599,In_697);
nor U1341 (N_1341,In_1859,In_969);
and U1342 (N_1342,In_1917,In_1719);
and U1343 (N_1343,In_476,In_609);
nor U1344 (N_1344,In_833,In_98);
and U1345 (N_1345,In_334,In_1746);
or U1346 (N_1346,In_73,In_1373);
nand U1347 (N_1347,In_15,In_887);
or U1348 (N_1348,In_1133,In_1180);
nand U1349 (N_1349,In_950,In_1451);
or U1350 (N_1350,In_1928,In_1292);
nand U1351 (N_1351,In_195,In_1271);
xnor U1352 (N_1352,In_797,In_427);
nor U1353 (N_1353,In_1711,In_1452);
nor U1354 (N_1354,In_1090,In_94);
and U1355 (N_1355,In_974,In_1593);
and U1356 (N_1356,In_920,In_1789);
nand U1357 (N_1357,In_767,In_60);
xnor U1358 (N_1358,In_6,In_66);
nand U1359 (N_1359,In_489,In_1383);
and U1360 (N_1360,In_1790,In_1631);
nor U1361 (N_1361,In_1619,In_219);
and U1362 (N_1362,In_727,In_820);
nor U1363 (N_1363,In_1777,In_383);
or U1364 (N_1364,In_633,In_2);
nor U1365 (N_1365,In_1526,In_1107);
and U1366 (N_1366,In_1001,In_423);
nor U1367 (N_1367,In_381,In_1370);
and U1368 (N_1368,In_534,In_1982);
or U1369 (N_1369,In_1079,In_1789);
and U1370 (N_1370,In_1904,In_1189);
and U1371 (N_1371,In_39,In_413);
nand U1372 (N_1372,In_1935,In_786);
and U1373 (N_1373,In_381,In_453);
nand U1374 (N_1374,In_492,In_944);
nor U1375 (N_1375,In_1678,In_1993);
or U1376 (N_1376,In_1694,In_1519);
or U1377 (N_1377,In_910,In_1179);
nand U1378 (N_1378,In_1393,In_272);
and U1379 (N_1379,In_1864,In_1381);
or U1380 (N_1380,In_518,In_1272);
and U1381 (N_1381,In_1770,In_601);
nor U1382 (N_1382,In_1177,In_129);
nor U1383 (N_1383,In_258,In_639);
nor U1384 (N_1384,In_1947,In_1451);
nand U1385 (N_1385,In_1945,In_1694);
nand U1386 (N_1386,In_1101,In_1477);
nand U1387 (N_1387,In_1703,In_475);
nand U1388 (N_1388,In_22,In_1888);
nand U1389 (N_1389,In_599,In_1858);
or U1390 (N_1390,In_1538,In_573);
and U1391 (N_1391,In_1967,In_383);
nand U1392 (N_1392,In_66,In_1843);
or U1393 (N_1393,In_1620,In_1582);
nand U1394 (N_1394,In_618,In_763);
nor U1395 (N_1395,In_1114,In_171);
nor U1396 (N_1396,In_1534,In_703);
and U1397 (N_1397,In_1714,In_523);
nor U1398 (N_1398,In_851,In_1830);
and U1399 (N_1399,In_1039,In_438);
and U1400 (N_1400,In_570,In_103);
nand U1401 (N_1401,In_1591,In_1837);
nor U1402 (N_1402,In_1118,In_595);
and U1403 (N_1403,In_904,In_716);
or U1404 (N_1404,In_571,In_773);
or U1405 (N_1405,In_783,In_1127);
nor U1406 (N_1406,In_1743,In_531);
nand U1407 (N_1407,In_1716,In_1511);
nand U1408 (N_1408,In_556,In_1201);
nand U1409 (N_1409,In_1461,In_262);
and U1410 (N_1410,In_1759,In_1813);
or U1411 (N_1411,In_1633,In_1696);
or U1412 (N_1412,In_1822,In_1156);
nand U1413 (N_1413,In_869,In_398);
or U1414 (N_1414,In_649,In_796);
nor U1415 (N_1415,In_612,In_1161);
nor U1416 (N_1416,In_703,In_368);
xor U1417 (N_1417,In_549,In_1469);
or U1418 (N_1418,In_1626,In_1484);
and U1419 (N_1419,In_341,In_162);
and U1420 (N_1420,In_685,In_247);
and U1421 (N_1421,In_880,In_1693);
and U1422 (N_1422,In_545,In_756);
nor U1423 (N_1423,In_1471,In_13);
and U1424 (N_1424,In_876,In_1562);
nand U1425 (N_1425,In_1808,In_322);
and U1426 (N_1426,In_596,In_560);
or U1427 (N_1427,In_1110,In_711);
or U1428 (N_1428,In_353,In_1803);
or U1429 (N_1429,In_947,In_1375);
nor U1430 (N_1430,In_840,In_1378);
nand U1431 (N_1431,In_979,In_418);
nor U1432 (N_1432,In_1981,In_865);
nand U1433 (N_1433,In_1919,In_1958);
nor U1434 (N_1434,In_669,In_382);
or U1435 (N_1435,In_598,In_139);
and U1436 (N_1436,In_1447,In_1625);
and U1437 (N_1437,In_1178,In_577);
nand U1438 (N_1438,In_471,In_984);
or U1439 (N_1439,In_1563,In_1920);
nand U1440 (N_1440,In_139,In_1540);
or U1441 (N_1441,In_398,In_761);
or U1442 (N_1442,In_1619,In_864);
nand U1443 (N_1443,In_1135,In_621);
nand U1444 (N_1444,In_761,In_1688);
or U1445 (N_1445,In_1358,In_1341);
nand U1446 (N_1446,In_76,In_1451);
nor U1447 (N_1447,In_1392,In_1291);
or U1448 (N_1448,In_694,In_1747);
nand U1449 (N_1449,In_1120,In_92);
and U1450 (N_1450,In_150,In_1460);
nor U1451 (N_1451,In_1981,In_1309);
and U1452 (N_1452,In_1176,In_1334);
nand U1453 (N_1453,In_1876,In_14);
nand U1454 (N_1454,In_764,In_1188);
nand U1455 (N_1455,In_373,In_1225);
nand U1456 (N_1456,In_605,In_1271);
nor U1457 (N_1457,In_729,In_1643);
and U1458 (N_1458,In_1011,In_1560);
nand U1459 (N_1459,In_1583,In_1329);
and U1460 (N_1460,In_1860,In_1598);
nand U1461 (N_1461,In_317,In_57);
and U1462 (N_1462,In_288,In_1117);
and U1463 (N_1463,In_1323,In_1229);
nand U1464 (N_1464,In_848,In_1491);
nand U1465 (N_1465,In_147,In_1034);
and U1466 (N_1466,In_1630,In_1167);
nand U1467 (N_1467,In_1195,In_351);
and U1468 (N_1468,In_1948,In_1837);
nand U1469 (N_1469,In_1028,In_1542);
nor U1470 (N_1470,In_1313,In_742);
and U1471 (N_1471,In_1089,In_1440);
nand U1472 (N_1472,In_925,In_1325);
nand U1473 (N_1473,In_1735,In_592);
nand U1474 (N_1474,In_1236,In_628);
and U1475 (N_1475,In_1022,In_784);
xnor U1476 (N_1476,In_138,In_706);
nor U1477 (N_1477,In_1916,In_1330);
or U1478 (N_1478,In_146,In_419);
or U1479 (N_1479,In_675,In_498);
nor U1480 (N_1480,In_1218,In_1685);
or U1481 (N_1481,In_1472,In_862);
nand U1482 (N_1482,In_1258,In_731);
and U1483 (N_1483,In_832,In_359);
or U1484 (N_1484,In_1656,In_1232);
nand U1485 (N_1485,In_32,In_376);
nor U1486 (N_1486,In_986,In_1192);
nand U1487 (N_1487,In_209,In_1136);
nor U1488 (N_1488,In_1569,In_1619);
nor U1489 (N_1489,In_1663,In_763);
nand U1490 (N_1490,In_1194,In_457);
xnor U1491 (N_1491,In_1488,In_695);
or U1492 (N_1492,In_849,In_1063);
nand U1493 (N_1493,In_1083,In_1227);
nor U1494 (N_1494,In_1987,In_58);
nand U1495 (N_1495,In_1747,In_1836);
nor U1496 (N_1496,In_1960,In_1596);
and U1497 (N_1497,In_1020,In_1632);
nand U1498 (N_1498,In_1188,In_1791);
nor U1499 (N_1499,In_1794,In_1934);
nor U1500 (N_1500,In_535,In_1819);
and U1501 (N_1501,In_407,In_944);
nor U1502 (N_1502,In_1324,In_896);
and U1503 (N_1503,In_1436,In_1771);
and U1504 (N_1504,In_14,In_936);
nor U1505 (N_1505,In_972,In_1891);
nand U1506 (N_1506,In_52,In_67);
nor U1507 (N_1507,In_229,In_781);
nor U1508 (N_1508,In_94,In_280);
or U1509 (N_1509,In_16,In_293);
and U1510 (N_1510,In_5,In_1212);
or U1511 (N_1511,In_76,In_130);
or U1512 (N_1512,In_792,In_1532);
or U1513 (N_1513,In_1973,In_25);
nor U1514 (N_1514,In_1532,In_932);
and U1515 (N_1515,In_1541,In_1569);
and U1516 (N_1516,In_1299,In_1021);
nor U1517 (N_1517,In_1181,In_974);
nand U1518 (N_1518,In_1604,In_1753);
nor U1519 (N_1519,In_45,In_1866);
nor U1520 (N_1520,In_737,In_373);
or U1521 (N_1521,In_1336,In_1357);
nor U1522 (N_1522,In_1834,In_430);
or U1523 (N_1523,In_353,In_1215);
nand U1524 (N_1524,In_506,In_1167);
and U1525 (N_1525,In_980,In_304);
or U1526 (N_1526,In_1416,In_1198);
nor U1527 (N_1527,In_1840,In_1509);
or U1528 (N_1528,In_1740,In_369);
nor U1529 (N_1529,In_1505,In_404);
nor U1530 (N_1530,In_1754,In_520);
nor U1531 (N_1531,In_6,In_760);
nand U1532 (N_1532,In_196,In_843);
nor U1533 (N_1533,In_375,In_699);
nor U1534 (N_1534,In_655,In_852);
and U1535 (N_1535,In_685,In_138);
or U1536 (N_1536,In_1195,In_122);
nand U1537 (N_1537,In_1148,In_1918);
or U1538 (N_1538,In_216,In_1305);
or U1539 (N_1539,In_1701,In_479);
nand U1540 (N_1540,In_1380,In_1738);
nor U1541 (N_1541,In_1260,In_1781);
nor U1542 (N_1542,In_1551,In_1269);
nor U1543 (N_1543,In_191,In_535);
and U1544 (N_1544,In_930,In_588);
and U1545 (N_1545,In_1308,In_1349);
or U1546 (N_1546,In_1641,In_1162);
nor U1547 (N_1547,In_647,In_943);
or U1548 (N_1548,In_835,In_1790);
nor U1549 (N_1549,In_14,In_1233);
and U1550 (N_1550,In_550,In_1805);
and U1551 (N_1551,In_1463,In_263);
and U1552 (N_1552,In_606,In_1342);
nor U1553 (N_1553,In_1387,In_658);
and U1554 (N_1554,In_1792,In_3);
or U1555 (N_1555,In_216,In_536);
nor U1556 (N_1556,In_996,In_1289);
nand U1557 (N_1557,In_1482,In_395);
and U1558 (N_1558,In_1814,In_1360);
and U1559 (N_1559,In_969,In_1788);
nor U1560 (N_1560,In_1449,In_1837);
or U1561 (N_1561,In_584,In_650);
and U1562 (N_1562,In_703,In_1549);
nor U1563 (N_1563,In_114,In_459);
nand U1564 (N_1564,In_1375,In_125);
nor U1565 (N_1565,In_1626,In_1986);
or U1566 (N_1566,In_1547,In_42);
and U1567 (N_1567,In_999,In_1514);
xor U1568 (N_1568,In_963,In_281);
nor U1569 (N_1569,In_1432,In_1474);
and U1570 (N_1570,In_54,In_1682);
and U1571 (N_1571,In_307,In_1859);
nand U1572 (N_1572,In_354,In_538);
nor U1573 (N_1573,In_30,In_63);
nand U1574 (N_1574,In_1292,In_549);
or U1575 (N_1575,In_606,In_1217);
nand U1576 (N_1576,In_1656,In_716);
and U1577 (N_1577,In_1605,In_489);
nand U1578 (N_1578,In_1561,In_293);
or U1579 (N_1579,In_407,In_374);
and U1580 (N_1580,In_1660,In_57);
nor U1581 (N_1581,In_623,In_1605);
nor U1582 (N_1582,In_1112,In_1034);
nor U1583 (N_1583,In_280,In_1313);
or U1584 (N_1584,In_1672,In_401);
nand U1585 (N_1585,In_1010,In_1663);
nand U1586 (N_1586,In_960,In_500);
nor U1587 (N_1587,In_674,In_1365);
nor U1588 (N_1588,In_1567,In_1802);
nor U1589 (N_1589,In_74,In_367);
or U1590 (N_1590,In_1270,In_1768);
nand U1591 (N_1591,In_907,In_369);
nor U1592 (N_1592,In_1516,In_724);
or U1593 (N_1593,In_1627,In_1087);
and U1594 (N_1594,In_382,In_1240);
and U1595 (N_1595,In_1693,In_1151);
nand U1596 (N_1596,In_111,In_863);
nand U1597 (N_1597,In_1408,In_570);
nand U1598 (N_1598,In_270,In_951);
nand U1599 (N_1599,In_1597,In_1021);
and U1600 (N_1600,In_506,In_351);
nor U1601 (N_1601,In_1337,In_564);
nand U1602 (N_1602,In_1746,In_309);
or U1603 (N_1603,In_713,In_1471);
nor U1604 (N_1604,In_246,In_589);
nand U1605 (N_1605,In_130,In_1203);
and U1606 (N_1606,In_785,In_983);
nor U1607 (N_1607,In_1096,In_1477);
or U1608 (N_1608,In_252,In_1889);
and U1609 (N_1609,In_1183,In_1663);
and U1610 (N_1610,In_321,In_1543);
nor U1611 (N_1611,In_1391,In_1985);
nand U1612 (N_1612,In_562,In_68);
nand U1613 (N_1613,In_1072,In_1989);
or U1614 (N_1614,In_1938,In_1863);
nor U1615 (N_1615,In_202,In_203);
and U1616 (N_1616,In_1125,In_83);
nor U1617 (N_1617,In_1110,In_1132);
nand U1618 (N_1618,In_649,In_584);
nand U1619 (N_1619,In_735,In_967);
nand U1620 (N_1620,In_662,In_1760);
nand U1621 (N_1621,In_1624,In_1562);
nand U1622 (N_1622,In_874,In_1233);
nor U1623 (N_1623,In_658,In_1105);
or U1624 (N_1624,In_1806,In_60);
or U1625 (N_1625,In_1980,In_131);
nor U1626 (N_1626,In_1352,In_1694);
nor U1627 (N_1627,In_747,In_1758);
nor U1628 (N_1628,In_306,In_98);
nand U1629 (N_1629,In_1415,In_219);
nand U1630 (N_1630,In_1618,In_1669);
nor U1631 (N_1631,In_1228,In_177);
and U1632 (N_1632,In_873,In_1983);
nand U1633 (N_1633,In_1076,In_1498);
and U1634 (N_1634,In_730,In_996);
nor U1635 (N_1635,In_1812,In_1434);
and U1636 (N_1636,In_1661,In_1070);
nor U1637 (N_1637,In_976,In_288);
nor U1638 (N_1638,In_409,In_1300);
nand U1639 (N_1639,In_1929,In_270);
and U1640 (N_1640,In_412,In_524);
nor U1641 (N_1641,In_1892,In_1413);
or U1642 (N_1642,In_771,In_1627);
and U1643 (N_1643,In_1556,In_165);
nor U1644 (N_1644,In_174,In_1034);
nand U1645 (N_1645,In_1324,In_1439);
nor U1646 (N_1646,In_293,In_1856);
and U1647 (N_1647,In_1774,In_637);
and U1648 (N_1648,In_1837,In_1592);
or U1649 (N_1649,In_1801,In_1965);
nand U1650 (N_1650,In_189,In_71);
nand U1651 (N_1651,In_930,In_236);
and U1652 (N_1652,In_398,In_299);
nand U1653 (N_1653,In_1673,In_1244);
nand U1654 (N_1654,In_912,In_1644);
nand U1655 (N_1655,In_1938,In_1239);
nor U1656 (N_1656,In_1438,In_762);
nor U1657 (N_1657,In_1388,In_853);
and U1658 (N_1658,In_1934,In_1372);
nand U1659 (N_1659,In_1337,In_529);
and U1660 (N_1660,In_1116,In_944);
nand U1661 (N_1661,In_1341,In_647);
and U1662 (N_1662,In_434,In_664);
or U1663 (N_1663,In_687,In_865);
nor U1664 (N_1664,In_357,In_1553);
nor U1665 (N_1665,In_848,In_1857);
nand U1666 (N_1666,In_486,In_300);
and U1667 (N_1667,In_1847,In_434);
nand U1668 (N_1668,In_15,In_1341);
nand U1669 (N_1669,In_1362,In_912);
or U1670 (N_1670,In_101,In_399);
nand U1671 (N_1671,In_825,In_1460);
and U1672 (N_1672,In_1168,In_227);
or U1673 (N_1673,In_1768,In_721);
or U1674 (N_1674,In_286,In_89);
xor U1675 (N_1675,In_1453,In_1958);
nand U1676 (N_1676,In_1305,In_769);
nand U1677 (N_1677,In_1705,In_1281);
nand U1678 (N_1678,In_1478,In_1128);
and U1679 (N_1679,In_1167,In_1670);
nor U1680 (N_1680,In_266,In_1498);
nand U1681 (N_1681,In_1820,In_1490);
nor U1682 (N_1682,In_1789,In_683);
nand U1683 (N_1683,In_298,In_1498);
xnor U1684 (N_1684,In_537,In_720);
nor U1685 (N_1685,In_1585,In_1248);
nand U1686 (N_1686,In_870,In_1105);
nand U1687 (N_1687,In_465,In_1870);
nand U1688 (N_1688,In_756,In_1966);
and U1689 (N_1689,In_1841,In_1648);
nand U1690 (N_1690,In_1795,In_590);
nor U1691 (N_1691,In_316,In_1131);
or U1692 (N_1692,In_982,In_1813);
nand U1693 (N_1693,In_892,In_487);
nand U1694 (N_1694,In_1024,In_122);
nand U1695 (N_1695,In_1405,In_1610);
nor U1696 (N_1696,In_1695,In_1148);
and U1697 (N_1697,In_1930,In_1807);
nor U1698 (N_1698,In_1489,In_1096);
nand U1699 (N_1699,In_1365,In_1443);
and U1700 (N_1700,In_1663,In_1433);
nor U1701 (N_1701,In_822,In_719);
or U1702 (N_1702,In_1486,In_676);
and U1703 (N_1703,In_1067,In_1411);
nor U1704 (N_1704,In_1952,In_1443);
nor U1705 (N_1705,In_920,In_1578);
nor U1706 (N_1706,In_753,In_773);
nor U1707 (N_1707,In_1168,In_671);
or U1708 (N_1708,In_703,In_1722);
nor U1709 (N_1709,In_1036,In_831);
or U1710 (N_1710,In_297,In_1445);
nor U1711 (N_1711,In_1566,In_233);
nand U1712 (N_1712,In_728,In_801);
and U1713 (N_1713,In_889,In_808);
or U1714 (N_1714,In_1625,In_902);
nand U1715 (N_1715,In_269,In_295);
nand U1716 (N_1716,In_1607,In_1503);
nand U1717 (N_1717,In_302,In_733);
nor U1718 (N_1718,In_717,In_1546);
nand U1719 (N_1719,In_377,In_259);
nand U1720 (N_1720,In_1407,In_1649);
or U1721 (N_1721,In_699,In_1858);
and U1722 (N_1722,In_1498,In_1816);
nor U1723 (N_1723,In_1242,In_1134);
nand U1724 (N_1724,In_775,In_1566);
and U1725 (N_1725,In_661,In_1668);
or U1726 (N_1726,In_1322,In_196);
nor U1727 (N_1727,In_846,In_88);
or U1728 (N_1728,In_615,In_1766);
nor U1729 (N_1729,In_693,In_605);
and U1730 (N_1730,In_908,In_1868);
and U1731 (N_1731,In_1334,In_385);
and U1732 (N_1732,In_490,In_805);
nor U1733 (N_1733,In_1879,In_1703);
nand U1734 (N_1734,In_1706,In_483);
nor U1735 (N_1735,In_137,In_1360);
and U1736 (N_1736,In_1373,In_1866);
nand U1737 (N_1737,In_1710,In_981);
or U1738 (N_1738,In_1092,In_1961);
nor U1739 (N_1739,In_237,In_1762);
nor U1740 (N_1740,In_178,In_927);
and U1741 (N_1741,In_1017,In_623);
nor U1742 (N_1742,In_1919,In_516);
or U1743 (N_1743,In_687,In_82);
and U1744 (N_1744,In_432,In_1586);
nor U1745 (N_1745,In_1734,In_1924);
or U1746 (N_1746,In_1508,In_1092);
or U1747 (N_1747,In_1328,In_983);
and U1748 (N_1748,In_1982,In_1556);
nor U1749 (N_1749,In_289,In_316);
nand U1750 (N_1750,In_1037,In_980);
nor U1751 (N_1751,In_14,In_997);
and U1752 (N_1752,In_375,In_1169);
nor U1753 (N_1753,In_1444,In_410);
or U1754 (N_1754,In_1333,In_856);
nor U1755 (N_1755,In_1600,In_276);
nor U1756 (N_1756,In_975,In_845);
nor U1757 (N_1757,In_1861,In_1737);
nand U1758 (N_1758,In_1317,In_407);
nor U1759 (N_1759,In_330,In_1486);
nor U1760 (N_1760,In_670,In_716);
and U1761 (N_1761,In_889,In_1225);
nor U1762 (N_1762,In_1029,In_1611);
nor U1763 (N_1763,In_1051,In_1374);
and U1764 (N_1764,In_1768,In_1196);
nor U1765 (N_1765,In_1166,In_1426);
nand U1766 (N_1766,In_947,In_1179);
or U1767 (N_1767,In_1906,In_947);
nor U1768 (N_1768,In_568,In_1913);
and U1769 (N_1769,In_1254,In_1115);
nand U1770 (N_1770,In_774,In_1400);
or U1771 (N_1771,In_1023,In_936);
nand U1772 (N_1772,In_304,In_422);
nand U1773 (N_1773,In_1402,In_693);
or U1774 (N_1774,In_1160,In_1184);
and U1775 (N_1775,In_1882,In_1011);
and U1776 (N_1776,In_1642,In_396);
or U1777 (N_1777,In_577,In_585);
or U1778 (N_1778,In_1187,In_523);
nand U1779 (N_1779,In_1762,In_1116);
nor U1780 (N_1780,In_282,In_877);
nand U1781 (N_1781,In_4,In_1698);
or U1782 (N_1782,In_204,In_1132);
nor U1783 (N_1783,In_1778,In_753);
nor U1784 (N_1784,In_620,In_269);
or U1785 (N_1785,In_1781,In_584);
or U1786 (N_1786,In_1479,In_618);
nand U1787 (N_1787,In_108,In_0);
or U1788 (N_1788,In_591,In_306);
nand U1789 (N_1789,In_1684,In_293);
xor U1790 (N_1790,In_926,In_441);
and U1791 (N_1791,In_1934,In_1454);
or U1792 (N_1792,In_172,In_496);
and U1793 (N_1793,In_1696,In_629);
and U1794 (N_1794,In_1882,In_1843);
nand U1795 (N_1795,In_1890,In_1995);
and U1796 (N_1796,In_136,In_1389);
nor U1797 (N_1797,In_549,In_688);
nand U1798 (N_1798,In_832,In_1790);
and U1799 (N_1799,In_1015,In_1036);
nand U1800 (N_1800,In_42,In_483);
nand U1801 (N_1801,In_671,In_639);
and U1802 (N_1802,In_1387,In_1037);
and U1803 (N_1803,In_368,In_1275);
and U1804 (N_1804,In_1327,In_663);
nand U1805 (N_1805,In_1202,In_1780);
nand U1806 (N_1806,In_1345,In_1533);
and U1807 (N_1807,In_1743,In_1992);
nor U1808 (N_1808,In_203,In_579);
and U1809 (N_1809,In_939,In_1983);
and U1810 (N_1810,In_1475,In_1423);
nand U1811 (N_1811,In_158,In_1921);
and U1812 (N_1812,In_1811,In_738);
nand U1813 (N_1813,In_508,In_186);
and U1814 (N_1814,In_979,In_601);
nor U1815 (N_1815,In_399,In_53);
and U1816 (N_1816,In_1895,In_1269);
nand U1817 (N_1817,In_52,In_194);
nor U1818 (N_1818,In_1744,In_1462);
nor U1819 (N_1819,In_1727,In_1568);
or U1820 (N_1820,In_1503,In_342);
and U1821 (N_1821,In_1778,In_1953);
and U1822 (N_1822,In_1536,In_1694);
nand U1823 (N_1823,In_921,In_894);
and U1824 (N_1824,In_1197,In_1563);
and U1825 (N_1825,In_1448,In_1358);
nand U1826 (N_1826,In_898,In_697);
nor U1827 (N_1827,In_1615,In_859);
and U1828 (N_1828,In_1795,In_546);
nand U1829 (N_1829,In_66,In_400);
or U1830 (N_1830,In_1390,In_169);
nor U1831 (N_1831,In_1151,In_828);
nand U1832 (N_1832,In_1131,In_946);
xor U1833 (N_1833,In_1133,In_1700);
nand U1834 (N_1834,In_899,In_1510);
and U1835 (N_1835,In_241,In_1653);
and U1836 (N_1836,In_901,In_1508);
nand U1837 (N_1837,In_119,In_730);
nand U1838 (N_1838,In_516,In_1098);
nor U1839 (N_1839,In_215,In_1487);
nand U1840 (N_1840,In_1663,In_984);
nor U1841 (N_1841,In_979,In_1366);
nand U1842 (N_1842,In_168,In_198);
and U1843 (N_1843,In_241,In_565);
nand U1844 (N_1844,In_1230,In_927);
nand U1845 (N_1845,In_1305,In_979);
nor U1846 (N_1846,In_1250,In_1378);
and U1847 (N_1847,In_107,In_30);
and U1848 (N_1848,In_1401,In_688);
and U1849 (N_1849,In_608,In_963);
nor U1850 (N_1850,In_527,In_1800);
nor U1851 (N_1851,In_1631,In_726);
nand U1852 (N_1852,In_1575,In_342);
nor U1853 (N_1853,In_579,In_616);
nor U1854 (N_1854,In_689,In_1419);
and U1855 (N_1855,In_861,In_808);
nand U1856 (N_1856,In_415,In_211);
nand U1857 (N_1857,In_94,In_1758);
and U1858 (N_1858,In_277,In_1922);
nand U1859 (N_1859,In_932,In_1937);
or U1860 (N_1860,In_269,In_1766);
nor U1861 (N_1861,In_1131,In_667);
nor U1862 (N_1862,In_278,In_1735);
nor U1863 (N_1863,In_1763,In_1205);
nor U1864 (N_1864,In_1980,In_1971);
and U1865 (N_1865,In_1657,In_1422);
nor U1866 (N_1866,In_1437,In_275);
nand U1867 (N_1867,In_1930,In_168);
nand U1868 (N_1868,In_1420,In_1586);
and U1869 (N_1869,In_1373,In_1042);
and U1870 (N_1870,In_150,In_638);
xnor U1871 (N_1871,In_1243,In_1351);
or U1872 (N_1872,In_1457,In_384);
and U1873 (N_1873,In_116,In_1870);
and U1874 (N_1874,In_430,In_76);
nor U1875 (N_1875,In_1077,In_1115);
or U1876 (N_1876,In_1235,In_818);
and U1877 (N_1877,In_1171,In_949);
and U1878 (N_1878,In_1928,In_1597);
or U1879 (N_1879,In_1611,In_610);
nor U1880 (N_1880,In_1499,In_1656);
and U1881 (N_1881,In_1220,In_1854);
or U1882 (N_1882,In_785,In_25);
nand U1883 (N_1883,In_1694,In_1107);
and U1884 (N_1884,In_969,In_406);
nand U1885 (N_1885,In_1446,In_1409);
nor U1886 (N_1886,In_533,In_1570);
nor U1887 (N_1887,In_564,In_724);
nor U1888 (N_1888,In_669,In_1768);
nand U1889 (N_1889,In_974,In_921);
and U1890 (N_1890,In_964,In_1831);
nand U1891 (N_1891,In_1874,In_118);
nor U1892 (N_1892,In_577,In_1478);
or U1893 (N_1893,In_1566,In_1092);
or U1894 (N_1894,In_37,In_1572);
nor U1895 (N_1895,In_595,In_890);
nor U1896 (N_1896,In_918,In_668);
or U1897 (N_1897,In_600,In_3);
nand U1898 (N_1898,In_653,In_238);
nand U1899 (N_1899,In_233,In_675);
or U1900 (N_1900,In_1440,In_1215);
and U1901 (N_1901,In_854,In_314);
or U1902 (N_1902,In_1490,In_1878);
and U1903 (N_1903,In_917,In_691);
nand U1904 (N_1904,In_571,In_1630);
nor U1905 (N_1905,In_1526,In_1387);
and U1906 (N_1906,In_742,In_872);
nand U1907 (N_1907,In_912,In_1717);
nand U1908 (N_1908,In_956,In_828);
nand U1909 (N_1909,In_343,In_1078);
nand U1910 (N_1910,In_969,In_394);
nand U1911 (N_1911,In_1046,In_265);
nor U1912 (N_1912,In_558,In_419);
and U1913 (N_1913,In_1096,In_1833);
and U1914 (N_1914,In_1587,In_280);
nand U1915 (N_1915,In_1548,In_1293);
and U1916 (N_1916,In_1082,In_1044);
or U1917 (N_1917,In_1086,In_1572);
nand U1918 (N_1918,In_1131,In_355);
and U1919 (N_1919,In_1737,In_19);
and U1920 (N_1920,In_1422,In_1114);
or U1921 (N_1921,In_1897,In_365);
and U1922 (N_1922,In_1351,In_74);
or U1923 (N_1923,In_1209,In_630);
nor U1924 (N_1924,In_638,In_1586);
nand U1925 (N_1925,In_1511,In_769);
and U1926 (N_1926,In_1753,In_1379);
or U1927 (N_1927,In_1682,In_1359);
nand U1928 (N_1928,In_1923,In_334);
nor U1929 (N_1929,In_1586,In_1500);
nand U1930 (N_1930,In_1814,In_1760);
nor U1931 (N_1931,In_381,In_66);
nor U1932 (N_1932,In_1283,In_360);
nor U1933 (N_1933,In_1189,In_1988);
and U1934 (N_1934,In_189,In_291);
and U1935 (N_1935,In_551,In_756);
nor U1936 (N_1936,In_994,In_82);
and U1937 (N_1937,In_852,In_230);
nand U1938 (N_1938,In_1434,In_1507);
and U1939 (N_1939,In_1917,In_1272);
nor U1940 (N_1940,In_93,In_604);
nor U1941 (N_1941,In_928,In_645);
and U1942 (N_1942,In_597,In_1166);
nand U1943 (N_1943,In_1705,In_1630);
or U1944 (N_1944,In_1429,In_1022);
nand U1945 (N_1945,In_1701,In_579);
nand U1946 (N_1946,In_321,In_68);
and U1947 (N_1947,In_893,In_524);
or U1948 (N_1948,In_707,In_1746);
nand U1949 (N_1949,In_1147,In_410);
and U1950 (N_1950,In_1587,In_1182);
or U1951 (N_1951,In_1569,In_1741);
or U1952 (N_1952,In_1857,In_1616);
or U1953 (N_1953,In_1487,In_1746);
or U1954 (N_1954,In_1168,In_1903);
nor U1955 (N_1955,In_1464,In_384);
or U1956 (N_1956,In_1970,In_1480);
nor U1957 (N_1957,In_679,In_259);
nand U1958 (N_1958,In_926,In_1398);
or U1959 (N_1959,In_1446,In_1092);
xnor U1960 (N_1960,In_615,In_153);
and U1961 (N_1961,In_243,In_518);
and U1962 (N_1962,In_19,In_590);
xnor U1963 (N_1963,In_883,In_1271);
nor U1964 (N_1964,In_1662,In_844);
or U1965 (N_1965,In_887,In_1601);
and U1966 (N_1966,In_354,In_1090);
nor U1967 (N_1967,In_798,In_1393);
or U1968 (N_1968,In_325,In_400);
nand U1969 (N_1969,In_393,In_1949);
nor U1970 (N_1970,In_333,In_342);
nor U1971 (N_1971,In_841,In_129);
or U1972 (N_1972,In_1872,In_1463);
and U1973 (N_1973,In_504,In_550);
and U1974 (N_1974,In_1869,In_405);
nor U1975 (N_1975,In_328,In_134);
and U1976 (N_1976,In_1696,In_1561);
and U1977 (N_1977,In_634,In_194);
nor U1978 (N_1978,In_21,In_1274);
nand U1979 (N_1979,In_339,In_117);
nor U1980 (N_1980,In_1531,In_1730);
nand U1981 (N_1981,In_1096,In_1418);
or U1982 (N_1982,In_1845,In_1275);
nor U1983 (N_1983,In_1008,In_1850);
and U1984 (N_1984,In_1513,In_1945);
or U1985 (N_1985,In_859,In_80);
nand U1986 (N_1986,In_170,In_1473);
or U1987 (N_1987,In_1746,In_406);
and U1988 (N_1988,In_1046,In_39);
and U1989 (N_1989,In_854,In_292);
nand U1990 (N_1990,In_789,In_1038);
and U1991 (N_1991,In_1605,In_1735);
or U1992 (N_1992,In_69,In_130);
nand U1993 (N_1993,In_1053,In_1949);
nor U1994 (N_1994,In_1733,In_354);
or U1995 (N_1995,In_248,In_1736);
nand U1996 (N_1996,In_223,In_299);
and U1997 (N_1997,In_536,In_892);
nor U1998 (N_1998,In_1021,In_1825);
nand U1999 (N_1999,In_1897,In_866);
and U2000 (N_2000,In_268,In_682);
or U2001 (N_2001,In_1480,In_42);
nand U2002 (N_2002,In_668,In_1906);
nor U2003 (N_2003,In_1311,In_621);
and U2004 (N_2004,In_1501,In_341);
and U2005 (N_2005,In_1570,In_735);
or U2006 (N_2006,In_1048,In_1252);
nor U2007 (N_2007,In_1554,In_1119);
and U2008 (N_2008,In_810,In_510);
nor U2009 (N_2009,In_1762,In_96);
or U2010 (N_2010,In_2,In_1309);
and U2011 (N_2011,In_938,In_428);
and U2012 (N_2012,In_998,In_573);
nor U2013 (N_2013,In_21,In_1692);
nor U2014 (N_2014,In_533,In_1133);
nand U2015 (N_2015,In_931,In_446);
and U2016 (N_2016,In_1601,In_1379);
nand U2017 (N_2017,In_952,In_53);
nor U2018 (N_2018,In_280,In_950);
nand U2019 (N_2019,In_673,In_216);
and U2020 (N_2020,In_641,In_1401);
nor U2021 (N_2021,In_1091,In_888);
or U2022 (N_2022,In_850,In_1887);
nor U2023 (N_2023,In_49,In_970);
nor U2024 (N_2024,In_1886,In_1290);
and U2025 (N_2025,In_1062,In_1203);
nand U2026 (N_2026,In_4,In_13);
nand U2027 (N_2027,In_733,In_1033);
nor U2028 (N_2028,In_1876,In_601);
nand U2029 (N_2029,In_1966,In_490);
nand U2030 (N_2030,In_767,In_261);
nor U2031 (N_2031,In_830,In_1601);
nand U2032 (N_2032,In_1369,In_179);
nand U2033 (N_2033,In_837,In_115);
and U2034 (N_2034,In_944,In_375);
and U2035 (N_2035,In_770,In_516);
xor U2036 (N_2036,In_900,In_1120);
and U2037 (N_2037,In_148,In_1810);
or U2038 (N_2038,In_1134,In_1020);
nand U2039 (N_2039,In_506,In_955);
nor U2040 (N_2040,In_1772,In_242);
nor U2041 (N_2041,In_739,In_944);
xor U2042 (N_2042,In_1848,In_1378);
or U2043 (N_2043,In_978,In_193);
and U2044 (N_2044,In_1766,In_1209);
nor U2045 (N_2045,In_967,In_1652);
nand U2046 (N_2046,In_527,In_1078);
nand U2047 (N_2047,In_373,In_1128);
and U2048 (N_2048,In_668,In_952);
and U2049 (N_2049,In_1335,In_732);
or U2050 (N_2050,In_837,In_427);
nor U2051 (N_2051,In_1322,In_272);
nand U2052 (N_2052,In_43,In_1968);
or U2053 (N_2053,In_1156,In_1812);
or U2054 (N_2054,In_1468,In_700);
or U2055 (N_2055,In_1279,In_1443);
or U2056 (N_2056,In_1024,In_963);
and U2057 (N_2057,In_686,In_1988);
nor U2058 (N_2058,In_1709,In_1058);
nand U2059 (N_2059,In_137,In_695);
or U2060 (N_2060,In_197,In_1548);
nand U2061 (N_2061,In_1757,In_229);
and U2062 (N_2062,In_583,In_293);
nor U2063 (N_2063,In_1598,In_1348);
nand U2064 (N_2064,In_1829,In_752);
or U2065 (N_2065,In_767,In_1797);
nor U2066 (N_2066,In_1619,In_41);
or U2067 (N_2067,In_1376,In_1381);
nand U2068 (N_2068,In_701,In_899);
nand U2069 (N_2069,In_1329,In_659);
or U2070 (N_2070,In_1506,In_644);
nand U2071 (N_2071,In_969,In_972);
nand U2072 (N_2072,In_202,In_1662);
nor U2073 (N_2073,In_1129,In_1061);
or U2074 (N_2074,In_275,In_837);
or U2075 (N_2075,In_839,In_1002);
or U2076 (N_2076,In_680,In_370);
xnor U2077 (N_2077,In_719,In_850);
nand U2078 (N_2078,In_1105,In_1506);
nand U2079 (N_2079,In_522,In_1547);
or U2080 (N_2080,In_1648,In_555);
and U2081 (N_2081,In_1566,In_1931);
or U2082 (N_2082,In_1351,In_1086);
or U2083 (N_2083,In_1124,In_288);
or U2084 (N_2084,In_1332,In_1351);
or U2085 (N_2085,In_1541,In_1818);
nand U2086 (N_2086,In_638,In_82);
and U2087 (N_2087,In_746,In_724);
or U2088 (N_2088,In_1254,In_1101);
and U2089 (N_2089,In_1180,In_1994);
or U2090 (N_2090,In_1324,In_432);
nor U2091 (N_2091,In_274,In_600);
nand U2092 (N_2092,In_1768,In_97);
and U2093 (N_2093,In_1891,In_467);
or U2094 (N_2094,In_957,In_1799);
nor U2095 (N_2095,In_1028,In_343);
nand U2096 (N_2096,In_298,In_922);
xor U2097 (N_2097,In_1082,In_891);
nand U2098 (N_2098,In_1278,In_155);
nand U2099 (N_2099,In_1025,In_1654);
nand U2100 (N_2100,In_356,In_527);
nand U2101 (N_2101,In_334,In_463);
nor U2102 (N_2102,In_1239,In_249);
nor U2103 (N_2103,In_421,In_1437);
or U2104 (N_2104,In_930,In_1230);
nand U2105 (N_2105,In_487,In_118);
nand U2106 (N_2106,In_1358,In_163);
and U2107 (N_2107,In_581,In_191);
or U2108 (N_2108,In_1324,In_886);
nor U2109 (N_2109,In_948,In_1827);
and U2110 (N_2110,In_910,In_1168);
xor U2111 (N_2111,In_1299,In_1298);
and U2112 (N_2112,In_1141,In_1980);
nand U2113 (N_2113,In_1353,In_1831);
nand U2114 (N_2114,In_1549,In_227);
nor U2115 (N_2115,In_336,In_1820);
nor U2116 (N_2116,In_1256,In_1254);
nand U2117 (N_2117,In_733,In_1643);
or U2118 (N_2118,In_1996,In_1321);
nand U2119 (N_2119,In_665,In_871);
and U2120 (N_2120,In_410,In_1877);
nand U2121 (N_2121,In_1711,In_407);
nor U2122 (N_2122,In_1969,In_410);
nor U2123 (N_2123,In_1176,In_290);
nand U2124 (N_2124,In_1398,In_1896);
or U2125 (N_2125,In_1114,In_1802);
or U2126 (N_2126,In_1063,In_1138);
nand U2127 (N_2127,In_1580,In_741);
or U2128 (N_2128,In_261,In_1258);
nor U2129 (N_2129,In_1526,In_1677);
or U2130 (N_2130,In_1400,In_436);
and U2131 (N_2131,In_864,In_41);
nor U2132 (N_2132,In_975,In_752);
and U2133 (N_2133,In_832,In_1889);
and U2134 (N_2134,In_882,In_876);
nand U2135 (N_2135,In_1616,In_141);
nand U2136 (N_2136,In_86,In_91);
nor U2137 (N_2137,In_194,In_1135);
nand U2138 (N_2138,In_5,In_1638);
or U2139 (N_2139,In_1439,In_507);
xor U2140 (N_2140,In_1173,In_1638);
nor U2141 (N_2141,In_590,In_580);
or U2142 (N_2142,In_574,In_1910);
nor U2143 (N_2143,In_1137,In_733);
and U2144 (N_2144,In_1023,In_1631);
nor U2145 (N_2145,In_144,In_1820);
and U2146 (N_2146,In_1639,In_672);
and U2147 (N_2147,In_302,In_1307);
or U2148 (N_2148,In_1516,In_1018);
nand U2149 (N_2149,In_1780,In_403);
or U2150 (N_2150,In_1929,In_1477);
nand U2151 (N_2151,In_749,In_522);
nor U2152 (N_2152,In_547,In_614);
xor U2153 (N_2153,In_1623,In_153);
or U2154 (N_2154,In_1945,In_359);
nand U2155 (N_2155,In_1618,In_555);
and U2156 (N_2156,In_901,In_56);
nor U2157 (N_2157,In_40,In_611);
and U2158 (N_2158,In_1482,In_1216);
nor U2159 (N_2159,In_932,In_1733);
nor U2160 (N_2160,In_1603,In_775);
nor U2161 (N_2161,In_1998,In_1817);
nand U2162 (N_2162,In_1103,In_425);
and U2163 (N_2163,In_509,In_1808);
nand U2164 (N_2164,In_590,In_1435);
and U2165 (N_2165,In_1218,In_1884);
or U2166 (N_2166,In_643,In_1747);
and U2167 (N_2167,In_940,In_1891);
nand U2168 (N_2168,In_1601,In_1424);
or U2169 (N_2169,In_570,In_1889);
nand U2170 (N_2170,In_954,In_1993);
or U2171 (N_2171,In_1603,In_1377);
and U2172 (N_2172,In_1554,In_258);
nor U2173 (N_2173,In_1991,In_1148);
or U2174 (N_2174,In_1893,In_693);
nor U2175 (N_2175,In_447,In_1745);
nand U2176 (N_2176,In_1808,In_907);
nand U2177 (N_2177,In_1615,In_95);
nor U2178 (N_2178,In_341,In_1382);
xnor U2179 (N_2179,In_444,In_1742);
or U2180 (N_2180,In_798,In_533);
or U2181 (N_2181,In_1402,In_899);
nor U2182 (N_2182,In_820,In_300);
and U2183 (N_2183,In_702,In_1045);
nand U2184 (N_2184,In_1500,In_219);
or U2185 (N_2185,In_1167,In_215);
nor U2186 (N_2186,In_618,In_264);
nor U2187 (N_2187,In_776,In_627);
or U2188 (N_2188,In_1277,In_538);
or U2189 (N_2189,In_1260,In_1389);
nand U2190 (N_2190,In_475,In_1385);
nand U2191 (N_2191,In_340,In_1852);
nor U2192 (N_2192,In_1425,In_1936);
nor U2193 (N_2193,In_95,In_1609);
nand U2194 (N_2194,In_1812,In_258);
nand U2195 (N_2195,In_592,In_672);
nand U2196 (N_2196,In_24,In_700);
nor U2197 (N_2197,In_854,In_198);
nand U2198 (N_2198,In_1983,In_1273);
nand U2199 (N_2199,In_1175,In_722);
or U2200 (N_2200,In_210,In_1480);
xnor U2201 (N_2201,In_1067,In_1460);
or U2202 (N_2202,In_512,In_124);
nor U2203 (N_2203,In_962,In_417);
nand U2204 (N_2204,In_1634,In_1973);
and U2205 (N_2205,In_429,In_934);
nand U2206 (N_2206,In_1876,In_509);
nand U2207 (N_2207,In_797,In_838);
or U2208 (N_2208,In_283,In_1868);
nand U2209 (N_2209,In_1679,In_484);
or U2210 (N_2210,In_918,In_294);
nand U2211 (N_2211,In_285,In_8);
and U2212 (N_2212,In_43,In_1652);
nand U2213 (N_2213,In_759,In_198);
and U2214 (N_2214,In_786,In_344);
nor U2215 (N_2215,In_1743,In_672);
nor U2216 (N_2216,In_830,In_1774);
nor U2217 (N_2217,In_881,In_121);
xnor U2218 (N_2218,In_1131,In_798);
nor U2219 (N_2219,In_339,In_140);
and U2220 (N_2220,In_964,In_300);
and U2221 (N_2221,In_494,In_1236);
or U2222 (N_2222,In_1851,In_362);
or U2223 (N_2223,In_1681,In_1253);
and U2224 (N_2224,In_471,In_261);
nand U2225 (N_2225,In_1688,In_934);
xnor U2226 (N_2226,In_174,In_1851);
or U2227 (N_2227,In_1697,In_1780);
or U2228 (N_2228,In_597,In_59);
nor U2229 (N_2229,In_343,In_629);
nand U2230 (N_2230,In_70,In_1358);
nor U2231 (N_2231,In_621,In_1530);
nor U2232 (N_2232,In_1489,In_977);
nand U2233 (N_2233,In_285,In_293);
nor U2234 (N_2234,In_659,In_992);
nand U2235 (N_2235,In_860,In_1973);
nor U2236 (N_2236,In_1408,In_233);
and U2237 (N_2237,In_531,In_1825);
and U2238 (N_2238,In_1665,In_642);
nor U2239 (N_2239,In_1126,In_627);
or U2240 (N_2240,In_1860,In_1434);
nor U2241 (N_2241,In_1292,In_1353);
nand U2242 (N_2242,In_1896,In_373);
and U2243 (N_2243,In_1408,In_1512);
xnor U2244 (N_2244,In_1343,In_605);
nand U2245 (N_2245,In_333,In_890);
and U2246 (N_2246,In_1516,In_112);
and U2247 (N_2247,In_46,In_1876);
or U2248 (N_2248,In_122,In_1859);
nor U2249 (N_2249,In_1797,In_276);
nand U2250 (N_2250,In_125,In_1948);
or U2251 (N_2251,In_476,In_1258);
nor U2252 (N_2252,In_1085,In_1131);
or U2253 (N_2253,In_1907,In_1057);
nand U2254 (N_2254,In_299,In_381);
nand U2255 (N_2255,In_1137,In_392);
nor U2256 (N_2256,In_644,In_1675);
nand U2257 (N_2257,In_842,In_628);
and U2258 (N_2258,In_291,In_1411);
nor U2259 (N_2259,In_1382,In_1683);
nor U2260 (N_2260,In_1637,In_101);
or U2261 (N_2261,In_270,In_1688);
and U2262 (N_2262,In_363,In_1012);
or U2263 (N_2263,In_936,In_1774);
nand U2264 (N_2264,In_1419,In_1545);
nor U2265 (N_2265,In_1540,In_1115);
nand U2266 (N_2266,In_1118,In_144);
nand U2267 (N_2267,In_664,In_288);
nor U2268 (N_2268,In_1613,In_938);
nand U2269 (N_2269,In_1812,In_521);
nor U2270 (N_2270,In_1724,In_721);
and U2271 (N_2271,In_1481,In_325);
nand U2272 (N_2272,In_557,In_856);
nand U2273 (N_2273,In_432,In_1738);
nand U2274 (N_2274,In_1449,In_775);
nor U2275 (N_2275,In_1251,In_1989);
and U2276 (N_2276,In_252,In_1413);
and U2277 (N_2277,In_178,In_878);
or U2278 (N_2278,In_398,In_797);
nor U2279 (N_2279,In_1743,In_1928);
nor U2280 (N_2280,In_359,In_1181);
and U2281 (N_2281,In_702,In_108);
nor U2282 (N_2282,In_196,In_838);
nand U2283 (N_2283,In_61,In_1907);
or U2284 (N_2284,In_581,In_1754);
and U2285 (N_2285,In_206,In_1970);
or U2286 (N_2286,In_759,In_1942);
nand U2287 (N_2287,In_591,In_933);
and U2288 (N_2288,In_127,In_1215);
nand U2289 (N_2289,In_53,In_866);
or U2290 (N_2290,In_1086,In_1901);
nand U2291 (N_2291,In_979,In_1671);
or U2292 (N_2292,In_1121,In_340);
or U2293 (N_2293,In_866,In_1548);
nor U2294 (N_2294,In_747,In_242);
nor U2295 (N_2295,In_312,In_1285);
and U2296 (N_2296,In_997,In_719);
and U2297 (N_2297,In_827,In_1805);
or U2298 (N_2298,In_1827,In_1339);
nor U2299 (N_2299,In_537,In_1801);
and U2300 (N_2300,In_1830,In_1668);
nor U2301 (N_2301,In_32,In_1472);
nand U2302 (N_2302,In_1675,In_1826);
nand U2303 (N_2303,In_1175,In_706);
nand U2304 (N_2304,In_897,In_1839);
or U2305 (N_2305,In_1377,In_1768);
and U2306 (N_2306,In_1120,In_1652);
or U2307 (N_2307,In_1645,In_1049);
or U2308 (N_2308,In_1716,In_907);
or U2309 (N_2309,In_1748,In_229);
or U2310 (N_2310,In_1388,In_257);
or U2311 (N_2311,In_1436,In_491);
or U2312 (N_2312,In_1332,In_1715);
nor U2313 (N_2313,In_705,In_485);
nand U2314 (N_2314,In_1897,In_1707);
nor U2315 (N_2315,In_1825,In_962);
or U2316 (N_2316,In_1630,In_1295);
nand U2317 (N_2317,In_1711,In_954);
nand U2318 (N_2318,In_1716,In_1622);
or U2319 (N_2319,In_1759,In_1369);
nand U2320 (N_2320,In_1047,In_765);
nor U2321 (N_2321,In_541,In_1115);
or U2322 (N_2322,In_1835,In_1125);
nor U2323 (N_2323,In_1566,In_30);
and U2324 (N_2324,In_248,In_1898);
nand U2325 (N_2325,In_205,In_1293);
and U2326 (N_2326,In_692,In_1433);
and U2327 (N_2327,In_1706,In_1532);
and U2328 (N_2328,In_1073,In_1853);
nand U2329 (N_2329,In_1888,In_1431);
nor U2330 (N_2330,In_1796,In_1145);
nand U2331 (N_2331,In_140,In_1760);
nand U2332 (N_2332,In_1318,In_1349);
and U2333 (N_2333,In_1486,In_105);
and U2334 (N_2334,In_1420,In_1662);
nor U2335 (N_2335,In_437,In_1566);
or U2336 (N_2336,In_1203,In_1357);
or U2337 (N_2337,In_10,In_353);
or U2338 (N_2338,In_506,In_753);
or U2339 (N_2339,In_311,In_1429);
and U2340 (N_2340,In_1864,In_1495);
nand U2341 (N_2341,In_1890,In_147);
nand U2342 (N_2342,In_376,In_1510);
or U2343 (N_2343,In_553,In_180);
and U2344 (N_2344,In_1264,In_637);
nor U2345 (N_2345,In_16,In_1832);
nand U2346 (N_2346,In_1863,In_1557);
nand U2347 (N_2347,In_1750,In_1719);
nand U2348 (N_2348,In_1721,In_1650);
or U2349 (N_2349,In_1146,In_1604);
nor U2350 (N_2350,In_1445,In_1341);
or U2351 (N_2351,In_800,In_717);
nor U2352 (N_2352,In_774,In_1247);
nand U2353 (N_2353,In_306,In_1833);
nor U2354 (N_2354,In_384,In_1354);
and U2355 (N_2355,In_1702,In_1493);
and U2356 (N_2356,In_1154,In_1768);
nand U2357 (N_2357,In_815,In_1253);
and U2358 (N_2358,In_1709,In_1172);
or U2359 (N_2359,In_1885,In_1945);
nor U2360 (N_2360,In_1355,In_712);
or U2361 (N_2361,In_348,In_252);
or U2362 (N_2362,In_1583,In_1393);
nand U2363 (N_2363,In_1614,In_1051);
nor U2364 (N_2364,In_382,In_1872);
and U2365 (N_2365,In_856,In_1086);
nor U2366 (N_2366,In_485,In_1298);
nand U2367 (N_2367,In_1381,In_124);
nor U2368 (N_2368,In_1693,In_381);
nor U2369 (N_2369,In_801,In_1955);
and U2370 (N_2370,In_1795,In_1560);
or U2371 (N_2371,In_897,In_1418);
nor U2372 (N_2372,In_1776,In_1907);
or U2373 (N_2373,In_270,In_1970);
or U2374 (N_2374,In_977,In_1579);
and U2375 (N_2375,In_441,In_791);
nor U2376 (N_2376,In_1546,In_1911);
nor U2377 (N_2377,In_426,In_1165);
nor U2378 (N_2378,In_1605,In_1928);
nand U2379 (N_2379,In_1557,In_846);
nor U2380 (N_2380,In_1097,In_430);
nand U2381 (N_2381,In_537,In_504);
nor U2382 (N_2382,In_1563,In_1136);
nor U2383 (N_2383,In_1925,In_895);
nand U2384 (N_2384,In_1198,In_1805);
nand U2385 (N_2385,In_501,In_1246);
nand U2386 (N_2386,In_559,In_151);
nor U2387 (N_2387,In_161,In_690);
nand U2388 (N_2388,In_1444,In_777);
and U2389 (N_2389,In_1520,In_693);
and U2390 (N_2390,In_954,In_765);
nor U2391 (N_2391,In_718,In_727);
nand U2392 (N_2392,In_909,In_1936);
nor U2393 (N_2393,In_83,In_1386);
nor U2394 (N_2394,In_1663,In_337);
or U2395 (N_2395,In_1188,In_1267);
nand U2396 (N_2396,In_876,In_1209);
nor U2397 (N_2397,In_865,In_1766);
nand U2398 (N_2398,In_1359,In_445);
nand U2399 (N_2399,In_1739,In_1203);
nor U2400 (N_2400,In_739,In_1330);
nor U2401 (N_2401,In_959,In_1376);
or U2402 (N_2402,In_242,In_1259);
nor U2403 (N_2403,In_215,In_282);
nor U2404 (N_2404,In_145,In_137);
and U2405 (N_2405,In_1685,In_1054);
nor U2406 (N_2406,In_695,In_1284);
or U2407 (N_2407,In_654,In_1260);
nand U2408 (N_2408,In_820,In_1339);
and U2409 (N_2409,In_634,In_1604);
nor U2410 (N_2410,In_488,In_1629);
nand U2411 (N_2411,In_458,In_1073);
or U2412 (N_2412,In_259,In_1192);
nor U2413 (N_2413,In_183,In_1344);
and U2414 (N_2414,In_1267,In_1795);
nor U2415 (N_2415,In_164,In_1334);
or U2416 (N_2416,In_391,In_254);
nor U2417 (N_2417,In_855,In_185);
or U2418 (N_2418,In_808,In_1539);
nor U2419 (N_2419,In_1092,In_1308);
and U2420 (N_2420,In_891,In_13);
nand U2421 (N_2421,In_1018,In_703);
nand U2422 (N_2422,In_1054,In_522);
nor U2423 (N_2423,In_24,In_348);
and U2424 (N_2424,In_226,In_1334);
and U2425 (N_2425,In_1477,In_1198);
nand U2426 (N_2426,In_1414,In_1096);
or U2427 (N_2427,In_1143,In_1102);
or U2428 (N_2428,In_211,In_1587);
nand U2429 (N_2429,In_959,In_14);
nor U2430 (N_2430,In_1482,In_726);
and U2431 (N_2431,In_1908,In_132);
or U2432 (N_2432,In_1944,In_1178);
nand U2433 (N_2433,In_1158,In_739);
nand U2434 (N_2434,In_1120,In_1360);
nor U2435 (N_2435,In_963,In_881);
nand U2436 (N_2436,In_1017,In_211);
nand U2437 (N_2437,In_274,In_669);
and U2438 (N_2438,In_1421,In_190);
or U2439 (N_2439,In_723,In_1361);
and U2440 (N_2440,In_363,In_942);
nor U2441 (N_2441,In_827,In_779);
nand U2442 (N_2442,In_758,In_1071);
and U2443 (N_2443,In_74,In_1941);
nand U2444 (N_2444,In_366,In_1502);
and U2445 (N_2445,In_461,In_532);
nand U2446 (N_2446,In_852,In_77);
nand U2447 (N_2447,In_1865,In_549);
nor U2448 (N_2448,In_127,In_1388);
or U2449 (N_2449,In_786,In_90);
nand U2450 (N_2450,In_909,In_681);
or U2451 (N_2451,In_274,In_1309);
or U2452 (N_2452,In_1276,In_1842);
xor U2453 (N_2453,In_785,In_1889);
or U2454 (N_2454,In_1650,In_559);
and U2455 (N_2455,In_156,In_1047);
nor U2456 (N_2456,In_827,In_1018);
nand U2457 (N_2457,In_453,In_1937);
or U2458 (N_2458,In_1905,In_675);
nor U2459 (N_2459,In_1313,In_1981);
nor U2460 (N_2460,In_299,In_33);
or U2461 (N_2461,In_494,In_1514);
nor U2462 (N_2462,In_1751,In_3);
and U2463 (N_2463,In_1657,In_177);
nor U2464 (N_2464,In_813,In_1579);
or U2465 (N_2465,In_1197,In_1921);
and U2466 (N_2466,In_1380,In_1516);
or U2467 (N_2467,In_1181,In_381);
nand U2468 (N_2468,In_1058,In_1409);
nor U2469 (N_2469,In_1327,In_710);
nand U2470 (N_2470,In_133,In_1650);
and U2471 (N_2471,In_1871,In_1260);
or U2472 (N_2472,In_1214,In_851);
nand U2473 (N_2473,In_613,In_152);
or U2474 (N_2474,In_993,In_1443);
nor U2475 (N_2475,In_795,In_790);
and U2476 (N_2476,In_436,In_723);
and U2477 (N_2477,In_1571,In_1980);
and U2478 (N_2478,In_1330,In_1776);
nor U2479 (N_2479,In_960,In_1600);
nor U2480 (N_2480,In_298,In_437);
nand U2481 (N_2481,In_1322,In_1361);
nand U2482 (N_2482,In_1667,In_963);
nand U2483 (N_2483,In_519,In_0);
nand U2484 (N_2484,In_997,In_214);
nor U2485 (N_2485,In_75,In_427);
nor U2486 (N_2486,In_1256,In_1223);
nor U2487 (N_2487,In_1076,In_1209);
or U2488 (N_2488,In_728,In_623);
nor U2489 (N_2489,In_198,In_1656);
nor U2490 (N_2490,In_288,In_1274);
and U2491 (N_2491,In_728,In_1552);
nor U2492 (N_2492,In_473,In_1472);
nor U2493 (N_2493,In_1631,In_1828);
nor U2494 (N_2494,In_1998,In_1150);
nor U2495 (N_2495,In_1801,In_1529);
nand U2496 (N_2496,In_560,In_1033);
nor U2497 (N_2497,In_1911,In_556);
and U2498 (N_2498,In_1539,In_1268);
and U2499 (N_2499,In_281,In_1956);
and U2500 (N_2500,In_1210,In_1041);
nand U2501 (N_2501,In_1187,In_1507);
nor U2502 (N_2502,In_833,In_1299);
or U2503 (N_2503,In_1980,In_1922);
nand U2504 (N_2504,In_391,In_1414);
and U2505 (N_2505,In_1599,In_346);
and U2506 (N_2506,In_1507,In_649);
nand U2507 (N_2507,In_1737,In_1297);
nor U2508 (N_2508,In_1336,In_1959);
and U2509 (N_2509,In_350,In_1602);
nor U2510 (N_2510,In_1206,In_831);
nor U2511 (N_2511,In_1971,In_1828);
and U2512 (N_2512,In_1974,In_1833);
or U2513 (N_2513,In_106,In_1264);
or U2514 (N_2514,In_321,In_1128);
or U2515 (N_2515,In_1084,In_1922);
nor U2516 (N_2516,In_1057,In_1903);
and U2517 (N_2517,In_235,In_99);
nand U2518 (N_2518,In_1261,In_1966);
or U2519 (N_2519,In_1599,In_541);
and U2520 (N_2520,In_564,In_699);
or U2521 (N_2521,In_1580,In_1436);
nor U2522 (N_2522,In_1756,In_1403);
nand U2523 (N_2523,In_1794,In_377);
and U2524 (N_2524,In_1156,In_14);
nor U2525 (N_2525,In_1944,In_41);
nor U2526 (N_2526,In_1773,In_296);
or U2527 (N_2527,In_1509,In_986);
or U2528 (N_2528,In_524,In_1394);
nor U2529 (N_2529,In_631,In_1038);
nand U2530 (N_2530,In_293,In_494);
nor U2531 (N_2531,In_1343,In_460);
nor U2532 (N_2532,In_1444,In_989);
and U2533 (N_2533,In_1702,In_2);
and U2534 (N_2534,In_1195,In_1758);
nor U2535 (N_2535,In_1702,In_788);
and U2536 (N_2536,In_332,In_1229);
nand U2537 (N_2537,In_1201,In_381);
nand U2538 (N_2538,In_1180,In_1798);
or U2539 (N_2539,In_1598,In_1961);
nor U2540 (N_2540,In_798,In_1633);
and U2541 (N_2541,In_145,In_1372);
and U2542 (N_2542,In_273,In_348);
nor U2543 (N_2543,In_1981,In_1214);
and U2544 (N_2544,In_792,In_952);
and U2545 (N_2545,In_667,In_1451);
or U2546 (N_2546,In_745,In_1936);
and U2547 (N_2547,In_1131,In_0);
or U2548 (N_2548,In_393,In_394);
nand U2549 (N_2549,In_1010,In_1266);
nand U2550 (N_2550,In_85,In_603);
xor U2551 (N_2551,In_1251,In_363);
nor U2552 (N_2552,In_1486,In_994);
nand U2553 (N_2553,In_24,In_34);
nor U2554 (N_2554,In_452,In_1865);
nand U2555 (N_2555,In_1380,In_535);
and U2556 (N_2556,In_1458,In_1032);
nor U2557 (N_2557,In_496,In_1505);
nor U2558 (N_2558,In_1757,In_528);
and U2559 (N_2559,In_833,In_352);
nor U2560 (N_2560,In_492,In_591);
or U2561 (N_2561,In_1250,In_1779);
nor U2562 (N_2562,In_1028,In_301);
xor U2563 (N_2563,In_1621,In_1816);
nor U2564 (N_2564,In_861,In_1623);
and U2565 (N_2565,In_1892,In_558);
and U2566 (N_2566,In_1628,In_1235);
nand U2567 (N_2567,In_1740,In_75);
or U2568 (N_2568,In_740,In_1923);
and U2569 (N_2569,In_12,In_1257);
and U2570 (N_2570,In_1751,In_505);
or U2571 (N_2571,In_1865,In_1615);
and U2572 (N_2572,In_1376,In_261);
nand U2573 (N_2573,In_552,In_763);
and U2574 (N_2574,In_717,In_1737);
nor U2575 (N_2575,In_1620,In_1307);
or U2576 (N_2576,In_307,In_1131);
or U2577 (N_2577,In_1309,In_504);
and U2578 (N_2578,In_1156,In_1548);
and U2579 (N_2579,In_1259,In_939);
nand U2580 (N_2580,In_1719,In_1801);
nand U2581 (N_2581,In_624,In_389);
or U2582 (N_2582,In_1012,In_15);
and U2583 (N_2583,In_1366,In_456);
nor U2584 (N_2584,In_1992,In_631);
nand U2585 (N_2585,In_697,In_1302);
or U2586 (N_2586,In_661,In_611);
nor U2587 (N_2587,In_42,In_1282);
or U2588 (N_2588,In_1371,In_645);
and U2589 (N_2589,In_1092,In_38);
or U2590 (N_2590,In_33,In_701);
xor U2591 (N_2591,In_1310,In_1782);
nand U2592 (N_2592,In_999,In_1117);
nor U2593 (N_2593,In_714,In_608);
nand U2594 (N_2594,In_360,In_1784);
nand U2595 (N_2595,In_847,In_421);
or U2596 (N_2596,In_1310,In_142);
nor U2597 (N_2597,In_1412,In_1190);
nor U2598 (N_2598,In_1676,In_755);
or U2599 (N_2599,In_32,In_1841);
or U2600 (N_2600,In_1417,In_405);
or U2601 (N_2601,In_207,In_1009);
and U2602 (N_2602,In_618,In_996);
nor U2603 (N_2603,In_1436,In_66);
nand U2604 (N_2604,In_1034,In_656);
and U2605 (N_2605,In_1324,In_734);
nor U2606 (N_2606,In_1556,In_480);
nand U2607 (N_2607,In_1774,In_1583);
nor U2608 (N_2608,In_18,In_1155);
and U2609 (N_2609,In_81,In_897);
nor U2610 (N_2610,In_1119,In_1555);
and U2611 (N_2611,In_1508,In_547);
nor U2612 (N_2612,In_277,In_1941);
nand U2613 (N_2613,In_191,In_1858);
or U2614 (N_2614,In_1184,In_1392);
nand U2615 (N_2615,In_1082,In_271);
xnor U2616 (N_2616,In_18,In_108);
nand U2617 (N_2617,In_1228,In_886);
nand U2618 (N_2618,In_1987,In_1886);
nor U2619 (N_2619,In_1334,In_1959);
nand U2620 (N_2620,In_84,In_1527);
or U2621 (N_2621,In_363,In_1299);
nand U2622 (N_2622,In_1843,In_1069);
xor U2623 (N_2623,In_496,In_1320);
nor U2624 (N_2624,In_544,In_1681);
and U2625 (N_2625,In_321,In_721);
nor U2626 (N_2626,In_1448,In_1395);
nor U2627 (N_2627,In_383,In_216);
and U2628 (N_2628,In_56,In_934);
or U2629 (N_2629,In_1047,In_137);
and U2630 (N_2630,In_46,In_177);
nor U2631 (N_2631,In_494,In_949);
nand U2632 (N_2632,In_1876,In_1691);
and U2633 (N_2633,In_1017,In_52);
or U2634 (N_2634,In_1792,In_1745);
and U2635 (N_2635,In_253,In_1322);
nand U2636 (N_2636,In_443,In_1482);
nand U2637 (N_2637,In_363,In_1508);
nand U2638 (N_2638,In_706,In_399);
nand U2639 (N_2639,In_1478,In_631);
or U2640 (N_2640,In_155,In_1859);
nand U2641 (N_2641,In_1495,In_612);
xor U2642 (N_2642,In_1539,In_1718);
nor U2643 (N_2643,In_1290,In_683);
nand U2644 (N_2644,In_1170,In_1627);
or U2645 (N_2645,In_1942,In_749);
or U2646 (N_2646,In_1111,In_758);
or U2647 (N_2647,In_968,In_580);
nor U2648 (N_2648,In_1150,In_192);
or U2649 (N_2649,In_1486,In_1904);
and U2650 (N_2650,In_1977,In_1710);
or U2651 (N_2651,In_1235,In_1915);
or U2652 (N_2652,In_319,In_1623);
nand U2653 (N_2653,In_231,In_1801);
nand U2654 (N_2654,In_856,In_306);
nor U2655 (N_2655,In_1620,In_1315);
nor U2656 (N_2656,In_1640,In_536);
or U2657 (N_2657,In_1530,In_1675);
and U2658 (N_2658,In_166,In_1875);
xor U2659 (N_2659,In_1724,In_63);
nand U2660 (N_2660,In_1936,In_1865);
nand U2661 (N_2661,In_467,In_701);
nor U2662 (N_2662,In_1317,In_1096);
or U2663 (N_2663,In_257,In_557);
nand U2664 (N_2664,In_1724,In_1834);
or U2665 (N_2665,In_1110,In_293);
nor U2666 (N_2666,In_948,In_213);
and U2667 (N_2667,In_675,In_973);
nor U2668 (N_2668,In_245,In_1495);
nor U2669 (N_2669,In_1289,In_426);
nor U2670 (N_2670,In_1334,In_1473);
or U2671 (N_2671,In_423,In_451);
or U2672 (N_2672,In_1708,In_1378);
nand U2673 (N_2673,In_394,In_456);
nand U2674 (N_2674,In_495,In_280);
and U2675 (N_2675,In_1765,In_502);
nor U2676 (N_2676,In_251,In_377);
xor U2677 (N_2677,In_1814,In_1822);
and U2678 (N_2678,In_340,In_1374);
and U2679 (N_2679,In_1034,In_430);
nand U2680 (N_2680,In_360,In_46);
nor U2681 (N_2681,In_619,In_659);
nand U2682 (N_2682,In_1638,In_1782);
and U2683 (N_2683,In_1760,In_1932);
xnor U2684 (N_2684,In_450,In_783);
nand U2685 (N_2685,In_1933,In_1999);
and U2686 (N_2686,In_864,In_564);
or U2687 (N_2687,In_193,In_1758);
or U2688 (N_2688,In_564,In_608);
or U2689 (N_2689,In_1948,In_798);
nor U2690 (N_2690,In_47,In_963);
nand U2691 (N_2691,In_81,In_357);
xor U2692 (N_2692,In_1776,In_839);
nor U2693 (N_2693,In_913,In_329);
nor U2694 (N_2694,In_1119,In_360);
nor U2695 (N_2695,In_732,In_274);
or U2696 (N_2696,In_335,In_1084);
nor U2697 (N_2697,In_1949,In_119);
nand U2698 (N_2698,In_1854,In_1707);
nor U2699 (N_2699,In_594,In_992);
nand U2700 (N_2700,In_1468,In_1594);
nor U2701 (N_2701,In_394,In_1002);
nand U2702 (N_2702,In_1420,In_978);
and U2703 (N_2703,In_1512,In_1957);
nor U2704 (N_2704,In_1873,In_891);
nor U2705 (N_2705,In_706,In_1563);
nand U2706 (N_2706,In_1466,In_1252);
or U2707 (N_2707,In_476,In_1826);
nor U2708 (N_2708,In_918,In_1493);
nor U2709 (N_2709,In_895,In_718);
or U2710 (N_2710,In_1218,In_1438);
and U2711 (N_2711,In_1045,In_76);
or U2712 (N_2712,In_531,In_528);
nand U2713 (N_2713,In_184,In_1758);
xor U2714 (N_2714,In_1719,In_1497);
and U2715 (N_2715,In_520,In_1164);
or U2716 (N_2716,In_1935,In_1985);
or U2717 (N_2717,In_899,In_876);
and U2718 (N_2718,In_1723,In_939);
nand U2719 (N_2719,In_890,In_686);
nand U2720 (N_2720,In_203,In_1651);
nand U2721 (N_2721,In_1403,In_1299);
nand U2722 (N_2722,In_345,In_587);
or U2723 (N_2723,In_584,In_1053);
and U2724 (N_2724,In_1952,In_1239);
and U2725 (N_2725,In_1449,In_197);
and U2726 (N_2726,In_1754,In_51);
nand U2727 (N_2727,In_948,In_214);
nand U2728 (N_2728,In_1787,In_278);
nand U2729 (N_2729,In_1571,In_1778);
or U2730 (N_2730,In_223,In_790);
and U2731 (N_2731,In_1107,In_585);
nand U2732 (N_2732,In_152,In_1772);
nand U2733 (N_2733,In_1606,In_552);
or U2734 (N_2734,In_741,In_272);
and U2735 (N_2735,In_430,In_1217);
or U2736 (N_2736,In_391,In_239);
nand U2737 (N_2737,In_757,In_723);
and U2738 (N_2738,In_89,In_1481);
nand U2739 (N_2739,In_493,In_690);
and U2740 (N_2740,In_855,In_369);
nand U2741 (N_2741,In_635,In_178);
nor U2742 (N_2742,In_1492,In_1743);
or U2743 (N_2743,In_519,In_54);
and U2744 (N_2744,In_1823,In_38);
nand U2745 (N_2745,In_729,In_576);
nand U2746 (N_2746,In_1038,In_442);
nand U2747 (N_2747,In_840,In_1893);
and U2748 (N_2748,In_1404,In_105);
nor U2749 (N_2749,In_1292,In_784);
or U2750 (N_2750,In_720,In_1227);
nor U2751 (N_2751,In_1224,In_1664);
and U2752 (N_2752,In_1364,In_177);
and U2753 (N_2753,In_346,In_392);
and U2754 (N_2754,In_1450,In_19);
and U2755 (N_2755,In_1187,In_1719);
nor U2756 (N_2756,In_1930,In_246);
nor U2757 (N_2757,In_1887,In_225);
nand U2758 (N_2758,In_1686,In_559);
or U2759 (N_2759,In_859,In_26);
and U2760 (N_2760,In_214,In_1231);
or U2761 (N_2761,In_6,In_885);
and U2762 (N_2762,In_1488,In_680);
nand U2763 (N_2763,In_594,In_1310);
nand U2764 (N_2764,In_187,In_740);
nand U2765 (N_2765,In_1818,In_1323);
nor U2766 (N_2766,In_1906,In_1364);
nor U2767 (N_2767,In_674,In_1443);
nand U2768 (N_2768,In_1898,In_1497);
and U2769 (N_2769,In_619,In_1928);
or U2770 (N_2770,In_1102,In_1960);
or U2771 (N_2771,In_624,In_1985);
and U2772 (N_2772,In_445,In_1464);
and U2773 (N_2773,In_434,In_1240);
or U2774 (N_2774,In_1593,In_1320);
or U2775 (N_2775,In_1956,In_1913);
or U2776 (N_2776,In_1594,In_448);
or U2777 (N_2777,In_1050,In_1644);
and U2778 (N_2778,In_1158,In_279);
and U2779 (N_2779,In_1728,In_22);
nand U2780 (N_2780,In_1969,In_764);
nand U2781 (N_2781,In_1955,In_17);
and U2782 (N_2782,In_423,In_806);
or U2783 (N_2783,In_974,In_1913);
nand U2784 (N_2784,In_368,In_1728);
and U2785 (N_2785,In_552,In_759);
nor U2786 (N_2786,In_1846,In_778);
nand U2787 (N_2787,In_1394,In_1975);
and U2788 (N_2788,In_1700,In_1890);
nor U2789 (N_2789,In_1032,In_1429);
nand U2790 (N_2790,In_483,In_1201);
nand U2791 (N_2791,In_402,In_1770);
nor U2792 (N_2792,In_40,In_1625);
and U2793 (N_2793,In_1942,In_590);
nand U2794 (N_2794,In_251,In_1265);
and U2795 (N_2795,In_1097,In_203);
nand U2796 (N_2796,In_407,In_1546);
or U2797 (N_2797,In_1243,In_307);
or U2798 (N_2798,In_426,In_794);
and U2799 (N_2799,In_1174,In_1659);
or U2800 (N_2800,In_1098,In_1675);
nor U2801 (N_2801,In_287,In_596);
and U2802 (N_2802,In_1319,In_916);
and U2803 (N_2803,In_1884,In_1878);
nor U2804 (N_2804,In_944,In_96);
nor U2805 (N_2805,In_1158,In_1432);
nor U2806 (N_2806,In_906,In_622);
nand U2807 (N_2807,In_318,In_570);
or U2808 (N_2808,In_1503,In_1146);
or U2809 (N_2809,In_847,In_154);
nor U2810 (N_2810,In_1576,In_1437);
nand U2811 (N_2811,In_1069,In_575);
or U2812 (N_2812,In_1242,In_776);
nor U2813 (N_2813,In_1901,In_68);
or U2814 (N_2814,In_297,In_1210);
and U2815 (N_2815,In_531,In_1384);
or U2816 (N_2816,In_1401,In_963);
or U2817 (N_2817,In_1666,In_370);
and U2818 (N_2818,In_59,In_1496);
nor U2819 (N_2819,In_780,In_1982);
nor U2820 (N_2820,In_1403,In_1074);
nand U2821 (N_2821,In_582,In_852);
and U2822 (N_2822,In_1224,In_1739);
and U2823 (N_2823,In_1808,In_231);
nand U2824 (N_2824,In_174,In_643);
nor U2825 (N_2825,In_630,In_1894);
nand U2826 (N_2826,In_489,In_1050);
and U2827 (N_2827,In_1297,In_754);
nand U2828 (N_2828,In_1623,In_1052);
or U2829 (N_2829,In_1171,In_1202);
nand U2830 (N_2830,In_1343,In_528);
or U2831 (N_2831,In_1327,In_1665);
or U2832 (N_2832,In_596,In_304);
or U2833 (N_2833,In_1015,In_759);
and U2834 (N_2834,In_344,In_1963);
or U2835 (N_2835,In_866,In_1910);
xnor U2836 (N_2836,In_119,In_1013);
nand U2837 (N_2837,In_216,In_457);
and U2838 (N_2838,In_1008,In_1941);
nor U2839 (N_2839,In_1326,In_807);
nand U2840 (N_2840,In_1773,In_630);
or U2841 (N_2841,In_11,In_704);
or U2842 (N_2842,In_476,In_187);
nand U2843 (N_2843,In_958,In_1596);
nor U2844 (N_2844,In_482,In_1124);
and U2845 (N_2845,In_777,In_432);
or U2846 (N_2846,In_50,In_724);
nand U2847 (N_2847,In_80,In_1337);
nand U2848 (N_2848,In_1958,In_461);
and U2849 (N_2849,In_631,In_1334);
nand U2850 (N_2850,In_1960,In_714);
nor U2851 (N_2851,In_1857,In_34);
nor U2852 (N_2852,In_1412,In_207);
nand U2853 (N_2853,In_1302,In_811);
nor U2854 (N_2854,In_669,In_1887);
nand U2855 (N_2855,In_858,In_1232);
nand U2856 (N_2856,In_789,In_149);
or U2857 (N_2857,In_1703,In_1442);
and U2858 (N_2858,In_1171,In_119);
nand U2859 (N_2859,In_979,In_1555);
nand U2860 (N_2860,In_1685,In_996);
and U2861 (N_2861,In_1701,In_1259);
xor U2862 (N_2862,In_817,In_1635);
nand U2863 (N_2863,In_1319,In_1760);
or U2864 (N_2864,In_623,In_195);
or U2865 (N_2865,In_565,In_1938);
and U2866 (N_2866,In_1644,In_1137);
and U2867 (N_2867,In_1501,In_1065);
nor U2868 (N_2868,In_361,In_127);
and U2869 (N_2869,In_104,In_1372);
and U2870 (N_2870,In_546,In_998);
and U2871 (N_2871,In_176,In_630);
and U2872 (N_2872,In_486,In_258);
and U2873 (N_2873,In_1348,In_1715);
and U2874 (N_2874,In_1091,In_1282);
nand U2875 (N_2875,In_1885,In_586);
and U2876 (N_2876,In_731,In_436);
xnor U2877 (N_2877,In_636,In_1687);
nor U2878 (N_2878,In_1005,In_582);
or U2879 (N_2879,In_104,In_398);
and U2880 (N_2880,In_1207,In_145);
or U2881 (N_2881,In_1078,In_429);
or U2882 (N_2882,In_1125,In_236);
and U2883 (N_2883,In_1356,In_1529);
and U2884 (N_2884,In_751,In_1304);
and U2885 (N_2885,In_614,In_1400);
nand U2886 (N_2886,In_616,In_1675);
nor U2887 (N_2887,In_1067,In_689);
nand U2888 (N_2888,In_514,In_1106);
nor U2889 (N_2889,In_476,In_1955);
nand U2890 (N_2890,In_413,In_1506);
or U2891 (N_2891,In_386,In_1542);
nand U2892 (N_2892,In_1096,In_539);
and U2893 (N_2893,In_792,In_464);
nor U2894 (N_2894,In_1246,In_1971);
and U2895 (N_2895,In_1282,In_34);
nand U2896 (N_2896,In_76,In_798);
nand U2897 (N_2897,In_658,In_680);
nor U2898 (N_2898,In_1778,In_621);
and U2899 (N_2899,In_195,In_703);
nand U2900 (N_2900,In_702,In_1076);
nor U2901 (N_2901,In_897,In_296);
nor U2902 (N_2902,In_1474,In_442);
nand U2903 (N_2903,In_81,In_395);
and U2904 (N_2904,In_1589,In_1523);
nor U2905 (N_2905,In_326,In_1039);
nor U2906 (N_2906,In_1896,In_764);
nand U2907 (N_2907,In_1848,In_917);
nor U2908 (N_2908,In_1467,In_205);
and U2909 (N_2909,In_1933,In_875);
and U2910 (N_2910,In_1614,In_1715);
and U2911 (N_2911,In_1741,In_1694);
or U2912 (N_2912,In_1264,In_110);
or U2913 (N_2913,In_932,In_1611);
nand U2914 (N_2914,In_1002,In_871);
nor U2915 (N_2915,In_1572,In_1326);
nor U2916 (N_2916,In_1891,In_310);
nor U2917 (N_2917,In_487,In_257);
nor U2918 (N_2918,In_1536,In_1569);
or U2919 (N_2919,In_662,In_1296);
and U2920 (N_2920,In_642,In_1254);
nor U2921 (N_2921,In_1639,In_1158);
nand U2922 (N_2922,In_654,In_1017);
and U2923 (N_2923,In_1464,In_1301);
nand U2924 (N_2924,In_1254,In_82);
nor U2925 (N_2925,In_1140,In_434);
and U2926 (N_2926,In_580,In_1709);
and U2927 (N_2927,In_1967,In_548);
and U2928 (N_2928,In_531,In_350);
nor U2929 (N_2929,In_903,In_963);
nand U2930 (N_2930,In_372,In_1645);
and U2931 (N_2931,In_1721,In_334);
and U2932 (N_2932,In_1160,In_300);
and U2933 (N_2933,In_1136,In_427);
nand U2934 (N_2934,In_1595,In_1089);
or U2935 (N_2935,In_1075,In_268);
nor U2936 (N_2936,In_764,In_217);
nand U2937 (N_2937,In_483,In_1993);
or U2938 (N_2938,In_739,In_453);
nor U2939 (N_2939,In_1850,In_1987);
nand U2940 (N_2940,In_1363,In_847);
nand U2941 (N_2941,In_1347,In_637);
and U2942 (N_2942,In_683,In_1101);
nor U2943 (N_2943,In_308,In_1008);
or U2944 (N_2944,In_451,In_962);
nor U2945 (N_2945,In_1257,In_1043);
and U2946 (N_2946,In_209,In_1719);
or U2947 (N_2947,In_777,In_495);
nand U2948 (N_2948,In_1403,In_1834);
or U2949 (N_2949,In_1514,In_962);
and U2950 (N_2950,In_1569,In_1295);
nor U2951 (N_2951,In_1144,In_1559);
nor U2952 (N_2952,In_1449,In_808);
nor U2953 (N_2953,In_279,In_897);
and U2954 (N_2954,In_1060,In_1156);
and U2955 (N_2955,In_1163,In_921);
and U2956 (N_2956,In_1618,In_404);
nor U2957 (N_2957,In_931,In_482);
nor U2958 (N_2958,In_1168,In_941);
and U2959 (N_2959,In_540,In_721);
nor U2960 (N_2960,In_565,In_1617);
nand U2961 (N_2961,In_436,In_545);
nor U2962 (N_2962,In_469,In_316);
and U2963 (N_2963,In_719,In_1709);
xnor U2964 (N_2964,In_631,In_330);
and U2965 (N_2965,In_1788,In_50);
and U2966 (N_2966,In_1503,In_8);
nor U2967 (N_2967,In_701,In_66);
or U2968 (N_2968,In_1168,In_731);
nor U2969 (N_2969,In_1543,In_1724);
nor U2970 (N_2970,In_1918,In_1745);
nand U2971 (N_2971,In_353,In_1042);
and U2972 (N_2972,In_1809,In_1044);
nor U2973 (N_2973,In_679,In_360);
or U2974 (N_2974,In_1536,In_688);
and U2975 (N_2975,In_292,In_1305);
nor U2976 (N_2976,In_1002,In_730);
nor U2977 (N_2977,In_910,In_600);
and U2978 (N_2978,In_1201,In_1474);
nand U2979 (N_2979,In_860,In_1830);
or U2980 (N_2980,In_860,In_684);
nor U2981 (N_2981,In_259,In_503);
or U2982 (N_2982,In_399,In_1923);
nand U2983 (N_2983,In_827,In_492);
nor U2984 (N_2984,In_716,In_1483);
nand U2985 (N_2985,In_672,In_1994);
or U2986 (N_2986,In_439,In_1453);
and U2987 (N_2987,In_683,In_1323);
or U2988 (N_2988,In_383,In_1123);
or U2989 (N_2989,In_1358,In_687);
and U2990 (N_2990,In_995,In_909);
or U2991 (N_2991,In_1533,In_725);
or U2992 (N_2992,In_71,In_1270);
nand U2993 (N_2993,In_465,In_1103);
nor U2994 (N_2994,In_1282,In_1817);
nand U2995 (N_2995,In_804,In_1147);
nand U2996 (N_2996,In_973,In_775);
nand U2997 (N_2997,In_1737,In_1047);
nor U2998 (N_2998,In_1329,In_878);
and U2999 (N_2999,In_427,In_1309);
nand U3000 (N_3000,In_710,In_275);
or U3001 (N_3001,In_1124,In_82);
nor U3002 (N_3002,In_36,In_682);
nor U3003 (N_3003,In_1651,In_1337);
or U3004 (N_3004,In_20,In_375);
nor U3005 (N_3005,In_1118,In_494);
and U3006 (N_3006,In_1262,In_1448);
and U3007 (N_3007,In_1971,In_861);
nor U3008 (N_3008,In_1476,In_205);
nand U3009 (N_3009,In_391,In_1439);
nor U3010 (N_3010,In_443,In_22);
nor U3011 (N_3011,In_1308,In_136);
nor U3012 (N_3012,In_1619,In_1310);
nand U3013 (N_3013,In_668,In_1720);
and U3014 (N_3014,In_935,In_726);
and U3015 (N_3015,In_1141,In_600);
and U3016 (N_3016,In_152,In_842);
and U3017 (N_3017,In_1484,In_1908);
nand U3018 (N_3018,In_1218,In_299);
nand U3019 (N_3019,In_639,In_424);
nand U3020 (N_3020,In_451,In_694);
or U3021 (N_3021,In_1601,In_1588);
and U3022 (N_3022,In_136,In_1687);
or U3023 (N_3023,In_1613,In_1705);
and U3024 (N_3024,In_1044,In_674);
nand U3025 (N_3025,In_1721,In_865);
nand U3026 (N_3026,In_825,In_122);
and U3027 (N_3027,In_1547,In_1474);
or U3028 (N_3028,In_646,In_1461);
and U3029 (N_3029,In_1940,In_1765);
nor U3030 (N_3030,In_301,In_927);
nor U3031 (N_3031,In_791,In_1375);
nor U3032 (N_3032,In_828,In_699);
nand U3033 (N_3033,In_361,In_1746);
or U3034 (N_3034,In_940,In_1704);
and U3035 (N_3035,In_652,In_1596);
and U3036 (N_3036,In_1398,In_615);
or U3037 (N_3037,In_1876,In_98);
or U3038 (N_3038,In_204,In_1604);
nand U3039 (N_3039,In_117,In_1910);
or U3040 (N_3040,In_1961,In_1735);
and U3041 (N_3041,In_1180,In_1857);
nand U3042 (N_3042,In_744,In_717);
nand U3043 (N_3043,In_1667,In_1904);
and U3044 (N_3044,In_1845,In_639);
nor U3045 (N_3045,In_1522,In_964);
nand U3046 (N_3046,In_18,In_1417);
or U3047 (N_3047,In_1381,In_1477);
nor U3048 (N_3048,In_1655,In_33);
or U3049 (N_3049,In_1665,In_1516);
or U3050 (N_3050,In_227,In_896);
nor U3051 (N_3051,In_1154,In_169);
or U3052 (N_3052,In_1294,In_1085);
and U3053 (N_3053,In_71,In_1125);
nand U3054 (N_3054,In_1213,In_1003);
nand U3055 (N_3055,In_15,In_1410);
nand U3056 (N_3056,In_154,In_1284);
and U3057 (N_3057,In_972,In_1419);
or U3058 (N_3058,In_1160,In_1999);
nor U3059 (N_3059,In_589,In_1758);
and U3060 (N_3060,In_869,In_1508);
or U3061 (N_3061,In_1348,In_1980);
nor U3062 (N_3062,In_1031,In_30);
and U3063 (N_3063,In_1701,In_637);
nand U3064 (N_3064,In_1207,In_178);
or U3065 (N_3065,In_941,In_1000);
nand U3066 (N_3066,In_1893,In_1132);
nor U3067 (N_3067,In_862,In_1081);
and U3068 (N_3068,In_1977,In_139);
or U3069 (N_3069,In_1346,In_1899);
or U3070 (N_3070,In_310,In_431);
nand U3071 (N_3071,In_1631,In_1560);
or U3072 (N_3072,In_1392,In_975);
or U3073 (N_3073,In_1930,In_114);
and U3074 (N_3074,In_405,In_563);
nor U3075 (N_3075,In_801,In_1365);
and U3076 (N_3076,In_86,In_1749);
nor U3077 (N_3077,In_1667,In_278);
nand U3078 (N_3078,In_419,In_1667);
nand U3079 (N_3079,In_710,In_497);
and U3080 (N_3080,In_1064,In_184);
and U3081 (N_3081,In_930,In_666);
nor U3082 (N_3082,In_165,In_82);
nor U3083 (N_3083,In_1463,In_1330);
and U3084 (N_3084,In_331,In_507);
nand U3085 (N_3085,In_696,In_1300);
nand U3086 (N_3086,In_1455,In_1340);
or U3087 (N_3087,In_1678,In_1644);
and U3088 (N_3088,In_1549,In_1681);
nand U3089 (N_3089,In_185,In_442);
and U3090 (N_3090,In_1709,In_1433);
or U3091 (N_3091,In_1292,In_1420);
nor U3092 (N_3092,In_1483,In_1755);
or U3093 (N_3093,In_1936,In_542);
nor U3094 (N_3094,In_198,In_853);
and U3095 (N_3095,In_564,In_1599);
nor U3096 (N_3096,In_492,In_134);
or U3097 (N_3097,In_1153,In_605);
nor U3098 (N_3098,In_1153,In_670);
nand U3099 (N_3099,In_1989,In_1629);
and U3100 (N_3100,In_1833,In_1276);
nor U3101 (N_3101,In_22,In_472);
and U3102 (N_3102,In_654,In_1815);
nand U3103 (N_3103,In_1064,In_1132);
nor U3104 (N_3104,In_1623,In_1844);
nor U3105 (N_3105,In_1095,In_180);
or U3106 (N_3106,In_1898,In_787);
or U3107 (N_3107,In_1146,In_4);
nor U3108 (N_3108,In_1522,In_268);
nor U3109 (N_3109,In_982,In_889);
and U3110 (N_3110,In_1338,In_1802);
nor U3111 (N_3111,In_103,In_819);
or U3112 (N_3112,In_730,In_807);
nor U3113 (N_3113,In_480,In_7);
and U3114 (N_3114,In_853,In_533);
nand U3115 (N_3115,In_986,In_339);
and U3116 (N_3116,In_1658,In_1233);
nand U3117 (N_3117,In_1965,In_1042);
nand U3118 (N_3118,In_977,In_491);
or U3119 (N_3119,In_1563,In_364);
or U3120 (N_3120,In_930,In_1718);
nor U3121 (N_3121,In_635,In_1351);
and U3122 (N_3122,In_310,In_483);
or U3123 (N_3123,In_217,In_1199);
nor U3124 (N_3124,In_1221,In_1676);
nor U3125 (N_3125,In_255,In_443);
nor U3126 (N_3126,In_1562,In_1742);
and U3127 (N_3127,In_1085,In_1948);
and U3128 (N_3128,In_1057,In_1296);
and U3129 (N_3129,In_870,In_1128);
or U3130 (N_3130,In_1199,In_172);
and U3131 (N_3131,In_1934,In_1104);
or U3132 (N_3132,In_1710,In_506);
or U3133 (N_3133,In_1533,In_1190);
nand U3134 (N_3134,In_291,In_1475);
xor U3135 (N_3135,In_1234,In_173);
and U3136 (N_3136,In_170,In_67);
and U3137 (N_3137,In_38,In_1761);
or U3138 (N_3138,In_786,In_811);
or U3139 (N_3139,In_1516,In_411);
nand U3140 (N_3140,In_1362,In_208);
and U3141 (N_3141,In_1172,In_1994);
or U3142 (N_3142,In_1764,In_1610);
and U3143 (N_3143,In_1711,In_1431);
and U3144 (N_3144,In_249,In_773);
or U3145 (N_3145,In_839,In_1191);
nand U3146 (N_3146,In_1229,In_1739);
nor U3147 (N_3147,In_1786,In_234);
nand U3148 (N_3148,In_893,In_40);
nor U3149 (N_3149,In_981,In_1644);
or U3150 (N_3150,In_1371,In_1822);
or U3151 (N_3151,In_681,In_379);
nor U3152 (N_3152,In_1797,In_720);
and U3153 (N_3153,In_536,In_655);
or U3154 (N_3154,In_1084,In_414);
or U3155 (N_3155,In_92,In_595);
nor U3156 (N_3156,In_777,In_668);
nand U3157 (N_3157,In_369,In_112);
nor U3158 (N_3158,In_1000,In_9);
nand U3159 (N_3159,In_1947,In_761);
nor U3160 (N_3160,In_775,In_31);
nand U3161 (N_3161,In_1280,In_1801);
nand U3162 (N_3162,In_1270,In_276);
nor U3163 (N_3163,In_830,In_1815);
nand U3164 (N_3164,In_523,In_1290);
nor U3165 (N_3165,In_1365,In_527);
or U3166 (N_3166,In_937,In_8);
nor U3167 (N_3167,In_1714,In_1874);
nand U3168 (N_3168,In_1106,In_1166);
and U3169 (N_3169,In_942,In_1534);
nand U3170 (N_3170,In_1117,In_1688);
and U3171 (N_3171,In_184,In_854);
and U3172 (N_3172,In_512,In_1014);
nor U3173 (N_3173,In_106,In_1852);
or U3174 (N_3174,In_686,In_1144);
and U3175 (N_3175,In_340,In_695);
nand U3176 (N_3176,In_139,In_1997);
nand U3177 (N_3177,In_1137,In_1209);
nand U3178 (N_3178,In_780,In_1211);
nand U3179 (N_3179,In_698,In_746);
or U3180 (N_3180,In_1284,In_1583);
or U3181 (N_3181,In_728,In_1312);
nor U3182 (N_3182,In_22,In_1733);
and U3183 (N_3183,In_1312,In_605);
or U3184 (N_3184,In_1495,In_568);
or U3185 (N_3185,In_1975,In_1844);
and U3186 (N_3186,In_1858,In_40);
nand U3187 (N_3187,In_1805,In_214);
and U3188 (N_3188,In_1051,In_343);
nor U3189 (N_3189,In_635,In_154);
nand U3190 (N_3190,In_275,In_1521);
and U3191 (N_3191,In_442,In_1061);
and U3192 (N_3192,In_268,In_1632);
nand U3193 (N_3193,In_1325,In_260);
or U3194 (N_3194,In_1725,In_389);
nor U3195 (N_3195,In_805,In_497);
nand U3196 (N_3196,In_408,In_1783);
nand U3197 (N_3197,In_1975,In_1824);
or U3198 (N_3198,In_1453,In_87);
and U3199 (N_3199,In_1222,In_1998);
or U3200 (N_3200,In_206,In_1816);
nand U3201 (N_3201,In_1875,In_24);
nand U3202 (N_3202,In_1732,In_1480);
or U3203 (N_3203,In_1155,In_1640);
and U3204 (N_3204,In_1898,In_1719);
or U3205 (N_3205,In_345,In_1410);
nor U3206 (N_3206,In_1715,In_1982);
and U3207 (N_3207,In_834,In_673);
nand U3208 (N_3208,In_1881,In_1337);
or U3209 (N_3209,In_644,In_1238);
nor U3210 (N_3210,In_368,In_216);
nor U3211 (N_3211,In_245,In_985);
nor U3212 (N_3212,In_1659,In_848);
nor U3213 (N_3213,In_1781,In_199);
nor U3214 (N_3214,In_1700,In_1275);
or U3215 (N_3215,In_1420,In_481);
and U3216 (N_3216,In_1395,In_917);
or U3217 (N_3217,In_936,In_1444);
and U3218 (N_3218,In_1725,In_334);
nand U3219 (N_3219,In_1323,In_771);
nor U3220 (N_3220,In_1152,In_1843);
nand U3221 (N_3221,In_1487,In_112);
and U3222 (N_3222,In_1758,In_1935);
or U3223 (N_3223,In_371,In_1661);
nand U3224 (N_3224,In_982,In_1720);
and U3225 (N_3225,In_1078,In_1926);
nor U3226 (N_3226,In_1120,In_1874);
nand U3227 (N_3227,In_1591,In_617);
or U3228 (N_3228,In_1443,In_17);
or U3229 (N_3229,In_1124,In_1263);
xor U3230 (N_3230,In_853,In_620);
and U3231 (N_3231,In_1540,In_433);
nor U3232 (N_3232,In_831,In_916);
nand U3233 (N_3233,In_593,In_1914);
and U3234 (N_3234,In_785,In_994);
and U3235 (N_3235,In_1426,In_271);
nand U3236 (N_3236,In_1087,In_250);
or U3237 (N_3237,In_527,In_1654);
or U3238 (N_3238,In_261,In_1786);
nor U3239 (N_3239,In_1182,In_1498);
nand U3240 (N_3240,In_1929,In_1460);
nand U3241 (N_3241,In_1021,In_1819);
or U3242 (N_3242,In_465,In_1134);
nand U3243 (N_3243,In_1396,In_1457);
or U3244 (N_3244,In_1436,In_1782);
or U3245 (N_3245,In_95,In_1083);
or U3246 (N_3246,In_1706,In_1039);
or U3247 (N_3247,In_544,In_1283);
and U3248 (N_3248,In_384,In_716);
nor U3249 (N_3249,In_682,In_48);
and U3250 (N_3250,In_556,In_839);
or U3251 (N_3251,In_1650,In_57);
or U3252 (N_3252,In_281,In_1039);
nand U3253 (N_3253,In_1815,In_126);
or U3254 (N_3254,In_552,In_1280);
or U3255 (N_3255,In_1444,In_508);
or U3256 (N_3256,In_1506,In_856);
or U3257 (N_3257,In_1419,In_848);
nor U3258 (N_3258,In_1759,In_1123);
nor U3259 (N_3259,In_232,In_1301);
nor U3260 (N_3260,In_1787,In_1062);
and U3261 (N_3261,In_1236,In_1151);
nor U3262 (N_3262,In_989,In_1172);
nor U3263 (N_3263,In_1494,In_1737);
and U3264 (N_3264,In_1712,In_177);
or U3265 (N_3265,In_1288,In_598);
nor U3266 (N_3266,In_493,In_1044);
and U3267 (N_3267,In_504,In_279);
nand U3268 (N_3268,In_1718,In_1793);
or U3269 (N_3269,In_1297,In_420);
nand U3270 (N_3270,In_114,In_1583);
and U3271 (N_3271,In_1513,In_1751);
and U3272 (N_3272,In_220,In_1564);
nor U3273 (N_3273,In_238,In_178);
or U3274 (N_3274,In_996,In_405);
nor U3275 (N_3275,In_1430,In_84);
nor U3276 (N_3276,In_1291,In_432);
or U3277 (N_3277,In_1555,In_1363);
and U3278 (N_3278,In_1599,In_895);
nand U3279 (N_3279,In_1689,In_1126);
or U3280 (N_3280,In_702,In_444);
or U3281 (N_3281,In_1768,In_1355);
nand U3282 (N_3282,In_690,In_1220);
nand U3283 (N_3283,In_1513,In_337);
nor U3284 (N_3284,In_1161,In_323);
nor U3285 (N_3285,In_491,In_1565);
nand U3286 (N_3286,In_1602,In_1327);
nor U3287 (N_3287,In_1142,In_115);
nor U3288 (N_3288,In_739,In_78);
nand U3289 (N_3289,In_1101,In_1743);
nand U3290 (N_3290,In_191,In_1836);
nor U3291 (N_3291,In_401,In_1938);
nor U3292 (N_3292,In_444,In_728);
or U3293 (N_3293,In_1563,In_1911);
or U3294 (N_3294,In_1309,In_1561);
and U3295 (N_3295,In_1949,In_800);
nor U3296 (N_3296,In_282,In_1410);
nor U3297 (N_3297,In_1826,In_942);
nand U3298 (N_3298,In_1040,In_171);
or U3299 (N_3299,In_51,In_1580);
and U3300 (N_3300,In_1858,In_528);
nor U3301 (N_3301,In_1620,In_1722);
nand U3302 (N_3302,In_600,In_451);
nand U3303 (N_3303,In_1366,In_593);
nand U3304 (N_3304,In_849,In_1663);
or U3305 (N_3305,In_656,In_55);
or U3306 (N_3306,In_280,In_1175);
nand U3307 (N_3307,In_1289,In_1817);
and U3308 (N_3308,In_1363,In_995);
or U3309 (N_3309,In_877,In_341);
and U3310 (N_3310,In_577,In_292);
or U3311 (N_3311,In_349,In_238);
and U3312 (N_3312,In_1420,In_1698);
and U3313 (N_3313,In_1115,In_1513);
nor U3314 (N_3314,In_706,In_1709);
and U3315 (N_3315,In_1659,In_345);
and U3316 (N_3316,In_1182,In_1321);
or U3317 (N_3317,In_1169,In_342);
or U3318 (N_3318,In_998,In_563);
xor U3319 (N_3319,In_368,In_478);
nor U3320 (N_3320,In_1145,In_614);
nor U3321 (N_3321,In_1935,In_1728);
nand U3322 (N_3322,In_256,In_856);
nor U3323 (N_3323,In_1261,In_255);
nor U3324 (N_3324,In_1224,In_1081);
and U3325 (N_3325,In_58,In_429);
nand U3326 (N_3326,In_150,In_1024);
nor U3327 (N_3327,In_1789,In_1597);
nand U3328 (N_3328,In_737,In_82);
nand U3329 (N_3329,In_1491,In_1116);
nand U3330 (N_3330,In_737,In_1194);
and U3331 (N_3331,In_705,In_1290);
nor U3332 (N_3332,In_625,In_286);
nand U3333 (N_3333,In_1845,In_1227);
or U3334 (N_3334,In_1592,In_874);
nand U3335 (N_3335,In_1594,In_1370);
or U3336 (N_3336,In_375,In_1797);
or U3337 (N_3337,In_310,In_1708);
or U3338 (N_3338,In_677,In_760);
or U3339 (N_3339,In_1430,In_1208);
and U3340 (N_3340,In_427,In_1696);
nand U3341 (N_3341,In_357,In_1359);
and U3342 (N_3342,In_904,In_1673);
or U3343 (N_3343,In_1848,In_849);
nand U3344 (N_3344,In_444,In_1690);
or U3345 (N_3345,In_464,In_861);
and U3346 (N_3346,In_1628,In_1041);
or U3347 (N_3347,In_1586,In_305);
or U3348 (N_3348,In_1439,In_1670);
or U3349 (N_3349,In_1398,In_1146);
or U3350 (N_3350,In_1511,In_698);
nand U3351 (N_3351,In_343,In_987);
and U3352 (N_3352,In_1919,In_800);
or U3353 (N_3353,In_1970,In_1921);
and U3354 (N_3354,In_1047,In_1005);
and U3355 (N_3355,In_11,In_830);
and U3356 (N_3356,In_65,In_1767);
or U3357 (N_3357,In_1649,In_373);
or U3358 (N_3358,In_665,In_119);
and U3359 (N_3359,In_1491,In_662);
nor U3360 (N_3360,In_1751,In_688);
nor U3361 (N_3361,In_1235,In_608);
nand U3362 (N_3362,In_788,In_652);
and U3363 (N_3363,In_1767,In_505);
nand U3364 (N_3364,In_1585,In_1056);
nand U3365 (N_3365,In_1442,In_1848);
nand U3366 (N_3366,In_110,In_471);
and U3367 (N_3367,In_207,In_219);
or U3368 (N_3368,In_1966,In_1883);
nand U3369 (N_3369,In_1135,In_1567);
nor U3370 (N_3370,In_425,In_1766);
nor U3371 (N_3371,In_974,In_718);
nand U3372 (N_3372,In_1095,In_793);
and U3373 (N_3373,In_679,In_504);
or U3374 (N_3374,In_139,In_1625);
and U3375 (N_3375,In_1386,In_96);
or U3376 (N_3376,In_1329,In_481);
and U3377 (N_3377,In_278,In_1911);
nand U3378 (N_3378,In_998,In_1443);
nand U3379 (N_3379,In_300,In_277);
nand U3380 (N_3380,In_344,In_1863);
and U3381 (N_3381,In_522,In_767);
or U3382 (N_3382,In_1296,In_1628);
and U3383 (N_3383,In_1153,In_1738);
and U3384 (N_3384,In_1638,In_786);
nand U3385 (N_3385,In_1840,In_1393);
or U3386 (N_3386,In_397,In_883);
or U3387 (N_3387,In_1199,In_277);
nor U3388 (N_3388,In_1802,In_589);
nor U3389 (N_3389,In_1757,In_1726);
and U3390 (N_3390,In_1585,In_361);
or U3391 (N_3391,In_897,In_1659);
nand U3392 (N_3392,In_1224,In_1581);
or U3393 (N_3393,In_755,In_653);
nand U3394 (N_3394,In_1564,In_724);
nand U3395 (N_3395,In_54,In_13);
nand U3396 (N_3396,In_973,In_1834);
nand U3397 (N_3397,In_1203,In_452);
nor U3398 (N_3398,In_1739,In_521);
and U3399 (N_3399,In_1928,In_1154);
nor U3400 (N_3400,In_342,In_865);
or U3401 (N_3401,In_1657,In_312);
or U3402 (N_3402,In_1583,In_233);
nor U3403 (N_3403,In_1532,In_696);
nand U3404 (N_3404,In_372,In_1301);
and U3405 (N_3405,In_1043,In_1016);
and U3406 (N_3406,In_1786,In_401);
nand U3407 (N_3407,In_73,In_1571);
nand U3408 (N_3408,In_1431,In_1595);
nor U3409 (N_3409,In_1954,In_471);
nand U3410 (N_3410,In_769,In_1604);
or U3411 (N_3411,In_512,In_1681);
nand U3412 (N_3412,In_1047,In_1748);
and U3413 (N_3413,In_1476,In_1639);
or U3414 (N_3414,In_931,In_855);
nand U3415 (N_3415,In_1599,In_1658);
xor U3416 (N_3416,In_124,In_527);
nor U3417 (N_3417,In_1951,In_1359);
and U3418 (N_3418,In_1179,In_836);
nor U3419 (N_3419,In_389,In_311);
nor U3420 (N_3420,In_406,In_1346);
and U3421 (N_3421,In_842,In_784);
and U3422 (N_3422,In_1800,In_675);
xnor U3423 (N_3423,In_1683,In_62);
and U3424 (N_3424,In_632,In_1912);
and U3425 (N_3425,In_1536,In_1283);
and U3426 (N_3426,In_174,In_523);
and U3427 (N_3427,In_1447,In_1584);
nand U3428 (N_3428,In_41,In_53);
or U3429 (N_3429,In_335,In_1197);
and U3430 (N_3430,In_1468,In_1983);
and U3431 (N_3431,In_1072,In_1945);
nor U3432 (N_3432,In_240,In_1868);
nor U3433 (N_3433,In_1313,In_1147);
or U3434 (N_3434,In_1042,In_1770);
and U3435 (N_3435,In_1972,In_1974);
nor U3436 (N_3436,In_1112,In_289);
or U3437 (N_3437,In_78,In_1372);
nand U3438 (N_3438,In_453,In_83);
and U3439 (N_3439,In_1740,In_610);
or U3440 (N_3440,In_240,In_1293);
nor U3441 (N_3441,In_1115,In_211);
nor U3442 (N_3442,In_364,In_1722);
nand U3443 (N_3443,In_246,In_159);
nor U3444 (N_3444,In_1937,In_1622);
nor U3445 (N_3445,In_869,In_394);
or U3446 (N_3446,In_1743,In_761);
nor U3447 (N_3447,In_1414,In_1675);
and U3448 (N_3448,In_814,In_1507);
or U3449 (N_3449,In_88,In_702);
and U3450 (N_3450,In_1515,In_691);
nand U3451 (N_3451,In_1013,In_649);
or U3452 (N_3452,In_1585,In_1602);
xnor U3453 (N_3453,In_1360,In_360);
xor U3454 (N_3454,In_245,In_1284);
or U3455 (N_3455,In_138,In_432);
and U3456 (N_3456,In_1394,In_1493);
or U3457 (N_3457,In_1439,In_634);
nor U3458 (N_3458,In_686,In_1242);
nand U3459 (N_3459,In_1286,In_1895);
nor U3460 (N_3460,In_35,In_196);
or U3461 (N_3461,In_1209,In_143);
and U3462 (N_3462,In_981,In_1036);
nor U3463 (N_3463,In_267,In_785);
nand U3464 (N_3464,In_1800,In_1289);
or U3465 (N_3465,In_1293,In_722);
nand U3466 (N_3466,In_166,In_1163);
or U3467 (N_3467,In_236,In_116);
nor U3468 (N_3468,In_206,In_1877);
or U3469 (N_3469,In_306,In_727);
or U3470 (N_3470,In_589,In_230);
nor U3471 (N_3471,In_427,In_726);
or U3472 (N_3472,In_381,In_690);
nand U3473 (N_3473,In_238,In_1682);
and U3474 (N_3474,In_1651,In_217);
nand U3475 (N_3475,In_1930,In_1922);
and U3476 (N_3476,In_914,In_1582);
nor U3477 (N_3477,In_1887,In_1700);
nor U3478 (N_3478,In_827,In_1383);
nor U3479 (N_3479,In_1710,In_1711);
and U3480 (N_3480,In_523,In_212);
or U3481 (N_3481,In_451,In_1284);
nand U3482 (N_3482,In_277,In_1365);
nor U3483 (N_3483,In_796,In_179);
nor U3484 (N_3484,In_1577,In_1622);
nor U3485 (N_3485,In_1400,In_1949);
or U3486 (N_3486,In_1055,In_1513);
and U3487 (N_3487,In_571,In_326);
xor U3488 (N_3488,In_701,In_1645);
or U3489 (N_3489,In_673,In_335);
and U3490 (N_3490,In_107,In_162);
and U3491 (N_3491,In_896,In_1895);
nor U3492 (N_3492,In_834,In_1638);
and U3493 (N_3493,In_1357,In_475);
nand U3494 (N_3494,In_802,In_1210);
and U3495 (N_3495,In_531,In_842);
and U3496 (N_3496,In_1552,In_1466);
xor U3497 (N_3497,In_336,In_1739);
nor U3498 (N_3498,In_618,In_1072);
or U3499 (N_3499,In_1964,In_258);
nor U3500 (N_3500,In_747,In_1581);
nor U3501 (N_3501,In_1978,In_1973);
or U3502 (N_3502,In_1415,In_1850);
or U3503 (N_3503,In_1503,In_1034);
nand U3504 (N_3504,In_696,In_454);
and U3505 (N_3505,In_1916,In_1339);
and U3506 (N_3506,In_549,In_1181);
nor U3507 (N_3507,In_1910,In_1566);
or U3508 (N_3508,In_630,In_907);
and U3509 (N_3509,In_745,In_988);
nand U3510 (N_3510,In_752,In_463);
nor U3511 (N_3511,In_777,In_866);
and U3512 (N_3512,In_1179,In_716);
nand U3513 (N_3513,In_1818,In_409);
nand U3514 (N_3514,In_1855,In_417);
nand U3515 (N_3515,In_538,In_564);
nor U3516 (N_3516,In_1527,In_965);
and U3517 (N_3517,In_2,In_348);
and U3518 (N_3518,In_1694,In_41);
or U3519 (N_3519,In_1858,In_1414);
nor U3520 (N_3520,In_1099,In_99);
nor U3521 (N_3521,In_165,In_107);
nand U3522 (N_3522,In_1924,In_139);
nand U3523 (N_3523,In_1072,In_1224);
or U3524 (N_3524,In_553,In_1123);
nor U3525 (N_3525,In_695,In_1262);
or U3526 (N_3526,In_1759,In_1518);
nand U3527 (N_3527,In_1322,In_915);
and U3528 (N_3528,In_1388,In_1204);
or U3529 (N_3529,In_432,In_1015);
or U3530 (N_3530,In_1803,In_101);
nor U3531 (N_3531,In_853,In_763);
nand U3532 (N_3532,In_1930,In_1377);
nand U3533 (N_3533,In_71,In_708);
nor U3534 (N_3534,In_814,In_1814);
and U3535 (N_3535,In_1177,In_356);
nor U3536 (N_3536,In_1060,In_1341);
nor U3537 (N_3537,In_628,In_329);
and U3538 (N_3538,In_1992,In_1462);
nor U3539 (N_3539,In_1570,In_345);
and U3540 (N_3540,In_1590,In_794);
nor U3541 (N_3541,In_1058,In_736);
and U3542 (N_3542,In_674,In_783);
or U3543 (N_3543,In_1607,In_1441);
nor U3544 (N_3544,In_1740,In_975);
or U3545 (N_3545,In_1976,In_1345);
nor U3546 (N_3546,In_881,In_689);
nor U3547 (N_3547,In_154,In_1977);
nor U3548 (N_3548,In_128,In_716);
nand U3549 (N_3549,In_1564,In_922);
nand U3550 (N_3550,In_616,In_295);
nand U3551 (N_3551,In_1896,In_54);
or U3552 (N_3552,In_1273,In_1511);
nor U3553 (N_3553,In_1797,In_586);
or U3554 (N_3554,In_1336,In_406);
or U3555 (N_3555,In_1952,In_1959);
or U3556 (N_3556,In_968,In_1101);
nand U3557 (N_3557,In_1042,In_275);
and U3558 (N_3558,In_722,In_1807);
or U3559 (N_3559,In_902,In_1102);
or U3560 (N_3560,In_958,In_61);
and U3561 (N_3561,In_431,In_1588);
and U3562 (N_3562,In_250,In_1663);
and U3563 (N_3563,In_915,In_1833);
nor U3564 (N_3564,In_428,In_1786);
nor U3565 (N_3565,In_1193,In_429);
nand U3566 (N_3566,In_1176,In_1931);
and U3567 (N_3567,In_1965,In_243);
or U3568 (N_3568,In_1431,In_1581);
or U3569 (N_3569,In_792,In_1205);
nand U3570 (N_3570,In_631,In_1045);
and U3571 (N_3571,In_1011,In_1410);
or U3572 (N_3572,In_1861,In_610);
nor U3573 (N_3573,In_1255,In_1346);
and U3574 (N_3574,In_192,In_1952);
nor U3575 (N_3575,In_722,In_913);
and U3576 (N_3576,In_513,In_798);
or U3577 (N_3577,In_1426,In_849);
nor U3578 (N_3578,In_1698,In_1760);
or U3579 (N_3579,In_346,In_1383);
nor U3580 (N_3580,In_1077,In_1337);
and U3581 (N_3581,In_1186,In_1537);
xnor U3582 (N_3582,In_413,In_36);
and U3583 (N_3583,In_101,In_888);
nor U3584 (N_3584,In_1865,In_1807);
nor U3585 (N_3585,In_1071,In_822);
and U3586 (N_3586,In_121,In_1633);
or U3587 (N_3587,In_451,In_781);
nand U3588 (N_3588,In_1290,In_542);
or U3589 (N_3589,In_1211,In_93);
nor U3590 (N_3590,In_663,In_937);
or U3591 (N_3591,In_17,In_1252);
nand U3592 (N_3592,In_1840,In_1054);
or U3593 (N_3593,In_847,In_1677);
and U3594 (N_3594,In_877,In_1390);
nand U3595 (N_3595,In_68,In_1585);
and U3596 (N_3596,In_1006,In_411);
nand U3597 (N_3597,In_646,In_842);
nand U3598 (N_3598,In_1022,In_1269);
or U3599 (N_3599,In_929,In_172);
and U3600 (N_3600,In_1637,In_1757);
nand U3601 (N_3601,In_1233,In_1642);
nand U3602 (N_3602,In_850,In_725);
or U3603 (N_3603,In_295,In_227);
nor U3604 (N_3604,In_1442,In_1069);
nand U3605 (N_3605,In_1518,In_1934);
and U3606 (N_3606,In_615,In_1745);
nor U3607 (N_3607,In_120,In_442);
or U3608 (N_3608,In_912,In_1929);
nor U3609 (N_3609,In_541,In_1385);
or U3610 (N_3610,In_975,In_1841);
or U3611 (N_3611,In_1467,In_1705);
nand U3612 (N_3612,In_1809,In_284);
nand U3613 (N_3613,In_1641,In_1943);
or U3614 (N_3614,In_726,In_1914);
nand U3615 (N_3615,In_678,In_1303);
or U3616 (N_3616,In_1513,In_1850);
nand U3617 (N_3617,In_845,In_1891);
and U3618 (N_3618,In_622,In_1368);
nand U3619 (N_3619,In_1387,In_1758);
or U3620 (N_3620,In_1890,In_500);
nand U3621 (N_3621,In_120,In_4);
and U3622 (N_3622,In_1078,In_162);
nor U3623 (N_3623,In_1262,In_79);
nor U3624 (N_3624,In_1889,In_1638);
or U3625 (N_3625,In_1590,In_674);
or U3626 (N_3626,In_1613,In_50);
nand U3627 (N_3627,In_1456,In_1512);
and U3628 (N_3628,In_1147,In_645);
and U3629 (N_3629,In_918,In_1424);
nand U3630 (N_3630,In_1874,In_864);
nor U3631 (N_3631,In_771,In_480);
nand U3632 (N_3632,In_449,In_287);
and U3633 (N_3633,In_588,In_1528);
or U3634 (N_3634,In_40,In_370);
and U3635 (N_3635,In_713,In_314);
nor U3636 (N_3636,In_123,In_1326);
or U3637 (N_3637,In_1035,In_1050);
or U3638 (N_3638,In_1368,In_658);
and U3639 (N_3639,In_687,In_1073);
nand U3640 (N_3640,In_285,In_1760);
or U3641 (N_3641,In_1468,In_650);
and U3642 (N_3642,In_128,In_1514);
or U3643 (N_3643,In_1184,In_1340);
and U3644 (N_3644,In_719,In_378);
nand U3645 (N_3645,In_835,In_1394);
or U3646 (N_3646,In_1948,In_1372);
or U3647 (N_3647,In_930,In_515);
nor U3648 (N_3648,In_181,In_113);
and U3649 (N_3649,In_457,In_1904);
and U3650 (N_3650,In_1570,In_939);
or U3651 (N_3651,In_555,In_1211);
or U3652 (N_3652,In_404,In_1605);
or U3653 (N_3653,In_1152,In_1625);
nor U3654 (N_3654,In_623,In_1877);
nand U3655 (N_3655,In_1451,In_1190);
nor U3656 (N_3656,In_1036,In_1310);
nand U3657 (N_3657,In_1073,In_1784);
nand U3658 (N_3658,In_210,In_1762);
nor U3659 (N_3659,In_1977,In_1900);
and U3660 (N_3660,In_319,In_1473);
nand U3661 (N_3661,In_1849,In_890);
nor U3662 (N_3662,In_1568,In_1706);
and U3663 (N_3663,In_1354,In_973);
or U3664 (N_3664,In_667,In_198);
nor U3665 (N_3665,In_1239,In_1944);
nand U3666 (N_3666,In_1454,In_1098);
xor U3667 (N_3667,In_1074,In_1757);
and U3668 (N_3668,In_719,In_1054);
nand U3669 (N_3669,In_34,In_1793);
nor U3670 (N_3670,In_123,In_1478);
and U3671 (N_3671,In_1909,In_1029);
nand U3672 (N_3672,In_1668,In_1096);
or U3673 (N_3673,In_1099,In_1156);
or U3674 (N_3674,In_772,In_1230);
nor U3675 (N_3675,In_360,In_639);
and U3676 (N_3676,In_802,In_1565);
nand U3677 (N_3677,In_1037,In_1251);
nor U3678 (N_3678,In_1788,In_501);
or U3679 (N_3679,In_1798,In_56);
nor U3680 (N_3680,In_103,In_1156);
or U3681 (N_3681,In_1086,In_1085);
nor U3682 (N_3682,In_1012,In_1959);
and U3683 (N_3683,In_965,In_235);
nand U3684 (N_3684,In_379,In_12);
and U3685 (N_3685,In_1015,In_948);
or U3686 (N_3686,In_1173,In_561);
or U3687 (N_3687,In_22,In_380);
or U3688 (N_3688,In_381,In_327);
nor U3689 (N_3689,In_818,In_0);
and U3690 (N_3690,In_1614,In_1241);
and U3691 (N_3691,In_1457,In_15);
and U3692 (N_3692,In_919,In_1304);
or U3693 (N_3693,In_689,In_1242);
and U3694 (N_3694,In_15,In_857);
nand U3695 (N_3695,In_517,In_1119);
nand U3696 (N_3696,In_734,In_285);
and U3697 (N_3697,In_476,In_1284);
nor U3698 (N_3698,In_1741,In_898);
nand U3699 (N_3699,In_1268,In_882);
nand U3700 (N_3700,In_199,In_1169);
nor U3701 (N_3701,In_958,In_1722);
nor U3702 (N_3702,In_1577,In_1286);
and U3703 (N_3703,In_1817,In_1740);
and U3704 (N_3704,In_1798,In_620);
and U3705 (N_3705,In_1948,In_1128);
or U3706 (N_3706,In_527,In_1724);
and U3707 (N_3707,In_1284,In_877);
or U3708 (N_3708,In_1111,In_353);
nand U3709 (N_3709,In_1807,In_532);
nand U3710 (N_3710,In_1770,In_1124);
and U3711 (N_3711,In_220,In_1420);
nand U3712 (N_3712,In_1487,In_1439);
xnor U3713 (N_3713,In_973,In_1185);
nand U3714 (N_3714,In_1884,In_1118);
or U3715 (N_3715,In_392,In_74);
nor U3716 (N_3716,In_1844,In_430);
nand U3717 (N_3717,In_1625,In_146);
nor U3718 (N_3718,In_495,In_1051);
and U3719 (N_3719,In_1866,In_917);
xor U3720 (N_3720,In_1692,In_1986);
nor U3721 (N_3721,In_1040,In_204);
or U3722 (N_3722,In_971,In_697);
and U3723 (N_3723,In_1022,In_1561);
nor U3724 (N_3724,In_1872,In_441);
nor U3725 (N_3725,In_544,In_135);
nor U3726 (N_3726,In_869,In_990);
or U3727 (N_3727,In_26,In_1122);
and U3728 (N_3728,In_1205,In_29);
or U3729 (N_3729,In_836,In_436);
nor U3730 (N_3730,In_1347,In_728);
or U3731 (N_3731,In_94,In_1122);
and U3732 (N_3732,In_66,In_212);
nand U3733 (N_3733,In_1657,In_1185);
nor U3734 (N_3734,In_439,In_1475);
or U3735 (N_3735,In_1124,In_162);
and U3736 (N_3736,In_1076,In_205);
nor U3737 (N_3737,In_236,In_1059);
nor U3738 (N_3738,In_337,In_316);
nand U3739 (N_3739,In_1573,In_459);
or U3740 (N_3740,In_851,In_95);
nand U3741 (N_3741,In_1442,In_837);
nor U3742 (N_3742,In_411,In_1332);
and U3743 (N_3743,In_841,In_683);
nor U3744 (N_3744,In_280,In_1635);
and U3745 (N_3745,In_942,In_927);
nor U3746 (N_3746,In_1892,In_408);
nor U3747 (N_3747,In_1100,In_481);
or U3748 (N_3748,In_68,In_1804);
nand U3749 (N_3749,In_1634,In_1224);
and U3750 (N_3750,In_860,In_957);
nand U3751 (N_3751,In_947,In_112);
or U3752 (N_3752,In_1384,In_780);
or U3753 (N_3753,In_1761,In_1620);
nand U3754 (N_3754,In_1915,In_833);
and U3755 (N_3755,In_81,In_107);
nand U3756 (N_3756,In_875,In_915);
or U3757 (N_3757,In_396,In_207);
nand U3758 (N_3758,In_118,In_1087);
nand U3759 (N_3759,In_580,In_313);
nand U3760 (N_3760,In_1029,In_1267);
or U3761 (N_3761,In_563,In_1424);
nand U3762 (N_3762,In_1561,In_1748);
nor U3763 (N_3763,In_1996,In_1385);
nor U3764 (N_3764,In_1871,In_1103);
or U3765 (N_3765,In_88,In_300);
and U3766 (N_3766,In_1467,In_188);
and U3767 (N_3767,In_1614,In_1340);
nand U3768 (N_3768,In_1264,In_1901);
and U3769 (N_3769,In_370,In_1007);
and U3770 (N_3770,In_231,In_890);
nand U3771 (N_3771,In_1442,In_1305);
nand U3772 (N_3772,In_1248,In_786);
and U3773 (N_3773,In_868,In_1098);
nand U3774 (N_3774,In_1747,In_1169);
nand U3775 (N_3775,In_1397,In_281);
and U3776 (N_3776,In_1238,In_1130);
nor U3777 (N_3777,In_516,In_1710);
nand U3778 (N_3778,In_1867,In_1420);
nor U3779 (N_3779,In_978,In_1321);
nor U3780 (N_3780,In_1297,In_896);
nor U3781 (N_3781,In_115,In_1158);
nand U3782 (N_3782,In_523,In_1916);
or U3783 (N_3783,In_157,In_1058);
nand U3784 (N_3784,In_999,In_532);
nand U3785 (N_3785,In_1343,In_888);
and U3786 (N_3786,In_865,In_1730);
or U3787 (N_3787,In_1939,In_1862);
or U3788 (N_3788,In_170,In_1205);
and U3789 (N_3789,In_1263,In_1092);
or U3790 (N_3790,In_1602,In_1678);
nor U3791 (N_3791,In_735,In_1018);
or U3792 (N_3792,In_467,In_1106);
nor U3793 (N_3793,In_1509,In_1732);
nand U3794 (N_3794,In_892,In_1710);
and U3795 (N_3795,In_292,In_1175);
nand U3796 (N_3796,In_436,In_770);
nand U3797 (N_3797,In_72,In_876);
nand U3798 (N_3798,In_1489,In_1329);
and U3799 (N_3799,In_1088,In_1386);
nand U3800 (N_3800,In_582,In_630);
and U3801 (N_3801,In_1578,In_617);
nor U3802 (N_3802,In_339,In_1806);
or U3803 (N_3803,In_1076,In_701);
and U3804 (N_3804,In_974,In_1101);
nor U3805 (N_3805,In_611,In_1155);
or U3806 (N_3806,In_1035,In_1019);
and U3807 (N_3807,In_204,In_1456);
nand U3808 (N_3808,In_991,In_533);
nor U3809 (N_3809,In_1192,In_769);
or U3810 (N_3810,In_619,In_312);
and U3811 (N_3811,In_1429,In_126);
nor U3812 (N_3812,In_725,In_622);
nor U3813 (N_3813,In_1298,In_1379);
or U3814 (N_3814,In_1065,In_1492);
nor U3815 (N_3815,In_1412,In_1893);
nor U3816 (N_3816,In_1617,In_956);
nor U3817 (N_3817,In_1267,In_227);
nand U3818 (N_3818,In_1596,In_888);
nand U3819 (N_3819,In_1200,In_75);
or U3820 (N_3820,In_145,In_1308);
nor U3821 (N_3821,In_1834,In_711);
nor U3822 (N_3822,In_636,In_1785);
nand U3823 (N_3823,In_209,In_277);
or U3824 (N_3824,In_1138,In_927);
nand U3825 (N_3825,In_1385,In_260);
nand U3826 (N_3826,In_1196,In_1890);
and U3827 (N_3827,In_968,In_892);
and U3828 (N_3828,In_253,In_594);
and U3829 (N_3829,In_683,In_285);
nor U3830 (N_3830,In_340,In_1051);
nor U3831 (N_3831,In_1442,In_725);
nand U3832 (N_3832,In_898,In_806);
and U3833 (N_3833,In_1538,In_298);
nand U3834 (N_3834,In_855,In_26);
or U3835 (N_3835,In_1185,In_150);
or U3836 (N_3836,In_952,In_1736);
and U3837 (N_3837,In_361,In_1398);
or U3838 (N_3838,In_1537,In_759);
and U3839 (N_3839,In_1137,In_7);
nor U3840 (N_3840,In_1985,In_465);
and U3841 (N_3841,In_860,In_1454);
nand U3842 (N_3842,In_1498,In_713);
and U3843 (N_3843,In_122,In_956);
nor U3844 (N_3844,In_248,In_227);
nor U3845 (N_3845,In_1134,In_1543);
nor U3846 (N_3846,In_1577,In_481);
nor U3847 (N_3847,In_1306,In_1725);
nand U3848 (N_3848,In_160,In_1944);
and U3849 (N_3849,In_1452,In_940);
nor U3850 (N_3850,In_1120,In_1367);
or U3851 (N_3851,In_1705,In_1060);
nand U3852 (N_3852,In_855,In_934);
nand U3853 (N_3853,In_1330,In_1055);
and U3854 (N_3854,In_1156,In_482);
nand U3855 (N_3855,In_835,In_1068);
and U3856 (N_3856,In_1604,In_1567);
or U3857 (N_3857,In_697,In_852);
nor U3858 (N_3858,In_1635,In_1499);
nor U3859 (N_3859,In_1212,In_1114);
or U3860 (N_3860,In_201,In_866);
nand U3861 (N_3861,In_80,In_1613);
or U3862 (N_3862,In_546,In_58);
nor U3863 (N_3863,In_1870,In_617);
nor U3864 (N_3864,In_1055,In_385);
nand U3865 (N_3865,In_388,In_643);
or U3866 (N_3866,In_407,In_1063);
and U3867 (N_3867,In_277,In_1404);
nor U3868 (N_3868,In_1252,In_820);
nand U3869 (N_3869,In_1341,In_1988);
nor U3870 (N_3870,In_664,In_539);
or U3871 (N_3871,In_1390,In_565);
or U3872 (N_3872,In_1715,In_1065);
and U3873 (N_3873,In_555,In_739);
or U3874 (N_3874,In_1828,In_490);
or U3875 (N_3875,In_752,In_1682);
nand U3876 (N_3876,In_1949,In_350);
or U3877 (N_3877,In_19,In_1572);
and U3878 (N_3878,In_545,In_452);
nand U3879 (N_3879,In_569,In_55);
or U3880 (N_3880,In_1157,In_1725);
and U3881 (N_3881,In_1854,In_1817);
nor U3882 (N_3882,In_193,In_1967);
and U3883 (N_3883,In_630,In_1134);
nand U3884 (N_3884,In_892,In_1727);
nand U3885 (N_3885,In_1576,In_4);
nand U3886 (N_3886,In_580,In_839);
and U3887 (N_3887,In_218,In_1301);
nand U3888 (N_3888,In_1208,In_1992);
nor U3889 (N_3889,In_354,In_1204);
nor U3890 (N_3890,In_868,In_293);
or U3891 (N_3891,In_449,In_1859);
and U3892 (N_3892,In_1556,In_774);
nor U3893 (N_3893,In_657,In_143);
nand U3894 (N_3894,In_400,In_1026);
or U3895 (N_3895,In_137,In_1054);
nor U3896 (N_3896,In_10,In_1847);
or U3897 (N_3897,In_762,In_1012);
nand U3898 (N_3898,In_744,In_99);
nor U3899 (N_3899,In_1905,In_1265);
nor U3900 (N_3900,In_918,In_1668);
or U3901 (N_3901,In_1014,In_849);
nor U3902 (N_3902,In_1863,In_1645);
nand U3903 (N_3903,In_49,In_1476);
or U3904 (N_3904,In_43,In_1546);
or U3905 (N_3905,In_152,In_1939);
nand U3906 (N_3906,In_1347,In_629);
and U3907 (N_3907,In_158,In_780);
or U3908 (N_3908,In_1200,In_1666);
nor U3909 (N_3909,In_791,In_1424);
nor U3910 (N_3910,In_1932,In_852);
or U3911 (N_3911,In_489,In_57);
nor U3912 (N_3912,In_1693,In_1046);
nand U3913 (N_3913,In_773,In_1198);
or U3914 (N_3914,In_653,In_1279);
or U3915 (N_3915,In_1295,In_1101);
nand U3916 (N_3916,In_1220,In_1440);
nand U3917 (N_3917,In_1958,In_554);
nor U3918 (N_3918,In_850,In_1556);
and U3919 (N_3919,In_878,In_1291);
and U3920 (N_3920,In_1242,In_88);
and U3921 (N_3921,In_893,In_1622);
or U3922 (N_3922,In_408,In_23);
or U3923 (N_3923,In_1775,In_969);
nor U3924 (N_3924,In_1252,In_97);
or U3925 (N_3925,In_1643,In_39);
and U3926 (N_3926,In_625,In_108);
nand U3927 (N_3927,In_1720,In_1295);
nor U3928 (N_3928,In_1462,In_193);
nor U3929 (N_3929,In_968,In_1635);
nand U3930 (N_3930,In_323,In_1740);
nor U3931 (N_3931,In_793,In_1534);
nand U3932 (N_3932,In_830,In_1418);
nor U3933 (N_3933,In_1668,In_1416);
or U3934 (N_3934,In_62,In_825);
nand U3935 (N_3935,In_710,In_1455);
and U3936 (N_3936,In_1731,In_1560);
nor U3937 (N_3937,In_1843,In_1012);
or U3938 (N_3938,In_1088,In_485);
and U3939 (N_3939,In_1819,In_494);
and U3940 (N_3940,In_1284,In_1105);
and U3941 (N_3941,In_1100,In_917);
nor U3942 (N_3942,In_993,In_1584);
nor U3943 (N_3943,In_110,In_1143);
nand U3944 (N_3944,In_1003,In_68);
nand U3945 (N_3945,In_1540,In_1958);
or U3946 (N_3946,In_1885,In_1683);
or U3947 (N_3947,In_1266,In_1097);
or U3948 (N_3948,In_1317,In_1686);
nor U3949 (N_3949,In_1344,In_1744);
and U3950 (N_3950,In_1324,In_1199);
nor U3951 (N_3951,In_1912,In_1535);
nor U3952 (N_3952,In_50,In_1493);
or U3953 (N_3953,In_1091,In_542);
and U3954 (N_3954,In_599,In_678);
and U3955 (N_3955,In_1121,In_1778);
and U3956 (N_3956,In_248,In_1711);
nand U3957 (N_3957,In_1084,In_1057);
nor U3958 (N_3958,In_3,In_1269);
and U3959 (N_3959,In_1230,In_162);
nand U3960 (N_3960,In_378,In_385);
and U3961 (N_3961,In_287,In_835);
nand U3962 (N_3962,In_1326,In_1096);
and U3963 (N_3963,In_1641,In_653);
or U3964 (N_3964,In_543,In_1930);
nor U3965 (N_3965,In_953,In_1929);
nand U3966 (N_3966,In_394,In_1254);
and U3967 (N_3967,In_502,In_539);
nand U3968 (N_3968,In_603,In_1872);
or U3969 (N_3969,In_7,In_380);
and U3970 (N_3970,In_62,In_747);
nand U3971 (N_3971,In_1513,In_2);
nand U3972 (N_3972,In_205,In_1370);
nand U3973 (N_3973,In_798,In_1358);
and U3974 (N_3974,In_867,In_532);
and U3975 (N_3975,In_959,In_1091);
nor U3976 (N_3976,In_1889,In_1208);
nor U3977 (N_3977,In_1032,In_32);
and U3978 (N_3978,In_955,In_1731);
and U3979 (N_3979,In_1904,In_1929);
or U3980 (N_3980,In_706,In_1881);
or U3981 (N_3981,In_1011,In_1091);
nand U3982 (N_3982,In_107,In_902);
nor U3983 (N_3983,In_1956,In_247);
nand U3984 (N_3984,In_766,In_658);
nand U3985 (N_3985,In_1796,In_1036);
nand U3986 (N_3986,In_790,In_1452);
nor U3987 (N_3987,In_999,In_130);
or U3988 (N_3988,In_1240,In_885);
nor U3989 (N_3989,In_107,In_1141);
or U3990 (N_3990,In_1561,In_58);
nor U3991 (N_3991,In_204,In_488);
or U3992 (N_3992,In_1500,In_936);
nor U3993 (N_3993,In_453,In_1253);
nand U3994 (N_3994,In_1499,In_1668);
nor U3995 (N_3995,In_1070,In_539);
and U3996 (N_3996,In_1374,In_649);
nand U3997 (N_3997,In_53,In_1371);
and U3998 (N_3998,In_1176,In_207);
and U3999 (N_3999,In_1960,In_1938);
nand U4000 (N_4000,In_1427,In_30);
or U4001 (N_4001,In_1159,In_1585);
and U4002 (N_4002,In_566,In_1599);
and U4003 (N_4003,In_1974,In_771);
nand U4004 (N_4004,In_1165,In_918);
or U4005 (N_4005,In_621,In_669);
or U4006 (N_4006,In_1724,In_1978);
nor U4007 (N_4007,In_1539,In_1716);
nand U4008 (N_4008,In_1424,In_1637);
and U4009 (N_4009,In_1293,In_1592);
or U4010 (N_4010,In_109,In_552);
or U4011 (N_4011,In_937,In_1454);
or U4012 (N_4012,In_538,In_829);
nor U4013 (N_4013,In_1452,In_529);
or U4014 (N_4014,In_1663,In_1049);
or U4015 (N_4015,In_1326,In_1520);
or U4016 (N_4016,In_500,In_1888);
nand U4017 (N_4017,In_1253,In_1204);
nand U4018 (N_4018,In_333,In_169);
and U4019 (N_4019,In_293,In_279);
and U4020 (N_4020,In_593,In_211);
nor U4021 (N_4021,In_445,In_1585);
and U4022 (N_4022,In_1872,In_1027);
or U4023 (N_4023,In_1967,In_1833);
nand U4024 (N_4024,In_1264,In_402);
nand U4025 (N_4025,In_950,In_1280);
nor U4026 (N_4026,In_630,In_1230);
nand U4027 (N_4027,In_653,In_1932);
nor U4028 (N_4028,In_1901,In_396);
and U4029 (N_4029,In_1161,In_1160);
nor U4030 (N_4030,In_1417,In_920);
nor U4031 (N_4031,In_1750,In_692);
nand U4032 (N_4032,In_51,In_1381);
nor U4033 (N_4033,In_39,In_1112);
nor U4034 (N_4034,In_295,In_458);
nor U4035 (N_4035,In_1649,In_1267);
nand U4036 (N_4036,In_42,In_1477);
or U4037 (N_4037,In_1385,In_463);
and U4038 (N_4038,In_682,In_353);
or U4039 (N_4039,In_1001,In_162);
and U4040 (N_4040,In_110,In_1882);
nand U4041 (N_4041,In_444,In_577);
or U4042 (N_4042,In_950,In_1737);
and U4043 (N_4043,In_1835,In_1218);
nor U4044 (N_4044,In_1928,In_1204);
nand U4045 (N_4045,In_1788,In_215);
nand U4046 (N_4046,In_1647,In_240);
and U4047 (N_4047,In_810,In_186);
or U4048 (N_4048,In_983,In_760);
nor U4049 (N_4049,In_1912,In_1980);
nand U4050 (N_4050,In_1674,In_118);
and U4051 (N_4051,In_1225,In_648);
nand U4052 (N_4052,In_740,In_515);
nand U4053 (N_4053,In_1907,In_1081);
or U4054 (N_4054,In_1908,In_622);
and U4055 (N_4055,In_1998,In_123);
nor U4056 (N_4056,In_1943,In_874);
nor U4057 (N_4057,In_1801,In_826);
or U4058 (N_4058,In_894,In_1020);
nor U4059 (N_4059,In_728,In_1528);
or U4060 (N_4060,In_1654,In_595);
or U4061 (N_4061,In_1127,In_1383);
or U4062 (N_4062,In_1732,In_1294);
or U4063 (N_4063,In_1189,In_835);
nand U4064 (N_4064,In_560,In_214);
nand U4065 (N_4065,In_1981,In_578);
nand U4066 (N_4066,In_1545,In_1782);
and U4067 (N_4067,In_1334,In_262);
nand U4068 (N_4068,In_324,In_80);
and U4069 (N_4069,In_1027,In_942);
nand U4070 (N_4070,In_1180,In_162);
xor U4071 (N_4071,In_624,In_318);
and U4072 (N_4072,In_124,In_1134);
nand U4073 (N_4073,In_179,In_1993);
and U4074 (N_4074,In_1462,In_661);
and U4075 (N_4075,In_799,In_498);
nand U4076 (N_4076,In_179,In_1596);
and U4077 (N_4077,In_1075,In_708);
and U4078 (N_4078,In_433,In_1726);
and U4079 (N_4079,In_194,In_1212);
nor U4080 (N_4080,In_965,In_1941);
or U4081 (N_4081,In_259,In_1029);
nand U4082 (N_4082,In_1222,In_643);
or U4083 (N_4083,In_723,In_366);
nor U4084 (N_4084,In_634,In_1610);
nor U4085 (N_4085,In_905,In_1831);
or U4086 (N_4086,In_716,In_1254);
and U4087 (N_4087,In_1938,In_577);
nand U4088 (N_4088,In_601,In_1250);
nand U4089 (N_4089,In_692,In_1786);
and U4090 (N_4090,In_1762,In_41);
and U4091 (N_4091,In_1108,In_1695);
nand U4092 (N_4092,In_1902,In_759);
and U4093 (N_4093,In_1141,In_195);
and U4094 (N_4094,In_1408,In_217);
nand U4095 (N_4095,In_1762,In_69);
or U4096 (N_4096,In_1157,In_193);
or U4097 (N_4097,In_640,In_915);
or U4098 (N_4098,In_956,In_500);
or U4099 (N_4099,In_491,In_874);
nand U4100 (N_4100,In_1875,In_485);
and U4101 (N_4101,In_17,In_29);
nand U4102 (N_4102,In_1974,In_477);
and U4103 (N_4103,In_446,In_1625);
and U4104 (N_4104,In_999,In_809);
nand U4105 (N_4105,In_1035,In_407);
and U4106 (N_4106,In_1461,In_1863);
or U4107 (N_4107,In_353,In_1167);
or U4108 (N_4108,In_1459,In_1112);
xnor U4109 (N_4109,In_1048,In_1794);
or U4110 (N_4110,In_1407,In_1697);
and U4111 (N_4111,In_169,In_1767);
nor U4112 (N_4112,In_1954,In_1358);
nand U4113 (N_4113,In_1875,In_244);
nand U4114 (N_4114,In_610,In_76);
or U4115 (N_4115,In_1499,In_1079);
and U4116 (N_4116,In_1023,In_1606);
and U4117 (N_4117,In_1315,In_856);
and U4118 (N_4118,In_727,In_1463);
or U4119 (N_4119,In_1244,In_1762);
and U4120 (N_4120,In_1740,In_1767);
xor U4121 (N_4121,In_1423,In_1373);
nor U4122 (N_4122,In_778,In_229);
nand U4123 (N_4123,In_813,In_1980);
nor U4124 (N_4124,In_1001,In_1841);
nor U4125 (N_4125,In_1039,In_1329);
nor U4126 (N_4126,In_1739,In_586);
or U4127 (N_4127,In_1562,In_982);
and U4128 (N_4128,In_243,In_1741);
nor U4129 (N_4129,In_836,In_1892);
and U4130 (N_4130,In_107,In_504);
and U4131 (N_4131,In_1684,In_1445);
nor U4132 (N_4132,In_219,In_1792);
or U4133 (N_4133,In_1230,In_452);
and U4134 (N_4134,In_1925,In_1013);
or U4135 (N_4135,In_1951,In_541);
nand U4136 (N_4136,In_1603,In_147);
nor U4137 (N_4137,In_352,In_1281);
nand U4138 (N_4138,In_989,In_1715);
nor U4139 (N_4139,In_1410,In_1792);
nand U4140 (N_4140,In_201,In_1000);
and U4141 (N_4141,In_560,In_1903);
nand U4142 (N_4142,In_706,In_514);
nor U4143 (N_4143,In_977,In_1760);
nor U4144 (N_4144,In_1652,In_10);
nand U4145 (N_4145,In_1651,In_1060);
or U4146 (N_4146,In_143,In_1520);
nand U4147 (N_4147,In_574,In_729);
or U4148 (N_4148,In_1012,In_1824);
nand U4149 (N_4149,In_659,In_755);
or U4150 (N_4150,In_349,In_286);
nand U4151 (N_4151,In_478,In_1978);
nand U4152 (N_4152,In_227,In_972);
or U4153 (N_4153,In_1901,In_689);
or U4154 (N_4154,In_840,In_605);
xor U4155 (N_4155,In_1252,In_1311);
nor U4156 (N_4156,In_783,In_907);
and U4157 (N_4157,In_1687,In_1346);
or U4158 (N_4158,In_1304,In_1595);
nor U4159 (N_4159,In_197,In_337);
nand U4160 (N_4160,In_204,In_1149);
nand U4161 (N_4161,In_1144,In_1219);
or U4162 (N_4162,In_314,In_1043);
nand U4163 (N_4163,In_1267,In_878);
or U4164 (N_4164,In_1858,In_725);
and U4165 (N_4165,In_1844,In_1143);
and U4166 (N_4166,In_1696,In_686);
and U4167 (N_4167,In_1837,In_1946);
nor U4168 (N_4168,In_1295,In_326);
or U4169 (N_4169,In_816,In_1873);
and U4170 (N_4170,In_1732,In_943);
and U4171 (N_4171,In_7,In_483);
and U4172 (N_4172,In_1920,In_736);
nand U4173 (N_4173,In_792,In_1323);
nand U4174 (N_4174,In_437,In_210);
and U4175 (N_4175,In_293,In_522);
nor U4176 (N_4176,In_1971,In_1739);
nor U4177 (N_4177,In_390,In_17);
and U4178 (N_4178,In_485,In_1187);
and U4179 (N_4179,In_637,In_1164);
nand U4180 (N_4180,In_1278,In_1780);
nor U4181 (N_4181,In_829,In_1092);
and U4182 (N_4182,In_1737,In_1670);
and U4183 (N_4183,In_462,In_1527);
and U4184 (N_4184,In_1899,In_1007);
nand U4185 (N_4185,In_668,In_1198);
nand U4186 (N_4186,In_681,In_1611);
or U4187 (N_4187,In_409,In_878);
and U4188 (N_4188,In_816,In_243);
nor U4189 (N_4189,In_541,In_1242);
nor U4190 (N_4190,In_1984,In_1154);
nand U4191 (N_4191,In_1897,In_563);
or U4192 (N_4192,In_671,In_1278);
or U4193 (N_4193,In_629,In_1936);
nand U4194 (N_4194,In_1357,In_265);
and U4195 (N_4195,In_398,In_1642);
nand U4196 (N_4196,In_1739,In_387);
or U4197 (N_4197,In_1576,In_514);
or U4198 (N_4198,In_1435,In_1039);
xnor U4199 (N_4199,In_1505,In_1496);
and U4200 (N_4200,In_114,In_329);
nor U4201 (N_4201,In_357,In_220);
nand U4202 (N_4202,In_1687,In_1683);
and U4203 (N_4203,In_1906,In_347);
nand U4204 (N_4204,In_291,In_987);
nand U4205 (N_4205,In_1288,In_1678);
nand U4206 (N_4206,In_1739,In_881);
nor U4207 (N_4207,In_1652,In_1446);
nor U4208 (N_4208,In_1164,In_377);
nor U4209 (N_4209,In_1347,In_1337);
nand U4210 (N_4210,In_98,In_1713);
nor U4211 (N_4211,In_1229,In_1039);
and U4212 (N_4212,In_1617,In_1683);
or U4213 (N_4213,In_621,In_476);
nand U4214 (N_4214,In_1287,In_909);
or U4215 (N_4215,In_350,In_1927);
or U4216 (N_4216,In_1105,In_905);
nor U4217 (N_4217,In_1600,In_1837);
and U4218 (N_4218,In_218,In_1252);
nor U4219 (N_4219,In_1329,In_944);
and U4220 (N_4220,In_1314,In_1441);
or U4221 (N_4221,In_1322,In_110);
and U4222 (N_4222,In_1380,In_72);
nor U4223 (N_4223,In_1572,In_160);
and U4224 (N_4224,In_1235,In_924);
and U4225 (N_4225,In_1291,In_1912);
nand U4226 (N_4226,In_618,In_949);
nor U4227 (N_4227,In_1193,In_514);
nand U4228 (N_4228,In_1328,In_330);
and U4229 (N_4229,In_1033,In_877);
nor U4230 (N_4230,In_175,In_678);
nor U4231 (N_4231,In_427,In_1682);
and U4232 (N_4232,In_1293,In_949);
nand U4233 (N_4233,In_1178,In_404);
nand U4234 (N_4234,In_9,In_239);
and U4235 (N_4235,In_176,In_893);
nor U4236 (N_4236,In_1995,In_726);
and U4237 (N_4237,In_602,In_1659);
or U4238 (N_4238,In_574,In_1486);
or U4239 (N_4239,In_1977,In_1534);
nor U4240 (N_4240,In_1144,In_1296);
and U4241 (N_4241,In_1526,In_471);
and U4242 (N_4242,In_1614,In_122);
nor U4243 (N_4243,In_867,In_715);
nand U4244 (N_4244,In_1402,In_269);
or U4245 (N_4245,In_32,In_37);
or U4246 (N_4246,In_1789,In_1632);
and U4247 (N_4247,In_1707,In_135);
and U4248 (N_4248,In_1832,In_1421);
nand U4249 (N_4249,In_200,In_1573);
nor U4250 (N_4250,In_966,In_804);
nor U4251 (N_4251,In_364,In_319);
nand U4252 (N_4252,In_621,In_1169);
and U4253 (N_4253,In_1415,In_293);
nor U4254 (N_4254,In_1382,In_601);
or U4255 (N_4255,In_901,In_1304);
nor U4256 (N_4256,In_883,In_1664);
and U4257 (N_4257,In_1054,In_1454);
nor U4258 (N_4258,In_1924,In_678);
nand U4259 (N_4259,In_1323,In_1748);
nand U4260 (N_4260,In_1792,In_1281);
nor U4261 (N_4261,In_119,In_1524);
or U4262 (N_4262,In_1070,In_1292);
nand U4263 (N_4263,In_1130,In_1744);
or U4264 (N_4264,In_1371,In_1423);
or U4265 (N_4265,In_602,In_860);
nand U4266 (N_4266,In_333,In_418);
and U4267 (N_4267,In_1302,In_1520);
nand U4268 (N_4268,In_1007,In_1943);
nor U4269 (N_4269,In_573,In_1667);
and U4270 (N_4270,In_1168,In_625);
nor U4271 (N_4271,In_1884,In_521);
or U4272 (N_4272,In_742,In_963);
or U4273 (N_4273,In_1693,In_1195);
nor U4274 (N_4274,In_655,In_608);
nor U4275 (N_4275,In_272,In_357);
and U4276 (N_4276,In_50,In_527);
and U4277 (N_4277,In_1544,In_155);
or U4278 (N_4278,In_1757,In_1015);
and U4279 (N_4279,In_364,In_136);
and U4280 (N_4280,In_1877,In_887);
or U4281 (N_4281,In_1828,In_1626);
and U4282 (N_4282,In_533,In_498);
nand U4283 (N_4283,In_1705,In_429);
and U4284 (N_4284,In_1271,In_1065);
nor U4285 (N_4285,In_1515,In_1116);
or U4286 (N_4286,In_1288,In_1108);
nor U4287 (N_4287,In_1699,In_998);
and U4288 (N_4288,In_31,In_845);
and U4289 (N_4289,In_476,In_1969);
nand U4290 (N_4290,In_1395,In_1338);
nor U4291 (N_4291,In_535,In_1270);
nor U4292 (N_4292,In_1472,In_558);
and U4293 (N_4293,In_446,In_1447);
nand U4294 (N_4294,In_36,In_1321);
or U4295 (N_4295,In_1601,In_816);
nor U4296 (N_4296,In_907,In_957);
nor U4297 (N_4297,In_708,In_72);
nand U4298 (N_4298,In_1648,In_925);
nand U4299 (N_4299,In_1285,In_219);
and U4300 (N_4300,In_1032,In_114);
nand U4301 (N_4301,In_1621,In_502);
nor U4302 (N_4302,In_1007,In_1128);
nor U4303 (N_4303,In_311,In_1797);
nand U4304 (N_4304,In_1523,In_1765);
or U4305 (N_4305,In_1343,In_874);
nor U4306 (N_4306,In_267,In_640);
and U4307 (N_4307,In_977,In_1194);
nor U4308 (N_4308,In_1976,In_279);
or U4309 (N_4309,In_1112,In_911);
nand U4310 (N_4310,In_324,In_1854);
nand U4311 (N_4311,In_797,In_1197);
or U4312 (N_4312,In_810,In_585);
and U4313 (N_4313,In_1525,In_558);
or U4314 (N_4314,In_862,In_1239);
nor U4315 (N_4315,In_1526,In_1435);
nand U4316 (N_4316,In_879,In_1936);
nand U4317 (N_4317,In_536,In_1422);
or U4318 (N_4318,In_1238,In_1791);
nor U4319 (N_4319,In_1586,In_852);
nor U4320 (N_4320,In_410,In_1578);
and U4321 (N_4321,In_1861,In_1162);
or U4322 (N_4322,In_208,In_761);
and U4323 (N_4323,In_1046,In_835);
nand U4324 (N_4324,In_172,In_853);
and U4325 (N_4325,In_150,In_1285);
and U4326 (N_4326,In_679,In_177);
nor U4327 (N_4327,In_1550,In_1251);
nor U4328 (N_4328,In_993,In_95);
nand U4329 (N_4329,In_1366,In_1305);
or U4330 (N_4330,In_1982,In_1943);
nand U4331 (N_4331,In_1200,In_1778);
nor U4332 (N_4332,In_1662,In_174);
or U4333 (N_4333,In_1977,In_1878);
nor U4334 (N_4334,In_1054,In_1926);
nand U4335 (N_4335,In_1869,In_1774);
or U4336 (N_4336,In_566,In_1656);
nor U4337 (N_4337,In_1270,In_687);
or U4338 (N_4338,In_1943,In_1784);
nand U4339 (N_4339,In_914,In_505);
nand U4340 (N_4340,In_1985,In_1076);
nand U4341 (N_4341,In_1103,In_1552);
nor U4342 (N_4342,In_730,In_603);
nor U4343 (N_4343,In_1881,In_1143);
nand U4344 (N_4344,In_1918,In_1218);
nor U4345 (N_4345,In_1588,In_2);
nand U4346 (N_4346,In_1577,In_1461);
and U4347 (N_4347,In_1671,In_659);
or U4348 (N_4348,In_415,In_880);
nor U4349 (N_4349,In_498,In_859);
or U4350 (N_4350,In_869,In_795);
xor U4351 (N_4351,In_684,In_1093);
or U4352 (N_4352,In_782,In_970);
or U4353 (N_4353,In_1224,In_1472);
nor U4354 (N_4354,In_482,In_1779);
and U4355 (N_4355,In_198,In_547);
and U4356 (N_4356,In_350,In_1251);
nor U4357 (N_4357,In_890,In_761);
nand U4358 (N_4358,In_1130,In_1981);
or U4359 (N_4359,In_1577,In_1738);
or U4360 (N_4360,In_1665,In_1432);
or U4361 (N_4361,In_917,In_1702);
nor U4362 (N_4362,In_1550,In_1861);
nor U4363 (N_4363,In_272,In_1712);
or U4364 (N_4364,In_296,In_133);
and U4365 (N_4365,In_1842,In_1081);
and U4366 (N_4366,In_449,In_1599);
nor U4367 (N_4367,In_1805,In_1342);
or U4368 (N_4368,In_1256,In_393);
nand U4369 (N_4369,In_1253,In_359);
nor U4370 (N_4370,In_14,In_1847);
or U4371 (N_4371,In_894,In_76);
nor U4372 (N_4372,In_1208,In_1193);
and U4373 (N_4373,In_1757,In_1461);
or U4374 (N_4374,In_159,In_1298);
or U4375 (N_4375,In_25,In_493);
nor U4376 (N_4376,In_839,In_486);
nand U4377 (N_4377,In_1832,In_588);
or U4378 (N_4378,In_722,In_1220);
or U4379 (N_4379,In_287,In_466);
or U4380 (N_4380,In_719,In_1316);
and U4381 (N_4381,In_1434,In_116);
and U4382 (N_4382,In_1281,In_1805);
and U4383 (N_4383,In_593,In_1283);
nand U4384 (N_4384,In_1510,In_1274);
nand U4385 (N_4385,In_1916,In_1341);
nand U4386 (N_4386,In_615,In_1041);
nor U4387 (N_4387,In_44,In_1495);
and U4388 (N_4388,In_972,In_302);
or U4389 (N_4389,In_1508,In_1264);
or U4390 (N_4390,In_411,In_1606);
or U4391 (N_4391,In_1865,In_1380);
nand U4392 (N_4392,In_1933,In_1428);
nor U4393 (N_4393,In_561,In_1019);
nor U4394 (N_4394,In_1894,In_1112);
and U4395 (N_4395,In_1430,In_571);
or U4396 (N_4396,In_852,In_1842);
nor U4397 (N_4397,In_1039,In_1256);
or U4398 (N_4398,In_1002,In_35);
or U4399 (N_4399,In_826,In_1604);
nor U4400 (N_4400,In_994,In_978);
or U4401 (N_4401,In_974,In_1965);
and U4402 (N_4402,In_446,In_719);
and U4403 (N_4403,In_662,In_710);
nand U4404 (N_4404,In_332,In_203);
or U4405 (N_4405,In_437,In_952);
or U4406 (N_4406,In_4,In_14);
or U4407 (N_4407,In_231,In_541);
or U4408 (N_4408,In_1033,In_579);
or U4409 (N_4409,In_1822,In_1285);
nand U4410 (N_4410,In_1038,In_1063);
and U4411 (N_4411,In_531,In_397);
nor U4412 (N_4412,In_1448,In_1420);
and U4413 (N_4413,In_1547,In_1571);
or U4414 (N_4414,In_1564,In_820);
and U4415 (N_4415,In_1609,In_1705);
nor U4416 (N_4416,In_657,In_159);
nand U4417 (N_4417,In_532,In_184);
nand U4418 (N_4418,In_231,In_1279);
nor U4419 (N_4419,In_290,In_1761);
nand U4420 (N_4420,In_729,In_1325);
nor U4421 (N_4421,In_1438,In_1693);
and U4422 (N_4422,In_1448,In_823);
nor U4423 (N_4423,In_43,In_1278);
or U4424 (N_4424,In_336,In_804);
nor U4425 (N_4425,In_1741,In_162);
xor U4426 (N_4426,In_270,In_1404);
nand U4427 (N_4427,In_816,In_957);
nor U4428 (N_4428,In_1138,In_1131);
nor U4429 (N_4429,In_774,In_658);
nor U4430 (N_4430,In_978,In_722);
and U4431 (N_4431,In_735,In_497);
and U4432 (N_4432,In_1211,In_1472);
or U4433 (N_4433,In_590,In_815);
or U4434 (N_4434,In_1698,In_135);
nor U4435 (N_4435,In_1624,In_196);
nor U4436 (N_4436,In_234,In_632);
nor U4437 (N_4437,In_1140,In_338);
nor U4438 (N_4438,In_126,In_641);
nand U4439 (N_4439,In_267,In_46);
or U4440 (N_4440,In_1160,In_1933);
nand U4441 (N_4441,In_278,In_752);
nor U4442 (N_4442,In_1749,In_980);
and U4443 (N_4443,In_1211,In_802);
or U4444 (N_4444,In_1186,In_1864);
nor U4445 (N_4445,In_118,In_495);
nand U4446 (N_4446,In_1058,In_772);
nand U4447 (N_4447,In_1116,In_1270);
nand U4448 (N_4448,In_52,In_1480);
nor U4449 (N_4449,In_1690,In_1170);
nor U4450 (N_4450,In_1712,In_121);
nand U4451 (N_4451,In_195,In_415);
and U4452 (N_4452,In_1610,In_1367);
or U4453 (N_4453,In_1267,In_564);
or U4454 (N_4454,In_694,In_1926);
nor U4455 (N_4455,In_556,In_1427);
nand U4456 (N_4456,In_723,In_424);
nand U4457 (N_4457,In_1899,In_678);
and U4458 (N_4458,In_1490,In_1489);
and U4459 (N_4459,In_1639,In_1334);
nor U4460 (N_4460,In_388,In_291);
xor U4461 (N_4461,In_607,In_122);
nand U4462 (N_4462,In_1460,In_1151);
nand U4463 (N_4463,In_695,In_525);
nand U4464 (N_4464,In_843,In_1833);
or U4465 (N_4465,In_1102,In_853);
and U4466 (N_4466,In_450,In_1247);
nor U4467 (N_4467,In_77,In_155);
nand U4468 (N_4468,In_745,In_436);
or U4469 (N_4469,In_1881,In_1062);
nor U4470 (N_4470,In_1781,In_1353);
and U4471 (N_4471,In_308,In_965);
nand U4472 (N_4472,In_177,In_267);
nand U4473 (N_4473,In_1158,In_1599);
nor U4474 (N_4474,In_1578,In_1530);
or U4475 (N_4475,In_1214,In_654);
or U4476 (N_4476,In_927,In_1037);
nor U4477 (N_4477,In_7,In_1479);
and U4478 (N_4478,In_655,In_541);
nor U4479 (N_4479,In_1647,In_334);
nor U4480 (N_4480,In_1071,In_901);
nor U4481 (N_4481,In_758,In_1689);
and U4482 (N_4482,In_1875,In_1990);
or U4483 (N_4483,In_1029,In_614);
and U4484 (N_4484,In_1111,In_818);
nor U4485 (N_4485,In_78,In_188);
nor U4486 (N_4486,In_1258,In_1447);
or U4487 (N_4487,In_47,In_1678);
or U4488 (N_4488,In_736,In_1128);
and U4489 (N_4489,In_1118,In_1892);
xor U4490 (N_4490,In_547,In_1570);
nor U4491 (N_4491,In_697,In_562);
or U4492 (N_4492,In_1871,In_740);
or U4493 (N_4493,In_911,In_1371);
nand U4494 (N_4494,In_71,In_352);
nand U4495 (N_4495,In_1180,In_1229);
or U4496 (N_4496,In_1804,In_321);
and U4497 (N_4497,In_15,In_910);
nand U4498 (N_4498,In_1742,In_1074);
and U4499 (N_4499,In_1780,In_72);
nand U4500 (N_4500,In_1409,In_206);
nand U4501 (N_4501,In_885,In_380);
nand U4502 (N_4502,In_1907,In_1649);
or U4503 (N_4503,In_1489,In_434);
nor U4504 (N_4504,In_1333,In_1243);
and U4505 (N_4505,In_1735,In_803);
and U4506 (N_4506,In_275,In_1972);
and U4507 (N_4507,In_545,In_838);
nor U4508 (N_4508,In_1540,In_1927);
nand U4509 (N_4509,In_184,In_219);
and U4510 (N_4510,In_110,In_392);
or U4511 (N_4511,In_1347,In_1060);
nand U4512 (N_4512,In_691,In_412);
or U4513 (N_4513,In_705,In_1704);
nor U4514 (N_4514,In_1812,In_1385);
or U4515 (N_4515,In_1994,In_73);
and U4516 (N_4516,In_1420,In_155);
nand U4517 (N_4517,In_1636,In_381);
or U4518 (N_4518,In_1645,In_483);
nand U4519 (N_4519,In_1789,In_1661);
nand U4520 (N_4520,In_466,In_1872);
and U4521 (N_4521,In_1670,In_931);
nor U4522 (N_4522,In_1533,In_1143);
nand U4523 (N_4523,In_1458,In_253);
nand U4524 (N_4524,In_825,In_1028);
nand U4525 (N_4525,In_1930,In_811);
nor U4526 (N_4526,In_1927,In_1591);
and U4527 (N_4527,In_1114,In_579);
and U4528 (N_4528,In_1627,In_32);
and U4529 (N_4529,In_118,In_584);
and U4530 (N_4530,In_1356,In_1690);
nand U4531 (N_4531,In_312,In_924);
and U4532 (N_4532,In_1841,In_1316);
xnor U4533 (N_4533,In_1756,In_1469);
or U4534 (N_4534,In_1900,In_458);
and U4535 (N_4535,In_1754,In_1201);
and U4536 (N_4536,In_1798,In_1291);
nand U4537 (N_4537,In_1873,In_1494);
nor U4538 (N_4538,In_1515,In_1750);
or U4539 (N_4539,In_811,In_385);
and U4540 (N_4540,In_935,In_1863);
nor U4541 (N_4541,In_625,In_190);
and U4542 (N_4542,In_533,In_1384);
nor U4543 (N_4543,In_1353,In_659);
or U4544 (N_4544,In_1480,In_171);
nor U4545 (N_4545,In_1476,In_470);
and U4546 (N_4546,In_1406,In_1356);
or U4547 (N_4547,In_1399,In_23);
and U4548 (N_4548,In_1576,In_1061);
and U4549 (N_4549,In_1732,In_1957);
nor U4550 (N_4550,In_140,In_884);
nor U4551 (N_4551,In_158,In_1044);
nor U4552 (N_4552,In_794,In_1957);
nor U4553 (N_4553,In_875,In_965);
nor U4554 (N_4554,In_1437,In_999);
or U4555 (N_4555,In_272,In_1459);
nand U4556 (N_4556,In_725,In_1841);
and U4557 (N_4557,In_542,In_1617);
nor U4558 (N_4558,In_1156,In_998);
nand U4559 (N_4559,In_1616,In_1629);
and U4560 (N_4560,In_1232,In_341);
or U4561 (N_4561,In_930,In_295);
nor U4562 (N_4562,In_1236,In_653);
nand U4563 (N_4563,In_1308,In_780);
nor U4564 (N_4564,In_962,In_825);
or U4565 (N_4565,In_476,In_788);
or U4566 (N_4566,In_1747,In_331);
and U4567 (N_4567,In_211,In_1757);
and U4568 (N_4568,In_241,In_448);
nand U4569 (N_4569,In_1385,In_1747);
nand U4570 (N_4570,In_376,In_944);
nand U4571 (N_4571,In_1646,In_248);
or U4572 (N_4572,In_197,In_1127);
and U4573 (N_4573,In_1423,In_795);
and U4574 (N_4574,In_1429,In_1838);
nand U4575 (N_4575,In_60,In_838);
nand U4576 (N_4576,In_342,In_442);
and U4577 (N_4577,In_494,In_1845);
or U4578 (N_4578,In_1271,In_1112);
nor U4579 (N_4579,In_1668,In_228);
nor U4580 (N_4580,In_485,In_1027);
or U4581 (N_4581,In_1955,In_244);
or U4582 (N_4582,In_243,In_1987);
nor U4583 (N_4583,In_1221,In_184);
or U4584 (N_4584,In_445,In_1438);
or U4585 (N_4585,In_259,In_216);
or U4586 (N_4586,In_330,In_1772);
and U4587 (N_4587,In_997,In_1812);
nand U4588 (N_4588,In_1559,In_1254);
or U4589 (N_4589,In_66,In_1688);
xnor U4590 (N_4590,In_430,In_1180);
nor U4591 (N_4591,In_1375,In_274);
nand U4592 (N_4592,In_507,In_68);
or U4593 (N_4593,In_794,In_137);
or U4594 (N_4594,In_1963,In_272);
and U4595 (N_4595,In_1325,In_296);
and U4596 (N_4596,In_892,In_1110);
nand U4597 (N_4597,In_1990,In_728);
and U4598 (N_4598,In_1644,In_1769);
or U4599 (N_4599,In_1406,In_1155);
nor U4600 (N_4600,In_1974,In_1752);
nor U4601 (N_4601,In_1734,In_1359);
or U4602 (N_4602,In_1748,In_1344);
nor U4603 (N_4603,In_483,In_1473);
nand U4604 (N_4604,In_526,In_1390);
nor U4605 (N_4605,In_1290,In_2);
and U4606 (N_4606,In_860,In_1900);
nor U4607 (N_4607,In_375,In_1675);
or U4608 (N_4608,In_665,In_378);
and U4609 (N_4609,In_568,In_383);
or U4610 (N_4610,In_1718,In_1443);
and U4611 (N_4611,In_1147,In_931);
and U4612 (N_4612,In_1199,In_1789);
nor U4613 (N_4613,In_1203,In_1201);
and U4614 (N_4614,In_660,In_1520);
nor U4615 (N_4615,In_1378,In_471);
and U4616 (N_4616,In_74,In_1657);
and U4617 (N_4617,In_682,In_1496);
nor U4618 (N_4618,In_542,In_1766);
and U4619 (N_4619,In_1961,In_1959);
nand U4620 (N_4620,In_1930,In_1508);
nand U4621 (N_4621,In_1772,In_1527);
and U4622 (N_4622,In_397,In_1170);
and U4623 (N_4623,In_1699,In_272);
nand U4624 (N_4624,In_882,In_1632);
and U4625 (N_4625,In_687,In_1998);
nand U4626 (N_4626,In_527,In_561);
nand U4627 (N_4627,In_260,In_1395);
nor U4628 (N_4628,In_1564,In_588);
or U4629 (N_4629,In_1645,In_770);
nand U4630 (N_4630,In_1052,In_1797);
and U4631 (N_4631,In_1978,In_672);
and U4632 (N_4632,In_643,In_1591);
nand U4633 (N_4633,In_1314,In_994);
nor U4634 (N_4634,In_1612,In_854);
nand U4635 (N_4635,In_1825,In_182);
nand U4636 (N_4636,In_1140,In_641);
nand U4637 (N_4637,In_1488,In_1992);
nand U4638 (N_4638,In_1309,In_44);
nor U4639 (N_4639,In_1981,In_971);
nand U4640 (N_4640,In_1463,In_696);
or U4641 (N_4641,In_1251,In_175);
nand U4642 (N_4642,In_1476,In_985);
or U4643 (N_4643,In_1842,In_1012);
or U4644 (N_4644,In_1141,In_550);
nand U4645 (N_4645,In_1891,In_851);
or U4646 (N_4646,In_642,In_54);
or U4647 (N_4647,In_1315,In_1645);
nor U4648 (N_4648,In_583,In_815);
nand U4649 (N_4649,In_849,In_338);
nor U4650 (N_4650,In_1662,In_1144);
and U4651 (N_4651,In_1649,In_1375);
nand U4652 (N_4652,In_193,In_1257);
nor U4653 (N_4653,In_1413,In_837);
and U4654 (N_4654,In_1834,In_1211);
and U4655 (N_4655,In_712,In_1307);
xnor U4656 (N_4656,In_1724,In_257);
and U4657 (N_4657,In_1907,In_249);
and U4658 (N_4658,In_1216,In_136);
nand U4659 (N_4659,In_74,In_1759);
nand U4660 (N_4660,In_1037,In_1469);
nand U4661 (N_4661,In_1435,In_176);
and U4662 (N_4662,In_307,In_1780);
or U4663 (N_4663,In_1398,In_51);
nor U4664 (N_4664,In_357,In_316);
or U4665 (N_4665,In_315,In_943);
or U4666 (N_4666,In_989,In_1560);
or U4667 (N_4667,In_1911,In_349);
nor U4668 (N_4668,In_361,In_1778);
nor U4669 (N_4669,In_1238,In_1665);
nand U4670 (N_4670,In_1458,In_1526);
nand U4671 (N_4671,In_1753,In_952);
and U4672 (N_4672,In_205,In_137);
nand U4673 (N_4673,In_424,In_1395);
and U4674 (N_4674,In_911,In_1631);
or U4675 (N_4675,In_1117,In_1686);
nand U4676 (N_4676,In_1695,In_380);
nor U4677 (N_4677,In_1303,In_817);
or U4678 (N_4678,In_641,In_7);
or U4679 (N_4679,In_1191,In_1106);
or U4680 (N_4680,In_1366,In_1603);
nor U4681 (N_4681,In_1635,In_1934);
nor U4682 (N_4682,In_745,In_901);
and U4683 (N_4683,In_1634,In_592);
nor U4684 (N_4684,In_1568,In_756);
nand U4685 (N_4685,In_1625,In_452);
and U4686 (N_4686,In_1128,In_1907);
nor U4687 (N_4687,In_1804,In_1947);
nor U4688 (N_4688,In_212,In_853);
nor U4689 (N_4689,In_1526,In_1204);
nor U4690 (N_4690,In_1723,In_1166);
nand U4691 (N_4691,In_1101,In_1561);
or U4692 (N_4692,In_574,In_700);
or U4693 (N_4693,In_1363,In_1010);
nor U4694 (N_4694,In_1147,In_1566);
nand U4695 (N_4695,In_1876,In_1029);
nor U4696 (N_4696,In_915,In_1223);
and U4697 (N_4697,In_686,In_1164);
nand U4698 (N_4698,In_1298,In_1270);
nor U4699 (N_4699,In_140,In_1790);
nand U4700 (N_4700,In_82,In_1058);
nand U4701 (N_4701,In_1876,In_1714);
nand U4702 (N_4702,In_1174,In_421);
nand U4703 (N_4703,In_1820,In_1257);
and U4704 (N_4704,In_1059,In_1013);
nand U4705 (N_4705,In_861,In_1444);
nor U4706 (N_4706,In_1593,In_773);
or U4707 (N_4707,In_1775,In_985);
and U4708 (N_4708,In_1344,In_89);
or U4709 (N_4709,In_1340,In_706);
and U4710 (N_4710,In_93,In_1960);
nor U4711 (N_4711,In_481,In_169);
and U4712 (N_4712,In_1757,In_633);
nand U4713 (N_4713,In_1888,In_314);
nand U4714 (N_4714,In_1926,In_486);
or U4715 (N_4715,In_787,In_1689);
and U4716 (N_4716,In_97,In_956);
nand U4717 (N_4717,In_1324,In_1445);
or U4718 (N_4718,In_409,In_907);
nand U4719 (N_4719,In_1740,In_1838);
nor U4720 (N_4720,In_683,In_257);
nor U4721 (N_4721,In_103,In_220);
xnor U4722 (N_4722,In_625,In_1508);
nor U4723 (N_4723,In_1552,In_1565);
xor U4724 (N_4724,In_1567,In_744);
and U4725 (N_4725,In_982,In_1596);
or U4726 (N_4726,In_1152,In_152);
nor U4727 (N_4727,In_19,In_1320);
or U4728 (N_4728,In_1628,In_1936);
nand U4729 (N_4729,In_1174,In_1067);
and U4730 (N_4730,In_833,In_548);
and U4731 (N_4731,In_1017,In_1151);
nand U4732 (N_4732,In_913,In_1322);
nand U4733 (N_4733,In_569,In_429);
and U4734 (N_4734,In_760,In_1016);
nor U4735 (N_4735,In_343,In_25);
nor U4736 (N_4736,In_1191,In_1963);
or U4737 (N_4737,In_108,In_10);
or U4738 (N_4738,In_942,In_1423);
nand U4739 (N_4739,In_703,In_1372);
or U4740 (N_4740,In_1968,In_1419);
nor U4741 (N_4741,In_1702,In_522);
or U4742 (N_4742,In_1698,In_633);
nor U4743 (N_4743,In_1275,In_493);
nor U4744 (N_4744,In_1783,In_299);
or U4745 (N_4745,In_1626,In_1318);
and U4746 (N_4746,In_820,In_1012);
and U4747 (N_4747,In_539,In_1830);
or U4748 (N_4748,In_788,In_872);
nand U4749 (N_4749,In_741,In_1984);
or U4750 (N_4750,In_1570,In_941);
nand U4751 (N_4751,In_451,In_1434);
or U4752 (N_4752,In_913,In_131);
nand U4753 (N_4753,In_1185,In_1381);
and U4754 (N_4754,In_1256,In_723);
and U4755 (N_4755,In_1499,In_808);
and U4756 (N_4756,In_1459,In_1990);
and U4757 (N_4757,In_673,In_1875);
or U4758 (N_4758,In_147,In_1978);
and U4759 (N_4759,In_1225,In_184);
and U4760 (N_4760,In_1637,In_1491);
and U4761 (N_4761,In_1916,In_1149);
nand U4762 (N_4762,In_914,In_1726);
and U4763 (N_4763,In_1437,In_480);
and U4764 (N_4764,In_9,In_368);
and U4765 (N_4765,In_697,In_346);
nor U4766 (N_4766,In_552,In_1231);
or U4767 (N_4767,In_595,In_1536);
nand U4768 (N_4768,In_688,In_1591);
and U4769 (N_4769,In_350,In_229);
nor U4770 (N_4770,In_1413,In_548);
or U4771 (N_4771,In_536,In_158);
nor U4772 (N_4772,In_1778,In_972);
or U4773 (N_4773,In_579,In_1354);
or U4774 (N_4774,In_558,In_218);
nand U4775 (N_4775,In_93,In_1426);
or U4776 (N_4776,In_1923,In_360);
or U4777 (N_4777,In_556,In_1367);
nand U4778 (N_4778,In_1856,In_576);
and U4779 (N_4779,In_589,In_378);
nor U4780 (N_4780,In_938,In_753);
nand U4781 (N_4781,In_244,In_258);
nor U4782 (N_4782,In_846,In_1581);
and U4783 (N_4783,In_904,In_1503);
nor U4784 (N_4784,In_1708,In_759);
and U4785 (N_4785,In_306,In_383);
nand U4786 (N_4786,In_467,In_466);
and U4787 (N_4787,In_643,In_1445);
nand U4788 (N_4788,In_1860,In_674);
nor U4789 (N_4789,In_249,In_372);
or U4790 (N_4790,In_842,In_672);
nor U4791 (N_4791,In_74,In_59);
and U4792 (N_4792,In_181,In_1708);
nor U4793 (N_4793,In_1849,In_517);
nor U4794 (N_4794,In_167,In_1095);
or U4795 (N_4795,In_804,In_442);
nand U4796 (N_4796,In_40,In_858);
or U4797 (N_4797,In_1262,In_618);
nor U4798 (N_4798,In_1898,In_796);
and U4799 (N_4799,In_1597,In_1397);
nor U4800 (N_4800,In_883,In_662);
and U4801 (N_4801,In_786,In_654);
and U4802 (N_4802,In_1025,In_1537);
nor U4803 (N_4803,In_1771,In_1243);
nor U4804 (N_4804,In_1230,In_1848);
and U4805 (N_4805,In_1640,In_1270);
or U4806 (N_4806,In_1928,In_378);
or U4807 (N_4807,In_639,In_1288);
or U4808 (N_4808,In_1249,In_487);
and U4809 (N_4809,In_1422,In_1656);
nand U4810 (N_4810,In_566,In_1074);
and U4811 (N_4811,In_1533,In_1702);
nor U4812 (N_4812,In_1324,In_1259);
and U4813 (N_4813,In_1943,In_1709);
xnor U4814 (N_4814,In_1220,In_103);
nor U4815 (N_4815,In_273,In_1141);
and U4816 (N_4816,In_656,In_1435);
and U4817 (N_4817,In_379,In_1503);
nand U4818 (N_4818,In_1321,In_1152);
or U4819 (N_4819,In_610,In_1678);
or U4820 (N_4820,In_1744,In_1571);
and U4821 (N_4821,In_88,In_1102);
and U4822 (N_4822,In_1955,In_60);
nand U4823 (N_4823,In_1295,In_1011);
nor U4824 (N_4824,In_383,In_1947);
nor U4825 (N_4825,In_1397,In_713);
nand U4826 (N_4826,In_685,In_1595);
or U4827 (N_4827,In_34,In_988);
nor U4828 (N_4828,In_543,In_74);
nand U4829 (N_4829,In_773,In_224);
nor U4830 (N_4830,In_451,In_1370);
nor U4831 (N_4831,In_932,In_52);
nand U4832 (N_4832,In_1665,In_251);
nor U4833 (N_4833,In_633,In_1652);
nand U4834 (N_4834,In_760,In_227);
nor U4835 (N_4835,In_1347,In_1630);
nand U4836 (N_4836,In_91,In_885);
and U4837 (N_4837,In_246,In_1033);
nand U4838 (N_4838,In_1500,In_450);
and U4839 (N_4839,In_1812,In_453);
nor U4840 (N_4840,In_997,In_131);
nand U4841 (N_4841,In_1138,In_1187);
nand U4842 (N_4842,In_945,In_1229);
or U4843 (N_4843,In_354,In_1083);
nor U4844 (N_4844,In_405,In_1203);
or U4845 (N_4845,In_151,In_173);
nand U4846 (N_4846,In_360,In_1093);
or U4847 (N_4847,In_1997,In_1277);
nand U4848 (N_4848,In_60,In_1324);
and U4849 (N_4849,In_501,In_1832);
or U4850 (N_4850,In_261,In_51);
nor U4851 (N_4851,In_1638,In_220);
nand U4852 (N_4852,In_669,In_1876);
and U4853 (N_4853,In_485,In_1530);
nand U4854 (N_4854,In_234,In_260);
nor U4855 (N_4855,In_1424,In_520);
nand U4856 (N_4856,In_44,In_1394);
nand U4857 (N_4857,In_1419,In_496);
and U4858 (N_4858,In_1150,In_330);
or U4859 (N_4859,In_439,In_1398);
or U4860 (N_4860,In_296,In_55);
or U4861 (N_4861,In_156,In_1538);
nand U4862 (N_4862,In_1187,In_185);
nor U4863 (N_4863,In_1771,In_1302);
nor U4864 (N_4864,In_1201,In_1370);
nor U4865 (N_4865,In_1424,In_1323);
and U4866 (N_4866,In_499,In_493);
and U4867 (N_4867,In_97,In_515);
xor U4868 (N_4868,In_1482,In_1551);
nor U4869 (N_4869,In_1489,In_1467);
nand U4870 (N_4870,In_738,In_1081);
nor U4871 (N_4871,In_612,In_305);
nand U4872 (N_4872,In_159,In_470);
nor U4873 (N_4873,In_493,In_1983);
nor U4874 (N_4874,In_304,In_1318);
nand U4875 (N_4875,In_1791,In_1073);
nand U4876 (N_4876,In_250,In_1198);
nand U4877 (N_4877,In_1075,In_1954);
and U4878 (N_4878,In_64,In_1836);
nand U4879 (N_4879,In_225,In_747);
and U4880 (N_4880,In_513,In_473);
nor U4881 (N_4881,In_418,In_824);
nor U4882 (N_4882,In_1750,In_1674);
nand U4883 (N_4883,In_410,In_40);
and U4884 (N_4884,In_1112,In_1367);
nor U4885 (N_4885,In_519,In_356);
nor U4886 (N_4886,In_819,In_1788);
nand U4887 (N_4887,In_143,In_377);
or U4888 (N_4888,In_1806,In_903);
and U4889 (N_4889,In_103,In_1769);
and U4890 (N_4890,In_295,In_485);
and U4891 (N_4891,In_1352,In_572);
or U4892 (N_4892,In_1066,In_383);
and U4893 (N_4893,In_347,In_816);
nor U4894 (N_4894,In_12,In_1709);
or U4895 (N_4895,In_1858,In_1095);
nand U4896 (N_4896,In_471,In_1833);
nand U4897 (N_4897,In_268,In_791);
and U4898 (N_4898,In_107,In_1253);
nor U4899 (N_4899,In_580,In_1662);
nand U4900 (N_4900,In_1322,In_769);
nor U4901 (N_4901,In_1553,In_1694);
nand U4902 (N_4902,In_1675,In_233);
or U4903 (N_4903,In_1417,In_739);
nand U4904 (N_4904,In_582,In_1371);
or U4905 (N_4905,In_928,In_1821);
or U4906 (N_4906,In_1890,In_1533);
nor U4907 (N_4907,In_1863,In_751);
nand U4908 (N_4908,In_1267,In_111);
nor U4909 (N_4909,In_1852,In_959);
or U4910 (N_4910,In_1229,In_585);
and U4911 (N_4911,In_1190,In_86);
nand U4912 (N_4912,In_1125,In_1662);
nand U4913 (N_4913,In_1865,In_775);
nand U4914 (N_4914,In_1348,In_1277);
nor U4915 (N_4915,In_84,In_289);
or U4916 (N_4916,In_523,In_1867);
nor U4917 (N_4917,In_640,In_691);
nand U4918 (N_4918,In_1854,In_821);
and U4919 (N_4919,In_1933,In_1462);
nor U4920 (N_4920,In_530,In_1903);
or U4921 (N_4921,In_1404,In_1946);
nand U4922 (N_4922,In_531,In_210);
nor U4923 (N_4923,In_1768,In_1278);
nand U4924 (N_4924,In_1085,In_114);
nand U4925 (N_4925,In_953,In_201);
and U4926 (N_4926,In_1992,In_616);
nand U4927 (N_4927,In_1815,In_86);
or U4928 (N_4928,In_189,In_973);
and U4929 (N_4929,In_1695,In_1387);
or U4930 (N_4930,In_1109,In_783);
nor U4931 (N_4931,In_1257,In_1428);
nor U4932 (N_4932,In_1296,In_1505);
nor U4933 (N_4933,In_1376,In_1641);
nor U4934 (N_4934,In_63,In_743);
nand U4935 (N_4935,In_541,In_259);
or U4936 (N_4936,In_1645,In_1148);
or U4937 (N_4937,In_363,In_1520);
xor U4938 (N_4938,In_1180,In_443);
nor U4939 (N_4939,In_1546,In_1583);
and U4940 (N_4940,In_624,In_511);
nand U4941 (N_4941,In_1103,In_647);
nor U4942 (N_4942,In_1271,In_42);
nand U4943 (N_4943,In_1429,In_908);
nor U4944 (N_4944,In_957,In_1739);
nand U4945 (N_4945,In_1144,In_1085);
or U4946 (N_4946,In_1491,In_974);
nor U4947 (N_4947,In_1805,In_418);
nor U4948 (N_4948,In_1382,In_1274);
or U4949 (N_4949,In_30,In_730);
and U4950 (N_4950,In_1265,In_1978);
nand U4951 (N_4951,In_1988,In_36);
nand U4952 (N_4952,In_419,In_1261);
or U4953 (N_4953,In_355,In_80);
or U4954 (N_4954,In_327,In_764);
nor U4955 (N_4955,In_349,In_850);
or U4956 (N_4956,In_682,In_1393);
and U4957 (N_4957,In_1111,In_1713);
nand U4958 (N_4958,In_1297,In_1752);
nand U4959 (N_4959,In_357,In_1046);
nor U4960 (N_4960,In_1036,In_96);
nand U4961 (N_4961,In_464,In_1203);
nor U4962 (N_4962,In_1360,In_1865);
or U4963 (N_4963,In_124,In_476);
and U4964 (N_4964,In_738,In_773);
nand U4965 (N_4965,In_522,In_935);
and U4966 (N_4966,In_1916,In_1162);
nand U4967 (N_4967,In_1656,In_231);
or U4968 (N_4968,In_1653,In_852);
or U4969 (N_4969,In_815,In_589);
or U4970 (N_4970,In_1051,In_1868);
and U4971 (N_4971,In_296,In_67);
nand U4972 (N_4972,In_557,In_1446);
nor U4973 (N_4973,In_1794,In_650);
nand U4974 (N_4974,In_338,In_1245);
nor U4975 (N_4975,In_968,In_11);
nor U4976 (N_4976,In_799,In_779);
nand U4977 (N_4977,In_1303,In_810);
or U4978 (N_4978,In_805,In_1891);
and U4979 (N_4979,In_1525,In_54);
and U4980 (N_4980,In_387,In_490);
nand U4981 (N_4981,In_1307,In_129);
or U4982 (N_4982,In_1144,In_203);
nor U4983 (N_4983,In_1442,In_1663);
nor U4984 (N_4984,In_1532,In_1977);
nor U4985 (N_4985,In_1157,In_641);
nand U4986 (N_4986,In_255,In_1403);
or U4987 (N_4987,In_473,In_1243);
or U4988 (N_4988,In_233,In_1093);
nand U4989 (N_4989,In_283,In_1817);
or U4990 (N_4990,In_444,In_251);
nor U4991 (N_4991,In_838,In_1821);
and U4992 (N_4992,In_1120,In_1552);
or U4993 (N_4993,In_185,In_1396);
and U4994 (N_4994,In_1511,In_382);
nand U4995 (N_4995,In_440,In_1854);
or U4996 (N_4996,In_1512,In_1393);
and U4997 (N_4997,In_1653,In_357);
nor U4998 (N_4998,In_624,In_1886);
nor U4999 (N_4999,In_1270,In_728);
or U5000 (N_5000,N_2445,N_3368);
nor U5001 (N_5001,N_4353,N_1330);
or U5002 (N_5002,N_1458,N_128);
and U5003 (N_5003,N_3315,N_2208);
nand U5004 (N_5004,N_3774,N_3538);
or U5005 (N_5005,N_4345,N_1114);
nand U5006 (N_5006,N_4973,N_436);
and U5007 (N_5007,N_3151,N_322);
nand U5008 (N_5008,N_3299,N_874);
and U5009 (N_5009,N_3044,N_2685);
xnor U5010 (N_5010,N_4179,N_1542);
or U5011 (N_5011,N_3174,N_3262);
nor U5012 (N_5012,N_234,N_2090);
and U5013 (N_5013,N_38,N_33);
and U5014 (N_5014,N_893,N_1573);
nand U5015 (N_5015,N_4857,N_1028);
nand U5016 (N_5016,N_2953,N_4934);
or U5017 (N_5017,N_1534,N_829);
nor U5018 (N_5018,N_2331,N_4758);
and U5019 (N_5019,N_2518,N_4062);
or U5020 (N_5020,N_2059,N_3935);
nand U5021 (N_5021,N_184,N_2880);
nor U5022 (N_5022,N_1996,N_4279);
nor U5023 (N_5023,N_1860,N_3693);
and U5024 (N_5024,N_3097,N_2310);
or U5025 (N_5025,N_3212,N_535);
nand U5026 (N_5026,N_2359,N_1570);
nand U5027 (N_5027,N_434,N_4595);
nand U5028 (N_5028,N_883,N_1313);
nor U5029 (N_5029,N_2302,N_1483);
nor U5030 (N_5030,N_3829,N_1641);
or U5031 (N_5031,N_4634,N_2329);
nor U5032 (N_5032,N_208,N_196);
or U5033 (N_5033,N_3851,N_1557);
nor U5034 (N_5034,N_3766,N_1985);
nor U5035 (N_5035,N_4391,N_1096);
nor U5036 (N_5036,N_4061,N_812);
nor U5037 (N_5037,N_2636,N_4892);
or U5038 (N_5038,N_4356,N_1283);
nand U5039 (N_5039,N_1648,N_4814);
or U5040 (N_5040,N_2525,N_4026);
nor U5041 (N_5041,N_4178,N_3127);
nor U5042 (N_5042,N_3796,N_2731);
nor U5043 (N_5043,N_4464,N_485);
and U5044 (N_5044,N_1270,N_204);
or U5045 (N_5045,N_2157,N_1060);
nand U5046 (N_5046,N_563,N_3028);
nand U5047 (N_5047,N_3780,N_3902);
nand U5048 (N_5048,N_3920,N_517);
or U5049 (N_5049,N_532,N_59);
or U5050 (N_5050,N_2749,N_578);
nor U5051 (N_5051,N_932,N_978);
nor U5052 (N_5052,N_2630,N_1245);
or U5053 (N_5053,N_3257,N_1309);
nor U5054 (N_5054,N_2999,N_4381);
and U5055 (N_5055,N_4565,N_2514);
or U5056 (N_5056,N_815,N_1740);
and U5057 (N_5057,N_2725,N_2714);
or U5058 (N_5058,N_3997,N_1590);
or U5059 (N_5059,N_2404,N_4905);
nand U5060 (N_5060,N_4534,N_4871);
or U5061 (N_5061,N_92,N_4710);
or U5062 (N_5062,N_3995,N_280);
xor U5063 (N_5063,N_826,N_2798);
and U5064 (N_5064,N_9,N_4306);
and U5065 (N_5065,N_401,N_2893);
and U5066 (N_5066,N_2479,N_1386);
and U5067 (N_5067,N_3624,N_2361);
and U5068 (N_5068,N_2146,N_2357);
nor U5069 (N_5069,N_4517,N_65);
nor U5070 (N_5070,N_415,N_1835);
or U5071 (N_5071,N_4006,N_199);
nand U5072 (N_5072,N_4466,N_1999);
or U5073 (N_5073,N_894,N_3053);
or U5074 (N_5074,N_3584,N_1861);
nand U5075 (N_5075,N_1136,N_319);
nand U5076 (N_5076,N_3977,N_3561);
xnor U5077 (N_5077,N_1705,N_1549);
nor U5078 (N_5078,N_304,N_3265);
or U5079 (N_5079,N_1672,N_2495);
or U5080 (N_5080,N_2571,N_2307);
or U5081 (N_5081,N_242,N_3704);
nor U5082 (N_5082,N_1525,N_887);
or U5083 (N_5083,N_4294,N_2784);
or U5084 (N_5084,N_2759,N_1919);
nand U5085 (N_5085,N_4716,N_3905);
or U5086 (N_5086,N_3122,N_1217);
nand U5087 (N_5087,N_1457,N_382);
and U5088 (N_5088,N_810,N_337);
or U5089 (N_5089,N_2425,N_3923);
nand U5090 (N_5090,N_1061,N_170);
xnor U5091 (N_5091,N_155,N_2552);
and U5092 (N_5092,N_3404,N_3399);
or U5093 (N_5093,N_3745,N_3638);
or U5094 (N_5094,N_2114,N_4722);
and U5095 (N_5095,N_3047,N_2596);
or U5096 (N_5096,N_808,N_4131);
nand U5097 (N_5097,N_4095,N_1250);
nand U5098 (N_5098,N_263,N_1156);
nor U5099 (N_5099,N_4352,N_4874);
or U5100 (N_5100,N_254,N_3732);
nor U5101 (N_5101,N_3447,N_198);
and U5102 (N_5102,N_1165,N_4756);
and U5103 (N_5103,N_3383,N_716);
nand U5104 (N_5104,N_2494,N_3654);
nor U5105 (N_5105,N_3585,N_406);
and U5106 (N_5106,N_3754,N_2997);
or U5107 (N_5107,N_10,N_2292);
nor U5108 (N_5108,N_3489,N_4024);
nand U5109 (N_5109,N_1361,N_1868);
nand U5110 (N_5110,N_570,N_1108);
nor U5111 (N_5111,N_1410,N_1888);
nor U5112 (N_5112,N_2619,N_1034);
and U5113 (N_5113,N_2073,N_2907);
and U5114 (N_5114,N_3221,N_853);
nand U5115 (N_5115,N_880,N_843);
and U5116 (N_5116,N_2794,N_2649);
xnor U5117 (N_5117,N_4937,N_3778);
nor U5118 (N_5118,N_4719,N_630);
or U5119 (N_5119,N_1427,N_2804);
nor U5120 (N_5120,N_4043,N_1703);
or U5121 (N_5121,N_3305,N_4658);
nor U5122 (N_5122,N_2177,N_4358);
nor U5123 (N_5123,N_3990,N_2720);
or U5124 (N_5124,N_1638,N_2593);
nor U5125 (N_5125,N_1463,N_3444);
or U5126 (N_5126,N_4745,N_4388);
nor U5127 (N_5127,N_2904,N_4718);
or U5128 (N_5128,N_4695,N_1857);
or U5129 (N_5129,N_1310,N_135);
nor U5130 (N_5130,N_1091,N_4056);
nor U5131 (N_5131,N_2344,N_2612);
or U5132 (N_5132,N_4673,N_742);
or U5133 (N_5133,N_470,N_4876);
nand U5134 (N_5134,N_3026,N_539);
nor U5135 (N_5135,N_2850,N_1097);
and U5136 (N_5136,N_2456,N_2155);
nand U5137 (N_5137,N_452,N_1223);
or U5138 (N_5138,N_425,N_407);
or U5139 (N_5139,N_456,N_2186);
nand U5140 (N_5140,N_4399,N_4834);
nand U5141 (N_5141,N_4766,N_4791);
nand U5142 (N_5142,N_2046,N_4980);
and U5143 (N_5143,N_3973,N_3093);
nor U5144 (N_5144,N_4645,N_3471);
and U5145 (N_5145,N_2278,N_423);
or U5146 (N_5146,N_3244,N_3750);
and U5147 (N_5147,N_4370,N_3901);
nand U5148 (N_5148,N_3854,N_4193);
nor U5149 (N_5149,N_1897,N_1571);
nor U5150 (N_5150,N_3335,N_3338);
xor U5151 (N_5151,N_841,N_992);
nand U5152 (N_5152,N_3464,N_3075);
or U5153 (N_5153,N_246,N_4096);
nand U5154 (N_5154,N_4480,N_4371);
and U5155 (N_5155,N_4495,N_4210);
or U5156 (N_5156,N_1013,N_3574);
nand U5157 (N_5157,N_938,N_1538);
nand U5158 (N_5158,N_2625,N_981);
nand U5159 (N_5159,N_4474,N_1170);
nor U5160 (N_5160,N_3862,N_1247);
or U5161 (N_5161,N_4,N_4623);
and U5162 (N_5162,N_4514,N_3481);
or U5163 (N_5163,N_1141,N_2451);
nand U5164 (N_5164,N_2283,N_4827);
nor U5165 (N_5165,N_1065,N_4962);
nor U5166 (N_5166,N_1986,N_3631);
nor U5167 (N_5167,N_4494,N_21);
and U5168 (N_5168,N_2573,N_3222);
nand U5169 (N_5169,N_685,N_4802);
or U5170 (N_5170,N_1294,N_1143);
or U5171 (N_5171,N_1948,N_2504);
nor U5172 (N_5172,N_2094,N_2860);
nand U5173 (N_5173,N_1117,N_437);
or U5174 (N_5174,N_2556,N_2449);
and U5175 (N_5175,N_2005,N_362);
and U5176 (N_5176,N_3791,N_1314);
nor U5177 (N_5177,N_2841,N_2528);
and U5178 (N_5178,N_1653,N_4203);
nand U5179 (N_5179,N_2818,N_2297);
or U5180 (N_5180,N_422,N_1788);
nor U5181 (N_5181,N_4038,N_596);
nor U5182 (N_5182,N_1846,N_1907);
nor U5183 (N_5183,N_1526,N_4420);
and U5184 (N_5184,N_1135,N_4487);
nor U5185 (N_5185,N_1295,N_4031);
nand U5186 (N_5186,N_4458,N_62);
nor U5187 (N_5187,N_3559,N_3996);
or U5188 (N_5188,N_2866,N_4740);
nand U5189 (N_5189,N_3485,N_1558);
nor U5190 (N_5190,N_232,N_4418);
or U5191 (N_5191,N_958,N_317);
nand U5192 (N_5192,N_2767,N_1654);
and U5193 (N_5193,N_595,N_2092);
and U5194 (N_5194,N_4106,N_600);
or U5195 (N_5195,N_4245,N_3168);
nor U5196 (N_5196,N_3915,N_1145);
nand U5197 (N_5197,N_1731,N_635);
nand U5198 (N_5198,N_3595,N_269);
or U5199 (N_5199,N_438,N_3325);
nand U5200 (N_5200,N_4460,N_1515);
nor U5201 (N_5201,N_136,N_4950);
or U5202 (N_5202,N_573,N_1406);
and U5203 (N_5203,N_230,N_3885);
and U5204 (N_5204,N_2032,N_1915);
nand U5205 (N_5205,N_2041,N_1190);
or U5206 (N_5206,N_753,N_4362);
or U5207 (N_5207,N_4894,N_3196);
and U5208 (N_5208,N_2864,N_3562);
nor U5209 (N_5209,N_378,N_1337);
and U5210 (N_5210,N_706,N_4259);
and U5211 (N_5211,N_4145,N_763);
and U5212 (N_5212,N_256,N_348);
or U5213 (N_5213,N_3579,N_2805);
nor U5214 (N_5214,N_1767,N_3301);
nor U5215 (N_5215,N_1658,N_409);
nor U5216 (N_5216,N_4948,N_367);
nor U5217 (N_5217,N_4800,N_1914);
nand U5218 (N_5218,N_1029,N_2311);
nand U5219 (N_5219,N_4676,N_3674);
nand U5220 (N_5220,N_4715,N_478);
and U5221 (N_5221,N_3435,N_2234);
nor U5222 (N_5222,N_4723,N_744);
and U5223 (N_5223,N_2959,N_1210);
and U5224 (N_5224,N_3869,N_3176);
nor U5225 (N_5225,N_2730,N_1299);
and U5226 (N_5226,N_2586,N_4515);
nor U5227 (N_5227,N_2658,N_849);
nand U5228 (N_5228,N_1485,N_3123);
or U5229 (N_5229,N_686,N_1104);
or U5230 (N_5230,N_3298,N_2611);
and U5231 (N_5231,N_3040,N_4152);
or U5232 (N_5232,N_2539,N_4562);
nor U5233 (N_5233,N_3879,N_4496);
nor U5234 (N_5234,N_4530,N_1784);
and U5235 (N_5235,N_2626,N_1886);
nand U5236 (N_5236,N_4700,N_2130);
xor U5237 (N_5237,N_440,N_2168);
nand U5238 (N_5238,N_3458,N_1043);
nor U5239 (N_5239,N_179,N_1875);
nor U5240 (N_5240,N_4955,N_4432);
nand U5241 (N_5241,N_3794,N_2640);
nor U5242 (N_5242,N_1883,N_661);
and U5243 (N_5243,N_498,N_2238);
nand U5244 (N_5244,N_2567,N_4153);
and U5245 (N_5245,N_2948,N_4180);
or U5246 (N_5246,N_2624,N_3492);
nor U5247 (N_5247,N_2915,N_1271);
or U5248 (N_5248,N_4188,N_2549);
nand U5249 (N_5249,N_3177,N_521);
or U5250 (N_5250,N_3119,N_3596);
nor U5251 (N_5251,N_399,N_3319);
nor U5252 (N_5252,N_2692,N_4198);
and U5253 (N_5253,N_2373,N_1514);
or U5254 (N_5254,N_1377,N_351);
xor U5255 (N_5255,N_231,N_987);
nor U5256 (N_5256,N_4709,N_3259);
and U5257 (N_5257,N_3455,N_457);
nor U5258 (N_5258,N_3645,N_780);
nand U5259 (N_5259,N_446,N_3252);
nor U5260 (N_5260,N_4606,N_2647);
nand U5261 (N_5261,N_2418,N_3573);
nor U5262 (N_5262,N_2162,N_2365);
nor U5263 (N_5263,N_2068,N_3353);
nand U5264 (N_5264,N_4521,N_377);
and U5265 (N_5265,N_3924,N_607);
and U5266 (N_5266,N_1578,N_3436);
nand U5267 (N_5267,N_3088,N_2763);
or U5268 (N_5268,N_4736,N_173);
nand U5269 (N_5269,N_4143,N_875);
nand U5270 (N_5270,N_2231,N_3022);
or U5271 (N_5271,N_4412,N_628);
nor U5272 (N_5272,N_140,N_3032);
nand U5273 (N_5273,N_145,N_1089);
and U5274 (N_5274,N_1216,N_4071);
nor U5275 (N_5275,N_166,N_1083);
nand U5276 (N_5276,N_4239,N_1496);
nand U5277 (N_5277,N_3872,N_3651);
nand U5278 (N_5278,N_3812,N_4271);
or U5279 (N_5279,N_814,N_4942);
or U5280 (N_5280,N_416,N_649);
nand U5281 (N_5281,N_2016,N_1470);
nor U5282 (N_5282,N_1338,N_1711);
and U5283 (N_5283,N_3466,N_1172);
nand U5284 (N_5284,N_3618,N_633);
and U5285 (N_5285,N_2751,N_1841);
nor U5286 (N_5286,N_4435,N_4342);
or U5287 (N_5287,N_286,N_3139);
or U5288 (N_5288,N_2239,N_2216);
nand U5289 (N_5289,N_4385,N_3856);
nand U5290 (N_5290,N_1805,N_2729);
and U5291 (N_5291,N_844,N_3999);
and U5292 (N_5292,N_2289,N_3684);
nand U5293 (N_5293,N_4256,N_2204);
nor U5294 (N_5294,N_366,N_2812);
and U5295 (N_5295,N_4073,N_268);
and U5296 (N_5296,N_2847,N_3472);
nand U5297 (N_5297,N_872,N_293);
nand U5298 (N_5298,N_4448,N_3577);
nand U5299 (N_5299,N_2657,N_2741);
or U5300 (N_5300,N_281,N_432);
nand U5301 (N_5301,N_1062,N_3217);
nor U5302 (N_5302,N_2064,N_2656);
nand U5303 (N_5303,N_1481,N_1808);
nand U5304 (N_5304,N_2437,N_2172);
or U5305 (N_5305,N_4215,N_683);
nor U5306 (N_5306,N_1021,N_1036);
or U5307 (N_5307,N_25,N_4251);
nor U5308 (N_5308,N_3179,N_2034);
nand U5309 (N_5309,N_1246,N_3895);
and U5310 (N_5310,N_945,N_610);
nor U5311 (N_5311,N_2367,N_4670);
nor U5312 (N_5312,N_395,N_3586);
and U5313 (N_5313,N_2050,N_3756);
and U5314 (N_5314,N_3340,N_2512);
nand U5315 (N_5315,N_560,N_3101);
or U5316 (N_5316,N_4675,N_4925);
nand U5317 (N_5317,N_2536,N_2591);
nor U5318 (N_5318,N_76,N_4126);
nor U5319 (N_5319,N_3509,N_2564);
and U5320 (N_5320,N_3083,N_1012);
and U5321 (N_5321,N_2855,N_4442);
and U5322 (N_5322,N_1824,N_3271);
or U5323 (N_5323,N_2927,N_4777);
or U5324 (N_5324,N_4255,N_1231);
nor U5325 (N_5325,N_3676,N_4309);
and U5326 (N_5326,N_751,N_4683);
nand U5327 (N_5327,N_1011,N_3475);
nor U5328 (N_5328,N_3017,N_4053);
nand U5329 (N_5329,N_3129,N_205);
and U5330 (N_5330,N_964,N_2453);
nor U5331 (N_5331,N_3229,N_29);
and U5332 (N_5332,N_4429,N_1370);
nand U5333 (N_5333,N_174,N_3884);
and U5334 (N_5334,N_2432,N_102);
nor U5335 (N_5335,N_1848,N_2533);
nand U5336 (N_5336,N_1090,N_4473);
nor U5337 (N_5337,N_3072,N_3647);
nand U5338 (N_5338,N_3925,N_2957);
xnor U5339 (N_5339,N_3591,N_3260);
nand U5340 (N_5340,N_2677,N_4561);
or U5341 (N_5341,N_4396,N_1630);
and U5342 (N_5342,N_493,N_4621);
and U5343 (N_5343,N_2088,N_17);
and U5344 (N_5344,N_3006,N_2853);
nor U5345 (N_5345,N_2538,N_3051);
nor U5346 (N_5346,N_4401,N_2808);
and U5347 (N_5347,N_969,N_3507);
nand U5348 (N_5348,N_2584,N_163);
nand U5349 (N_5349,N_2403,N_3133);
nand U5350 (N_5350,N_91,N_1042);
or U5351 (N_5351,N_1844,N_3109);
and U5352 (N_5352,N_836,N_183);
nand U5353 (N_5353,N_1635,N_2985);
and U5354 (N_5354,N_1344,N_408);
and U5355 (N_5355,N_2515,N_2682);
and U5356 (N_5356,N_2315,N_1288);
or U5357 (N_5357,N_3891,N_1580);
nor U5358 (N_5358,N_4292,N_4235);
or U5359 (N_5359,N_4949,N_1939);
or U5360 (N_5360,N_4619,N_1823);
nor U5361 (N_5361,N_1044,N_599);
nor U5362 (N_5362,N_4246,N_424);
xnor U5363 (N_5363,N_4602,N_4105);
nor U5364 (N_5364,N_2127,N_2594);
or U5365 (N_5365,N_2683,N_1292);
nand U5366 (N_5366,N_3437,N_1119);
nand U5367 (N_5367,N_2883,N_813);
nor U5368 (N_5368,N_1284,N_3822);
nand U5369 (N_5369,N_3300,N_4818);
and U5370 (N_5370,N_902,N_1656);
or U5371 (N_5371,N_1945,N_3570);
and U5372 (N_5372,N_1148,N_764);
or U5373 (N_5373,N_3148,N_307);
nor U5374 (N_5374,N_335,N_2977);
nand U5375 (N_5375,N_2223,N_1647);
or U5376 (N_5376,N_2415,N_2668);
or U5377 (N_5377,N_2503,N_4360);
nand U5378 (N_5378,N_1388,N_4705);
or U5379 (N_5379,N_387,N_701);
nor U5380 (N_5380,N_3132,N_2220);
nor U5381 (N_5381,N_3959,N_1780);
or U5382 (N_5382,N_2422,N_2551);
and U5383 (N_5383,N_2387,N_326);
nand U5384 (N_5384,N_2643,N_2752);
nand U5385 (N_5385,N_4632,N_3427);
and U5386 (N_5386,N_889,N_2711);
nand U5387 (N_5387,N_914,N_299);
nor U5388 (N_5388,N_1955,N_4446);
and U5389 (N_5389,N_2305,N_698);
or U5390 (N_5390,N_3204,N_4733);
nor U5391 (N_5391,N_990,N_1430);
nand U5392 (N_5392,N_2230,N_1432);
and U5393 (N_5393,N_4783,N_4017);
nor U5394 (N_5394,N_13,N_704);
nand U5395 (N_5395,N_2378,N_2994);
nor U5396 (N_5396,N_3571,N_1191);
nor U5397 (N_5397,N_1686,N_143);
and U5398 (N_5398,N_703,N_555);
nand U5399 (N_5399,N_3663,N_1679);
or U5400 (N_5400,N_508,N_4574);
nand U5401 (N_5401,N_4826,N_3508);
nand U5402 (N_5402,N_3728,N_1959);
nor U5403 (N_5403,N_4679,N_4486);
xor U5404 (N_5404,N_360,N_3598);
nor U5405 (N_5405,N_3825,N_3166);
nand U5406 (N_5406,N_122,N_3276);
and U5407 (N_5407,N_1462,N_1379);
nand U5408 (N_5408,N_4626,N_3459);
and U5409 (N_5409,N_4859,N_386);
nand U5410 (N_5410,N_2398,N_4540);
and U5411 (N_5411,N_2644,N_4076);
or U5412 (N_5412,N_4406,N_916);
or U5413 (N_5413,N_4118,N_4384);
nor U5414 (N_5414,N_585,N_3327);
nor U5415 (N_5415,N_4582,N_1278);
and U5416 (N_5416,N_711,N_4628);
or U5417 (N_5417,N_3701,N_3978);
nand U5418 (N_5418,N_3374,N_1152);
nand U5419 (N_5419,N_19,N_4433);
and U5420 (N_5420,N_1659,N_329);
or U5421 (N_5421,N_855,N_3033);
nor U5422 (N_5422,N_627,N_638);
nor U5423 (N_5423,N_3543,N_3474);
nand U5424 (N_5424,N_2910,N_4436);
and U5425 (N_5425,N_4421,N_612);
nor U5426 (N_5426,N_2793,N_1080);
nand U5427 (N_5427,N_3253,N_2136);
nor U5428 (N_5428,N_3566,N_777);
nand U5429 (N_5429,N_4699,N_2074);
nand U5430 (N_5430,N_1545,N_2859);
nand U5431 (N_5431,N_2213,N_3410);
nand U5432 (N_5432,N_1963,N_1650);
nand U5433 (N_5433,N_2832,N_420);
and U5434 (N_5434,N_3429,N_2086);
or U5435 (N_5435,N_1277,N_2576);
or U5436 (N_5436,N_1921,N_2782);
or U5437 (N_5437,N_4763,N_860);
nor U5438 (N_5438,N_4267,N_4354);
nand U5439 (N_5439,N_3324,N_1990);
and U5440 (N_5440,N_88,N_3289);
and U5441 (N_5441,N_1768,N_2955);
nand U5442 (N_5442,N_3084,N_3930);
and U5443 (N_5443,N_3776,N_4469);
nand U5444 (N_5444,N_97,N_1842);
xnor U5445 (N_5445,N_2326,N_1567);
nand U5446 (N_5446,N_2330,N_1023);
nand U5447 (N_5447,N_591,N_3557);
or U5448 (N_5448,N_379,N_1159);
or U5449 (N_5449,N_3548,N_3483);
nand U5450 (N_5450,N_4539,N_1508);
and U5451 (N_5451,N_3535,N_3066);
and U5452 (N_5452,N_2700,N_516);
or U5453 (N_5453,N_3453,N_3671);
or U5454 (N_5454,N_4694,N_2060);
or U5455 (N_5455,N_684,N_3733);
and U5456 (N_5456,N_156,N_3295);
or U5457 (N_5457,N_2868,N_821);
nand U5458 (N_5458,N_2975,N_4021);
nand U5459 (N_5459,N_1287,N_4008);
and U5460 (N_5460,N_3894,N_3232);
nor U5461 (N_5461,N_2116,N_2627);
and U5462 (N_5462,N_3734,N_4302);
nor U5463 (N_5463,N_3981,N_977);
or U5464 (N_5464,N_4046,N_1750);
nand U5465 (N_5465,N_2147,N_106);
or U5466 (N_5466,N_3108,N_2488);
nand U5467 (N_5467,N_4732,N_3904);
nand U5468 (N_5468,N_3161,N_3608);
and U5469 (N_5469,N_939,N_4990);
or U5470 (N_5470,N_157,N_2062);
or U5471 (N_5471,N_4701,N_4638);
and U5472 (N_5472,N_3515,N_1282);
and U5473 (N_5473,N_2820,N_3782);
nor U5474 (N_5474,N_4727,N_1642);
and U5475 (N_5475,N_4033,N_2412);
or U5476 (N_5476,N_4347,N_1164);
nand U5477 (N_5477,N_3401,N_3802);
nand U5478 (N_5478,N_679,N_2608);
nor U5479 (N_5479,N_490,N_225);
or U5480 (N_5480,N_4842,N_3580);
and U5481 (N_5481,N_116,N_2651);
or U5482 (N_5482,N_581,N_3567);
and U5483 (N_5483,N_854,N_1499);
and U5484 (N_5484,N_4091,N_511);
or U5485 (N_5485,N_3149,N_2471);
and U5486 (N_5486,N_2544,N_1418);
nand U5487 (N_5487,N_4049,N_4535);
nand U5488 (N_5488,N_3405,N_2641);
or U5489 (N_5489,N_3355,N_1975);
nor U5490 (N_5490,N_4924,N_2843);
nor U5491 (N_5491,N_586,N_4513);
or U5492 (N_5492,N_3422,N_295);
or U5493 (N_5493,N_3815,N_1890);
or U5494 (N_5494,N_4069,N_1139);
nor U5495 (N_5495,N_2195,N_3100);
nand U5496 (N_5496,N_168,N_1826);
nand U5497 (N_5497,N_1436,N_736);
nor U5498 (N_5498,N_4417,N_3773);
nor U5499 (N_5499,N_383,N_4112);
or U5500 (N_5500,N_1372,N_1208);
nor U5501 (N_5501,N_2560,N_512);
nand U5502 (N_5502,N_4693,N_734);
or U5503 (N_5503,N_1866,N_819);
nor U5504 (N_5504,N_725,N_4324);
or U5505 (N_5505,N_1252,N_3560);
or U5506 (N_5506,N_4493,N_2835);
or U5507 (N_5507,N_4268,N_3589);
or U5508 (N_5508,N_1204,N_1285);
xor U5509 (N_5509,N_724,N_3758);
nand U5510 (N_5510,N_3424,N_2849);
nor U5511 (N_5511,N_4058,N_3980);
nor U5512 (N_5512,N_2267,N_4136);
nor U5513 (N_5513,N_3376,N_1810);
nor U5514 (N_5514,N_4672,N_39);
nor U5515 (N_5515,N_2779,N_1892);
nand U5516 (N_5516,N_2296,N_212);
and U5517 (N_5517,N_1429,N_2795);
and U5518 (N_5518,N_4790,N_1887);
nand U5519 (N_5519,N_3594,N_435);
nand U5520 (N_5520,N_3739,N_3012);
nor U5521 (N_5521,N_4314,N_2486);
and U5522 (N_5522,N_3683,N_2894);
nand U5523 (N_5523,N_192,N_3070);
and U5524 (N_5524,N_2395,N_4277);
nand U5525 (N_5525,N_2634,N_1049);
nand U5526 (N_5526,N_729,N_352);
and U5527 (N_5527,N_3991,N_741);
and U5528 (N_5528,N_126,N_354);
nor U5529 (N_5529,N_1193,N_1431);
or U5530 (N_5530,N_2746,N_2704);
or U5531 (N_5531,N_3803,N_770);
and U5532 (N_5532,N_3781,N_4372);
and U5533 (N_5533,N_4798,N_1966);
nor U5534 (N_5534,N_2941,N_1974);
or U5535 (N_5535,N_4537,N_748);
and U5536 (N_5536,N_1908,N_4221);
and U5537 (N_5537,N_1497,N_613);
xor U5538 (N_5538,N_4440,N_1220);
or U5539 (N_5539,N_2423,N_4951);
and U5540 (N_5540,N_3800,N_3394);
and U5541 (N_5541,N_2770,N_4724);
nor U5542 (N_5542,N_2566,N_864);
or U5543 (N_5543,N_2117,N_4116);
nor U5544 (N_5544,N_1550,N_1079);
or U5545 (N_5545,N_3344,N_2635);
and U5546 (N_5546,N_2246,N_851);
nor U5547 (N_5547,N_1614,N_4375);
nor U5548 (N_5548,N_4726,N_1205);
and U5549 (N_5549,N_3352,N_2645);
and U5550 (N_5550,N_2385,N_4443);
and U5551 (N_5551,N_2722,N_306);
nand U5552 (N_5552,N_2984,N_2210);
nand U5553 (N_5553,N_1577,N_3219);
or U5554 (N_5554,N_2582,N_2534);
or U5555 (N_5555,N_3117,N_4964);
or U5556 (N_5556,N_898,N_3198);
nor U5557 (N_5557,N_1618,N_1645);
nand U5558 (N_5558,N_258,N_873);
nand U5559 (N_5559,N_2595,N_2664);
nand U5560 (N_5560,N_265,N_3351);
nor U5561 (N_5561,N_4663,N_4484);
nand U5562 (N_5562,N_1770,N_3049);
or U5563 (N_5563,N_3349,N_4822);
or U5564 (N_5564,N_4079,N_4249);
nor U5565 (N_5565,N_3023,N_2708);
nor U5566 (N_5566,N_4836,N_624);
and U5567 (N_5567,N_3686,N_738);
and U5568 (N_5568,N_1140,N_7);
nor U5569 (N_5569,N_1318,N_4148);
nand U5570 (N_5570,N_828,N_4407);
nor U5571 (N_5571,N_2192,N_4927);
or U5572 (N_5572,N_2971,N_479);
or U5573 (N_5573,N_552,N_3581);
nand U5574 (N_5574,N_740,N_876);
and U5575 (N_5575,N_3656,N_99);
nor U5576 (N_5576,N_3922,N_865);
nand U5577 (N_5577,N_4797,N_655);
nor U5578 (N_5578,N_3860,N_2733);
nand U5579 (N_5579,N_3477,N_3411);
nor U5580 (N_5580,N_4500,N_2998);
nor U5581 (N_5581,N_3974,N_4004);
or U5582 (N_5582,N_1596,N_20);
nor U5583 (N_5583,N_1437,N_4533);
or U5584 (N_5584,N_1195,N_1964);
nand U5585 (N_5585,N_3789,N_1976);
nand U5586 (N_5586,N_3290,N_3539);
or U5587 (N_5587,N_4479,N_4788);
or U5588 (N_5588,N_260,N_111);
and U5589 (N_5589,N_4133,N_3003);
or U5590 (N_5590,N_4451,N_2198);
or U5591 (N_5591,N_3278,N_54);
nor U5592 (N_5592,N_3669,N_3824);
and U5593 (N_5593,N_358,N_915);
nor U5594 (N_5594,N_4346,N_4739);
and U5595 (N_5595,N_3971,N_4002);
nor U5596 (N_5596,N_2945,N_3450);
and U5597 (N_5597,N_1815,N_3388);
or U5598 (N_5598,N_1747,N_1173);
nor U5599 (N_5599,N_1275,N_1434);
nand U5600 (N_5600,N_4276,N_338);
or U5601 (N_5601,N_886,N_222);
nand U5602 (N_5602,N_2557,N_2235);
and U5603 (N_5603,N_2960,N_2602);
nand U5604 (N_5604,N_2099,N_3738);
nand U5605 (N_5605,N_1077,N_4899);
nor U5606 (N_5606,N_3081,N_2055);
nand U5607 (N_5607,N_1151,N_2067);
or U5608 (N_5608,N_1925,N_1859);
or U5609 (N_5609,N_3592,N_2021);
or U5610 (N_5610,N_235,N_2650);
nor U5611 (N_5611,N_1521,N_4817);
nand U5612 (N_5612,N_67,N_86);
nand U5613 (N_5613,N_428,N_4639);
or U5614 (N_5614,N_4839,N_3673);
nand U5615 (N_5615,N_4444,N_3857);
nor U5616 (N_5616,N_897,N_3587);
nand U5617 (N_5617,N_4080,N_1068);
or U5618 (N_5618,N_2732,N_4731);
nor U5619 (N_5619,N_1196,N_2141);
nor U5620 (N_5620,N_1734,N_4258);
and U5621 (N_5621,N_2426,N_3961);
nand U5622 (N_5622,N_2211,N_2477);
and U5623 (N_5623,N_1735,N_676);
nand U5624 (N_5624,N_4050,N_224);
or U5625 (N_5625,N_846,N_4281);
and U5626 (N_5626,N_1411,N_3220);
nor U5627 (N_5627,N_441,N_4671);
and U5628 (N_5628,N_1535,N_3367);
or U5629 (N_5629,N_100,N_1185);
and U5630 (N_5630,N_976,N_2085);
and U5631 (N_5631,N_1840,N_792);
or U5632 (N_5632,N_568,N_101);
and U5633 (N_5633,N_2616,N_3329);
nand U5634 (N_5634,N_831,N_660);
nand U5635 (N_5635,N_2040,N_2266);
and U5636 (N_5636,N_1778,N_2115);
nand U5637 (N_5637,N_4856,N_1174);
and U5638 (N_5638,N_623,N_1513);
or U5639 (N_5639,N_4953,N_3425);
or U5640 (N_5640,N_3926,N_4917);
and U5641 (N_5641,N_1069,N_3408);
nor U5642 (N_5642,N_4858,N_1527);
or U5643 (N_5643,N_1637,N_4481);
or U5644 (N_5644,N_3621,N_4902);
nand U5645 (N_5645,N_3498,N_4204);
and U5646 (N_5646,N_3960,N_4720);
and U5647 (N_5647,N_1358,N_2181);
or U5648 (N_5648,N_650,N_1257);
nand U5649 (N_5649,N_2293,N_1038);
and U5650 (N_5650,N_264,N_866);
nor U5651 (N_5651,N_4983,N_3644);
or U5652 (N_5652,N_14,N_2699);
or U5653 (N_5653,N_721,N_187);
nor U5654 (N_5654,N_1460,N_2838);
xor U5655 (N_5655,N_845,N_3966);
and U5656 (N_5656,N_3502,N_1594);
nand U5657 (N_5657,N_1423,N_4967);
or U5658 (N_5658,N_1994,N_2194);
nand U5659 (N_5659,N_1599,N_2530);
nor U5660 (N_5660,N_4339,N_1753);
nand U5661 (N_5661,N_691,N_4083);
nor U5662 (N_5662,N_1884,N_2338);
or U5663 (N_5663,N_4060,N_4146);
nand U5664 (N_5664,N_4243,N_4068);
nand U5665 (N_5665,N_2137,N_2947);
or U5666 (N_5666,N_81,N_1793);
nor U5667 (N_5667,N_4875,N_1063);
and U5668 (N_5668,N_4551,N_267);
or U5669 (N_5669,N_2459,N_1326);
nand U5670 (N_5670,N_2031,N_1585);
nand U5671 (N_5671,N_840,N_3691);
nand U5672 (N_5672,N_3821,N_161);
nand U5673 (N_5673,N_1180,N_1825);
and U5674 (N_5674,N_2813,N_4159);
and U5675 (N_5675,N_237,N_3238);
nor U5676 (N_5676,N_2084,N_4627);
and U5677 (N_5677,N_3415,N_4904);
nand U5678 (N_5678,N_1255,N_835);
nand U5679 (N_5679,N_2781,N_3223);
and U5680 (N_5680,N_4092,N_1749);
nor U5681 (N_5681,N_2342,N_1903);
and U5682 (N_5682,N_1487,N_4958);
xor U5683 (N_5683,N_1506,N_4378);
nand U5684 (N_5684,N_1830,N_2222);
or U5685 (N_5685,N_3460,N_1248);
nand U5686 (N_5686,N_4725,N_3568);
or U5687 (N_5687,N_4828,N_283);
nand U5688 (N_5688,N_4223,N_820);
or U5689 (N_5689,N_1522,N_2674);
nor U5690 (N_5690,N_2837,N_1607);
and U5691 (N_5691,N_2333,N_4684);
nor U5692 (N_5692,N_1723,N_1891);
nor U5693 (N_5693,N_2098,N_4508);
nor U5694 (N_5694,N_2930,N_1608);
or U5695 (N_5695,N_300,N_500);
or U5696 (N_5696,N_2681,N_364);
nor U5697 (N_5697,N_1009,N_2968);
nand U5698 (N_5698,N_261,N_3964);
nand U5699 (N_5699,N_4975,N_2811);
and U5700 (N_5700,N_2066,N_3231);
nor U5701 (N_5701,N_2207,N_1369);
nand U5702 (N_5702,N_3092,N_2473);
nand U5703 (N_5703,N_51,N_3180);
or U5704 (N_5704,N_2986,N_647);
nor U5705 (N_5705,N_3725,N_3942);
nand U5706 (N_5706,N_3115,N_2159);
and U5707 (N_5707,N_4222,N_2680);
and U5708 (N_5708,N_1562,N_2316);
nand U5709 (N_5709,N_1965,N_4018);
or U5710 (N_5710,N_3178,N_1307);
or U5711 (N_5711,N_2462,N_986);
or U5712 (N_5712,N_2701,N_2603);
or U5713 (N_5713,N_1507,N_4270);
nand U5714 (N_5714,N_3440,N_637);
nor U5715 (N_5715,N_4999,N_4845);
or U5716 (N_5716,N_3934,N_2491);
nor U5717 (N_5717,N_2498,N_483);
nand U5718 (N_5718,N_1092,N_4233);
and U5719 (N_5719,N_4714,N_3634);
nor U5720 (N_5720,N_3818,N_687);
or U5721 (N_5721,N_2938,N_967);
nand U5722 (N_5722,N_4007,N_3722);
nand U5723 (N_5723,N_2932,N_991);
and U5724 (N_5724,N_652,N_2191);
nand U5725 (N_5725,N_1509,N_1364);
nand U5726 (N_5726,N_1801,N_75);
and U5727 (N_5727,N_524,N_3706);
nand U5728 (N_5728,N_3903,N_737);
nor U5729 (N_5729,N_4933,N_2097);
and U5730 (N_5730,N_3529,N_1911);
and U5731 (N_5731,N_3830,N_47);
or U5732 (N_5732,N_903,N_2607);
and U5733 (N_5733,N_911,N_3378);
nand U5734 (N_5734,N_467,N_321);
and U5735 (N_5735,N_4355,N_3797);
or U5736 (N_5736,N_2007,N_4408);
nand U5737 (N_5737,N_947,N_132);
nor U5738 (N_5738,N_4185,N_1493);
nor U5739 (N_5739,N_23,N_4125);
or U5740 (N_5740,N_910,N_1213);
and U5741 (N_5741,N_3696,N_3848);
nor U5742 (N_5742,N_954,N_1572);
or U5743 (N_5743,N_2898,N_3152);
nand U5744 (N_5744,N_4931,N_1448);
xnor U5745 (N_5745,N_3147,N_1909);
or U5746 (N_5746,N_4556,N_4410);
or U5747 (N_5747,N_2718,N_1563);
nand U5748 (N_5748,N_3470,N_4334);
or U5749 (N_5749,N_3670,N_4301);
nor U5750 (N_5750,N_1234,N_2766);
and U5751 (N_5751,N_1566,N_4164);
nor U5752 (N_5752,N_1188,N_4113);
nor U5753 (N_5753,N_104,N_296);
nor U5754 (N_5754,N_1981,N_2169);
and U5755 (N_5755,N_2243,N_3927);
nor U5756 (N_5756,N_907,N_2642);
or U5757 (N_5757,N_3392,N_767);
or U5758 (N_5758,N_4690,N_3469);
or U5759 (N_5759,N_4109,N_529);
or U5760 (N_5760,N_3762,N_899);
or U5761 (N_5761,N_2863,N_4832);
or U5762 (N_5762,N_4465,N_4119);
nor U5763 (N_5763,N_4605,N_1315);
and U5764 (N_5764,N_3116,N_3909);
or U5765 (N_5765,N_4503,N_839);
or U5766 (N_5766,N_1343,N_985);
or U5767 (N_5767,N_3014,N_4819);
nand U5768 (N_5768,N_3866,N_3556);
and U5769 (N_5769,N_3658,N_663);
and U5770 (N_5770,N_688,N_994);
nor U5771 (N_5771,N_2870,N_2240);
nand U5772 (N_5772,N_3784,N_206);
and U5773 (N_5773,N_3685,N_4184);
nor U5774 (N_5774,N_1529,N_2424);
and U5775 (N_5775,N_1241,N_396);
nor U5776 (N_5776,N_3544,N_2577);
nand U5777 (N_5777,N_137,N_4527);
or U5778 (N_5778,N_779,N_3396);
nand U5779 (N_5779,N_1992,N_245);
or U5780 (N_5780,N_4231,N_707);
nor U5781 (N_5781,N_1777,N_2877);
or U5782 (N_5782,N_2775,N_1776);
nand U5783 (N_5783,N_1662,N_469);
nand U5784 (N_5784,N_3449,N_2970);
or U5785 (N_5785,N_2030,N_1345);
nor U5786 (N_5786,N_2940,N_3678);
nor U5787 (N_5787,N_3664,N_811);
or U5788 (N_5788,N_2830,N_2372);
or U5789 (N_5789,N_951,N_2973);
nor U5790 (N_5790,N_4988,N_3986);
and U5791 (N_5791,N_662,N_949);
and U5792 (N_5792,N_2184,N_4320);
nor U5793 (N_5793,N_1733,N_720);
or U5794 (N_5794,N_710,N_3813);
nor U5795 (N_5795,N_1484,N_1149);
and U5796 (N_5796,N_2600,N_4124);
nand U5797 (N_5797,N_3307,N_417);
or U5798 (N_5798,N_2416,N_4209);
nor U5799 (N_5799,N_2933,N_1833);
nor U5800 (N_5800,N_3173,N_1564);
and U5801 (N_5801,N_2056,N_404);
and U5802 (N_5802,N_4603,N_3167);
nand U5803 (N_5803,N_2723,N_1243);
nor U5804 (N_5804,N_2303,N_4173);
and U5805 (N_5805,N_1895,N_2807);
nor U5806 (N_5806,N_941,N_1237);
nand U5807 (N_5807,N_1748,N_2547);
nor U5808 (N_5808,N_774,N_3692);
and U5809 (N_5809,N_1206,N_1867);
nand U5810 (N_5810,N_3372,N_4000);
nand U5811 (N_5811,N_4289,N_1189);
nand U5812 (N_5812,N_2761,N_3695);
nor U5813 (N_5813,N_3192,N_3135);
nor U5814 (N_5814,N_850,N_499);
nand U5815 (N_5815,N_2075,N_2070);
and U5816 (N_5816,N_3735,N_4776);
and U5817 (N_5817,N_4274,N_31);
and U5818 (N_5818,N_2468,N_347);
or U5819 (N_5819,N_1098,N_2982);
nand U5820 (N_5820,N_4285,N_4037);
and U5821 (N_5821,N_291,N_2043);
nand U5822 (N_5822,N_3749,N_4728);
xor U5823 (N_5823,N_228,N_1633);
and U5824 (N_5824,N_2815,N_1905);
nand U5825 (N_5825,N_2317,N_3015);
and U5826 (N_5826,N_693,N_3690);
and U5827 (N_5827,N_3334,N_557);
nand U5828 (N_5828,N_2360,N_1371);
or U5829 (N_5829,N_2414,N_4891);
nand U5830 (N_5830,N_2306,N_130);
or U5831 (N_5831,N_447,N_4449);
nand U5832 (N_5832,N_3318,N_2819);
nand U5833 (N_5833,N_3779,N_85);
or U5834 (N_5834,N_4563,N_2814);
and U5835 (N_5835,N_2531,N_4266);
or U5836 (N_5836,N_657,N_3709);
nor U5837 (N_5837,N_2011,N_4335);
nor U5838 (N_5838,N_530,N_3530);
and U5839 (N_5839,N_2587,N_1904);
or U5840 (N_5840,N_2384,N_2284);
or U5841 (N_5841,N_3407,N_689);
and U5842 (N_5842,N_4290,N_3333);
nor U5843 (N_5843,N_1839,N_4938);
nor U5844 (N_5844,N_2991,N_4573);
nor U5845 (N_5845,N_2145,N_448);
or U5846 (N_5846,N_1639,N_4969);
nor U5847 (N_5847,N_2899,N_2112);
and U5848 (N_5848,N_670,N_616);
or U5849 (N_5849,N_936,N_1612);
nand U5850 (N_5850,N_1779,N_3605);
or U5851 (N_5851,N_3245,N_489);
nor U5852 (N_5852,N_1177,N_1311);
nor U5853 (N_5853,N_1461,N_3025);
nand U5854 (N_5854,N_2457,N_3569);
or U5855 (N_5855,N_2693,N_4831);
nand U5856 (N_5856,N_803,N_4946);
or U5857 (N_5857,N_2747,N_2406);
nor U5858 (N_5858,N_1451,N_3919);
nor U5859 (N_5859,N_4217,N_1874);
or U5860 (N_5860,N_1916,N_3314);
nand U5861 (N_5861,N_3639,N_4377);
and U5862 (N_5862,N_1924,N_2967);
or U5863 (N_5863,N_3657,N_1811);
and U5864 (N_5864,N_4415,N_0);
and U5865 (N_5865,N_2065,N_4880);
and U5866 (N_5866,N_2138,N_791);
and U5867 (N_5867,N_1407,N_2487);
nor U5868 (N_5868,N_4321,N_4020);
and U5869 (N_5869,N_3233,N_2541);
nand U5870 (N_5870,N_2442,N_1321);
or U5871 (N_5871,N_1456,N_2706);
and U5872 (N_5872,N_2840,N_2102);
nor U5873 (N_5873,N_3847,N_4862);
nor U5874 (N_5874,N_1286,N_3234);
or U5875 (N_5875,N_3128,N_882);
nor U5876 (N_5876,N_642,N_412);
and U5877 (N_5877,N_2803,N_4250);
or U5878 (N_5878,N_2281,N_2911);
nor U5879 (N_5879,N_1856,N_1665);
and U5880 (N_5880,N_653,N_1327);
nor U5881 (N_5881,N_2679,N_1122);
and U5882 (N_5882,N_2943,N_2738);
or U5883 (N_5883,N_2087,N_138);
or U5884 (N_5884,N_3059,N_3104);
nand U5885 (N_5885,N_3614,N_2697);
and U5886 (N_5886,N_4208,N_807);
and U5887 (N_5887,N_2862,N_4064);
and U5888 (N_5888,N_4330,N_1592);
nand U5889 (N_5889,N_4640,N_1920);
nand U5890 (N_5890,N_859,N_2049);
or U5891 (N_5891,N_1128,N_3306);
or U5892 (N_5892,N_453,N_4852);
nor U5893 (N_5893,N_389,N_4405);
nand U5894 (N_5894,N_3342,N_4538);
nor U5895 (N_5895,N_3432,N_4074);
nand U5896 (N_5896,N_618,N_3160);
nor U5897 (N_5897,N_3303,N_3597);
and U5898 (N_5898,N_4557,N_1071);
nor U5899 (N_5899,N_1126,N_3182);
nor U5900 (N_5900,N_2012,N_3363);
nor U5901 (N_5901,N_1899,N_2052);
and U5902 (N_5902,N_2153,N_4803);
nand U5903 (N_5903,N_2077,N_3274);
nor U5904 (N_5904,N_117,N_1629);
or U5905 (N_5905,N_90,N_4422);
nand U5906 (N_5906,N_2769,N_3550);
and U5907 (N_5907,N_619,N_1469);
nand U5908 (N_5908,N_4789,N_1473);
nor U5909 (N_5909,N_4956,N_1802);
nand U5910 (N_5910,N_1673,N_2485);
and U5911 (N_5911,N_3578,N_4601);
or U5912 (N_5912,N_2563,N_3946);
nor U5913 (N_5913,N_2605,N_3486);
nand U5914 (N_5914,N_636,N_574);
or U5915 (N_5915,N_491,N_4511);
and U5916 (N_5916,N_1031,N_3970);
and U5917 (N_5917,N_357,N_4630);
nor U5918 (N_5918,N_4741,N_1067);
or U5919 (N_5919,N_4580,N_2029);
and U5920 (N_5920,N_1531,N_2253);
or U5921 (N_5921,N_4781,N_36);
and U5922 (N_5922,N_1845,N_2054);
nand U5923 (N_5923,N_1584,N_3433);
or U5924 (N_5924,N_3718,N_1256);
nand U5925 (N_5925,N_2233,N_4896);
nor U5926 (N_5926,N_2834,N_2413);
and U5927 (N_5927,N_4552,N_1626);
nor U5928 (N_5928,N_3949,N_1103);
nor U5929 (N_5929,N_3698,N_565);
or U5930 (N_5930,N_4122,N_4077);
nand U5931 (N_5931,N_2772,N_1229);
or U5932 (N_5932,N_2374,N_1254);
or U5933 (N_5933,N_4382,N_2824);
or U5934 (N_5934,N_3810,N_1301);
and U5935 (N_5935,N_3058,N_3018);
and U5936 (N_5936,N_2241,N_1968);
nor U5937 (N_5937,N_1688,N_4103);
or U5938 (N_5938,N_4331,N_1619);
nand U5939 (N_5939,N_2579,N_2865);
nand U5940 (N_5940,N_1969,N_180);
and U5941 (N_5941,N_3876,N_1773);
and U5942 (N_5942,N_1233,N_4520);
or U5943 (N_5943,N_3130,N_1240);
nor U5944 (N_5944,N_3360,N_4841);
or U5945 (N_5945,N_3304,N_320);
and U5946 (N_5946,N_3246,N_4742);
nand U5947 (N_5947,N_3256,N_57);
nand U5948 (N_5948,N_4230,N_2170);
nor U5949 (N_5949,N_278,N_3864);
and U5950 (N_5950,N_3240,N_2076);
nor U5951 (N_5951,N_999,N_4165);
nor U5952 (N_5952,N_257,N_2371);
nand U5953 (N_5953,N_1799,N_3452);
or U5954 (N_5954,N_963,N_4241);
or U5955 (N_5955,N_391,N_2369);
nand U5956 (N_5956,N_3937,N_4889);
nand U5957 (N_5957,N_2314,N_606);
nand U5958 (N_5958,N_4746,N_1352);
or U5959 (N_5959,N_4009,N_41);
nand U5960 (N_5960,N_2057,N_1202);
or U5961 (N_5961,N_4903,N_3284);
nand U5962 (N_5962,N_2785,N_4772);
or U5963 (N_5963,N_4795,N_118);
nand U5964 (N_5964,N_2458,N_3512);
or U5965 (N_5965,N_3713,N_3888);
or U5966 (N_5966,N_4082,N_4291);
or U5967 (N_5967,N_3514,N_1852);
or U5968 (N_5968,N_2916,N_3199);
nand U5969 (N_5969,N_2328,N_72);
nor U5970 (N_5970,N_4523,N_4642);
and U5971 (N_5971,N_2937,N_4176);
or U5972 (N_5972,N_1355,N_1082);
and U5973 (N_5973,N_997,N_1380);
and U5974 (N_5974,N_602,N_22);
and U5975 (N_5975,N_781,N_1769);
or U5976 (N_5976,N_528,N_3998);
and U5977 (N_5977,N_2750,N_2492);
or U5978 (N_5978,N_146,N_4631);
nor U5979 (N_5979,N_4947,N_4940);
or U5980 (N_5980,N_2776,N_2000);
nor U5981 (N_5981,N_3035,N_3759);
and U5982 (N_5982,N_1360,N_4383);
or U5983 (N_5983,N_4264,N_4468);
or U5984 (N_5984,N_2110,N_2511);
nor U5985 (N_5985,N_18,N_671);
nand U5986 (N_5986,N_1455,N_4317);
or U5987 (N_5987,N_2340,N_3430);
nor U5988 (N_5988,N_390,N_4752);
nand U5989 (N_5989,N_4322,N_3145);
nor U5990 (N_5990,N_3826,N_418);
nor U5991 (N_5991,N_646,N_4808);
and U5992 (N_5992,N_1803,N_3216);
nor U5993 (N_5993,N_2672,N_3416);
nand U5994 (N_5994,N_556,N_4374);
and U5995 (N_5995,N_1120,N_995);
nand U5996 (N_5996,N_1498,N_2470);
nor U5997 (N_5997,N_2298,N_867);
nand U5998 (N_5998,N_4288,N_2332);
nand U5999 (N_5999,N_2572,N_2128);
and U6000 (N_6000,N_3125,N_1724);
nor U6001 (N_6001,N_1742,N_1045);
and U6002 (N_6002,N_1817,N_519);
and U6003 (N_6003,N_1007,N_3703);
and U6004 (N_6004,N_4965,N_3849);
nand U6005 (N_6005,N_1664,N_4005);
or U6006 (N_6006,N_2161,N_3375);
nor U6007 (N_6007,N_1967,N_4211);
or U6008 (N_6008,N_4438,N_2245);
nor U6009 (N_6009,N_2263,N_1759);
nor U6010 (N_6010,N_4863,N_3002);
and U6011 (N_6011,N_2312,N_1242);
nor U6012 (N_6012,N_722,N_1438);
nor U6013 (N_6013,N_569,N_2956);
or U6014 (N_6014,N_1095,N_2044);
nand U6015 (N_6015,N_4655,N_2724);
and U6016 (N_6016,N_1881,N_1628);
and U6017 (N_6017,N_4478,N_1131);
nor U6018 (N_6018,N_1923,N_1962);
nor U6019 (N_6019,N_2816,N_1927);
and U6020 (N_6020,N_3506,N_4323);
nor U6021 (N_6021,N_4167,N_1086);
or U6022 (N_6022,N_3945,N_4086);
nor U6023 (N_6023,N_1383,N_2606);
nand U6024 (N_6024,N_1782,N_2914);
nand U6025 (N_6025,N_1561,N_4691);
nand U6026 (N_6026,N_2817,N_3316);
nor U6027 (N_6027,N_2022,N_3627);
and U6028 (N_6028,N_1184,N_4228);
nor U6029 (N_6029,N_4757,N_4813);
or U6030 (N_6030,N_1587,N_169);
nor U6031 (N_6031,N_1998,N_735);
nor U6032 (N_6032,N_988,N_571);
or U6033 (N_6033,N_2269,N_2673);
nor U6034 (N_6034,N_4102,N_2800);
and U6035 (N_6035,N_922,N_3060);
nor U6036 (N_6036,N_1583,N_4492);
nor U6037 (N_6037,N_1625,N_2981);
and U6038 (N_6038,N_2846,N_233);
nand U6039 (N_6039,N_2348,N_3273);
or U6040 (N_6040,N_342,N_2926);
nand U6041 (N_6041,N_2952,N_1744);
nand U6042 (N_6042,N_1528,N_3255);
and U6043 (N_6043,N_3011,N_1951);
or U6044 (N_6044,N_2581,N_2013);
nor U6045 (N_6045,N_4350,N_4936);
nor U6046 (N_6046,N_2150,N_1953);
and U6047 (N_6047,N_426,N_3279);
or U6048 (N_6048,N_481,N_3765);
and U6049 (N_6049,N_1346,N_3519);
nor U6050 (N_6050,N_4893,N_4702);
nor U6051 (N_6051,N_2443,N_3038);
nor U6052 (N_6052,N_2124,N_4641);
nand U6053 (N_6053,N_2368,N_1351);
nor U6054 (N_6054,N_1876,N_1093);
nand U6055 (N_6055,N_558,N_211);
nand U6056 (N_6056,N_4598,N_3076);
or U6057 (N_6057,N_4216,N_290);
or U6058 (N_6058,N_4907,N_1730);
nand U6059 (N_6059,N_3845,N_4625);
nand U6060 (N_6060,N_4041,N_863);
nand U6061 (N_6061,N_149,N_2882);
and U6062 (N_6062,N_215,N_2710);
nor U6063 (N_6063,N_1402,N_940);
and U6064 (N_6064,N_1931,N_3534);
nand U6065 (N_6065,N_3194,N_4943);
nand U6066 (N_6066,N_487,N_227);
or U6067 (N_6067,N_4287,N_804);
nor U6068 (N_6068,N_2185,N_3193);
or U6069 (N_6069,N_515,N_3911);
or U6070 (N_6070,N_833,N_4870);
nand U6071 (N_6071,N_4644,N_4483);
or U6072 (N_6072,N_2771,N_213);
nor U6073 (N_6073,N_1072,N_3347);
nand U6074 (N_6074,N_4773,N_185);
nor U6075 (N_6075,N_2520,N_1132);
nand U6076 (N_6076,N_4376,N_4780);
nand U6077 (N_6077,N_1678,N_110);
or U6078 (N_6078,N_355,N_838);
or U6079 (N_6079,N_3056,N_3185);
nand U6080 (N_6080,N_4708,N_1363);
nand U6081 (N_6081,N_4594,N_3140);
nor U6082 (N_6082,N_3418,N_1480);
nand U6083 (N_6083,N_1544,N_2179);
nand U6084 (N_6084,N_4622,N_1512);
nand U6085 (N_6085,N_723,N_4504);
xnor U6086 (N_6086,N_1322,N_3154);
and U6087 (N_6087,N_617,N_346);
nor U6088 (N_6088,N_1878,N_393);
and U6089 (N_6089,N_3792,N_2546);
nand U6090 (N_6090,N_476,N_402);
nand U6091 (N_6091,N_4974,N_2753);
and U6092 (N_6092,N_1598,N_1812);
nand U6093 (N_6093,N_2202,N_3031);
nand U6094 (N_6094,N_3126,N_2480);
and U6095 (N_6095,N_1057,N_1537);
nor U6096 (N_6096,N_1439,N_4806);
nor U6097 (N_6097,N_1676,N_1792);
nand U6098 (N_6098,N_4441,N_3954);
and U6099 (N_6099,N_4507,N_3790);
and U6100 (N_6100,N_4001,N_3241);
and U6101 (N_6101,N_4760,N_2896);
and U6102 (N_6102,N_747,N_247);
nand U6103 (N_6103,N_3751,N_1758);
nand U6104 (N_6104,N_4843,N_2583);
nand U6105 (N_6105,N_2201,N_1922);
and U6106 (N_6106,N_1713,N_2285);
and U6107 (N_6107,N_2962,N_2653);
nand U6108 (N_6108,N_105,N_1382);
and U6109 (N_6109,N_1693,N_4237);
or U6110 (N_6110,N_1627,N_2980);
or U6111 (N_6111,N_4698,N_4729);
or U6112 (N_6112,N_2628,N_3899);
and U6113 (N_6113,N_4088,N_310);
nand U6114 (N_6114,N_3215,N_1581);
or U6115 (N_6115,N_582,N_1087);
nand U6116 (N_6116,N_2493,N_3753);
and U6117 (N_6117,N_3743,N_1863);
or U6118 (N_6118,N_4067,N_3827);
or U6119 (N_6119,N_1707,N_2247);
and U6120 (N_6120,N_4171,N_1674);
nor U6121 (N_6121,N_848,N_2313);
nor U6122 (N_6122,N_1405,N_2178);
nand U6123 (N_6123,N_1983,N_4932);
nor U6124 (N_6124,N_3906,N_279);
xor U6125 (N_6125,N_1631,N_4197);
nor U6126 (N_6126,N_298,N_3214);
nand U6127 (N_6127,N_1991,N_2949);
and U6128 (N_6128,N_1026,N_4688);
and U6129 (N_6129,N_4168,N_2219);
or U6130 (N_6130,N_4575,N_3846);
or U6131 (N_6131,N_2678,N_1541);
or U6132 (N_6132,N_142,N_2799);
nor U6133 (N_6133,N_1002,N_2);
nand U6134 (N_6134,N_4156,N_2778);
or U6135 (N_6135,N_2881,N_3034);
nor U6136 (N_6136,N_1829,N_3172);
or U6137 (N_6137,N_209,N_4915);
nand U6138 (N_6138,N_4613,N_4357);
nand U6139 (N_6139,N_3029,N_1467);
nand U6140 (N_6140,N_2149,N_4510);
or U6141 (N_6141,N_2382,N_2496);
or U6142 (N_6142,N_4633,N_984);
or U6143 (N_6143,N_3069,N_43);
nand U6144 (N_6144,N_3707,N_4137);
nand U6145 (N_6145,N_2696,N_1391);
nor U6146 (N_6146,N_1906,N_1047);
or U6147 (N_6147,N_3111,N_4608);
or U6148 (N_6148,N_3456,N_2575);
nor U6149 (N_6149,N_4365,N_2411);
and U6150 (N_6150,N_4296,N_4807);
or U6151 (N_6151,N_750,N_4140);
nand U6152 (N_6152,N_2101,N_472);
or U6153 (N_6153,N_4734,N_3576);
nor U6154 (N_6154,N_4162,N_4989);
nand U6155 (N_6155,N_4452,N_4366);
nand U6156 (N_6156,N_564,N_4456);
nor U6157 (N_6157,N_4447,N_1543);
nand U6158 (N_6158,N_609,N_2905);
nand U6159 (N_6159,N_2199,N_1880);
nand U6160 (N_6160,N_2091,N_1160);
nand U6161 (N_6161,N_1828,N_4387);
nor U6162 (N_6162,N_993,N_2791);
nand U6163 (N_6163,N_3612,N_1134);
nor U6164 (N_6164,N_2652,N_2639);
and U6165 (N_6165,N_1634,N_2250);
nand U6166 (N_6166,N_3667,N_2754);
nand U6167 (N_6167,N_3391,N_2633);
nor U6168 (N_6168,N_1409,N_3878);
and U6169 (N_6169,N_3321,N_4090);
and U6170 (N_6170,N_3,N_761);
nand U6171 (N_6171,N_297,N_1154);
nand U6172 (N_6172,N_2879,N_1593);
and U6173 (N_6173,N_4248,N_3680);
nor U6174 (N_6174,N_3371,N_965);
xnor U6175 (N_6175,N_4793,N_3833);
nand U6176 (N_6176,N_3917,N_3249);
nand U6177 (N_6177,N_495,N_4970);
or U6178 (N_6178,N_4121,N_1374);
nor U6179 (N_6179,N_2388,N_2622);
or U6180 (N_6180,N_411,N_4786);
nand U6181 (N_6181,N_3263,N_1116);
nand U6182 (N_6182,N_758,N_2659);
and U6183 (N_6183,N_2200,N_891);
nand U6184 (N_6184,N_2780,N_2206);
nor U6185 (N_6185,N_2568,N_2509);
or U6186 (N_6186,N_3604,N_3642);
nor U6187 (N_6187,N_1517,N_1142);
nand U6188 (N_6188,N_4471,N_2666);
and U6189 (N_6189,N_605,N_3880);
and U6190 (N_6190,N_4900,N_1576);
and U6191 (N_6191,N_1111,N_3855);
nor U6192 (N_6192,N_109,N_2018);
nor U6193 (N_6193,N_2829,N_1879);
and U6194 (N_6194,N_4138,N_3649);
or U6195 (N_6195,N_4260,N_3623);
nand U6196 (N_6196,N_405,N_4609);
and U6197 (N_6197,N_2254,N_905);
nor U6198 (N_6198,N_4099,N_3712);
nor U6199 (N_6199,N_1791,N_6);
and U6200 (N_6200,N_523,N_2823);
or U6201 (N_6201,N_4030,N_2045);
nand U6202 (N_6202,N_2654,N_3258);
and U6203 (N_6203,N_2004,N_1445);
nor U6204 (N_6204,N_622,N_380);
nand U6205 (N_6205,N_700,N_3400);
nor U6206 (N_6206,N_1666,N_3250);
or U6207 (N_6207,N_666,N_1064);
and U6208 (N_6208,N_289,N_1917);
nand U6209 (N_6209,N_468,N_4577);
or U6210 (N_6210,N_3893,N_4850);
xor U6211 (N_6211,N_1609,N_1014);
or U6212 (N_6212,N_2103,N_2337);
nand U6213 (N_6213,N_4993,N_2394);
and U6214 (N_6214,N_1524,N_1279);
and U6215 (N_6215,N_1375,N_3293);
nor U6216 (N_6216,N_4393,N_2051);
nor U6217 (N_6217,N_1972,N_2901);
and U6218 (N_6218,N_1291,N_4717);
nand U6219 (N_6219,N_3957,N_3853);
or U6220 (N_6220,N_1396,N_4130);
or U6221 (N_6221,N_2167,N_3134);
and U6222 (N_6222,N_1230,N_2125);
nand U6223 (N_6223,N_374,N_1946);
nand U6224 (N_6224,N_3521,N_1258);
and U6225 (N_6225,N_1357,N_3907);
or U6226 (N_6226,N_3841,N_1712);
or U6227 (N_6227,N_766,N_1054);
or U6228 (N_6228,N_2609,N_2972);
nand U6229 (N_6229,N_1055,N_2540);
and U6230 (N_6230,N_8,N_4703);
and U6231 (N_6231,N_3496,N_400);
xor U6232 (N_6232,N_3163,N_2106);
or U6233 (N_6233,N_2037,N_2839);
or U6234 (N_6234,N_413,N_1312);
or U6235 (N_6235,N_3085,N_2483);
or U6236 (N_6236,N_154,N_2434);
or U6237 (N_6237,N_4583,N_1251);
nor U6238 (N_6238,N_4191,N_3121);
or U6239 (N_6239,N_4369,N_3001);
and U6240 (N_6240,N_794,N_3080);
and U6241 (N_6241,N_1124,N_112);
nand U6242 (N_6242,N_4386,N_3213);
or U6243 (N_6243,N_2646,N_2987);
and U6244 (N_6244,N_3476,N_1400);
and U6245 (N_6245,N_1589,N_1212);
nand U6246 (N_6246,N_2321,N_1425);
nand U6247 (N_6247,N_1006,N_786);
nand U6248 (N_6248,N_868,N_2694);
nand U6249 (N_6249,N_503,N_1847);
nand U6250 (N_6250,N_4823,N_1435);
and U6251 (N_6251,N_1056,N_3601);
nand U6252 (N_6252,N_4359,N_194);
or U6253 (N_6253,N_3811,N_34);
nor U6254 (N_6254,N_115,N_690);
and U6255 (N_6255,N_4849,N_3041);
and U6256 (N_6256,N_1168,N_3761);
nor U6257 (N_6257,N_749,N_151);
or U6258 (N_6258,N_3882,N_799);
nor U6259 (N_6259,N_4571,N_2108);
and U6260 (N_6260,N_3281,N_1671);
or U6261 (N_6261,N_1249,N_2884);
or U6262 (N_6262,N_4035,N_3500);
nor U6263 (N_6263,N_1214,N_1877);
nand U6264 (N_6264,N_3681,N_601);
nor U6265 (N_6265,N_3842,N_996);
or U6266 (N_6266,N_4522,N_1024);
nand U6267 (N_6267,N_1422,N_879);
nand U6268 (N_6268,N_159,N_1035);
or U6269 (N_6269,N_3402,N_3294);
nand U6270 (N_6270,N_309,N_4921);
nand U6271 (N_6271,N_3871,N_3549);
or U6272 (N_6272,N_3010,N_3607);
or U6273 (N_6273,N_1336,N_4810);
xnor U6274 (N_6274,N_4431,N_4163);
or U6275 (N_6275,N_133,N_966);
or U6276 (N_6276,N_2993,N_768);
nand U6277 (N_6277,N_3863,N_3850);
or U6278 (N_6278,N_3764,N_3343);
or U6279 (N_6279,N_1472,N_302);
or U6280 (N_6280,N_4572,N_1329);
nor U6281 (N_6281,N_2886,N_4172);
or U6282 (N_6282,N_3982,N_4669);
nor U6283 (N_6283,N_4926,N_1616);
or U6284 (N_6284,N_4055,N_1579);
nand U6285 (N_6285,N_3763,N_3102);
or U6286 (N_6286,N_1450,N_1918);
xnor U6287 (N_6287,N_832,N_449);
and U6288 (N_6288,N_3112,N_3931);
and U6289 (N_6289,N_4332,N_4120);
nand U6290 (N_6290,N_4867,N_4304);
nand U6291 (N_6291,N_970,N_1547);
nand U6292 (N_6292,N_451,N_2113);
nor U6293 (N_6293,N_4647,N_429);
and U6294 (N_6294,N_2082,N_466);
nor U6295 (N_6295,N_4590,N_3700);
or U6296 (N_6296,N_200,N_4524);
or U6297 (N_6297,N_4860,N_3962);
nor U6298 (N_6298,N_785,N_4886);
or U6299 (N_6299,N_2936,N_4599);
and U6300 (N_6300,N_3181,N_1787);
and U6301 (N_6301,N_473,N_514);
nor U6302 (N_6302,N_1272,N_2190);
nor U6303 (N_6303,N_1617,N_2695);
nor U6304 (N_6304,N_344,N_4253);
nand U6305 (N_6305,N_1854,N_3443);
nor U6306 (N_6306,N_2550,N_2909);
nand U6307 (N_6307,N_2786,N_4939);
and U6308 (N_6308,N_3807,N_2203);
and U6309 (N_6309,N_4189,N_1147);
and U6310 (N_6310,N_2822,N_4978);
and U6311 (N_6311,N_3558,N_1995);
or U6312 (N_6312,N_4307,N_1133);
and U6313 (N_6313,N_2454,N_626);
nor U6314 (N_6314,N_1178,N_4426);
or U6315 (N_6315,N_392,N_1424);
nand U6316 (N_6316,N_2019,N_1215);
and U6317 (N_6317,N_238,N_3287);
or U6318 (N_6318,N_2464,N_3320);
nand U6319 (N_6319,N_3617,N_2756);
nor U6320 (N_6320,N_3118,N_3955);
nor U6321 (N_6321,N_4134,N_30);
or U6322 (N_6322,N_522,N_1050);
nand U6323 (N_6323,N_953,N_709);
or U6324 (N_6324,N_3242,N_195);
or U6325 (N_6325,N_2828,N_3419);
or U6326 (N_6326,N_2709,N_74);
nor U6327 (N_6327,N_1813,N_125);
nor U6328 (N_6328,N_4263,N_4512);
and U6329 (N_6329,N_4170,N_906);
and U6330 (N_6330,N_4654,N_731);
and U6331 (N_6331,N_4984,N_4935);
or U6332 (N_6332,N_3030,N_431);
and U6333 (N_6333,N_1221,N_3175);
nand U6334 (N_6334,N_1855,N_1960);
and U6335 (N_6335,N_2308,N_61);
or U6336 (N_6336,N_52,N_1709);
nand U6337 (N_6337,N_1980,N_4298);
nand U6338 (N_6338,N_1790,N_4966);
nand U6339 (N_6339,N_1944,N_4025);
and U6340 (N_6340,N_695,N_2320);
and U6341 (N_6341,N_3247,N_4445);
nor U6342 (N_6342,N_323,N_3985);
or U6343 (N_6343,N_285,N_551);
nand U6344 (N_6344,N_2244,N_2558);
nor U6345 (N_6345,N_4457,N_4066);
nor U6346 (N_6346,N_3687,N_2737);
nor U6347 (N_6347,N_680,N_370);
nand U6348 (N_6348,N_1316,N_757);
and U6349 (N_6349,N_3144,N_2346);
nor U6350 (N_6350,N_3583,N_4453);
nand U6351 (N_6351,N_2225,N_4747);
nor U6352 (N_6352,N_1052,N_4796);
or U6353 (N_6353,N_3626,N_201);
nor U6354 (N_6354,N_789,N_3479);
nand U6355 (N_6355,N_1171,N_4662);
or U6356 (N_6356,N_3071,N_892);
or U6357 (N_6357,N_3501,N_4110);
or U6358 (N_6358,N_1746,N_2565);
or U6359 (N_6359,N_4299,N_1459);
nor U6360 (N_6360,N_332,N_2845);
or U6361 (N_6361,N_1468,N_2721);
or U6362 (N_6362,N_3020,N_1511);
nand U6363 (N_6363,N_3043,N_2792);
nand U6364 (N_6364,N_559,N_1894);
or U6365 (N_6365,N_694,N_2324);
nand U6366 (N_6366,N_732,N_4971);
nand U6367 (N_6367,N_4127,N_900);
nand U6368 (N_6368,N_4914,N_3808);
and U6369 (N_6369,N_896,N_1913);
or U6370 (N_6370,N_2120,N_4578);
nand U6371 (N_6371,N_4261,N_4805);
or U6372 (N_6372,N_2618,N_3089);
nand U6373 (N_6373,N_4398,N_4825);
nand U6374 (N_6374,N_2917,N_756);
and U6375 (N_6375,N_2047,N_2482);
or U6376 (N_6376,N_1532,N_103);
nor U6377 (N_6377,N_1738,N_856);
or U6378 (N_6378,N_2561,N_3575);
and U6379 (N_6379,N_4689,N_2545);
xnor U6380 (N_6380,N_3224,N_3350);
nor U6381 (N_6381,N_305,N_3504);
nor U6382 (N_6382,N_678,N_273);
nand U6383 (N_6383,N_1902,N_3210);
or U6384 (N_6384,N_2402,N_4318);
nor U6385 (N_6385,N_3008,N_492);
nand U6386 (N_6386,N_1265,N_634);
and U6387 (N_6387,N_4462,N_2079);
or U6388 (N_6388,N_1756,N_4558);
nand U6389 (N_6389,N_3042,N_2912);
nor U6390 (N_6390,N_3814,N_4224);
nor U6391 (N_6391,N_2335,N_594);
nand U6392 (N_6392,N_2764,N_3171);
nand U6393 (N_6393,N_164,N_3254);
and U6394 (N_6394,N_2702,N_4908);
or U6395 (N_6395,N_1491,N_2351);
and U6396 (N_6396,N_2954,N_1465);
nand U6397 (N_6397,N_4753,N_2270);
nor U6398 (N_6398,N_4380,N_3131);
or U6399 (N_6399,N_2341,N_3077);
and U6400 (N_6400,N_2992,N_760);
nor U6401 (N_6401,N_1690,N_3036);
nand U6402 (N_6402,N_1016,N_3892);
nor U6403 (N_6403,N_3615,N_253);
nor U6404 (N_6404,N_4402,N_191);
nand U6405 (N_6405,N_3292,N_318);
or U6406 (N_6406,N_2867,N_1476);
or U6407 (N_6407,N_2925,N_4057);
nor U6408 (N_6408,N_4311,N_1834);
and U6409 (N_6409,N_4160,N_1870);
and U6410 (N_6410,N_2667,N_2687);
nand U6411 (N_6411,N_4589,N_1728);
nor U6412 (N_6412,N_1,N_4336);
and U6413 (N_6413,N_2122,N_3553);
and U6414 (N_6414,N_2358,N_3317);
and U6415 (N_6415,N_4039,N_974);
and U6416 (N_6416,N_4036,N_4767);
or U6417 (N_6417,N_3799,N_2096);
and U6418 (N_6418,N_2268,N_1032);
and U6419 (N_6419,N_553,N_795);
nor U6420 (N_6420,N_2015,N_1236);
nor U6421 (N_6421,N_1603,N_1041);
and U6422 (N_6422,N_762,N_3913);
nor U6423 (N_6423,N_2588,N_68);
and U6424 (N_6424,N_3526,N_4252);
and U6425 (N_6425,N_3438,N_2543);
nor U6426 (N_6426,N_912,N_2740);
or U6427 (N_6427,N_282,N_1426);
and U6428 (N_6428,N_4280,N_3195);
and U6429 (N_6429,N_3730,N_1789);
nand U6430 (N_6430,N_3105,N_2671);
or U6431 (N_6431,N_554,N_433);
and U6432 (N_6432,N_1464,N_3736);
or U6433 (N_6433,N_3520,N_2950);
nand U6434 (N_6434,N_2484,N_1421);
and U6435 (N_6435,N_1412,N_1076);
and U6436 (N_6436,N_3620,N_913);
nor U6437 (N_6437,N_1179,N_4650);
nor U6438 (N_6438,N_4275,N_2762);
or U6439 (N_6439,N_1167,N_3770);
xnor U6440 (N_6440,N_463,N_1620);
nand U6441 (N_6441,N_4544,N_3640);
nor U6442 (N_6442,N_4548,N_2513);
nor U6443 (N_6443,N_2183,N_696);
nor U6444 (N_6444,N_4202,N_2969);
or U6445 (N_6445,N_1615,N_3395);
and U6446 (N_6446,N_1466,N_2397);
nor U6447 (N_6447,N_3045,N_3478);
nand U6448 (N_6448,N_3269,N_3748);
nor U6449 (N_6449,N_4023,N_583);
or U6450 (N_6450,N_4847,N_2918);
nand U6451 (N_6451,N_2891,N_3633);
nor U6452 (N_6452,N_4735,N_4555);
and U6453 (N_6453,N_2410,N_1273);
and U6454 (N_6454,N_1843,N_926);
and U6455 (N_6455,N_4273,N_2662);
and U6456 (N_6456,N_877,N_2876);
or U6457 (N_6457,N_3426,N_2255);
or U6458 (N_6458,N_3599,N_3721);
xor U6459 (N_6459,N_359,N_4506);
and U6460 (N_6460,N_4329,N_800);
nand U6461 (N_6461,N_1764,N_3348);
nor U6462 (N_6462,N_1910,N_4668);
and U6463 (N_6463,N_3702,N_471);
or U6464 (N_6464,N_2100,N_4765);
nor U6465 (N_6465,N_113,N_3694);
nand U6466 (N_6466,N_1510,N_1809);
or U6467 (N_6467,N_2364,N_3065);
and U6468 (N_6468,N_3379,N_1797);
nor U6469 (N_6469,N_927,N_4653);
nand U6470 (N_6470,N_2500,N_3183);
and U6471 (N_6471,N_3786,N_2535);
and U6472 (N_6472,N_1798,N_4368);
or U6473 (N_6473,N_3019,N_4108);
nor U6474 (N_6474,N_1264,N_2260);
or U6475 (N_6475,N_4987,N_2173);
or U6476 (N_6476,N_160,N_2033);
or U6477 (N_6477,N_2139,N_3189);
or U6478 (N_6478,N_4541,N_3752);
or U6479 (N_6479,N_2135,N_1862);
nand U6480 (N_6480,N_3533,N_3582);
nor U6481 (N_6481,N_4916,N_1621);
or U6482 (N_6482,N_1390,N_4920);
nor U6483 (N_6483,N_4878,N_3330);
nand U6484 (N_6484,N_239,N_189);
nor U6485 (N_6485,N_1146,N_1105);
nor U6486 (N_6486,N_4300,N_745);
and U6487 (N_6487,N_4229,N_929);
or U6488 (N_6488,N_2433,N_4470);
nand U6489 (N_6489,N_182,N_1175);
or U6490 (N_6490,N_4584,N_71);
or U6491 (N_6491,N_3137,N_4667);
nand U6492 (N_6492,N_2620,N_2474);
and U6493 (N_6493,N_4890,N_4785);
and U6494 (N_6494,N_603,N_144);
and U6495 (N_6495,N_3000,N_2921);
nor U6496 (N_6496,N_4139,N_1198);
nand U6497 (N_6497,N_2133,N_4855);
nor U6498 (N_6498,N_933,N_1320);
nand U6499 (N_6499,N_3096,N_3106);
or U6500 (N_6500,N_4195,N_2532);
or U6501 (N_6501,N_4754,N_983);
nor U6502 (N_6502,N_590,N_3747);
nand U6503 (N_6503,N_513,N_427);
nand U6504 (N_6504,N_4611,N_1837);
and U6505 (N_6505,N_4463,N_3648);
nand U6506 (N_6506,N_2391,N_3635);
nand U6507 (N_6507,N_1471,N_444);
nor U6508 (N_6508,N_1404,N_262);
and U6509 (N_6509,N_2218,N_3768);
and U6510 (N_6510,N_2072,N_1715);
nand U6511 (N_6511,N_2553,N_2890);
and U6512 (N_6512,N_3852,N_3113);
or U6513 (N_6513,N_1979,N_3202);
or U6514 (N_6514,N_2529,N_3843);
and U6515 (N_6515,N_2143,N_2083);
xor U6516 (N_6516,N_2023,N_3107);
nand U6517 (N_6517,N_778,N_3397);
and U6518 (N_6518,N_301,N_3465);
nor U6519 (N_6519,N_477,N_4129);
nor U6520 (N_6520,N_2354,N_2892);
nor U6521 (N_6521,N_1643,N_518);
nor U6522 (N_6522,N_908,N_593);
nand U6523 (N_6523,N_1030,N_4529);
or U6524 (N_6524,N_2903,N_3356);
nand U6525 (N_6525,N_288,N_534);
or U6526 (N_6526,N_2274,N_783);
and U6527 (N_6527,N_2123,N_1340);
nor U6528 (N_6528,N_2258,N_4149);
nor U6529 (N_6529,N_3938,N_2436);
nor U6530 (N_6530,N_3155,N_1763);
nand U6531 (N_6531,N_2288,N_4681);
and U6532 (N_6532,N_2221,N_4337);
and U6533 (N_6533,N_361,N_739);
nand U6534 (N_6534,N_4363,N_1266);
xnor U6535 (N_6535,N_2585,N_4150);
nor U6536 (N_6536,N_4303,N_2979);
and U6537 (N_6537,N_3057,N_3711);
and U6538 (N_6538,N_4142,N_2758);
nor U6539 (N_6539,N_2242,N_1048);
nor U6540 (N_6540,N_2352,N_1938);
nor U6541 (N_6541,N_2420,N_3110);
and U6542 (N_6542,N_203,N_1670);
nand U6543 (N_6543,N_1555,N_4546);
nand U6544 (N_6544,N_2944,N_925);
nand U6545 (N_6545,N_2282,N_3563);
nand U6546 (N_6546,N_3039,N_4954);
nand U6547 (N_6547,N_825,N_1331);
nand U6548 (N_6548,N_3552,N_1554);
and U6549 (N_6549,N_1718,N_2063);
and U6550 (N_6550,N_188,N_1033);
nor U6551 (N_6551,N_3243,N_1161);
or U6552 (N_6552,N_2438,N_4636);
and U6553 (N_6553,N_2401,N_3205);
and U6554 (N_6554,N_4677,N_4861);
nand U6555 (N_6555,N_3048,N_2014);
or U6556 (N_6556,N_935,N_3336);
and U6557 (N_6557,N_4254,N_1685);
nor U6558 (N_6558,N_277,N_4674);
nand U6559 (N_6559,N_252,N_1110);
nand U6560 (N_6560,N_3932,N_3190);
and U6561 (N_6561,N_4794,N_2765);
and U6562 (N_6562,N_1520,N_3206);
nand U6563 (N_6563,N_3883,N_1192);
or U6564 (N_6564,N_1772,N_1395);
or U6565 (N_6565,N_509,N_1127);
nor U6566 (N_6566,N_2810,N_566);
nand U6567 (N_6567,N_70,N_4238);
or U6568 (N_6568,N_266,N_917);
nand U6569 (N_6569,N_3079,N_2475);
or U6570 (N_6570,N_3610,N_1970);
or U6571 (N_6571,N_3230,N_2006);
nand U6572 (N_6572,N_1094,N_496);
nor U6573 (N_6573,N_3380,N_1401);
and U6574 (N_6574,N_1200,N_3063);
nor U6575 (N_6575,N_3941,N_4242);
nand U6576 (N_6576,N_1893,N_2516);
nor U6577 (N_6577,N_3054,N_46);
nor U6578 (N_6578,N_3414,N_4519);
nor U6579 (N_6579,N_3377,N_2768);
nand U6580 (N_6580,N_1935,N_3641);
and U6581 (N_6581,N_1486,N_1368);
nand U6582 (N_6582,N_4615,N_784);
nor U6583 (N_6583,N_497,N_2821);
nor U6584 (N_6584,N_4778,N_885);
nor U6585 (N_6585,N_2836,N_3769);
and U6586 (N_6586,N_3064,N_1419);
and U6587 (N_6587,N_3373,N_1454);
nand U6588 (N_6588,N_2613,N_2789);
and U6589 (N_6589,N_3609,N_1347);
nor U6590 (N_6590,N_1163,N_1118);
and U6591 (N_6591,N_3668,N_2489);
nand U6592 (N_6592,N_1636,N_1073);
or U6593 (N_6593,N_4588,N_313);
nand U6594 (N_6594,N_77,N_1900);
or U6595 (N_6595,N_4661,N_549);
nor U6596 (N_6596,N_4225,N_3473);
or U6597 (N_6597,N_3153,N_2966);
nor U6598 (N_6598,N_2300,N_2717);
or U6599 (N_6599,N_1492,N_73);
nand U6600 (N_6600,N_3516,N_3016);
nand U6601 (N_6601,N_3688,N_1015);
and U6602 (N_6602,N_960,N_537);
and U6603 (N_6603,N_2623,N_1475);
nand U6604 (N_6604,N_644,N_3103);
or U6605 (N_6605,N_2227,N_713);
nor U6606 (N_6606,N_2323,N_312);
nand U6607 (N_6607,N_1757,N_3389);
nand U6608 (N_6608,N_3967,N_4048);
nand U6609 (N_6609,N_982,N_2719);
and U6610 (N_6610,N_1760,N_1800);
nand U6611 (N_6611,N_4425,N_3201);
nand U6612 (N_6612,N_4501,N_2889);
nand U6613 (N_6613,N_2559,N_4340);
nand U6614 (N_6614,N_430,N_4003);
nand U6615 (N_6615,N_4961,N_1997);
nand U6616 (N_6616,N_3200,N_40);
or U6617 (N_6617,N_1741,N_715);
nand U6618 (N_6618,N_665,N_1155);
or U6619 (N_6619,N_272,N_1203);
or U6620 (N_6620,N_2188,N_1121);
and U6621 (N_6621,N_4196,N_2069);
or U6622 (N_6622,N_4885,N_3311);
and U6623 (N_6623,N_2570,N_4866);
nand U6624 (N_6624,N_345,N_2939);
or U6625 (N_6625,N_365,N_2467);
or U6626 (N_6626,N_1632,N_4879);
nand U6627 (N_6627,N_4174,N_1745);
nand U6628 (N_6628,N_942,N_3887);
nor U6629 (N_6629,N_1408,N_4923);
nand U6630 (N_6630,N_3197,N_1936);
and U6631 (N_6631,N_4423,N_946);
nor U6632 (N_6632,N_3602,N_878);
nor U6633 (N_6633,N_2287,N_3138);
nor U6634 (N_6634,N_2632,N_980);
nor U6635 (N_6635,N_3939,N_2366);
or U6636 (N_6636,N_2440,N_3819);
xor U6637 (N_6637,N_1416,N_1182);
nor U6638 (N_6638,N_2748,N_2160);
nand U6639 (N_6639,N_158,N_3793);
xnor U6640 (N_6640,N_1348,N_4151);
nand U6641 (N_6641,N_3381,N_1717);
nand U6642 (N_6642,N_2827,N_4135);
nand U6643 (N_6643,N_2377,N_3291);
nor U6644 (N_6644,N_3896,N_464);
or U6645 (N_6645,N_4319,N_3235);
nand U6646 (N_6646,N_44,N_4593);
or U6647 (N_6647,N_4488,N_3921);
nand U6648 (N_6648,N_1901,N_1253);
or U6649 (N_6649,N_746,N_4992);
nand U6650 (N_6650,N_486,N_3503);
nor U6651 (N_6651,N_4265,N_3801);
and U6652 (N_6652,N_4591,N_3918);
nor U6653 (N_6653,N_904,N_2963);
and U6654 (N_6654,N_629,N_3004);
or U6655 (N_6655,N_2193,N_919);
nand U6656 (N_6656,N_1479,N_3150);
or U6657 (N_6657,N_3666,N_1349);
and U6658 (N_6658,N_2165,N_3522);
nand U6659 (N_6659,N_1075,N_1317);
and U6660 (N_6660,N_1183,N_1958);
nand U6661 (N_6661,N_4430,N_1441);
or U6662 (N_6662,N_3451,N_82);
or U6663 (N_6663,N_4439,N_2104);
and U6664 (N_6664,N_4604,N_3337);
or U6665 (N_6665,N_1807,N_1224);
nor U6666 (N_6666,N_1710,N_1003);
nor U6667 (N_6667,N_2760,N_4844);
or U6668 (N_6668,N_1359,N_4713);
or U6669 (N_6669,N_4065,N_2617);
nand U6670 (N_6670,N_971,N_4532);
and U6671 (N_6671,N_4607,N_2874);
nand U6672 (N_6672,N_162,N_3365);
nor U6673 (N_6673,N_1194,N_3629);
or U6674 (N_6674,N_336,N_1088);
or U6675 (N_6675,N_1851,N_1452);
nor U6676 (N_6676,N_3141,N_1130);
and U6677 (N_6677,N_114,N_240);
nor U6678 (N_6678,N_445,N_42);
nor U6679 (N_6679,N_1714,N_2048);
and U6680 (N_6680,N_2774,N_2322);
nor U6681 (N_6681,N_656,N_2290);
nand U6682 (N_6682,N_1582,N_3546);
and U6683 (N_6683,N_3757,N_4490);
nor U6684 (N_6684,N_3078,N_4226);
and U6685 (N_6685,N_4379,N_3499);
nor U6686 (N_6686,N_1211,N_2809);
xor U6687 (N_6687,N_3951,N_3297);
or U6688 (N_6688,N_488,N_1197);
nand U6689 (N_6689,N_275,N_3094);
nand U6690 (N_6690,N_4568,N_376);
nor U6691 (N_6691,N_505,N_1053);
nor U6692 (N_6692,N_504,N_3874);
and U6693 (N_6693,N_2107,N_1774);
nand U6694 (N_6694,N_316,N_510);
nor U6695 (N_6695,N_3537,N_2665);
and U6696 (N_6696,N_1754,N_3357);
nor U6697 (N_6697,N_4697,N_589);
and U6698 (N_6698,N_1941,N_3518);
nand U6699 (N_6699,N_4569,N_4373);
nor U6700 (N_6700,N_3007,N_2205);
nand U6701 (N_6701,N_2187,N_4804);
and U6702 (N_6702,N_597,N_802);
and U6703 (N_6703,N_1176,N_4183);
and U6704 (N_6704,N_1226,N_1303);
nor U6705 (N_6705,N_1930,N_2355);
and U6706 (N_6706,N_2705,N_1447);
nand U6707 (N_6707,N_2214,N_1896);
nand U6708 (N_6708,N_3536,N_2396);
nand U6709 (N_6709,N_202,N_3239);
nor U6710 (N_6710,N_4175,N_975);
and U6711 (N_6711,N_4081,N_1341);
nand U6712 (N_6712,N_3037,N_2469);
or U6713 (N_6713,N_3948,N_3308);
or U6714 (N_6714,N_2028,N_2256);
nand U6715 (N_6715,N_3310,N_373);
or U6716 (N_6716,N_172,N_1235);
or U6717 (N_6717,N_3326,N_3697);
and U6718 (N_6718,N_55,N_4107);
and U6719 (N_6719,N_2152,N_4812);
and U6720 (N_6720,N_4761,N_1604);
and U6721 (N_6721,N_2924,N_4247);
and U6722 (N_6722,N_1037,N_89);
nor U6723 (N_6723,N_120,N_4411);
nand U6724 (N_6724,N_2009,N_2988);
or U6725 (N_6725,N_2983,N_2291);
or U6726 (N_6726,N_2363,N_2703);
nor U6727 (N_6727,N_1482,N_4327);
nor U6728 (N_6728,N_4811,N_79);
and U6729 (N_6729,N_3875,N_793);
and U6730 (N_6730,N_2419,N_167);
nand U6731 (N_6731,N_4295,N_4161);
nor U6732 (N_6732,N_1940,N_2506);
nand U6733 (N_6733,N_4872,N_1477);
or U6734 (N_6734,N_2409,N_625);
nor U6735 (N_6735,N_3742,N_3457);
nor U6736 (N_6736,N_3881,N_1074);
nand U6737 (N_6737,N_1417,N_94);
nor U6738 (N_6738,N_4147,N_64);
and U6739 (N_6739,N_4454,N_333);
or U6740 (N_6740,N_2236,N_3963);
nor U6741 (N_6741,N_699,N_2272);
or U6742 (N_6742,N_2299,N_858);
and U6743 (N_6743,N_1646,N_1644);
nand U6744 (N_6744,N_881,N_4648);
or U6745 (N_6745,N_181,N_2249);
nand U6746 (N_6746,N_1929,N_4887);
nor U6747 (N_6747,N_2264,N_3434);
nor U6748 (N_6748,N_2589,N_943);
nor U6749 (N_6749,N_4559,N_1684);
nor U6750 (N_6750,N_4141,N_1394);
and U6751 (N_6751,N_1677,N_1500);
nand U6752 (N_6752,N_2497,N_3969);
and U6753 (N_6753,N_2189,N_1138);
nand U6754 (N_6754,N_3714,N_4283);
or U6755 (N_6755,N_4128,N_1339);
nor U6756 (N_6756,N_718,N_3288);
nand U6757 (N_6757,N_2598,N_3528);
nand U6758 (N_6758,N_870,N_4840);
or U6759 (N_6759,N_1385,N_2275);
or U6760 (N_6760,N_3588,N_27);
nand U6761 (N_6761,N_2325,N_2265);
or U6762 (N_6762,N_4968,N_4762);
nor U6763 (N_6763,N_226,N_540);
or U6764 (N_6764,N_4909,N_1274);
nand U6765 (N_6765,N_4547,N_3046);
nand U6766 (N_6766,N_577,N_4059);
or U6767 (N_6767,N_3726,N_1150);
nand U6768 (N_6768,N_244,N_2712);
nand U6769 (N_6769,N_2790,N_1752);
xnor U6770 (N_6770,N_4394,N_2460);
nand U6771 (N_6771,N_1384,N_2421);
or U6772 (N_6772,N_11,N_2343);
and U6773 (N_6773,N_4829,N_772);
or U6774 (N_6774,N_2379,N_2166);
or U6775 (N_6775,N_4737,N_798);
nor U6776 (N_6776,N_4286,N_248);
nand U6777 (N_6777,N_1125,N_3366);
or U6778 (N_6778,N_375,N_2669);
nor U6779 (N_6779,N_3228,N_2908);
nand U6780 (N_6780,N_3979,N_1025);
nor U6781 (N_6781,N_4392,N_1296);
nor U6782 (N_6782,N_1943,N_3209);
nor U6783 (N_6783,N_1084,N_1699);
nor U6784 (N_6784,N_1070,N_3143);
nor U6785 (N_6785,N_1478,N_4100);
nand U6786 (N_6786,N_1398,N_4182);
nand U6787 (N_6787,N_4898,N_4706);
or U6788 (N_6788,N_675,N_1158);
nand U6789 (N_6789,N_584,N_1350);
or U6790 (N_6790,N_3403,N_1882);
or U6791 (N_6791,N_3296,N_934);
or U6792 (N_6792,N_2574,N_641);
or U6793 (N_6793,N_930,N_3159);
and U6794 (N_6794,N_2851,N_2861);
nand U6795 (N_6795,N_4945,N_2461);
or U6796 (N_6796,N_1551,N_4227);
nor U6797 (N_6797,N_4692,N_83);
nor U6798 (N_6798,N_1850,N_2347);
nand U6799 (N_6799,N_2081,N_1503);
or U6800 (N_6800,N_3052,N_2508);
and U6801 (N_6801,N_458,N_3409);
nor U6802 (N_6802,N_4489,N_3413);
nor U6803 (N_6803,N_3510,N_1356);
or U6804 (N_6804,N_4282,N_3660);
or U6805 (N_6805,N_2510,N_1819);
and U6806 (N_6806,N_334,N_1444);
and U6807 (N_6807,N_759,N_1397);
and U6808 (N_6808,N_3328,N_1804);
and U6809 (N_6809,N_3332,N_475);
or U6810 (N_6810,N_3832,N_2897);
xnor U6811 (N_6811,N_3839,N_587);
nor U6812 (N_6812,N_4846,N_3992);
nand U6813 (N_6813,N_2777,N_4930);
and U6814 (N_6814,N_127,N_2562);
nand U6815 (N_6815,N_2142,N_1937);
or U6816 (N_6816,N_1504,N_4390);
nor U6817 (N_6817,N_1739,N_2336);
or U6818 (N_6818,N_314,N_3541);
and U6819 (N_6819,N_2555,N_4751);
nor U6820 (N_6820,N_3387,N_2906);
or U6821 (N_6821,N_207,N_773);
and U6822 (N_6822,N_3417,N_2691);
nand U6823 (N_6823,N_2757,N_890);
nor U6824 (N_6824,N_2431,N_2134);
and U6825 (N_6825,N_4994,N_968);
nor U6826 (N_6826,N_3441,N_3302);
nand U6827 (N_6827,N_4084,N_3772);
and U6828 (N_6828,N_2739,N_1366);
and U6829 (N_6829,N_60,N_4711);
nand U6830 (N_6830,N_790,N_4868);
nor U6831 (N_6831,N_343,N_1565);
and U6832 (N_6832,N_325,N_4848);
or U6833 (N_6833,N_2271,N_1869);
or U6834 (N_6834,N_1600,N_3828);
or U6835 (N_6835,N_2519,N_3867);
or U6836 (N_6836,N_84,N_4651);
nand U6837 (N_6837,N_1228,N_640);
or U6838 (N_6838,N_1319,N_2061);
nand U6839 (N_6839,N_3672,N_2728);
nand U6840 (N_6840,N_177,N_561);
nand U6841 (N_6841,N_371,N_2111);
and U6842 (N_6842,N_1952,N_2648);
or U6843 (N_6843,N_2989,N_659);
nor U6844 (N_6844,N_4201,N_1548);
xnor U6845 (N_6845,N_1696,N_1663);
nor U6846 (N_6846,N_2389,N_2370);
and U6847 (N_6847,N_797,N_884);
or U6848 (N_6848,N_1928,N_4678);
nand U6849 (N_6849,N_4998,N_421);
nor U6850 (N_6850,N_480,N_4755);
nand U6851 (N_6851,N_4166,N_1017);
and U6852 (N_6852,N_4895,N_1232);
nor U6853 (N_6853,N_1806,N_4278);
and U6854 (N_6854,N_2405,N_3861);
nand U6855 (N_6855,N_4649,N_2465);
nor U6856 (N_6856,N_4089,N_1668);
nor U6857 (N_6857,N_3777,N_1721);
and U6858 (N_6858,N_673,N_219);
and U6859 (N_6859,N_1605,N_3675);
nand U6860 (N_6860,N_957,N_1988);
nand U6861 (N_6861,N_3719,N_719);
xnor U6862 (N_6862,N_3323,N_501);
and U6863 (N_6863,N_1691,N_937);
or U6864 (N_6864,N_3531,N_1727);
nand U6865 (N_6865,N_2614,N_3741);
or U6866 (N_6866,N_4696,N_1058);
nor U6867 (N_6867,N_2393,N_482);
nand U6868 (N_6868,N_3074,N_474);
or U6869 (N_6869,N_830,N_455);
nand U6870 (N_6870,N_3662,N_575);
nor U6871 (N_6871,N_2755,N_3062);
nand U6872 (N_6872,N_2025,N_3050);
and U6873 (N_6873,N_1020,N_4853);
nor U6874 (N_6874,N_1716,N_4078);
nand U6875 (N_6875,N_2450,N_643);
xor U6876 (N_6876,N_1244,N_3491);
nand U6877 (N_6877,N_1680,N_4117);
nand U6878 (N_6878,N_3227,N_3341);
or U6879 (N_6879,N_462,N_4770);
nor U6880 (N_6880,N_2171,N_4232);
nand U6881 (N_6881,N_3910,N_1559);
or U6882 (N_6882,N_4389,N_632);
nor U6883 (N_6883,N_4986,N_2441);
nor U6884 (N_6884,N_410,N_4450);
nand U6885 (N_6885,N_2232,N_129);
nand U6886 (N_6886,N_3865,N_4787);
nand U6887 (N_6887,N_80,N_2262);
nand U6888 (N_6888,N_952,N_1546);
nor U6889 (N_6889,N_3820,N_2521);
nand U6890 (N_6890,N_3547,N_3346);
nor U6891 (N_6891,N_631,N_1449);
nor U6892 (N_6892,N_3760,N_4509);
nor U6893 (N_6893,N_1078,N_3737);
and U6894 (N_6894,N_4220,N_4054);
or U6895 (N_6895,N_4505,N_1682);
and U6896 (N_6896,N_1027,N_1821);
and U6897 (N_6897,N_857,N_2027);
xnor U6898 (N_6898,N_1783,N_2345);
or U6899 (N_6899,N_1898,N_2380);
nand U6900 (N_6900,N_1586,N_4612);
or U6901 (N_6901,N_1269,N_4316);
and U6902 (N_6902,N_2931,N_2965);
nand U6903 (N_6903,N_2852,N_3226);
nor U6904 (N_6904,N_806,N_2446);
nand U6905 (N_6905,N_1765,N_4022);
nand U6906 (N_6906,N_2126,N_3840);
and U6907 (N_6907,N_2554,N_1100);
nand U6908 (N_6908,N_1305,N_2499);
and U6909 (N_6909,N_3082,N_3565);
nor U6910 (N_6910,N_538,N_3908);
and U6911 (N_6911,N_3487,N_1832);
or U6912 (N_6912,N_4219,N_4010);
nand U6913 (N_6913,N_4045,N_3359);
nand U6914 (N_6914,N_4919,N_2215);
and U6915 (N_6915,N_2858,N_705);
nor U6916 (N_6916,N_4764,N_4234);
or U6917 (N_6917,N_53,N_4750);
nand U6918 (N_6918,N_3665,N_961);
nor U6919 (N_6919,N_2001,N_2885);
and U6920 (N_6920,N_2131,N_414);
and U6921 (N_6921,N_3448,N_2038);
nand U6922 (N_6922,N_4414,N_4815);
nor U6923 (N_6923,N_2599,N_4257);
nand U6924 (N_6924,N_2742,N_2523);
or U6925 (N_6925,N_315,N_4312);
and U6926 (N_6926,N_303,N_837);
or U6927 (N_6927,N_2182,N_3237);
and U6928 (N_6928,N_349,N_3886);
or U6929 (N_6929,N_274,N_1818);
or U6930 (N_6930,N_869,N_1655);
nor U6931 (N_6931,N_119,N_1597);
nand U6932 (N_6932,N_3715,N_3156);
or U6933 (N_6933,N_1706,N_2478);
or U6934 (N_6934,N_3275,N_4576);
or U6935 (N_6935,N_2661,N_2399);
and U6936 (N_6936,N_3142,N_1129);
or U6937 (N_6937,N_4477,N_2990);
or U6938 (N_6938,N_1814,N_190);
or U6939 (N_6939,N_2946,N_2490);
nand U6940 (N_6940,N_66,N_4721);
and U6941 (N_6941,N_3600,N_979);
nor U6942 (N_6942,N_536,N_1300);
or U6943 (N_6943,N_1066,N_923);
and U6944 (N_6944,N_4744,N_419);
nand U6945 (N_6945,N_1822,N_2294);
nand U6946 (N_6946,N_1575,N_4877);
nand U6947 (N_6947,N_484,N_1853);
and U6948 (N_6948,N_2976,N_3169);
nor U6949 (N_6949,N_4536,N_2277);
nand U6950 (N_6950,N_1225,N_271);
nor U6951 (N_6951,N_3831,N_3746);
or U6952 (N_6952,N_3309,N_1302);
and U6953 (N_6953,N_4941,N_4912);
nor U6954 (N_6954,N_3055,N_465);
and U6955 (N_6955,N_2228,N_3868);
and U6956 (N_6956,N_918,N_2212);
and U6957 (N_6957,N_2922,N_363);
nor U6958 (N_6958,N_541,N_1702);
or U6959 (N_6959,N_356,N_340);
nand U6960 (N_6960,N_817,N_3236);
nor U6961 (N_6961,N_4775,N_1387);
nand U6962 (N_6962,N_533,N_1761);
nor U6963 (N_6963,N_1732,N_4051);
and U6964 (N_6964,N_220,N_4614);
and U6965 (N_6965,N_3787,N_1501);
and U6966 (N_6966,N_2920,N_175);
or U6967 (N_6967,N_4579,N_294);
nand U6968 (N_6968,N_805,N_1308);
or U6969 (N_6969,N_2448,N_4864);
nand U6970 (N_6970,N_1989,N_4587);
and U6971 (N_6971,N_3322,N_4610);
nand U6972 (N_6972,N_2592,N_3976);
and U6973 (N_6973,N_3208,N_4526);
and U6974 (N_6974,N_2727,N_3987);
or U6975 (N_6975,N_1112,N_308);
nor U6976 (N_6976,N_1373,N_4101);
or U6977 (N_6977,N_4883,N_3280);
nand U6978 (N_6978,N_4097,N_1376);
and U6979 (N_6979,N_1186,N_3988);
and U6980 (N_6980,N_2684,N_1323);
or U6981 (N_6981,N_2008,N_1207);
nor U6982 (N_6982,N_96,N_726);
nand U6983 (N_6983,N_909,N_4707);
nor U6984 (N_6984,N_3897,N_2248);
nor U6985 (N_6985,N_4123,N_3984);
and U6986 (N_6986,N_4656,N_4029);
nor U6987 (N_6987,N_2713,N_2745);
nor U6988 (N_6988,N_3929,N_1227);
nand U6989 (N_6989,N_3968,N_131);
nand U6990 (N_6990,N_3157,N_3953);
xnor U6991 (N_6991,N_1099,N_28);
nand U6992 (N_6992,N_1622,N_3505);
or U6993 (N_6993,N_4586,N_178);
and U6994 (N_6994,N_3723,N_4957);
and U6995 (N_6995,N_1040,N_3994);
and U6996 (N_6996,N_3785,N_4052);
and U6997 (N_6997,N_2144,N_134);
nor U6998 (N_6998,N_669,N_3511);
and U6999 (N_6999,N_4525,N_3950);
or U7000 (N_7000,N_1957,N_2224);
or U7001 (N_7001,N_2502,N_3061);
nor U7002 (N_7002,N_3983,N_26);
or U7003 (N_7003,N_4313,N_4629);
and U7004 (N_7004,N_368,N_755);
nor U7005 (N_7005,N_4199,N_3158);
and U7006 (N_7006,N_459,N_2435);
nor U7007 (N_7007,N_2833,N_3313);
nand U7008 (N_7008,N_2226,N_525);
nand U7009 (N_7009,N_4564,N_1353);
nor U7010 (N_7010,N_3900,N_4620);
nand U7011 (N_7011,N_4824,N_2597);
or U7012 (N_7012,N_3710,N_2196);
nor U7013 (N_7013,N_2872,N_1560);
or U7014 (N_7014,N_1414,N_4428);
nor U7015 (N_7015,N_388,N_888);
nand U7016 (N_7016,N_531,N_2690);
nand U7017 (N_7017,N_330,N_1181);
and U7018 (N_7018,N_733,N_4344);
nand U7019 (N_7019,N_2237,N_3699);
and U7020 (N_7020,N_2349,N_580);
or U7021 (N_7021,N_3916,N_3270);
nor U7022 (N_7022,N_49,N_221);
nor U7023 (N_7023,N_3689,N_1849);
nand U7024 (N_7024,N_4749,N_1737);
and U7025 (N_7025,N_4155,N_1539);
or U7026 (N_7026,N_1000,N_608);
or U7027 (N_7027,N_3947,N_2158);
and U7028 (N_7028,N_3358,N_3716);
nor U7029 (N_7029,N_153,N_2698);
or U7030 (N_7030,N_1871,N_3312);
and U7031 (N_7031,N_1781,N_2156);
nor U7032 (N_7032,N_241,N_4269);
and U7033 (N_7033,N_4809,N_3873);
nand U7034 (N_7034,N_3362,N_259);
nand U7035 (N_7035,N_2010,N_216);
nand U7036 (N_7036,N_4833,N_620);
nand U7037 (N_7037,N_3188,N_1692);
nand U7038 (N_7038,N_2842,N_12);
nor U7039 (N_7039,N_372,N_4996);
nor U7040 (N_7040,N_4333,N_3406);
and U7041 (N_7041,N_4042,N_921);
nor U7042 (N_7042,N_3540,N_439);
nor U7043 (N_7043,N_2856,N_1794);
and U7044 (N_7044,N_287,N_2180);
or U7045 (N_7045,N_3423,N_3805);
or U7046 (N_7046,N_1652,N_1262);
and U7047 (N_7047,N_4455,N_1328);
nor U7048 (N_7048,N_4169,N_4646);
or U7049 (N_7049,N_4297,N_2670);
and U7050 (N_7050,N_3364,N_847);
or U7051 (N_7051,N_4771,N_4485);
and U7052 (N_7052,N_3944,N_1954);
or U7053 (N_7053,N_4187,N_4343);
nor U7054 (N_7054,N_1297,N_2286);
nor U7055 (N_7055,N_2707,N_2318);
nor U7056 (N_7056,N_4543,N_2522);
nor U7057 (N_7057,N_928,N_1601);
nand U7058 (N_7058,N_311,N_1298);
nand U7059 (N_7059,N_3124,N_1553);
or U7060 (N_7060,N_4212,N_1755);
nor U7061 (N_7061,N_1885,N_2229);
nand U7062 (N_7062,N_2688,N_3788);
and U7063 (N_7063,N_2176,N_4157);
nand U7064 (N_7064,N_3480,N_4985);
or U7065 (N_7065,N_2974,N_3488);
nor U7066 (N_7066,N_4461,N_460);
nor U7067 (N_7067,N_4497,N_4348);
and U7068 (N_7068,N_3616,N_645);
nor U7069 (N_7069,N_1085,N_4884);
xor U7070 (N_7070,N_284,N_2080);
nand U7071 (N_7071,N_4098,N_3898);
nand U7072 (N_7072,N_1443,N_3087);
nor U7073 (N_7073,N_3727,N_2844);
xnor U7074 (N_7074,N_1681,N_3203);
nor U7075 (N_7075,N_147,N_989);
or U7076 (N_7076,N_1018,N_2507);
and U7077 (N_7077,N_3283,N_1399);
and U7078 (N_7078,N_2002,N_3267);
nor U7079 (N_7079,N_1533,N_3740);
and U7080 (N_7080,N_545,N_3554);
nand U7081 (N_7081,N_108,N_165);
nor U7082 (N_7082,N_1518,N_2569);
nand U7083 (N_7083,N_2951,N_818);
and U7084 (N_7084,N_4560,N_3495);
nor U7085 (N_7085,N_4888,N_2408);
nand U7086 (N_7086,N_3859,N_4851);
and U7087 (N_7087,N_520,N_4730);
and U7088 (N_7088,N_3184,N_3005);
nor U7089 (N_7089,N_3463,N_4666);
nand U7090 (N_7090,N_2580,N_2806);
and U7091 (N_7091,N_2900,N_3653);
and U7092 (N_7092,N_4349,N_1495);
or U7093 (N_7093,N_4472,N_1169);
and U7094 (N_7094,N_4070,N_1263);
and U7095 (N_7095,N_2121,N_3630);
xor U7096 (N_7096,N_4738,N_1008);
or U7097 (N_7097,N_920,N_1505);
nor U7098 (N_7098,N_4104,N_4821);
or U7099 (N_7099,N_4186,N_1858);
nor U7100 (N_7100,N_3838,N_950);
nor U7101 (N_7101,N_4660,N_2071);
nor U7102 (N_7102,N_3439,N_3339);
nor U7103 (N_7103,N_1289,N_4047);
nand U7104 (N_7104,N_2174,N_1153);
or U7105 (N_7105,N_1786,N_2660);
nand U7106 (N_7106,N_1640,N_3795);
and U7107 (N_7107,N_3461,N_4424);
nand U7108 (N_7108,N_579,N_3705);
xor U7109 (N_7109,N_3659,N_3532);
nand U7110 (N_7110,N_2517,N_2744);
or U7111 (N_7111,N_2020,N_1335);
or U7112 (N_7112,N_48,N_2430);
or U7113 (N_7113,N_4596,N_1816);
or U7114 (N_7114,N_2273,N_4704);
nor U7115 (N_7115,N_2334,N_717);
nand U7116 (N_7116,N_1978,N_1569);
and U7117 (N_7117,N_3067,N_3225);
and U7118 (N_7118,N_1649,N_1836);
and U7119 (N_7119,N_1342,N_1795);
and U7120 (N_7120,N_1218,N_4293);
nand U7121 (N_7121,N_2439,N_2428);
and U7122 (N_7122,N_2217,N_3956);
nor U7123 (N_7123,N_3090,N_924);
nand U7124 (N_7124,N_1942,N_1719);
or U7125 (N_7125,N_3421,N_1162);
or U7126 (N_7126,N_2140,N_562);
nor U7127 (N_7127,N_2078,N_15);
nand U7128 (N_7128,N_1971,N_664);
or U7129 (N_7129,N_3767,N_4869);
or U7130 (N_7130,N_3545,N_3467);
nand U7131 (N_7131,N_769,N_4911);
or U7132 (N_7132,N_32,N_1393);
or U7133 (N_7133,N_588,N_3484);
nand U7134 (N_7134,N_3165,N_1661);
nor U7135 (N_7135,N_4114,N_255);
or U7136 (N_7136,N_728,N_4972);
or U7137 (N_7137,N_2175,N_3603);
nand U7138 (N_7138,N_1109,N_4341);
nor U7139 (N_7139,N_4592,N_4019);
nand U7140 (N_7140,N_1831,N_4545);
nor U7141 (N_7141,N_3628,N_788);
and U7142 (N_7142,N_834,N_4427);
nor U7143 (N_7143,N_4338,N_250);
nor U7144 (N_7144,N_3643,N_1389);
nor U7145 (N_7145,N_1523,N_852);
and U7146 (N_7146,N_4310,N_217);
nor U7147 (N_7147,N_2686,N_3218);
nor U7148 (N_7148,N_2356,N_3989);
and U7149 (N_7149,N_1019,N_1949);
nand U7150 (N_7150,N_4361,N_4976);
or U7151 (N_7151,N_1519,N_2024);
nand U7152 (N_7152,N_4181,N_1651);
and U7153 (N_7153,N_1137,N_827);
nor U7154 (N_7154,N_223,N_2058);
nand U7155 (N_7155,N_3914,N_1725);
and U7156 (N_7156,N_3724,N_2978);
and U7157 (N_7157,N_1238,N_4566);
and U7158 (N_7158,N_3187,N_327);
or U7159 (N_7159,N_3611,N_787);
nand U7160 (N_7160,N_3564,N_1106);
or U7161 (N_7161,N_2279,N_3207);
nor U7162 (N_7162,N_4305,N_3720);
nand U7163 (N_7163,N_4014,N_328);
or U7164 (N_7164,N_1552,N_4015);
nor U7165 (N_7165,N_2035,N_2629);
nor U7166 (N_7166,N_2295,N_4567);
and U7167 (N_7167,N_2003,N_3958);
and U7168 (N_7168,N_1613,N_3393);
and U7169 (N_7169,N_3482,N_2902);
and U7170 (N_7170,N_4906,N_4929);
nand U7171 (N_7171,N_2455,N_2888);
nor U7172 (N_7172,N_249,N_107);
and U7173 (N_7173,N_1354,N_3555);
or U7174 (N_7174,N_4498,N_3428);
or U7175 (N_7175,N_4207,N_2383);
and U7176 (N_7176,N_1984,N_2542);
nor U7177 (N_7177,N_2526,N_1872);
nor U7178 (N_7178,N_1413,N_214);
nor U7179 (N_7179,N_4491,N_3823);
nor U7180 (N_7180,N_4190,N_1675);
nor U7181 (N_7181,N_3542,N_4910);
nand U7182 (N_7182,N_4158,N_1704);
or U7183 (N_7183,N_2964,N_1695);
nand U7184 (N_7184,N_369,N_576);
xor U7185 (N_7185,N_251,N_1698);
nand U7186 (N_7186,N_3442,N_1536);
or U7187 (N_7187,N_1446,N_2537);
or U7188 (N_7188,N_2129,N_1687);
or U7189 (N_7189,N_2604,N_3369);
nor U7190 (N_7190,N_809,N_572);
nand U7191 (N_7191,N_4240,N_1144);
nor U7192 (N_7192,N_2427,N_2407);
nor U7193 (N_7193,N_776,N_4028);
or U7194 (N_7194,N_2148,N_3264);
nor U7195 (N_7195,N_2689,N_1222);
nand U7196 (N_7196,N_4400,N_3783);
and U7197 (N_7197,N_4664,N_4467);
nand U7198 (N_7198,N_2452,N_4115);
nand U7199 (N_7199,N_3099,N_461);
nand U7200 (N_7200,N_1912,N_2105);
or U7201 (N_7201,N_712,N_4782);
nand U7202 (N_7202,N_1623,N_1306);
and U7203 (N_7203,N_3806,N_403);
or U7204 (N_7204,N_3933,N_3162);
nand U7205 (N_7205,N_2301,N_2869);
nand U7206 (N_7206,N_171,N_2017);
and U7207 (N_7207,N_1474,N_1081);
or U7208 (N_7208,N_4682,N_3836);
or U7209 (N_7209,N_2259,N_1669);
nand U7210 (N_7210,N_3816,N_548);
nor U7211 (N_7211,N_871,N_1820);
or U7212 (N_7212,N_3382,N_3682);
nor U7213 (N_7213,N_3114,N_3266);
or U7214 (N_7214,N_4244,N_4769);
or U7215 (N_7215,N_3912,N_4531);
nand U7216 (N_7216,N_1720,N_2788);
or U7217 (N_7217,N_3965,N_4982);
nor U7218 (N_7218,N_931,N_2895);
or U7219 (N_7219,N_236,N_697);
xnor U7220 (N_7220,N_1864,N_4032);
nand U7221 (N_7221,N_1290,N_765);
or U7222 (N_7222,N_2463,N_16);
nand U7223 (N_7223,N_2392,N_1001);
nand U7224 (N_7224,N_998,N_2734);
and U7225 (N_7225,N_1568,N_1494);
and U7226 (N_7226,N_4928,N_1115);
nand U7227 (N_7227,N_2802,N_2638);
or U7228 (N_7228,N_4838,N_3804);
nor U7229 (N_7229,N_324,N_4581);
nor U7230 (N_7230,N_4085,N_962);
nor U7231 (N_7231,N_1624,N_4499);
nand U7232 (N_7232,N_3632,N_1838);
nor U7233 (N_7233,N_4518,N_730);
nor U7234 (N_7234,N_1280,N_4554);
and U7235 (N_7235,N_4262,N_2942);
nor U7236 (N_7236,N_442,N_2675);
nand U7237 (N_7237,N_35,N_1602);
nor U7238 (N_7238,N_4854,N_1433);
nand U7239 (N_7239,N_1926,N_2995);
or U7240 (N_7240,N_1046,N_4194);
nor U7241 (N_7241,N_2362,N_1022);
or U7242 (N_7242,N_141,N_339);
or U7243 (N_7243,N_1201,N_58);
and U7244 (N_7244,N_1051,N_816);
and U7245 (N_7245,N_4177,N_681);
or U7246 (N_7246,N_4315,N_2787);
and U7247 (N_7247,N_1332,N_385);
nor U7248 (N_7248,N_526,N_3261);
nor U7249 (N_7249,N_1516,N_2501);
and U7250 (N_7250,N_3590,N_4837);
or U7251 (N_7251,N_3277,N_4665);
nor U7252 (N_7252,N_972,N_3993);
or U7253 (N_7253,N_1611,N_1281);
or U7254 (N_7254,N_2164,N_2655);
nor U7255 (N_7255,N_3146,N_3729);
nor U7256 (N_7256,N_3622,N_1102);
nand U7257 (N_7257,N_1762,N_2304);
nand U7258 (N_7258,N_973,N_1428);
nor U7259 (N_7259,N_397,N_4012);
nor U7260 (N_7260,N_547,N_4981);
or U7261 (N_7261,N_3858,N_3877);
or U7262 (N_7262,N_1700,N_3798);
nand U7263 (N_7263,N_2923,N_822);
nand U7264 (N_7264,N_3345,N_2875);
or U7265 (N_7265,N_210,N_4409);
nor U7266 (N_7266,N_3251,N_3073);
and U7267 (N_7267,N_3170,N_1199);
and U7268 (N_7268,N_3398,N_2036);
or U7269 (N_7269,N_63,N_4034);
nor U7270 (N_7270,N_4897,N_677);
or U7271 (N_7271,N_1950,N_50);
nand U7272 (N_7272,N_682,N_614);
nor U7273 (N_7273,N_4960,N_4549);
or U7274 (N_7274,N_1334,N_4768);
and U7275 (N_7275,N_3928,N_152);
nor U7276 (N_7276,N_3361,N_56);
and U7277 (N_7277,N_2878,N_5);
nand U7278 (N_7278,N_4550,N_331);
and U7279 (N_7279,N_1362,N_1403);
nand U7280 (N_7280,N_3834,N_4094);
or U7281 (N_7281,N_3021,N_3775);
and U7282 (N_7282,N_1004,N_4963);
and U7283 (N_7283,N_801,N_69);
nand U7284 (N_7284,N_2676,N_4476);
and U7285 (N_7285,N_2353,N_2958);
or U7286 (N_7286,N_454,N_3708);
and U7287 (N_7287,N_4617,N_3679);
and U7288 (N_7288,N_955,N_782);
nand U7289 (N_7289,N_639,N_121);
nand U7290 (N_7290,N_3527,N_3091);
nor U7291 (N_7291,N_3525,N_4979);
nand U7292 (N_7292,N_3655,N_4459);
nor U7293 (N_7293,N_4865,N_654);
or U7294 (N_7294,N_4528,N_4419);
or U7295 (N_7295,N_3524,N_3285);
nor U7296 (N_7296,N_2053,N_4395);
and U7297 (N_7297,N_2773,N_4213);
or U7298 (N_7298,N_37,N_3494);
or U7299 (N_7299,N_2309,N_1610);
nor U7300 (N_7300,N_752,N_3809);
nand U7301 (N_7301,N_3384,N_3837);
and U7302 (N_7302,N_796,N_2715);
and U7303 (N_7303,N_148,N_3468);
and U7304 (N_7304,N_1502,N_2276);
and U7305 (N_7305,N_4326,N_1276);
nand U7306 (N_7306,N_2663,N_3164);
or U7307 (N_7307,N_4397,N_4977);
nand U7308 (N_7308,N_4743,N_2252);
and U7309 (N_7309,N_1219,N_3386);
and U7310 (N_7310,N_124,N_1934);
nand U7311 (N_7311,N_1933,N_2319);
nor U7312 (N_7312,N_4830,N_901);
nand U7313 (N_7313,N_3731,N_2726);
nand U7314 (N_7314,N_4404,N_3889);
or U7315 (N_7315,N_4367,N_4044);
nand U7316 (N_7316,N_292,N_4901);
nor U7317 (N_7317,N_4236,N_1488);
or U7318 (N_7318,N_2610,N_708);
or U7319 (N_7319,N_1827,N_4553);
or U7320 (N_7320,N_3646,N_4686);
nand U7321 (N_7321,N_4328,N_2637);
nand U7322 (N_7322,N_2736,N_4272);
nor U7323 (N_7323,N_3490,N_2417);
nor U7324 (N_7324,N_2578,N_1701);
and U7325 (N_7325,N_3637,N_502);
nor U7326 (N_7326,N_3454,N_1606);
nor U7327 (N_7327,N_2961,N_1304);
and U7328 (N_7328,N_4214,N_4759);
and U7329 (N_7329,N_3282,N_4111);
nor U7330 (N_7330,N_2505,N_2466);
nand U7331 (N_7331,N_4072,N_3744);
nand U7332 (N_7332,N_2854,N_507);
or U7333 (N_7333,N_2386,N_862);
nor U7334 (N_7334,N_381,N_1325);
and U7335 (N_7335,N_3354,N_1993);
nor U7336 (N_7336,N_2350,N_4881);
and U7337 (N_7337,N_4637,N_4624);
nor U7338 (N_7338,N_3211,N_4063);
nand U7339 (N_7339,N_4774,N_714);
nand U7340 (N_7340,N_3606,N_3943);
nor U7341 (N_7341,N_2826,N_3636);
and U7342 (N_7342,N_674,N_2615);
nor U7343 (N_7343,N_550,N_3412);
nand U7344 (N_7344,N_2118,N_2280);
or U7345 (N_7345,N_3095,N_2375);
or U7346 (N_7346,N_4516,N_78);
and U7347 (N_7347,N_3331,N_2919);
nand U7348 (N_7348,N_2996,N_1743);
nor U7349 (N_7349,N_4308,N_1556);
and U7350 (N_7350,N_3755,N_2524);
nand U7351 (N_7351,N_87,N_4685);
xnor U7352 (N_7352,N_443,N_546);
nand U7353 (N_7353,N_3272,N_1490);
nor U7354 (N_7354,N_754,N_4585);
nand U7355 (N_7355,N_193,N_2797);
or U7356 (N_7356,N_4413,N_4502);
and U7357 (N_7357,N_621,N_4659);
nor U7358 (N_7358,N_176,N_3446);
and U7359 (N_7359,N_3186,N_1694);
nand U7360 (N_7360,N_4712,N_611);
nor U7361 (N_7361,N_2743,N_1101);
nor U7362 (N_7362,N_1530,N_450);
and U7363 (N_7363,N_3717,N_1293);
and U7364 (N_7364,N_1574,N_823);
nor U7365 (N_7365,N_2476,N_1865);
xor U7366 (N_7366,N_842,N_4635);
or U7367 (N_7367,N_4801,N_543);
nand U7368 (N_7368,N_2929,N_3661);
xnor U7369 (N_7369,N_3370,N_2257);
nand U7370 (N_7370,N_3952,N_1961);
nor U7371 (N_7371,N_4570,N_2934);
or U7372 (N_7372,N_3613,N_2026);
and U7373 (N_7373,N_1932,N_2848);
nand U7374 (N_7374,N_3890,N_4144);
nand U7375 (N_7375,N_1889,N_1771);
nor U7376 (N_7376,N_743,N_1442);
nand U7377 (N_7377,N_2095,N_1736);
and U7378 (N_7378,N_2601,N_1726);
nand U7379 (N_7379,N_1123,N_4192);
nand U7380 (N_7380,N_1261,N_2089);
nand U7381 (N_7381,N_2716,N_1107);
xor U7382 (N_7382,N_3972,N_1595);
nor U7383 (N_7383,N_648,N_2871);
xnor U7384 (N_7384,N_4799,N_2197);
and U7385 (N_7385,N_186,N_4542);
or U7386 (N_7386,N_592,N_3390);
or U7387 (N_7387,N_692,N_2447);
nor U7388 (N_7388,N_4351,N_1540);
nor U7389 (N_7389,N_384,N_944);
nand U7390 (N_7390,N_1873,N_1657);
and U7391 (N_7391,N_3835,N_3013);
nand U7392 (N_7392,N_1440,N_4093);
and U7393 (N_7393,N_2039,N_2154);
and U7394 (N_7394,N_506,N_4416);
or U7395 (N_7395,N_1324,N_494);
and U7396 (N_7396,N_4132,N_2376);
nor U7397 (N_7397,N_4013,N_3268);
nor U7398 (N_7398,N_4922,N_2590);
or U7399 (N_7399,N_4657,N_4816);
and U7400 (N_7400,N_527,N_1775);
and U7401 (N_7401,N_2339,N_4882);
and U7402 (N_7402,N_658,N_2913);
or U7403 (N_7403,N_3497,N_45);
nor U7404 (N_7404,N_668,N_1378);
nor U7405 (N_7405,N_2548,N_4040);
or U7406 (N_7406,N_1982,N_4680);
nor U7407 (N_7407,N_98,N_672);
or U7408 (N_7408,N_4364,N_2381);
or U7409 (N_7409,N_3385,N_2857);
nand U7410 (N_7410,N_598,N_243);
or U7411 (N_7411,N_1039,N_3024);
nand U7412 (N_7412,N_702,N_1987);
nand U7413 (N_7413,N_1977,N_2209);
nor U7414 (N_7414,N_1766,N_2132);
and U7415 (N_7415,N_4835,N_2935);
nand U7416 (N_7416,N_1113,N_1059);
or U7417 (N_7417,N_861,N_1660);
or U7418 (N_7418,N_959,N_3098);
and U7419 (N_7419,N_4913,N_3248);
nor U7420 (N_7420,N_2163,N_2042);
nand U7421 (N_7421,N_4997,N_4200);
nor U7422 (N_7422,N_2831,N_2261);
and U7423 (N_7423,N_4027,N_24);
nor U7424 (N_7424,N_727,N_651);
or U7425 (N_7425,N_4779,N_3523);
or U7426 (N_7426,N_4792,N_4952);
nand U7427 (N_7427,N_3817,N_4687);
and U7428 (N_7428,N_775,N_3191);
and U7429 (N_7429,N_3619,N_1751);
nand U7430 (N_7430,N_1683,N_2928);
nor U7431 (N_7431,N_4959,N_3517);
and U7432 (N_7432,N_123,N_3650);
or U7433 (N_7433,N_1333,N_2873);
nand U7434 (N_7434,N_4995,N_3445);
or U7435 (N_7435,N_3120,N_2251);
or U7436 (N_7436,N_3493,N_1708);
nor U7437 (N_7437,N_4205,N_4652);
or U7438 (N_7438,N_1260,N_3462);
nand U7439 (N_7439,N_4011,N_3551);
and U7440 (N_7440,N_4475,N_895);
nand U7441 (N_7441,N_1973,N_567);
or U7442 (N_7442,N_4820,N_3844);
nand U7443 (N_7443,N_1697,N_667);
nand U7444 (N_7444,N_3420,N_1239);
and U7445 (N_7445,N_3027,N_4784);
nor U7446 (N_7446,N_1415,N_4206);
nand U7447 (N_7447,N_3593,N_615);
nand U7448 (N_7448,N_2151,N_4016);
or U7449 (N_7449,N_3086,N_2481);
nor U7450 (N_7450,N_4991,N_1367);
nand U7451 (N_7451,N_1268,N_4482);
and U7452 (N_7452,N_270,N_394);
or U7453 (N_7453,N_1381,N_2796);
or U7454 (N_7454,N_3513,N_3286);
and U7455 (N_7455,N_2887,N_1956);
and U7456 (N_7456,N_1259,N_542);
nor U7457 (N_7457,N_1729,N_2109);
and U7458 (N_7458,N_150,N_93);
and U7459 (N_7459,N_4618,N_2390);
nand U7460 (N_7460,N_2735,N_2825);
or U7461 (N_7461,N_2429,N_1591);
nor U7462 (N_7462,N_276,N_4434);
xnor U7463 (N_7463,N_398,N_544);
or U7464 (N_7464,N_771,N_353);
or U7465 (N_7465,N_1689,N_4218);
or U7466 (N_7466,N_3652,N_218);
nand U7467 (N_7467,N_3136,N_2527);
nor U7468 (N_7468,N_3677,N_2444);
nor U7469 (N_7469,N_1209,N_3068);
nand U7470 (N_7470,N_2327,N_956);
nor U7471 (N_7471,N_3940,N_3870);
nor U7472 (N_7472,N_229,N_2783);
nand U7473 (N_7473,N_3936,N_2621);
and U7474 (N_7474,N_1489,N_4600);
or U7475 (N_7475,N_139,N_4748);
nor U7476 (N_7476,N_4325,N_1267);
nand U7477 (N_7477,N_2801,N_1010);
and U7478 (N_7478,N_4437,N_604);
nand U7479 (N_7479,N_1947,N_3975);
xnor U7480 (N_7480,N_1420,N_1453);
nor U7481 (N_7481,N_2472,N_2631);
and U7482 (N_7482,N_2400,N_1796);
nor U7483 (N_7483,N_4616,N_1157);
nand U7484 (N_7484,N_4087,N_4918);
and U7485 (N_7485,N_4873,N_1785);
and U7486 (N_7486,N_1005,N_4284);
nand U7487 (N_7487,N_1588,N_3771);
nor U7488 (N_7488,N_2093,N_1392);
nor U7489 (N_7489,N_948,N_4643);
nor U7490 (N_7490,N_2119,N_3431);
nor U7491 (N_7491,N_4403,N_1722);
and U7492 (N_7492,N_197,N_4597);
nor U7493 (N_7493,N_4944,N_3572);
and U7494 (N_7494,N_1667,N_95);
or U7495 (N_7495,N_341,N_3625);
and U7496 (N_7496,N_824,N_1187);
and U7497 (N_7497,N_350,N_3009);
and U7498 (N_7498,N_1166,N_4075);
nand U7499 (N_7499,N_1365,N_4154);
or U7500 (N_7500,N_1170,N_574);
nor U7501 (N_7501,N_601,N_3724);
or U7502 (N_7502,N_4236,N_3007);
nor U7503 (N_7503,N_56,N_4099);
nand U7504 (N_7504,N_3780,N_980);
nand U7505 (N_7505,N_1526,N_1221);
and U7506 (N_7506,N_4536,N_4723);
and U7507 (N_7507,N_4240,N_1773);
nand U7508 (N_7508,N_549,N_4075);
or U7509 (N_7509,N_2514,N_115);
or U7510 (N_7510,N_2290,N_1308);
and U7511 (N_7511,N_2042,N_891);
nand U7512 (N_7512,N_2727,N_3836);
and U7513 (N_7513,N_685,N_2991);
or U7514 (N_7514,N_1904,N_643);
and U7515 (N_7515,N_4066,N_455);
and U7516 (N_7516,N_802,N_751);
or U7517 (N_7517,N_830,N_2573);
and U7518 (N_7518,N_60,N_4494);
and U7519 (N_7519,N_1314,N_2211);
nand U7520 (N_7520,N_641,N_2044);
xnor U7521 (N_7521,N_1142,N_857);
nand U7522 (N_7522,N_4364,N_3416);
or U7523 (N_7523,N_2995,N_2285);
and U7524 (N_7524,N_4498,N_2712);
or U7525 (N_7525,N_2639,N_2965);
nor U7526 (N_7526,N_954,N_3342);
nand U7527 (N_7527,N_4572,N_4530);
nor U7528 (N_7528,N_4542,N_1584);
nand U7529 (N_7529,N_1786,N_1070);
nor U7530 (N_7530,N_3429,N_400);
and U7531 (N_7531,N_1549,N_1318);
or U7532 (N_7532,N_3301,N_1407);
nor U7533 (N_7533,N_2079,N_518);
and U7534 (N_7534,N_1094,N_4789);
nand U7535 (N_7535,N_948,N_472);
and U7536 (N_7536,N_4093,N_2563);
and U7537 (N_7537,N_117,N_1643);
nand U7538 (N_7538,N_4523,N_2852);
nand U7539 (N_7539,N_1405,N_4951);
or U7540 (N_7540,N_487,N_4117);
and U7541 (N_7541,N_4157,N_949);
or U7542 (N_7542,N_592,N_1109);
and U7543 (N_7543,N_1096,N_622);
and U7544 (N_7544,N_2030,N_155);
and U7545 (N_7545,N_267,N_3571);
and U7546 (N_7546,N_533,N_231);
or U7547 (N_7547,N_4702,N_3952);
nor U7548 (N_7548,N_4341,N_3486);
or U7549 (N_7549,N_2190,N_2662);
and U7550 (N_7550,N_2260,N_2351);
nor U7551 (N_7551,N_3548,N_161);
or U7552 (N_7552,N_388,N_3177);
or U7553 (N_7553,N_1228,N_4371);
or U7554 (N_7554,N_910,N_2197);
and U7555 (N_7555,N_4345,N_3568);
or U7556 (N_7556,N_1652,N_4986);
or U7557 (N_7557,N_4426,N_2992);
nor U7558 (N_7558,N_2383,N_4087);
or U7559 (N_7559,N_1640,N_3141);
nor U7560 (N_7560,N_4673,N_2274);
and U7561 (N_7561,N_3037,N_593);
and U7562 (N_7562,N_2422,N_2502);
or U7563 (N_7563,N_2775,N_3781);
nor U7564 (N_7564,N_4009,N_1416);
and U7565 (N_7565,N_4306,N_4050);
nand U7566 (N_7566,N_1852,N_842);
nand U7567 (N_7567,N_3029,N_3022);
or U7568 (N_7568,N_3758,N_1091);
nand U7569 (N_7569,N_2575,N_1858);
nand U7570 (N_7570,N_325,N_2518);
nor U7571 (N_7571,N_290,N_222);
or U7572 (N_7572,N_4067,N_1487);
nor U7573 (N_7573,N_2630,N_3026);
or U7574 (N_7574,N_2000,N_374);
and U7575 (N_7575,N_2513,N_2136);
nand U7576 (N_7576,N_2667,N_2780);
nor U7577 (N_7577,N_2939,N_4387);
nor U7578 (N_7578,N_4546,N_4407);
and U7579 (N_7579,N_71,N_1419);
nand U7580 (N_7580,N_624,N_3213);
or U7581 (N_7581,N_3126,N_197);
and U7582 (N_7582,N_3562,N_1869);
nor U7583 (N_7583,N_3378,N_3529);
nand U7584 (N_7584,N_2909,N_3269);
and U7585 (N_7585,N_4824,N_4420);
or U7586 (N_7586,N_655,N_3123);
nor U7587 (N_7587,N_3299,N_303);
and U7588 (N_7588,N_1956,N_1763);
nor U7589 (N_7589,N_1358,N_4158);
nand U7590 (N_7590,N_4976,N_4198);
nand U7591 (N_7591,N_115,N_29);
nand U7592 (N_7592,N_564,N_959);
and U7593 (N_7593,N_903,N_79);
nand U7594 (N_7594,N_4023,N_3812);
or U7595 (N_7595,N_3620,N_4864);
or U7596 (N_7596,N_1488,N_2343);
nand U7597 (N_7597,N_4535,N_4888);
or U7598 (N_7598,N_2921,N_3247);
nor U7599 (N_7599,N_1873,N_1504);
or U7600 (N_7600,N_4734,N_2428);
nand U7601 (N_7601,N_1852,N_939);
nand U7602 (N_7602,N_4921,N_3063);
and U7603 (N_7603,N_4397,N_3955);
nor U7604 (N_7604,N_2105,N_3594);
or U7605 (N_7605,N_4264,N_3373);
and U7606 (N_7606,N_3003,N_4545);
nor U7607 (N_7607,N_42,N_2754);
nand U7608 (N_7608,N_2030,N_4066);
nand U7609 (N_7609,N_1277,N_1707);
or U7610 (N_7610,N_1108,N_1683);
nand U7611 (N_7611,N_1897,N_1596);
and U7612 (N_7612,N_4268,N_1976);
or U7613 (N_7613,N_3043,N_4057);
and U7614 (N_7614,N_2153,N_2156);
and U7615 (N_7615,N_856,N_3334);
and U7616 (N_7616,N_1596,N_779);
or U7617 (N_7617,N_89,N_1771);
nor U7618 (N_7618,N_3420,N_2082);
nand U7619 (N_7619,N_360,N_4598);
or U7620 (N_7620,N_4441,N_4619);
and U7621 (N_7621,N_3493,N_2744);
nor U7622 (N_7622,N_3751,N_3011);
and U7623 (N_7623,N_2107,N_1112);
nand U7624 (N_7624,N_2571,N_2085);
and U7625 (N_7625,N_3092,N_3281);
nand U7626 (N_7626,N_1530,N_663);
nor U7627 (N_7627,N_4650,N_3072);
and U7628 (N_7628,N_4034,N_4878);
nor U7629 (N_7629,N_4884,N_3289);
and U7630 (N_7630,N_675,N_3341);
nor U7631 (N_7631,N_3930,N_3422);
or U7632 (N_7632,N_2914,N_2313);
nor U7633 (N_7633,N_1675,N_91);
nor U7634 (N_7634,N_1740,N_4050);
or U7635 (N_7635,N_4476,N_4810);
and U7636 (N_7636,N_1481,N_1684);
and U7637 (N_7637,N_3686,N_2336);
nand U7638 (N_7638,N_307,N_3985);
nor U7639 (N_7639,N_1329,N_3608);
and U7640 (N_7640,N_2393,N_2552);
and U7641 (N_7641,N_4190,N_4111);
or U7642 (N_7642,N_2662,N_1474);
or U7643 (N_7643,N_2802,N_4211);
or U7644 (N_7644,N_3110,N_144);
xnor U7645 (N_7645,N_9,N_1966);
and U7646 (N_7646,N_4207,N_741);
nor U7647 (N_7647,N_648,N_1484);
and U7648 (N_7648,N_3443,N_909);
nand U7649 (N_7649,N_3611,N_3001);
nand U7650 (N_7650,N_4687,N_1234);
and U7651 (N_7651,N_4534,N_2798);
nand U7652 (N_7652,N_2581,N_312);
or U7653 (N_7653,N_489,N_4967);
and U7654 (N_7654,N_1458,N_2578);
and U7655 (N_7655,N_3025,N_3511);
or U7656 (N_7656,N_4813,N_4908);
or U7657 (N_7657,N_3915,N_2465);
or U7658 (N_7658,N_3975,N_3230);
nor U7659 (N_7659,N_2247,N_2179);
nand U7660 (N_7660,N_3989,N_4397);
xor U7661 (N_7661,N_2938,N_3281);
nand U7662 (N_7662,N_4488,N_1767);
nor U7663 (N_7663,N_3343,N_4886);
nand U7664 (N_7664,N_469,N_3173);
or U7665 (N_7665,N_4315,N_2941);
or U7666 (N_7666,N_3965,N_267);
and U7667 (N_7667,N_635,N_1317);
nor U7668 (N_7668,N_734,N_2873);
nor U7669 (N_7669,N_3732,N_2344);
nand U7670 (N_7670,N_671,N_1703);
and U7671 (N_7671,N_1154,N_3052);
xor U7672 (N_7672,N_4432,N_4995);
and U7673 (N_7673,N_277,N_732);
and U7674 (N_7674,N_2310,N_3769);
or U7675 (N_7675,N_2908,N_1507);
and U7676 (N_7676,N_4371,N_4859);
nand U7677 (N_7677,N_972,N_4968);
and U7678 (N_7678,N_1215,N_782);
nand U7679 (N_7679,N_3992,N_4679);
and U7680 (N_7680,N_2953,N_4288);
nand U7681 (N_7681,N_3394,N_4586);
nand U7682 (N_7682,N_3234,N_4460);
nor U7683 (N_7683,N_4438,N_2978);
or U7684 (N_7684,N_3926,N_4973);
nor U7685 (N_7685,N_4677,N_3113);
nor U7686 (N_7686,N_254,N_2026);
and U7687 (N_7687,N_3642,N_4561);
and U7688 (N_7688,N_4068,N_2521);
or U7689 (N_7689,N_4879,N_255);
or U7690 (N_7690,N_4640,N_4973);
nor U7691 (N_7691,N_1047,N_270);
and U7692 (N_7692,N_1191,N_3476);
or U7693 (N_7693,N_3607,N_913);
nand U7694 (N_7694,N_4986,N_2169);
nand U7695 (N_7695,N_2680,N_3863);
or U7696 (N_7696,N_1594,N_514);
and U7697 (N_7697,N_4873,N_3709);
nor U7698 (N_7698,N_3617,N_4648);
nand U7699 (N_7699,N_588,N_2620);
nand U7700 (N_7700,N_394,N_938);
and U7701 (N_7701,N_519,N_2651);
nor U7702 (N_7702,N_1666,N_3161);
and U7703 (N_7703,N_2149,N_593);
nor U7704 (N_7704,N_3032,N_3079);
nor U7705 (N_7705,N_2041,N_4199);
or U7706 (N_7706,N_4762,N_774);
and U7707 (N_7707,N_4369,N_4958);
and U7708 (N_7708,N_1871,N_2533);
nand U7709 (N_7709,N_456,N_758);
and U7710 (N_7710,N_1996,N_2963);
nand U7711 (N_7711,N_3848,N_3603);
nand U7712 (N_7712,N_3423,N_1065);
nor U7713 (N_7713,N_3711,N_2029);
nor U7714 (N_7714,N_3115,N_3930);
and U7715 (N_7715,N_583,N_2511);
nand U7716 (N_7716,N_2315,N_3733);
or U7717 (N_7717,N_212,N_1106);
nand U7718 (N_7718,N_2666,N_3783);
or U7719 (N_7719,N_748,N_3536);
and U7720 (N_7720,N_4668,N_3873);
nor U7721 (N_7721,N_4513,N_565);
and U7722 (N_7722,N_1069,N_3624);
nor U7723 (N_7723,N_2195,N_3610);
nand U7724 (N_7724,N_2413,N_2927);
nand U7725 (N_7725,N_4436,N_2956);
nand U7726 (N_7726,N_1473,N_4740);
nor U7727 (N_7727,N_4994,N_649);
nor U7728 (N_7728,N_2019,N_4361);
nand U7729 (N_7729,N_87,N_1409);
xnor U7730 (N_7730,N_3949,N_3831);
nor U7731 (N_7731,N_3574,N_3782);
or U7732 (N_7732,N_2790,N_3971);
nand U7733 (N_7733,N_1523,N_857);
nand U7734 (N_7734,N_343,N_1472);
nor U7735 (N_7735,N_2494,N_1789);
and U7736 (N_7736,N_4406,N_3420);
nor U7737 (N_7737,N_1169,N_1507);
nor U7738 (N_7738,N_1177,N_1116);
or U7739 (N_7739,N_176,N_3224);
nand U7740 (N_7740,N_1884,N_3945);
or U7741 (N_7741,N_683,N_1898);
and U7742 (N_7742,N_885,N_2918);
nand U7743 (N_7743,N_3565,N_1070);
nand U7744 (N_7744,N_3606,N_1145);
or U7745 (N_7745,N_1908,N_1458);
nor U7746 (N_7746,N_583,N_2075);
or U7747 (N_7747,N_3547,N_3549);
nor U7748 (N_7748,N_4945,N_1444);
nand U7749 (N_7749,N_1496,N_4673);
or U7750 (N_7750,N_2851,N_2592);
nand U7751 (N_7751,N_2831,N_4130);
nor U7752 (N_7752,N_3339,N_2948);
nor U7753 (N_7753,N_3178,N_3059);
and U7754 (N_7754,N_3832,N_2553);
nor U7755 (N_7755,N_2106,N_432);
nand U7756 (N_7756,N_3060,N_2861);
or U7757 (N_7757,N_1673,N_4406);
and U7758 (N_7758,N_4184,N_3218);
and U7759 (N_7759,N_987,N_134);
or U7760 (N_7760,N_1692,N_775);
nand U7761 (N_7761,N_1483,N_1827);
or U7762 (N_7762,N_693,N_4722);
and U7763 (N_7763,N_2658,N_718);
and U7764 (N_7764,N_3266,N_325);
nor U7765 (N_7765,N_4574,N_2571);
nor U7766 (N_7766,N_4035,N_346);
or U7767 (N_7767,N_1715,N_3519);
and U7768 (N_7768,N_575,N_4224);
nand U7769 (N_7769,N_83,N_2575);
nand U7770 (N_7770,N_784,N_741);
and U7771 (N_7771,N_1236,N_127);
nand U7772 (N_7772,N_3916,N_2676);
nand U7773 (N_7773,N_4193,N_1330);
nand U7774 (N_7774,N_2421,N_1551);
nand U7775 (N_7775,N_2471,N_2191);
or U7776 (N_7776,N_4064,N_4151);
nand U7777 (N_7777,N_1994,N_602);
nor U7778 (N_7778,N_1741,N_1040);
nor U7779 (N_7779,N_299,N_1853);
or U7780 (N_7780,N_77,N_3282);
or U7781 (N_7781,N_3561,N_973);
or U7782 (N_7782,N_25,N_138);
nand U7783 (N_7783,N_1341,N_2786);
nand U7784 (N_7784,N_3737,N_4647);
or U7785 (N_7785,N_3120,N_298);
nand U7786 (N_7786,N_4660,N_523);
or U7787 (N_7787,N_3912,N_14);
and U7788 (N_7788,N_1949,N_173);
nor U7789 (N_7789,N_1363,N_3528);
or U7790 (N_7790,N_1696,N_4965);
nor U7791 (N_7791,N_2683,N_1142);
nor U7792 (N_7792,N_1838,N_3521);
or U7793 (N_7793,N_3439,N_4911);
nand U7794 (N_7794,N_2301,N_1844);
nand U7795 (N_7795,N_4379,N_4468);
and U7796 (N_7796,N_3658,N_716);
and U7797 (N_7797,N_2956,N_1769);
nor U7798 (N_7798,N_2296,N_3766);
or U7799 (N_7799,N_1580,N_3677);
nor U7800 (N_7800,N_2852,N_1899);
or U7801 (N_7801,N_805,N_971);
nand U7802 (N_7802,N_3976,N_282);
nor U7803 (N_7803,N_3535,N_2659);
nor U7804 (N_7804,N_749,N_4553);
nand U7805 (N_7805,N_2172,N_3448);
nand U7806 (N_7806,N_3983,N_1220);
xnor U7807 (N_7807,N_2386,N_4853);
nand U7808 (N_7808,N_2330,N_2524);
or U7809 (N_7809,N_1021,N_3956);
nand U7810 (N_7810,N_2079,N_3873);
nand U7811 (N_7811,N_2111,N_1630);
nor U7812 (N_7812,N_4326,N_1411);
nor U7813 (N_7813,N_1658,N_537);
or U7814 (N_7814,N_3246,N_848);
nor U7815 (N_7815,N_27,N_3604);
and U7816 (N_7816,N_2724,N_4581);
nor U7817 (N_7817,N_231,N_2818);
nand U7818 (N_7818,N_1788,N_1029);
xor U7819 (N_7819,N_219,N_2847);
nor U7820 (N_7820,N_2473,N_1098);
and U7821 (N_7821,N_780,N_1913);
and U7822 (N_7822,N_1860,N_2181);
and U7823 (N_7823,N_4238,N_3379);
nor U7824 (N_7824,N_1490,N_912);
nor U7825 (N_7825,N_998,N_4218);
or U7826 (N_7826,N_2219,N_434);
nor U7827 (N_7827,N_413,N_2618);
nand U7828 (N_7828,N_4249,N_651);
nor U7829 (N_7829,N_1956,N_2799);
nand U7830 (N_7830,N_3130,N_3128);
or U7831 (N_7831,N_1925,N_3533);
and U7832 (N_7832,N_4526,N_908);
nand U7833 (N_7833,N_3499,N_126);
nand U7834 (N_7834,N_276,N_3924);
nand U7835 (N_7835,N_4805,N_3002);
nor U7836 (N_7836,N_4270,N_2898);
nand U7837 (N_7837,N_3609,N_3888);
and U7838 (N_7838,N_3403,N_2164);
or U7839 (N_7839,N_622,N_4047);
nand U7840 (N_7840,N_1417,N_3468);
or U7841 (N_7841,N_1177,N_225);
nor U7842 (N_7842,N_4671,N_2385);
nand U7843 (N_7843,N_566,N_4303);
and U7844 (N_7844,N_829,N_3438);
nand U7845 (N_7845,N_1649,N_2694);
or U7846 (N_7846,N_552,N_4196);
nand U7847 (N_7847,N_1103,N_3637);
nor U7848 (N_7848,N_447,N_1095);
and U7849 (N_7849,N_4735,N_1061);
and U7850 (N_7850,N_3108,N_1695);
and U7851 (N_7851,N_2247,N_2584);
or U7852 (N_7852,N_170,N_1785);
nand U7853 (N_7853,N_4838,N_236);
nor U7854 (N_7854,N_421,N_21);
nand U7855 (N_7855,N_3622,N_1779);
nor U7856 (N_7856,N_2605,N_1037);
nor U7857 (N_7857,N_108,N_2999);
nor U7858 (N_7858,N_4081,N_3623);
nor U7859 (N_7859,N_1030,N_2483);
or U7860 (N_7860,N_831,N_905);
nor U7861 (N_7861,N_3775,N_231);
and U7862 (N_7862,N_3013,N_3299);
nand U7863 (N_7863,N_4379,N_1512);
or U7864 (N_7864,N_2630,N_4430);
nor U7865 (N_7865,N_1033,N_2241);
and U7866 (N_7866,N_1663,N_3558);
and U7867 (N_7867,N_428,N_4157);
and U7868 (N_7868,N_142,N_1846);
or U7869 (N_7869,N_2758,N_2992);
or U7870 (N_7870,N_2174,N_1461);
nor U7871 (N_7871,N_4376,N_2815);
or U7872 (N_7872,N_4881,N_3054);
nor U7873 (N_7873,N_1196,N_329);
xnor U7874 (N_7874,N_2920,N_4122);
and U7875 (N_7875,N_1633,N_4351);
or U7876 (N_7876,N_1282,N_2965);
nand U7877 (N_7877,N_3166,N_1213);
nand U7878 (N_7878,N_1655,N_1198);
nor U7879 (N_7879,N_4239,N_3414);
nand U7880 (N_7880,N_3985,N_3742);
nand U7881 (N_7881,N_3775,N_4889);
nand U7882 (N_7882,N_2444,N_603);
nand U7883 (N_7883,N_2673,N_2231);
or U7884 (N_7884,N_4644,N_2716);
nor U7885 (N_7885,N_761,N_3013);
nand U7886 (N_7886,N_61,N_96);
or U7887 (N_7887,N_102,N_362);
or U7888 (N_7888,N_3518,N_3007);
nand U7889 (N_7889,N_2846,N_3797);
nand U7890 (N_7890,N_4555,N_1957);
and U7891 (N_7891,N_2041,N_618);
and U7892 (N_7892,N_3708,N_2844);
and U7893 (N_7893,N_4816,N_267);
and U7894 (N_7894,N_4402,N_558);
and U7895 (N_7895,N_1751,N_4488);
nand U7896 (N_7896,N_924,N_2816);
nand U7897 (N_7897,N_4242,N_1859);
or U7898 (N_7898,N_1991,N_394);
and U7899 (N_7899,N_420,N_1104);
or U7900 (N_7900,N_4400,N_1832);
nor U7901 (N_7901,N_1930,N_3555);
nor U7902 (N_7902,N_1429,N_1140);
and U7903 (N_7903,N_3307,N_861);
and U7904 (N_7904,N_595,N_1133);
or U7905 (N_7905,N_4387,N_4786);
nand U7906 (N_7906,N_981,N_1256);
nor U7907 (N_7907,N_303,N_2157);
nor U7908 (N_7908,N_944,N_3809);
nor U7909 (N_7909,N_564,N_2221);
and U7910 (N_7910,N_2052,N_3969);
nor U7911 (N_7911,N_2286,N_40);
nor U7912 (N_7912,N_2116,N_526);
or U7913 (N_7913,N_416,N_3604);
nand U7914 (N_7914,N_3736,N_4877);
or U7915 (N_7915,N_2236,N_1917);
nand U7916 (N_7916,N_65,N_4977);
nor U7917 (N_7917,N_3209,N_2814);
or U7918 (N_7918,N_3352,N_4521);
and U7919 (N_7919,N_4594,N_2172);
and U7920 (N_7920,N_2330,N_3854);
and U7921 (N_7921,N_3099,N_3118);
nand U7922 (N_7922,N_1025,N_4582);
nor U7923 (N_7923,N_676,N_4492);
nor U7924 (N_7924,N_1617,N_1714);
xnor U7925 (N_7925,N_46,N_3591);
and U7926 (N_7926,N_3536,N_4535);
nand U7927 (N_7927,N_3427,N_727);
nor U7928 (N_7928,N_3001,N_1656);
nor U7929 (N_7929,N_351,N_3939);
and U7930 (N_7930,N_1845,N_1083);
nand U7931 (N_7931,N_3518,N_2264);
and U7932 (N_7932,N_1160,N_912);
nand U7933 (N_7933,N_2738,N_4306);
nand U7934 (N_7934,N_310,N_638);
or U7935 (N_7935,N_3317,N_4548);
nand U7936 (N_7936,N_2217,N_230);
or U7937 (N_7937,N_2942,N_2499);
or U7938 (N_7938,N_4416,N_29);
and U7939 (N_7939,N_549,N_1438);
and U7940 (N_7940,N_1144,N_628);
and U7941 (N_7941,N_4000,N_3907);
and U7942 (N_7942,N_2997,N_2702);
nand U7943 (N_7943,N_1652,N_4160);
and U7944 (N_7944,N_3513,N_863);
and U7945 (N_7945,N_3176,N_3258);
or U7946 (N_7946,N_202,N_4505);
nor U7947 (N_7947,N_1828,N_585);
and U7948 (N_7948,N_2746,N_4916);
nand U7949 (N_7949,N_4867,N_2974);
or U7950 (N_7950,N_2943,N_4229);
nor U7951 (N_7951,N_2181,N_1783);
nand U7952 (N_7952,N_4049,N_601);
nor U7953 (N_7953,N_2522,N_4618);
nor U7954 (N_7954,N_4918,N_3745);
nand U7955 (N_7955,N_1129,N_1872);
and U7956 (N_7956,N_2280,N_2313);
or U7957 (N_7957,N_406,N_2192);
or U7958 (N_7958,N_3247,N_1315);
nor U7959 (N_7959,N_3618,N_221);
or U7960 (N_7960,N_4825,N_855);
nor U7961 (N_7961,N_2698,N_3044);
nand U7962 (N_7962,N_1542,N_3081);
and U7963 (N_7963,N_3133,N_4442);
or U7964 (N_7964,N_506,N_2442);
nand U7965 (N_7965,N_1684,N_1750);
and U7966 (N_7966,N_3519,N_3263);
nand U7967 (N_7967,N_2327,N_3057);
nand U7968 (N_7968,N_4354,N_2060);
xor U7969 (N_7969,N_1538,N_1337);
nor U7970 (N_7970,N_2738,N_1846);
and U7971 (N_7971,N_1096,N_3827);
or U7972 (N_7972,N_395,N_1583);
nor U7973 (N_7973,N_3994,N_149);
nor U7974 (N_7974,N_553,N_3509);
nand U7975 (N_7975,N_3900,N_2626);
or U7976 (N_7976,N_2238,N_4823);
and U7977 (N_7977,N_3892,N_1357);
nand U7978 (N_7978,N_2488,N_1593);
or U7979 (N_7979,N_2250,N_483);
nand U7980 (N_7980,N_2707,N_1764);
and U7981 (N_7981,N_4990,N_3870);
nand U7982 (N_7982,N_3225,N_4880);
nand U7983 (N_7983,N_3263,N_2236);
or U7984 (N_7984,N_2448,N_1461);
nand U7985 (N_7985,N_3218,N_3560);
and U7986 (N_7986,N_3430,N_4693);
nand U7987 (N_7987,N_1057,N_1572);
or U7988 (N_7988,N_2982,N_4583);
nand U7989 (N_7989,N_3319,N_3732);
nand U7990 (N_7990,N_622,N_4577);
and U7991 (N_7991,N_2428,N_1945);
nand U7992 (N_7992,N_3590,N_4563);
nor U7993 (N_7993,N_1554,N_4790);
and U7994 (N_7994,N_1712,N_2469);
nand U7995 (N_7995,N_3355,N_2339);
nand U7996 (N_7996,N_574,N_189);
nor U7997 (N_7997,N_2301,N_1794);
and U7998 (N_7998,N_1891,N_4190);
and U7999 (N_7999,N_3571,N_1993);
nand U8000 (N_8000,N_1139,N_3909);
and U8001 (N_8001,N_954,N_991);
nand U8002 (N_8002,N_943,N_952);
nand U8003 (N_8003,N_3584,N_926);
nand U8004 (N_8004,N_2303,N_2430);
nor U8005 (N_8005,N_4470,N_554);
nand U8006 (N_8006,N_4225,N_765);
or U8007 (N_8007,N_625,N_936);
and U8008 (N_8008,N_3110,N_2695);
nor U8009 (N_8009,N_3220,N_3674);
nand U8010 (N_8010,N_4961,N_3729);
nand U8011 (N_8011,N_4546,N_3505);
nor U8012 (N_8012,N_3899,N_1951);
nand U8013 (N_8013,N_3206,N_4916);
and U8014 (N_8014,N_1075,N_741);
nand U8015 (N_8015,N_3398,N_1699);
nor U8016 (N_8016,N_3278,N_4559);
and U8017 (N_8017,N_3713,N_524);
or U8018 (N_8018,N_2045,N_2420);
and U8019 (N_8019,N_2984,N_1787);
nor U8020 (N_8020,N_1963,N_4145);
nor U8021 (N_8021,N_2368,N_1761);
nor U8022 (N_8022,N_1201,N_2652);
nand U8023 (N_8023,N_1200,N_4351);
and U8024 (N_8024,N_4203,N_4738);
or U8025 (N_8025,N_574,N_4352);
nor U8026 (N_8026,N_2584,N_3368);
nor U8027 (N_8027,N_2685,N_2741);
and U8028 (N_8028,N_2576,N_1590);
nand U8029 (N_8029,N_78,N_769);
nor U8030 (N_8030,N_3693,N_3840);
and U8031 (N_8031,N_3917,N_4131);
nand U8032 (N_8032,N_4604,N_3740);
nor U8033 (N_8033,N_544,N_4608);
nor U8034 (N_8034,N_461,N_4506);
and U8035 (N_8035,N_2753,N_1687);
and U8036 (N_8036,N_2530,N_571);
nor U8037 (N_8037,N_3138,N_4725);
or U8038 (N_8038,N_2071,N_1315);
or U8039 (N_8039,N_3355,N_2494);
nor U8040 (N_8040,N_289,N_523);
nand U8041 (N_8041,N_532,N_3713);
nand U8042 (N_8042,N_596,N_193);
and U8043 (N_8043,N_2433,N_378);
or U8044 (N_8044,N_2024,N_3833);
or U8045 (N_8045,N_690,N_189);
or U8046 (N_8046,N_1435,N_2223);
or U8047 (N_8047,N_2139,N_3179);
and U8048 (N_8048,N_4432,N_771);
and U8049 (N_8049,N_584,N_2980);
and U8050 (N_8050,N_4712,N_1039);
and U8051 (N_8051,N_2295,N_3911);
nand U8052 (N_8052,N_4828,N_2328);
nor U8053 (N_8053,N_3507,N_4368);
nand U8054 (N_8054,N_923,N_1000);
nor U8055 (N_8055,N_4167,N_4838);
nor U8056 (N_8056,N_1139,N_3723);
nand U8057 (N_8057,N_3961,N_4074);
or U8058 (N_8058,N_1221,N_2321);
nand U8059 (N_8059,N_1978,N_4162);
and U8060 (N_8060,N_1736,N_932);
or U8061 (N_8061,N_1614,N_1946);
and U8062 (N_8062,N_3731,N_4024);
nor U8063 (N_8063,N_3964,N_2777);
and U8064 (N_8064,N_3901,N_28);
nor U8065 (N_8065,N_1697,N_547);
nand U8066 (N_8066,N_4098,N_3937);
and U8067 (N_8067,N_4160,N_3381);
nor U8068 (N_8068,N_332,N_1489);
nand U8069 (N_8069,N_1764,N_1189);
nand U8070 (N_8070,N_302,N_1116);
and U8071 (N_8071,N_2184,N_4570);
nor U8072 (N_8072,N_1645,N_3777);
nor U8073 (N_8073,N_1431,N_1536);
nor U8074 (N_8074,N_1194,N_2372);
nor U8075 (N_8075,N_4833,N_2993);
or U8076 (N_8076,N_2836,N_3935);
nand U8077 (N_8077,N_1376,N_199);
and U8078 (N_8078,N_3288,N_4651);
nor U8079 (N_8079,N_4291,N_249);
nand U8080 (N_8080,N_2385,N_1629);
or U8081 (N_8081,N_265,N_569);
xnor U8082 (N_8082,N_2271,N_2698);
and U8083 (N_8083,N_4174,N_2575);
nor U8084 (N_8084,N_726,N_3976);
and U8085 (N_8085,N_964,N_3350);
or U8086 (N_8086,N_2806,N_1681);
or U8087 (N_8087,N_3329,N_3514);
and U8088 (N_8088,N_2041,N_4946);
nor U8089 (N_8089,N_4063,N_3131);
or U8090 (N_8090,N_1398,N_1425);
nand U8091 (N_8091,N_1356,N_1929);
or U8092 (N_8092,N_1855,N_4413);
or U8093 (N_8093,N_2242,N_2142);
and U8094 (N_8094,N_2622,N_218);
and U8095 (N_8095,N_1744,N_4054);
xnor U8096 (N_8096,N_3256,N_1432);
nand U8097 (N_8097,N_2503,N_4445);
nor U8098 (N_8098,N_3065,N_4920);
nor U8099 (N_8099,N_1205,N_3508);
and U8100 (N_8100,N_2790,N_687);
nand U8101 (N_8101,N_4702,N_2054);
nand U8102 (N_8102,N_1539,N_819);
xnor U8103 (N_8103,N_4592,N_3687);
or U8104 (N_8104,N_3193,N_1497);
or U8105 (N_8105,N_1838,N_3147);
nor U8106 (N_8106,N_3305,N_3500);
or U8107 (N_8107,N_162,N_3082);
and U8108 (N_8108,N_1106,N_3703);
or U8109 (N_8109,N_3056,N_2564);
xnor U8110 (N_8110,N_2980,N_3654);
or U8111 (N_8111,N_3614,N_1411);
or U8112 (N_8112,N_4908,N_3769);
and U8113 (N_8113,N_3617,N_4374);
nand U8114 (N_8114,N_857,N_928);
nand U8115 (N_8115,N_3573,N_4745);
and U8116 (N_8116,N_2070,N_2594);
nand U8117 (N_8117,N_309,N_4005);
nor U8118 (N_8118,N_1313,N_4581);
nand U8119 (N_8119,N_2115,N_4314);
or U8120 (N_8120,N_2764,N_53);
nand U8121 (N_8121,N_4411,N_2382);
and U8122 (N_8122,N_463,N_1460);
nor U8123 (N_8123,N_3117,N_1138);
nand U8124 (N_8124,N_296,N_949);
nand U8125 (N_8125,N_163,N_4876);
and U8126 (N_8126,N_2120,N_2010);
or U8127 (N_8127,N_2664,N_1452);
nand U8128 (N_8128,N_2898,N_527);
or U8129 (N_8129,N_84,N_1798);
nor U8130 (N_8130,N_3061,N_4006);
nor U8131 (N_8131,N_4030,N_1836);
nand U8132 (N_8132,N_2480,N_2110);
nor U8133 (N_8133,N_4703,N_4011);
or U8134 (N_8134,N_2081,N_2077);
and U8135 (N_8135,N_373,N_1261);
nand U8136 (N_8136,N_911,N_3558);
or U8137 (N_8137,N_611,N_4235);
or U8138 (N_8138,N_4640,N_2963);
nand U8139 (N_8139,N_1065,N_1574);
nand U8140 (N_8140,N_2073,N_3660);
nor U8141 (N_8141,N_3435,N_4882);
nand U8142 (N_8142,N_4747,N_2698);
nor U8143 (N_8143,N_4956,N_4951);
nor U8144 (N_8144,N_3434,N_3509);
nor U8145 (N_8145,N_1340,N_1536);
and U8146 (N_8146,N_1366,N_265);
and U8147 (N_8147,N_4790,N_4552);
nand U8148 (N_8148,N_3178,N_178);
nand U8149 (N_8149,N_4628,N_4709);
nor U8150 (N_8150,N_1459,N_2320);
and U8151 (N_8151,N_1801,N_3948);
nand U8152 (N_8152,N_1673,N_4551);
nand U8153 (N_8153,N_1038,N_2296);
xnor U8154 (N_8154,N_2556,N_2161);
nor U8155 (N_8155,N_4372,N_4655);
nor U8156 (N_8156,N_859,N_2961);
nand U8157 (N_8157,N_3694,N_606);
nand U8158 (N_8158,N_3244,N_4687);
nand U8159 (N_8159,N_966,N_664);
nor U8160 (N_8160,N_3784,N_2703);
nand U8161 (N_8161,N_3026,N_1926);
and U8162 (N_8162,N_3256,N_667);
nor U8163 (N_8163,N_2303,N_3455);
or U8164 (N_8164,N_3539,N_848);
or U8165 (N_8165,N_2408,N_2047);
or U8166 (N_8166,N_4017,N_3309);
nor U8167 (N_8167,N_4779,N_4199);
and U8168 (N_8168,N_4589,N_3755);
or U8169 (N_8169,N_1831,N_1163);
nand U8170 (N_8170,N_2792,N_2687);
nand U8171 (N_8171,N_2295,N_6);
or U8172 (N_8172,N_282,N_2778);
nor U8173 (N_8173,N_3012,N_3281);
nor U8174 (N_8174,N_826,N_946);
and U8175 (N_8175,N_2312,N_4942);
or U8176 (N_8176,N_3543,N_672);
and U8177 (N_8177,N_4302,N_1100);
nor U8178 (N_8178,N_2387,N_1774);
and U8179 (N_8179,N_4487,N_4536);
xnor U8180 (N_8180,N_2895,N_3501);
and U8181 (N_8181,N_4745,N_2717);
nand U8182 (N_8182,N_4961,N_2597);
or U8183 (N_8183,N_4403,N_4238);
nand U8184 (N_8184,N_1535,N_3055);
or U8185 (N_8185,N_1784,N_1857);
nand U8186 (N_8186,N_950,N_2001);
nor U8187 (N_8187,N_4198,N_2267);
and U8188 (N_8188,N_3093,N_3990);
and U8189 (N_8189,N_4516,N_173);
nor U8190 (N_8190,N_3272,N_2664);
or U8191 (N_8191,N_2470,N_1825);
nor U8192 (N_8192,N_2387,N_1762);
or U8193 (N_8193,N_282,N_2578);
and U8194 (N_8194,N_1835,N_1924);
nor U8195 (N_8195,N_3717,N_1290);
nor U8196 (N_8196,N_70,N_669);
nor U8197 (N_8197,N_3519,N_2538);
or U8198 (N_8198,N_3639,N_2620);
nand U8199 (N_8199,N_2119,N_3863);
nand U8200 (N_8200,N_2429,N_2712);
and U8201 (N_8201,N_2882,N_1658);
nand U8202 (N_8202,N_342,N_2720);
nor U8203 (N_8203,N_4440,N_4477);
nor U8204 (N_8204,N_2319,N_4870);
nand U8205 (N_8205,N_1069,N_3197);
or U8206 (N_8206,N_1804,N_295);
or U8207 (N_8207,N_2791,N_3756);
or U8208 (N_8208,N_4923,N_2307);
nand U8209 (N_8209,N_2435,N_4007);
nand U8210 (N_8210,N_2689,N_4347);
and U8211 (N_8211,N_4687,N_3035);
nand U8212 (N_8212,N_1540,N_4716);
nand U8213 (N_8213,N_3875,N_4932);
and U8214 (N_8214,N_609,N_4031);
and U8215 (N_8215,N_3302,N_4662);
nor U8216 (N_8216,N_632,N_777);
xnor U8217 (N_8217,N_3365,N_2624);
nor U8218 (N_8218,N_3115,N_1143);
nor U8219 (N_8219,N_3652,N_2476);
and U8220 (N_8220,N_2201,N_1674);
or U8221 (N_8221,N_3106,N_1762);
nand U8222 (N_8222,N_3890,N_653);
and U8223 (N_8223,N_3975,N_31);
nand U8224 (N_8224,N_2264,N_4987);
and U8225 (N_8225,N_4300,N_4826);
nor U8226 (N_8226,N_3416,N_4064);
and U8227 (N_8227,N_2344,N_1983);
or U8228 (N_8228,N_4012,N_3484);
nand U8229 (N_8229,N_3138,N_405);
and U8230 (N_8230,N_494,N_4031);
or U8231 (N_8231,N_2235,N_4316);
nand U8232 (N_8232,N_2017,N_435);
nor U8233 (N_8233,N_644,N_2651);
and U8234 (N_8234,N_1579,N_1983);
nand U8235 (N_8235,N_1701,N_734);
and U8236 (N_8236,N_4654,N_1612);
nand U8237 (N_8237,N_4712,N_2538);
or U8238 (N_8238,N_3292,N_4020);
nand U8239 (N_8239,N_962,N_2899);
nand U8240 (N_8240,N_2957,N_4929);
xnor U8241 (N_8241,N_1515,N_2561);
or U8242 (N_8242,N_1284,N_162);
nor U8243 (N_8243,N_4525,N_1059);
or U8244 (N_8244,N_105,N_2241);
or U8245 (N_8245,N_3965,N_2051);
or U8246 (N_8246,N_3639,N_1889);
and U8247 (N_8247,N_1928,N_3465);
nand U8248 (N_8248,N_2723,N_2394);
and U8249 (N_8249,N_2923,N_1773);
nor U8250 (N_8250,N_879,N_893);
nor U8251 (N_8251,N_4829,N_246);
and U8252 (N_8252,N_3915,N_1520);
nand U8253 (N_8253,N_308,N_4433);
nand U8254 (N_8254,N_2628,N_1872);
and U8255 (N_8255,N_2479,N_3368);
nor U8256 (N_8256,N_284,N_2065);
and U8257 (N_8257,N_1366,N_1578);
nand U8258 (N_8258,N_437,N_374);
and U8259 (N_8259,N_4629,N_1572);
nand U8260 (N_8260,N_2148,N_1181);
and U8261 (N_8261,N_4451,N_336);
or U8262 (N_8262,N_4306,N_1354);
nand U8263 (N_8263,N_1928,N_4411);
and U8264 (N_8264,N_3275,N_1813);
or U8265 (N_8265,N_3147,N_2800);
nor U8266 (N_8266,N_1451,N_261);
or U8267 (N_8267,N_4998,N_3886);
nand U8268 (N_8268,N_1692,N_1477);
or U8269 (N_8269,N_4769,N_109);
and U8270 (N_8270,N_3828,N_292);
or U8271 (N_8271,N_2818,N_586);
or U8272 (N_8272,N_4963,N_993);
nor U8273 (N_8273,N_2275,N_3874);
nor U8274 (N_8274,N_3843,N_1762);
nand U8275 (N_8275,N_3150,N_4503);
nor U8276 (N_8276,N_3697,N_2997);
and U8277 (N_8277,N_236,N_2970);
nand U8278 (N_8278,N_2662,N_194);
and U8279 (N_8279,N_1035,N_583);
nor U8280 (N_8280,N_4971,N_3281);
and U8281 (N_8281,N_4942,N_1953);
nor U8282 (N_8282,N_1493,N_3789);
nor U8283 (N_8283,N_3436,N_2619);
or U8284 (N_8284,N_4401,N_1978);
nor U8285 (N_8285,N_2222,N_2531);
nand U8286 (N_8286,N_1372,N_4106);
nor U8287 (N_8287,N_4968,N_2810);
nor U8288 (N_8288,N_4160,N_1361);
or U8289 (N_8289,N_2302,N_2594);
nor U8290 (N_8290,N_2096,N_35);
or U8291 (N_8291,N_3807,N_277);
or U8292 (N_8292,N_1503,N_1065);
or U8293 (N_8293,N_4515,N_4353);
nor U8294 (N_8294,N_2255,N_2043);
nand U8295 (N_8295,N_2503,N_3071);
or U8296 (N_8296,N_2385,N_2979);
nand U8297 (N_8297,N_4260,N_218);
nand U8298 (N_8298,N_1651,N_1338);
nand U8299 (N_8299,N_1523,N_4766);
nor U8300 (N_8300,N_1949,N_1417);
nor U8301 (N_8301,N_3528,N_1137);
nor U8302 (N_8302,N_2036,N_717);
or U8303 (N_8303,N_2187,N_902);
nor U8304 (N_8304,N_997,N_2034);
and U8305 (N_8305,N_1751,N_2539);
and U8306 (N_8306,N_3032,N_2203);
or U8307 (N_8307,N_1715,N_2654);
nor U8308 (N_8308,N_2070,N_1553);
nand U8309 (N_8309,N_223,N_2032);
and U8310 (N_8310,N_4434,N_4643);
nand U8311 (N_8311,N_4945,N_1918);
or U8312 (N_8312,N_588,N_4679);
nand U8313 (N_8313,N_3511,N_838);
nand U8314 (N_8314,N_505,N_669);
nand U8315 (N_8315,N_3498,N_2718);
nand U8316 (N_8316,N_4473,N_1880);
or U8317 (N_8317,N_1518,N_3460);
and U8318 (N_8318,N_3435,N_2163);
nand U8319 (N_8319,N_761,N_2631);
and U8320 (N_8320,N_1405,N_88);
or U8321 (N_8321,N_1234,N_1059);
and U8322 (N_8322,N_4262,N_443);
nand U8323 (N_8323,N_2919,N_514);
and U8324 (N_8324,N_4506,N_1991);
and U8325 (N_8325,N_3063,N_1267);
nor U8326 (N_8326,N_4272,N_2289);
or U8327 (N_8327,N_2395,N_2447);
nand U8328 (N_8328,N_211,N_1581);
nor U8329 (N_8329,N_2660,N_477);
or U8330 (N_8330,N_126,N_395);
nand U8331 (N_8331,N_3471,N_3467);
nand U8332 (N_8332,N_3687,N_1806);
nor U8333 (N_8333,N_1763,N_3501);
and U8334 (N_8334,N_485,N_1412);
or U8335 (N_8335,N_4145,N_2500);
nor U8336 (N_8336,N_4384,N_1840);
and U8337 (N_8337,N_4665,N_345);
and U8338 (N_8338,N_4004,N_2534);
or U8339 (N_8339,N_911,N_4361);
or U8340 (N_8340,N_3471,N_1290);
or U8341 (N_8341,N_1412,N_3992);
or U8342 (N_8342,N_2738,N_2778);
nand U8343 (N_8343,N_2854,N_3614);
and U8344 (N_8344,N_2864,N_2283);
nand U8345 (N_8345,N_2981,N_1506);
nor U8346 (N_8346,N_365,N_1106);
and U8347 (N_8347,N_1529,N_868);
or U8348 (N_8348,N_826,N_1527);
and U8349 (N_8349,N_1917,N_4180);
and U8350 (N_8350,N_4197,N_2631);
nor U8351 (N_8351,N_4589,N_3031);
or U8352 (N_8352,N_662,N_1867);
or U8353 (N_8353,N_1108,N_4577);
nor U8354 (N_8354,N_1492,N_1915);
nor U8355 (N_8355,N_2952,N_2947);
nand U8356 (N_8356,N_570,N_4587);
and U8357 (N_8357,N_3689,N_2300);
and U8358 (N_8358,N_1017,N_1472);
or U8359 (N_8359,N_174,N_889);
nand U8360 (N_8360,N_1518,N_2264);
and U8361 (N_8361,N_4147,N_4263);
or U8362 (N_8362,N_2411,N_132);
or U8363 (N_8363,N_2491,N_2108);
or U8364 (N_8364,N_1886,N_908);
nor U8365 (N_8365,N_3689,N_796);
or U8366 (N_8366,N_1614,N_3290);
nor U8367 (N_8367,N_4931,N_2394);
nor U8368 (N_8368,N_3407,N_4354);
nor U8369 (N_8369,N_2144,N_4052);
nor U8370 (N_8370,N_4972,N_3150);
xnor U8371 (N_8371,N_3109,N_1085);
or U8372 (N_8372,N_647,N_4889);
or U8373 (N_8373,N_1472,N_829);
and U8374 (N_8374,N_3588,N_3833);
nor U8375 (N_8375,N_3766,N_4607);
and U8376 (N_8376,N_2879,N_3461);
and U8377 (N_8377,N_4899,N_1222);
and U8378 (N_8378,N_3196,N_4517);
nor U8379 (N_8379,N_2800,N_2996);
nand U8380 (N_8380,N_3540,N_1217);
nand U8381 (N_8381,N_4910,N_418);
and U8382 (N_8382,N_3998,N_3);
and U8383 (N_8383,N_750,N_1914);
xnor U8384 (N_8384,N_465,N_2750);
nor U8385 (N_8385,N_1105,N_1600);
and U8386 (N_8386,N_1749,N_1485);
and U8387 (N_8387,N_339,N_4301);
and U8388 (N_8388,N_4675,N_1575);
nand U8389 (N_8389,N_1512,N_2736);
or U8390 (N_8390,N_1657,N_3079);
nand U8391 (N_8391,N_4362,N_1204);
and U8392 (N_8392,N_3507,N_3540);
or U8393 (N_8393,N_4898,N_1850);
or U8394 (N_8394,N_1493,N_3379);
nand U8395 (N_8395,N_3634,N_2388);
nand U8396 (N_8396,N_1108,N_1717);
nor U8397 (N_8397,N_2215,N_953);
nor U8398 (N_8398,N_3426,N_4922);
and U8399 (N_8399,N_3120,N_4355);
xor U8400 (N_8400,N_904,N_4057);
nand U8401 (N_8401,N_2827,N_4027);
and U8402 (N_8402,N_4862,N_1311);
or U8403 (N_8403,N_3326,N_700);
or U8404 (N_8404,N_3149,N_2627);
nand U8405 (N_8405,N_2248,N_3184);
nor U8406 (N_8406,N_1022,N_4426);
nand U8407 (N_8407,N_726,N_4644);
nand U8408 (N_8408,N_2771,N_2633);
and U8409 (N_8409,N_232,N_1644);
or U8410 (N_8410,N_1007,N_3956);
nor U8411 (N_8411,N_1477,N_178);
and U8412 (N_8412,N_3131,N_2920);
nor U8413 (N_8413,N_975,N_4275);
and U8414 (N_8414,N_4764,N_614);
and U8415 (N_8415,N_1717,N_3785);
or U8416 (N_8416,N_109,N_2718);
nor U8417 (N_8417,N_1466,N_1329);
or U8418 (N_8418,N_2136,N_4247);
nor U8419 (N_8419,N_149,N_1187);
or U8420 (N_8420,N_3889,N_4860);
nand U8421 (N_8421,N_2665,N_1544);
or U8422 (N_8422,N_61,N_938);
nand U8423 (N_8423,N_3824,N_4543);
or U8424 (N_8424,N_2077,N_2593);
or U8425 (N_8425,N_958,N_1867);
and U8426 (N_8426,N_343,N_3912);
nor U8427 (N_8427,N_2522,N_2826);
or U8428 (N_8428,N_1155,N_1432);
nor U8429 (N_8429,N_2272,N_2756);
or U8430 (N_8430,N_890,N_3771);
or U8431 (N_8431,N_4508,N_2100);
nand U8432 (N_8432,N_4977,N_3928);
or U8433 (N_8433,N_971,N_2266);
nor U8434 (N_8434,N_3816,N_663);
nand U8435 (N_8435,N_243,N_680);
and U8436 (N_8436,N_486,N_1474);
nor U8437 (N_8437,N_2355,N_2275);
and U8438 (N_8438,N_2279,N_3465);
nor U8439 (N_8439,N_3025,N_3766);
and U8440 (N_8440,N_3413,N_3724);
or U8441 (N_8441,N_2928,N_1687);
or U8442 (N_8442,N_352,N_3450);
and U8443 (N_8443,N_746,N_1348);
nor U8444 (N_8444,N_213,N_4262);
or U8445 (N_8445,N_4110,N_4358);
and U8446 (N_8446,N_3019,N_3693);
nor U8447 (N_8447,N_1184,N_2348);
nand U8448 (N_8448,N_1202,N_338);
nor U8449 (N_8449,N_4960,N_2684);
or U8450 (N_8450,N_3105,N_1244);
nor U8451 (N_8451,N_4222,N_3742);
nor U8452 (N_8452,N_4131,N_2591);
and U8453 (N_8453,N_460,N_908);
or U8454 (N_8454,N_1939,N_1900);
nor U8455 (N_8455,N_4410,N_1497);
and U8456 (N_8456,N_1438,N_3445);
or U8457 (N_8457,N_3585,N_2187);
nand U8458 (N_8458,N_779,N_582);
nor U8459 (N_8459,N_2701,N_4118);
xnor U8460 (N_8460,N_1458,N_3668);
nand U8461 (N_8461,N_1261,N_4328);
and U8462 (N_8462,N_3415,N_1870);
or U8463 (N_8463,N_2314,N_2395);
nand U8464 (N_8464,N_310,N_4078);
or U8465 (N_8465,N_1620,N_3319);
or U8466 (N_8466,N_4520,N_3162);
nand U8467 (N_8467,N_3066,N_2831);
and U8468 (N_8468,N_4448,N_1020);
and U8469 (N_8469,N_2477,N_595);
nor U8470 (N_8470,N_638,N_2776);
nand U8471 (N_8471,N_1493,N_270);
and U8472 (N_8472,N_4037,N_4828);
and U8473 (N_8473,N_937,N_4605);
nor U8474 (N_8474,N_2079,N_3673);
and U8475 (N_8475,N_3014,N_2335);
nor U8476 (N_8476,N_431,N_609);
nand U8477 (N_8477,N_267,N_3802);
nand U8478 (N_8478,N_4830,N_1007);
nand U8479 (N_8479,N_3848,N_2022);
nand U8480 (N_8480,N_733,N_1476);
nand U8481 (N_8481,N_3683,N_3563);
and U8482 (N_8482,N_4858,N_4219);
nand U8483 (N_8483,N_2541,N_3897);
and U8484 (N_8484,N_2474,N_134);
or U8485 (N_8485,N_3509,N_4479);
nand U8486 (N_8486,N_4993,N_2431);
nand U8487 (N_8487,N_2204,N_4196);
nand U8488 (N_8488,N_2555,N_3315);
nand U8489 (N_8489,N_3546,N_2868);
nand U8490 (N_8490,N_3919,N_2738);
nand U8491 (N_8491,N_894,N_4489);
and U8492 (N_8492,N_710,N_3492);
and U8493 (N_8493,N_4400,N_2008);
nand U8494 (N_8494,N_4177,N_41);
nand U8495 (N_8495,N_4424,N_1353);
nor U8496 (N_8496,N_2462,N_3212);
or U8497 (N_8497,N_4626,N_598);
nand U8498 (N_8498,N_4920,N_3816);
nand U8499 (N_8499,N_2008,N_2102);
nor U8500 (N_8500,N_3397,N_905);
or U8501 (N_8501,N_2856,N_4949);
nor U8502 (N_8502,N_3358,N_4075);
xor U8503 (N_8503,N_1003,N_3470);
nand U8504 (N_8504,N_2603,N_1237);
nand U8505 (N_8505,N_1959,N_1774);
or U8506 (N_8506,N_556,N_4723);
or U8507 (N_8507,N_2564,N_831);
xor U8508 (N_8508,N_1750,N_244);
and U8509 (N_8509,N_3900,N_1737);
or U8510 (N_8510,N_914,N_4394);
nand U8511 (N_8511,N_368,N_1012);
nor U8512 (N_8512,N_1787,N_1285);
nor U8513 (N_8513,N_3999,N_2565);
and U8514 (N_8514,N_843,N_2669);
nand U8515 (N_8515,N_2025,N_4360);
nor U8516 (N_8516,N_4924,N_4099);
or U8517 (N_8517,N_73,N_941);
or U8518 (N_8518,N_890,N_2206);
or U8519 (N_8519,N_3298,N_2964);
and U8520 (N_8520,N_4298,N_4719);
or U8521 (N_8521,N_3579,N_3942);
nor U8522 (N_8522,N_3212,N_879);
and U8523 (N_8523,N_2995,N_2897);
and U8524 (N_8524,N_874,N_4060);
nor U8525 (N_8525,N_2584,N_4283);
nand U8526 (N_8526,N_601,N_1242);
nor U8527 (N_8527,N_3147,N_3945);
nand U8528 (N_8528,N_4947,N_3814);
or U8529 (N_8529,N_1785,N_2794);
or U8530 (N_8530,N_519,N_4233);
and U8531 (N_8531,N_3568,N_2455);
or U8532 (N_8532,N_3462,N_3155);
and U8533 (N_8533,N_915,N_958);
nor U8534 (N_8534,N_911,N_882);
or U8535 (N_8535,N_1391,N_3973);
or U8536 (N_8536,N_4909,N_1532);
and U8537 (N_8537,N_451,N_1486);
and U8538 (N_8538,N_1811,N_4236);
nand U8539 (N_8539,N_2959,N_354);
and U8540 (N_8540,N_4378,N_3932);
xnor U8541 (N_8541,N_3597,N_609);
or U8542 (N_8542,N_420,N_1668);
nand U8543 (N_8543,N_3216,N_2776);
and U8544 (N_8544,N_3355,N_2707);
nand U8545 (N_8545,N_257,N_2818);
nand U8546 (N_8546,N_1982,N_1150);
and U8547 (N_8547,N_3450,N_2961);
or U8548 (N_8548,N_2161,N_2836);
nor U8549 (N_8549,N_2181,N_1887);
and U8550 (N_8550,N_854,N_1342);
or U8551 (N_8551,N_2309,N_1063);
nand U8552 (N_8552,N_1372,N_4740);
nand U8553 (N_8553,N_3209,N_810);
or U8554 (N_8554,N_2390,N_4653);
nor U8555 (N_8555,N_4221,N_2010);
or U8556 (N_8556,N_3766,N_1837);
or U8557 (N_8557,N_1120,N_981);
and U8558 (N_8558,N_4101,N_2006);
and U8559 (N_8559,N_1021,N_4335);
nor U8560 (N_8560,N_4860,N_3651);
nor U8561 (N_8561,N_547,N_569);
and U8562 (N_8562,N_2730,N_4415);
nor U8563 (N_8563,N_165,N_4517);
nor U8564 (N_8564,N_1301,N_102);
and U8565 (N_8565,N_4352,N_2771);
or U8566 (N_8566,N_3616,N_3978);
and U8567 (N_8567,N_2319,N_2794);
or U8568 (N_8568,N_50,N_2770);
and U8569 (N_8569,N_2924,N_2784);
and U8570 (N_8570,N_3130,N_1759);
nand U8571 (N_8571,N_1981,N_559);
and U8572 (N_8572,N_3958,N_4098);
or U8573 (N_8573,N_4803,N_4212);
nor U8574 (N_8574,N_3394,N_250);
nor U8575 (N_8575,N_1845,N_533);
nand U8576 (N_8576,N_132,N_4606);
nand U8577 (N_8577,N_446,N_1247);
nand U8578 (N_8578,N_899,N_468);
and U8579 (N_8579,N_3316,N_4930);
nand U8580 (N_8580,N_4167,N_4100);
and U8581 (N_8581,N_3040,N_3390);
nand U8582 (N_8582,N_2835,N_993);
nor U8583 (N_8583,N_4120,N_987);
and U8584 (N_8584,N_3074,N_317);
nand U8585 (N_8585,N_1752,N_2202);
nand U8586 (N_8586,N_2491,N_1358);
or U8587 (N_8587,N_2836,N_924);
nor U8588 (N_8588,N_1878,N_250);
nand U8589 (N_8589,N_99,N_2440);
and U8590 (N_8590,N_1408,N_2302);
nand U8591 (N_8591,N_3802,N_465);
nor U8592 (N_8592,N_158,N_2412);
nor U8593 (N_8593,N_3092,N_1295);
nor U8594 (N_8594,N_3646,N_2071);
or U8595 (N_8595,N_4184,N_395);
nand U8596 (N_8596,N_1054,N_3847);
nand U8597 (N_8597,N_2256,N_1309);
nand U8598 (N_8598,N_748,N_3095);
nor U8599 (N_8599,N_82,N_2588);
nor U8600 (N_8600,N_4121,N_936);
or U8601 (N_8601,N_4796,N_399);
nor U8602 (N_8602,N_3744,N_4536);
and U8603 (N_8603,N_1808,N_1240);
nor U8604 (N_8604,N_738,N_2579);
and U8605 (N_8605,N_2990,N_2421);
nand U8606 (N_8606,N_1417,N_3147);
nand U8607 (N_8607,N_4401,N_2603);
nor U8608 (N_8608,N_1710,N_794);
nor U8609 (N_8609,N_1565,N_2949);
xor U8610 (N_8610,N_2021,N_1978);
nor U8611 (N_8611,N_683,N_2517);
and U8612 (N_8612,N_1426,N_383);
nand U8613 (N_8613,N_2878,N_3315);
nand U8614 (N_8614,N_1098,N_2855);
nor U8615 (N_8615,N_2492,N_1159);
nand U8616 (N_8616,N_4230,N_4126);
and U8617 (N_8617,N_3672,N_42);
or U8618 (N_8618,N_4982,N_380);
nand U8619 (N_8619,N_3370,N_1963);
and U8620 (N_8620,N_2615,N_4168);
nor U8621 (N_8621,N_3911,N_4032);
or U8622 (N_8622,N_2016,N_3273);
nor U8623 (N_8623,N_163,N_918);
or U8624 (N_8624,N_3338,N_1128);
nand U8625 (N_8625,N_885,N_3971);
nand U8626 (N_8626,N_3926,N_3595);
nor U8627 (N_8627,N_4211,N_1102);
or U8628 (N_8628,N_470,N_3983);
nor U8629 (N_8629,N_1392,N_1050);
or U8630 (N_8630,N_1865,N_4653);
and U8631 (N_8631,N_2386,N_4210);
nand U8632 (N_8632,N_4979,N_723);
or U8633 (N_8633,N_4306,N_4015);
and U8634 (N_8634,N_290,N_4840);
nand U8635 (N_8635,N_1719,N_2507);
and U8636 (N_8636,N_4709,N_383);
nand U8637 (N_8637,N_2472,N_2183);
nor U8638 (N_8638,N_2503,N_1644);
and U8639 (N_8639,N_4684,N_1308);
nand U8640 (N_8640,N_4850,N_1023);
nand U8641 (N_8641,N_649,N_1140);
or U8642 (N_8642,N_554,N_553);
or U8643 (N_8643,N_660,N_488);
or U8644 (N_8644,N_3104,N_4525);
and U8645 (N_8645,N_2975,N_1958);
and U8646 (N_8646,N_39,N_3581);
or U8647 (N_8647,N_3702,N_1431);
nor U8648 (N_8648,N_4276,N_3885);
nand U8649 (N_8649,N_2416,N_1488);
or U8650 (N_8650,N_3755,N_149);
or U8651 (N_8651,N_1619,N_2148);
or U8652 (N_8652,N_369,N_2443);
nor U8653 (N_8653,N_3024,N_2758);
or U8654 (N_8654,N_264,N_4963);
or U8655 (N_8655,N_1657,N_2695);
and U8656 (N_8656,N_776,N_2156);
nand U8657 (N_8657,N_4679,N_4782);
and U8658 (N_8658,N_4989,N_658);
nor U8659 (N_8659,N_3518,N_3113);
and U8660 (N_8660,N_615,N_4831);
nand U8661 (N_8661,N_423,N_717);
nor U8662 (N_8662,N_3357,N_1997);
nor U8663 (N_8663,N_4434,N_4581);
nand U8664 (N_8664,N_2810,N_1124);
nand U8665 (N_8665,N_2619,N_1498);
nand U8666 (N_8666,N_2355,N_1206);
and U8667 (N_8667,N_546,N_735);
nand U8668 (N_8668,N_3107,N_3385);
nor U8669 (N_8669,N_267,N_1813);
or U8670 (N_8670,N_1832,N_4467);
nand U8671 (N_8671,N_413,N_4890);
or U8672 (N_8672,N_824,N_1597);
nor U8673 (N_8673,N_999,N_1979);
or U8674 (N_8674,N_2799,N_3567);
or U8675 (N_8675,N_1577,N_473);
nand U8676 (N_8676,N_1605,N_4522);
nand U8677 (N_8677,N_3515,N_2700);
nor U8678 (N_8678,N_2707,N_3229);
nor U8679 (N_8679,N_1800,N_2520);
nand U8680 (N_8680,N_1254,N_798);
xor U8681 (N_8681,N_275,N_3637);
nand U8682 (N_8682,N_90,N_831);
nand U8683 (N_8683,N_291,N_4326);
and U8684 (N_8684,N_3180,N_2597);
or U8685 (N_8685,N_4446,N_1966);
and U8686 (N_8686,N_4232,N_3133);
nor U8687 (N_8687,N_4828,N_3670);
nor U8688 (N_8688,N_1029,N_983);
nor U8689 (N_8689,N_536,N_1271);
nand U8690 (N_8690,N_4987,N_7);
and U8691 (N_8691,N_1966,N_1893);
nor U8692 (N_8692,N_3109,N_303);
xnor U8693 (N_8693,N_366,N_4003);
nand U8694 (N_8694,N_603,N_2876);
and U8695 (N_8695,N_1850,N_121);
and U8696 (N_8696,N_2802,N_2128);
or U8697 (N_8697,N_642,N_3890);
nand U8698 (N_8698,N_1399,N_3282);
and U8699 (N_8699,N_1289,N_2397);
nand U8700 (N_8700,N_2833,N_3642);
nand U8701 (N_8701,N_3772,N_3722);
or U8702 (N_8702,N_1229,N_483);
nand U8703 (N_8703,N_2531,N_626);
and U8704 (N_8704,N_172,N_4960);
or U8705 (N_8705,N_4657,N_930);
and U8706 (N_8706,N_1037,N_2087);
nor U8707 (N_8707,N_1717,N_271);
nand U8708 (N_8708,N_1164,N_2764);
nor U8709 (N_8709,N_889,N_2527);
or U8710 (N_8710,N_1290,N_664);
nand U8711 (N_8711,N_411,N_1051);
and U8712 (N_8712,N_4444,N_3790);
or U8713 (N_8713,N_4497,N_4652);
or U8714 (N_8714,N_2453,N_3125);
nand U8715 (N_8715,N_1826,N_134);
nor U8716 (N_8716,N_2031,N_1785);
nor U8717 (N_8717,N_4537,N_3534);
nor U8718 (N_8718,N_2936,N_1809);
or U8719 (N_8719,N_1152,N_4271);
and U8720 (N_8720,N_1510,N_2623);
and U8721 (N_8721,N_1129,N_4062);
nand U8722 (N_8722,N_4950,N_4451);
and U8723 (N_8723,N_4364,N_1395);
and U8724 (N_8724,N_2963,N_144);
or U8725 (N_8725,N_3513,N_2549);
nand U8726 (N_8726,N_3891,N_2704);
nand U8727 (N_8727,N_1423,N_3001);
or U8728 (N_8728,N_4525,N_4939);
and U8729 (N_8729,N_3843,N_483);
or U8730 (N_8730,N_46,N_3965);
nand U8731 (N_8731,N_3562,N_1222);
nand U8732 (N_8732,N_919,N_1640);
nor U8733 (N_8733,N_1644,N_4127);
and U8734 (N_8734,N_4916,N_428);
and U8735 (N_8735,N_2922,N_1226);
nor U8736 (N_8736,N_2199,N_1875);
nand U8737 (N_8737,N_2509,N_3200);
nand U8738 (N_8738,N_434,N_1971);
and U8739 (N_8739,N_3904,N_1730);
and U8740 (N_8740,N_2689,N_2050);
nor U8741 (N_8741,N_2638,N_3798);
and U8742 (N_8742,N_853,N_2316);
or U8743 (N_8743,N_3030,N_4340);
nand U8744 (N_8744,N_3421,N_725);
or U8745 (N_8745,N_2558,N_320);
or U8746 (N_8746,N_590,N_1732);
nor U8747 (N_8747,N_2441,N_1473);
nand U8748 (N_8748,N_530,N_39);
nand U8749 (N_8749,N_312,N_2363);
and U8750 (N_8750,N_3446,N_1612);
or U8751 (N_8751,N_4376,N_1548);
or U8752 (N_8752,N_1742,N_560);
or U8753 (N_8753,N_3105,N_388);
nand U8754 (N_8754,N_2099,N_4464);
or U8755 (N_8755,N_2921,N_962);
nor U8756 (N_8756,N_814,N_4897);
nand U8757 (N_8757,N_1982,N_105);
or U8758 (N_8758,N_795,N_4265);
nor U8759 (N_8759,N_3618,N_1140);
and U8760 (N_8760,N_75,N_3699);
and U8761 (N_8761,N_4324,N_2356);
and U8762 (N_8762,N_2527,N_4881);
and U8763 (N_8763,N_3740,N_854);
and U8764 (N_8764,N_2934,N_1535);
and U8765 (N_8765,N_921,N_442);
and U8766 (N_8766,N_1795,N_4004);
nor U8767 (N_8767,N_4842,N_2470);
and U8768 (N_8768,N_415,N_4601);
or U8769 (N_8769,N_4743,N_1829);
or U8770 (N_8770,N_3020,N_1633);
nand U8771 (N_8771,N_3188,N_1192);
and U8772 (N_8772,N_4989,N_285);
nand U8773 (N_8773,N_1784,N_2332);
nor U8774 (N_8774,N_3520,N_3710);
nand U8775 (N_8775,N_3776,N_4619);
xnor U8776 (N_8776,N_2329,N_110);
or U8777 (N_8777,N_2642,N_2967);
or U8778 (N_8778,N_693,N_2015);
nand U8779 (N_8779,N_347,N_3838);
or U8780 (N_8780,N_2558,N_1721);
or U8781 (N_8781,N_1333,N_2700);
and U8782 (N_8782,N_2127,N_1219);
or U8783 (N_8783,N_3589,N_3448);
nor U8784 (N_8784,N_2458,N_2822);
nor U8785 (N_8785,N_152,N_1066);
nor U8786 (N_8786,N_368,N_255);
nand U8787 (N_8787,N_528,N_4202);
nand U8788 (N_8788,N_2777,N_2743);
nand U8789 (N_8789,N_113,N_4392);
nand U8790 (N_8790,N_2069,N_4931);
nand U8791 (N_8791,N_3261,N_3640);
or U8792 (N_8792,N_2981,N_845);
xnor U8793 (N_8793,N_3594,N_2878);
or U8794 (N_8794,N_2520,N_4495);
or U8795 (N_8795,N_595,N_4344);
or U8796 (N_8796,N_4259,N_4576);
and U8797 (N_8797,N_531,N_1501);
and U8798 (N_8798,N_2339,N_2405);
nor U8799 (N_8799,N_3907,N_1230);
nand U8800 (N_8800,N_2271,N_204);
nor U8801 (N_8801,N_121,N_2213);
xor U8802 (N_8802,N_2659,N_1068);
nand U8803 (N_8803,N_2352,N_2573);
nand U8804 (N_8804,N_4672,N_99);
nor U8805 (N_8805,N_2019,N_681);
or U8806 (N_8806,N_3497,N_1010);
or U8807 (N_8807,N_3063,N_639);
or U8808 (N_8808,N_1379,N_2467);
or U8809 (N_8809,N_4753,N_4999);
nor U8810 (N_8810,N_3746,N_1504);
or U8811 (N_8811,N_1437,N_465);
and U8812 (N_8812,N_4275,N_421);
and U8813 (N_8813,N_4020,N_2584);
or U8814 (N_8814,N_4293,N_4821);
and U8815 (N_8815,N_267,N_3016);
or U8816 (N_8816,N_386,N_504);
nor U8817 (N_8817,N_3609,N_4975);
and U8818 (N_8818,N_479,N_32);
and U8819 (N_8819,N_112,N_1306);
nand U8820 (N_8820,N_3516,N_2931);
or U8821 (N_8821,N_1361,N_2829);
or U8822 (N_8822,N_4228,N_3633);
or U8823 (N_8823,N_340,N_4939);
nor U8824 (N_8824,N_3715,N_3334);
nand U8825 (N_8825,N_2342,N_4275);
nor U8826 (N_8826,N_2280,N_4910);
nor U8827 (N_8827,N_3702,N_2816);
or U8828 (N_8828,N_1441,N_2962);
nor U8829 (N_8829,N_831,N_192);
and U8830 (N_8830,N_3198,N_3878);
and U8831 (N_8831,N_467,N_3546);
nor U8832 (N_8832,N_1728,N_3824);
and U8833 (N_8833,N_3998,N_4883);
and U8834 (N_8834,N_2808,N_3264);
and U8835 (N_8835,N_3053,N_1775);
nor U8836 (N_8836,N_3570,N_1417);
nor U8837 (N_8837,N_4307,N_17);
nand U8838 (N_8838,N_2198,N_2323);
nand U8839 (N_8839,N_3354,N_2585);
or U8840 (N_8840,N_553,N_1152);
nand U8841 (N_8841,N_332,N_219);
or U8842 (N_8842,N_236,N_4558);
and U8843 (N_8843,N_2804,N_3709);
nand U8844 (N_8844,N_3887,N_3115);
and U8845 (N_8845,N_603,N_1380);
nand U8846 (N_8846,N_4287,N_1660);
or U8847 (N_8847,N_2459,N_3977);
and U8848 (N_8848,N_787,N_557);
nor U8849 (N_8849,N_2214,N_4056);
and U8850 (N_8850,N_2842,N_2824);
nand U8851 (N_8851,N_4013,N_4262);
nand U8852 (N_8852,N_3100,N_2512);
nor U8853 (N_8853,N_4850,N_3747);
or U8854 (N_8854,N_2506,N_1528);
nor U8855 (N_8855,N_2919,N_596);
xor U8856 (N_8856,N_2686,N_3478);
nor U8857 (N_8857,N_1781,N_4682);
nor U8858 (N_8858,N_3653,N_3897);
nor U8859 (N_8859,N_1888,N_1060);
nand U8860 (N_8860,N_4373,N_2866);
nand U8861 (N_8861,N_3047,N_3070);
or U8862 (N_8862,N_3695,N_1988);
and U8863 (N_8863,N_281,N_2646);
nor U8864 (N_8864,N_456,N_1945);
and U8865 (N_8865,N_1892,N_4488);
and U8866 (N_8866,N_2788,N_159);
nand U8867 (N_8867,N_2555,N_4934);
nor U8868 (N_8868,N_326,N_2186);
nand U8869 (N_8869,N_3480,N_958);
nor U8870 (N_8870,N_3179,N_4386);
nand U8871 (N_8871,N_3577,N_1797);
nor U8872 (N_8872,N_362,N_1810);
nand U8873 (N_8873,N_3914,N_4181);
nand U8874 (N_8874,N_2812,N_4753);
nor U8875 (N_8875,N_3193,N_4372);
or U8876 (N_8876,N_1544,N_1495);
or U8877 (N_8877,N_727,N_4873);
nor U8878 (N_8878,N_462,N_1094);
and U8879 (N_8879,N_3208,N_4246);
or U8880 (N_8880,N_3754,N_320);
nor U8881 (N_8881,N_4666,N_2031);
or U8882 (N_8882,N_2557,N_2750);
nand U8883 (N_8883,N_4310,N_4398);
and U8884 (N_8884,N_3508,N_2561);
and U8885 (N_8885,N_226,N_1826);
nand U8886 (N_8886,N_1658,N_3906);
nand U8887 (N_8887,N_1493,N_3135);
nand U8888 (N_8888,N_404,N_3280);
or U8889 (N_8889,N_3528,N_4261);
and U8890 (N_8890,N_3398,N_2831);
and U8891 (N_8891,N_4239,N_4178);
or U8892 (N_8892,N_3968,N_2898);
nor U8893 (N_8893,N_4386,N_1386);
nor U8894 (N_8894,N_3984,N_602);
and U8895 (N_8895,N_2394,N_1992);
nor U8896 (N_8896,N_4414,N_4189);
or U8897 (N_8897,N_2933,N_1066);
nor U8898 (N_8898,N_622,N_1219);
or U8899 (N_8899,N_667,N_1978);
or U8900 (N_8900,N_2842,N_4315);
or U8901 (N_8901,N_4417,N_664);
nand U8902 (N_8902,N_4617,N_466);
nor U8903 (N_8903,N_475,N_555);
or U8904 (N_8904,N_4806,N_3540);
or U8905 (N_8905,N_3246,N_3795);
or U8906 (N_8906,N_3782,N_1802);
nand U8907 (N_8907,N_3440,N_597);
nor U8908 (N_8908,N_157,N_3995);
nor U8909 (N_8909,N_2922,N_4745);
or U8910 (N_8910,N_2709,N_981);
nor U8911 (N_8911,N_3582,N_3809);
or U8912 (N_8912,N_2789,N_2822);
and U8913 (N_8913,N_4278,N_4086);
nand U8914 (N_8914,N_3864,N_1034);
and U8915 (N_8915,N_2935,N_4359);
nor U8916 (N_8916,N_4275,N_2195);
and U8917 (N_8917,N_584,N_1550);
nand U8918 (N_8918,N_4227,N_1543);
and U8919 (N_8919,N_3834,N_1797);
and U8920 (N_8920,N_2498,N_4153);
and U8921 (N_8921,N_4402,N_3651);
or U8922 (N_8922,N_4019,N_3009);
and U8923 (N_8923,N_1367,N_3836);
nor U8924 (N_8924,N_1703,N_1723);
and U8925 (N_8925,N_236,N_1389);
and U8926 (N_8926,N_1964,N_2814);
and U8927 (N_8927,N_2650,N_2589);
and U8928 (N_8928,N_4605,N_2801);
nor U8929 (N_8929,N_408,N_3008);
nand U8930 (N_8930,N_3279,N_2859);
and U8931 (N_8931,N_2848,N_3593);
nor U8932 (N_8932,N_4817,N_2247);
nand U8933 (N_8933,N_1563,N_2716);
nand U8934 (N_8934,N_120,N_3071);
nor U8935 (N_8935,N_2567,N_1172);
nand U8936 (N_8936,N_2200,N_2844);
and U8937 (N_8937,N_2279,N_765);
nor U8938 (N_8938,N_3989,N_2511);
nand U8939 (N_8939,N_2553,N_3849);
and U8940 (N_8940,N_2981,N_4767);
nor U8941 (N_8941,N_4727,N_1929);
nand U8942 (N_8942,N_4040,N_2546);
or U8943 (N_8943,N_3424,N_372);
nand U8944 (N_8944,N_1537,N_3340);
nor U8945 (N_8945,N_3332,N_3727);
and U8946 (N_8946,N_4336,N_4637);
nand U8947 (N_8947,N_2570,N_2794);
nand U8948 (N_8948,N_4375,N_2182);
or U8949 (N_8949,N_2435,N_573);
and U8950 (N_8950,N_4240,N_2002);
or U8951 (N_8951,N_4444,N_4075);
and U8952 (N_8952,N_738,N_96);
or U8953 (N_8953,N_2411,N_142);
nand U8954 (N_8954,N_595,N_4927);
or U8955 (N_8955,N_465,N_2369);
nor U8956 (N_8956,N_4719,N_1338);
and U8957 (N_8957,N_3971,N_105);
nand U8958 (N_8958,N_2663,N_4586);
nand U8959 (N_8959,N_2825,N_1063);
nand U8960 (N_8960,N_1224,N_326);
nor U8961 (N_8961,N_4654,N_632);
or U8962 (N_8962,N_1831,N_4833);
nand U8963 (N_8963,N_1091,N_4158);
and U8964 (N_8964,N_1752,N_915);
nor U8965 (N_8965,N_4434,N_3225);
nand U8966 (N_8966,N_2634,N_979);
nand U8967 (N_8967,N_1653,N_2174);
or U8968 (N_8968,N_495,N_497);
nand U8969 (N_8969,N_1280,N_2551);
or U8970 (N_8970,N_3717,N_152);
and U8971 (N_8971,N_4032,N_1349);
and U8972 (N_8972,N_1754,N_4461);
nand U8973 (N_8973,N_4183,N_2018);
or U8974 (N_8974,N_1543,N_3329);
nand U8975 (N_8975,N_3696,N_1914);
and U8976 (N_8976,N_3901,N_523);
and U8977 (N_8977,N_2333,N_3995);
nor U8978 (N_8978,N_875,N_2246);
and U8979 (N_8979,N_3178,N_1201);
and U8980 (N_8980,N_2556,N_1511);
nand U8981 (N_8981,N_1569,N_3647);
and U8982 (N_8982,N_2755,N_3001);
nor U8983 (N_8983,N_560,N_3623);
nor U8984 (N_8984,N_3103,N_1098);
nand U8985 (N_8985,N_655,N_652);
nand U8986 (N_8986,N_3560,N_4014);
and U8987 (N_8987,N_3737,N_3952);
and U8988 (N_8988,N_4645,N_1967);
and U8989 (N_8989,N_1105,N_1849);
or U8990 (N_8990,N_2858,N_4591);
nor U8991 (N_8991,N_4874,N_3432);
nand U8992 (N_8992,N_1781,N_2697);
or U8993 (N_8993,N_1813,N_1012);
or U8994 (N_8994,N_1560,N_3241);
or U8995 (N_8995,N_1093,N_1574);
nor U8996 (N_8996,N_4654,N_1599);
and U8997 (N_8997,N_4726,N_3993);
and U8998 (N_8998,N_3795,N_1220);
nand U8999 (N_8999,N_1520,N_2904);
nand U9000 (N_9000,N_1867,N_1960);
nand U9001 (N_9001,N_3734,N_4441);
and U9002 (N_9002,N_4198,N_3103);
xor U9003 (N_9003,N_3217,N_1552);
nand U9004 (N_9004,N_1981,N_1079);
nor U9005 (N_9005,N_4782,N_3035);
nor U9006 (N_9006,N_1003,N_1218);
nand U9007 (N_9007,N_4746,N_40);
or U9008 (N_9008,N_2471,N_1543);
nor U9009 (N_9009,N_4504,N_556);
and U9010 (N_9010,N_2769,N_4747);
nand U9011 (N_9011,N_696,N_722);
and U9012 (N_9012,N_3926,N_2704);
and U9013 (N_9013,N_1514,N_4388);
nand U9014 (N_9014,N_2470,N_3464);
nand U9015 (N_9015,N_4465,N_2882);
and U9016 (N_9016,N_3599,N_3960);
nor U9017 (N_9017,N_461,N_4432);
or U9018 (N_9018,N_1524,N_2437);
or U9019 (N_9019,N_3095,N_4508);
and U9020 (N_9020,N_3212,N_3735);
nor U9021 (N_9021,N_381,N_4797);
and U9022 (N_9022,N_1845,N_1990);
nor U9023 (N_9023,N_1237,N_3769);
nor U9024 (N_9024,N_4601,N_4432);
and U9025 (N_9025,N_707,N_1412);
or U9026 (N_9026,N_3096,N_820);
nand U9027 (N_9027,N_1571,N_1711);
and U9028 (N_9028,N_3073,N_3184);
nand U9029 (N_9029,N_1153,N_3747);
nand U9030 (N_9030,N_2287,N_1645);
and U9031 (N_9031,N_2448,N_142);
nor U9032 (N_9032,N_3327,N_3863);
and U9033 (N_9033,N_814,N_1694);
nand U9034 (N_9034,N_3831,N_3513);
and U9035 (N_9035,N_3122,N_190);
and U9036 (N_9036,N_2745,N_1828);
nor U9037 (N_9037,N_2393,N_4411);
and U9038 (N_9038,N_866,N_323);
nand U9039 (N_9039,N_3028,N_1284);
nand U9040 (N_9040,N_1500,N_4149);
nand U9041 (N_9041,N_4754,N_3195);
or U9042 (N_9042,N_2462,N_1462);
nor U9043 (N_9043,N_44,N_4449);
and U9044 (N_9044,N_2982,N_455);
nor U9045 (N_9045,N_1634,N_3677);
and U9046 (N_9046,N_582,N_4085);
nor U9047 (N_9047,N_2826,N_4012);
nand U9048 (N_9048,N_3796,N_3878);
or U9049 (N_9049,N_949,N_2026);
nor U9050 (N_9050,N_872,N_1261);
nor U9051 (N_9051,N_3558,N_1855);
nor U9052 (N_9052,N_1783,N_1461);
and U9053 (N_9053,N_2107,N_1318);
nor U9054 (N_9054,N_2894,N_1147);
nor U9055 (N_9055,N_4666,N_4252);
nor U9056 (N_9056,N_24,N_4882);
or U9057 (N_9057,N_1201,N_504);
or U9058 (N_9058,N_2740,N_2883);
and U9059 (N_9059,N_3457,N_3996);
nand U9060 (N_9060,N_84,N_4614);
nand U9061 (N_9061,N_2391,N_3583);
and U9062 (N_9062,N_1116,N_3258);
nand U9063 (N_9063,N_1181,N_936);
and U9064 (N_9064,N_4320,N_900);
or U9065 (N_9065,N_752,N_60);
or U9066 (N_9066,N_1929,N_3568);
or U9067 (N_9067,N_3837,N_4904);
nor U9068 (N_9068,N_1690,N_4812);
nor U9069 (N_9069,N_1527,N_2869);
nor U9070 (N_9070,N_1336,N_1155);
nor U9071 (N_9071,N_1550,N_4628);
and U9072 (N_9072,N_3681,N_4819);
nand U9073 (N_9073,N_1418,N_847);
or U9074 (N_9074,N_1832,N_3750);
nand U9075 (N_9075,N_1790,N_3146);
nand U9076 (N_9076,N_178,N_3876);
or U9077 (N_9077,N_1689,N_299);
nand U9078 (N_9078,N_2303,N_314);
nor U9079 (N_9079,N_4411,N_1484);
nand U9080 (N_9080,N_1501,N_3560);
nand U9081 (N_9081,N_4901,N_906);
and U9082 (N_9082,N_2069,N_217);
nor U9083 (N_9083,N_1865,N_3318);
and U9084 (N_9084,N_1765,N_1808);
nand U9085 (N_9085,N_594,N_1180);
and U9086 (N_9086,N_3975,N_4759);
nand U9087 (N_9087,N_3267,N_252);
and U9088 (N_9088,N_1749,N_2766);
and U9089 (N_9089,N_3572,N_77);
nor U9090 (N_9090,N_2081,N_2603);
nor U9091 (N_9091,N_2309,N_4407);
nand U9092 (N_9092,N_3138,N_3140);
nand U9093 (N_9093,N_855,N_2861);
nor U9094 (N_9094,N_2567,N_936);
or U9095 (N_9095,N_4399,N_832);
nand U9096 (N_9096,N_4332,N_2001);
and U9097 (N_9097,N_1547,N_1083);
and U9098 (N_9098,N_2373,N_1105);
or U9099 (N_9099,N_1267,N_1377);
or U9100 (N_9100,N_3665,N_3641);
and U9101 (N_9101,N_3113,N_3079);
or U9102 (N_9102,N_2421,N_2776);
and U9103 (N_9103,N_1914,N_838);
nand U9104 (N_9104,N_1131,N_779);
and U9105 (N_9105,N_595,N_578);
nor U9106 (N_9106,N_571,N_3095);
nand U9107 (N_9107,N_2803,N_965);
or U9108 (N_9108,N_3388,N_4141);
or U9109 (N_9109,N_3728,N_4172);
and U9110 (N_9110,N_4056,N_769);
nor U9111 (N_9111,N_57,N_145);
or U9112 (N_9112,N_4430,N_2675);
and U9113 (N_9113,N_4974,N_2297);
and U9114 (N_9114,N_2746,N_1069);
or U9115 (N_9115,N_3000,N_3124);
and U9116 (N_9116,N_3907,N_2171);
and U9117 (N_9117,N_1177,N_3833);
nor U9118 (N_9118,N_228,N_4671);
nand U9119 (N_9119,N_160,N_4291);
and U9120 (N_9120,N_625,N_2281);
nor U9121 (N_9121,N_2472,N_2352);
or U9122 (N_9122,N_1293,N_3636);
nand U9123 (N_9123,N_3786,N_3106);
and U9124 (N_9124,N_1308,N_420);
and U9125 (N_9125,N_1492,N_4328);
nand U9126 (N_9126,N_958,N_1276);
nand U9127 (N_9127,N_375,N_2625);
and U9128 (N_9128,N_1398,N_2639);
nor U9129 (N_9129,N_3917,N_2887);
nor U9130 (N_9130,N_4585,N_4203);
nand U9131 (N_9131,N_4082,N_2423);
nand U9132 (N_9132,N_3365,N_4562);
or U9133 (N_9133,N_2635,N_4043);
nor U9134 (N_9134,N_4901,N_1559);
nor U9135 (N_9135,N_3549,N_1196);
and U9136 (N_9136,N_2480,N_4689);
or U9137 (N_9137,N_4978,N_636);
xor U9138 (N_9138,N_2,N_169);
or U9139 (N_9139,N_2989,N_2803);
nor U9140 (N_9140,N_11,N_495);
and U9141 (N_9141,N_2082,N_1318);
nand U9142 (N_9142,N_1903,N_1765);
nor U9143 (N_9143,N_597,N_177);
nand U9144 (N_9144,N_1557,N_2738);
nor U9145 (N_9145,N_687,N_2754);
nand U9146 (N_9146,N_3981,N_4718);
and U9147 (N_9147,N_2172,N_354);
nand U9148 (N_9148,N_3595,N_3511);
and U9149 (N_9149,N_3490,N_996);
or U9150 (N_9150,N_3661,N_4189);
and U9151 (N_9151,N_2194,N_838);
nor U9152 (N_9152,N_4171,N_4814);
nand U9153 (N_9153,N_1434,N_3801);
and U9154 (N_9154,N_4714,N_2604);
nor U9155 (N_9155,N_3993,N_477);
or U9156 (N_9156,N_3719,N_4574);
or U9157 (N_9157,N_2346,N_3811);
nand U9158 (N_9158,N_4910,N_1173);
nor U9159 (N_9159,N_55,N_1279);
and U9160 (N_9160,N_3471,N_3348);
nand U9161 (N_9161,N_4927,N_1515);
and U9162 (N_9162,N_4310,N_4328);
or U9163 (N_9163,N_987,N_2287);
or U9164 (N_9164,N_356,N_2845);
nor U9165 (N_9165,N_4020,N_943);
nand U9166 (N_9166,N_4274,N_1213);
or U9167 (N_9167,N_3489,N_4132);
or U9168 (N_9168,N_2158,N_170);
nor U9169 (N_9169,N_1008,N_3493);
or U9170 (N_9170,N_2623,N_2574);
or U9171 (N_9171,N_881,N_4506);
and U9172 (N_9172,N_3853,N_2600);
nand U9173 (N_9173,N_2885,N_3897);
or U9174 (N_9174,N_2578,N_3065);
nand U9175 (N_9175,N_1356,N_2294);
nand U9176 (N_9176,N_2,N_3984);
nand U9177 (N_9177,N_2998,N_1319);
or U9178 (N_9178,N_742,N_1512);
nor U9179 (N_9179,N_1387,N_4067);
xnor U9180 (N_9180,N_827,N_3547);
nand U9181 (N_9181,N_4890,N_4525);
and U9182 (N_9182,N_4314,N_4194);
nand U9183 (N_9183,N_3183,N_833);
or U9184 (N_9184,N_2720,N_2814);
or U9185 (N_9185,N_4797,N_3082);
nand U9186 (N_9186,N_4630,N_4617);
or U9187 (N_9187,N_4968,N_2500);
and U9188 (N_9188,N_4448,N_4037);
nor U9189 (N_9189,N_891,N_2570);
xor U9190 (N_9190,N_93,N_4582);
nor U9191 (N_9191,N_1289,N_3546);
or U9192 (N_9192,N_1681,N_1348);
nor U9193 (N_9193,N_1235,N_18);
nand U9194 (N_9194,N_2439,N_799);
nor U9195 (N_9195,N_834,N_1357);
and U9196 (N_9196,N_4040,N_4881);
and U9197 (N_9197,N_4671,N_343);
nand U9198 (N_9198,N_1862,N_66);
nand U9199 (N_9199,N_452,N_3955);
nor U9200 (N_9200,N_4032,N_4484);
or U9201 (N_9201,N_3836,N_2459);
or U9202 (N_9202,N_4880,N_306);
nor U9203 (N_9203,N_2127,N_3813);
nand U9204 (N_9204,N_2823,N_2213);
nand U9205 (N_9205,N_1230,N_4460);
and U9206 (N_9206,N_1350,N_1432);
nand U9207 (N_9207,N_3046,N_2966);
nor U9208 (N_9208,N_2386,N_776);
and U9209 (N_9209,N_4401,N_631);
and U9210 (N_9210,N_487,N_1594);
and U9211 (N_9211,N_2832,N_1441);
or U9212 (N_9212,N_4751,N_3793);
or U9213 (N_9213,N_626,N_962);
nand U9214 (N_9214,N_4644,N_456);
nor U9215 (N_9215,N_3601,N_1036);
nor U9216 (N_9216,N_3917,N_2684);
nor U9217 (N_9217,N_1402,N_3188);
nor U9218 (N_9218,N_880,N_1433);
nor U9219 (N_9219,N_772,N_3016);
nor U9220 (N_9220,N_2834,N_850);
nor U9221 (N_9221,N_2854,N_4291);
or U9222 (N_9222,N_3157,N_2654);
nor U9223 (N_9223,N_328,N_2144);
nor U9224 (N_9224,N_3560,N_719);
and U9225 (N_9225,N_3705,N_99);
xor U9226 (N_9226,N_3388,N_568);
nand U9227 (N_9227,N_3019,N_4626);
or U9228 (N_9228,N_477,N_501);
nor U9229 (N_9229,N_2174,N_257);
nand U9230 (N_9230,N_4215,N_734);
nand U9231 (N_9231,N_2325,N_2827);
or U9232 (N_9232,N_3031,N_1717);
nand U9233 (N_9233,N_3256,N_3656);
or U9234 (N_9234,N_3542,N_2799);
nor U9235 (N_9235,N_4070,N_4335);
nor U9236 (N_9236,N_2491,N_2057);
or U9237 (N_9237,N_1019,N_2984);
nand U9238 (N_9238,N_985,N_2836);
or U9239 (N_9239,N_2725,N_849);
nand U9240 (N_9240,N_2204,N_4663);
or U9241 (N_9241,N_4569,N_3377);
nor U9242 (N_9242,N_2918,N_286);
and U9243 (N_9243,N_4432,N_2142);
nor U9244 (N_9244,N_3242,N_3872);
or U9245 (N_9245,N_3775,N_130);
or U9246 (N_9246,N_882,N_2468);
and U9247 (N_9247,N_3486,N_4038);
nor U9248 (N_9248,N_1709,N_3109);
nor U9249 (N_9249,N_3526,N_2424);
nand U9250 (N_9250,N_4556,N_3308);
and U9251 (N_9251,N_3972,N_3757);
xnor U9252 (N_9252,N_479,N_1602);
nand U9253 (N_9253,N_3661,N_3185);
or U9254 (N_9254,N_449,N_2891);
and U9255 (N_9255,N_1355,N_2444);
nand U9256 (N_9256,N_4228,N_156);
and U9257 (N_9257,N_887,N_507);
nand U9258 (N_9258,N_4400,N_4183);
nand U9259 (N_9259,N_4113,N_2572);
nor U9260 (N_9260,N_1212,N_810);
nor U9261 (N_9261,N_4075,N_674);
nor U9262 (N_9262,N_1054,N_4987);
or U9263 (N_9263,N_1155,N_2919);
or U9264 (N_9264,N_4542,N_3848);
nand U9265 (N_9265,N_4749,N_1288);
nor U9266 (N_9266,N_3288,N_4089);
nand U9267 (N_9267,N_4415,N_3466);
nor U9268 (N_9268,N_4360,N_1200);
and U9269 (N_9269,N_4410,N_4448);
and U9270 (N_9270,N_2795,N_3168);
nand U9271 (N_9271,N_2213,N_1328);
and U9272 (N_9272,N_1675,N_2317);
and U9273 (N_9273,N_2314,N_1752);
or U9274 (N_9274,N_533,N_4798);
nand U9275 (N_9275,N_1355,N_314);
or U9276 (N_9276,N_1008,N_2540);
xor U9277 (N_9277,N_137,N_4820);
and U9278 (N_9278,N_3264,N_1992);
and U9279 (N_9279,N_3745,N_1542);
or U9280 (N_9280,N_2926,N_3436);
nand U9281 (N_9281,N_154,N_445);
and U9282 (N_9282,N_2539,N_4893);
nand U9283 (N_9283,N_2474,N_2987);
nand U9284 (N_9284,N_3132,N_3997);
or U9285 (N_9285,N_3372,N_1626);
nor U9286 (N_9286,N_4142,N_1578);
nor U9287 (N_9287,N_12,N_2411);
and U9288 (N_9288,N_203,N_3985);
nand U9289 (N_9289,N_479,N_3163);
nor U9290 (N_9290,N_1262,N_4556);
or U9291 (N_9291,N_780,N_2913);
and U9292 (N_9292,N_2830,N_386);
nand U9293 (N_9293,N_728,N_2909);
nand U9294 (N_9294,N_703,N_4548);
or U9295 (N_9295,N_948,N_1938);
or U9296 (N_9296,N_2263,N_1562);
nand U9297 (N_9297,N_2356,N_1590);
nor U9298 (N_9298,N_4474,N_145);
nor U9299 (N_9299,N_3451,N_227);
and U9300 (N_9300,N_2315,N_4677);
nand U9301 (N_9301,N_4460,N_2706);
or U9302 (N_9302,N_671,N_4531);
or U9303 (N_9303,N_315,N_1250);
nand U9304 (N_9304,N_4137,N_640);
and U9305 (N_9305,N_4653,N_4442);
or U9306 (N_9306,N_3011,N_1107);
and U9307 (N_9307,N_4783,N_512);
or U9308 (N_9308,N_1234,N_1681);
nor U9309 (N_9309,N_3559,N_2708);
nand U9310 (N_9310,N_570,N_1799);
nand U9311 (N_9311,N_3027,N_1347);
nand U9312 (N_9312,N_1625,N_2631);
or U9313 (N_9313,N_1469,N_4928);
nor U9314 (N_9314,N_445,N_771);
nor U9315 (N_9315,N_3376,N_1100);
nand U9316 (N_9316,N_3291,N_3835);
and U9317 (N_9317,N_1796,N_332);
and U9318 (N_9318,N_4439,N_3907);
nand U9319 (N_9319,N_1256,N_4744);
nand U9320 (N_9320,N_3545,N_4266);
nor U9321 (N_9321,N_2038,N_3835);
or U9322 (N_9322,N_433,N_2987);
or U9323 (N_9323,N_1333,N_3470);
nor U9324 (N_9324,N_3449,N_725);
and U9325 (N_9325,N_1485,N_3754);
nor U9326 (N_9326,N_3910,N_381);
nor U9327 (N_9327,N_4107,N_4066);
nor U9328 (N_9328,N_3047,N_3256);
nand U9329 (N_9329,N_4184,N_858);
or U9330 (N_9330,N_636,N_3500);
and U9331 (N_9331,N_3897,N_3995);
or U9332 (N_9332,N_2101,N_1144);
nand U9333 (N_9333,N_3929,N_3204);
nor U9334 (N_9334,N_4604,N_3590);
xnor U9335 (N_9335,N_2903,N_143);
nand U9336 (N_9336,N_2557,N_2623);
nor U9337 (N_9337,N_3283,N_3661);
nand U9338 (N_9338,N_3440,N_510);
and U9339 (N_9339,N_1879,N_2958);
and U9340 (N_9340,N_2879,N_4573);
and U9341 (N_9341,N_1921,N_663);
nor U9342 (N_9342,N_3082,N_3436);
and U9343 (N_9343,N_4412,N_587);
nor U9344 (N_9344,N_1031,N_1123);
or U9345 (N_9345,N_4995,N_1296);
nor U9346 (N_9346,N_1119,N_3925);
nor U9347 (N_9347,N_199,N_4121);
nor U9348 (N_9348,N_2433,N_4869);
nand U9349 (N_9349,N_1120,N_1586);
or U9350 (N_9350,N_1307,N_4671);
or U9351 (N_9351,N_223,N_1857);
or U9352 (N_9352,N_923,N_4065);
nor U9353 (N_9353,N_3326,N_1682);
or U9354 (N_9354,N_633,N_19);
nand U9355 (N_9355,N_1564,N_3703);
or U9356 (N_9356,N_4300,N_3762);
and U9357 (N_9357,N_1057,N_718);
nor U9358 (N_9358,N_165,N_1439);
and U9359 (N_9359,N_3357,N_2150);
or U9360 (N_9360,N_2164,N_3551);
and U9361 (N_9361,N_3622,N_1180);
or U9362 (N_9362,N_4712,N_3415);
and U9363 (N_9363,N_1556,N_3012);
nand U9364 (N_9364,N_2393,N_4180);
nor U9365 (N_9365,N_3028,N_1799);
and U9366 (N_9366,N_3810,N_3563);
nand U9367 (N_9367,N_350,N_4177);
and U9368 (N_9368,N_2975,N_2509);
nor U9369 (N_9369,N_2368,N_1192);
or U9370 (N_9370,N_4799,N_3710);
and U9371 (N_9371,N_2692,N_496);
nor U9372 (N_9372,N_2372,N_3174);
or U9373 (N_9373,N_1299,N_4292);
nor U9374 (N_9374,N_1856,N_811);
and U9375 (N_9375,N_3020,N_4934);
or U9376 (N_9376,N_2220,N_4549);
nand U9377 (N_9377,N_992,N_708);
and U9378 (N_9378,N_1096,N_4986);
and U9379 (N_9379,N_4020,N_951);
nor U9380 (N_9380,N_1738,N_3387);
nor U9381 (N_9381,N_3166,N_2739);
nor U9382 (N_9382,N_4115,N_1355);
nand U9383 (N_9383,N_3855,N_1202);
and U9384 (N_9384,N_3015,N_1403);
nand U9385 (N_9385,N_256,N_841);
or U9386 (N_9386,N_4688,N_1934);
and U9387 (N_9387,N_40,N_1494);
or U9388 (N_9388,N_2004,N_1328);
or U9389 (N_9389,N_2781,N_3531);
or U9390 (N_9390,N_2744,N_4196);
nand U9391 (N_9391,N_4573,N_1279);
or U9392 (N_9392,N_268,N_3603);
and U9393 (N_9393,N_3118,N_1675);
or U9394 (N_9394,N_628,N_4044);
or U9395 (N_9395,N_828,N_3615);
and U9396 (N_9396,N_3955,N_823);
and U9397 (N_9397,N_4304,N_3244);
nor U9398 (N_9398,N_3570,N_623);
or U9399 (N_9399,N_2426,N_3126);
nor U9400 (N_9400,N_2588,N_4998);
nand U9401 (N_9401,N_4163,N_266);
or U9402 (N_9402,N_4204,N_1999);
nand U9403 (N_9403,N_1796,N_4966);
nor U9404 (N_9404,N_2470,N_4963);
or U9405 (N_9405,N_475,N_1060);
or U9406 (N_9406,N_1905,N_513);
or U9407 (N_9407,N_3489,N_4834);
or U9408 (N_9408,N_3412,N_1159);
and U9409 (N_9409,N_4569,N_4643);
and U9410 (N_9410,N_1586,N_2102);
nor U9411 (N_9411,N_742,N_4247);
or U9412 (N_9412,N_2667,N_1506);
nand U9413 (N_9413,N_4386,N_1819);
or U9414 (N_9414,N_3815,N_4856);
and U9415 (N_9415,N_4738,N_4700);
nor U9416 (N_9416,N_1275,N_2325);
or U9417 (N_9417,N_587,N_2923);
or U9418 (N_9418,N_514,N_2468);
and U9419 (N_9419,N_1604,N_3167);
nand U9420 (N_9420,N_4054,N_3014);
or U9421 (N_9421,N_4852,N_1549);
or U9422 (N_9422,N_1843,N_3062);
nor U9423 (N_9423,N_4336,N_1108);
and U9424 (N_9424,N_4462,N_1500);
and U9425 (N_9425,N_2902,N_2458);
or U9426 (N_9426,N_2295,N_3841);
nand U9427 (N_9427,N_2418,N_3217);
nor U9428 (N_9428,N_1967,N_3496);
nor U9429 (N_9429,N_1956,N_1261);
and U9430 (N_9430,N_3647,N_2157);
and U9431 (N_9431,N_4030,N_1967);
and U9432 (N_9432,N_4807,N_2386);
nor U9433 (N_9433,N_2878,N_4424);
nand U9434 (N_9434,N_935,N_3148);
or U9435 (N_9435,N_4257,N_4956);
or U9436 (N_9436,N_3285,N_4145);
or U9437 (N_9437,N_4237,N_3644);
nor U9438 (N_9438,N_1392,N_2590);
and U9439 (N_9439,N_3384,N_592);
nand U9440 (N_9440,N_1190,N_669);
and U9441 (N_9441,N_4144,N_3891);
nand U9442 (N_9442,N_4582,N_3463);
nand U9443 (N_9443,N_4978,N_4942);
or U9444 (N_9444,N_2139,N_4298);
or U9445 (N_9445,N_4125,N_1426);
and U9446 (N_9446,N_4608,N_958);
nor U9447 (N_9447,N_2508,N_2269);
nand U9448 (N_9448,N_3267,N_1819);
nand U9449 (N_9449,N_4874,N_3854);
nand U9450 (N_9450,N_3133,N_2541);
or U9451 (N_9451,N_4714,N_3791);
nand U9452 (N_9452,N_4490,N_3537);
nor U9453 (N_9453,N_4386,N_2500);
nand U9454 (N_9454,N_3898,N_2455);
nor U9455 (N_9455,N_3069,N_1768);
nand U9456 (N_9456,N_4336,N_2487);
and U9457 (N_9457,N_1268,N_4239);
and U9458 (N_9458,N_3334,N_467);
nand U9459 (N_9459,N_3944,N_1585);
or U9460 (N_9460,N_2377,N_3128);
nor U9461 (N_9461,N_4502,N_1131);
or U9462 (N_9462,N_3330,N_2100);
nor U9463 (N_9463,N_3732,N_3256);
nor U9464 (N_9464,N_2568,N_1692);
xnor U9465 (N_9465,N_4062,N_304);
or U9466 (N_9466,N_4333,N_4425);
nand U9467 (N_9467,N_4635,N_119);
and U9468 (N_9468,N_4060,N_543);
and U9469 (N_9469,N_2256,N_4384);
nor U9470 (N_9470,N_2730,N_4883);
and U9471 (N_9471,N_1464,N_3448);
nor U9472 (N_9472,N_2397,N_682);
or U9473 (N_9473,N_1671,N_3323);
and U9474 (N_9474,N_3282,N_1326);
or U9475 (N_9475,N_1341,N_1195);
nor U9476 (N_9476,N_4769,N_3951);
or U9477 (N_9477,N_3178,N_181);
or U9478 (N_9478,N_2388,N_468);
nor U9479 (N_9479,N_577,N_4889);
nand U9480 (N_9480,N_3851,N_1919);
or U9481 (N_9481,N_1479,N_309);
and U9482 (N_9482,N_786,N_3115);
nand U9483 (N_9483,N_2180,N_3912);
or U9484 (N_9484,N_4744,N_3274);
nor U9485 (N_9485,N_4721,N_589);
and U9486 (N_9486,N_4427,N_4052);
nand U9487 (N_9487,N_4114,N_2577);
nand U9488 (N_9488,N_985,N_2397);
nand U9489 (N_9489,N_671,N_233);
nand U9490 (N_9490,N_3565,N_86);
nor U9491 (N_9491,N_1825,N_2372);
or U9492 (N_9492,N_2102,N_4188);
nor U9493 (N_9493,N_2699,N_3829);
or U9494 (N_9494,N_2833,N_4355);
or U9495 (N_9495,N_3376,N_1610);
or U9496 (N_9496,N_3724,N_2446);
xnor U9497 (N_9497,N_1663,N_4614);
nor U9498 (N_9498,N_1246,N_44);
or U9499 (N_9499,N_4709,N_4571);
and U9500 (N_9500,N_4032,N_3201);
nor U9501 (N_9501,N_1706,N_3922);
or U9502 (N_9502,N_424,N_2464);
and U9503 (N_9503,N_1204,N_2415);
or U9504 (N_9504,N_2673,N_859);
nand U9505 (N_9505,N_990,N_2104);
or U9506 (N_9506,N_2490,N_1493);
or U9507 (N_9507,N_2248,N_2347);
nand U9508 (N_9508,N_3226,N_2480);
nand U9509 (N_9509,N_2865,N_4592);
or U9510 (N_9510,N_3382,N_1859);
nor U9511 (N_9511,N_3486,N_3602);
or U9512 (N_9512,N_74,N_140);
nand U9513 (N_9513,N_1818,N_2719);
nor U9514 (N_9514,N_1956,N_4020);
and U9515 (N_9515,N_859,N_2808);
or U9516 (N_9516,N_4980,N_4267);
nor U9517 (N_9517,N_194,N_1855);
and U9518 (N_9518,N_2790,N_3654);
nor U9519 (N_9519,N_4939,N_114);
or U9520 (N_9520,N_1403,N_2397);
nand U9521 (N_9521,N_4180,N_3041);
nand U9522 (N_9522,N_1175,N_1892);
and U9523 (N_9523,N_3106,N_734);
and U9524 (N_9524,N_756,N_4534);
nor U9525 (N_9525,N_3711,N_4456);
nor U9526 (N_9526,N_1002,N_2236);
or U9527 (N_9527,N_3820,N_3453);
nor U9528 (N_9528,N_4150,N_3888);
nor U9529 (N_9529,N_4485,N_4549);
nor U9530 (N_9530,N_3588,N_1086);
and U9531 (N_9531,N_1980,N_4965);
nand U9532 (N_9532,N_1682,N_910);
and U9533 (N_9533,N_2453,N_4266);
and U9534 (N_9534,N_1163,N_4801);
nand U9535 (N_9535,N_4468,N_1459);
nor U9536 (N_9536,N_4285,N_1169);
nor U9537 (N_9537,N_2145,N_4000);
or U9538 (N_9538,N_3774,N_1820);
or U9539 (N_9539,N_1926,N_1477);
and U9540 (N_9540,N_4656,N_807);
nor U9541 (N_9541,N_3142,N_2631);
and U9542 (N_9542,N_2473,N_4132);
nand U9543 (N_9543,N_1682,N_1999);
or U9544 (N_9544,N_4362,N_431);
or U9545 (N_9545,N_3178,N_4383);
nor U9546 (N_9546,N_4163,N_3229);
nor U9547 (N_9547,N_4705,N_322);
nand U9548 (N_9548,N_4578,N_1942);
nor U9549 (N_9549,N_3378,N_3169);
or U9550 (N_9550,N_293,N_102);
and U9551 (N_9551,N_993,N_2977);
or U9552 (N_9552,N_4685,N_3244);
nor U9553 (N_9553,N_2379,N_4764);
nand U9554 (N_9554,N_4033,N_4480);
nor U9555 (N_9555,N_4221,N_3736);
xor U9556 (N_9556,N_2706,N_350);
and U9557 (N_9557,N_2149,N_936);
and U9558 (N_9558,N_773,N_4407);
nor U9559 (N_9559,N_2835,N_3415);
or U9560 (N_9560,N_3017,N_1379);
and U9561 (N_9561,N_2519,N_2912);
nand U9562 (N_9562,N_928,N_1340);
or U9563 (N_9563,N_4078,N_2124);
nor U9564 (N_9564,N_3403,N_37);
and U9565 (N_9565,N_2547,N_1733);
nand U9566 (N_9566,N_333,N_2344);
nand U9567 (N_9567,N_4155,N_3652);
and U9568 (N_9568,N_2000,N_2512);
and U9569 (N_9569,N_1594,N_3941);
and U9570 (N_9570,N_3433,N_2143);
and U9571 (N_9571,N_2817,N_1144);
nand U9572 (N_9572,N_2352,N_1860);
nor U9573 (N_9573,N_1955,N_2004);
or U9574 (N_9574,N_3136,N_1481);
nand U9575 (N_9575,N_4658,N_1049);
nor U9576 (N_9576,N_3259,N_721);
nor U9577 (N_9577,N_97,N_1981);
and U9578 (N_9578,N_3539,N_3409);
and U9579 (N_9579,N_2227,N_1873);
and U9580 (N_9580,N_4870,N_2183);
xnor U9581 (N_9581,N_419,N_3296);
nor U9582 (N_9582,N_3546,N_3403);
nor U9583 (N_9583,N_3344,N_2872);
xor U9584 (N_9584,N_1765,N_579);
nand U9585 (N_9585,N_2707,N_3589);
or U9586 (N_9586,N_2244,N_996);
nand U9587 (N_9587,N_1317,N_3321);
or U9588 (N_9588,N_2531,N_572);
nand U9589 (N_9589,N_1872,N_4213);
nand U9590 (N_9590,N_3931,N_4632);
nand U9591 (N_9591,N_647,N_1576);
or U9592 (N_9592,N_4791,N_4752);
or U9593 (N_9593,N_2221,N_246);
and U9594 (N_9594,N_924,N_2140);
or U9595 (N_9595,N_2177,N_268);
or U9596 (N_9596,N_4499,N_3533);
nor U9597 (N_9597,N_938,N_746);
nand U9598 (N_9598,N_3187,N_1901);
nand U9599 (N_9599,N_4547,N_4909);
or U9600 (N_9600,N_2128,N_498);
and U9601 (N_9601,N_934,N_2913);
nand U9602 (N_9602,N_3848,N_1080);
nand U9603 (N_9603,N_3464,N_4522);
and U9604 (N_9604,N_809,N_4829);
or U9605 (N_9605,N_3642,N_1138);
or U9606 (N_9606,N_226,N_1239);
nor U9607 (N_9607,N_3094,N_111);
nor U9608 (N_9608,N_2526,N_4445);
or U9609 (N_9609,N_3336,N_909);
nor U9610 (N_9610,N_2000,N_1366);
nor U9611 (N_9611,N_1167,N_3699);
and U9612 (N_9612,N_1358,N_4796);
and U9613 (N_9613,N_4619,N_4573);
nor U9614 (N_9614,N_1859,N_4408);
or U9615 (N_9615,N_2387,N_1849);
or U9616 (N_9616,N_774,N_1802);
nor U9617 (N_9617,N_2877,N_3284);
nand U9618 (N_9618,N_2622,N_1838);
or U9619 (N_9619,N_2842,N_3502);
nor U9620 (N_9620,N_1535,N_2153);
nand U9621 (N_9621,N_275,N_2680);
or U9622 (N_9622,N_4767,N_2939);
and U9623 (N_9623,N_816,N_2518);
and U9624 (N_9624,N_4368,N_390);
nand U9625 (N_9625,N_421,N_2386);
nand U9626 (N_9626,N_4283,N_580);
nor U9627 (N_9627,N_2572,N_3350);
nor U9628 (N_9628,N_706,N_1440);
or U9629 (N_9629,N_348,N_2855);
or U9630 (N_9630,N_1149,N_2604);
and U9631 (N_9631,N_3298,N_3770);
or U9632 (N_9632,N_2839,N_2810);
nand U9633 (N_9633,N_3642,N_692);
or U9634 (N_9634,N_3711,N_1780);
and U9635 (N_9635,N_2962,N_3993);
nor U9636 (N_9636,N_723,N_550);
nor U9637 (N_9637,N_1349,N_2982);
or U9638 (N_9638,N_4228,N_2848);
or U9639 (N_9639,N_2860,N_3095);
and U9640 (N_9640,N_3624,N_1882);
nor U9641 (N_9641,N_895,N_3735);
and U9642 (N_9642,N_1826,N_3001);
or U9643 (N_9643,N_4276,N_4680);
nand U9644 (N_9644,N_3901,N_3355);
nand U9645 (N_9645,N_899,N_716);
nor U9646 (N_9646,N_3453,N_356);
and U9647 (N_9647,N_2372,N_267);
and U9648 (N_9648,N_917,N_4789);
nand U9649 (N_9649,N_4950,N_1404);
or U9650 (N_9650,N_4096,N_1525);
nand U9651 (N_9651,N_1565,N_1650);
and U9652 (N_9652,N_3492,N_4589);
nor U9653 (N_9653,N_3021,N_2019);
nor U9654 (N_9654,N_936,N_3860);
and U9655 (N_9655,N_1697,N_3218);
or U9656 (N_9656,N_4159,N_4395);
nor U9657 (N_9657,N_1981,N_1912);
and U9658 (N_9658,N_1954,N_922);
and U9659 (N_9659,N_2296,N_2117);
and U9660 (N_9660,N_2788,N_132);
nor U9661 (N_9661,N_595,N_4403);
nand U9662 (N_9662,N_546,N_181);
or U9663 (N_9663,N_1944,N_3101);
nor U9664 (N_9664,N_3040,N_1382);
or U9665 (N_9665,N_1188,N_1935);
or U9666 (N_9666,N_2541,N_4841);
or U9667 (N_9667,N_3691,N_654);
nand U9668 (N_9668,N_1146,N_900);
nand U9669 (N_9669,N_3500,N_316);
or U9670 (N_9670,N_4960,N_522);
or U9671 (N_9671,N_1731,N_4039);
or U9672 (N_9672,N_3006,N_2905);
and U9673 (N_9673,N_324,N_667);
nor U9674 (N_9674,N_281,N_2580);
or U9675 (N_9675,N_3998,N_869);
or U9676 (N_9676,N_4184,N_2448);
or U9677 (N_9677,N_756,N_3599);
and U9678 (N_9678,N_4136,N_2790);
nand U9679 (N_9679,N_1002,N_3119);
nand U9680 (N_9680,N_4397,N_4974);
or U9681 (N_9681,N_395,N_3927);
nand U9682 (N_9682,N_2716,N_2147);
or U9683 (N_9683,N_453,N_412);
or U9684 (N_9684,N_477,N_3249);
or U9685 (N_9685,N_936,N_2044);
nor U9686 (N_9686,N_4220,N_2032);
and U9687 (N_9687,N_3326,N_3489);
nand U9688 (N_9688,N_171,N_1613);
or U9689 (N_9689,N_932,N_160);
nand U9690 (N_9690,N_191,N_4420);
xnor U9691 (N_9691,N_539,N_4933);
nand U9692 (N_9692,N_2502,N_1440);
and U9693 (N_9693,N_4382,N_1753);
and U9694 (N_9694,N_686,N_3568);
or U9695 (N_9695,N_1266,N_2075);
or U9696 (N_9696,N_3598,N_1317);
and U9697 (N_9697,N_2237,N_2742);
and U9698 (N_9698,N_4573,N_1181);
or U9699 (N_9699,N_2711,N_3471);
or U9700 (N_9700,N_658,N_4549);
and U9701 (N_9701,N_3873,N_1479);
or U9702 (N_9702,N_3941,N_575);
or U9703 (N_9703,N_1840,N_2353);
nand U9704 (N_9704,N_334,N_4213);
nor U9705 (N_9705,N_4078,N_1627);
and U9706 (N_9706,N_3124,N_4366);
nand U9707 (N_9707,N_2979,N_4400);
nand U9708 (N_9708,N_3561,N_1740);
or U9709 (N_9709,N_2008,N_4925);
and U9710 (N_9710,N_3071,N_2475);
nor U9711 (N_9711,N_4630,N_4806);
or U9712 (N_9712,N_4225,N_1319);
nand U9713 (N_9713,N_4217,N_1030);
and U9714 (N_9714,N_4581,N_1007);
nor U9715 (N_9715,N_2860,N_1751);
and U9716 (N_9716,N_3156,N_4633);
or U9717 (N_9717,N_3898,N_4951);
nand U9718 (N_9718,N_4814,N_2974);
nand U9719 (N_9719,N_3425,N_3122);
or U9720 (N_9720,N_4808,N_2602);
and U9721 (N_9721,N_4407,N_4274);
nand U9722 (N_9722,N_2960,N_961);
and U9723 (N_9723,N_3246,N_1091);
nand U9724 (N_9724,N_1569,N_4821);
or U9725 (N_9725,N_2272,N_2345);
nand U9726 (N_9726,N_1468,N_906);
nor U9727 (N_9727,N_660,N_4339);
or U9728 (N_9728,N_500,N_4207);
nand U9729 (N_9729,N_246,N_3964);
or U9730 (N_9730,N_1546,N_2071);
nand U9731 (N_9731,N_2107,N_2850);
or U9732 (N_9732,N_594,N_3058);
or U9733 (N_9733,N_1198,N_3981);
and U9734 (N_9734,N_4456,N_1635);
nand U9735 (N_9735,N_209,N_104);
or U9736 (N_9736,N_3491,N_256);
or U9737 (N_9737,N_1032,N_561);
nor U9738 (N_9738,N_313,N_3077);
nor U9739 (N_9739,N_2886,N_1848);
nand U9740 (N_9740,N_2052,N_1053);
nor U9741 (N_9741,N_1369,N_2315);
nor U9742 (N_9742,N_3874,N_184);
or U9743 (N_9743,N_4155,N_4694);
nor U9744 (N_9744,N_3305,N_138);
nand U9745 (N_9745,N_1095,N_4390);
nor U9746 (N_9746,N_2924,N_1260);
or U9747 (N_9747,N_1346,N_1409);
nand U9748 (N_9748,N_1124,N_3411);
nor U9749 (N_9749,N_4576,N_1000);
nand U9750 (N_9750,N_1489,N_1251);
and U9751 (N_9751,N_3596,N_4558);
and U9752 (N_9752,N_4900,N_3532);
nand U9753 (N_9753,N_1079,N_3790);
or U9754 (N_9754,N_675,N_3229);
nand U9755 (N_9755,N_143,N_232);
and U9756 (N_9756,N_2754,N_3934);
and U9757 (N_9757,N_4669,N_2459);
nand U9758 (N_9758,N_1312,N_4945);
nand U9759 (N_9759,N_1721,N_1308);
nor U9760 (N_9760,N_4027,N_1336);
nand U9761 (N_9761,N_4960,N_4276);
nor U9762 (N_9762,N_1512,N_431);
and U9763 (N_9763,N_990,N_2540);
nor U9764 (N_9764,N_4133,N_4045);
nor U9765 (N_9765,N_377,N_4394);
or U9766 (N_9766,N_4291,N_4419);
nor U9767 (N_9767,N_2521,N_1720);
and U9768 (N_9768,N_1287,N_205);
and U9769 (N_9769,N_2741,N_1659);
or U9770 (N_9770,N_435,N_1744);
nor U9771 (N_9771,N_1458,N_4035);
nor U9772 (N_9772,N_1884,N_1671);
and U9773 (N_9773,N_1195,N_4756);
and U9774 (N_9774,N_2124,N_3041);
nand U9775 (N_9775,N_1337,N_4808);
or U9776 (N_9776,N_525,N_3763);
or U9777 (N_9777,N_749,N_1656);
and U9778 (N_9778,N_3097,N_4572);
or U9779 (N_9779,N_2784,N_2762);
nor U9780 (N_9780,N_4270,N_1588);
nor U9781 (N_9781,N_1711,N_3442);
nor U9782 (N_9782,N_948,N_1003);
nand U9783 (N_9783,N_1848,N_1983);
nand U9784 (N_9784,N_1254,N_1040);
nand U9785 (N_9785,N_4960,N_1922);
and U9786 (N_9786,N_3941,N_4620);
or U9787 (N_9787,N_1019,N_223);
nand U9788 (N_9788,N_3783,N_2985);
or U9789 (N_9789,N_3611,N_4298);
or U9790 (N_9790,N_749,N_1262);
nor U9791 (N_9791,N_1873,N_3220);
and U9792 (N_9792,N_3481,N_172);
nor U9793 (N_9793,N_2482,N_3132);
and U9794 (N_9794,N_2793,N_3167);
or U9795 (N_9795,N_1673,N_2521);
nand U9796 (N_9796,N_4942,N_187);
nand U9797 (N_9797,N_1283,N_4603);
or U9798 (N_9798,N_2511,N_1895);
nand U9799 (N_9799,N_4311,N_9);
nand U9800 (N_9800,N_57,N_2313);
nand U9801 (N_9801,N_3915,N_4009);
nor U9802 (N_9802,N_4968,N_2534);
nand U9803 (N_9803,N_4890,N_3243);
nor U9804 (N_9804,N_4519,N_4650);
or U9805 (N_9805,N_3931,N_1743);
and U9806 (N_9806,N_1525,N_2256);
nand U9807 (N_9807,N_4714,N_2561);
nor U9808 (N_9808,N_1960,N_154);
nor U9809 (N_9809,N_2991,N_4322);
nor U9810 (N_9810,N_3,N_1225);
nand U9811 (N_9811,N_1356,N_2587);
or U9812 (N_9812,N_3638,N_1453);
nand U9813 (N_9813,N_4281,N_4473);
nand U9814 (N_9814,N_1122,N_1599);
nand U9815 (N_9815,N_2313,N_2725);
nor U9816 (N_9816,N_1004,N_2689);
and U9817 (N_9817,N_628,N_3799);
or U9818 (N_9818,N_3456,N_1818);
nand U9819 (N_9819,N_1862,N_869);
nor U9820 (N_9820,N_4461,N_4959);
and U9821 (N_9821,N_2843,N_1855);
or U9822 (N_9822,N_2538,N_1937);
and U9823 (N_9823,N_3485,N_2025);
and U9824 (N_9824,N_4271,N_4516);
xnor U9825 (N_9825,N_2223,N_2016);
or U9826 (N_9826,N_2453,N_1934);
and U9827 (N_9827,N_3669,N_2027);
or U9828 (N_9828,N_2661,N_791);
nand U9829 (N_9829,N_2497,N_43);
nor U9830 (N_9830,N_489,N_3632);
nand U9831 (N_9831,N_3277,N_833);
nand U9832 (N_9832,N_3884,N_1080);
or U9833 (N_9833,N_4310,N_3661);
or U9834 (N_9834,N_3471,N_3983);
and U9835 (N_9835,N_4683,N_4316);
and U9836 (N_9836,N_616,N_1329);
nor U9837 (N_9837,N_3994,N_3191);
and U9838 (N_9838,N_1183,N_1059);
or U9839 (N_9839,N_4975,N_3376);
nand U9840 (N_9840,N_3032,N_4023);
or U9841 (N_9841,N_1029,N_1851);
nand U9842 (N_9842,N_1254,N_1709);
and U9843 (N_9843,N_2961,N_3570);
nand U9844 (N_9844,N_3368,N_3459);
and U9845 (N_9845,N_321,N_3707);
nand U9846 (N_9846,N_1344,N_3768);
or U9847 (N_9847,N_2174,N_3570);
nand U9848 (N_9848,N_824,N_2944);
and U9849 (N_9849,N_2589,N_3414);
or U9850 (N_9850,N_4059,N_2467);
or U9851 (N_9851,N_4732,N_529);
nand U9852 (N_9852,N_4917,N_3652);
nand U9853 (N_9853,N_4624,N_2201);
and U9854 (N_9854,N_2185,N_3450);
and U9855 (N_9855,N_4400,N_1402);
nand U9856 (N_9856,N_3319,N_200);
nand U9857 (N_9857,N_171,N_3402);
and U9858 (N_9858,N_1852,N_2798);
nand U9859 (N_9859,N_3932,N_1942);
or U9860 (N_9860,N_4368,N_905);
nand U9861 (N_9861,N_4500,N_3107);
nor U9862 (N_9862,N_1873,N_2193);
or U9863 (N_9863,N_4309,N_495);
or U9864 (N_9864,N_2653,N_1779);
and U9865 (N_9865,N_4478,N_2953);
nor U9866 (N_9866,N_3946,N_3859);
or U9867 (N_9867,N_301,N_3069);
and U9868 (N_9868,N_2806,N_1965);
nor U9869 (N_9869,N_3215,N_4132);
or U9870 (N_9870,N_2652,N_3009);
nor U9871 (N_9871,N_4310,N_2755);
and U9872 (N_9872,N_451,N_3070);
nor U9873 (N_9873,N_4935,N_4348);
nor U9874 (N_9874,N_3543,N_1643);
nor U9875 (N_9875,N_1268,N_2029);
and U9876 (N_9876,N_3871,N_229);
nor U9877 (N_9877,N_1517,N_3993);
and U9878 (N_9878,N_410,N_774);
or U9879 (N_9879,N_2024,N_2143);
nand U9880 (N_9880,N_2790,N_3682);
and U9881 (N_9881,N_2847,N_2161);
and U9882 (N_9882,N_3755,N_1379);
nand U9883 (N_9883,N_4160,N_4429);
nor U9884 (N_9884,N_3031,N_3366);
or U9885 (N_9885,N_3812,N_200);
nor U9886 (N_9886,N_2658,N_2148);
nand U9887 (N_9887,N_4360,N_4564);
and U9888 (N_9888,N_888,N_2877);
nor U9889 (N_9889,N_2295,N_2398);
nand U9890 (N_9890,N_547,N_3014);
or U9891 (N_9891,N_927,N_3829);
nand U9892 (N_9892,N_4053,N_2417);
and U9893 (N_9893,N_801,N_2777);
or U9894 (N_9894,N_4279,N_2170);
or U9895 (N_9895,N_724,N_240);
xnor U9896 (N_9896,N_2861,N_4928);
nor U9897 (N_9897,N_1758,N_4167);
and U9898 (N_9898,N_1516,N_4746);
nand U9899 (N_9899,N_3373,N_2697);
nand U9900 (N_9900,N_34,N_1242);
nor U9901 (N_9901,N_1350,N_1090);
nand U9902 (N_9902,N_4353,N_3407);
or U9903 (N_9903,N_2660,N_1860);
or U9904 (N_9904,N_2872,N_1817);
or U9905 (N_9905,N_499,N_804);
nand U9906 (N_9906,N_1621,N_331);
or U9907 (N_9907,N_747,N_1334);
nor U9908 (N_9908,N_1303,N_4505);
xor U9909 (N_9909,N_2930,N_2680);
nand U9910 (N_9910,N_791,N_149);
nor U9911 (N_9911,N_3111,N_1565);
or U9912 (N_9912,N_3431,N_4535);
or U9913 (N_9913,N_2354,N_4154);
nor U9914 (N_9914,N_2660,N_3743);
nand U9915 (N_9915,N_1358,N_4387);
or U9916 (N_9916,N_728,N_1372);
nor U9917 (N_9917,N_545,N_2970);
or U9918 (N_9918,N_2021,N_1171);
and U9919 (N_9919,N_4769,N_4092);
or U9920 (N_9920,N_1218,N_453);
or U9921 (N_9921,N_4536,N_2914);
and U9922 (N_9922,N_4610,N_4979);
nor U9923 (N_9923,N_4553,N_4973);
nand U9924 (N_9924,N_4979,N_2921);
or U9925 (N_9925,N_3879,N_34);
nor U9926 (N_9926,N_1760,N_4226);
and U9927 (N_9927,N_408,N_4342);
nand U9928 (N_9928,N_4642,N_637);
nor U9929 (N_9929,N_3595,N_1491);
nand U9930 (N_9930,N_789,N_1575);
and U9931 (N_9931,N_3704,N_1264);
nor U9932 (N_9932,N_749,N_3404);
and U9933 (N_9933,N_4973,N_416);
nand U9934 (N_9934,N_1351,N_4458);
or U9935 (N_9935,N_4502,N_1792);
or U9936 (N_9936,N_2143,N_4765);
and U9937 (N_9937,N_1556,N_14);
and U9938 (N_9938,N_4948,N_3044);
or U9939 (N_9939,N_1517,N_4559);
and U9940 (N_9940,N_3622,N_1457);
nand U9941 (N_9941,N_2030,N_1127);
or U9942 (N_9942,N_4038,N_4149);
and U9943 (N_9943,N_910,N_1556);
and U9944 (N_9944,N_2079,N_2285);
and U9945 (N_9945,N_3417,N_918);
nand U9946 (N_9946,N_1437,N_4740);
and U9947 (N_9947,N_2002,N_1429);
or U9948 (N_9948,N_3584,N_3844);
nor U9949 (N_9949,N_367,N_4967);
or U9950 (N_9950,N_4859,N_3994);
nor U9951 (N_9951,N_1604,N_4854);
nor U9952 (N_9952,N_990,N_245);
nor U9953 (N_9953,N_4219,N_4437);
and U9954 (N_9954,N_621,N_4776);
and U9955 (N_9955,N_2808,N_682);
or U9956 (N_9956,N_1411,N_1362);
nor U9957 (N_9957,N_3170,N_4793);
and U9958 (N_9958,N_230,N_643);
and U9959 (N_9959,N_3973,N_612);
and U9960 (N_9960,N_2110,N_2939);
nand U9961 (N_9961,N_464,N_2130);
nand U9962 (N_9962,N_2199,N_351);
or U9963 (N_9963,N_3132,N_2776);
nand U9964 (N_9964,N_2892,N_393);
nor U9965 (N_9965,N_2981,N_2786);
nand U9966 (N_9966,N_3103,N_2284);
or U9967 (N_9967,N_2863,N_4930);
and U9968 (N_9968,N_2630,N_490);
nand U9969 (N_9969,N_3166,N_109);
nand U9970 (N_9970,N_2056,N_2372);
or U9971 (N_9971,N_286,N_3930);
and U9972 (N_9972,N_3456,N_1508);
nor U9973 (N_9973,N_1272,N_2744);
nand U9974 (N_9974,N_2977,N_694);
or U9975 (N_9975,N_4862,N_980);
or U9976 (N_9976,N_682,N_3385);
or U9977 (N_9977,N_3185,N_2589);
nand U9978 (N_9978,N_4056,N_734);
nand U9979 (N_9979,N_2180,N_3923);
nor U9980 (N_9980,N_4315,N_1286);
nor U9981 (N_9981,N_140,N_1750);
or U9982 (N_9982,N_1998,N_1170);
nand U9983 (N_9983,N_1835,N_1412);
nand U9984 (N_9984,N_1725,N_2801);
nor U9985 (N_9985,N_3234,N_3584);
and U9986 (N_9986,N_1907,N_1523);
nor U9987 (N_9987,N_4674,N_2013);
or U9988 (N_9988,N_4932,N_3383);
or U9989 (N_9989,N_729,N_1858);
or U9990 (N_9990,N_3524,N_2944);
and U9991 (N_9991,N_2001,N_4313);
nor U9992 (N_9992,N_673,N_2238);
nor U9993 (N_9993,N_4593,N_1147);
nor U9994 (N_9994,N_2086,N_1992);
nor U9995 (N_9995,N_1797,N_4003);
nor U9996 (N_9996,N_3668,N_2560);
nor U9997 (N_9997,N_4696,N_3749);
nand U9998 (N_9998,N_493,N_488);
and U9999 (N_9999,N_714,N_3855);
nor U10000 (N_10000,N_6596,N_7373);
or U10001 (N_10001,N_8235,N_5168);
or U10002 (N_10002,N_6362,N_7124);
or U10003 (N_10003,N_7548,N_5220);
nor U10004 (N_10004,N_9909,N_9913);
nor U10005 (N_10005,N_7767,N_5929);
nand U10006 (N_10006,N_7953,N_9427);
nand U10007 (N_10007,N_9880,N_8499);
nor U10008 (N_10008,N_9044,N_9529);
nand U10009 (N_10009,N_5225,N_6508);
nor U10010 (N_10010,N_6083,N_6529);
nor U10011 (N_10011,N_9174,N_8801);
nor U10012 (N_10012,N_5192,N_6289);
and U10013 (N_10013,N_9714,N_6949);
and U10014 (N_10014,N_8110,N_7570);
nor U10015 (N_10015,N_9741,N_7540);
nor U10016 (N_10016,N_5141,N_6991);
nor U10017 (N_10017,N_6907,N_5412);
nand U10018 (N_10018,N_8470,N_5780);
nor U10019 (N_10019,N_8089,N_9452);
nor U10020 (N_10020,N_6293,N_9480);
nand U10021 (N_10021,N_8493,N_9651);
nor U10022 (N_10022,N_9989,N_7948);
nor U10023 (N_10023,N_7376,N_6214);
or U10024 (N_10024,N_7895,N_9080);
nand U10025 (N_10025,N_7592,N_5006);
nand U10026 (N_10026,N_5932,N_9484);
or U10027 (N_10027,N_6054,N_5848);
or U10028 (N_10028,N_9949,N_9816);
nor U10029 (N_10029,N_6900,N_5745);
and U10030 (N_10030,N_5510,N_8805);
nand U10031 (N_10031,N_6252,N_6910);
and U10032 (N_10032,N_5113,N_6635);
nand U10033 (N_10033,N_7831,N_8619);
and U10034 (N_10034,N_8646,N_7112);
and U10035 (N_10035,N_9306,N_5421);
nor U10036 (N_10036,N_7572,N_8196);
and U10037 (N_10037,N_5472,N_5718);
nand U10038 (N_10038,N_5495,N_5404);
nand U10039 (N_10039,N_6776,N_8552);
and U10040 (N_10040,N_9984,N_9338);
nand U10041 (N_10041,N_5728,N_6905);
and U10042 (N_10042,N_8520,N_6786);
nor U10043 (N_10043,N_7947,N_9744);
nor U10044 (N_10044,N_7941,N_5329);
nor U10045 (N_10045,N_9551,N_8635);
nand U10046 (N_10046,N_5456,N_5528);
or U10047 (N_10047,N_7626,N_6393);
nor U10048 (N_10048,N_8239,N_5761);
and U10049 (N_10049,N_7232,N_7900);
or U10050 (N_10050,N_7510,N_5673);
nand U10051 (N_10051,N_5099,N_7068);
or U10052 (N_10052,N_7099,N_8905);
nor U10053 (N_10053,N_9535,N_5531);
and U10054 (N_10054,N_8639,N_7575);
or U10055 (N_10055,N_8878,N_5633);
nor U10056 (N_10056,N_5652,N_5631);
and U10057 (N_10057,N_5077,N_6833);
and U10058 (N_10058,N_5224,N_7425);
and U10059 (N_10059,N_9898,N_9593);
nand U10060 (N_10060,N_9790,N_5590);
or U10061 (N_10061,N_8178,N_9942);
and U10062 (N_10062,N_5587,N_7738);
and U10063 (N_10063,N_8935,N_6963);
or U10064 (N_10064,N_7054,N_9148);
nand U10065 (N_10065,N_8651,N_7455);
nor U10066 (N_10066,N_7633,N_6025);
nand U10067 (N_10067,N_6583,N_6008);
xor U10068 (N_10068,N_6241,N_8741);
or U10069 (N_10069,N_8773,N_6139);
nor U10070 (N_10070,N_5488,N_9724);
and U10071 (N_10071,N_7913,N_9681);
and U10072 (N_10072,N_5010,N_8155);
and U10073 (N_10073,N_5609,N_5941);
or U10074 (N_10074,N_6480,N_7549);
and U10075 (N_10075,N_6816,N_7166);
nand U10076 (N_10076,N_8461,N_6960);
nand U10077 (N_10077,N_5945,N_7008);
nor U10078 (N_10078,N_7389,N_5847);
and U10079 (N_10079,N_5616,N_9615);
nand U10080 (N_10080,N_8133,N_9751);
and U10081 (N_10081,N_9515,N_8414);
nand U10082 (N_10082,N_9738,N_8477);
nor U10083 (N_10083,N_8015,N_5038);
nand U10084 (N_10084,N_8980,N_6673);
or U10085 (N_10085,N_6953,N_9396);
and U10086 (N_10086,N_5557,N_6923);
or U10087 (N_10087,N_5452,N_7466);
nor U10088 (N_10088,N_8377,N_6416);
nand U10089 (N_10089,N_9934,N_6533);
or U10090 (N_10090,N_8299,N_5982);
nand U10091 (N_10091,N_9394,N_6282);
or U10092 (N_10092,N_5835,N_9386);
nand U10093 (N_10093,N_6917,N_6858);
or U10094 (N_10094,N_5800,N_7266);
nand U10095 (N_10095,N_8127,N_5730);
or U10096 (N_10096,N_6494,N_8753);
or U10097 (N_10097,N_5123,N_9550);
or U10098 (N_10098,N_5551,N_7140);
nor U10099 (N_10099,N_8230,N_9178);
nand U10100 (N_10100,N_8843,N_5623);
nand U10101 (N_10101,N_7305,N_8778);
and U10102 (N_10102,N_9666,N_9585);
nor U10103 (N_10103,N_6836,N_5217);
and U10104 (N_10104,N_6660,N_5555);
nand U10105 (N_10105,N_7826,N_9848);
xor U10106 (N_10106,N_6514,N_9892);
or U10107 (N_10107,N_7384,N_6137);
xor U10108 (N_10108,N_7639,N_6348);
and U10109 (N_10109,N_8537,N_8571);
nor U10110 (N_10110,N_9628,N_9004);
nor U10111 (N_10111,N_9123,N_7370);
and U10112 (N_10112,N_8433,N_6202);
nor U10113 (N_10113,N_5216,N_9111);
and U10114 (N_10114,N_6688,N_9041);
or U10115 (N_10115,N_6754,N_6271);
and U10116 (N_10116,N_6796,N_8623);
or U10117 (N_10117,N_5361,N_9289);
nand U10118 (N_10118,N_9654,N_6722);
or U10119 (N_10119,N_7462,N_9693);
or U10120 (N_10120,N_6893,N_6195);
nand U10121 (N_10121,N_7434,N_6255);
or U10122 (N_10122,N_8146,N_9150);
nand U10123 (N_10123,N_6043,N_7878);
and U10124 (N_10124,N_8519,N_9699);
and U10125 (N_10125,N_7977,N_6110);
and U10126 (N_10126,N_7753,N_5271);
and U10127 (N_10127,N_8601,N_7302);
nand U10128 (N_10128,N_7984,N_9166);
nor U10129 (N_10129,N_5622,N_6570);
or U10130 (N_10130,N_5773,N_9937);
nor U10131 (N_10131,N_6421,N_5397);
nand U10132 (N_10132,N_7331,N_5459);
and U10133 (N_10133,N_7970,N_8478);
and U10134 (N_10134,N_7696,N_6445);
nor U10135 (N_10135,N_5081,N_8047);
and U10136 (N_10136,N_9733,N_8175);
nor U10137 (N_10137,N_8349,N_9800);
or U10138 (N_10138,N_8294,N_7689);
or U10139 (N_10139,N_8347,N_6151);
or U10140 (N_10140,N_5339,N_8914);
and U10141 (N_10141,N_5749,N_5502);
nor U10142 (N_10142,N_8279,N_9182);
nor U10143 (N_10143,N_9927,N_9846);
nand U10144 (N_10144,N_7100,N_6857);
nand U10145 (N_10145,N_9031,N_8247);
or U10146 (N_10146,N_7388,N_5065);
nand U10147 (N_10147,N_5177,N_6048);
nor U10148 (N_10148,N_9808,N_7141);
and U10149 (N_10149,N_7902,N_5428);
or U10150 (N_10150,N_8617,N_6033);
nor U10151 (N_10151,N_6321,N_5444);
nand U10152 (N_10152,N_6668,N_7629);
nor U10153 (N_10153,N_8541,N_9948);
and U10154 (N_10154,N_6211,N_9778);
and U10155 (N_10155,N_5732,N_9684);
and U10156 (N_10156,N_7892,N_7855);
nand U10157 (N_10157,N_5267,N_6361);
nand U10158 (N_10158,N_8565,N_9587);
nand U10159 (N_10159,N_5525,N_7824);
xor U10160 (N_10160,N_5764,N_9385);
nor U10161 (N_10161,N_8290,N_5788);
and U10162 (N_10162,N_7194,N_9655);
or U10163 (N_10163,N_5309,N_5666);
and U10164 (N_10164,N_9656,N_7092);
and U10165 (N_10165,N_5526,N_8380);
nand U10166 (N_10166,N_6004,N_8119);
nand U10167 (N_10167,N_5147,N_5593);
or U10168 (N_10168,N_8798,N_5599);
or U10169 (N_10169,N_9798,N_6178);
nor U10170 (N_10170,N_6274,N_9955);
and U10171 (N_10171,N_6505,N_5056);
nor U10172 (N_10172,N_8486,N_5839);
and U10173 (N_10173,N_7918,N_9036);
and U10174 (N_10174,N_6853,N_8013);
nor U10175 (N_10175,N_8403,N_5713);
nor U10176 (N_10176,N_6653,N_5506);
nor U10177 (N_10177,N_6962,N_6888);
and U10178 (N_10178,N_5205,N_9265);
and U10179 (N_10179,N_5176,N_7555);
nor U10180 (N_10180,N_6469,N_5111);
and U10181 (N_10181,N_5034,N_8694);
nor U10182 (N_10182,N_5658,N_5376);
nor U10183 (N_10183,N_6777,N_8123);
nor U10184 (N_10184,N_8592,N_8131);
nand U10185 (N_10185,N_8944,N_5659);
nor U10186 (N_10186,N_8543,N_9904);
or U10187 (N_10187,N_8720,N_7714);
and U10188 (N_10188,N_9033,N_6801);
and U10189 (N_10189,N_7085,N_5246);
or U10190 (N_10190,N_6657,N_7760);
nand U10191 (N_10191,N_6984,N_6109);
and U10192 (N_10192,N_8803,N_6895);
nor U10193 (N_10193,N_6709,N_5569);
nand U10194 (N_10194,N_6671,N_7833);
or U10195 (N_10195,N_5247,N_8032);
and U10196 (N_10196,N_9809,N_8802);
and U10197 (N_10197,N_9956,N_7227);
and U10198 (N_10198,N_8590,N_8823);
nand U10199 (N_10199,N_8771,N_9102);
and U10200 (N_10200,N_7410,N_5942);
and U10201 (N_10201,N_9154,N_7143);
nand U10202 (N_10202,N_5364,N_7414);
nor U10203 (N_10203,N_5200,N_8615);
and U10204 (N_10204,N_6436,N_7508);
and U10205 (N_10205,N_8305,N_9418);
nor U10206 (N_10206,N_8036,N_5490);
nand U10207 (N_10207,N_8585,N_6001);
nor U10208 (N_10208,N_6028,N_9364);
nand U10209 (N_10209,N_6503,N_9944);
or U10210 (N_10210,N_8974,N_9629);
or U10211 (N_10211,N_9826,N_6000);
or U10212 (N_10212,N_8197,N_9345);
nand U10213 (N_10213,N_9737,N_9595);
nand U10214 (N_10214,N_5621,N_9363);
or U10215 (N_10215,N_9965,N_8763);
nand U10216 (N_10216,N_6546,N_8557);
nand U10217 (N_10217,N_6523,N_7197);
and U10218 (N_10218,N_6180,N_9392);
or U10219 (N_10219,N_9918,N_7547);
and U10220 (N_10220,N_7939,N_6153);
or U10221 (N_10221,N_8733,N_6471);
and U10222 (N_10222,N_9572,N_9627);
or U10223 (N_10223,N_6248,N_9841);
or U10224 (N_10224,N_9131,N_8917);
nand U10225 (N_10225,N_7774,N_9683);
or U10226 (N_10226,N_9725,N_8472);
nor U10227 (N_10227,N_6056,N_5004);
nor U10228 (N_10228,N_9505,N_9433);
or U10229 (N_10229,N_6041,N_9181);
nor U10230 (N_10230,N_9114,N_9717);
nor U10231 (N_10231,N_8715,N_7125);
and U10232 (N_10232,N_7418,N_8017);
nor U10233 (N_10233,N_5273,N_6820);
nand U10234 (N_10234,N_8467,N_8388);
and U10235 (N_10235,N_8528,N_7887);
and U10236 (N_10236,N_9488,N_5119);
nand U10237 (N_10237,N_6017,N_6579);
and U10238 (N_10238,N_7215,N_6415);
or U10239 (N_10239,N_9482,N_9916);
or U10240 (N_10240,N_6597,N_7867);
nand U10241 (N_10241,N_7568,N_8689);
and U10242 (N_10242,N_8220,N_8855);
and U10243 (N_10243,N_8242,N_8150);
or U10244 (N_10244,N_9066,N_8469);
nor U10245 (N_10245,N_8208,N_8986);
and U10246 (N_10246,N_8597,N_9795);
and U10247 (N_10247,N_5831,N_6342);
and U10248 (N_10248,N_7239,N_9255);
nor U10249 (N_10249,N_6954,N_7451);
nor U10250 (N_10250,N_7643,N_6213);
nor U10251 (N_10251,N_8393,N_6881);
nand U10252 (N_10252,N_7603,N_5933);
and U10253 (N_10253,N_9623,N_7890);
or U10254 (N_10254,N_8384,N_7365);
nor U10255 (N_10255,N_9202,N_8834);
nor U10256 (N_10256,N_9228,N_7993);
nand U10257 (N_10257,N_6427,N_8492);
and U10258 (N_10258,N_8337,N_6283);
nor U10259 (N_10259,N_7556,N_7228);
or U10260 (N_10260,N_6740,N_8756);
and U10261 (N_10261,N_7914,N_5377);
and U10262 (N_10262,N_9141,N_7704);
or U10263 (N_10263,N_7796,N_9569);
or U10264 (N_10264,N_8460,N_8121);
and U10265 (N_10265,N_7539,N_7981);
nor U10266 (N_10266,N_5044,N_6735);
or U10267 (N_10267,N_8832,N_5771);
or U10268 (N_10268,N_5998,N_6485);
or U10269 (N_10269,N_9945,N_8484);
or U10270 (N_10270,N_5861,N_6846);
or U10271 (N_10271,N_9384,N_8028);
and U10272 (N_10272,N_8359,N_7357);
or U10273 (N_10273,N_6639,N_8656);
nand U10274 (N_10274,N_8475,N_7298);
nand U10275 (N_10275,N_9539,N_6080);
nor U10276 (N_10276,N_5285,N_7048);
nand U10277 (N_10277,N_7505,N_8732);
and U10278 (N_10278,N_5331,N_5640);
and U10279 (N_10279,N_5539,N_9491);
and U10280 (N_10280,N_6852,N_7135);
nand U10281 (N_10281,N_9755,N_5386);
nor U10282 (N_10282,N_7579,N_9715);
nor U10283 (N_10283,N_5908,N_6383);
nand U10284 (N_10284,N_9653,N_5524);
or U10285 (N_10285,N_8903,N_6114);
nand U10286 (N_10286,N_5068,N_5729);
or U10287 (N_10287,N_6473,N_8099);
nand U10288 (N_10288,N_5212,N_6179);
or U10289 (N_10289,N_7148,N_9722);
nor U10290 (N_10290,N_6284,N_8668);
and U10291 (N_10291,N_9436,N_5035);
nand U10292 (N_10292,N_9037,N_7369);
and U10293 (N_10293,N_8943,N_7992);
nor U10294 (N_10294,N_9251,N_5282);
nor U10295 (N_10295,N_8016,N_5234);
nand U10296 (N_10296,N_5867,N_8244);
or U10297 (N_10297,N_7624,N_5442);
and U10298 (N_10298,N_7108,N_6059);
nand U10299 (N_10299,N_8971,N_6423);
nor U10300 (N_10300,N_8125,N_6357);
nand U10301 (N_10301,N_5134,N_5978);
nand U10302 (N_10302,N_6968,N_7938);
nor U10303 (N_10303,N_9940,N_9409);
nor U10304 (N_10304,N_8923,N_5008);
or U10305 (N_10305,N_9294,N_8824);
or U10306 (N_10306,N_7881,N_9872);
nand U10307 (N_10307,N_7631,N_7296);
and U10308 (N_10308,N_9865,N_5326);
or U10309 (N_10309,N_9618,N_5030);
nand U10310 (N_10310,N_7946,N_5135);
and U10311 (N_10311,N_8077,N_8648);
nand U10312 (N_10312,N_9007,N_9602);
and U10313 (N_10313,N_5612,N_8727);
nor U10314 (N_10314,N_8961,N_9512);
nor U10315 (N_10315,N_9967,N_7743);
nand U10316 (N_10316,N_7002,N_9132);
or U10317 (N_10317,N_6199,N_6868);
nor U10318 (N_10318,N_6340,N_6363);
nand U10319 (N_10319,N_7276,N_6078);
or U10320 (N_10320,N_7080,N_9663);
and U10321 (N_10321,N_5668,N_8796);
and U10322 (N_10322,N_6101,N_5603);
nand U10323 (N_10323,N_5855,N_8630);
nor U10324 (N_10324,N_6859,N_9526);
or U10325 (N_10325,N_8082,N_5284);
nand U10326 (N_10326,N_8872,N_7628);
and U10327 (N_10327,N_6064,N_8516);
nand U10328 (N_10328,N_8456,N_5228);
nor U10329 (N_10329,N_5950,N_6049);
and U10330 (N_10330,N_9946,N_7289);
and U10331 (N_10331,N_8454,N_8049);
and U10332 (N_10332,N_7820,N_7072);
nand U10333 (N_10333,N_8088,N_9827);
xor U10334 (N_10334,N_6159,N_9175);
or U10335 (N_10335,N_9270,N_5464);
nor U10336 (N_10336,N_7485,N_5100);
and U10337 (N_10337,N_9692,N_5214);
and U10338 (N_10338,N_6337,N_5450);
nor U10339 (N_10339,N_7105,N_7793);
nand U10340 (N_10340,N_7091,N_7907);
nand U10341 (N_10341,N_7996,N_7898);
or U10342 (N_10342,N_8613,N_9701);
nor U10343 (N_10343,N_9375,N_5682);
or U10344 (N_10344,N_5893,N_5074);
or U10345 (N_10345,N_9443,N_5317);
xor U10346 (N_10346,N_6094,N_8309);
or U10347 (N_10347,N_9072,N_7687);
or U10348 (N_10348,N_6980,N_5804);
nor U10349 (N_10349,N_9720,N_5070);
nor U10350 (N_10350,N_8936,N_7581);
nor U10351 (N_10351,N_7545,N_6990);
nand U10352 (N_10352,N_6455,N_9838);
or U10353 (N_10353,N_5744,N_7392);
and U10354 (N_10354,N_5253,N_8404);
nor U10355 (N_10355,N_9533,N_7374);
or U10356 (N_10356,N_5532,N_5431);
nand U10357 (N_10357,N_8334,N_9914);
nand U10358 (N_10358,N_6850,N_6057);
nand U10359 (N_10359,N_5232,N_9532);
nor U10360 (N_10360,N_6322,N_5811);
and U10361 (N_10361,N_5476,N_8394);
nand U10362 (N_10362,N_7612,N_5915);
nand U10363 (N_10363,N_6175,N_9911);
nor U10364 (N_10364,N_9110,N_6693);
nand U10365 (N_10365,N_7870,N_6650);
nor U10366 (N_10366,N_6120,N_8106);
nand U10367 (N_10367,N_6752,N_8268);
nand U10368 (N_10368,N_5249,N_7901);
and U10369 (N_10369,N_6769,N_8241);
or U10370 (N_10370,N_9679,N_6560);
or U10371 (N_10371,N_6612,N_7983);
and U10372 (N_10372,N_5142,N_9038);
or U10373 (N_10373,N_7912,N_6634);
and U10374 (N_10374,N_6860,N_8417);
nand U10375 (N_10375,N_9428,N_5521);
nand U10376 (N_10376,N_7372,N_6897);
and U10377 (N_10377,N_8779,N_7066);
nor U10378 (N_10378,N_7347,N_9691);
nor U10379 (N_10379,N_6005,N_7223);
or U10380 (N_10380,N_9735,N_8857);
nor U10381 (N_10381,N_7001,N_9027);
nor U10382 (N_10382,N_5211,N_5333);
nand U10383 (N_10383,N_6728,N_5629);
or U10384 (N_10384,N_9917,N_5693);
and U10385 (N_10385,N_7644,N_8233);
or U10386 (N_10386,N_7187,N_9746);
nand U10387 (N_10387,N_8819,N_6988);
nor U10388 (N_10388,N_7611,N_7720);
and U10389 (N_10389,N_8023,N_9857);
and U10390 (N_10390,N_9307,N_7730);
or U10391 (N_10391,N_7103,N_5426);
or U10392 (N_10392,N_5434,N_5422);
xnor U10393 (N_10393,N_6349,N_6746);
nand U10394 (N_10394,N_7514,N_6484);
nor U10395 (N_10395,N_9964,N_6975);
and U10396 (N_10396,N_9009,N_5257);
nand U10397 (N_10397,N_6931,N_9835);
nand U10398 (N_10398,N_5832,N_8907);
or U10399 (N_10399,N_8511,N_9630);
or U10400 (N_10400,N_7569,N_6593);
nand U10401 (N_10401,N_8224,N_8530);
nand U10402 (N_10402,N_8722,N_8285);
and U10403 (N_10403,N_9264,N_6924);
and U10404 (N_10404,N_7731,N_6997);
nand U10405 (N_10405,N_6036,N_6594);
nor U10406 (N_10406,N_6228,N_7963);
nor U10407 (N_10407,N_5115,N_9951);
nor U10408 (N_10408,N_9634,N_8940);
and U10409 (N_10409,N_8289,N_8594);
nand U10410 (N_10410,N_5605,N_5864);
and U10411 (N_10411,N_9355,N_5449);
and U10412 (N_10412,N_9574,N_6664);
or U10413 (N_10413,N_9130,N_5678);
nand U10414 (N_10414,N_9069,N_9299);
nor U10415 (N_10415,N_7708,N_9406);
nand U10416 (N_10416,N_5302,N_6744);
nor U10417 (N_10417,N_8743,N_6959);
and U10418 (N_10418,N_5890,N_5988);
nand U10419 (N_10419,N_6067,N_7649);
nor U10420 (N_10420,N_5344,N_7079);
nor U10421 (N_10421,N_7034,N_6144);
and U10422 (N_10422,N_9843,N_7747);
nor U10423 (N_10423,N_9943,N_9643);
nor U10424 (N_10424,N_8225,N_7529);
or U10425 (N_10425,N_8654,N_6877);
and U10426 (N_10426,N_5938,N_8343);
nor U10427 (N_10427,N_5983,N_9839);
nand U10428 (N_10428,N_9960,N_7356);
and U10429 (N_10429,N_6206,N_5703);
nor U10430 (N_10430,N_9567,N_8055);
nand U10431 (N_10431,N_8395,N_9779);
nand U10432 (N_10432,N_5436,N_5063);
nor U10433 (N_10433,N_5101,N_7111);
nor U10434 (N_10434,N_6136,N_6075);
and U10435 (N_10435,N_9584,N_9382);
and U10436 (N_10436,N_8117,N_6768);
nor U10437 (N_10437,N_9985,N_8702);
or U10438 (N_10438,N_5189,N_8717);
nand U10439 (N_10439,N_5316,N_6173);
nor U10440 (N_10440,N_7192,N_5304);
and U10441 (N_10441,N_6684,N_9250);
nand U10442 (N_10442,N_8793,N_6767);
nand U10443 (N_10443,N_9248,N_6148);
nor U10444 (N_10444,N_5834,N_6551);
nand U10445 (N_10445,N_8092,N_5306);
nand U10446 (N_10446,N_9050,N_6802);
nor U10447 (N_10447,N_6675,N_6239);
nand U10448 (N_10448,N_8628,N_8994);
or U10449 (N_10449,N_9117,N_7674);
nand U10450 (N_10450,N_8262,N_8981);
and U10451 (N_10451,N_6243,N_7284);
nand U10452 (N_10452,N_8153,N_5467);
nand U10453 (N_10453,N_8351,N_9026);
nand U10454 (N_10454,N_7903,N_6176);
nand U10455 (N_10455,N_8817,N_8988);
nand U10456 (N_10456,N_6230,N_9035);
nand U10457 (N_10457,N_7952,N_8072);
nand U10458 (N_10458,N_5385,N_7083);
and U10459 (N_10459,N_8218,N_9668);
or U10460 (N_10460,N_7333,N_6805);
and U10461 (N_10461,N_8479,N_7813);
nand U10462 (N_10462,N_5440,N_6609);
nor U10463 (N_10463,N_9499,N_9052);
or U10464 (N_10464,N_7709,N_9136);
or U10465 (N_10465,N_8589,N_8222);
nand U10466 (N_10466,N_8671,N_5482);
or U10467 (N_10467,N_9576,N_6755);
or U10468 (N_10468,N_7229,N_8256);
or U10469 (N_10469,N_5454,N_9979);
and U10470 (N_10470,N_7443,N_5453);
or U10471 (N_10471,N_7828,N_6135);
or U10472 (N_10472,N_6944,N_5705);
nor U10473 (N_10473,N_5512,N_6130);
nor U10474 (N_10474,N_8288,N_5592);
nor U10475 (N_10475,N_7620,N_8647);
nand U10476 (N_10476,N_5810,N_5158);
nor U10477 (N_10477,N_8664,N_8205);
or U10478 (N_10478,N_7551,N_7562);
or U10479 (N_10479,N_8443,N_9308);
and U10480 (N_10480,N_9465,N_5507);
or U10481 (N_10481,N_9998,N_7698);
or U10482 (N_10482,N_9145,N_9098);
nand U10483 (N_10483,N_9177,N_5584);
nor U10484 (N_10484,N_5020,N_6575);
and U10485 (N_10485,N_5420,N_9146);
and U10486 (N_10486,N_5727,N_5033);
and U10487 (N_10487,N_6902,N_9899);
nor U10488 (N_10488,N_6536,N_9680);
or U10489 (N_10489,N_6809,N_5536);
nand U10490 (N_10490,N_9451,N_7646);
and U10491 (N_10491,N_5628,N_9993);
or U10492 (N_10492,N_9811,N_5994);
and U10493 (N_10493,N_9407,N_5213);
or U10494 (N_10494,N_9401,N_5611);
nor U10495 (N_10495,N_7464,N_6463);
or U10496 (N_10496,N_6003,N_7859);
or U10497 (N_10497,N_6527,N_5279);
nand U10498 (N_10498,N_7557,N_8397);
and U10499 (N_10499,N_6224,N_5350);
nor U10500 (N_10500,N_5617,N_8626);
or U10501 (N_10501,N_7145,N_5563);
nand U10502 (N_10502,N_5719,N_5545);
and U10503 (N_10503,N_6627,N_6652);
or U10504 (N_10504,N_9119,N_5527);
nand U10505 (N_10505,N_7801,N_8749);
nand U10506 (N_10506,N_9820,N_5486);
or U10507 (N_10507,N_6045,N_7653);
nor U10508 (N_10508,N_9700,N_5916);
and U10509 (N_10509,N_8536,N_7257);
nand U10510 (N_10510,N_7172,N_5849);
or U10511 (N_10511,N_8789,N_5297);
or U10512 (N_10512,N_8984,N_7173);
nor U10513 (N_10513,N_7470,N_7537);
or U10514 (N_10514,N_5263,N_6294);
nand U10515 (N_10515,N_5071,N_9245);
or U10516 (N_10516,N_5875,N_7673);
and U10517 (N_10517,N_7408,N_8570);
or U10518 (N_10518,N_9344,N_5126);
xor U10519 (N_10519,N_6738,N_5921);
or U10520 (N_10520,N_5708,N_6345);
nand U10521 (N_10521,N_6764,N_8042);
or U10522 (N_10522,N_5425,N_8711);
and U10523 (N_10523,N_6411,N_6194);
nor U10524 (N_10524,N_9817,N_6861);
nand U10525 (N_10525,N_8658,N_5489);
nor U10526 (N_10526,N_9890,N_8742);
nor U10527 (N_10527,N_7291,N_9510);
nor U10528 (N_10528,N_8161,N_6989);
nand U10529 (N_10529,N_8967,N_9365);
or U10530 (N_10530,N_5466,N_7437);
or U10531 (N_10531,N_8071,N_5144);
nor U10532 (N_10532,N_7661,N_6882);
and U10533 (N_10533,N_8396,N_7515);
nor U10534 (N_10534,N_8572,N_7538);
or U10535 (N_10535,N_7049,N_9350);
and U10536 (N_10536,N_9970,N_7615);
and U10537 (N_10537,N_6373,N_5173);
or U10538 (N_10538,N_8159,N_6966);
and U10539 (N_10539,N_5405,N_5777);
and U10540 (N_10540,N_5974,N_7536);
nor U10541 (N_10541,N_5438,N_5962);
and U10542 (N_10542,N_5806,N_7886);
or U10543 (N_10543,N_6800,N_9754);
nor U10544 (N_10544,N_6624,N_7800);
or U10545 (N_10545,N_6187,N_8770);
nand U10546 (N_10546,N_7057,N_7989);
nand U10547 (N_10547,N_7608,N_9767);
nor U10548 (N_10548,N_9939,N_9087);
or U10549 (N_10549,N_9874,N_6659);
nor U10550 (N_10550,N_6557,N_7899);
and U10551 (N_10551,N_6319,N_9929);
and U10552 (N_10552,N_9813,N_6763);
nand U10553 (N_10553,N_9424,N_8296);
or U10554 (N_10554,N_5127,N_9391);
nor U10555 (N_10555,N_8833,N_6945);
nor U10556 (N_10556,N_7829,N_7823);
nand U10557 (N_10557,N_8100,N_9354);
nand U10558 (N_10558,N_8533,N_9973);
nand U10559 (N_10559,N_8321,N_7183);
nand U10560 (N_10560,N_7204,N_5383);
nor U10561 (N_10561,N_8385,N_5586);
nand U10562 (N_10562,N_8415,N_8738);
or U10563 (N_10563,N_8735,N_9685);
or U10564 (N_10564,N_6864,N_6814);
and U10565 (N_10565,N_6544,N_6280);
nor U10566 (N_10566,N_8157,N_8579);
nand U10567 (N_10567,N_8338,N_9362);
nor U10568 (N_10568,N_6715,N_5258);
nor U10569 (N_10569,N_9047,N_8525);
nand U10570 (N_10570,N_7561,N_7330);
and U10571 (N_10571,N_9487,N_9608);
or U10572 (N_10572,N_6843,N_7439);
nand U10573 (N_10573,N_5045,N_9658);
nand U10574 (N_10574,N_5935,N_5995);
or U10575 (N_10575,N_7402,N_8044);
nor U10576 (N_10576,N_6867,N_7118);
or U10577 (N_10577,N_5349,N_7047);
nor U10578 (N_10578,N_6216,N_6308);
and U10579 (N_10579,N_8489,N_8132);
nor U10580 (N_10580,N_6188,N_9235);
nand U10581 (N_10581,N_9103,N_8922);
nor U10582 (N_10582,N_6721,N_5597);
or U10583 (N_10583,N_6026,N_9977);
and U10584 (N_10584,N_7225,N_5163);
and U10585 (N_10585,N_7834,N_6678);
nand U10586 (N_10586,N_8487,N_9208);
and U10587 (N_10587,N_9200,N_8781);
nand U10588 (N_10588,N_8582,N_7945);
and U10589 (N_10589,N_8266,N_6060);
nor U10590 (N_10590,N_8972,N_8286);
nand U10591 (N_10591,N_5360,N_8708);
and U10592 (N_10592,N_7283,N_6555);
nand U10593 (N_10593,N_8567,N_6940);
nor U10594 (N_10594,N_8746,N_9695);
xor U10595 (N_10595,N_7805,N_9012);
nand U10596 (N_10596,N_5649,N_7883);
and U10597 (N_10597,N_8670,N_9280);
or U10598 (N_10598,N_9868,N_9115);
or U10599 (N_10599,N_5348,N_9081);
nand U10600 (N_10600,N_6788,N_9675);
or U10601 (N_10601,N_7028,N_6063);
or U10602 (N_10602,N_5060,N_6222);
and U10603 (N_10603,N_6649,N_6567);
and U10604 (N_10604,N_6190,N_5330);
nand U10605 (N_10605,N_6716,N_6762);
nor U10606 (N_10606,N_7078,N_5416);
nor U10607 (N_10607,N_8811,N_7146);
or U10608 (N_10608,N_7911,N_6588);
nor U10609 (N_10609,N_7695,N_8090);
nand U10610 (N_10610,N_9560,N_8019);
or U10611 (N_10611,N_5278,N_8620);
or U10612 (N_10612,N_5533,N_9331);
nor U10613 (N_10613,N_7432,N_8437);
nand U10614 (N_10614,N_5747,N_5918);
nand U10615 (N_10615,N_6712,N_8680);
nand U10616 (N_10616,N_6519,N_7393);
nor U10617 (N_10617,N_8008,N_5443);
nand U10618 (N_10618,N_9522,N_9224);
and U10619 (N_10619,N_5310,N_8598);
nand U10620 (N_10620,N_9043,N_8457);
nand U10621 (N_10621,N_5615,N_7189);
and U10622 (N_10622,N_9797,N_8737);
nor U10623 (N_10623,N_9635,N_9127);
nor U10624 (N_10624,N_7167,N_9840);
xor U10625 (N_10625,N_7512,N_5357);
nand U10626 (N_10626,N_5992,N_9084);
nand U10627 (N_10627,N_7258,N_9060);
or U10628 (N_10628,N_6916,N_8893);
and U10629 (N_10629,N_8118,N_5856);
and U10630 (N_10630,N_8381,N_8510);
nand U10631 (N_10631,N_5307,N_9573);
or U10632 (N_10632,N_7580,N_6079);
or U10633 (N_10633,N_6951,N_7679);
nor U10634 (N_10634,N_6601,N_7525);
and U10635 (N_10635,N_6182,N_5083);
and U10636 (N_10636,N_6128,N_9739);
nand U10637 (N_10637,N_9924,N_5517);
or U10638 (N_10638,N_7463,N_8164);
and U10639 (N_10639,N_8807,N_6264);
nand U10640 (N_10640,N_8560,N_7270);
and U10641 (N_10641,N_6146,N_8229);
nand U10642 (N_10642,N_9886,N_6540);
nand U10643 (N_10643,N_8933,N_5971);
nor U10644 (N_10644,N_6845,N_8221);
nand U10645 (N_10645,N_6014,N_8734);
or U10646 (N_10646,N_9372,N_9342);
or U10647 (N_10647,N_7500,N_6442);
nand U10648 (N_10648,N_5641,N_7488);
and U10649 (N_10649,N_7498,N_6405);
or U10650 (N_10650,N_6840,N_5255);
nor U10651 (N_10651,N_8750,N_5265);
and U10652 (N_10652,N_9140,N_5825);
and U10653 (N_10653,N_6726,N_9075);
and U10654 (N_10654,N_8600,N_7882);
or U10655 (N_10655,N_5743,N_8465);
nor U10656 (N_10656,N_6915,N_7323);
nand U10657 (N_10657,N_8911,N_7995);
and U10658 (N_10658,N_5648,N_8825);
and U10659 (N_10659,N_7277,N_9545);
or U10660 (N_10660,N_6921,N_6103);
nor U10661 (N_10661,N_5032,N_8996);
or U10662 (N_10662,N_9020,N_8663);
or U10663 (N_10663,N_8596,N_5763);
and U10664 (N_10664,N_6019,N_7755);
or U10665 (N_10665,N_5779,N_8200);
and U10666 (N_10666,N_5675,N_9748);
nand U10667 (N_10667,N_8970,N_5724);
or U10668 (N_10668,N_6623,N_5508);
nand U10669 (N_10669,N_9853,N_5949);
or U10670 (N_10670,N_6610,N_5860);
or U10671 (N_10671,N_5391,N_7184);
and U10672 (N_10672,N_5784,N_8688);
and U10673 (N_10673,N_7974,N_8762);
nor U10674 (N_10674,N_6667,N_6122);
nor U10675 (N_10675,N_9896,N_7521);
nand U10676 (N_10676,N_5429,N_7104);
and U10677 (N_10677,N_6183,N_8854);
nand U10678 (N_10678,N_9266,N_9854);
or U10679 (N_10679,N_8542,N_9758);
and U10680 (N_10680,N_8495,N_5735);
or U10681 (N_10681,N_9191,N_9711);
nor U10682 (N_10682,N_5955,N_5733);
nor U10683 (N_10683,N_5359,N_8026);
nand U10684 (N_10684,N_8160,N_9135);
or U10685 (N_10685,N_6105,N_6313);
or U10686 (N_10686,N_7741,N_8897);
nor U10687 (N_10687,N_6619,N_9555);
and U10688 (N_10688,N_7110,N_9719);
or U10689 (N_10689,N_9513,N_9784);
or U10690 (N_10690,N_9184,N_9837);
xnor U10691 (N_10691,N_9063,N_6212);
and U10692 (N_10692,N_5911,N_8087);
nor U10693 (N_10693,N_5996,N_7897);
and U10694 (N_10694,N_9262,N_6365);
nor U10695 (N_10695,N_5923,N_5064);
or U10696 (N_10696,N_9152,N_5792);
nand U10697 (N_10697,N_8184,N_6317);
nor U10698 (N_10698,N_8012,N_8983);
or U10699 (N_10699,N_8518,N_9291);
nor U10700 (N_10700,N_6310,N_6192);
nor U10701 (N_10701,N_9855,N_9614);
nor U10702 (N_10702,N_6620,N_9124);
or U10703 (N_10703,N_6651,N_6834);
or U10704 (N_10704,N_9204,N_5589);
nand U10705 (N_10705,N_7036,N_7958);
nor U10706 (N_10706,N_5690,N_8482);
or U10707 (N_10707,N_9229,N_8172);
nor U10708 (N_10708,N_8223,N_9336);
and U10709 (N_10709,N_9337,N_6052);
nor U10710 (N_10710,N_6142,N_6071);
nand U10711 (N_10711,N_7045,N_5084);
and U10712 (N_10712,N_9650,N_9187);
nor U10713 (N_10713,N_6598,N_8990);
nor U10714 (N_10714,N_6571,N_8660);
and U10715 (N_10715,N_7164,N_6670);
and U10716 (N_10716,N_9232,N_8010);
nor U10717 (N_10717,N_6061,N_9805);
nor U10718 (N_10718,N_7541,N_6440);
nor U10719 (N_10719,N_6300,N_8250);
or U10720 (N_10720,N_7282,N_9402);
or U10721 (N_10721,N_6022,N_5031);
nand U10722 (N_10722,N_7349,N_5850);
or U10723 (N_10723,N_8043,N_9445);
or U10724 (N_10724,N_6225,N_5807);
nor U10725 (N_10725,N_9665,N_8278);
and U10726 (N_10726,N_9997,N_7670);
nand U10727 (N_10727,N_5156,N_6808);
and U10728 (N_10728,N_8644,N_8886);
nor U10729 (N_10729,N_9822,N_7632);
or U10730 (N_10730,N_7852,N_7170);
or U10731 (N_10731,N_7522,N_9952);
or U10732 (N_10732,N_8627,N_9622);
xor U10733 (N_10733,N_7242,N_8846);
or U10734 (N_10734,N_9466,N_8344);
nor U10735 (N_10735,N_6171,N_6880);
or U10736 (N_10736,N_6538,N_8692);
nand U10737 (N_10737,N_7809,N_6177);
nand U10738 (N_10738,N_8871,N_9538);
and U10739 (N_10739,N_8104,N_6464);
nand U10740 (N_10740,N_6265,N_8190);
nor U10741 (N_10741,N_6474,N_9812);
nand U10742 (N_10742,N_6233,N_6096);
or U10743 (N_10743,N_9895,N_5492);
or U10744 (N_10744,N_7532,N_7723);
nand U10745 (N_10745,N_7053,N_9173);
nor U10746 (N_10746,N_7915,N_8539);
and U10747 (N_10747,N_5248,N_8445);
nand U10748 (N_10748,N_5876,N_5854);
and U10749 (N_10749,N_9537,N_5388);
nor U10750 (N_10750,N_7922,N_8942);
and U10751 (N_10751,N_7904,N_7591);
nand U10752 (N_10752,N_5313,N_7676);
and U10753 (N_10753,N_5179,N_9434);
nand U10754 (N_10754,N_5023,N_5245);
nand U10755 (N_10755,N_6196,N_7493);
nor U10756 (N_10756,N_6160,N_7101);
nor U10757 (N_10757,N_6254,N_7383);
nand U10758 (N_10758,N_7378,N_7685);
and U10759 (N_10759,N_8306,N_6269);
and U10760 (N_10760,N_8939,N_7097);
or U10761 (N_10761,N_8625,N_7788);
nor U10762 (N_10762,N_5959,N_6244);
nand U10763 (N_10763,N_8097,N_6268);
nand U10764 (N_10764,N_7052,N_9968);
or U10765 (N_10765,N_7642,N_6035);
and U10766 (N_10766,N_6781,N_9478);
nor U10767 (N_10767,N_7814,N_7093);
nor U10768 (N_10768,N_6577,N_7971);
or U10769 (N_10769,N_6347,N_9226);
or U10770 (N_10770,N_6112,N_5251);
and U10771 (N_10771,N_7116,N_5671);
nor U10772 (N_10772,N_6042,N_9479);
or U10773 (N_10773,N_7245,N_7732);
nand U10774 (N_10774,N_8887,N_5627);
or U10775 (N_10775,N_8054,N_8764);
nand U10776 (N_10776,N_8599,N_9871);
or U10777 (N_10777,N_5095,N_5053);
nand U10778 (N_10778,N_8453,N_6832);
nor U10779 (N_10779,N_9374,N_8039);
or U10780 (N_10780,N_5981,N_7560);
nor U10781 (N_10781,N_6710,N_7441);
or U10782 (N_10782,N_5948,N_6640);
nor U10783 (N_10783,N_8207,N_5878);
nor U10784 (N_10784,N_5817,N_8696);
or U10785 (N_10785,N_5351,N_9753);
and U10786 (N_10786,N_8103,N_5534);
or U10787 (N_10787,N_7790,N_7856);
nand U10788 (N_10788,N_9870,N_9164);
and U10789 (N_10789,N_5027,N_5845);
and U10790 (N_10790,N_8797,N_8063);
nor U10791 (N_10791,N_8504,N_9351);
nor U10792 (N_10792,N_7766,N_8555);
nor U10793 (N_10793,N_5751,N_5644);
or U10794 (N_10794,N_8853,N_7987);
or U10795 (N_10795,N_6645,N_8455);
nand U10796 (N_10796,N_5706,N_5303);
or U10797 (N_10797,N_9783,N_8399);
nor U10798 (N_10798,N_9334,N_8193);
nor U10799 (N_10799,N_9557,N_5150);
nor U10800 (N_10800,N_9323,N_8745);
or U10801 (N_10801,N_7705,N_8361);
and U10802 (N_10802,N_7029,N_6119);
nor U10803 (N_10803,N_8149,N_5927);
and U10804 (N_10804,N_9432,N_7304);
nand U10805 (N_10805,N_7991,N_5635);
and U10806 (N_10806,N_7775,N_9366);
nand U10807 (N_10807,N_5905,N_5116);
nand U10808 (N_10808,N_7482,N_5120);
or U10809 (N_10809,N_9819,N_6498);
nand U10810 (N_10810,N_6479,N_9706);
nand U10811 (N_10811,N_9543,N_9049);
nor U10812 (N_10812,N_5130,N_6821);
nand U10813 (N_10813,N_8341,N_7051);
nor U10814 (N_10814,N_8881,N_8879);
and U10815 (N_10815,N_7966,N_9716);
nor U10816 (N_10816,N_8892,N_5193);
nand U10817 (N_10817,N_6302,N_8920);
nand U10818 (N_10818,N_9024,N_5107);
or U10819 (N_10819,N_6406,N_9577);
nand U10820 (N_10820,N_6306,N_9771);
nor U10821 (N_10821,N_5821,N_9781);
and U10822 (N_10822,N_6326,N_5714);
nor U10823 (N_10823,N_5409,N_9077);
nand U10824 (N_10824,N_5325,N_9100);
and U10825 (N_10825,N_5889,N_6285);
nor U10826 (N_10826,N_8201,N_5975);
nand U10827 (N_10827,N_5109,N_5174);
nor U10828 (N_10828,N_7776,N_7598);
and U10829 (N_10829,N_9211,N_7397);
and U10830 (N_10830,N_5519,N_7605);
nand U10831 (N_10831,N_6168,N_7645);
nand U10832 (N_10832,N_7131,N_6311);
nand U10833 (N_10833,N_6757,N_6874);
nor U10834 (N_10834,N_5491,N_5538);
nand U10835 (N_10835,N_9238,N_6098);
and U10836 (N_10836,N_8419,N_7893);
or U10837 (N_10837,N_7986,N_9358);
and U10838 (N_10838,N_8975,N_6751);
nor U10839 (N_10839,N_6314,N_9782);
or U10840 (N_10840,N_6672,N_9321);
nand U10841 (N_10841,N_5826,N_7200);
and U10842 (N_10842,N_9455,N_6507);
nand U10843 (N_10843,N_8009,N_9531);
or U10844 (N_10844,N_7162,N_6426);
or U10845 (N_10845,N_7122,N_7126);
nor U10846 (N_10846,N_8431,N_5881);
nand U10847 (N_10847,N_7363,N_8283);
and U10848 (N_10848,N_7861,N_5280);
nor U10849 (N_10849,N_6044,N_6542);
nor U10850 (N_10850,N_9850,N_9568);
or U10851 (N_10851,N_5789,N_7863);
and U10852 (N_10852,N_8496,N_9552);
nand U10853 (N_10853,N_7233,N_5841);
nor U10854 (N_10854,N_9859,N_6013);
and U10855 (N_10855,N_5993,N_6376);
nor U10856 (N_10856,N_5299,N_9897);
nor U10857 (N_10857,N_7354,N_9190);
nand U10858 (N_10858,N_7528,N_8701);
nand U10859 (N_10859,N_7406,N_7652);
nand U10860 (N_10860,N_5169,N_8884);
nor U10861 (N_10861,N_9186,N_7558);
nand U10862 (N_10862,N_7456,N_6730);
nand U10863 (N_10863,N_7272,N_9417);
nand U10864 (N_10864,N_7254,N_9607);
and U10865 (N_10865,N_7179,N_8476);
nor U10866 (N_10866,N_5146,N_9006);
and U10867 (N_10867,N_9335,N_9796);
and U10868 (N_10868,N_8227,N_5373);
or U10869 (N_10869,N_9718,N_5194);
or U10870 (N_10870,N_8929,N_7310);
and U10871 (N_10871,N_8471,N_7191);
nand U10872 (N_10872,N_7426,N_6665);
or U10873 (N_10873,N_9768,N_5514);
nor U10874 (N_10874,N_9011,N_5371);
nand U10875 (N_10875,N_6143,N_6375);
or U10876 (N_10876,N_8095,N_6185);
nand U10877 (N_10877,N_7967,N_8851);
and U10878 (N_10878,N_8513,N_9303);
nand U10879 (N_10879,N_6287,N_6617);
and U10880 (N_10880,N_7317,N_6490);
and U10881 (N_10881,N_7119,N_7460);
nor U10882 (N_10882,N_8375,N_9931);
and U10883 (N_10883,N_7244,N_7497);
and U10884 (N_10884,N_7807,N_5481);
and U10885 (N_10885,N_9745,N_5151);
nand U10886 (N_10886,N_7312,N_8360);
nand U10887 (N_10887,N_6446,N_8407);
and U10888 (N_10888,N_5556,N_5154);
nor U10889 (N_10889,N_9274,N_8429);
nor U10890 (N_10890,N_5124,N_9832);
and U10891 (N_10891,N_6681,N_8067);
and U10892 (N_10892,N_7816,N_5186);
or U10893 (N_10893,N_9267,N_5149);
nor U10894 (N_10894,N_6088,N_7761);
xnor U10895 (N_10895,N_9547,N_9169);
nand U10896 (N_10896,N_5320,N_8517);
nor U10897 (N_10897,N_9378,N_8629);
or U10898 (N_10898,N_9189,N_7748);
nand U10899 (N_10899,N_7350,N_5697);
nor U10900 (N_10900,N_9108,N_9082);
nand U10901 (N_10901,N_8751,N_5182);
or U10902 (N_10902,N_6708,N_5160);
or U10903 (N_10903,N_7346,N_7546);
nand U10904 (N_10904,N_8695,N_6790);
nor U10905 (N_10905,N_5473,N_5776);
or U10906 (N_10906,N_8481,N_6106);
and U10907 (N_10907,N_9941,N_6069);
or U10908 (N_10908,N_7854,N_6541);
nand U10909 (N_10909,N_6303,N_8747);
and U10910 (N_10910,N_7594,N_8177);
or U10911 (N_10911,N_8216,N_5883);
and U10912 (N_10912,N_6625,N_5296);
nor U10913 (N_10913,N_8083,N_8263);
nor U10914 (N_10914,N_7074,N_7874);
and U10915 (N_10915,N_9988,N_9774);
and U10916 (N_10916,N_6456,N_6747);
nand U10917 (N_10917,N_5197,N_8603);
nand U10918 (N_10918,N_8780,N_6537);
nand U10919 (N_10919,N_6799,N_9097);
or U10920 (N_10920,N_7037,N_8739);
nand U10921 (N_10921,N_9523,N_8693);
and U10922 (N_10922,N_8606,N_7020);
nor U10923 (N_10923,N_7906,N_6535);
and U10924 (N_10924,N_6174,N_7217);
and U10925 (N_10925,N_7067,N_6262);
nor U10926 (N_10926,N_9669,N_6437);
nor U10927 (N_10927,N_6669,N_6548);
nor U10928 (N_10928,N_7208,N_5516);
nor U10929 (N_10929,N_9613,N_8965);
nor U10930 (N_10930,N_6158,N_8451);
nor U10931 (N_10931,N_5822,N_9113);
nor U10932 (N_10932,N_5112,N_8096);
nand U10933 (N_10933,N_9824,N_5018);
nor U10934 (N_10934,N_7416,N_6618);
and U10935 (N_10935,N_7399,N_6165);
and U10936 (N_10936,N_8342,N_5270);
nor U10937 (N_10937,N_7884,N_7096);
or U10938 (N_10938,N_8217,N_8562);
xor U10939 (N_10939,N_5058,N_6549);
and U10940 (N_10940,N_5000,N_5722);
and U10941 (N_10941,N_9453,N_7780);
nor U10942 (N_10942,N_5223,N_6690);
and U10943 (N_10943,N_7005,N_7770);
or U10944 (N_10944,N_5686,N_9167);
or U10945 (N_10945,N_9125,N_5387);
nor U10946 (N_10946,N_7662,N_5953);
nand U10947 (N_10947,N_5638,N_6655);
and U10948 (N_10948,N_6993,N_7022);
nor U10949 (N_10949,N_9408,N_6930);
or U10950 (N_10950,N_6969,N_5866);
or U10951 (N_10951,N_7476,N_8937);
or U10952 (N_10952,N_7715,N_6191);
or U10953 (N_10953,N_9054,N_8809);
nor U10954 (N_10954,N_9360,N_6157);
or U10955 (N_10955,N_9093,N_6305);
nand U10956 (N_10956,N_8398,N_9990);
nand U10957 (N_10957,N_6732,N_6648);
and U10958 (N_10958,N_7481,N_8261);
nand U10959 (N_10959,N_6704,N_7081);
nand U10960 (N_10960,N_5670,N_6761);
nor U10961 (N_10961,N_7447,N_7004);
nand U10962 (N_10962,N_7803,N_8550);
nor U10963 (N_10963,N_5322,N_8957);
and U10964 (N_10964,N_5954,N_5660);
or U10965 (N_10965,N_6547,N_7023);
or U10966 (N_10966,N_5382,N_7499);
nand U10967 (N_10967,N_6247,N_8800);
and U10968 (N_10968,N_9258,N_7319);
xnor U10969 (N_10969,N_9227,N_7934);
nor U10970 (N_10970,N_5572,N_7407);
nor U10971 (N_10971,N_5783,N_9017);
or U10972 (N_10972,N_8086,N_7585);
nand U10973 (N_10973,N_8955,N_8271);
nand U10974 (N_10974,N_7177,N_8427);
and U10975 (N_10975,N_8035,N_5090);
nand U10976 (N_10976,N_6502,N_6295);
xnor U10977 (N_10977,N_9736,N_5610);
or U10978 (N_10978,N_5723,N_7916);
nor U10979 (N_10979,N_7213,N_8633);
nand U10980 (N_10980,N_9494,N_9104);
nand U10981 (N_10981,N_5483,N_7106);
or U10982 (N_10982,N_6429,N_9013);
or U10983 (N_10983,N_6942,N_8491);
nor U10984 (N_10984,N_6118,N_5085);
nor U10985 (N_10985,N_8162,N_5157);
or U10986 (N_10986,N_7190,N_6878);
nand U10987 (N_10987,N_8502,N_5873);
and U10988 (N_10988,N_9548,N_6251);
and U10989 (N_10989,N_7366,N_6370);
and U10990 (N_10990,N_5451,N_6273);
and U10991 (N_10991,N_5986,N_7771);
nand U10992 (N_10992,N_5402,N_9373);
nor U10993 (N_10993,N_5645,N_7075);
nand U10994 (N_10994,N_7359,N_7371);
or U10995 (N_10995,N_8219,N_9239);
nor U10996 (N_10996,N_7928,N_6702);
nor U10997 (N_10997,N_6070,N_5830);
nand U10998 (N_10998,N_5114,N_5580);
nand U10999 (N_10999,N_7290,N_6528);
nand U11000 (N_11000,N_9188,N_6378);
nand U11001 (N_11001,N_8085,N_6169);
or U11002 (N_11002,N_9987,N_6922);
or U11003 (N_11003,N_9553,N_8062);
nor U11004 (N_11004,N_6509,N_9831);
or U11005 (N_11005,N_9974,N_7015);
and U11006 (N_11006,N_5281,N_9233);
nor U11007 (N_11007,N_5511,N_9252);
nand U11008 (N_11008,N_8882,N_8426);
nand U11009 (N_11009,N_7931,N_6615);
and U11010 (N_11010,N_5437,N_9646);
or U11011 (N_11011,N_5602,N_6844);
xor U11012 (N_11012,N_8932,N_8483);
and U11013 (N_11013,N_9277,N_6828);
nand U11014 (N_11014,N_6892,N_6654);
nor U11015 (N_11015,N_9441,N_5288);
nor U11016 (N_11016,N_6558,N_8390);
or U11017 (N_11017,N_7665,N_7998);
or U11018 (N_11018,N_8759,N_9246);
nand U11019 (N_11019,N_5522,N_5759);
xnor U11020 (N_11020,N_9025,N_9397);
nand U11021 (N_11021,N_6258,N_9423);
and U11022 (N_11022,N_7762,N_8418);
or U11023 (N_11023,N_8498,N_7739);
and U11024 (N_11024,N_8143,N_7043);
nor U11025 (N_11025,N_8048,N_9371);
nor U11026 (N_11026,N_7949,N_8370);
or U11027 (N_11027,N_9991,N_9022);
nor U11028 (N_11028,N_7427,N_9051);
and U11029 (N_11029,N_6443,N_7872);
and U11030 (N_11030,N_8636,N_5003);
nand U11031 (N_11031,N_7518,N_8553);
nor U11032 (N_11032,N_9559,N_8820);
and U11033 (N_11033,N_5846,N_7930);
or U11034 (N_11034,N_5054,N_5289);
nor U11035 (N_11035,N_9288,N_6616);
nor U11036 (N_11036,N_6420,N_6713);
or U11037 (N_11037,N_5075,N_6899);
nand U11038 (N_11038,N_7513,N_5272);
nor U11039 (N_11039,N_5677,N_6172);
and U11040 (N_11040,N_8991,N_5222);
nand U11041 (N_11041,N_9742,N_6073);
and U11042 (N_11042,N_9147,N_9625);
nand U11043 (N_11043,N_8505,N_9324);
nand U11044 (N_11044,N_9777,N_6576);
or U11045 (N_11045,N_8346,N_8204);
and U11046 (N_11046,N_6778,N_8069);
nor U11047 (N_11047,N_5740,N_5813);
nor U11048 (N_11048,N_9875,N_6830);
and U11049 (N_11049,N_7453,N_9357);
and U11050 (N_11050,N_9276,N_7026);
nand U11051 (N_11051,N_7142,N_7182);
or U11052 (N_11052,N_9959,N_7921);
or U11053 (N_11053,N_7355,N_5695);
nor U11054 (N_11054,N_5001,N_9091);
and U11055 (N_11055,N_8228,N_5122);
nor U11056 (N_11056,N_6613,N_5088);
and U11057 (N_11057,N_7055,N_5015);
nand U11058 (N_11058,N_7121,N_7495);
nor U11059 (N_11059,N_7656,N_8078);
or U11060 (N_11060,N_9370,N_6219);
or U11061 (N_11061,N_7163,N_6741);
and U11062 (N_11062,N_7050,N_5977);
nand U11063 (N_11063,N_7924,N_7573);
nand U11064 (N_11064,N_6745,N_6518);
and U11065 (N_11065,N_5544,N_5606);
and U11066 (N_11066,N_9645,N_8198);
or U11067 (N_11067,N_9861,N_9761);
and U11068 (N_11068,N_9348,N_9884);
and U11069 (N_11069,N_7386,N_5801);
nor U11070 (N_11070,N_5181,N_7630);
nand U11071 (N_11071,N_8729,N_8863);
or U11072 (N_11072,N_6705,N_5715);
nand U11073 (N_11073,N_5568,N_7138);
nand U11074 (N_11074,N_8938,N_8018);
nand U11075 (N_11075,N_9541,N_6927);
and U11076 (N_11076,N_5089,N_5550);
or U11077 (N_11077,N_9490,N_9501);
and U11078 (N_11078,N_5501,N_5688);
or U11079 (N_11079,N_8838,N_5892);
nand U11080 (N_11080,N_6381,N_8408);
or U11081 (N_11081,N_9347,N_8894);
nand U11082 (N_11082,N_9697,N_9446);
nand U11083 (N_11083,N_6948,N_7889);
nor U11084 (N_11084,N_8726,N_7785);
nor U11085 (N_11085,N_8551,N_9483);
or U11086 (N_11086,N_7553,N_6346);
or U11087 (N_11087,N_9852,N_6600);
and U11088 (N_11088,N_6066,N_9183);
or U11089 (N_11089,N_5484,N_7821);
nand U11090 (N_11090,N_9029,N_5891);
or U11091 (N_11091,N_8316,N_5736);
nor U11092 (N_11092,N_7678,N_9802);
and U11093 (N_11093,N_8765,N_5879);
and U11094 (N_11094,N_9016,N_6734);
nor U11095 (N_11095,N_5840,N_9194);
nand U11096 (N_11096,N_5435,N_7309);
and U11097 (N_11097,N_5292,N_7199);
nor U11098 (N_11098,N_8076,N_6099);
or U11099 (N_11099,N_9143,N_7593);
and U11100 (N_11100,N_5549,N_5958);
nor U11101 (N_11101,N_6501,N_8829);
nand U11102 (N_11102,N_5312,N_9591);
nand U11103 (N_11103,N_9708,N_8046);
nand U11104 (N_11104,N_7877,N_6460);
and U11105 (N_11105,N_9616,N_7375);
or U11106 (N_11106,N_8785,N_7917);
nand U11107 (N_11107,N_9449,N_5092);
or U11108 (N_11108,N_5354,N_6824);
nor U11109 (N_11109,N_5138,N_9379);
and U11110 (N_11110,N_7454,N_8186);
xnor U11111 (N_11111,N_9862,N_7461);
nand U11112 (N_11112,N_8852,N_8166);
or U11113 (N_11113,N_6150,N_8621);
or U11114 (N_11114,N_7590,N_6454);
and U11115 (N_11115,N_9214,N_9161);
nand U11116 (N_11116,N_7271,N_6841);
nand U11117 (N_11117,N_9429,N_5906);
nand U11118 (N_11118,N_9014,N_5017);
nand U11119 (N_11119,N_9575,N_8757);
nor U11120 (N_11120,N_9319,N_8014);
nor U11121 (N_11121,N_8168,N_9196);
nor U11122 (N_11122,N_9558,N_9925);
nand U11123 (N_11123,N_5600,N_5823);
and U11124 (N_11124,N_7297,N_9562);
or U11125 (N_11125,N_5934,N_5485);
nand U11126 (N_11126,N_5203,N_9687);
nand U11127 (N_11127,N_6338,N_5262);
nor U11128 (N_11128,N_5022,N_9223);
or U11129 (N_11129,N_6691,N_9296);
and U11130 (N_11130,N_5250,N_5972);
nor U11131 (N_11131,N_6226,N_6410);
or U11132 (N_11132,N_6027,N_5341);
and U11133 (N_11133,N_9707,N_8642);
nor U11134 (N_11134,N_6872,N_7519);
nor U11135 (N_11135,N_7431,N_9508);
nand U11136 (N_11136,N_8108,N_6249);
and U11137 (N_11137,N_8569,N_8135);
nand U11138 (N_11138,N_6204,N_8698);
or U11139 (N_11139,N_9906,N_6911);
and U11140 (N_11140,N_9295,N_7287);
or U11141 (N_11141,N_8170,N_7452);
nand U11142 (N_11142,N_5515,N_5964);
and U11143 (N_11143,N_8450,N_7060);
or U11144 (N_11144,N_6677,N_7294);
nor U11145 (N_11145,N_5973,N_7795);
or U11146 (N_11146,N_5324,N_7822);
nand U11147 (N_11147,N_9305,N_7061);
or U11148 (N_11148,N_8915,N_7256);
and U11149 (N_11149,N_8410,N_6685);
nand U11150 (N_11150,N_7216,N_8662);
nor U11151 (N_11151,N_9068,N_7264);
nor U11152 (N_11152,N_8645,N_9171);
nand U11153 (N_11153,N_7869,N_9869);
nor U11154 (N_11154,N_8068,N_8357);
nor U11155 (N_11155,N_5795,N_7379);
and U11156 (N_11156,N_8327,N_5040);
and U11157 (N_11157,N_6952,N_5766);
and U11158 (N_11158,N_8292,N_5768);
nand U11159 (N_11159,N_9328,N_6766);
nor U11160 (N_11160,N_6432,N_5865);
or U11161 (N_11161,N_5554,N_6956);
and U11162 (N_11162,N_7692,N_6586);
and U11163 (N_11163,N_9001,N_7944);
nor U11164 (N_11164,N_7564,N_9540);
nand U11165 (N_11165,N_6018,N_9603);
and U11166 (N_11166,N_5882,N_5794);
nor U11167 (N_11167,N_6330,N_6466);
nand U11168 (N_11168,N_8401,N_8766);
nand U11169 (N_11169,N_7115,N_5578);
nor U11170 (N_11170,N_5244,N_7677);
or U11171 (N_11171,N_5793,N_8916);
and U11172 (N_11172,N_8371,N_5979);
nor U11173 (N_11173,N_7390,N_6396);
and U11174 (N_11174,N_7251,N_9376);
and U11175 (N_11175,N_9172,N_6272);
nand U11176 (N_11176,N_8209,N_7578);
and U11177 (N_11177,N_7248,N_8775);
and U11178 (N_11178,N_7321,N_5901);
and U11179 (N_11179,N_8007,N_6007);
and U11180 (N_11180,N_5353,N_5165);
and U11181 (N_11181,N_6385,N_7584);
nor U11182 (N_11182,N_6789,N_9254);
nor U11183 (N_11183,N_8231,N_9240);
nor U11184 (N_11184,N_9325,N_6996);
nor U11185 (N_11185,N_5805,N_7011);
nand U11186 (N_11186,N_6318,N_9657);
and U11187 (N_11187,N_7086,N_8608);
and U11188 (N_11188,N_6929,N_5799);
or U11189 (N_11189,N_6587,N_8124);
nand U11190 (N_11190,N_6444,N_8307);
nand U11191 (N_11191,N_9624,N_5335);
nor U11192 (N_11192,N_9873,N_5227);
nor U11193 (N_11193,N_5468,N_7847);
and U11194 (N_11194,N_9995,N_6925);
and U11195 (N_11195,N_6267,N_9454);
nor U11196 (N_11196,N_6435,N_5028);
and U11197 (N_11197,N_7024,N_9520);
and U11198 (N_11198,N_9292,N_9611);
or U11199 (N_11199,N_6015,N_7136);
nand U11200 (N_11200,N_8577,N_6884);
or U11201 (N_11201,N_6215,N_6992);
or U11202 (N_11202,N_9983,N_9023);
and U11203 (N_11203,N_9673,N_8272);
or U11204 (N_11204,N_6827,N_7607);
or U11205 (N_11205,N_6771,N_8685);
nor U11206 (N_11206,N_8022,N_5399);
and U11207 (N_11207,N_8826,N_5025);
nor U11208 (N_11208,N_9867,N_8951);
or U11209 (N_11209,N_7044,N_5131);
nand U11210 (N_11210,N_9592,N_9930);
nor U11211 (N_11211,N_5888,N_6407);
nor U11212 (N_11212,N_6384,N_7234);
nor U11213 (N_11213,N_6281,N_7285);
or U11214 (N_11214,N_6483,N_6737);
or U11215 (N_11215,N_5726,N_6002);
or U11216 (N_11216,N_8441,N_5358);
nand U11217 (N_11217,N_7534,N_8206);
or U11218 (N_11218,N_5132,N_8269);
nor U11219 (N_11219,N_5493,N_9234);
nand U11220 (N_11220,N_9157,N_8033);
nand U11221 (N_11221,N_9810,N_7690);
nand U11222 (N_11222,N_7159,N_6350);
nand U11223 (N_11223,N_9582,N_7132);
nand U11224 (N_11224,N_9976,N_9542);
nand U11225 (N_11225,N_5969,N_8580);
or U11226 (N_11226,N_8930,N_8705);
nor U11227 (N_11227,N_6276,N_8945);
nor U11228 (N_11228,N_6797,N_8659);
and U11229 (N_11229,N_9493,N_7985);
nor U11230 (N_11230,N_9315,N_9444);
nand U11231 (N_11231,N_7601,N_7445);
or U11232 (N_11232,N_8898,N_9420);
nor U11233 (N_11233,N_6032,N_9039);
nand U11234 (N_11234,N_5863,N_7756);
nor U11235 (N_11235,N_9207,N_8081);
and U11236 (N_11236,N_5195,N_5161);
or U11237 (N_11237,N_8109,N_8293);
and U11238 (N_11238,N_9581,N_8257);
nor U11239 (N_11239,N_6516,N_5400);
nand U11240 (N_11240,N_6973,N_5770);
nand U11241 (N_11241,N_9133,N_6452);
nor U11242 (N_11242,N_6946,N_7668);
nor U11243 (N_11243,N_7880,N_9858);
nor U11244 (N_11244,N_5803,N_5445);
and U11245 (N_11245,N_5607,N_6873);
nor U11246 (N_11246,N_7329,N_9318);
nor U11247 (N_11247,N_9953,N_6581);
nand U11248 (N_11248,N_6773,N_5796);
nand U11249 (N_11249,N_5121,N_7133);
nand U11250 (N_11250,N_9058,N_9275);
and U11251 (N_11251,N_6795,N_6979);
and U11252 (N_11252,N_9138,N_7494);
nand U11253 (N_11253,N_5774,N_5368);
or U11254 (N_11254,N_8356,N_6534);
nand U11255 (N_11255,N_5447,N_9564);
and U11256 (N_11256,N_9316,N_6127);
and U11257 (N_11257,N_8810,N_7307);
nand U11258 (N_11258,N_9791,N_9549);
nand U11259 (N_11259,N_9099,N_8466);
or U11260 (N_11260,N_6475,N_9411);
and U11261 (N_11261,N_7400,N_6093);
and U11262 (N_11262,N_5716,N_9554);
or U11263 (N_11263,N_7694,N_9021);
nand U11264 (N_11264,N_5647,N_6316);
nand U11265 (N_11265,N_8707,N_6717);
or U11266 (N_11266,N_9156,N_7604);
xnor U11267 (N_11267,N_6457,N_7804);
nor U11268 (N_11268,N_9814,N_7076);
and U11269 (N_11269,N_6978,N_7700);
or U11270 (N_11270,N_7113,N_8973);
and U11271 (N_11271,N_8910,N_7012);
or U11272 (N_11272,N_9310,N_6161);
or U11273 (N_11273,N_9823,N_7292);
and U11274 (N_11274,N_9762,N_8947);
xor U11275 (N_11275,N_9419,N_9095);
or U11276 (N_11276,N_7318,N_6034);
nor U11277 (N_11277,N_6100,N_6637);
or U11278 (N_11278,N_6366,N_9475);
or U11279 (N_11279,N_5782,N_5717);
or U11280 (N_11280,N_7919,N_5108);
nor U11281 (N_11281,N_9920,N_8755);
and U11282 (N_11282,N_6379,N_8744);
nor U11283 (N_11283,N_6904,N_8060);
or U11284 (N_11284,N_8245,N_8335);
and U11285 (N_11285,N_9008,N_8549);
or U11286 (N_11286,N_7477,N_8376);
or U11287 (N_11287,N_9473,N_7071);
and U11288 (N_11288,N_9298,N_9619);
and U11289 (N_11289,N_7637,N_5159);
and U11290 (N_11290,N_9461,N_9412);
or U11291 (N_11291,N_7862,N_7391);
nand U11292 (N_11292,N_9682,N_6037);
and U11293 (N_11293,N_5833,N_7273);
and U11294 (N_11294,N_8314,N_9972);
and U11295 (N_11295,N_8232,N_5520);
or U11296 (N_11296,N_8348,N_8953);
or U11297 (N_11297,N_5639,N_5898);
nand U11298 (N_11298,N_5700,N_8576);
and U11299 (N_11299,N_5336,N_9170);
and U11300 (N_11300,N_8730,N_7675);
nor U11301 (N_11301,N_5558,N_7025);
or U11302 (N_11302,N_6699,N_6999);
and U11303 (N_11303,N_8666,N_7139);
nand U11304 (N_11304,N_6994,N_9048);
or U11305 (N_11305,N_8736,N_7688);
nand U11306 (N_11306,N_5650,N_6967);
nand U11307 (N_11307,N_9891,N_7006);
nand U11308 (N_11308,N_8837,N_6072);
nand U11309 (N_11309,N_9788,N_8098);
and U11310 (N_11310,N_6561,N_7411);
nand U11311 (N_11311,N_9259,N_7669);
and U11312 (N_11312,N_7237,N_6894);
nor U11313 (N_11313,N_8369,N_6403);
nor U11314 (N_11314,N_9221,N_6500);
nand U11315 (N_11315,N_6622,N_7810);
nand U11316 (N_11316,N_7210,N_9456);
or U11317 (N_11317,N_8860,N_5166);
or U11318 (N_11318,N_8328,N_6582);
and U11319 (N_11319,N_7419,N_7246);
nor U11320 (N_11320,N_8790,N_6291);
nor U11321 (N_11321,N_9071,N_7446);
nand U11322 (N_11322,N_9284,N_9521);
and U11323 (N_11323,N_8425,N_6870);
and U11324 (N_11324,N_8421,N_9472);
nor U11325 (N_11325,N_7710,N_6656);
nor U11326 (N_11326,N_5014,N_5720);
nand U11327 (N_11327,N_8522,N_7910);
and U11328 (N_11328,N_7252,N_6076);
and U11329 (N_11329,N_9003,N_5239);
xor U11330 (N_11330,N_7327,N_5415);
or U11331 (N_11331,N_7909,N_8226);
or U11332 (N_11332,N_6676,N_6724);
or U11333 (N_11333,N_9546,N_9860);
nand U11334 (N_11334,N_8716,N_8883);
or U11335 (N_11335,N_8515,N_6412);
or U11336 (N_11336,N_8287,N_8141);
or U11337 (N_11337,N_7777,N_8535);
nand U11338 (N_11338,N_8962,N_6643);
nor U11339 (N_11339,N_6259,N_5734);
and U11340 (N_11340,N_5323,N_8449);
and U11341 (N_11341,N_6297,N_5579);
and U11342 (N_11342,N_6837,N_8003);
and U11343 (N_11343,N_7858,N_9887);
or U11344 (N_11344,N_7503,N_8927);
or U11345 (N_11345,N_9019,N_7422);
nand U11346 (N_11346,N_7600,N_9763);
or U11347 (N_11347,N_8669,N_5667);
or U11348 (N_11348,N_9121,N_7316);
or U11349 (N_11349,N_7681,N_8836);
nand U11350 (N_11350,N_8584,N_5104);
and U11351 (N_11351,N_6599,N_8769);
nand U11352 (N_11352,N_8684,N_6810);
nand U11353 (N_11353,N_5664,N_5370);
and U11354 (N_11354,N_8637,N_5689);
nand U11355 (N_11355,N_9900,N_7864);
or U11356 (N_11356,N_6123,N_7475);
or U11357 (N_11357,N_8333,N_8001);
xor U11358 (N_11358,N_8926,N_9422);
xor U11359 (N_11359,N_9273,N_5461);
or U11360 (N_11360,N_7920,N_7523);
nand U11361 (N_11361,N_7483,N_5853);
nor U11362 (N_11362,N_9883,N_5989);
and U11363 (N_11363,N_9504,N_7089);
nand U11364 (N_11364,N_6315,N_5828);
or U11365 (N_11365,N_6351,N_6394);
and U11366 (N_11366,N_6632,N_6126);
and U11367 (N_11367,N_8277,N_8061);
nand U11368 (N_11368,N_7959,N_5005);
nand U11369 (N_11369,N_5970,N_8480);
nor U11370 (N_11370,N_8675,N_9980);
and U11371 (N_11371,N_8574,N_8556);
nor U11372 (N_11372,N_8828,N_7471);
or U11373 (N_11373,N_7701,N_9343);
xor U11374 (N_11374,N_6486,N_9339);
nor U11375 (N_11375,N_5681,N_6278);
or U11376 (N_11376,N_6141,N_5960);
and U11377 (N_11377,N_6731,N_6826);
nor U11378 (N_11378,N_6883,N_9747);
and U11379 (N_11379,N_9464,N_5642);
nand U11380 (N_11380,N_7789,N_8423);
nor U11381 (N_11381,N_7635,N_9830);
and U11382 (N_11382,N_5417,N_9312);
nand U11383 (N_11383,N_5093,N_6531);
nor U11384 (N_11384,N_7976,N_5583);
nor U11385 (N_11385,N_8494,N_8358);
nor U11386 (N_11386,N_5594,N_7241);
nand U11387 (N_11387,N_7360,N_7325);
nor U11388 (N_11388,N_6783,N_5535);
nand U11389 (N_11389,N_6391,N_6205);
nor U11390 (N_11390,N_9775,N_5419);
or U11391 (N_11391,N_6074,N_8888);
nor U11392 (N_11392,N_5042,N_5384);
nand U11393 (N_11393,N_8158,N_5542);
or U11394 (N_11394,N_8861,N_8612);
or U11395 (N_11395,N_5537,N_7114);
or U11396 (N_11396,N_6386,N_8372);
nor U11397 (N_11397,N_9743,N_9881);
nor U11398 (N_11398,N_7621,N_5984);
nor U11399 (N_11399,N_5226,N_7428);
and U11400 (N_11400,N_8024,N_8275);
or U11401 (N_11401,N_7876,N_6866);
nand U11402 (N_11402,N_8350,N_5541);
nand U11403 (N_11403,N_7436,N_8767);
and U11404 (N_11404,N_5218,N_6481);
nand U11405 (N_11405,N_9346,N_6725);
nor U11406 (N_11406,N_6886,N_8004);
nor U11407 (N_11407,N_8507,N_5570);
and U11408 (N_11408,N_5939,N_5662);
xor U11409 (N_11409,N_5380,N_8331);
and U11410 (N_11410,N_9440,N_6125);
and U11411 (N_11411,N_8167,N_8312);
nand U11412 (N_11412,N_6928,N_7726);
or U11413 (N_11413,N_5052,N_6058);
or U11414 (N_11414,N_6753,N_7838);
nand U11415 (N_11415,N_9586,N_9388);
and U11416 (N_11416,N_8139,N_6038);
nor U11417 (N_11417,N_7832,N_8679);
and U11418 (N_11418,N_7950,N_8215);
nand U11419 (N_11419,N_7250,N_9476);
nand U11420 (N_11420,N_8700,N_9361);
nand U11421 (N_11421,N_9320,N_6920);
or U11422 (N_11422,N_5957,N_7259);
nor U11423 (N_11423,N_6428,N_8138);
nor U11424 (N_11424,N_9430,N_9950);
nand U11425 (N_11425,N_9509,N_8295);
or U11426 (N_11426,N_7672,N_6606);
xor U11427 (N_11427,N_7176,N_9849);
and U11428 (N_11428,N_8203,N_9530);
and U11429 (N_11429,N_5148,N_7885);
nand U11430 (N_11430,N_9638,N_8564);
nor U11431 (N_11431,N_9894,N_8977);
nor U11432 (N_11432,N_9142,N_7361);
or U11433 (N_11433,N_6232,N_5613);
nand U11434 (N_11434,N_8816,N_7301);
or U11435 (N_11435,N_6298,N_6792);
and U11436 (N_11436,N_6666,N_8979);
nor U11437 (N_11437,N_8420,N_8265);
and U11438 (N_11438,N_7003,N_8436);
and U11439 (N_11439,N_5140,N_7334);
or U11440 (N_11440,N_6323,N_7473);
xnor U11441 (N_11441,N_9231,N_7150);
nor U11442 (N_11442,N_9387,N_6686);
or U11443 (N_11443,N_9804,N_8462);
and U11444 (N_11444,N_7896,N_6765);
and U11445 (N_11445,N_9061,N_6749);
nor U11446 (N_11446,N_9040,N_6355);
and U11447 (N_11447,N_7787,N_7181);
and U11448 (N_11448,N_9112,N_8602);
nor U11449 (N_11449,N_8249,N_6395);
nor U11450 (N_11450,N_7818,N_6156);
nor U11451 (N_11451,N_6589,N_5769);
nand U11452 (N_11452,N_9144,N_6369);
or U11453 (N_11453,N_6091,N_7962);
nand U11454 (N_11454,N_8276,N_7550);
and U11455 (N_11455,N_9193,N_6181);
nor U11456 (N_11456,N_6257,N_9727);
nor U11457 (N_11457,N_6515,N_7574);
nor U11458 (N_11458,N_7423,N_8434);
and U11459 (N_11459,N_9828,N_9863);
and U11460 (N_11460,N_9460,N_7429);
nand U11461 (N_11461,N_7438,N_8214);
or U11462 (N_11462,N_6354,N_8500);
and U11463 (N_11463,N_5167,N_8841);
and U11464 (N_11464,N_5079,N_7736);
nor U11465 (N_11465,N_7320,N_9247);
nand U11466 (N_11466,N_7087,N_7394);
nor U11467 (N_11467,N_8554,N_8332);
nor U11468 (N_11468,N_5637,N_9570);
or U11469 (N_11469,N_6217,N_7127);
nand U11470 (N_11470,N_5201,N_6774);
nor U11471 (N_11471,N_6608,N_7888);
and U11472 (N_11472,N_9064,N_6009);
nand U11473 (N_11473,N_6476,N_9978);
nor U11474 (N_11474,N_7351,N_5256);
and U11475 (N_11475,N_6324,N_7745);
nand U11476 (N_11476,N_8442,N_6197);
nor U11477 (N_11477,N_7666,N_7474);
nor U11478 (N_11478,N_6559,N_5204);
nor U11479 (N_11479,N_9729,N_8187);
and U11480 (N_11480,N_6865,N_8822);
and U11481 (N_11481,N_6849,N_6573);
and U11482 (N_11482,N_9786,N_7588);
and U11483 (N_11483,N_5857,N_5500);
or U11484 (N_11484,N_7719,N_6937);
or U11485 (N_11485,N_6950,N_5601);
nor U11486 (N_11486,N_8152,N_8900);
and U11487 (N_11487,N_9056,N_8531);
nor U11488 (N_11488,N_6238,N_6592);
and U11489 (N_11489,N_6296,N_5366);
or U11490 (N_11490,N_6425,N_5007);
and U11491 (N_11491,N_7894,N_5367);
and U11492 (N_11492,N_9750,N_7699);
or U11493 (N_11493,N_8723,N_8791);
and U11494 (N_11494,N_5013,N_7152);
nor U11495 (N_11495,N_7435,N_9789);
or U11496 (N_11496,N_9359,N_6081);
or U11497 (N_11497,N_8432,N_6343);
and U11498 (N_11498,N_5240,N_5619);
nor U11499 (N_11499,N_5567,N_9525);
or U11500 (N_11500,N_9414,N_9237);
nor U11501 (N_11501,N_5904,N_5375);
nor U11502 (N_11502,N_6696,N_5291);
and U11503 (N_11503,N_8246,N_8709);
nor U11504 (N_11504,N_8448,N_7396);
xor U11505 (N_11505,N_6602,N_5634);
and U11506 (N_11506,N_9598,N_9851);
nor U11507 (N_11507,N_6371,N_6499);
nand U11508 (N_11508,N_6163,N_6647);
nand U11509 (N_11509,N_7802,N_8310);
or U11510 (N_11510,N_7398,N_6461);
or U11511 (N_11511,N_9601,N_8622);
and U11512 (N_11512,N_7073,N_8473);
nand U11513 (N_11513,N_8835,N_6246);
and U11514 (N_11514,N_8148,N_7507);
nor U11515 (N_11515,N_5029,N_5608);
and U11516 (N_11516,N_8687,N_5072);
nor U11517 (N_11517,N_8503,N_9519);
nor U11518 (N_11518,N_5765,N_7960);
and U11519 (N_11519,N_8921,N_7313);
and U11520 (N_11520,N_5321,N_6263);
or U11521 (N_11521,N_9137,N_5460);
or U11522 (N_11522,N_8534,N_5190);
nand U11523 (N_11523,N_5738,N_9760);
nand U11524 (N_11524,N_8126,N_7634);
nor U11525 (N_11525,N_6270,N_9785);
nor U11526 (N_11526,N_6595,N_7261);
or U11527 (N_11527,N_8345,N_9205);
and U11528 (N_11528,N_8301,N_9000);
and U11529 (N_11529,N_9278,N_6149);
nand U11530 (N_11530,N_8830,N_6903);
or U11531 (N_11531,N_7979,N_9116);
and U11532 (N_11532,N_7566,N_8034);
nand U11533 (N_11533,N_5767,N_9664);
nand U11534 (N_11534,N_7778,N_5087);
and U11535 (N_11535,N_8339,N_5630);
and U11536 (N_11536,N_9671,N_6400);
nor U11537 (N_11537,N_5787,N_9015);
nand U11538 (N_11538,N_5011,N_7154);
or U11539 (N_11539,N_8025,N_7721);
nand U11540 (N_11540,N_8992,N_5816);
and U11541 (N_11541,N_5475,N_8568);
xnor U11542 (N_11542,N_5604,N_9947);
or U11543 (N_11543,N_5390,N_9926);
nor U11544 (N_11544,N_8144,N_5571);
and U11545 (N_11545,N_5374,N_9309);
nor U11546 (N_11546,N_9192,N_5742);
nor U11547 (N_11547,N_5073,N_9893);
nor U11548 (N_11548,N_7303,N_6021);
nor U11549 (N_11549,N_7195,N_6871);
and U11550 (N_11550,N_6692,N_7657);
and U11551 (N_11551,N_5196,N_8497);
nand U11552 (N_11552,N_7840,N_7504);
or U11553 (N_11553,N_6133,N_5187);
nor U11554 (N_11554,N_8712,N_8011);
nor U11555 (N_11555,N_7404,N_6439);
nor U11556 (N_11556,N_6290,N_6851);
or U11557 (N_11557,N_8941,N_7120);
or U11558 (N_11558,N_8721,N_8102);
or U11559 (N_11559,N_6822,N_8538);
xnor U11560 (N_11560,N_6662,N_7155);
or U11561 (N_11561,N_9090,N_9561);
and U11562 (N_11562,N_8956,N_8428);
and U11563 (N_11563,N_8368,N_8387);
and U11564 (N_11564,N_7647,N_6329);
nand U11565 (N_11565,N_6784,N_7424);
nor U11566 (N_11566,N_9992,N_7968);
or U11567 (N_11567,N_8676,N_6424);
nand U11568 (N_11568,N_7098,N_6642);
nor U11569 (N_11569,N_8329,N_7489);
or U11570 (N_11570,N_7433,N_6614);
or U11571 (N_11571,N_6628,N_6848);
or U11572 (N_11572,N_8136,N_8074);
nor U11573 (N_11573,N_6727,N_9395);
and U11574 (N_11574,N_7185,N_8710);
and U11575 (N_11575,N_9604,N_7367);
nand U11576 (N_11576,N_9910,N_6839);
and U11577 (N_11577,N_5184,N_6184);
and U11578 (N_11578,N_7088,N_9731);
nor U11579 (N_11579,N_7797,N_7990);
and U11580 (N_11580,N_6458,N_6145);
and U11581 (N_11581,N_7032,N_5401);
and U11582 (N_11582,N_6082,N_6938);
xnor U11583 (N_11583,N_7322,N_5772);
xor U11584 (N_11584,N_5665,N_8234);
xnor U11585 (N_11585,N_8891,N_5999);
nand U11586 (N_11586,N_8258,N_5824);
and U11587 (N_11587,N_7339,N_5207);
nor U11588 (N_11588,N_9369,N_7128);
or U11589 (N_11589,N_7752,N_8844);
and U11590 (N_11590,N_7094,N_7224);
nand U11591 (N_11591,N_7792,N_8330);
or U11592 (N_11592,N_7211,N_6943);
nand U11593 (N_11593,N_7214,N_9641);
nand U11594 (N_11594,N_5055,N_7524);
nand U11595 (N_11595,N_9219,N_8129);
or U11596 (N_11596,N_9876,N_5553);
nand U11597 (N_11597,N_8889,N_7364);
or U11598 (N_11598,N_8378,N_7844);
nand U11599 (N_11599,N_8978,N_9726);
or U11600 (N_11600,N_9094,N_8064);
nand U11601 (N_11601,N_9163,N_6304);
and U11602 (N_11602,N_7516,N_9471);
nand U11603 (N_11603,N_7144,N_8949);
and U11604 (N_11604,N_6152,N_6286);
nand U11605 (N_11605,N_7623,N_5790);
nand U11606 (N_11606,N_9986,N_6380);
nand U11607 (N_11607,N_5505,N_8084);
nand U11608 (N_11608,N_8199,N_8699);
or U11609 (N_11609,N_9073,N_7247);
nor U11610 (N_11610,N_6408,N_5328);
nand U11611 (N_11611,N_9971,N_7286);
or U11612 (N_11612,N_7444,N_6995);
nor U11613 (N_11613,N_5494,N_8508);
or U11614 (N_11614,N_6957,N_8768);
or U11615 (N_11615,N_8365,N_9495);
and U11616 (N_11616,N_8928,N_9210);
nor U11617 (N_11617,N_9462,N_6663);
nand U11618 (N_11618,N_6382,N_8506);
or U11619 (N_11619,N_6633,N_5427);
and U11620 (N_11620,N_5540,N_6053);
or U11621 (N_11621,N_5356,N_8194);
nor U11622 (N_11622,N_6739,N_5721);
nand U11623 (N_11623,N_5311,N_7554);
or U11624 (N_11624,N_8093,N_7440);
nand U11625 (N_11625,N_5172,N_6419);
or U11626 (N_11626,N_9678,N_9002);
and U11627 (N_11627,N_7936,N_8386);
nor U11628 (N_11628,N_9769,N_9469);
and U11629 (N_11629,N_9179,N_8681);
nand U11630 (N_11630,N_6275,N_7465);
nor U11631 (N_11631,N_7964,N_5365);
nor U11632 (N_11632,N_6250,N_8452);
or U11633 (N_11633,N_9151,N_7683);
and U11634 (N_11634,N_6793,N_9821);
and U11635 (N_11635,N_6812,N_9485);
nor U11636 (N_11636,N_8683,N_8847);
nor U11637 (N_11637,N_8463,N_6390);
nand U11638 (N_11638,N_8137,N_6352);
and U11639 (N_11639,N_6974,N_8029);
and U11640 (N_11640,N_6585,N_8632);
or U11641 (N_11641,N_6089,N_8514);
and U11642 (N_11642,N_8005,N_9107);
nor U11643 (N_11643,N_9902,N_7843);
and U11644 (N_11644,N_5943,N_9905);
and U11645 (N_11645,N_6465,N_7484);
nand U11646 (N_11646,N_8673,N_6891);
nor U11647 (N_11647,N_9399,N_5781);
and U11648 (N_11648,N_7583,N_5097);
or U11649 (N_11649,N_9982,N_9301);
nor U11650 (N_11650,N_5275,N_7691);
and U11651 (N_11651,N_6167,N_6511);
nor U11652 (N_11652,N_6193,N_8950);
nor U11653 (N_11653,N_7027,N_8383);
and U11654 (N_11654,N_5997,N_6985);
nor U11655 (N_11655,N_7281,N_8438);
or U11656 (N_11656,N_5691,N_5314);
and U11657 (N_11657,N_8547,N_8389);
or U11658 (N_11658,N_9410,N_9888);
and U11659 (N_11659,N_9437,N_8409);
and U11660 (N_11660,N_6288,N_5424);
and U11661 (N_11661,N_6970,N_8634);
nand U11662 (N_11662,N_8041,N_5012);
nor U11663 (N_11663,N_9329,N_8873);
and U11664 (N_11664,N_7352,N_9877);
nor U11665 (N_11665,N_8151,N_7857);
or U11666 (N_11666,N_7982,N_9647);
nand U11667 (N_11667,N_6972,N_6341);
nor U11668 (N_11668,N_9212,N_7614);
nor U11669 (N_11669,N_5711,N_8874);
and U11670 (N_11670,N_5487,N_6320);
nand U11671 (N_11671,N_8650,N_6569);
nand U11672 (N_11672,N_8808,N_7750);
nand U11673 (N_11673,N_5576,N_6935);
xnor U11674 (N_11674,N_6981,N_7207);
and U11675 (N_11675,N_9963,N_9089);
or U11676 (N_11676,N_8840,N_5036);
or U11677 (N_11677,N_7153,N_7478);
nand U11678 (N_11678,N_7942,N_5318);
nor U11679 (N_11679,N_7786,N_6155);
nor U11680 (N_11680,N_7905,N_9713);
or U11681 (N_11681,N_7240,N_5546);
or U11682 (N_11682,N_5902,N_5725);
or U11683 (N_11683,N_5343,N_9400);
nand U11684 (N_11684,N_9677,N_8901);
and U11685 (N_11685,N_7596,N_6240);
nor U11686 (N_11686,N_8281,N_9272);
or U11687 (N_11687,N_9213,N_8845);
or U11688 (N_11688,N_8251,N_9317);
nand U11689 (N_11689,N_7749,N_6798);
nand U11690 (N_11690,N_8183,N_9932);
or U11691 (N_11691,N_6543,N_8253);
and U11692 (N_11692,N_6818,N_7836);
and U11693 (N_11693,N_6309,N_5591);
and U11694 (N_11694,N_6591,N_5548);
or U11695 (N_11695,N_8611,N_5241);
nand U11696 (N_11696,N_9806,N_8869);
and U11697 (N_11697,N_9477,N_8813);
nand U11698 (N_11698,N_7382,N_7842);
and U11699 (N_11699,N_6772,N_7348);
nor U11700 (N_11700,N_6644,N_8754);
and U11701 (N_11701,N_7267,N_9829);
or U11702 (N_11702,N_6703,N_8964);
nor U11703 (N_11703,N_9435,N_7509);
or U11704 (N_11704,N_6977,N_6680);
or U11705 (N_11705,N_5254,N_6896);
and U11706 (N_11706,N_8320,N_8114);
nor U11707 (N_11707,N_6807,N_6493);
and U11708 (N_11708,N_6447,N_5712);
or U11709 (N_11709,N_9770,N_9938);
nand U11710 (N_11710,N_5661,N_5698);
nor U11711 (N_11711,N_5598,N_9415);
and U11712 (N_11712,N_8057,N_5403);
nor U11713 (N_11713,N_9882,N_6164);
or U11714 (N_11714,N_7017,N_5393);
nor U11715 (N_11715,N_6467,N_7123);
nand U11716 (N_11716,N_9481,N_5868);
or U11717 (N_11717,N_6901,N_7506);
nor U11718 (N_11718,N_9162,N_8211);
and U11719 (N_11719,N_6604,N_5175);
and U11720 (N_11720,N_5050,N_6207);
and U11721 (N_11721,N_9994,N_7759);
nor U11722 (N_11722,N_7430,N_7511);
or U11723 (N_11723,N_7157,N_5171);
or U11724 (N_11724,N_7222,N_5757);
nor U11725 (N_11725,N_6909,N_5754);
or U11726 (N_11726,N_8788,N_6189);
and U11727 (N_11727,N_9649,N_6719);
nor U11728 (N_11728,N_8273,N_8963);
or U11729 (N_11729,N_9333,N_5922);
nand U11730 (N_11730,N_8091,N_9106);
nor U11731 (N_11731,N_5305,N_5797);
or U11732 (N_11732,N_5096,N_8302);
and U11733 (N_11733,N_5143,N_8459);
nor U11734 (N_11734,N_9028,N_8691);
or U11735 (N_11735,N_8512,N_5692);
nor U11736 (N_11736,N_6550,N_9290);
nor U11737 (N_11737,N_6312,N_5407);
or U11738 (N_11738,N_7651,N_6108);
and U11739 (N_11739,N_5897,N_6987);
nor U11740 (N_11740,N_7520,N_7274);
and U11741 (N_11741,N_5872,N_9468);
and U11742 (N_11742,N_7975,N_5618);
nor U11743 (N_11743,N_8319,N_8458);
or U11744 (N_11744,N_5976,N_9636);
or U11745 (N_11745,N_5210,N_9118);
nor U11746 (N_11746,N_6578,N_6353);
and U11747 (N_11747,N_6065,N_5869);
or U11748 (N_11748,N_9709,N_9752);
nand U11749 (N_11749,N_6115,N_6791);
and U11750 (N_11750,N_7033,N_5748);
and U11751 (N_11751,N_8890,N_8925);
nor U11752 (N_11752,N_5009,N_9907);
nor U11753 (N_11753,N_8725,N_6636);
nor U11754 (N_11754,N_8761,N_5951);
or U11755 (N_11755,N_9803,N_9721);
nand U11756 (N_11756,N_9518,N_6590);
nor U11757 (N_11757,N_7344,N_9659);
or U11758 (N_11758,N_8704,N_7955);
or U11759 (N_11759,N_9149,N_8322);
nand U11760 (N_11760,N_6934,N_7819);
nor U11761 (N_11761,N_9730,N_8112);
and U11762 (N_11762,N_6626,N_9215);
and U11763 (N_11763,N_8405,N_7268);
and U11764 (N_11764,N_6638,N_8899);
or U11765 (N_11765,N_7599,N_8859);
nand U11766 (N_11766,N_7817,N_6030);
nor U11767 (N_11767,N_6714,N_8020);
or U11768 (N_11768,N_7218,N_8145);
or U11769 (N_11769,N_9153,N_7713);
nand U11770 (N_11770,N_6520,N_8189);
nor U11771 (N_11771,N_9936,N_7468);
nand U11772 (N_11772,N_7667,N_7873);
nor U11773 (N_11773,N_9652,N_5504);
or U11774 (N_11774,N_6706,N_7107);
and U11775 (N_11775,N_9168,N_7130);
xnor U11776 (N_11776,N_5389,N_9962);
nor U11777 (N_11777,N_9300,N_6862);
xnor U11778 (N_11778,N_5327,N_5760);
nor U11779 (N_11779,N_6919,N_5573);
xnor U11780 (N_11780,N_5562,N_8080);
or U11781 (N_11781,N_5900,N_9688);
nand U11782 (N_11782,N_9847,N_5396);
nor U11783 (N_11783,N_9218,N_6687);
and U11784 (N_11784,N_9672,N_9122);
or U11785 (N_11785,N_6006,N_6170);
nor U11786 (N_11786,N_8179,N_6242);
and U11787 (N_11787,N_6825,N_9878);
nand U11788 (N_11788,N_9139,N_6504);
and U11789 (N_11789,N_8173,N_5530);
or U11790 (N_11790,N_6811,N_7609);
nand U11791 (N_11791,N_9088,N_8191);
nor U11792 (N_11792,N_6441,N_5091);
nor U11793 (N_11793,N_8075,N_7927);
nand U11794 (N_11794,N_9413,N_7954);
or U11795 (N_11795,N_9818,N_8267);
nand U11796 (N_11796,N_6611,N_6890);
and U11797 (N_11797,N_5752,N_5701);
nor U11798 (N_11798,N_7811,N_5274);
nand U11799 (N_11799,N_5946,N_8652);
or U11800 (N_11800,N_6495,N_5676);
and U11801 (N_11801,N_8038,N_5221);
nand U11802 (N_11802,N_6517,N_6779);
or U11803 (N_11803,N_5684,N_5448);
nand U11804 (N_11804,N_6253,N_9728);
nor U11805 (N_11805,N_7926,N_5129);
and U11806 (N_11806,N_9901,N_5575);
or U11807 (N_11807,N_7582,N_7293);
nand U11808 (N_11808,N_9528,N_7221);
and U11809 (N_11809,N_5477,N_6817);
and U11810 (N_11810,N_6564,N_5051);
nor U11811 (N_11811,N_7659,N_9610);
and U11812 (N_11812,N_9617,N_7718);
nor U11813 (N_11813,N_9486,N_7219);
nand U11814 (N_11814,N_5884,N_7205);
and U11815 (N_11815,N_7655,N_5215);
or U11816 (N_11816,N_5413,N_9935);
or U11817 (N_11817,N_8027,N_8748);
and U11818 (N_11818,N_6682,N_7794);
and U11819 (N_11819,N_9263,N_8181);
nand U11820 (N_11820,N_6819,N_7526);
or U11821 (N_11821,N_7851,N_9590);
or U11822 (N_11822,N_9511,N_5952);
nor U11823 (N_11823,N_9352,N_9176);
or U11824 (N_11824,N_6842,N_7932);
and U11825 (N_11825,N_9999,N_6332);
and U11826 (N_11826,N_8954,N_5105);
nor U11827 (N_11827,N_7328,N_6526);
nor U11828 (N_11828,N_8931,N_8315);
or U11829 (N_11829,N_9160,N_8050);
and U11830 (N_11830,N_9981,N_9326);
nand U11831 (N_11831,N_9961,N_8147);
nor U11832 (N_11832,N_5582,N_7188);
and U11833 (N_11833,N_5837,N_8896);
nand U11834 (N_11834,N_9689,N_5656);
and U11835 (N_11835,N_8902,N_7039);
or U11836 (N_11836,N_7450,N_5276);
and U11837 (N_11837,N_7340,N_7697);
and U11838 (N_11838,N_6574,N_5209);
and U11839 (N_11839,N_5188,N_8544);
and U11840 (N_11840,N_6087,N_6804);
nand U11841 (N_11841,N_7542,N_7243);
nand U11842 (N_11842,N_6770,N_7686);
nor U11843 (N_11843,N_7636,N_6218);
nand U11844 (N_11844,N_6545,N_5260);
nor U11845 (N_11845,N_9220,N_8786);
or U11846 (N_11846,N_8300,N_9260);
nor U11847 (N_11847,N_6401,N_8850);
nand U11848 (N_11848,N_7567,N_7783);
and U11849 (N_11849,N_6939,N_6051);
or U11850 (N_11850,N_5332,N_6307);
and U11851 (N_11851,N_8875,N_8993);
nor U11852 (N_11852,N_9101,N_7062);
and U11853 (N_11853,N_8868,N_6237);
or U11854 (N_11854,N_9919,N_5585);
or U11855 (N_11855,N_9261,N_5643);
nor U11856 (N_11856,N_5936,N_7830);
nor U11857 (N_11857,N_5653,N_5547);
and U11858 (N_11858,N_7171,N_8180);
or U11859 (N_11859,N_6525,N_7848);
nor U11860 (N_11860,N_5277,N_6986);
xnor U11861 (N_11861,N_7754,N_6409);
nor U11862 (N_11862,N_5145,N_8918);
nor U11863 (N_11863,N_9380,N_7773);
nand U11864 (N_11864,N_9764,N_9383);
and U11865 (N_11865,N_5410,N_9332);
and U11866 (N_11866,N_7706,N_7671);
and U11867 (N_11867,N_6236,N_5066);
or U11868 (N_11868,N_5625,N_6603);
or U11869 (N_11869,N_9640,N_9866);
or U11870 (N_11870,N_9349,N_9474);
nand U11871 (N_11871,N_5624,N_6229);
and U11872 (N_11872,N_5944,N_7744);
and U11873 (N_11873,N_5940,N_9597);
nand U11874 (N_11874,N_7812,N_6339);
nand U11875 (N_11875,N_6965,N_6679);
and U11876 (N_11876,N_9642,N_8238);
nor U11877 (N_11877,N_8908,N_6430);
nor U11878 (N_11878,N_6875,N_9442);
nor U11879 (N_11879,N_8059,N_9966);
or U11880 (N_11880,N_6856,N_7235);
nand U11881 (N_11881,N_7193,N_8237);
and U11882 (N_11882,N_5394,N_9165);
or U11883 (N_11883,N_9327,N_7765);
nand U11884 (N_11884,N_9216,N_6468);
and U11885 (N_11885,N_8661,N_5704);
or U11886 (N_11886,N_8827,N_6780);
nand U11887 (N_11887,N_5363,N_5372);
nand U11888 (N_11888,N_8842,N_7923);
or U11889 (N_11889,N_7712,N_8524);
nand U11890 (N_11890,N_9356,N_9500);
nor U11891 (N_11891,N_9458,N_6552);
and U11892 (N_11892,N_8128,N_6658);
or U11893 (N_11893,N_5086,N_8724);
and U11894 (N_11894,N_6723,N_5125);
xor U11895 (N_11895,N_8079,N_7654);
or U11896 (N_11896,N_9242,N_9923);
nor U11897 (N_11897,N_9034,N_9070);
and U11898 (N_11898,N_9431,N_5513);
and U11899 (N_11899,N_7231,N_7160);
or U11900 (N_11900,N_7326,N_7009);
nand U11901 (N_11901,N_7527,N_7622);
nor U11902 (N_11902,N_6388,N_5046);
nand U11903 (N_11903,N_7865,N_8313);
nand U11904 (N_11904,N_8849,N_6539);
nand U11905 (N_11905,N_9197,N_9908);
xor U11906 (N_11906,N_9199,N_5078);
or U11907 (N_11907,N_5152,N_5355);
nand U11908 (N_11908,N_5191,N_8581);
or U11909 (N_11909,N_9596,N_8188);
and U11910 (N_11910,N_7306,N_6084);
nand U11911 (N_11911,N_9780,N_5899);
or U11912 (N_11912,N_9457,N_9271);
nand U11913 (N_11913,N_7230,N_9660);
nand U11914 (N_11914,N_5798,N_6621);
nand U11915 (N_11915,N_8030,N_5392);
nand U11916 (N_11916,N_5441,N_6046);
or U11917 (N_11917,N_9954,N_5208);
nor U11918 (N_11918,N_6756,N_5755);
or U11919 (N_11919,N_5503,N_6492);
or U11920 (N_11920,N_5710,N_7260);
nor U11921 (N_11921,N_6131,N_9046);
or U11922 (N_11922,N_9694,N_5233);
or U11923 (N_11923,N_5651,N_6932);
nand U11924 (N_11924,N_5243,N_6016);
nor U11925 (N_11925,N_7925,N_7409);
or U11926 (N_11926,N_7729,N_5614);
nand U11927 (N_11927,N_5543,N_9612);
and U11928 (N_11928,N_9195,N_9912);
nor U11929 (N_11929,N_9516,N_5920);
or U11930 (N_11930,N_7969,N_8367);
nand U11931 (N_11931,N_9772,N_7129);
nand U11932 (N_11932,N_6491,N_9632);
and U11933 (N_11933,N_6231,N_9644);
nor U11934 (N_11934,N_9958,N_6971);
nor U11935 (N_11935,N_8115,N_7165);
and U11936 (N_11936,N_9032,N_8587);
or U11937 (N_11937,N_7269,N_6433);
and U11938 (N_11938,N_7458,N_7742);
nand U11939 (N_11939,N_7879,N_7059);
or U11940 (N_11940,N_6450,N_5886);
nor U11941 (N_11941,N_9450,N_7980);
and U11942 (N_11942,N_5470,N_8176);
nand U11943 (N_11943,N_6823,N_5293);
nand U11944 (N_11944,N_9109,N_6010);
or U11945 (N_11945,N_9497,N_6998);
or U11946 (N_11946,N_9079,N_9667);
nand U11947 (N_11947,N_7353,N_7825);
and U11948 (N_11948,N_9588,N_8366);
and U11949 (N_11949,N_8353,N_6085);
or U11950 (N_11950,N_5286,N_6831);
or U11951 (N_11951,N_6040,N_5439);
or U11952 (N_11952,N_9969,N_5786);
or U11953 (N_11953,N_9563,N_7956);
nor U11954 (N_11954,N_9793,N_8792);
and U11955 (N_11955,N_8784,N_6477);
nand U11956 (N_11956,N_5596,N_5446);
and U11957 (N_11957,N_6068,N_7134);
nand U11958 (N_11958,N_6266,N_8521);
nand U11959 (N_11959,N_7860,N_6506);
nor U11960 (N_11960,N_6277,N_7641);
and U11961 (N_11961,N_6775,N_8804);
nand U11962 (N_11962,N_5669,N_5827);
nor U11963 (N_11963,N_7368,N_8831);
nor U11964 (N_11964,N_7314,N_6854);
and U11965 (N_11965,N_8444,N_7533);
or U11966 (N_11966,N_7220,N_5895);
and U11967 (N_11967,N_6208,N_8783);
or U11968 (N_11968,N_7871,N_9975);
and U11969 (N_11969,N_7362,N_9055);
nand U11970 (N_11970,N_8880,N_9340);
or U11971 (N_11971,N_8968,N_8906);
and U11972 (N_11972,N_7180,N_6399);
nand U11973 (N_11973,N_5235,N_9921);
and U11974 (N_11974,N_7151,N_5802);
and U11975 (N_11975,N_6358,N_9686);
or U11976 (N_11976,N_7933,N_5731);
and U11977 (N_11977,N_5919,N_7769);
nand U11978 (N_11978,N_7203,N_8864);
nor U11979 (N_11979,N_9698,N_5694);
nand U11980 (N_11980,N_5308,N_5559);
or U11981 (N_11981,N_9180,N_7849);
or U11982 (N_11982,N_9690,N_6090);
nor U11983 (N_11983,N_5762,N_5819);
and U11984 (N_11984,N_8105,N_8248);
and U11985 (N_11985,N_8440,N_5985);
nand U11986 (N_11986,N_8752,N_9230);
or U11987 (N_11987,N_6024,N_5836);
nor U11988 (N_11988,N_8913,N_6367);
and U11989 (N_11989,N_8056,N_5219);
or U11990 (N_11990,N_8559,N_6889);
nand U11991 (N_11991,N_7935,N_5903);
nand U11992 (N_11992,N_6700,N_8501);
nor U11993 (N_11993,N_8593,N_9074);
or U11994 (N_11994,N_5696,N_6086);
or U11995 (N_11995,N_8605,N_8140);
and U11996 (N_11996,N_9134,N_9470);
nand U11997 (N_11997,N_8406,N_5098);
nand U11998 (N_11998,N_5398,N_7957);
nor U11999 (N_11999,N_5016,N_9626);
or U12000 (N_12000,N_8182,N_9256);
and U12001 (N_12001,N_9217,N_9062);
nand U12002 (N_12002,N_6077,N_9885);
xnor U12003 (N_12003,N_8304,N_6720);
nor U12004 (N_12004,N_7077,N_7619);
nand U12005 (N_12005,N_7737,N_5657);
nor U12006 (N_12006,N_8430,N_8291);
nand U12007 (N_12007,N_6116,N_8174);
or U12008 (N_12008,N_9314,N_8649);
nand U12009 (N_12009,N_8120,N_9065);
and U12010 (N_12010,N_5455,N_7149);
nor U12011 (N_12011,N_7943,N_6983);
or U12012 (N_12012,N_7875,N_7387);
nand U12013 (N_12013,N_7492,N_7065);
or U12014 (N_12014,N_5523,N_7412);
or U12015 (N_12015,N_6107,N_8912);
xor U12016 (N_12016,N_7784,N_9631);
and U12017 (N_12017,N_8284,N_5237);
or U12018 (N_12018,N_8526,N_8677);
nand U12019 (N_12019,N_6279,N_7835);
and U12020 (N_12020,N_5907,N_5202);
nor U12021 (N_12021,N_9128,N_8546);
nand U12022 (N_12022,N_8355,N_5266);
or U12023 (N_12023,N_5924,N_8446);
and U12024 (N_12024,N_8987,N_8545);
nor U12025 (N_12025,N_8731,N_6299);
and U12026 (N_12026,N_5082,N_8464);
or U12027 (N_12027,N_6863,N_7161);
and U12028 (N_12028,N_6785,N_5785);
or U12029 (N_12029,N_6758,N_6554);
and U12030 (N_12030,N_6760,N_7951);
nand U12031 (N_12031,N_9605,N_6947);
or U12032 (N_12032,N_7175,N_6887);
and U12033 (N_12033,N_9389,N_5560);
nand U12034 (N_12034,N_6260,N_7202);
and U12035 (N_12035,N_5153,N_8142);
and U12036 (N_12036,N_7664,N_8653);
nor U12037 (N_12037,N_8814,N_8858);
nand U12038 (N_12038,N_6210,N_9825);
and U12039 (N_12039,N_5352,N_7315);
and U12040 (N_12040,N_7640,N_7758);
nor U12041 (N_12041,N_5966,N_9589);
nor U12042 (N_12042,N_7280,N_8610);
and U12043 (N_12043,N_5080,N_9996);
nor U12044 (N_12044,N_6414,N_5963);
nand U12045 (N_12045,N_8411,N_8909);
nor U12046 (N_12046,N_8667,N_5457);
nor U12047 (N_12047,N_7058,N_9670);
nand U12048 (N_12048,N_5229,N_6701);
nand U12049 (N_12049,N_9766,N_7442);
or U12050 (N_12050,N_6221,N_8924);
nor U12051 (N_12051,N_8999,N_5369);
and U12052 (N_12052,N_8760,N_6497);
nor U12053 (N_12053,N_9732,N_5913);
or U12054 (N_12054,N_8782,N_6565);
nor U12055 (N_12055,N_7781,N_7965);
nor U12056 (N_12056,N_6711,N_6936);
and U12057 (N_12057,N_6562,N_5909);
or U12058 (N_12058,N_6223,N_8210);
xor U12059 (N_12059,N_6976,N_5620);
nand U12060 (N_12060,N_7929,N_9856);
nor U12061 (N_12061,N_9287,N_5041);
nor U12062 (N_12062,N_9390,N_9524);
nand U12063 (N_12063,N_5340,N_8326);
and U12064 (N_12064,N_6389,N_5465);
and U12065 (N_12065,N_9438,N_6459);
nand U12066 (N_12066,N_6914,N_5930);
nand U12067 (N_12067,N_7650,N_7209);
and U12068 (N_12068,N_7472,N_9269);
and U12069 (N_12069,N_9244,N_7663);
nand U12070 (N_12070,N_9421,N_7014);
and U12071 (N_12071,N_9620,N_8297);
nor U12072 (N_12072,N_7035,N_7648);
nor U12073 (N_12073,N_7937,N_5683);
nor U12074 (N_12074,N_5885,N_7343);
nor U12075 (N_12075,N_6630,N_7332);
and U12076 (N_12076,N_7725,N_5315);
or U12077 (N_12077,N_9281,N_7617);
nand U12078 (N_12078,N_7469,N_5462);
or U12079 (N_12079,N_5756,N_8212);
and U12080 (N_12080,N_9621,N_7716);
nand U12081 (N_12081,N_5707,N_7413);
nand U12082 (N_12082,N_8154,N_6104);
or U12083 (N_12083,N_5851,N_5155);
and U12084 (N_12084,N_5896,N_6631);
or U12085 (N_12085,N_6417,N_7616);
nand U12086 (N_12086,N_8607,N_8280);
nand U12087 (N_12087,N_5862,N_5687);
and U12088 (N_12088,N_9283,N_7082);
nor U12089 (N_12089,N_5739,N_6134);
or U12090 (N_12090,N_8094,N_7186);
or U12091 (N_12091,N_6835,N_7702);
nand U12092 (N_12092,N_6478,N_5838);
nand U12093 (N_12093,N_8821,N_5577);
nor U12094 (N_12094,N_5814,N_5791);
and U12095 (N_12095,N_5067,N_7610);
or U12096 (N_12096,N_8058,N_7253);
nand U12097 (N_12097,N_8776,N_5471);
or U12098 (N_12098,N_8474,N_9293);
nor U12099 (N_12099,N_6607,N_9498);
nor U12100 (N_12100,N_7449,N_5301);
and U12101 (N_12101,N_5750,N_8740);
nand U12102 (N_12102,N_6117,N_6855);
nor U12103 (N_12103,N_9661,N_8718);
nor U12104 (N_12104,N_7768,N_6422);
nand U12105 (N_12105,N_7999,N_8614);
or U12106 (N_12106,N_7908,N_5418);
nand U12107 (N_12107,N_5430,N_7703);
xor U12108 (N_12108,N_5478,N_8877);
and U12109 (N_12109,N_8794,N_9928);
nor U12110 (N_12110,N_8392,N_9609);
and U12111 (N_12111,N_8848,N_9489);
nor U12112 (N_12112,N_5937,N_8958);
and U12113 (N_12113,N_9915,N_7559);
and U12114 (N_12114,N_7845,N_9341);
nor U12115 (N_12115,N_5039,N_6524);
nor U12116 (N_12116,N_6553,N_7746);
and U12117 (N_12117,N_8113,N_6377);
nand U12118 (N_12118,N_8966,N_6697);
nor U12119 (N_12119,N_6097,N_8374);
and U12120 (N_12120,N_6209,N_5469);
and U12121 (N_12121,N_6055,N_8959);
and U12122 (N_12122,N_8952,N_7866);
and U12123 (N_12123,N_7000,N_8998);
and U12124 (N_12124,N_7018,N_5049);
and U12125 (N_12125,N_9633,N_5561);
and U12126 (N_12126,N_8318,N_8213);
nor U12127 (N_12127,N_8631,N_6470);
nor U12128 (N_12128,N_5408,N_8609);
or U12129 (N_12129,N_5496,N_6462);
xnor U12130 (N_12130,N_5912,N_8870);
nor U12131 (N_12131,N_7563,N_7064);
or U12132 (N_12132,N_8163,N_9426);
or U12133 (N_12133,N_6512,N_5133);
and U12134 (N_12134,N_6689,N_7178);
nor U12135 (N_12135,N_9759,N_9889);
nor U12136 (N_12136,N_9085,N_6646);
or U12137 (N_12137,N_8540,N_8422);
and U12138 (N_12138,N_8548,N_7479);
or U12139 (N_12139,N_7808,N_5062);
and U12140 (N_12140,N_9710,N_8298);
nand U12141 (N_12141,N_5626,N_5737);
or U12142 (N_12142,N_5259,N_8678);
and U12143 (N_12143,N_7727,N_6364);
nor U12144 (N_12144,N_5414,N_7278);
nor U12145 (N_12145,N_7717,N_5178);
and U12146 (N_12146,N_8948,N_7415);
and U12147 (N_12147,N_7682,N_9833);
nand U12148 (N_12148,N_7070,N_7457);
and U12149 (N_12149,N_7236,N_8325);
and U12150 (N_12150,N_9517,N_6958);
nor U12151 (N_12151,N_6200,N_6510);
and U12152 (N_12152,N_9536,N_8866);
nor U12153 (N_12153,N_6047,N_8111);
nor U12154 (N_12154,N_6121,N_6563);
and U12155 (N_12155,N_8509,N_8976);
nor U12156 (N_12156,N_8254,N_9253);
or U12157 (N_12157,N_5117,N_6530);
nor U12158 (N_12158,N_5362,N_9534);
nand U12159 (N_12159,N_8488,N_5300);
or U12160 (N_12160,N_9203,N_6186);
nor U12161 (N_12161,N_5057,N_9105);
and U12162 (N_12162,N_8728,N_5059);
nand U12163 (N_12163,N_7016,N_6629);
nor U12164 (N_12164,N_5588,N_8895);
and U12165 (N_12165,N_8202,N_7174);
nor U12166 (N_12166,N_9637,N_7311);
nand U12167 (N_12167,N_8997,N_9377);
nor U12168 (N_12168,N_7587,N_5709);
and U12169 (N_12169,N_9367,N_5775);
nand U12170 (N_12170,N_5928,N_8000);
nor U12171 (N_12171,N_7198,N_8818);
and U12172 (N_12172,N_7586,N_5574);
nand U12173 (N_12173,N_6344,N_6220);
nand U12174 (N_12174,N_6434,N_9282);
nand U12175 (N_12175,N_8274,N_9834);
and U12176 (N_12176,N_8682,N_9185);
nor U12177 (N_12177,N_7158,N_9393);
nand U12178 (N_12178,N_7046,N_9398);
nor U12179 (N_12179,N_8037,N_8686);
nor U12180 (N_12180,N_6029,N_5199);
and U12181 (N_12181,N_8391,N_6743);
or U12182 (N_12182,N_6482,N_9571);
and U12183 (N_12183,N_7618,N_5118);
nand U12184 (N_12184,N_6847,N_5268);
and U12185 (N_12185,N_5980,N_7597);
nor U12186 (N_12186,N_5261,N_8101);
or U12187 (N_12187,N_5252,N_7019);
nor U12188 (N_12188,N_7868,N_9756);
nand U12189 (N_12189,N_8373,N_9158);
and U12190 (N_12190,N_5474,N_5206);
or U12191 (N_12191,N_9502,N_6413);
or U12192 (N_12192,N_8107,N_8116);
nor U12193 (N_12193,N_9579,N_7168);
or U12194 (N_12194,N_7764,N_8264);
or U12195 (N_12195,N_5238,N_6360);
or U12196 (N_12196,N_6898,N_7395);
and U12197 (N_12197,N_7156,N_8876);
nor U12198 (N_12198,N_5679,N_9740);
nand U12199 (N_12199,N_7041,N_8485);
nor U12200 (N_12200,N_6256,N_5808);
and U12201 (N_12201,N_6876,N_7201);
and U12202 (N_12202,N_8066,N_8165);
or U12203 (N_12203,N_8714,N_6803);
nor U12204 (N_12204,N_7972,N_9879);
nand U12205 (N_12205,N_5870,N_5965);
nor U12206 (N_12206,N_9304,N_9209);
or U12207 (N_12207,N_9243,N_7606);
nand U12208 (N_12208,N_8638,N_7839);
nor U12209 (N_12209,N_9057,N_7117);
nand U12210 (N_12210,N_8985,N_8719);
nand U12211 (N_12211,N_8532,N_7530);
nor U12212 (N_12212,N_8578,N_8561);
and U12213 (N_12213,N_8563,N_5395);
nand U12214 (N_12214,N_5674,N_8447);
and U12215 (N_12215,N_6154,N_5663);
nor U12216 (N_12216,N_6359,N_6829);
and U12217 (N_12217,N_7013,N_9313);
or U12218 (N_12218,N_9594,N_6572);
or U12219 (N_12219,N_6261,N_6605);
nand U12220 (N_12220,N_8787,N_8643);
nand U12221 (N_12221,N_7798,N_7891);
and U12222 (N_12222,N_8697,N_8468);
and U12223 (N_12223,N_9042,N_8252);
or U12224 (N_12224,N_7417,N_7337);
nor U12225 (N_12225,N_5871,N_7263);
nor U12226 (N_12226,N_6964,N_5103);
and U12227 (N_12227,N_6333,N_6372);
nor U12228 (N_12228,N_6328,N_8255);
nand U12229 (N_12229,N_7961,N_6140);
or U12230 (N_12230,N_5106,N_6111);
or U12231 (N_12231,N_9078,N_6431);
nor U12232 (N_12232,N_6235,N_5968);
or U12233 (N_12233,N_5646,N_5346);
nor U12234 (N_12234,N_6398,N_9368);
nor U12235 (N_12235,N_6227,N_6913);
or U12236 (N_12236,N_9712,N_8774);
or U12237 (N_12237,N_7779,N_9757);
nor U12238 (N_12238,N_5859,N_8192);
and U12239 (N_12239,N_5685,N_6869);
nor U12240 (N_12240,N_5967,N_8566);
or U12241 (N_12241,N_9765,N_8583);
or U12242 (N_12242,N_8308,N_6641);
nand U12243 (N_12243,N_9702,N_5139);
nor U12244 (N_12244,N_6397,N_6488);
and U12245 (N_12245,N_6532,N_6368);
nand U12246 (N_12246,N_5529,N_8640);
nand U12247 (N_12247,N_8065,N_8195);
and U12248 (N_12248,N_9787,N_5294);
nand U12249 (N_12249,N_8363,N_5818);
nor U12250 (N_12250,N_8527,N_7486);
and U12251 (N_12251,N_7806,N_7308);
and U12252 (N_12252,N_8240,N_8703);
nand U12253 (N_12253,N_7595,N_8795);
and U12254 (N_12254,N_6356,N_6815);
or U12255 (N_12255,N_6203,N_7680);
or U12256 (N_12256,N_6113,N_6522);
or U12257 (N_12257,N_5433,N_6487);
nor U12258 (N_12258,N_8303,N_8657);
nand U12259 (N_12259,N_8354,N_6496);
nand U12260 (N_12260,N_9285,N_8758);
or U12261 (N_12261,N_9005,N_9206);
or U12262 (N_12262,N_9045,N_8236);
nand U12263 (N_12263,N_8815,N_8031);
nand U12264 (N_12264,N_9257,N_6733);
and U12265 (N_12265,N_8259,N_6301);
nand U12266 (N_12266,N_8523,N_6556);
nand U12267 (N_12267,N_6327,N_7381);
nor U12268 (N_12268,N_9225,N_8558);
or U12269 (N_12269,N_5423,N_6695);
nand U12270 (N_12270,N_9198,N_7684);
nor U12271 (N_12271,N_6661,N_7837);
and U12272 (N_12272,N_9059,N_5379);
or U12273 (N_12273,N_6292,N_8904);
or U12274 (N_12274,N_7262,N_5319);
nor U12275 (N_12275,N_8665,N_7711);
nand U12276 (N_12276,N_5381,N_8772);
nor U12277 (N_12277,N_8490,N_9703);
nor U12278 (N_12278,N_8243,N_8052);
nand U12279 (N_12279,N_9801,N_5874);
and U12280 (N_12280,N_8919,N_8260);
nand U12281 (N_12281,N_6011,N_5069);
or U12282 (N_12282,N_5987,N_5094);
and U12283 (N_12283,N_8672,N_7448);
nand U12284 (N_12284,N_9957,N_8336);
and U12285 (N_12285,N_8706,N_7249);
xnor U12286 (N_12286,N_6806,N_6879);
nand U12287 (N_12287,N_8073,N_5741);
nand U12288 (N_12288,N_9903,N_7238);
or U12289 (N_12289,N_5858,N_7571);
nand U12290 (N_12290,N_6718,N_8655);
nor U12291 (N_12291,N_6787,N_7342);
nor U12292 (N_12292,N_8402,N_5956);
or U12293 (N_12293,N_7846,N_6674);
nor U12294 (N_12294,N_9096,N_9330);
or U12295 (N_12295,N_9018,N_7345);
and U12296 (N_12296,N_6201,N_9496);
or U12297 (N_12297,N_7196,N_9662);
nand U12298 (N_12298,N_8946,N_5509);
nand U12299 (N_12299,N_7722,N_9268);
and U12300 (N_12300,N_8641,N_8169);
or U12301 (N_12301,N_6031,N_7467);
or U12302 (N_12302,N_6933,N_9639);
nor U12303 (N_12303,N_8379,N_7535);
nand U12304 (N_12304,N_7265,N_9241);
nand U12305 (N_12305,N_8400,N_7385);
or U12306 (N_12306,N_6918,N_8969);
nor U12307 (N_12307,N_5463,N_6736);
or U12308 (N_12308,N_6404,N_9723);
or U12309 (N_12309,N_9447,N_8591);
or U12310 (N_12310,N_7988,N_7576);
and U12311 (N_12311,N_5162,N_5295);
and U12312 (N_12312,N_9705,N_6335);
nand U12313 (N_12313,N_5076,N_7288);
and U12314 (N_12314,N_9492,N_5914);
and U12315 (N_12315,N_6906,N_5342);
or U12316 (N_12316,N_5298,N_9566);
or U12317 (N_12317,N_5019,N_7627);
or U12318 (N_12318,N_9381,N_5290);
and U12319 (N_12319,N_7275,N_9126);
or U12320 (N_12320,N_6912,N_9459);
or U12321 (N_12321,N_5498,N_7850);
nor U12322 (N_12322,N_6147,N_7063);
nor U12323 (N_12323,N_9311,N_8674);
nand U12324 (N_12324,N_6941,N_9425);
nand U12325 (N_12325,N_9514,N_9302);
and U12326 (N_12326,N_9799,N_9279);
or U12327 (N_12327,N_9201,N_5552);
nor U12328 (N_12328,N_5672,N_9776);
or U12329 (N_12329,N_7040,N_5991);
and U12330 (N_12330,N_9010,N_6453);
nor U12331 (N_12331,N_8311,N_7341);
nor U12332 (N_12332,N_7031,N_9448);
or U12333 (N_12333,N_7095,N_5947);
nand U12334 (N_12334,N_5844,N_7380);
nor U12335 (N_12335,N_6331,N_6742);
nor U12336 (N_12336,N_5843,N_5164);
or U12337 (N_12337,N_5564,N_7137);
and U12338 (N_12338,N_8588,N_5137);
or U12339 (N_12339,N_7707,N_8134);
and U12340 (N_12340,N_5231,N_5815);
nor U12341 (N_12341,N_8002,N_8171);
nor U12342 (N_12342,N_6885,N_9922);
nand U12343 (N_12343,N_9674,N_8053);
and U12344 (N_12344,N_7226,N_8624);
and U12345 (N_12345,N_7940,N_9648);
and U12346 (N_12346,N_6449,N_7589);
nand U12347 (N_12347,N_8382,N_6584);
and U12348 (N_12348,N_6012,N_7279);
and U12349 (N_12349,N_5110,N_9696);
nand U12350 (N_12350,N_6050,N_7517);
nand U12351 (N_12351,N_9844,N_6039);
and U12352 (N_12352,N_9933,N_6782);
nor U12353 (N_12353,N_6198,N_7543);
nand U12354 (N_12354,N_7638,N_7038);
or U12355 (N_12355,N_7480,N_5136);
and U12356 (N_12356,N_8352,N_8156);
or U12357 (N_12357,N_8021,N_6438);
nand U12358 (N_12358,N_8989,N_6095);
nand U12359 (N_12359,N_7338,N_7577);
nand U12360 (N_12360,N_7010,N_6418);
or U12361 (N_12361,N_9322,N_7102);
or U12362 (N_12362,N_5345,N_7042);
and U12363 (N_12363,N_5021,N_7502);
nand U12364 (N_12364,N_9580,N_7212);
or U12365 (N_12365,N_7169,N_9527);
or U12366 (N_12366,N_9076,N_6334);
xor U12367 (N_12367,N_5518,N_5566);
nand U12368 (N_12368,N_9155,N_5910);
or U12369 (N_12369,N_9792,N_6961);
nand U12370 (N_12370,N_5746,N_5829);
nor U12371 (N_12371,N_5185,N_5283);
or U12372 (N_12372,N_8839,N_9467);
or U12373 (N_12373,N_8130,N_8586);
and U12374 (N_12374,N_7069,N_9086);
or U12375 (N_12375,N_8573,N_7997);
nand U12376 (N_12376,N_5043,N_7827);
or U12377 (N_12377,N_6245,N_6402);
nor U12378 (N_12378,N_7496,N_7299);
or U12379 (N_12379,N_5480,N_6955);
and U12380 (N_12380,N_7109,N_7734);
and U12381 (N_12381,N_7459,N_9353);
nand U12382 (N_12382,N_9807,N_5287);
nand U12383 (N_12383,N_8960,N_5812);
nand U12384 (N_12384,N_7487,N_6448);
nor U12385 (N_12385,N_6566,N_8529);
and U12386 (N_12386,N_8006,N_9749);
nor U12387 (N_12387,N_7613,N_8439);
or U12388 (N_12388,N_8070,N_6336);
nand U12389 (N_12389,N_6580,N_6020);
or U12390 (N_12390,N_9129,N_5411);
and U12391 (N_12391,N_8885,N_9286);
or U12392 (N_12392,N_9704,N_6166);
nor U12393 (N_12393,N_6568,N_6838);
nor U12394 (N_12394,N_6794,N_5242);
nand U12395 (N_12395,N_5334,N_9544);
nand U12396 (N_12396,N_6694,N_9503);
nand U12397 (N_12397,N_6982,N_5753);
nand U12398 (N_12398,N_8324,N_6387);
and U12399 (N_12399,N_8317,N_7147);
or U12400 (N_12400,N_5264,N_7007);
and U12401 (N_12401,N_8413,N_6138);
nand U12402 (N_12402,N_6472,N_5961);
nor U12403 (N_12403,N_7295,N_9599);
nor U12404 (N_12404,N_5990,N_6023);
and U12405 (N_12405,N_5925,N_6092);
nor U12406 (N_12406,N_5406,N_6729);
nor U12407 (N_12407,N_6513,N_7565);
nor U12408 (N_12408,N_6374,N_7403);
or U12409 (N_12409,N_5778,N_6707);
or U12410 (N_12410,N_8934,N_5565);
or U12411 (N_12411,N_8323,N_9836);
nand U12412 (N_12412,N_9676,N_5047);
and U12413 (N_12413,N_9053,N_6234);
nand U12414 (N_12414,N_5820,N_9463);
or U12415 (N_12415,N_5654,N_8595);
nand U12416 (N_12416,N_8604,N_5337);
nor U12417 (N_12417,N_5887,N_9405);
or U12418 (N_12418,N_9416,N_8812);
nor U12419 (N_12419,N_7090,N_8416);
and U12420 (N_12420,N_7735,N_6748);
nand U12421 (N_12421,N_5499,N_7405);
or U12422 (N_12422,N_5002,N_6521);
and U12423 (N_12423,N_8412,N_8282);
nor U12424 (N_12424,N_5877,N_8713);
nand U12425 (N_12425,N_5632,N_9507);
or U12426 (N_12426,N_7531,N_6325);
nand U12427 (N_12427,N_6062,N_9600);
or U12428 (N_12428,N_9842,N_5458);
or U12429 (N_12429,N_7994,N_9249);
nand U12430 (N_12430,N_7490,N_9578);
nand U12431 (N_12431,N_8435,N_9845);
or U12432 (N_12432,N_6759,N_5037);
and U12433 (N_12433,N_7841,N_7255);
nand U12434 (N_12434,N_5581,N_5170);
and U12435 (N_12435,N_5026,N_8040);
xnor U12436 (N_12436,N_7728,N_8690);
nor U12437 (N_12437,N_8982,N_9734);
and U12438 (N_12438,N_5917,N_5198);
nand U12439 (N_12439,N_9236,N_6451);
or U12440 (N_12440,N_5347,N_7625);
nor U12441 (N_12441,N_7358,N_7693);
nand U12442 (N_12442,N_5269,N_5183);
nor U12443 (N_12443,N_9404,N_7501);
or U12444 (N_12444,N_8777,N_7853);
nand U12445 (N_12445,N_8364,N_9815);
or U12446 (N_12446,N_9583,N_7552);
nor U12447 (N_12447,N_6132,N_6102);
nand U12448 (N_12448,N_7978,N_7815);
and U12449 (N_12449,N_8362,N_7791);
nand U12450 (N_12450,N_5338,N_7763);
nand U12451 (N_12451,N_8856,N_9606);
nand U12452 (N_12452,N_9092,N_5024);
nor U12453 (N_12453,N_6162,N_6926);
nor U12454 (N_12454,N_7021,N_8799);
nor U12455 (N_12455,N_7421,N_9403);
and U12456 (N_12456,N_7733,N_5926);
or U12457 (N_12457,N_7336,N_5236);
nand U12458 (N_12458,N_8995,N_6813);
and U12459 (N_12459,N_7420,N_9773);
or U12460 (N_12460,N_5595,N_5699);
nand U12461 (N_12461,N_7206,N_5061);
nand U12462 (N_12462,N_7401,N_8270);
nand U12463 (N_12463,N_8340,N_9030);
nand U12464 (N_12464,N_8122,N_8051);
nor U12465 (N_12465,N_6124,N_8618);
nand U12466 (N_12466,N_7544,N_9439);
nand U12467 (N_12467,N_6908,N_6489);
nor U12468 (N_12468,N_5180,N_9120);
nand U12469 (N_12469,N_7799,N_5680);
nand U12470 (N_12470,N_8865,N_7757);
nand U12471 (N_12471,N_6129,N_6698);
xor U12472 (N_12472,N_9794,N_5852);
and U12473 (N_12473,N_5758,N_6750);
or U12474 (N_12474,N_5655,N_7973);
nor U12475 (N_12475,N_7324,N_8045);
nand U12476 (N_12476,N_7658,N_9556);
nand U12477 (N_12477,N_7602,N_7300);
nand U12478 (N_12478,N_7491,N_8185);
nor U12479 (N_12479,N_7335,N_9565);
or U12480 (N_12480,N_5842,N_6392);
nand U12481 (N_12481,N_8424,N_9222);
or U12482 (N_12482,N_9067,N_8616);
and U12483 (N_12483,N_7084,N_9506);
nor U12484 (N_12484,N_7772,N_8806);
nor U12485 (N_12485,N_5230,N_5048);
nor U12486 (N_12486,N_7056,N_9083);
and U12487 (N_12487,N_9159,N_5702);
nand U12488 (N_12488,N_8862,N_9864);
nor U12489 (N_12489,N_7724,N_7740);
xor U12490 (N_12490,N_7782,N_5636);
and U12491 (N_12491,N_6683,N_5378);
or U12492 (N_12492,N_8575,N_8867);
and U12493 (N_12493,N_5128,N_5102);
and U12494 (N_12494,N_7030,N_5809);
nor U12495 (N_12495,N_5894,N_5880);
and U12496 (N_12496,N_5432,N_5931);
or U12497 (N_12497,N_7660,N_5497);
and U12498 (N_12498,N_5479,N_7377);
nor U12499 (N_12499,N_7751,N_9297);
or U12500 (N_12500,N_9791,N_7868);
or U12501 (N_12501,N_8565,N_9175);
nand U12502 (N_12502,N_7142,N_9196);
nand U12503 (N_12503,N_6929,N_5669);
nand U12504 (N_12504,N_5354,N_9590);
nor U12505 (N_12505,N_7477,N_8377);
nor U12506 (N_12506,N_7177,N_6169);
and U12507 (N_12507,N_5865,N_8685);
or U12508 (N_12508,N_9277,N_9084);
nand U12509 (N_12509,N_5461,N_5264);
or U12510 (N_12510,N_6761,N_8733);
nand U12511 (N_12511,N_7216,N_8236);
nand U12512 (N_12512,N_5892,N_8612);
or U12513 (N_12513,N_5601,N_8299);
nand U12514 (N_12514,N_9553,N_5723);
and U12515 (N_12515,N_6310,N_6375);
and U12516 (N_12516,N_6761,N_5793);
nor U12517 (N_12517,N_7956,N_7993);
or U12518 (N_12518,N_7066,N_9324);
nor U12519 (N_12519,N_6529,N_9102);
or U12520 (N_12520,N_5773,N_8210);
or U12521 (N_12521,N_8211,N_7240);
nor U12522 (N_12522,N_7955,N_9360);
and U12523 (N_12523,N_7717,N_7333);
and U12524 (N_12524,N_5343,N_5631);
and U12525 (N_12525,N_9465,N_7338);
nor U12526 (N_12526,N_7158,N_6417);
nor U12527 (N_12527,N_8267,N_6171);
nand U12528 (N_12528,N_6121,N_9620);
and U12529 (N_12529,N_9067,N_5882);
and U12530 (N_12530,N_9435,N_6994);
or U12531 (N_12531,N_5843,N_8366);
and U12532 (N_12532,N_9596,N_7558);
and U12533 (N_12533,N_9728,N_5830);
nand U12534 (N_12534,N_6652,N_6308);
nand U12535 (N_12535,N_5753,N_7304);
or U12536 (N_12536,N_6817,N_5720);
nor U12537 (N_12537,N_9163,N_6246);
nand U12538 (N_12538,N_6174,N_6722);
nor U12539 (N_12539,N_7216,N_9847);
and U12540 (N_12540,N_5204,N_6896);
nor U12541 (N_12541,N_8238,N_8594);
nor U12542 (N_12542,N_6138,N_6710);
nor U12543 (N_12543,N_9796,N_9042);
nand U12544 (N_12544,N_9018,N_7025);
nand U12545 (N_12545,N_9313,N_8351);
and U12546 (N_12546,N_8497,N_9043);
or U12547 (N_12547,N_5729,N_5010);
nand U12548 (N_12548,N_7509,N_5257);
nand U12549 (N_12549,N_6323,N_5208);
nand U12550 (N_12550,N_7535,N_9352);
and U12551 (N_12551,N_9532,N_7437);
nand U12552 (N_12552,N_8914,N_8581);
nor U12553 (N_12553,N_5366,N_7306);
or U12554 (N_12554,N_6021,N_9215);
or U12555 (N_12555,N_5588,N_8602);
or U12556 (N_12556,N_5190,N_6136);
nor U12557 (N_12557,N_8296,N_5806);
nand U12558 (N_12558,N_6035,N_8102);
nand U12559 (N_12559,N_9797,N_6023);
nor U12560 (N_12560,N_8346,N_9542);
or U12561 (N_12561,N_9757,N_7289);
nand U12562 (N_12562,N_8516,N_8233);
and U12563 (N_12563,N_7621,N_5777);
nor U12564 (N_12564,N_7447,N_8993);
nand U12565 (N_12565,N_6094,N_8022);
nand U12566 (N_12566,N_6403,N_5155);
or U12567 (N_12567,N_7655,N_6802);
nor U12568 (N_12568,N_9758,N_7056);
nor U12569 (N_12569,N_5292,N_8917);
or U12570 (N_12570,N_5754,N_6205);
and U12571 (N_12571,N_6871,N_7712);
nand U12572 (N_12572,N_8905,N_9995);
and U12573 (N_12573,N_6874,N_8779);
nand U12574 (N_12574,N_5658,N_8705);
nand U12575 (N_12575,N_9425,N_7443);
nand U12576 (N_12576,N_9429,N_9956);
nor U12577 (N_12577,N_9994,N_6142);
and U12578 (N_12578,N_5688,N_6501);
and U12579 (N_12579,N_9469,N_8341);
and U12580 (N_12580,N_6616,N_6337);
and U12581 (N_12581,N_9944,N_9741);
or U12582 (N_12582,N_9482,N_9953);
nor U12583 (N_12583,N_6500,N_8595);
nor U12584 (N_12584,N_5828,N_8861);
and U12585 (N_12585,N_8246,N_5581);
nand U12586 (N_12586,N_5071,N_7834);
nand U12587 (N_12587,N_8699,N_5088);
or U12588 (N_12588,N_8425,N_6948);
or U12589 (N_12589,N_7017,N_6745);
nor U12590 (N_12590,N_9750,N_6919);
nor U12591 (N_12591,N_7110,N_9658);
and U12592 (N_12592,N_5781,N_5632);
or U12593 (N_12593,N_6489,N_9567);
or U12594 (N_12594,N_9099,N_5554);
nand U12595 (N_12595,N_6116,N_8230);
or U12596 (N_12596,N_8328,N_5236);
nor U12597 (N_12597,N_5844,N_6825);
or U12598 (N_12598,N_8684,N_7333);
or U12599 (N_12599,N_7299,N_7315);
and U12600 (N_12600,N_9052,N_7140);
and U12601 (N_12601,N_9157,N_6362);
nor U12602 (N_12602,N_6592,N_6992);
or U12603 (N_12603,N_5854,N_6110);
nand U12604 (N_12604,N_5683,N_9934);
xnor U12605 (N_12605,N_8703,N_5200);
nor U12606 (N_12606,N_5031,N_5605);
nand U12607 (N_12607,N_5957,N_9873);
and U12608 (N_12608,N_8192,N_8397);
nand U12609 (N_12609,N_6422,N_5209);
nor U12610 (N_12610,N_5234,N_9459);
nand U12611 (N_12611,N_8326,N_9006);
or U12612 (N_12612,N_8625,N_9032);
nor U12613 (N_12613,N_9240,N_8559);
nor U12614 (N_12614,N_9259,N_7045);
or U12615 (N_12615,N_7138,N_5574);
nand U12616 (N_12616,N_6882,N_8952);
nand U12617 (N_12617,N_8538,N_5971);
nor U12618 (N_12618,N_9102,N_8195);
or U12619 (N_12619,N_9792,N_5455);
and U12620 (N_12620,N_9466,N_7058);
and U12621 (N_12621,N_7289,N_7779);
and U12622 (N_12622,N_5331,N_8903);
nand U12623 (N_12623,N_5835,N_9424);
nand U12624 (N_12624,N_6125,N_9285);
nand U12625 (N_12625,N_7563,N_6924);
and U12626 (N_12626,N_8715,N_9243);
nor U12627 (N_12627,N_9855,N_7019);
nor U12628 (N_12628,N_6338,N_8101);
or U12629 (N_12629,N_7715,N_7983);
or U12630 (N_12630,N_7753,N_9064);
and U12631 (N_12631,N_5692,N_9316);
and U12632 (N_12632,N_6019,N_9537);
nand U12633 (N_12633,N_7991,N_9766);
or U12634 (N_12634,N_7256,N_6191);
or U12635 (N_12635,N_8999,N_6786);
nor U12636 (N_12636,N_5420,N_7490);
and U12637 (N_12637,N_9926,N_9633);
nor U12638 (N_12638,N_5167,N_6454);
or U12639 (N_12639,N_5232,N_8715);
nor U12640 (N_12640,N_8591,N_7186);
nor U12641 (N_12641,N_9509,N_5346);
nor U12642 (N_12642,N_5566,N_9540);
and U12643 (N_12643,N_6736,N_5344);
and U12644 (N_12644,N_8928,N_8343);
nor U12645 (N_12645,N_6127,N_8006);
xor U12646 (N_12646,N_6362,N_8235);
and U12647 (N_12647,N_8818,N_9610);
or U12648 (N_12648,N_8248,N_6843);
or U12649 (N_12649,N_6293,N_5527);
or U12650 (N_12650,N_7821,N_6474);
nor U12651 (N_12651,N_7431,N_9768);
or U12652 (N_12652,N_6113,N_7264);
nand U12653 (N_12653,N_9468,N_8498);
and U12654 (N_12654,N_8787,N_8963);
nand U12655 (N_12655,N_7649,N_7254);
nand U12656 (N_12656,N_5831,N_9674);
nand U12657 (N_12657,N_5577,N_7147);
and U12658 (N_12658,N_9207,N_5352);
or U12659 (N_12659,N_5082,N_8538);
xnor U12660 (N_12660,N_7846,N_9850);
or U12661 (N_12661,N_5478,N_9379);
nand U12662 (N_12662,N_6272,N_7009);
and U12663 (N_12663,N_5942,N_6140);
nor U12664 (N_12664,N_9529,N_6616);
and U12665 (N_12665,N_5973,N_9293);
nor U12666 (N_12666,N_5772,N_7989);
or U12667 (N_12667,N_8986,N_8141);
and U12668 (N_12668,N_7172,N_9761);
or U12669 (N_12669,N_6966,N_5512);
nand U12670 (N_12670,N_5203,N_7165);
nor U12671 (N_12671,N_5657,N_5509);
and U12672 (N_12672,N_9719,N_5510);
nor U12673 (N_12673,N_7153,N_5214);
or U12674 (N_12674,N_6625,N_7051);
nor U12675 (N_12675,N_9221,N_6222);
or U12676 (N_12676,N_6401,N_9733);
and U12677 (N_12677,N_9090,N_7435);
nand U12678 (N_12678,N_7564,N_7421);
nand U12679 (N_12679,N_8364,N_9019);
nor U12680 (N_12680,N_7497,N_6817);
and U12681 (N_12681,N_7963,N_9506);
or U12682 (N_12682,N_5878,N_5636);
and U12683 (N_12683,N_5135,N_5208);
nand U12684 (N_12684,N_7084,N_9154);
nor U12685 (N_12685,N_9122,N_6022);
or U12686 (N_12686,N_7783,N_9164);
nor U12687 (N_12687,N_9644,N_9194);
nand U12688 (N_12688,N_8532,N_8536);
and U12689 (N_12689,N_8485,N_5356);
or U12690 (N_12690,N_7825,N_6013);
nor U12691 (N_12691,N_5838,N_5784);
or U12692 (N_12692,N_6239,N_7413);
xnor U12693 (N_12693,N_6394,N_5213);
and U12694 (N_12694,N_6141,N_6208);
nor U12695 (N_12695,N_9716,N_6522);
nand U12696 (N_12696,N_9831,N_7274);
or U12697 (N_12697,N_5208,N_7438);
nand U12698 (N_12698,N_5635,N_7355);
and U12699 (N_12699,N_8017,N_7528);
and U12700 (N_12700,N_6899,N_7568);
nor U12701 (N_12701,N_5761,N_7903);
or U12702 (N_12702,N_6974,N_7473);
and U12703 (N_12703,N_8416,N_5942);
nand U12704 (N_12704,N_9641,N_5002);
or U12705 (N_12705,N_9179,N_7599);
or U12706 (N_12706,N_7025,N_8378);
and U12707 (N_12707,N_5147,N_9293);
and U12708 (N_12708,N_9536,N_9025);
nor U12709 (N_12709,N_6615,N_8271);
nor U12710 (N_12710,N_8134,N_6658);
or U12711 (N_12711,N_5436,N_8437);
nor U12712 (N_12712,N_5042,N_6385);
nand U12713 (N_12713,N_7735,N_5890);
nor U12714 (N_12714,N_8807,N_5246);
and U12715 (N_12715,N_6723,N_7560);
nor U12716 (N_12716,N_6723,N_5876);
and U12717 (N_12717,N_9600,N_9918);
nor U12718 (N_12718,N_5314,N_5647);
and U12719 (N_12719,N_5170,N_7079);
nand U12720 (N_12720,N_7697,N_5735);
or U12721 (N_12721,N_8040,N_8258);
nand U12722 (N_12722,N_7900,N_7582);
nand U12723 (N_12723,N_9667,N_6876);
nor U12724 (N_12724,N_9611,N_6783);
and U12725 (N_12725,N_8873,N_6313);
and U12726 (N_12726,N_9402,N_5423);
and U12727 (N_12727,N_7160,N_6722);
nor U12728 (N_12728,N_9051,N_5206);
and U12729 (N_12729,N_9760,N_5657);
and U12730 (N_12730,N_7788,N_5340);
nand U12731 (N_12731,N_5832,N_7347);
and U12732 (N_12732,N_5690,N_5855);
nor U12733 (N_12733,N_6324,N_5493);
nor U12734 (N_12734,N_8153,N_5930);
or U12735 (N_12735,N_5356,N_6298);
nand U12736 (N_12736,N_7405,N_6655);
nor U12737 (N_12737,N_7601,N_6456);
and U12738 (N_12738,N_5177,N_7418);
and U12739 (N_12739,N_7157,N_7673);
and U12740 (N_12740,N_6242,N_8222);
or U12741 (N_12741,N_9812,N_5958);
and U12742 (N_12742,N_9380,N_9543);
or U12743 (N_12743,N_9649,N_7416);
nand U12744 (N_12744,N_6585,N_6902);
nand U12745 (N_12745,N_5958,N_6683);
or U12746 (N_12746,N_8003,N_6143);
nor U12747 (N_12747,N_5335,N_8253);
or U12748 (N_12748,N_5340,N_8990);
nor U12749 (N_12749,N_6819,N_8095);
and U12750 (N_12750,N_8191,N_8839);
nand U12751 (N_12751,N_5072,N_8542);
nand U12752 (N_12752,N_6965,N_9430);
and U12753 (N_12753,N_8409,N_9819);
and U12754 (N_12754,N_5930,N_9471);
and U12755 (N_12755,N_9147,N_8698);
nand U12756 (N_12756,N_6570,N_6352);
nand U12757 (N_12757,N_6620,N_6871);
nor U12758 (N_12758,N_8905,N_8997);
or U12759 (N_12759,N_6936,N_5533);
and U12760 (N_12760,N_6957,N_7327);
nand U12761 (N_12761,N_9876,N_5367);
and U12762 (N_12762,N_5449,N_8282);
or U12763 (N_12763,N_8509,N_7186);
or U12764 (N_12764,N_7860,N_9229);
nand U12765 (N_12765,N_6934,N_5375);
or U12766 (N_12766,N_8262,N_9435);
and U12767 (N_12767,N_5887,N_8163);
nor U12768 (N_12768,N_7771,N_7509);
nand U12769 (N_12769,N_7789,N_9949);
nand U12770 (N_12770,N_7333,N_5071);
and U12771 (N_12771,N_6486,N_5642);
and U12772 (N_12772,N_6788,N_6748);
and U12773 (N_12773,N_6236,N_9566);
xnor U12774 (N_12774,N_9550,N_7827);
xnor U12775 (N_12775,N_6662,N_9536);
and U12776 (N_12776,N_7029,N_8465);
and U12777 (N_12777,N_7623,N_6171);
or U12778 (N_12778,N_9553,N_5550);
and U12779 (N_12779,N_7616,N_6207);
and U12780 (N_12780,N_9590,N_8988);
nor U12781 (N_12781,N_6354,N_7564);
nand U12782 (N_12782,N_5055,N_5324);
nor U12783 (N_12783,N_8494,N_5757);
nor U12784 (N_12784,N_5177,N_7085);
nand U12785 (N_12785,N_9549,N_8334);
nor U12786 (N_12786,N_8087,N_9298);
or U12787 (N_12787,N_7956,N_8677);
nor U12788 (N_12788,N_5514,N_6791);
nand U12789 (N_12789,N_6136,N_9035);
and U12790 (N_12790,N_5309,N_7532);
or U12791 (N_12791,N_9854,N_5070);
or U12792 (N_12792,N_8638,N_7844);
or U12793 (N_12793,N_8567,N_9603);
nand U12794 (N_12794,N_7223,N_8331);
and U12795 (N_12795,N_5996,N_8473);
and U12796 (N_12796,N_6564,N_7288);
and U12797 (N_12797,N_7751,N_9121);
and U12798 (N_12798,N_8916,N_7554);
nor U12799 (N_12799,N_5182,N_6579);
or U12800 (N_12800,N_8418,N_8382);
nor U12801 (N_12801,N_7836,N_5184);
nand U12802 (N_12802,N_9938,N_8182);
or U12803 (N_12803,N_7772,N_5998);
and U12804 (N_12804,N_7494,N_6523);
and U12805 (N_12805,N_7336,N_7562);
nor U12806 (N_12806,N_9309,N_9582);
and U12807 (N_12807,N_5303,N_9478);
nand U12808 (N_12808,N_5485,N_6886);
or U12809 (N_12809,N_6670,N_6789);
nor U12810 (N_12810,N_5401,N_9914);
or U12811 (N_12811,N_6472,N_8967);
and U12812 (N_12812,N_7845,N_7689);
and U12813 (N_12813,N_7715,N_6261);
nor U12814 (N_12814,N_5694,N_5705);
nor U12815 (N_12815,N_7308,N_8099);
nand U12816 (N_12816,N_9427,N_6262);
or U12817 (N_12817,N_6470,N_8491);
nor U12818 (N_12818,N_9520,N_6519);
nand U12819 (N_12819,N_6938,N_7803);
nor U12820 (N_12820,N_9792,N_9681);
or U12821 (N_12821,N_8559,N_7292);
or U12822 (N_12822,N_7061,N_9011);
and U12823 (N_12823,N_8106,N_5570);
or U12824 (N_12824,N_5811,N_8542);
nand U12825 (N_12825,N_7710,N_5975);
and U12826 (N_12826,N_7487,N_7949);
nor U12827 (N_12827,N_9274,N_9074);
nor U12828 (N_12828,N_8261,N_5877);
or U12829 (N_12829,N_6283,N_7018);
nor U12830 (N_12830,N_6389,N_7282);
nand U12831 (N_12831,N_5337,N_9809);
xor U12832 (N_12832,N_7296,N_7922);
and U12833 (N_12833,N_7202,N_7108);
nor U12834 (N_12834,N_9235,N_9720);
and U12835 (N_12835,N_9276,N_9056);
nor U12836 (N_12836,N_6370,N_9066);
nor U12837 (N_12837,N_5870,N_6061);
nand U12838 (N_12838,N_6425,N_8937);
nor U12839 (N_12839,N_5036,N_8785);
nor U12840 (N_12840,N_7381,N_9642);
and U12841 (N_12841,N_9929,N_7204);
and U12842 (N_12842,N_5360,N_7740);
or U12843 (N_12843,N_8104,N_8262);
nand U12844 (N_12844,N_6868,N_6404);
or U12845 (N_12845,N_5276,N_5079);
nand U12846 (N_12846,N_6399,N_5917);
nor U12847 (N_12847,N_7208,N_8950);
and U12848 (N_12848,N_6616,N_8245);
nand U12849 (N_12849,N_8337,N_9827);
or U12850 (N_12850,N_8467,N_9194);
or U12851 (N_12851,N_9900,N_8865);
nand U12852 (N_12852,N_5656,N_8898);
nor U12853 (N_12853,N_8616,N_7524);
nand U12854 (N_12854,N_6247,N_5156);
and U12855 (N_12855,N_6957,N_8266);
nand U12856 (N_12856,N_9616,N_6251);
nand U12857 (N_12857,N_9481,N_5247);
and U12858 (N_12858,N_6880,N_5687);
nand U12859 (N_12859,N_9676,N_6560);
or U12860 (N_12860,N_6131,N_6717);
nand U12861 (N_12861,N_7950,N_6176);
nand U12862 (N_12862,N_7204,N_9707);
and U12863 (N_12863,N_5147,N_6781);
or U12864 (N_12864,N_6176,N_5008);
nand U12865 (N_12865,N_9323,N_8201);
and U12866 (N_12866,N_6858,N_6875);
or U12867 (N_12867,N_7474,N_5446);
nor U12868 (N_12868,N_6930,N_7505);
nor U12869 (N_12869,N_8631,N_7732);
and U12870 (N_12870,N_8335,N_8000);
nand U12871 (N_12871,N_5930,N_6401);
or U12872 (N_12872,N_6282,N_5572);
nand U12873 (N_12873,N_9139,N_6324);
or U12874 (N_12874,N_9497,N_9858);
xnor U12875 (N_12875,N_8406,N_5004);
or U12876 (N_12876,N_8747,N_8773);
or U12877 (N_12877,N_5510,N_8425);
nor U12878 (N_12878,N_8883,N_6352);
nand U12879 (N_12879,N_9612,N_5513);
or U12880 (N_12880,N_7121,N_7551);
and U12881 (N_12881,N_8461,N_9975);
or U12882 (N_12882,N_7517,N_8832);
and U12883 (N_12883,N_9217,N_8588);
nand U12884 (N_12884,N_9127,N_9371);
nand U12885 (N_12885,N_9931,N_6337);
nand U12886 (N_12886,N_8518,N_5759);
nand U12887 (N_12887,N_5604,N_7524);
nand U12888 (N_12888,N_7523,N_7012);
nand U12889 (N_12889,N_8710,N_5109);
nand U12890 (N_12890,N_9398,N_7895);
and U12891 (N_12891,N_5065,N_7548);
and U12892 (N_12892,N_7228,N_7734);
nor U12893 (N_12893,N_6145,N_6639);
nand U12894 (N_12894,N_5371,N_5153);
nor U12895 (N_12895,N_5355,N_6861);
and U12896 (N_12896,N_7497,N_7375);
and U12897 (N_12897,N_8833,N_7396);
and U12898 (N_12898,N_5552,N_7996);
nand U12899 (N_12899,N_6280,N_5053);
or U12900 (N_12900,N_6799,N_8697);
nor U12901 (N_12901,N_5537,N_9205);
or U12902 (N_12902,N_5069,N_8154);
nand U12903 (N_12903,N_6340,N_9636);
and U12904 (N_12904,N_9995,N_9244);
nor U12905 (N_12905,N_6520,N_5891);
or U12906 (N_12906,N_6144,N_5201);
and U12907 (N_12907,N_9212,N_8312);
or U12908 (N_12908,N_7520,N_9571);
and U12909 (N_12909,N_6848,N_9978);
or U12910 (N_12910,N_5469,N_5446);
nor U12911 (N_12911,N_5270,N_6025);
or U12912 (N_12912,N_9596,N_9729);
nand U12913 (N_12913,N_8599,N_6574);
and U12914 (N_12914,N_8253,N_8305);
or U12915 (N_12915,N_9226,N_6059);
nand U12916 (N_12916,N_8702,N_9697);
nand U12917 (N_12917,N_6245,N_6828);
nor U12918 (N_12918,N_9627,N_8457);
nor U12919 (N_12919,N_8383,N_9991);
nand U12920 (N_12920,N_8271,N_6195);
nor U12921 (N_12921,N_5859,N_5391);
and U12922 (N_12922,N_5664,N_6261);
nor U12923 (N_12923,N_6660,N_6934);
nor U12924 (N_12924,N_9211,N_5045);
nor U12925 (N_12925,N_5633,N_8256);
or U12926 (N_12926,N_7982,N_8196);
and U12927 (N_12927,N_8713,N_9716);
or U12928 (N_12928,N_5773,N_7435);
nand U12929 (N_12929,N_8235,N_8270);
or U12930 (N_12930,N_5483,N_7544);
nor U12931 (N_12931,N_5967,N_8983);
or U12932 (N_12932,N_5967,N_6274);
and U12933 (N_12933,N_7349,N_5715);
nand U12934 (N_12934,N_5179,N_5678);
nand U12935 (N_12935,N_5141,N_8915);
and U12936 (N_12936,N_6987,N_6381);
or U12937 (N_12937,N_5591,N_5566);
nor U12938 (N_12938,N_8987,N_6146);
or U12939 (N_12939,N_5346,N_8831);
and U12940 (N_12940,N_8011,N_6752);
nand U12941 (N_12941,N_8340,N_6191);
or U12942 (N_12942,N_6170,N_6272);
or U12943 (N_12943,N_9428,N_7461);
nor U12944 (N_12944,N_5396,N_5674);
nor U12945 (N_12945,N_5404,N_5381);
nand U12946 (N_12946,N_7535,N_7968);
nand U12947 (N_12947,N_8287,N_9903);
nand U12948 (N_12948,N_5082,N_5090);
nand U12949 (N_12949,N_7151,N_7331);
or U12950 (N_12950,N_5706,N_6713);
nand U12951 (N_12951,N_6619,N_7446);
and U12952 (N_12952,N_8435,N_5262);
nor U12953 (N_12953,N_9312,N_9803);
nand U12954 (N_12954,N_5009,N_7543);
nor U12955 (N_12955,N_9364,N_7890);
nor U12956 (N_12956,N_9479,N_9639);
and U12957 (N_12957,N_5706,N_9188);
or U12958 (N_12958,N_6416,N_9609);
and U12959 (N_12959,N_6117,N_9568);
nor U12960 (N_12960,N_5226,N_7204);
nor U12961 (N_12961,N_8526,N_7772);
and U12962 (N_12962,N_5456,N_9837);
and U12963 (N_12963,N_8110,N_7754);
or U12964 (N_12964,N_6336,N_6987);
and U12965 (N_12965,N_9129,N_5562);
and U12966 (N_12966,N_7902,N_9559);
nand U12967 (N_12967,N_6299,N_6665);
nor U12968 (N_12968,N_9383,N_6181);
or U12969 (N_12969,N_7835,N_5398);
nand U12970 (N_12970,N_9481,N_6126);
or U12971 (N_12971,N_7630,N_8681);
nor U12972 (N_12972,N_9901,N_7722);
nand U12973 (N_12973,N_5575,N_9090);
and U12974 (N_12974,N_5918,N_6292);
nor U12975 (N_12975,N_9105,N_7901);
and U12976 (N_12976,N_7672,N_8819);
and U12977 (N_12977,N_5952,N_6083);
and U12978 (N_12978,N_7351,N_7349);
nor U12979 (N_12979,N_6550,N_7542);
or U12980 (N_12980,N_9612,N_7302);
and U12981 (N_12981,N_8156,N_8674);
or U12982 (N_12982,N_8180,N_8362);
and U12983 (N_12983,N_7543,N_8910);
nand U12984 (N_12984,N_9156,N_7823);
nand U12985 (N_12985,N_8148,N_5147);
nand U12986 (N_12986,N_9372,N_7561);
and U12987 (N_12987,N_9146,N_8059);
nor U12988 (N_12988,N_6316,N_7695);
nand U12989 (N_12989,N_9308,N_8890);
nand U12990 (N_12990,N_9111,N_7413);
nor U12991 (N_12991,N_9518,N_6919);
nor U12992 (N_12992,N_9605,N_5561);
nor U12993 (N_12993,N_8984,N_7711);
nand U12994 (N_12994,N_5055,N_9346);
or U12995 (N_12995,N_9935,N_5266);
and U12996 (N_12996,N_5284,N_7409);
and U12997 (N_12997,N_8383,N_8175);
nor U12998 (N_12998,N_9700,N_9823);
nand U12999 (N_12999,N_6395,N_6388);
and U13000 (N_13000,N_6438,N_8592);
and U13001 (N_13001,N_7473,N_9571);
nand U13002 (N_13002,N_6017,N_9096);
nor U13003 (N_13003,N_6019,N_7845);
or U13004 (N_13004,N_9328,N_6957);
and U13005 (N_13005,N_7166,N_6892);
or U13006 (N_13006,N_8916,N_7908);
nor U13007 (N_13007,N_7770,N_8075);
or U13008 (N_13008,N_5347,N_7150);
nor U13009 (N_13009,N_6983,N_5306);
nor U13010 (N_13010,N_5147,N_6786);
nand U13011 (N_13011,N_6902,N_6904);
nor U13012 (N_13012,N_6620,N_9953);
nor U13013 (N_13013,N_5092,N_5619);
nand U13014 (N_13014,N_8054,N_5914);
nor U13015 (N_13015,N_9415,N_9906);
or U13016 (N_13016,N_5538,N_9119);
and U13017 (N_13017,N_7240,N_7878);
nand U13018 (N_13018,N_7246,N_8139);
and U13019 (N_13019,N_8098,N_8292);
and U13020 (N_13020,N_7747,N_5149);
nor U13021 (N_13021,N_7936,N_8115);
nor U13022 (N_13022,N_7466,N_5970);
xor U13023 (N_13023,N_8582,N_9993);
nor U13024 (N_13024,N_8695,N_6862);
or U13025 (N_13025,N_9645,N_8572);
nor U13026 (N_13026,N_5745,N_9924);
and U13027 (N_13027,N_7274,N_9787);
nand U13028 (N_13028,N_6667,N_7639);
nor U13029 (N_13029,N_8622,N_9135);
nor U13030 (N_13030,N_8449,N_7682);
and U13031 (N_13031,N_7313,N_9883);
or U13032 (N_13032,N_8018,N_9037);
nand U13033 (N_13033,N_7720,N_7183);
nor U13034 (N_13034,N_7575,N_7889);
and U13035 (N_13035,N_7865,N_7710);
or U13036 (N_13036,N_6998,N_7528);
or U13037 (N_13037,N_8137,N_8256);
nor U13038 (N_13038,N_8275,N_9900);
nor U13039 (N_13039,N_8282,N_6191);
nand U13040 (N_13040,N_6343,N_6244);
nand U13041 (N_13041,N_5435,N_8916);
nor U13042 (N_13042,N_7231,N_9270);
nand U13043 (N_13043,N_9849,N_5841);
nor U13044 (N_13044,N_8396,N_8896);
and U13045 (N_13045,N_6611,N_6839);
nand U13046 (N_13046,N_9344,N_7965);
and U13047 (N_13047,N_8853,N_9744);
nor U13048 (N_13048,N_8105,N_9261);
or U13049 (N_13049,N_5863,N_8164);
nand U13050 (N_13050,N_8914,N_8757);
nand U13051 (N_13051,N_8184,N_8609);
nor U13052 (N_13052,N_8268,N_8337);
and U13053 (N_13053,N_7872,N_6160);
nor U13054 (N_13054,N_5956,N_8005);
or U13055 (N_13055,N_5776,N_7075);
and U13056 (N_13056,N_5414,N_8639);
or U13057 (N_13057,N_6524,N_8511);
nand U13058 (N_13058,N_7921,N_8581);
nand U13059 (N_13059,N_8590,N_5056);
nor U13060 (N_13060,N_9963,N_6980);
or U13061 (N_13061,N_9887,N_6809);
or U13062 (N_13062,N_6317,N_7078);
or U13063 (N_13063,N_5649,N_5152);
nor U13064 (N_13064,N_8383,N_6811);
and U13065 (N_13065,N_8582,N_8765);
nor U13066 (N_13066,N_8099,N_5503);
nand U13067 (N_13067,N_7406,N_6918);
and U13068 (N_13068,N_9859,N_9494);
or U13069 (N_13069,N_9904,N_8433);
nor U13070 (N_13070,N_6174,N_6556);
nand U13071 (N_13071,N_8925,N_8450);
nor U13072 (N_13072,N_8125,N_6898);
or U13073 (N_13073,N_8599,N_7660);
nand U13074 (N_13074,N_5476,N_6142);
and U13075 (N_13075,N_6044,N_7682);
nor U13076 (N_13076,N_5341,N_8119);
nand U13077 (N_13077,N_9865,N_6810);
nand U13078 (N_13078,N_9379,N_7186);
nor U13079 (N_13079,N_5332,N_7452);
or U13080 (N_13080,N_7902,N_5794);
and U13081 (N_13081,N_7403,N_7174);
nor U13082 (N_13082,N_9324,N_9128);
and U13083 (N_13083,N_9816,N_8367);
or U13084 (N_13084,N_7473,N_5150);
nor U13085 (N_13085,N_8069,N_6269);
nand U13086 (N_13086,N_8338,N_5464);
nand U13087 (N_13087,N_9847,N_9652);
nor U13088 (N_13088,N_8475,N_5268);
or U13089 (N_13089,N_7395,N_9711);
nand U13090 (N_13090,N_8880,N_5846);
and U13091 (N_13091,N_7975,N_5937);
nor U13092 (N_13092,N_8640,N_9907);
and U13093 (N_13093,N_9068,N_7323);
or U13094 (N_13094,N_8314,N_9725);
or U13095 (N_13095,N_9724,N_6482);
and U13096 (N_13096,N_8154,N_8894);
and U13097 (N_13097,N_6398,N_6835);
nand U13098 (N_13098,N_7443,N_6689);
nor U13099 (N_13099,N_5663,N_9936);
xor U13100 (N_13100,N_5090,N_7651);
and U13101 (N_13101,N_5212,N_5374);
nor U13102 (N_13102,N_5449,N_5697);
nand U13103 (N_13103,N_7986,N_8799);
nor U13104 (N_13104,N_9603,N_6558);
or U13105 (N_13105,N_5561,N_6566);
nor U13106 (N_13106,N_5292,N_8281);
and U13107 (N_13107,N_8191,N_7822);
or U13108 (N_13108,N_7799,N_7752);
and U13109 (N_13109,N_7762,N_5382);
and U13110 (N_13110,N_5174,N_5721);
or U13111 (N_13111,N_8618,N_7994);
nand U13112 (N_13112,N_5105,N_6797);
nor U13113 (N_13113,N_7758,N_5056);
nand U13114 (N_13114,N_7406,N_6696);
or U13115 (N_13115,N_7132,N_8545);
nand U13116 (N_13116,N_7046,N_5167);
nand U13117 (N_13117,N_5673,N_7296);
nor U13118 (N_13118,N_6515,N_6245);
or U13119 (N_13119,N_8851,N_5981);
nand U13120 (N_13120,N_6807,N_9960);
nand U13121 (N_13121,N_5275,N_7893);
nand U13122 (N_13122,N_7408,N_8645);
and U13123 (N_13123,N_8341,N_6458);
or U13124 (N_13124,N_9160,N_5841);
or U13125 (N_13125,N_5008,N_5568);
and U13126 (N_13126,N_6232,N_6449);
nand U13127 (N_13127,N_5030,N_7264);
or U13128 (N_13128,N_6057,N_9512);
nand U13129 (N_13129,N_9285,N_5387);
nor U13130 (N_13130,N_7775,N_8796);
nand U13131 (N_13131,N_8911,N_7422);
and U13132 (N_13132,N_5756,N_8415);
or U13133 (N_13133,N_6016,N_6539);
or U13134 (N_13134,N_8234,N_9821);
and U13135 (N_13135,N_8418,N_9414);
xor U13136 (N_13136,N_6585,N_7282);
and U13137 (N_13137,N_5883,N_8058);
or U13138 (N_13138,N_8853,N_7883);
xnor U13139 (N_13139,N_6862,N_5655);
and U13140 (N_13140,N_5929,N_8979);
nand U13141 (N_13141,N_6471,N_8914);
and U13142 (N_13142,N_9011,N_7630);
or U13143 (N_13143,N_5523,N_8065);
or U13144 (N_13144,N_7329,N_6579);
or U13145 (N_13145,N_6565,N_6012);
nor U13146 (N_13146,N_5046,N_7368);
nor U13147 (N_13147,N_8275,N_5488);
nor U13148 (N_13148,N_9088,N_5779);
nor U13149 (N_13149,N_9149,N_5402);
nor U13150 (N_13150,N_8248,N_9121);
nor U13151 (N_13151,N_9528,N_9724);
nor U13152 (N_13152,N_5738,N_6096);
nor U13153 (N_13153,N_7726,N_9746);
nand U13154 (N_13154,N_8600,N_7520);
nor U13155 (N_13155,N_9136,N_7663);
nor U13156 (N_13156,N_9983,N_8109);
and U13157 (N_13157,N_8873,N_7604);
nand U13158 (N_13158,N_9203,N_7904);
nand U13159 (N_13159,N_5055,N_9180);
or U13160 (N_13160,N_8416,N_6908);
nor U13161 (N_13161,N_6514,N_7278);
nand U13162 (N_13162,N_6673,N_6078);
or U13163 (N_13163,N_7057,N_6012);
nand U13164 (N_13164,N_6175,N_8515);
or U13165 (N_13165,N_5294,N_6272);
or U13166 (N_13166,N_9988,N_5315);
and U13167 (N_13167,N_8811,N_8385);
or U13168 (N_13168,N_5411,N_8979);
xor U13169 (N_13169,N_8866,N_5548);
nor U13170 (N_13170,N_5968,N_7121);
or U13171 (N_13171,N_5304,N_7520);
or U13172 (N_13172,N_7969,N_7624);
nand U13173 (N_13173,N_5778,N_7642);
nand U13174 (N_13174,N_9597,N_5261);
nor U13175 (N_13175,N_6740,N_7514);
and U13176 (N_13176,N_7085,N_6801);
xnor U13177 (N_13177,N_7603,N_7037);
and U13178 (N_13178,N_8620,N_7590);
and U13179 (N_13179,N_6539,N_6923);
or U13180 (N_13180,N_9154,N_7514);
and U13181 (N_13181,N_7425,N_8235);
xnor U13182 (N_13182,N_6600,N_5676);
nor U13183 (N_13183,N_8514,N_5377);
or U13184 (N_13184,N_8564,N_7483);
nor U13185 (N_13185,N_8130,N_9975);
nand U13186 (N_13186,N_7625,N_5585);
or U13187 (N_13187,N_5572,N_5025);
and U13188 (N_13188,N_9035,N_5277);
nand U13189 (N_13189,N_9122,N_6915);
nor U13190 (N_13190,N_9059,N_9490);
and U13191 (N_13191,N_5691,N_8946);
nor U13192 (N_13192,N_6289,N_8480);
nand U13193 (N_13193,N_6062,N_7825);
or U13194 (N_13194,N_9879,N_7541);
and U13195 (N_13195,N_9465,N_9861);
or U13196 (N_13196,N_5328,N_7308);
and U13197 (N_13197,N_9127,N_6847);
and U13198 (N_13198,N_9383,N_8549);
and U13199 (N_13199,N_8990,N_9563);
and U13200 (N_13200,N_8149,N_5469);
nand U13201 (N_13201,N_6336,N_7889);
or U13202 (N_13202,N_9243,N_8372);
nand U13203 (N_13203,N_9050,N_5296);
or U13204 (N_13204,N_6382,N_5678);
nor U13205 (N_13205,N_6849,N_8088);
nand U13206 (N_13206,N_7264,N_5115);
and U13207 (N_13207,N_9285,N_5286);
and U13208 (N_13208,N_5854,N_5965);
nand U13209 (N_13209,N_6351,N_8533);
and U13210 (N_13210,N_7029,N_7044);
or U13211 (N_13211,N_8397,N_8907);
and U13212 (N_13212,N_9448,N_6327);
nand U13213 (N_13213,N_7115,N_9540);
or U13214 (N_13214,N_8925,N_7720);
nand U13215 (N_13215,N_6425,N_6323);
and U13216 (N_13216,N_8212,N_5014);
nand U13217 (N_13217,N_9488,N_7139);
or U13218 (N_13218,N_6013,N_6607);
or U13219 (N_13219,N_7130,N_7464);
nor U13220 (N_13220,N_5144,N_7549);
and U13221 (N_13221,N_8831,N_7900);
nor U13222 (N_13222,N_8386,N_5460);
or U13223 (N_13223,N_9923,N_5538);
or U13224 (N_13224,N_8660,N_7597);
nor U13225 (N_13225,N_9813,N_7894);
and U13226 (N_13226,N_6318,N_5281);
nor U13227 (N_13227,N_8713,N_6266);
nor U13228 (N_13228,N_6456,N_9595);
nor U13229 (N_13229,N_9190,N_7534);
nand U13230 (N_13230,N_5482,N_8907);
and U13231 (N_13231,N_6595,N_9173);
and U13232 (N_13232,N_6169,N_7973);
nand U13233 (N_13233,N_5722,N_7837);
nor U13234 (N_13234,N_9780,N_9402);
nor U13235 (N_13235,N_7558,N_7098);
or U13236 (N_13236,N_9366,N_6905);
nor U13237 (N_13237,N_9084,N_7477);
nand U13238 (N_13238,N_5273,N_8893);
or U13239 (N_13239,N_7218,N_6046);
nor U13240 (N_13240,N_6843,N_9137);
or U13241 (N_13241,N_7662,N_6849);
and U13242 (N_13242,N_7086,N_6605);
nand U13243 (N_13243,N_6199,N_8266);
and U13244 (N_13244,N_8964,N_5916);
or U13245 (N_13245,N_8299,N_9944);
nor U13246 (N_13246,N_5673,N_9589);
nor U13247 (N_13247,N_8369,N_5920);
xor U13248 (N_13248,N_8903,N_5126);
nand U13249 (N_13249,N_6196,N_6255);
nor U13250 (N_13250,N_7311,N_8511);
nor U13251 (N_13251,N_8980,N_9599);
or U13252 (N_13252,N_8482,N_6078);
or U13253 (N_13253,N_7181,N_8168);
nor U13254 (N_13254,N_7888,N_6300);
or U13255 (N_13255,N_5740,N_8874);
and U13256 (N_13256,N_5254,N_7026);
xor U13257 (N_13257,N_5705,N_5462);
or U13258 (N_13258,N_5407,N_9028);
nor U13259 (N_13259,N_9274,N_8948);
and U13260 (N_13260,N_9501,N_5136);
nand U13261 (N_13261,N_5322,N_8181);
or U13262 (N_13262,N_8612,N_9107);
nand U13263 (N_13263,N_8189,N_8245);
or U13264 (N_13264,N_7182,N_7882);
and U13265 (N_13265,N_7284,N_6888);
nand U13266 (N_13266,N_8697,N_6466);
or U13267 (N_13267,N_9014,N_8148);
nand U13268 (N_13268,N_9472,N_5576);
or U13269 (N_13269,N_5315,N_5310);
nand U13270 (N_13270,N_6861,N_5225);
or U13271 (N_13271,N_6062,N_7629);
nor U13272 (N_13272,N_5194,N_8717);
or U13273 (N_13273,N_9620,N_8184);
and U13274 (N_13274,N_7404,N_6810);
and U13275 (N_13275,N_5292,N_7274);
nor U13276 (N_13276,N_6452,N_8480);
nand U13277 (N_13277,N_9219,N_5014);
nand U13278 (N_13278,N_9299,N_7497);
nor U13279 (N_13279,N_8779,N_7891);
and U13280 (N_13280,N_9752,N_8317);
nor U13281 (N_13281,N_6313,N_6718);
nor U13282 (N_13282,N_6250,N_8091);
nor U13283 (N_13283,N_6681,N_6921);
nor U13284 (N_13284,N_6728,N_8283);
or U13285 (N_13285,N_5800,N_5962);
and U13286 (N_13286,N_9923,N_8436);
and U13287 (N_13287,N_5893,N_7405);
and U13288 (N_13288,N_5885,N_5663);
or U13289 (N_13289,N_9743,N_5395);
nor U13290 (N_13290,N_5383,N_5493);
and U13291 (N_13291,N_6299,N_6309);
nor U13292 (N_13292,N_5875,N_9969);
or U13293 (N_13293,N_7502,N_6454);
and U13294 (N_13294,N_9532,N_5310);
nand U13295 (N_13295,N_6092,N_8135);
nor U13296 (N_13296,N_7992,N_9458);
and U13297 (N_13297,N_9173,N_8929);
and U13298 (N_13298,N_9174,N_6387);
nand U13299 (N_13299,N_5805,N_7502);
nor U13300 (N_13300,N_7017,N_8925);
nand U13301 (N_13301,N_5146,N_5194);
and U13302 (N_13302,N_7879,N_7012);
or U13303 (N_13303,N_7083,N_6666);
nor U13304 (N_13304,N_6173,N_8024);
nor U13305 (N_13305,N_7879,N_7692);
nand U13306 (N_13306,N_6541,N_6955);
nor U13307 (N_13307,N_5665,N_8532);
nor U13308 (N_13308,N_7816,N_9171);
nand U13309 (N_13309,N_8769,N_6631);
nand U13310 (N_13310,N_7640,N_6479);
nand U13311 (N_13311,N_6700,N_5309);
or U13312 (N_13312,N_7371,N_6718);
or U13313 (N_13313,N_7074,N_9734);
or U13314 (N_13314,N_6967,N_9743);
nand U13315 (N_13315,N_8676,N_7410);
nor U13316 (N_13316,N_9889,N_9550);
and U13317 (N_13317,N_5081,N_5008);
or U13318 (N_13318,N_5680,N_8095);
and U13319 (N_13319,N_7695,N_7839);
nor U13320 (N_13320,N_7745,N_6774);
or U13321 (N_13321,N_9191,N_7921);
nor U13322 (N_13322,N_9889,N_7410);
or U13323 (N_13323,N_8893,N_6040);
nor U13324 (N_13324,N_7334,N_5531);
and U13325 (N_13325,N_8997,N_8271);
and U13326 (N_13326,N_6867,N_6106);
or U13327 (N_13327,N_7601,N_9469);
or U13328 (N_13328,N_7173,N_6476);
or U13329 (N_13329,N_7038,N_9732);
and U13330 (N_13330,N_5007,N_8832);
or U13331 (N_13331,N_9719,N_7305);
nor U13332 (N_13332,N_9022,N_8164);
and U13333 (N_13333,N_7522,N_5426);
nand U13334 (N_13334,N_9948,N_8747);
nand U13335 (N_13335,N_8728,N_9995);
nand U13336 (N_13336,N_6252,N_6662);
or U13337 (N_13337,N_9636,N_6270);
and U13338 (N_13338,N_5961,N_7104);
nor U13339 (N_13339,N_5031,N_7856);
nor U13340 (N_13340,N_5692,N_9257);
nand U13341 (N_13341,N_9115,N_8935);
nor U13342 (N_13342,N_6913,N_5428);
or U13343 (N_13343,N_8576,N_9715);
or U13344 (N_13344,N_9798,N_5046);
nand U13345 (N_13345,N_8257,N_9998);
and U13346 (N_13346,N_6326,N_7398);
and U13347 (N_13347,N_7632,N_5724);
and U13348 (N_13348,N_8741,N_8858);
or U13349 (N_13349,N_9917,N_9107);
and U13350 (N_13350,N_5974,N_7625);
nor U13351 (N_13351,N_8522,N_5068);
xor U13352 (N_13352,N_7446,N_6993);
nand U13353 (N_13353,N_6081,N_6188);
nand U13354 (N_13354,N_9991,N_5517);
nand U13355 (N_13355,N_9983,N_8025);
and U13356 (N_13356,N_8754,N_7170);
and U13357 (N_13357,N_8982,N_6609);
and U13358 (N_13358,N_9974,N_9903);
or U13359 (N_13359,N_7450,N_8926);
and U13360 (N_13360,N_9308,N_5493);
nand U13361 (N_13361,N_9404,N_6834);
and U13362 (N_13362,N_9009,N_9174);
and U13363 (N_13363,N_6920,N_6437);
or U13364 (N_13364,N_8261,N_8629);
nor U13365 (N_13365,N_7543,N_7488);
nor U13366 (N_13366,N_6228,N_5729);
and U13367 (N_13367,N_9138,N_9307);
and U13368 (N_13368,N_7131,N_7649);
nor U13369 (N_13369,N_6207,N_8961);
nor U13370 (N_13370,N_5713,N_5702);
nor U13371 (N_13371,N_6368,N_8801);
and U13372 (N_13372,N_7994,N_5346);
and U13373 (N_13373,N_5743,N_6608);
xnor U13374 (N_13374,N_8323,N_9720);
nor U13375 (N_13375,N_8880,N_7386);
or U13376 (N_13376,N_5779,N_7978);
nor U13377 (N_13377,N_7440,N_8727);
and U13378 (N_13378,N_5424,N_9679);
or U13379 (N_13379,N_8953,N_9568);
or U13380 (N_13380,N_7822,N_7380);
or U13381 (N_13381,N_7697,N_8602);
and U13382 (N_13382,N_9292,N_5870);
and U13383 (N_13383,N_5632,N_7276);
nand U13384 (N_13384,N_6810,N_7701);
nor U13385 (N_13385,N_8459,N_6976);
or U13386 (N_13386,N_9014,N_9699);
and U13387 (N_13387,N_7179,N_8135);
or U13388 (N_13388,N_9064,N_9634);
nand U13389 (N_13389,N_6069,N_9363);
and U13390 (N_13390,N_6426,N_6247);
nor U13391 (N_13391,N_5390,N_7399);
and U13392 (N_13392,N_8197,N_5884);
and U13393 (N_13393,N_7577,N_6482);
nand U13394 (N_13394,N_7186,N_5549);
nor U13395 (N_13395,N_8322,N_5288);
or U13396 (N_13396,N_5116,N_9866);
nand U13397 (N_13397,N_8144,N_8606);
and U13398 (N_13398,N_6992,N_9184);
nand U13399 (N_13399,N_6999,N_5841);
or U13400 (N_13400,N_7565,N_9224);
nor U13401 (N_13401,N_6609,N_8097);
or U13402 (N_13402,N_9307,N_5356);
nand U13403 (N_13403,N_7427,N_9528);
nor U13404 (N_13404,N_5294,N_8690);
or U13405 (N_13405,N_8755,N_6263);
and U13406 (N_13406,N_9067,N_6063);
nand U13407 (N_13407,N_7188,N_9341);
and U13408 (N_13408,N_7609,N_5509);
xor U13409 (N_13409,N_9212,N_9208);
nand U13410 (N_13410,N_6961,N_7743);
and U13411 (N_13411,N_8428,N_8992);
nand U13412 (N_13412,N_7823,N_5930);
nor U13413 (N_13413,N_7474,N_5885);
nand U13414 (N_13414,N_5985,N_6014);
nor U13415 (N_13415,N_9138,N_7313);
or U13416 (N_13416,N_7130,N_7237);
nor U13417 (N_13417,N_6259,N_5761);
or U13418 (N_13418,N_8449,N_5571);
and U13419 (N_13419,N_9289,N_5629);
and U13420 (N_13420,N_9255,N_5751);
or U13421 (N_13421,N_8159,N_5574);
and U13422 (N_13422,N_7014,N_6744);
nand U13423 (N_13423,N_8748,N_7129);
or U13424 (N_13424,N_9036,N_9622);
and U13425 (N_13425,N_8875,N_6841);
or U13426 (N_13426,N_9804,N_6324);
or U13427 (N_13427,N_5866,N_8474);
or U13428 (N_13428,N_5136,N_8242);
and U13429 (N_13429,N_9665,N_7165);
and U13430 (N_13430,N_7298,N_5677);
or U13431 (N_13431,N_5227,N_5099);
and U13432 (N_13432,N_5460,N_9510);
nand U13433 (N_13433,N_5062,N_5403);
nand U13434 (N_13434,N_5518,N_6512);
nor U13435 (N_13435,N_7444,N_8149);
nand U13436 (N_13436,N_5504,N_8898);
or U13437 (N_13437,N_6559,N_5081);
nand U13438 (N_13438,N_8543,N_9557);
nor U13439 (N_13439,N_9154,N_9612);
or U13440 (N_13440,N_6981,N_7695);
or U13441 (N_13441,N_9205,N_6497);
and U13442 (N_13442,N_6803,N_5425);
and U13443 (N_13443,N_9930,N_6546);
nor U13444 (N_13444,N_8742,N_9678);
and U13445 (N_13445,N_6213,N_7816);
and U13446 (N_13446,N_7662,N_7742);
or U13447 (N_13447,N_8356,N_6721);
nor U13448 (N_13448,N_9841,N_9869);
or U13449 (N_13449,N_6189,N_7723);
or U13450 (N_13450,N_5706,N_8033);
nor U13451 (N_13451,N_6201,N_9970);
and U13452 (N_13452,N_6653,N_5585);
or U13453 (N_13453,N_7617,N_9508);
nand U13454 (N_13454,N_7902,N_9472);
nor U13455 (N_13455,N_6266,N_9326);
and U13456 (N_13456,N_7996,N_6758);
and U13457 (N_13457,N_9050,N_5894);
nor U13458 (N_13458,N_5178,N_5286);
nor U13459 (N_13459,N_7214,N_6569);
nand U13460 (N_13460,N_5405,N_8731);
nand U13461 (N_13461,N_6851,N_5610);
or U13462 (N_13462,N_8542,N_7649);
nor U13463 (N_13463,N_5651,N_6819);
and U13464 (N_13464,N_9316,N_8544);
or U13465 (N_13465,N_6217,N_8571);
or U13466 (N_13466,N_8003,N_5234);
or U13467 (N_13467,N_5667,N_8780);
nand U13468 (N_13468,N_7386,N_9047);
and U13469 (N_13469,N_8859,N_9044);
nand U13470 (N_13470,N_7882,N_8079);
and U13471 (N_13471,N_7413,N_8553);
nand U13472 (N_13472,N_6976,N_7627);
or U13473 (N_13473,N_8664,N_6042);
nand U13474 (N_13474,N_6602,N_8861);
and U13475 (N_13475,N_7629,N_9974);
nor U13476 (N_13476,N_7404,N_6228);
and U13477 (N_13477,N_9338,N_6097);
nor U13478 (N_13478,N_7618,N_7049);
or U13479 (N_13479,N_6614,N_8352);
and U13480 (N_13480,N_8313,N_8152);
nand U13481 (N_13481,N_8464,N_7543);
or U13482 (N_13482,N_5247,N_7186);
nand U13483 (N_13483,N_7586,N_5580);
or U13484 (N_13484,N_5089,N_7230);
nand U13485 (N_13485,N_8623,N_7944);
and U13486 (N_13486,N_8730,N_7885);
or U13487 (N_13487,N_9711,N_7937);
or U13488 (N_13488,N_5411,N_5240);
nor U13489 (N_13489,N_6582,N_7771);
nand U13490 (N_13490,N_7998,N_7426);
and U13491 (N_13491,N_8774,N_5193);
nand U13492 (N_13492,N_5110,N_9724);
nor U13493 (N_13493,N_5993,N_7708);
or U13494 (N_13494,N_6928,N_6208);
nor U13495 (N_13495,N_5437,N_6951);
and U13496 (N_13496,N_5190,N_8692);
nor U13497 (N_13497,N_8833,N_5223);
nor U13498 (N_13498,N_7824,N_9996);
or U13499 (N_13499,N_7268,N_6180);
and U13500 (N_13500,N_5695,N_7800);
and U13501 (N_13501,N_5537,N_6238);
nand U13502 (N_13502,N_5181,N_6811);
nor U13503 (N_13503,N_6683,N_6224);
or U13504 (N_13504,N_6832,N_8550);
and U13505 (N_13505,N_7780,N_8875);
nor U13506 (N_13506,N_6950,N_9327);
or U13507 (N_13507,N_9729,N_5347);
and U13508 (N_13508,N_8540,N_7197);
and U13509 (N_13509,N_7021,N_7212);
nand U13510 (N_13510,N_8148,N_9953);
and U13511 (N_13511,N_5359,N_5554);
and U13512 (N_13512,N_7836,N_8251);
and U13513 (N_13513,N_8371,N_7761);
and U13514 (N_13514,N_5442,N_9642);
nor U13515 (N_13515,N_7730,N_9017);
and U13516 (N_13516,N_8348,N_7032);
nand U13517 (N_13517,N_6096,N_7020);
nor U13518 (N_13518,N_6260,N_8444);
or U13519 (N_13519,N_8249,N_5670);
or U13520 (N_13520,N_8250,N_8727);
and U13521 (N_13521,N_9367,N_7305);
nand U13522 (N_13522,N_5574,N_9285);
nor U13523 (N_13523,N_8507,N_8367);
and U13524 (N_13524,N_6105,N_8030);
and U13525 (N_13525,N_6020,N_6599);
and U13526 (N_13526,N_8275,N_5996);
and U13527 (N_13527,N_5184,N_6326);
and U13528 (N_13528,N_6014,N_9454);
or U13529 (N_13529,N_6638,N_9844);
nor U13530 (N_13530,N_8181,N_7571);
or U13531 (N_13531,N_8525,N_5724);
nand U13532 (N_13532,N_7386,N_9972);
or U13533 (N_13533,N_7238,N_7837);
xnor U13534 (N_13534,N_8931,N_5604);
or U13535 (N_13535,N_9145,N_5200);
or U13536 (N_13536,N_5191,N_6485);
nand U13537 (N_13537,N_9607,N_6101);
and U13538 (N_13538,N_5754,N_6630);
and U13539 (N_13539,N_5765,N_8469);
and U13540 (N_13540,N_7696,N_9941);
nor U13541 (N_13541,N_6127,N_6290);
nor U13542 (N_13542,N_9156,N_5355);
nand U13543 (N_13543,N_9834,N_9557);
or U13544 (N_13544,N_5310,N_5644);
and U13545 (N_13545,N_6715,N_6451);
nor U13546 (N_13546,N_7982,N_6750);
nor U13547 (N_13547,N_5616,N_9952);
xnor U13548 (N_13548,N_9430,N_7434);
nor U13549 (N_13549,N_6804,N_9052);
nand U13550 (N_13550,N_7013,N_5671);
or U13551 (N_13551,N_6225,N_7008);
nand U13552 (N_13552,N_6747,N_9051);
nor U13553 (N_13553,N_5440,N_8873);
and U13554 (N_13554,N_8623,N_9262);
nand U13555 (N_13555,N_5599,N_5737);
nor U13556 (N_13556,N_7189,N_7818);
nor U13557 (N_13557,N_7741,N_8362);
and U13558 (N_13558,N_7755,N_6691);
nand U13559 (N_13559,N_5881,N_5549);
and U13560 (N_13560,N_6955,N_6886);
and U13561 (N_13561,N_6057,N_9469);
or U13562 (N_13562,N_8473,N_6388);
nor U13563 (N_13563,N_8693,N_9773);
or U13564 (N_13564,N_6468,N_6619);
and U13565 (N_13565,N_6251,N_9135);
nor U13566 (N_13566,N_8698,N_8207);
or U13567 (N_13567,N_7298,N_9625);
or U13568 (N_13568,N_6175,N_7714);
or U13569 (N_13569,N_8602,N_6746);
nand U13570 (N_13570,N_7490,N_8313);
nor U13571 (N_13571,N_7684,N_6595);
or U13572 (N_13572,N_6162,N_7401);
and U13573 (N_13573,N_6083,N_6548);
or U13574 (N_13574,N_9831,N_8065);
and U13575 (N_13575,N_9594,N_8010);
nor U13576 (N_13576,N_8383,N_6270);
nor U13577 (N_13577,N_8615,N_6496);
or U13578 (N_13578,N_9026,N_6401);
nor U13579 (N_13579,N_7923,N_6619);
and U13580 (N_13580,N_5055,N_9193);
or U13581 (N_13581,N_9008,N_5170);
nor U13582 (N_13582,N_9968,N_7038);
nand U13583 (N_13583,N_7350,N_6568);
and U13584 (N_13584,N_5875,N_5968);
nor U13585 (N_13585,N_5838,N_8083);
or U13586 (N_13586,N_6289,N_7568);
and U13587 (N_13587,N_6593,N_5201);
nor U13588 (N_13588,N_5647,N_8426);
nor U13589 (N_13589,N_7610,N_5915);
nor U13590 (N_13590,N_8255,N_6468);
or U13591 (N_13591,N_9207,N_9774);
or U13592 (N_13592,N_8860,N_8250);
and U13593 (N_13593,N_7789,N_7612);
or U13594 (N_13594,N_9544,N_6984);
and U13595 (N_13595,N_9676,N_8856);
nor U13596 (N_13596,N_9245,N_8041);
nor U13597 (N_13597,N_8611,N_9903);
or U13598 (N_13598,N_9407,N_8023);
and U13599 (N_13599,N_6988,N_9684);
and U13600 (N_13600,N_5030,N_5979);
nand U13601 (N_13601,N_7188,N_5193);
nand U13602 (N_13602,N_6173,N_8574);
and U13603 (N_13603,N_7228,N_8653);
nand U13604 (N_13604,N_9094,N_6405);
nor U13605 (N_13605,N_8353,N_8481);
or U13606 (N_13606,N_9424,N_6214);
and U13607 (N_13607,N_6607,N_8715);
and U13608 (N_13608,N_8122,N_9881);
and U13609 (N_13609,N_8924,N_8907);
and U13610 (N_13610,N_7018,N_6917);
nand U13611 (N_13611,N_6442,N_7188);
or U13612 (N_13612,N_5205,N_9919);
nor U13613 (N_13613,N_9321,N_8582);
nor U13614 (N_13614,N_5465,N_6714);
or U13615 (N_13615,N_8704,N_8982);
or U13616 (N_13616,N_8675,N_6834);
or U13617 (N_13617,N_5629,N_5657);
nand U13618 (N_13618,N_8442,N_5471);
and U13619 (N_13619,N_5305,N_9292);
nand U13620 (N_13620,N_7082,N_6796);
or U13621 (N_13621,N_8099,N_8496);
or U13622 (N_13622,N_8518,N_9386);
or U13623 (N_13623,N_6301,N_9368);
nor U13624 (N_13624,N_9051,N_6314);
nor U13625 (N_13625,N_6476,N_5040);
or U13626 (N_13626,N_5957,N_7941);
nand U13627 (N_13627,N_7440,N_6323);
or U13628 (N_13628,N_6106,N_6095);
or U13629 (N_13629,N_7421,N_6836);
nor U13630 (N_13630,N_6479,N_5678);
and U13631 (N_13631,N_6037,N_8070);
and U13632 (N_13632,N_9283,N_9837);
or U13633 (N_13633,N_8825,N_7201);
nor U13634 (N_13634,N_6617,N_8351);
nor U13635 (N_13635,N_7855,N_5585);
nand U13636 (N_13636,N_5424,N_6664);
nor U13637 (N_13637,N_8484,N_5195);
or U13638 (N_13638,N_6439,N_6911);
nand U13639 (N_13639,N_7666,N_9672);
or U13640 (N_13640,N_6334,N_8640);
and U13641 (N_13641,N_7921,N_9429);
nor U13642 (N_13642,N_7744,N_5311);
nand U13643 (N_13643,N_8160,N_8174);
nor U13644 (N_13644,N_8032,N_6204);
or U13645 (N_13645,N_6979,N_5073);
and U13646 (N_13646,N_5755,N_9459);
or U13647 (N_13647,N_8613,N_8292);
nor U13648 (N_13648,N_6033,N_5956);
nand U13649 (N_13649,N_9035,N_9613);
nor U13650 (N_13650,N_8191,N_8146);
nor U13651 (N_13651,N_5468,N_8837);
and U13652 (N_13652,N_7653,N_6543);
nand U13653 (N_13653,N_9915,N_5432);
nor U13654 (N_13654,N_8756,N_5641);
nor U13655 (N_13655,N_8225,N_6294);
nand U13656 (N_13656,N_5393,N_9203);
or U13657 (N_13657,N_8640,N_9986);
nand U13658 (N_13658,N_8010,N_8141);
or U13659 (N_13659,N_9047,N_9546);
and U13660 (N_13660,N_5947,N_8437);
or U13661 (N_13661,N_6950,N_6408);
or U13662 (N_13662,N_6727,N_7000);
or U13663 (N_13663,N_9775,N_9749);
nand U13664 (N_13664,N_9434,N_5145);
nor U13665 (N_13665,N_6578,N_6780);
and U13666 (N_13666,N_6913,N_7307);
nor U13667 (N_13667,N_6940,N_9118);
and U13668 (N_13668,N_8621,N_7719);
and U13669 (N_13669,N_9700,N_8067);
nand U13670 (N_13670,N_6221,N_5631);
or U13671 (N_13671,N_9499,N_8681);
and U13672 (N_13672,N_5603,N_5027);
and U13673 (N_13673,N_6452,N_9824);
or U13674 (N_13674,N_7161,N_8855);
nor U13675 (N_13675,N_6494,N_6148);
or U13676 (N_13676,N_8872,N_6602);
or U13677 (N_13677,N_8386,N_9208);
and U13678 (N_13678,N_9048,N_8061);
and U13679 (N_13679,N_8559,N_9698);
nor U13680 (N_13680,N_8916,N_7317);
nor U13681 (N_13681,N_7760,N_8421);
nand U13682 (N_13682,N_8448,N_6857);
or U13683 (N_13683,N_9391,N_6695);
and U13684 (N_13684,N_5887,N_9423);
nand U13685 (N_13685,N_5711,N_9676);
and U13686 (N_13686,N_7531,N_6436);
or U13687 (N_13687,N_5174,N_8272);
nand U13688 (N_13688,N_9249,N_9818);
nand U13689 (N_13689,N_5194,N_6229);
or U13690 (N_13690,N_6223,N_7605);
or U13691 (N_13691,N_5186,N_9033);
and U13692 (N_13692,N_9310,N_7120);
nand U13693 (N_13693,N_5004,N_8158);
or U13694 (N_13694,N_5759,N_7866);
and U13695 (N_13695,N_9307,N_9501);
nand U13696 (N_13696,N_5627,N_5094);
nor U13697 (N_13697,N_7093,N_7408);
or U13698 (N_13698,N_5762,N_9769);
or U13699 (N_13699,N_8648,N_8741);
nor U13700 (N_13700,N_5788,N_5457);
nand U13701 (N_13701,N_5833,N_9338);
or U13702 (N_13702,N_7375,N_5212);
and U13703 (N_13703,N_7906,N_6492);
nor U13704 (N_13704,N_5326,N_5580);
nor U13705 (N_13705,N_9617,N_9945);
nand U13706 (N_13706,N_6348,N_8452);
or U13707 (N_13707,N_8945,N_6818);
and U13708 (N_13708,N_5378,N_7132);
nand U13709 (N_13709,N_7966,N_5678);
nor U13710 (N_13710,N_9788,N_6542);
or U13711 (N_13711,N_9875,N_8875);
nor U13712 (N_13712,N_9090,N_6461);
or U13713 (N_13713,N_8363,N_5771);
and U13714 (N_13714,N_9663,N_9445);
nand U13715 (N_13715,N_9110,N_8463);
or U13716 (N_13716,N_9823,N_6891);
or U13717 (N_13717,N_6747,N_8594);
nand U13718 (N_13718,N_5553,N_7952);
nor U13719 (N_13719,N_6989,N_8065);
nor U13720 (N_13720,N_9721,N_6065);
or U13721 (N_13721,N_7910,N_5063);
or U13722 (N_13722,N_6096,N_6952);
nor U13723 (N_13723,N_8674,N_6265);
nor U13724 (N_13724,N_8071,N_7025);
and U13725 (N_13725,N_9405,N_6702);
nand U13726 (N_13726,N_9488,N_9995);
nand U13727 (N_13727,N_5337,N_7273);
or U13728 (N_13728,N_7953,N_5460);
nand U13729 (N_13729,N_9564,N_6979);
or U13730 (N_13730,N_9130,N_5276);
nor U13731 (N_13731,N_8606,N_5661);
nor U13732 (N_13732,N_9603,N_8983);
nand U13733 (N_13733,N_7759,N_6962);
nand U13734 (N_13734,N_9841,N_8015);
or U13735 (N_13735,N_5109,N_8469);
and U13736 (N_13736,N_6115,N_6675);
nand U13737 (N_13737,N_8709,N_6533);
nand U13738 (N_13738,N_9959,N_9673);
nor U13739 (N_13739,N_6211,N_9426);
nand U13740 (N_13740,N_5265,N_8938);
nand U13741 (N_13741,N_5730,N_7101);
nor U13742 (N_13742,N_7786,N_7067);
nand U13743 (N_13743,N_8423,N_6996);
and U13744 (N_13744,N_7149,N_6642);
or U13745 (N_13745,N_5206,N_5327);
nand U13746 (N_13746,N_9578,N_9805);
or U13747 (N_13747,N_8734,N_6931);
nand U13748 (N_13748,N_7545,N_8852);
and U13749 (N_13749,N_8457,N_9942);
nor U13750 (N_13750,N_7741,N_5874);
nand U13751 (N_13751,N_7538,N_7447);
nor U13752 (N_13752,N_5718,N_6044);
nor U13753 (N_13753,N_5960,N_7489);
and U13754 (N_13754,N_7051,N_5265);
or U13755 (N_13755,N_9279,N_6583);
and U13756 (N_13756,N_5240,N_7784);
and U13757 (N_13757,N_5757,N_6196);
nor U13758 (N_13758,N_5208,N_8262);
nor U13759 (N_13759,N_5120,N_7203);
nand U13760 (N_13760,N_7988,N_6556);
or U13761 (N_13761,N_6669,N_9451);
nor U13762 (N_13762,N_7861,N_5856);
nor U13763 (N_13763,N_5254,N_7278);
nor U13764 (N_13764,N_7356,N_9038);
nand U13765 (N_13765,N_6687,N_6986);
and U13766 (N_13766,N_5777,N_8444);
nand U13767 (N_13767,N_9946,N_6428);
nand U13768 (N_13768,N_9546,N_7147);
nor U13769 (N_13769,N_5481,N_8218);
xnor U13770 (N_13770,N_5016,N_7310);
or U13771 (N_13771,N_6511,N_9685);
or U13772 (N_13772,N_9877,N_5205);
or U13773 (N_13773,N_9100,N_7002);
and U13774 (N_13774,N_9204,N_5679);
nor U13775 (N_13775,N_9001,N_9738);
nor U13776 (N_13776,N_9060,N_7999);
and U13777 (N_13777,N_6937,N_7649);
or U13778 (N_13778,N_7983,N_6864);
nand U13779 (N_13779,N_5453,N_9313);
or U13780 (N_13780,N_9875,N_9575);
nor U13781 (N_13781,N_8377,N_7324);
nand U13782 (N_13782,N_6757,N_8475);
nand U13783 (N_13783,N_5033,N_8462);
nand U13784 (N_13784,N_9898,N_6290);
and U13785 (N_13785,N_5060,N_7982);
nand U13786 (N_13786,N_9913,N_9620);
nand U13787 (N_13787,N_5659,N_7460);
and U13788 (N_13788,N_5925,N_5778);
nand U13789 (N_13789,N_9343,N_8729);
nand U13790 (N_13790,N_6482,N_5445);
nor U13791 (N_13791,N_7263,N_8315);
or U13792 (N_13792,N_6467,N_6133);
or U13793 (N_13793,N_5069,N_9218);
nor U13794 (N_13794,N_6224,N_9950);
or U13795 (N_13795,N_5266,N_7201);
or U13796 (N_13796,N_9985,N_6412);
or U13797 (N_13797,N_9304,N_6885);
or U13798 (N_13798,N_8832,N_5242);
nand U13799 (N_13799,N_6010,N_9506);
or U13800 (N_13800,N_6706,N_6360);
and U13801 (N_13801,N_7931,N_7789);
and U13802 (N_13802,N_7325,N_7922);
nor U13803 (N_13803,N_6220,N_5092);
and U13804 (N_13804,N_6383,N_9207);
and U13805 (N_13805,N_9078,N_5052);
and U13806 (N_13806,N_8280,N_9728);
nand U13807 (N_13807,N_8121,N_7584);
nand U13808 (N_13808,N_9899,N_9808);
nand U13809 (N_13809,N_5801,N_6714);
nand U13810 (N_13810,N_8708,N_5775);
nand U13811 (N_13811,N_5634,N_9275);
and U13812 (N_13812,N_8671,N_5833);
or U13813 (N_13813,N_7122,N_9329);
or U13814 (N_13814,N_9606,N_6793);
nor U13815 (N_13815,N_6705,N_8136);
or U13816 (N_13816,N_9980,N_9621);
nand U13817 (N_13817,N_8052,N_5130);
or U13818 (N_13818,N_6318,N_7040);
nand U13819 (N_13819,N_7100,N_8689);
nor U13820 (N_13820,N_9339,N_8225);
nor U13821 (N_13821,N_7063,N_6581);
nand U13822 (N_13822,N_9014,N_7917);
or U13823 (N_13823,N_6701,N_5858);
nand U13824 (N_13824,N_9257,N_7067);
and U13825 (N_13825,N_8819,N_5959);
and U13826 (N_13826,N_6817,N_8828);
nand U13827 (N_13827,N_8196,N_8020);
and U13828 (N_13828,N_8346,N_7858);
nand U13829 (N_13829,N_8928,N_7246);
or U13830 (N_13830,N_8988,N_6699);
nor U13831 (N_13831,N_9948,N_9098);
nand U13832 (N_13832,N_7293,N_9922);
nor U13833 (N_13833,N_7860,N_6160);
nand U13834 (N_13834,N_7842,N_7227);
and U13835 (N_13835,N_5175,N_7855);
nand U13836 (N_13836,N_7563,N_9830);
nor U13837 (N_13837,N_9629,N_7974);
and U13838 (N_13838,N_8563,N_8175);
or U13839 (N_13839,N_6432,N_5624);
nor U13840 (N_13840,N_6457,N_9349);
xnor U13841 (N_13841,N_8665,N_9632);
and U13842 (N_13842,N_9609,N_5688);
nor U13843 (N_13843,N_9907,N_6535);
or U13844 (N_13844,N_8352,N_7505);
nand U13845 (N_13845,N_9638,N_7607);
nand U13846 (N_13846,N_5614,N_8420);
and U13847 (N_13847,N_9425,N_8868);
nand U13848 (N_13848,N_5723,N_7322);
nor U13849 (N_13849,N_5865,N_7207);
or U13850 (N_13850,N_7672,N_7048);
xor U13851 (N_13851,N_8279,N_6220);
nand U13852 (N_13852,N_9729,N_8840);
nor U13853 (N_13853,N_9222,N_8276);
nand U13854 (N_13854,N_9346,N_5889);
nor U13855 (N_13855,N_5648,N_6327);
nor U13856 (N_13856,N_6574,N_9368);
nand U13857 (N_13857,N_7185,N_5795);
nor U13858 (N_13858,N_8682,N_9249);
and U13859 (N_13859,N_6733,N_7813);
and U13860 (N_13860,N_9733,N_7859);
and U13861 (N_13861,N_8842,N_5318);
nor U13862 (N_13862,N_5335,N_7882);
and U13863 (N_13863,N_9723,N_8150);
nand U13864 (N_13864,N_6474,N_9476);
and U13865 (N_13865,N_8478,N_9083);
nand U13866 (N_13866,N_8379,N_7263);
nor U13867 (N_13867,N_6453,N_6394);
nand U13868 (N_13868,N_7723,N_5549);
or U13869 (N_13869,N_7960,N_7704);
or U13870 (N_13870,N_8396,N_5963);
nand U13871 (N_13871,N_9304,N_9613);
nor U13872 (N_13872,N_9788,N_9871);
nand U13873 (N_13873,N_7225,N_9037);
xor U13874 (N_13874,N_5783,N_6023);
nor U13875 (N_13875,N_5642,N_9909);
or U13876 (N_13876,N_9446,N_9294);
nand U13877 (N_13877,N_7470,N_8467);
nand U13878 (N_13878,N_9138,N_8411);
nor U13879 (N_13879,N_7893,N_7163);
or U13880 (N_13880,N_8473,N_6062);
nor U13881 (N_13881,N_8529,N_7138);
nor U13882 (N_13882,N_8172,N_8376);
or U13883 (N_13883,N_7975,N_6118);
and U13884 (N_13884,N_8219,N_5478);
or U13885 (N_13885,N_8900,N_9450);
or U13886 (N_13886,N_8070,N_5539);
and U13887 (N_13887,N_8719,N_7230);
nor U13888 (N_13888,N_6193,N_9283);
nand U13889 (N_13889,N_7340,N_7995);
nor U13890 (N_13890,N_9608,N_9206);
xor U13891 (N_13891,N_9989,N_7826);
and U13892 (N_13892,N_9994,N_9177);
or U13893 (N_13893,N_9196,N_7221);
and U13894 (N_13894,N_9051,N_5292);
nand U13895 (N_13895,N_7397,N_5118);
xor U13896 (N_13896,N_9707,N_5420);
or U13897 (N_13897,N_9456,N_7247);
or U13898 (N_13898,N_6645,N_8973);
nor U13899 (N_13899,N_5365,N_8047);
or U13900 (N_13900,N_8090,N_5447);
and U13901 (N_13901,N_5952,N_5633);
or U13902 (N_13902,N_6903,N_5058);
and U13903 (N_13903,N_5161,N_9965);
or U13904 (N_13904,N_9357,N_9020);
xor U13905 (N_13905,N_6936,N_8369);
nor U13906 (N_13906,N_5043,N_6033);
nand U13907 (N_13907,N_8349,N_6872);
nor U13908 (N_13908,N_7091,N_8547);
and U13909 (N_13909,N_7155,N_8173);
xor U13910 (N_13910,N_7074,N_6929);
or U13911 (N_13911,N_8350,N_5150);
or U13912 (N_13912,N_6442,N_8672);
and U13913 (N_13913,N_7584,N_8142);
nand U13914 (N_13914,N_9615,N_9540);
and U13915 (N_13915,N_7688,N_7873);
and U13916 (N_13916,N_8686,N_9814);
nand U13917 (N_13917,N_7005,N_8739);
and U13918 (N_13918,N_7901,N_6224);
and U13919 (N_13919,N_5765,N_5823);
or U13920 (N_13920,N_8226,N_9228);
nor U13921 (N_13921,N_6855,N_8175);
nand U13922 (N_13922,N_8811,N_8883);
or U13923 (N_13923,N_6482,N_9731);
nor U13924 (N_13924,N_6161,N_9083);
nand U13925 (N_13925,N_5280,N_6739);
and U13926 (N_13926,N_7093,N_6694);
and U13927 (N_13927,N_9738,N_7533);
or U13928 (N_13928,N_8188,N_6904);
nor U13929 (N_13929,N_8137,N_9305);
nand U13930 (N_13930,N_9913,N_8427);
and U13931 (N_13931,N_5189,N_9686);
nand U13932 (N_13932,N_6761,N_7230);
nor U13933 (N_13933,N_9068,N_7500);
and U13934 (N_13934,N_7712,N_8953);
or U13935 (N_13935,N_7286,N_9333);
nand U13936 (N_13936,N_9717,N_9377);
or U13937 (N_13937,N_6535,N_6220);
or U13938 (N_13938,N_8595,N_7368);
or U13939 (N_13939,N_9850,N_9214);
nor U13940 (N_13940,N_9840,N_9081);
and U13941 (N_13941,N_6252,N_8290);
nor U13942 (N_13942,N_6264,N_9569);
or U13943 (N_13943,N_9616,N_8744);
or U13944 (N_13944,N_7038,N_6401);
or U13945 (N_13945,N_5185,N_7284);
nor U13946 (N_13946,N_8574,N_5224);
nand U13947 (N_13947,N_7612,N_8700);
and U13948 (N_13948,N_5124,N_6639);
or U13949 (N_13949,N_6894,N_5306);
and U13950 (N_13950,N_5780,N_8278);
xor U13951 (N_13951,N_5075,N_6139);
or U13952 (N_13952,N_8040,N_8927);
nor U13953 (N_13953,N_7139,N_5245);
nand U13954 (N_13954,N_7592,N_9316);
nor U13955 (N_13955,N_6385,N_5113);
nor U13956 (N_13956,N_6016,N_6438);
nor U13957 (N_13957,N_9777,N_9285);
and U13958 (N_13958,N_5605,N_5521);
and U13959 (N_13959,N_5517,N_6268);
nor U13960 (N_13960,N_6808,N_8931);
or U13961 (N_13961,N_9680,N_7481);
or U13962 (N_13962,N_9430,N_7049);
nand U13963 (N_13963,N_6276,N_9931);
and U13964 (N_13964,N_7505,N_6243);
nand U13965 (N_13965,N_7378,N_9744);
and U13966 (N_13966,N_8322,N_5193);
nand U13967 (N_13967,N_6733,N_5451);
nor U13968 (N_13968,N_9014,N_9096);
nand U13969 (N_13969,N_6704,N_7904);
nand U13970 (N_13970,N_8928,N_8767);
or U13971 (N_13971,N_6848,N_7120);
or U13972 (N_13972,N_5038,N_9795);
and U13973 (N_13973,N_7339,N_6527);
nand U13974 (N_13974,N_6566,N_8635);
nor U13975 (N_13975,N_7605,N_7331);
nand U13976 (N_13976,N_5308,N_6066);
nor U13977 (N_13977,N_7895,N_5866);
or U13978 (N_13978,N_6124,N_7234);
or U13979 (N_13979,N_6121,N_9884);
or U13980 (N_13980,N_8892,N_7753);
nor U13981 (N_13981,N_8614,N_9069);
nor U13982 (N_13982,N_8081,N_5149);
nand U13983 (N_13983,N_5687,N_5012);
nor U13984 (N_13984,N_8123,N_5190);
nand U13985 (N_13985,N_5643,N_9367);
or U13986 (N_13986,N_6558,N_6210);
nor U13987 (N_13987,N_6157,N_5396);
or U13988 (N_13988,N_7015,N_5754);
nand U13989 (N_13989,N_8310,N_8634);
and U13990 (N_13990,N_9060,N_6662);
or U13991 (N_13991,N_5193,N_5914);
or U13992 (N_13992,N_7687,N_5652);
or U13993 (N_13993,N_7303,N_9053);
nand U13994 (N_13994,N_9144,N_7702);
or U13995 (N_13995,N_8457,N_6887);
nor U13996 (N_13996,N_8058,N_6834);
and U13997 (N_13997,N_8956,N_9460);
or U13998 (N_13998,N_5579,N_9270);
or U13999 (N_13999,N_9117,N_6736);
nor U14000 (N_14000,N_6419,N_7940);
nor U14001 (N_14001,N_5047,N_9445);
or U14002 (N_14002,N_5626,N_8571);
nand U14003 (N_14003,N_5139,N_9864);
or U14004 (N_14004,N_8882,N_5032);
and U14005 (N_14005,N_9768,N_7156);
nor U14006 (N_14006,N_8238,N_9559);
nor U14007 (N_14007,N_5437,N_6715);
nor U14008 (N_14008,N_8701,N_7094);
and U14009 (N_14009,N_7682,N_9871);
and U14010 (N_14010,N_9136,N_8289);
nand U14011 (N_14011,N_8346,N_9703);
and U14012 (N_14012,N_5013,N_7583);
nor U14013 (N_14013,N_5174,N_6553);
nor U14014 (N_14014,N_9596,N_5994);
and U14015 (N_14015,N_6847,N_5693);
or U14016 (N_14016,N_9467,N_8228);
or U14017 (N_14017,N_7995,N_6449);
xor U14018 (N_14018,N_7013,N_5582);
nor U14019 (N_14019,N_5456,N_9991);
nor U14020 (N_14020,N_9289,N_9744);
nor U14021 (N_14021,N_6549,N_7653);
nor U14022 (N_14022,N_8653,N_6615);
nor U14023 (N_14023,N_8867,N_6355);
and U14024 (N_14024,N_6117,N_6544);
or U14025 (N_14025,N_5226,N_9701);
or U14026 (N_14026,N_6410,N_9076);
or U14027 (N_14027,N_7757,N_7283);
or U14028 (N_14028,N_6235,N_9198);
and U14029 (N_14029,N_5363,N_9448);
nand U14030 (N_14030,N_6921,N_6020);
nor U14031 (N_14031,N_9507,N_7123);
or U14032 (N_14032,N_9054,N_7597);
and U14033 (N_14033,N_6443,N_6065);
xor U14034 (N_14034,N_5148,N_7738);
or U14035 (N_14035,N_6452,N_7069);
or U14036 (N_14036,N_5897,N_6084);
nand U14037 (N_14037,N_7517,N_6706);
nand U14038 (N_14038,N_6089,N_7920);
or U14039 (N_14039,N_7378,N_8337);
or U14040 (N_14040,N_9969,N_8809);
nand U14041 (N_14041,N_6675,N_8062);
or U14042 (N_14042,N_5950,N_8086);
nor U14043 (N_14043,N_9452,N_5578);
or U14044 (N_14044,N_8317,N_7017);
nor U14045 (N_14045,N_7944,N_9525);
nor U14046 (N_14046,N_8333,N_7545);
and U14047 (N_14047,N_5783,N_5057);
xnor U14048 (N_14048,N_7228,N_6994);
nor U14049 (N_14049,N_6437,N_9345);
nor U14050 (N_14050,N_9697,N_6858);
or U14051 (N_14051,N_5806,N_5013);
and U14052 (N_14052,N_5639,N_8430);
nand U14053 (N_14053,N_7827,N_9941);
nand U14054 (N_14054,N_7379,N_7121);
and U14055 (N_14055,N_5869,N_5277);
and U14056 (N_14056,N_5096,N_6851);
nand U14057 (N_14057,N_6592,N_8677);
nor U14058 (N_14058,N_9856,N_8576);
and U14059 (N_14059,N_5253,N_5689);
and U14060 (N_14060,N_5733,N_8077);
nor U14061 (N_14061,N_7208,N_7759);
nand U14062 (N_14062,N_8770,N_7313);
nor U14063 (N_14063,N_6897,N_5186);
and U14064 (N_14064,N_5221,N_5259);
and U14065 (N_14065,N_9103,N_9728);
nor U14066 (N_14066,N_5551,N_6713);
nand U14067 (N_14067,N_8259,N_8397);
or U14068 (N_14068,N_7302,N_9741);
nand U14069 (N_14069,N_9855,N_8707);
or U14070 (N_14070,N_9641,N_6771);
and U14071 (N_14071,N_9813,N_8701);
nor U14072 (N_14072,N_7190,N_5383);
nor U14073 (N_14073,N_5507,N_9146);
or U14074 (N_14074,N_7684,N_9828);
and U14075 (N_14075,N_8487,N_6256);
nand U14076 (N_14076,N_5534,N_5787);
nor U14077 (N_14077,N_7314,N_5300);
nor U14078 (N_14078,N_6401,N_8587);
nand U14079 (N_14079,N_5287,N_8045);
nand U14080 (N_14080,N_7104,N_6796);
or U14081 (N_14081,N_9916,N_6642);
nor U14082 (N_14082,N_8625,N_8773);
nand U14083 (N_14083,N_7792,N_8498);
and U14084 (N_14084,N_5385,N_8876);
nor U14085 (N_14085,N_8382,N_6668);
and U14086 (N_14086,N_9067,N_8236);
nand U14087 (N_14087,N_6338,N_6816);
or U14088 (N_14088,N_8440,N_8645);
nand U14089 (N_14089,N_7934,N_5230);
and U14090 (N_14090,N_9159,N_6651);
nand U14091 (N_14091,N_9944,N_6018);
nor U14092 (N_14092,N_6150,N_8186);
nor U14093 (N_14093,N_8118,N_8603);
or U14094 (N_14094,N_9927,N_9945);
and U14095 (N_14095,N_9909,N_8068);
or U14096 (N_14096,N_9310,N_6794);
and U14097 (N_14097,N_7238,N_6707);
nor U14098 (N_14098,N_5223,N_7791);
or U14099 (N_14099,N_6642,N_6852);
nand U14100 (N_14100,N_5635,N_5469);
nand U14101 (N_14101,N_9454,N_5819);
or U14102 (N_14102,N_9785,N_7825);
nand U14103 (N_14103,N_8587,N_6304);
or U14104 (N_14104,N_6420,N_9755);
nand U14105 (N_14105,N_9955,N_7405);
nor U14106 (N_14106,N_8168,N_7165);
nor U14107 (N_14107,N_8461,N_9080);
or U14108 (N_14108,N_6646,N_6949);
or U14109 (N_14109,N_9816,N_6646);
and U14110 (N_14110,N_6762,N_5069);
or U14111 (N_14111,N_9044,N_8232);
nand U14112 (N_14112,N_7009,N_7917);
and U14113 (N_14113,N_5486,N_6321);
nor U14114 (N_14114,N_6623,N_9105);
and U14115 (N_14115,N_5126,N_7030);
nand U14116 (N_14116,N_8136,N_7201);
nor U14117 (N_14117,N_6606,N_9464);
or U14118 (N_14118,N_6567,N_7266);
nand U14119 (N_14119,N_7193,N_5007);
or U14120 (N_14120,N_7921,N_6654);
and U14121 (N_14121,N_5707,N_9473);
or U14122 (N_14122,N_5503,N_5837);
or U14123 (N_14123,N_9051,N_7253);
nand U14124 (N_14124,N_8767,N_6395);
and U14125 (N_14125,N_5428,N_5026);
or U14126 (N_14126,N_5046,N_8108);
or U14127 (N_14127,N_7123,N_8751);
or U14128 (N_14128,N_9323,N_6190);
nor U14129 (N_14129,N_5590,N_8337);
and U14130 (N_14130,N_5562,N_7318);
or U14131 (N_14131,N_6550,N_5734);
nor U14132 (N_14132,N_9106,N_8252);
or U14133 (N_14133,N_7525,N_8273);
and U14134 (N_14134,N_6349,N_5349);
nand U14135 (N_14135,N_8514,N_9399);
nor U14136 (N_14136,N_8717,N_5313);
and U14137 (N_14137,N_7676,N_8823);
nor U14138 (N_14138,N_6052,N_8837);
and U14139 (N_14139,N_6751,N_6809);
nand U14140 (N_14140,N_6772,N_6485);
nor U14141 (N_14141,N_5247,N_5636);
nand U14142 (N_14142,N_5543,N_6067);
nand U14143 (N_14143,N_5049,N_7817);
nand U14144 (N_14144,N_7367,N_5320);
nand U14145 (N_14145,N_5033,N_6820);
nand U14146 (N_14146,N_6982,N_9801);
and U14147 (N_14147,N_9290,N_5499);
or U14148 (N_14148,N_7890,N_7796);
nor U14149 (N_14149,N_9116,N_6659);
nand U14150 (N_14150,N_9365,N_9780);
xnor U14151 (N_14151,N_6950,N_6928);
nand U14152 (N_14152,N_6700,N_5902);
and U14153 (N_14153,N_5701,N_5931);
or U14154 (N_14154,N_7643,N_7996);
nor U14155 (N_14155,N_7016,N_8886);
nand U14156 (N_14156,N_6564,N_7500);
nand U14157 (N_14157,N_5870,N_7242);
or U14158 (N_14158,N_6701,N_6364);
or U14159 (N_14159,N_6296,N_6355);
nor U14160 (N_14160,N_6899,N_7980);
and U14161 (N_14161,N_6286,N_5220);
and U14162 (N_14162,N_5732,N_9553);
or U14163 (N_14163,N_8011,N_6316);
nand U14164 (N_14164,N_9159,N_7982);
nand U14165 (N_14165,N_6155,N_8115);
or U14166 (N_14166,N_5039,N_8949);
and U14167 (N_14167,N_6588,N_9876);
or U14168 (N_14168,N_5359,N_5647);
or U14169 (N_14169,N_6312,N_6412);
or U14170 (N_14170,N_8757,N_8055);
and U14171 (N_14171,N_9469,N_6382);
nand U14172 (N_14172,N_6024,N_8232);
or U14173 (N_14173,N_5197,N_6393);
nor U14174 (N_14174,N_5482,N_8693);
or U14175 (N_14175,N_5454,N_9800);
nor U14176 (N_14176,N_6387,N_9288);
or U14177 (N_14177,N_5488,N_8516);
or U14178 (N_14178,N_9692,N_7431);
and U14179 (N_14179,N_7737,N_9378);
or U14180 (N_14180,N_9250,N_8012);
nand U14181 (N_14181,N_5142,N_9024);
or U14182 (N_14182,N_5387,N_9803);
nand U14183 (N_14183,N_7536,N_8304);
nor U14184 (N_14184,N_9856,N_8050);
and U14185 (N_14185,N_8229,N_6674);
nand U14186 (N_14186,N_9564,N_6015);
nand U14187 (N_14187,N_9423,N_5584);
or U14188 (N_14188,N_6356,N_7876);
or U14189 (N_14189,N_7776,N_6492);
and U14190 (N_14190,N_8282,N_9467);
and U14191 (N_14191,N_5899,N_9793);
nand U14192 (N_14192,N_9340,N_7478);
and U14193 (N_14193,N_7146,N_5581);
nand U14194 (N_14194,N_9285,N_6510);
nand U14195 (N_14195,N_5866,N_8840);
and U14196 (N_14196,N_8840,N_6657);
or U14197 (N_14197,N_5182,N_8282);
and U14198 (N_14198,N_9300,N_8198);
nor U14199 (N_14199,N_6454,N_5615);
nand U14200 (N_14200,N_6390,N_5465);
nand U14201 (N_14201,N_5294,N_7487);
and U14202 (N_14202,N_9520,N_8420);
and U14203 (N_14203,N_9482,N_5005);
nand U14204 (N_14204,N_7820,N_5648);
nand U14205 (N_14205,N_9399,N_7865);
nand U14206 (N_14206,N_9538,N_8319);
or U14207 (N_14207,N_7494,N_9736);
or U14208 (N_14208,N_6997,N_5291);
or U14209 (N_14209,N_5264,N_9885);
and U14210 (N_14210,N_5744,N_5281);
nor U14211 (N_14211,N_9410,N_6255);
nor U14212 (N_14212,N_9975,N_9283);
and U14213 (N_14213,N_7995,N_9324);
nor U14214 (N_14214,N_7378,N_6349);
or U14215 (N_14215,N_5908,N_5005);
or U14216 (N_14216,N_6786,N_8155);
and U14217 (N_14217,N_7502,N_6478);
nor U14218 (N_14218,N_6095,N_5186);
or U14219 (N_14219,N_7107,N_9955);
nand U14220 (N_14220,N_6371,N_7097);
or U14221 (N_14221,N_8966,N_8951);
or U14222 (N_14222,N_8825,N_7658);
and U14223 (N_14223,N_7812,N_8154);
and U14224 (N_14224,N_5443,N_5647);
nand U14225 (N_14225,N_8493,N_9249);
nand U14226 (N_14226,N_9379,N_7686);
nor U14227 (N_14227,N_8877,N_8376);
or U14228 (N_14228,N_6565,N_7307);
nor U14229 (N_14229,N_6653,N_9626);
nand U14230 (N_14230,N_5549,N_5069);
or U14231 (N_14231,N_8548,N_6424);
nand U14232 (N_14232,N_9865,N_6440);
nand U14233 (N_14233,N_5323,N_5373);
or U14234 (N_14234,N_8871,N_8939);
nand U14235 (N_14235,N_6265,N_6434);
or U14236 (N_14236,N_9825,N_5246);
nor U14237 (N_14237,N_9085,N_9991);
or U14238 (N_14238,N_6782,N_9460);
nand U14239 (N_14239,N_9277,N_5351);
nor U14240 (N_14240,N_6427,N_6170);
nor U14241 (N_14241,N_5353,N_6785);
or U14242 (N_14242,N_5378,N_5857);
nand U14243 (N_14243,N_8305,N_5893);
nand U14244 (N_14244,N_8019,N_7088);
or U14245 (N_14245,N_5651,N_8916);
nor U14246 (N_14246,N_8820,N_8065);
nor U14247 (N_14247,N_7506,N_6682);
or U14248 (N_14248,N_9031,N_9245);
nor U14249 (N_14249,N_8463,N_5980);
nor U14250 (N_14250,N_9671,N_5548);
or U14251 (N_14251,N_5208,N_5578);
or U14252 (N_14252,N_8129,N_7982);
and U14253 (N_14253,N_9930,N_7666);
nand U14254 (N_14254,N_9913,N_6363);
nand U14255 (N_14255,N_8901,N_8341);
nor U14256 (N_14256,N_7190,N_8203);
nand U14257 (N_14257,N_6405,N_9592);
or U14258 (N_14258,N_6028,N_9854);
nand U14259 (N_14259,N_9627,N_9199);
and U14260 (N_14260,N_5269,N_5605);
nor U14261 (N_14261,N_7324,N_8595);
and U14262 (N_14262,N_8759,N_6390);
and U14263 (N_14263,N_9781,N_5931);
nor U14264 (N_14264,N_5204,N_7066);
nand U14265 (N_14265,N_8450,N_9412);
nor U14266 (N_14266,N_5678,N_8325);
nor U14267 (N_14267,N_5716,N_6757);
or U14268 (N_14268,N_7581,N_5748);
nand U14269 (N_14269,N_6974,N_9071);
nand U14270 (N_14270,N_5509,N_7281);
or U14271 (N_14271,N_9282,N_9930);
or U14272 (N_14272,N_5237,N_8927);
nand U14273 (N_14273,N_9881,N_7425);
and U14274 (N_14274,N_7592,N_7366);
and U14275 (N_14275,N_7622,N_7173);
nand U14276 (N_14276,N_7484,N_9937);
nand U14277 (N_14277,N_9612,N_9049);
or U14278 (N_14278,N_6810,N_8891);
and U14279 (N_14279,N_9969,N_8356);
nand U14280 (N_14280,N_8652,N_6901);
and U14281 (N_14281,N_8894,N_9970);
or U14282 (N_14282,N_6486,N_8373);
and U14283 (N_14283,N_9148,N_7370);
or U14284 (N_14284,N_5869,N_8988);
and U14285 (N_14285,N_6655,N_9314);
or U14286 (N_14286,N_8743,N_6866);
nor U14287 (N_14287,N_6333,N_7202);
and U14288 (N_14288,N_6080,N_9637);
nand U14289 (N_14289,N_9229,N_6010);
and U14290 (N_14290,N_5890,N_7818);
nand U14291 (N_14291,N_8429,N_7215);
nand U14292 (N_14292,N_5234,N_9557);
nor U14293 (N_14293,N_6608,N_5043);
and U14294 (N_14294,N_6628,N_5623);
nor U14295 (N_14295,N_9551,N_5030);
or U14296 (N_14296,N_6382,N_7324);
and U14297 (N_14297,N_8576,N_5372);
and U14298 (N_14298,N_7862,N_6053);
and U14299 (N_14299,N_6078,N_6710);
or U14300 (N_14300,N_6345,N_9674);
nor U14301 (N_14301,N_5703,N_8790);
and U14302 (N_14302,N_9529,N_6468);
and U14303 (N_14303,N_9848,N_6343);
and U14304 (N_14304,N_5034,N_7004);
and U14305 (N_14305,N_5161,N_6322);
and U14306 (N_14306,N_6362,N_5209);
or U14307 (N_14307,N_9965,N_6676);
or U14308 (N_14308,N_8853,N_7425);
nor U14309 (N_14309,N_6969,N_5014);
nand U14310 (N_14310,N_6951,N_9618);
nand U14311 (N_14311,N_9792,N_5654);
and U14312 (N_14312,N_8547,N_6662);
and U14313 (N_14313,N_5466,N_5903);
nand U14314 (N_14314,N_9116,N_8328);
or U14315 (N_14315,N_6269,N_8136);
or U14316 (N_14316,N_8171,N_8427);
or U14317 (N_14317,N_7513,N_6676);
nand U14318 (N_14318,N_8567,N_9463);
and U14319 (N_14319,N_6677,N_6832);
nand U14320 (N_14320,N_6094,N_7884);
and U14321 (N_14321,N_8766,N_6695);
and U14322 (N_14322,N_9259,N_8818);
or U14323 (N_14323,N_9823,N_9019);
or U14324 (N_14324,N_7670,N_9419);
or U14325 (N_14325,N_5349,N_9260);
nor U14326 (N_14326,N_6152,N_8928);
nand U14327 (N_14327,N_6429,N_6304);
or U14328 (N_14328,N_9340,N_5925);
nor U14329 (N_14329,N_6847,N_9993);
nand U14330 (N_14330,N_7304,N_8053);
nor U14331 (N_14331,N_8711,N_9960);
or U14332 (N_14332,N_8130,N_6041);
or U14333 (N_14333,N_6737,N_9544);
and U14334 (N_14334,N_9902,N_9468);
nor U14335 (N_14335,N_8003,N_7717);
and U14336 (N_14336,N_8282,N_9795);
or U14337 (N_14337,N_8167,N_6600);
and U14338 (N_14338,N_8272,N_8394);
or U14339 (N_14339,N_9578,N_5334);
and U14340 (N_14340,N_6002,N_5991);
nor U14341 (N_14341,N_9240,N_8435);
nand U14342 (N_14342,N_6233,N_7156);
or U14343 (N_14343,N_5364,N_7859);
nor U14344 (N_14344,N_7393,N_9487);
nand U14345 (N_14345,N_9851,N_5316);
or U14346 (N_14346,N_6238,N_9683);
and U14347 (N_14347,N_6734,N_9027);
and U14348 (N_14348,N_6735,N_6885);
nor U14349 (N_14349,N_6449,N_5438);
or U14350 (N_14350,N_7092,N_6551);
or U14351 (N_14351,N_9421,N_7527);
nand U14352 (N_14352,N_9989,N_6050);
or U14353 (N_14353,N_5176,N_9918);
nand U14354 (N_14354,N_6833,N_6193);
and U14355 (N_14355,N_7572,N_8742);
nand U14356 (N_14356,N_7984,N_8084);
nor U14357 (N_14357,N_8412,N_9450);
nand U14358 (N_14358,N_8911,N_7811);
and U14359 (N_14359,N_8893,N_6654);
and U14360 (N_14360,N_5274,N_8083);
and U14361 (N_14361,N_7423,N_9199);
nand U14362 (N_14362,N_5890,N_9374);
nor U14363 (N_14363,N_5946,N_6348);
nand U14364 (N_14364,N_7272,N_7108);
nor U14365 (N_14365,N_5640,N_6592);
and U14366 (N_14366,N_5342,N_7560);
nand U14367 (N_14367,N_6540,N_8492);
nand U14368 (N_14368,N_7606,N_8673);
or U14369 (N_14369,N_5941,N_8074);
nor U14370 (N_14370,N_9830,N_6751);
or U14371 (N_14371,N_9785,N_8044);
or U14372 (N_14372,N_6101,N_5152);
nor U14373 (N_14373,N_6127,N_7538);
or U14374 (N_14374,N_7182,N_9399);
nor U14375 (N_14375,N_7917,N_9495);
and U14376 (N_14376,N_7372,N_7220);
nand U14377 (N_14377,N_9744,N_5167);
and U14378 (N_14378,N_7038,N_7486);
or U14379 (N_14379,N_8490,N_5326);
or U14380 (N_14380,N_8391,N_9652);
nor U14381 (N_14381,N_7781,N_9845);
and U14382 (N_14382,N_7751,N_7641);
and U14383 (N_14383,N_8257,N_6207);
nor U14384 (N_14384,N_6109,N_6066);
nor U14385 (N_14385,N_5443,N_5949);
or U14386 (N_14386,N_6634,N_7607);
or U14387 (N_14387,N_8700,N_8118);
and U14388 (N_14388,N_8382,N_6393);
or U14389 (N_14389,N_5840,N_9677);
nor U14390 (N_14390,N_7283,N_9668);
or U14391 (N_14391,N_9821,N_9318);
nor U14392 (N_14392,N_5188,N_8112);
nor U14393 (N_14393,N_8773,N_8551);
nor U14394 (N_14394,N_8288,N_9192);
nand U14395 (N_14395,N_7358,N_5718);
xnor U14396 (N_14396,N_5701,N_5114);
nor U14397 (N_14397,N_9423,N_8367);
nand U14398 (N_14398,N_9317,N_6912);
or U14399 (N_14399,N_6085,N_5972);
or U14400 (N_14400,N_5030,N_8127);
and U14401 (N_14401,N_7234,N_5811);
nor U14402 (N_14402,N_7641,N_8794);
nand U14403 (N_14403,N_6451,N_8989);
and U14404 (N_14404,N_7290,N_9252);
nand U14405 (N_14405,N_5293,N_5800);
and U14406 (N_14406,N_7635,N_8919);
or U14407 (N_14407,N_6499,N_5223);
and U14408 (N_14408,N_6518,N_6995);
or U14409 (N_14409,N_7321,N_5304);
and U14410 (N_14410,N_7802,N_5702);
and U14411 (N_14411,N_9683,N_7289);
or U14412 (N_14412,N_6432,N_8197);
nand U14413 (N_14413,N_9574,N_6314);
or U14414 (N_14414,N_7329,N_6945);
or U14415 (N_14415,N_6834,N_8663);
nor U14416 (N_14416,N_5216,N_5455);
or U14417 (N_14417,N_9582,N_6976);
nand U14418 (N_14418,N_5971,N_7369);
or U14419 (N_14419,N_7376,N_7048);
and U14420 (N_14420,N_7306,N_6935);
or U14421 (N_14421,N_8488,N_5356);
or U14422 (N_14422,N_9627,N_8003);
nand U14423 (N_14423,N_6155,N_5178);
or U14424 (N_14424,N_8902,N_9326);
xor U14425 (N_14425,N_5141,N_7840);
nand U14426 (N_14426,N_6250,N_8183);
nand U14427 (N_14427,N_5777,N_7990);
nand U14428 (N_14428,N_7809,N_6372);
nand U14429 (N_14429,N_6602,N_6148);
xnor U14430 (N_14430,N_6406,N_9295);
nand U14431 (N_14431,N_5953,N_8491);
and U14432 (N_14432,N_8518,N_7418);
nor U14433 (N_14433,N_8365,N_5092);
nand U14434 (N_14434,N_5837,N_5571);
and U14435 (N_14435,N_6541,N_8416);
and U14436 (N_14436,N_9104,N_5120);
or U14437 (N_14437,N_8645,N_6290);
nand U14438 (N_14438,N_9911,N_5722);
nand U14439 (N_14439,N_7504,N_8798);
nor U14440 (N_14440,N_6154,N_8511);
nor U14441 (N_14441,N_7604,N_8117);
or U14442 (N_14442,N_5938,N_5051);
nor U14443 (N_14443,N_6166,N_8218);
nor U14444 (N_14444,N_9689,N_9871);
nor U14445 (N_14445,N_5697,N_7520);
nand U14446 (N_14446,N_6477,N_5576);
and U14447 (N_14447,N_7114,N_5116);
nand U14448 (N_14448,N_5309,N_5877);
or U14449 (N_14449,N_8710,N_7636);
nor U14450 (N_14450,N_7387,N_9094);
or U14451 (N_14451,N_7737,N_7891);
and U14452 (N_14452,N_6436,N_7511);
nor U14453 (N_14453,N_9981,N_6085);
and U14454 (N_14454,N_7905,N_7840);
nand U14455 (N_14455,N_9897,N_6280);
and U14456 (N_14456,N_9525,N_8253);
and U14457 (N_14457,N_6914,N_7592);
nor U14458 (N_14458,N_5389,N_6438);
or U14459 (N_14459,N_7574,N_5988);
nand U14460 (N_14460,N_7143,N_8591);
or U14461 (N_14461,N_5807,N_9471);
and U14462 (N_14462,N_6976,N_6802);
or U14463 (N_14463,N_7081,N_9522);
or U14464 (N_14464,N_8289,N_8286);
xnor U14465 (N_14465,N_9006,N_6547);
or U14466 (N_14466,N_6255,N_9245);
nor U14467 (N_14467,N_6157,N_9492);
or U14468 (N_14468,N_5231,N_5957);
or U14469 (N_14469,N_8956,N_9967);
or U14470 (N_14470,N_8135,N_8693);
nor U14471 (N_14471,N_7070,N_6112);
or U14472 (N_14472,N_9603,N_5131);
nor U14473 (N_14473,N_9563,N_7247);
nand U14474 (N_14474,N_9163,N_9458);
nand U14475 (N_14475,N_8354,N_7393);
or U14476 (N_14476,N_6247,N_6202);
nand U14477 (N_14477,N_5074,N_8133);
nand U14478 (N_14478,N_8388,N_5422);
or U14479 (N_14479,N_8447,N_7755);
nor U14480 (N_14480,N_9063,N_6926);
and U14481 (N_14481,N_5350,N_8548);
nor U14482 (N_14482,N_6382,N_5455);
nor U14483 (N_14483,N_8853,N_6735);
nor U14484 (N_14484,N_7334,N_5485);
or U14485 (N_14485,N_9045,N_9462);
nand U14486 (N_14486,N_5864,N_6011);
and U14487 (N_14487,N_8304,N_8003);
nand U14488 (N_14488,N_5848,N_8467);
nor U14489 (N_14489,N_8983,N_7624);
or U14490 (N_14490,N_6226,N_6827);
nand U14491 (N_14491,N_7960,N_7214);
or U14492 (N_14492,N_8699,N_6596);
or U14493 (N_14493,N_6782,N_8492);
nor U14494 (N_14494,N_9736,N_9306);
nor U14495 (N_14495,N_5809,N_8164);
or U14496 (N_14496,N_6961,N_6088);
nand U14497 (N_14497,N_8113,N_7875);
and U14498 (N_14498,N_6284,N_9077);
and U14499 (N_14499,N_6342,N_8793);
or U14500 (N_14500,N_5222,N_5292);
or U14501 (N_14501,N_6376,N_9715);
or U14502 (N_14502,N_5018,N_9500);
and U14503 (N_14503,N_9346,N_9911);
nand U14504 (N_14504,N_6610,N_9455);
nand U14505 (N_14505,N_6587,N_6214);
nand U14506 (N_14506,N_6535,N_8888);
nor U14507 (N_14507,N_5765,N_8538);
and U14508 (N_14508,N_8939,N_5700);
nand U14509 (N_14509,N_8701,N_7614);
and U14510 (N_14510,N_8656,N_8764);
or U14511 (N_14511,N_7078,N_6674);
nor U14512 (N_14512,N_6168,N_5217);
nor U14513 (N_14513,N_8999,N_8193);
nand U14514 (N_14514,N_8687,N_9816);
nor U14515 (N_14515,N_8369,N_6296);
nor U14516 (N_14516,N_7107,N_6817);
nand U14517 (N_14517,N_7330,N_5136);
nor U14518 (N_14518,N_6162,N_8964);
nor U14519 (N_14519,N_7279,N_8085);
and U14520 (N_14520,N_5229,N_9403);
or U14521 (N_14521,N_8120,N_8969);
and U14522 (N_14522,N_6063,N_5149);
nor U14523 (N_14523,N_9330,N_9827);
nand U14524 (N_14524,N_5414,N_5622);
or U14525 (N_14525,N_5365,N_8547);
or U14526 (N_14526,N_9460,N_7316);
xor U14527 (N_14527,N_9287,N_8051);
nand U14528 (N_14528,N_7866,N_6448);
nand U14529 (N_14529,N_9025,N_9674);
nand U14530 (N_14530,N_8808,N_9507);
nand U14531 (N_14531,N_5669,N_7341);
and U14532 (N_14532,N_5727,N_7995);
and U14533 (N_14533,N_8170,N_7236);
and U14534 (N_14534,N_9895,N_8886);
nand U14535 (N_14535,N_8259,N_6198);
and U14536 (N_14536,N_8732,N_5054);
nand U14537 (N_14537,N_9922,N_9258);
nor U14538 (N_14538,N_8314,N_6485);
and U14539 (N_14539,N_5528,N_7307);
or U14540 (N_14540,N_7045,N_8188);
or U14541 (N_14541,N_9309,N_7409);
and U14542 (N_14542,N_6397,N_5613);
or U14543 (N_14543,N_9920,N_9428);
nor U14544 (N_14544,N_8058,N_7666);
and U14545 (N_14545,N_5324,N_8939);
and U14546 (N_14546,N_6711,N_8068);
and U14547 (N_14547,N_9726,N_9207);
and U14548 (N_14548,N_8160,N_9774);
and U14549 (N_14549,N_6096,N_7825);
xor U14550 (N_14550,N_8443,N_9853);
and U14551 (N_14551,N_7855,N_6902);
nor U14552 (N_14552,N_8909,N_8776);
nor U14553 (N_14553,N_5340,N_9637);
nand U14554 (N_14554,N_5021,N_9871);
nor U14555 (N_14555,N_5732,N_6689);
nand U14556 (N_14556,N_6317,N_7333);
and U14557 (N_14557,N_5971,N_9677);
or U14558 (N_14558,N_5344,N_9156);
nand U14559 (N_14559,N_9037,N_5214);
or U14560 (N_14560,N_6087,N_8678);
and U14561 (N_14561,N_9171,N_5605);
and U14562 (N_14562,N_8423,N_6362);
and U14563 (N_14563,N_9416,N_9873);
nand U14564 (N_14564,N_6950,N_9994);
nor U14565 (N_14565,N_8649,N_6880);
or U14566 (N_14566,N_6647,N_9400);
or U14567 (N_14567,N_5701,N_8902);
nor U14568 (N_14568,N_7563,N_6889);
and U14569 (N_14569,N_6986,N_8932);
and U14570 (N_14570,N_9566,N_7575);
nor U14571 (N_14571,N_5296,N_6763);
xor U14572 (N_14572,N_5501,N_8575);
nor U14573 (N_14573,N_9805,N_8640);
nor U14574 (N_14574,N_9901,N_5928);
nand U14575 (N_14575,N_8868,N_8719);
and U14576 (N_14576,N_8364,N_5888);
and U14577 (N_14577,N_6872,N_5002);
or U14578 (N_14578,N_8079,N_5754);
nand U14579 (N_14579,N_9550,N_7704);
or U14580 (N_14580,N_8923,N_7304);
nand U14581 (N_14581,N_7508,N_6532);
nor U14582 (N_14582,N_6876,N_9919);
nand U14583 (N_14583,N_6438,N_8720);
or U14584 (N_14584,N_7751,N_8640);
and U14585 (N_14585,N_7015,N_6166);
or U14586 (N_14586,N_8935,N_5891);
nor U14587 (N_14587,N_5701,N_7449);
or U14588 (N_14588,N_5583,N_8100);
nand U14589 (N_14589,N_7567,N_9766);
nor U14590 (N_14590,N_6212,N_5613);
or U14591 (N_14591,N_9667,N_7006);
and U14592 (N_14592,N_7572,N_6268);
and U14593 (N_14593,N_9638,N_8865);
nor U14594 (N_14594,N_7065,N_6654);
nand U14595 (N_14595,N_7988,N_9658);
and U14596 (N_14596,N_6279,N_7786);
nand U14597 (N_14597,N_7970,N_9920);
or U14598 (N_14598,N_5089,N_8934);
nor U14599 (N_14599,N_7238,N_6360);
or U14600 (N_14600,N_6823,N_9534);
and U14601 (N_14601,N_6528,N_9048);
or U14602 (N_14602,N_6415,N_5770);
or U14603 (N_14603,N_7112,N_6652);
or U14604 (N_14604,N_5824,N_8980);
or U14605 (N_14605,N_7868,N_6793);
and U14606 (N_14606,N_6817,N_7526);
nand U14607 (N_14607,N_8829,N_9390);
nor U14608 (N_14608,N_8683,N_6324);
nor U14609 (N_14609,N_7864,N_5344);
nor U14610 (N_14610,N_5372,N_7387);
and U14611 (N_14611,N_7656,N_9431);
nand U14612 (N_14612,N_8615,N_8934);
or U14613 (N_14613,N_7248,N_8347);
or U14614 (N_14614,N_7134,N_7315);
nor U14615 (N_14615,N_7270,N_9096);
and U14616 (N_14616,N_5538,N_9797);
nor U14617 (N_14617,N_9809,N_6524);
nor U14618 (N_14618,N_8431,N_7763);
nor U14619 (N_14619,N_6938,N_8509);
or U14620 (N_14620,N_6590,N_8875);
nor U14621 (N_14621,N_5444,N_5993);
nor U14622 (N_14622,N_8189,N_8304);
and U14623 (N_14623,N_6517,N_8052);
and U14624 (N_14624,N_7005,N_9940);
nor U14625 (N_14625,N_8567,N_7502);
nand U14626 (N_14626,N_9915,N_8360);
nor U14627 (N_14627,N_6773,N_9503);
or U14628 (N_14628,N_8182,N_5371);
nor U14629 (N_14629,N_5999,N_9607);
and U14630 (N_14630,N_7488,N_9487);
nor U14631 (N_14631,N_5165,N_9341);
xor U14632 (N_14632,N_8288,N_8236);
and U14633 (N_14633,N_8776,N_8553);
nand U14634 (N_14634,N_6413,N_8656);
or U14635 (N_14635,N_9593,N_5231);
nand U14636 (N_14636,N_9592,N_6835);
nor U14637 (N_14637,N_8933,N_9438);
and U14638 (N_14638,N_9188,N_9807);
nor U14639 (N_14639,N_7295,N_6081);
nand U14640 (N_14640,N_6672,N_7518);
and U14641 (N_14641,N_9415,N_5801);
or U14642 (N_14642,N_6651,N_8252);
nand U14643 (N_14643,N_7033,N_5845);
nor U14644 (N_14644,N_9239,N_7494);
or U14645 (N_14645,N_7285,N_6456);
or U14646 (N_14646,N_7471,N_9554);
or U14647 (N_14647,N_5592,N_7049);
and U14648 (N_14648,N_9751,N_9503);
nand U14649 (N_14649,N_9951,N_7312);
nor U14650 (N_14650,N_6131,N_8412);
nor U14651 (N_14651,N_7546,N_9194);
nor U14652 (N_14652,N_5382,N_7592);
or U14653 (N_14653,N_5842,N_8429);
nand U14654 (N_14654,N_5764,N_7314);
nor U14655 (N_14655,N_5217,N_6047);
or U14656 (N_14656,N_5855,N_8787);
and U14657 (N_14657,N_8068,N_6663);
nor U14658 (N_14658,N_7719,N_7019);
and U14659 (N_14659,N_7555,N_7629);
nor U14660 (N_14660,N_6875,N_7632);
nand U14661 (N_14661,N_8713,N_8887);
or U14662 (N_14662,N_5960,N_6637);
or U14663 (N_14663,N_6389,N_6305);
nor U14664 (N_14664,N_7100,N_7964);
nand U14665 (N_14665,N_6963,N_5853);
or U14666 (N_14666,N_8624,N_6462);
nand U14667 (N_14667,N_5307,N_9213);
or U14668 (N_14668,N_6561,N_8756);
and U14669 (N_14669,N_6544,N_7967);
nand U14670 (N_14670,N_5636,N_8391);
and U14671 (N_14671,N_6822,N_8798);
nand U14672 (N_14672,N_6330,N_9712);
and U14673 (N_14673,N_7202,N_8754);
nand U14674 (N_14674,N_6898,N_5068);
nand U14675 (N_14675,N_7816,N_5260);
nand U14676 (N_14676,N_7385,N_7125);
nand U14677 (N_14677,N_5146,N_8424);
nand U14678 (N_14678,N_9590,N_6698);
nor U14679 (N_14679,N_5334,N_7114);
and U14680 (N_14680,N_6890,N_8142);
nand U14681 (N_14681,N_9405,N_6897);
nor U14682 (N_14682,N_9967,N_8388);
and U14683 (N_14683,N_6536,N_5965);
nor U14684 (N_14684,N_8236,N_7564);
nor U14685 (N_14685,N_9246,N_5802);
and U14686 (N_14686,N_9798,N_9218);
xor U14687 (N_14687,N_9111,N_9613);
nor U14688 (N_14688,N_5775,N_8487);
and U14689 (N_14689,N_9338,N_6066);
or U14690 (N_14690,N_5456,N_8027);
and U14691 (N_14691,N_7095,N_7285);
nand U14692 (N_14692,N_7134,N_5760);
and U14693 (N_14693,N_6902,N_6479);
nor U14694 (N_14694,N_5557,N_8857);
nand U14695 (N_14695,N_5356,N_8633);
nand U14696 (N_14696,N_8180,N_7160);
nand U14697 (N_14697,N_8543,N_5811);
and U14698 (N_14698,N_8964,N_9297);
or U14699 (N_14699,N_8263,N_7341);
and U14700 (N_14700,N_6087,N_9655);
nor U14701 (N_14701,N_8310,N_6004);
nand U14702 (N_14702,N_8133,N_8290);
nand U14703 (N_14703,N_9804,N_9655);
or U14704 (N_14704,N_7441,N_5792);
and U14705 (N_14705,N_5321,N_7210);
or U14706 (N_14706,N_5794,N_5303);
nand U14707 (N_14707,N_8351,N_9308);
and U14708 (N_14708,N_6244,N_9243);
nor U14709 (N_14709,N_5731,N_9240);
and U14710 (N_14710,N_8457,N_5582);
nor U14711 (N_14711,N_9298,N_5314);
nand U14712 (N_14712,N_6083,N_9465);
nor U14713 (N_14713,N_7382,N_9854);
nor U14714 (N_14714,N_6767,N_5712);
or U14715 (N_14715,N_8712,N_9788);
nor U14716 (N_14716,N_6938,N_7835);
or U14717 (N_14717,N_8529,N_8293);
nor U14718 (N_14718,N_6361,N_6625);
nand U14719 (N_14719,N_8303,N_6963);
or U14720 (N_14720,N_9786,N_8230);
nand U14721 (N_14721,N_8121,N_9929);
or U14722 (N_14722,N_7840,N_5269);
nand U14723 (N_14723,N_5528,N_7295);
and U14724 (N_14724,N_9306,N_7809);
or U14725 (N_14725,N_6092,N_5627);
or U14726 (N_14726,N_7292,N_7477);
and U14727 (N_14727,N_9335,N_9662);
and U14728 (N_14728,N_6349,N_6975);
and U14729 (N_14729,N_5323,N_9801);
and U14730 (N_14730,N_6236,N_5625);
nand U14731 (N_14731,N_5455,N_6232);
and U14732 (N_14732,N_6820,N_5821);
nand U14733 (N_14733,N_9678,N_8126);
and U14734 (N_14734,N_7728,N_5487);
nor U14735 (N_14735,N_8605,N_7299);
or U14736 (N_14736,N_5832,N_8103);
and U14737 (N_14737,N_5624,N_9041);
or U14738 (N_14738,N_6634,N_8395);
nor U14739 (N_14739,N_9370,N_6871);
nand U14740 (N_14740,N_9140,N_8453);
or U14741 (N_14741,N_5861,N_8214);
or U14742 (N_14742,N_6763,N_9609);
nor U14743 (N_14743,N_9429,N_7122);
and U14744 (N_14744,N_7249,N_7161);
nand U14745 (N_14745,N_9074,N_7512);
nand U14746 (N_14746,N_8496,N_9648);
nor U14747 (N_14747,N_8540,N_7983);
and U14748 (N_14748,N_5647,N_7251);
nor U14749 (N_14749,N_7078,N_9610);
xnor U14750 (N_14750,N_7403,N_9933);
nor U14751 (N_14751,N_9259,N_9678);
or U14752 (N_14752,N_5844,N_9849);
or U14753 (N_14753,N_6814,N_9671);
or U14754 (N_14754,N_5560,N_8242);
or U14755 (N_14755,N_8636,N_6414);
nand U14756 (N_14756,N_9962,N_6363);
xor U14757 (N_14757,N_6067,N_7935);
and U14758 (N_14758,N_8393,N_5573);
or U14759 (N_14759,N_8002,N_9906);
nor U14760 (N_14760,N_6687,N_9071);
and U14761 (N_14761,N_8077,N_6520);
and U14762 (N_14762,N_7819,N_5579);
and U14763 (N_14763,N_7879,N_6493);
or U14764 (N_14764,N_7238,N_6902);
and U14765 (N_14765,N_5667,N_9955);
and U14766 (N_14766,N_7623,N_5236);
and U14767 (N_14767,N_8355,N_5916);
nor U14768 (N_14768,N_5651,N_7429);
or U14769 (N_14769,N_8815,N_6890);
nand U14770 (N_14770,N_5323,N_6731);
nor U14771 (N_14771,N_5756,N_5641);
and U14772 (N_14772,N_9312,N_5243);
and U14773 (N_14773,N_6925,N_9511);
nand U14774 (N_14774,N_5421,N_8600);
nand U14775 (N_14775,N_6814,N_7834);
nand U14776 (N_14776,N_5072,N_8373);
nor U14777 (N_14777,N_7180,N_9387);
and U14778 (N_14778,N_8685,N_7462);
and U14779 (N_14779,N_5917,N_5477);
nor U14780 (N_14780,N_5105,N_7606);
and U14781 (N_14781,N_8122,N_5125);
nor U14782 (N_14782,N_6171,N_9911);
nor U14783 (N_14783,N_6917,N_5647);
nand U14784 (N_14784,N_9360,N_5815);
nor U14785 (N_14785,N_8848,N_7416);
and U14786 (N_14786,N_5919,N_7633);
or U14787 (N_14787,N_9088,N_5317);
and U14788 (N_14788,N_8348,N_5450);
nand U14789 (N_14789,N_6451,N_7326);
and U14790 (N_14790,N_7716,N_5528);
nor U14791 (N_14791,N_6097,N_6770);
nand U14792 (N_14792,N_9654,N_6417);
nor U14793 (N_14793,N_6164,N_9709);
nor U14794 (N_14794,N_7190,N_9603);
nor U14795 (N_14795,N_5502,N_7268);
nor U14796 (N_14796,N_9356,N_8786);
or U14797 (N_14797,N_6721,N_8988);
and U14798 (N_14798,N_7337,N_7825);
or U14799 (N_14799,N_5997,N_6466);
nand U14800 (N_14800,N_7071,N_6666);
nor U14801 (N_14801,N_6498,N_8769);
and U14802 (N_14802,N_5540,N_8492);
or U14803 (N_14803,N_9587,N_8273);
and U14804 (N_14804,N_5433,N_5802);
nand U14805 (N_14805,N_8527,N_7116);
or U14806 (N_14806,N_9603,N_8827);
or U14807 (N_14807,N_5141,N_7513);
nand U14808 (N_14808,N_8713,N_8957);
nand U14809 (N_14809,N_6815,N_9475);
or U14810 (N_14810,N_9725,N_6680);
or U14811 (N_14811,N_7564,N_5108);
and U14812 (N_14812,N_8100,N_9241);
nor U14813 (N_14813,N_7861,N_9340);
nor U14814 (N_14814,N_8625,N_6554);
or U14815 (N_14815,N_7883,N_5494);
or U14816 (N_14816,N_9210,N_5244);
nor U14817 (N_14817,N_6280,N_7368);
or U14818 (N_14818,N_9526,N_9396);
and U14819 (N_14819,N_9900,N_8586);
nand U14820 (N_14820,N_9210,N_9248);
nor U14821 (N_14821,N_9252,N_8035);
nor U14822 (N_14822,N_6067,N_9401);
and U14823 (N_14823,N_5746,N_8048);
nand U14824 (N_14824,N_8214,N_6411);
nor U14825 (N_14825,N_8644,N_6205);
and U14826 (N_14826,N_6305,N_5297);
and U14827 (N_14827,N_6105,N_7801);
nand U14828 (N_14828,N_6979,N_5334);
nor U14829 (N_14829,N_5420,N_8534);
or U14830 (N_14830,N_6683,N_7473);
nand U14831 (N_14831,N_6347,N_9672);
or U14832 (N_14832,N_7134,N_5624);
nand U14833 (N_14833,N_7486,N_6267);
nand U14834 (N_14834,N_6947,N_7530);
and U14835 (N_14835,N_8482,N_6039);
or U14836 (N_14836,N_6273,N_5754);
nand U14837 (N_14837,N_8219,N_9935);
or U14838 (N_14838,N_7767,N_6873);
nand U14839 (N_14839,N_6543,N_5875);
or U14840 (N_14840,N_6506,N_5625);
nand U14841 (N_14841,N_6296,N_8984);
and U14842 (N_14842,N_8601,N_7645);
nor U14843 (N_14843,N_9869,N_9936);
and U14844 (N_14844,N_9846,N_7828);
nand U14845 (N_14845,N_8062,N_7733);
and U14846 (N_14846,N_8489,N_8628);
nor U14847 (N_14847,N_9552,N_8649);
or U14848 (N_14848,N_6702,N_8209);
or U14849 (N_14849,N_5704,N_6248);
nor U14850 (N_14850,N_7425,N_6821);
or U14851 (N_14851,N_6649,N_9020);
nor U14852 (N_14852,N_7521,N_8468);
or U14853 (N_14853,N_9447,N_9177);
nand U14854 (N_14854,N_7225,N_8846);
nor U14855 (N_14855,N_8795,N_6430);
nor U14856 (N_14856,N_6538,N_9259);
nor U14857 (N_14857,N_9225,N_7328);
nor U14858 (N_14858,N_7523,N_9840);
or U14859 (N_14859,N_7656,N_8719);
and U14860 (N_14860,N_9638,N_8316);
nor U14861 (N_14861,N_6289,N_6176);
and U14862 (N_14862,N_9058,N_5222);
nor U14863 (N_14863,N_7825,N_5666);
nand U14864 (N_14864,N_7974,N_9458);
or U14865 (N_14865,N_8707,N_6750);
nor U14866 (N_14866,N_6573,N_6484);
and U14867 (N_14867,N_5623,N_7594);
or U14868 (N_14868,N_5987,N_6854);
or U14869 (N_14869,N_9105,N_8600);
or U14870 (N_14870,N_7986,N_9479);
or U14871 (N_14871,N_8547,N_9724);
nand U14872 (N_14872,N_8698,N_5586);
nor U14873 (N_14873,N_5297,N_8738);
nand U14874 (N_14874,N_9214,N_5341);
or U14875 (N_14875,N_9941,N_5086);
nor U14876 (N_14876,N_9839,N_8818);
nand U14877 (N_14877,N_7021,N_6869);
and U14878 (N_14878,N_9039,N_5389);
or U14879 (N_14879,N_9914,N_5369);
nor U14880 (N_14880,N_9984,N_9923);
nand U14881 (N_14881,N_7260,N_7606);
nor U14882 (N_14882,N_7125,N_5751);
nor U14883 (N_14883,N_8139,N_9263);
or U14884 (N_14884,N_8877,N_5484);
nor U14885 (N_14885,N_8978,N_9680);
nor U14886 (N_14886,N_7545,N_9111);
and U14887 (N_14887,N_6372,N_5545);
nand U14888 (N_14888,N_8661,N_9311);
xor U14889 (N_14889,N_7697,N_9485);
nor U14890 (N_14890,N_7061,N_7092);
or U14891 (N_14891,N_6108,N_5898);
nor U14892 (N_14892,N_9561,N_6630);
and U14893 (N_14893,N_6086,N_5457);
or U14894 (N_14894,N_7469,N_6979);
or U14895 (N_14895,N_8281,N_8444);
and U14896 (N_14896,N_7292,N_9342);
and U14897 (N_14897,N_5365,N_7850);
nor U14898 (N_14898,N_9399,N_5182);
and U14899 (N_14899,N_9653,N_8888);
nand U14900 (N_14900,N_8969,N_7156);
or U14901 (N_14901,N_9487,N_6990);
and U14902 (N_14902,N_5808,N_8772);
or U14903 (N_14903,N_7534,N_8326);
nor U14904 (N_14904,N_7954,N_9437);
nand U14905 (N_14905,N_8430,N_7589);
nand U14906 (N_14906,N_7185,N_5648);
and U14907 (N_14907,N_9297,N_9106);
and U14908 (N_14908,N_5940,N_9385);
nand U14909 (N_14909,N_7807,N_8858);
nand U14910 (N_14910,N_7657,N_6120);
nand U14911 (N_14911,N_7200,N_7457);
or U14912 (N_14912,N_9414,N_6497);
nand U14913 (N_14913,N_6190,N_5424);
and U14914 (N_14914,N_8277,N_7211);
nand U14915 (N_14915,N_7924,N_8448);
or U14916 (N_14916,N_8375,N_8500);
and U14917 (N_14917,N_6054,N_7188);
or U14918 (N_14918,N_9977,N_6983);
or U14919 (N_14919,N_8616,N_9978);
nand U14920 (N_14920,N_7533,N_8679);
and U14921 (N_14921,N_8834,N_7406);
and U14922 (N_14922,N_5634,N_5525);
xor U14923 (N_14923,N_5599,N_7742);
nand U14924 (N_14924,N_6645,N_5855);
nand U14925 (N_14925,N_7019,N_8179);
and U14926 (N_14926,N_9075,N_8601);
nor U14927 (N_14927,N_5541,N_9426);
or U14928 (N_14928,N_7066,N_7346);
and U14929 (N_14929,N_5583,N_7829);
nor U14930 (N_14930,N_8578,N_9198);
or U14931 (N_14931,N_9782,N_6931);
and U14932 (N_14932,N_7115,N_8003);
nor U14933 (N_14933,N_6906,N_5617);
nand U14934 (N_14934,N_7802,N_8913);
nand U14935 (N_14935,N_7575,N_5618);
and U14936 (N_14936,N_8966,N_6301);
or U14937 (N_14937,N_8523,N_6571);
or U14938 (N_14938,N_8385,N_8321);
or U14939 (N_14939,N_5574,N_9679);
nor U14940 (N_14940,N_5195,N_5201);
and U14941 (N_14941,N_5220,N_5868);
and U14942 (N_14942,N_9362,N_5873);
and U14943 (N_14943,N_5503,N_7709);
nor U14944 (N_14944,N_5471,N_5198);
or U14945 (N_14945,N_6030,N_5370);
nor U14946 (N_14946,N_6283,N_9406);
or U14947 (N_14947,N_7913,N_8776);
or U14948 (N_14948,N_7124,N_7226);
nor U14949 (N_14949,N_8646,N_9482);
nor U14950 (N_14950,N_8781,N_7049);
or U14951 (N_14951,N_8088,N_7066);
nand U14952 (N_14952,N_9799,N_8016);
nand U14953 (N_14953,N_9988,N_9073);
nor U14954 (N_14954,N_9326,N_5410);
nand U14955 (N_14955,N_9527,N_8153);
and U14956 (N_14956,N_9962,N_5287);
nand U14957 (N_14957,N_6517,N_6142);
nand U14958 (N_14958,N_8767,N_6658);
nand U14959 (N_14959,N_5920,N_9336);
nand U14960 (N_14960,N_5100,N_6315);
nor U14961 (N_14961,N_7885,N_8687);
or U14962 (N_14962,N_9974,N_9228);
or U14963 (N_14963,N_5889,N_8612);
or U14964 (N_14964,N_8030,N_6113);
and U14965 (N_14965,N_5603,N_9705);
or U14966 (N_14966,N_9543,N_8000);
and U14967 (N_14967,N_6654,N_9427);
nor U14968 (N_14968,N_9661,N_7067);
and U14969 (N_14969,N_7408,N_7836);
or U14970 (N_14970,N_8212,N_6641);
and U14971 (N_14971,N_8911,N_5044);
or U14972 (N_14972,N_8264,N_9366);
or U14973 (N_14973,N_5638,N_7658);
or U14974 (N_14974,N_6254,N_6239);
nor U14975 (N_14975,N_6754,N_7714);
nand U14976 (N_14976,N_7181,N_6909);
nor U14977 (N_14977,N_7356,N_5103);
or U14978 (N_14978,N_5403,N_9273);
nand U14979 (N_14979,N_9811,N_8991);
or U14980 (N_14980,N_8571,N_9590);
or U14981 (N_14981,N_5887,N_9698);
nand U14982 (N_14982,N_5552,N_6438);
nand U14983 (N_14983,N_5410,N_6734);
nand U14984 (N_14984,N_6294,N_9359);
nor U14985 (N_14985,N_6711,N_6462);
or U14986 (N_14986,N_5435,N_5347);
or U14987 (N_14987,N_6589,N_9880);
and U14988 (N_14988,N_9293,N_8741);
nor U14989 (N_14989,N_9265,N_7828);
nand U14990 (N_14990,N_8744,N_5520);
or U14991 (N_14991,N_8768,N_6761);
or U14992 (N_14992,N_8080,N_6122);
nand U14993 (N_14993,N_8824,N_6666);
nand U14994 (N_14994,N_5433,N_5805);
or U14995 (N_14995,N_6562,N_6794);
nor U14996 (N_14996,N_5923,N_6642);
or U14997 (N_14997,N_9899,N_5343);
nand U14998 (N_14998,N_6983,N_5970);
or U14999 (N_14999,N_5102,N_6313);
nand U15000 (N_15000,N_13635,N_12819);
and U15001 (N_15001,N_13419,N_11498);
xor U15002 (N_15002,N_10408,N_10520);
and U15003 (N_15003,N_12793,N_11025);
and U15004 (N_15004,N_10400,N_12883);
or U15005 (N_15005,N_14563,N_12243);
and U15006 (N_15006,N_11570,N_13256);
and U15007 (N_15007,N_11728,N_13325);
nor U15008 (N_15008,N_14099,N_13455);
and U15009 (N_15009,N_12119,N_11780);
or U15010 (N_15010,N_10468,N_12513);
and U15011 (N_15011,N_14538,N_11963);
nand U15012 (N_15012,N_13890,N_11612);
nor U15013 (N_15013,N_12671,N_11341);
and U15014 (N_15014,N_10279,N_11052);
and U15015 (N_15015,N_13286,N_11461);
nand U15016 (N_15016,N_14978,N_11924);
and U15017 (N_15017,N_14699,N_13672);
and U15018 (N_15018,N_10594,N_14742);
or U15019 (N_15019,N_12955,N_13856);
or U15020 (N_15020,N_13211,N_10623);
xor U15021 (N_15021,N_12845,N_10919);
nor U15022 (N_15022,N_11663,N_10569);
nand U15023 (N_15023,N_12804,N_10316);
nor U15024 (N_15024,N_13513,N_13497);
and U15025 (N_15025,N_14012,N_14565);
nor U15026 (N_15026,N_12407,N_13449);
nand U15027 (N_15027,N_11426,N_14349);
and U15028 (N_15028,N_14910,N_11578);
nand U15029 (N_15029,N_11708,N_14104);
and U15030 (N_15030,N_11907,N_12928);
nand U15031 (N_15031,N_10150,N_13245);
nor U15032 (N_15032,N_10430,N_10626);
and U15033 (N_15033,N_11109,N_10972);
nand U15034 (N_15034,N_13451,N_13422);
and U15035 (N_15035,N_12189,N_13039);
or U15036 (N_15036,N_10374,N_11378);
or U15037 (N_15037,N_11914,N_13399);
nand U15038 (N_15038,N_14945,N_14931);
and U15039 (N_15039,N_10806,N_12163);
nor U15040 (N_15040,N_13876,N_13309);
nor U15041 (N_15041,N_11683,N_11597);
nor U15042 (N_15042,N_10779,N_12875);
nor U15043 (N_15043,N_11418,N_13779);
nor U15044 (N_15044,N_10656,N_10578);
or U15045 (N_15045,N_14835,N_10431);
or U15046 (N_15046,N_14250,N_11503);
and U15047 (N_15047,N_11806,N_13444);
nand U15048 (N_15048,N_13116,N_14124);
and U15049 (N_15049,N_13602,N_11958);
nor U15050 (N_15050,N_13210,N_12543);
and U15051 (N_15051,N_13804,N_14050);
nand U15052 (N_15052,N_10717,N_10151);
or U15053 (N_15053,N_12584,N_11697);
nand U15054 (N_15054,N_10356,N_11591);
or U15055 (N_15055,N_12601,N_13137);
or U15056 (N_15056,N_14290,N_14069);
and U15057 (N_15057,N_14571,N_11118);
and U15058 (N_15058,N_13695,N_12923);
nand U15059 (N_15059,N_10928,N_12102);
or U15060 (N_15060,N_12185,N_13459);
and U15061 (N_15061,N_13749,N_13769);
and U15062 (N_15062,N_12772,N_10551);
nand U15063 (N_15063,N_13660,N_11156);
xor U15064 (N_15064,N_13202,N_14287);
and U15065 (N_15065,N_11234,N_12290);
nor U15066 (N_15066,N_12881,N_12559);
or U15067 (N_15067,N_13611,N_11759);
and U15068 (N_15068,N_13648,N_12794);
or U15069 (N_15069,N_13280,N_14786);
or U15070 (N_15070,N_12729,N_12609);
nor U15071 (N_15071,N_11363,N_14583);
or U15072 (N_15072,N_14119,N_13281);
nor U15073 (N_15073,N_11230,N_12203);
or U15074 (N_15074,N_14589,N_12944);
and U15075 (N_15075,N_10525,N_12703);
or U15076 (N_15076,N_13029,N_14371);
nand U15077 (N_15077,N_11559,N_14464);
and U15078 (N_15078,N_14638,N_14698);
nand U15079 (N_15079,N_13035,N_13884);
or U15080 (N_15080,N_12504,N_12977);
nand U15081 (N_15081,N_12791,N_14007);
and U15082 (N_15082,N_13500,N_14856);
xnor U15083 (N_15083,N_11615,N_11482);
nor U15084 (N_15084,N_11389,N_13011);
and U15085 (N_15085,N_10305,N_11198);
and U15086 (N_15086,N_11420,N_14015);
or U15087 (N_15087,N_11167,N_11055);
nand U15088 (N_15088,N_14787,N_10961);
and U15089 (N_15089,N_10250,N_13369);
nand U15090 (N_15090,N_11676,N_14550);
or U15091 (N_15091,N_11154,N_14803);
nor U15092 (N_15092,N_14614,N_12635);
or U15093 (N_15093,N_10591,N_11732);
and U15094 (N_15094,N_13199,N_11462);
nand U15095 (N_15095,N_14259,N_10503);
and U15096 (N_15096,N_10954,N_14804);
nor U15097 (N_15097,N_13299,N_11117);
or U15098 (N_15098,N_13244,N_11931);
nand U15099 (N_15099,N_13456,N_10653);
or U15100 (N_15100,N_14768,N_11529);
nor U15101 (N_15101,N_10963,N_12694);
or U15102 (N_15102,N_11543,N_10969);
and U15103 (N_15103,N_10882,N_12331);
and U15104 (N_15104,N_10071,N_12452);
nand U15105 (N_15105,N_11816,N_11011);
nor U15106 (N_15106,N_13662,N_13151);
or U15107 (N_15107,N_12877,N_11454);
or U15108 (N_15108,N_10583,N_11565);
or U15109 (N_15109,N_11768,N_11553);
or U15110 (N_15110,N_12376,N_10877);
nand U15111 (N_15111,N_13208,N_12567);
or U15112 (N_15112,N_14416,N_11065);
nand U15113 (N_15113,N_14096,N_10489);
and U15114 (N_15114,N_14561,N_13697);
nor U15115 (N_15115,N_10289,N_14721);
nor U15116 (N_15116,N_12956,N_13327);
xnor U15117 (N_15117,N_10548,N_14204);
nand U15118 (N_15118,N_10792,N_12117);
nand U15119 (N_15119,N_10115,N_13903);
and U15120 (N_15120,N_14067,N_13331);
or U15121 (N_15121,N_11743,N_11797);
or U15122 (N_15122,N_10690,N_13366);
or U15123 (N_15123,N_10738,N_14309);
nor U15124 (N_15124,N_11374,N_13512);
or U15125 (N_15125,N_12523,N_14516);
nor U15126 (N_15126,N_10276,N_13825);
or U15127 (N_15127,N_12488,N_12850);
or U15128 (N_15128,N_13814,N_11416);
nor U15129 (N_15129,N_14273,N_11369);
nand U15130 (N_15130,N_14210,N_12186);
or U15131 (N_15131,N_11210,N_10642);
or U15132 (N_15132,N_12045,N_13507);
or U15133 (N_15133,N_12582,N_10444);
and U15134 (N_15134,N_13488,N_14381);
and U15135 (N_15135,N_10308,N_10080);
nand U15136 (N_15136,N_12428,N_11532);
nor U15137 (N_15137,N_11906,N_12071);
xnor U15138 (N_15138,N_11904,N_10934);
and U15139 (N_15139,N_13720,N_11355);
or U15140 (N_15140,N_10202,N_12183);
or U15141 (N_15141,N_13810,N_13114);
and U15142 (N_15142,N_12140,N_12372);
or U15143 (N_15143,N_14556,N_12404);
or U15144 (N_15144,N_13462,N_13384);
nand U15145 (N_15145,N_13382,N_12992);
and U15146 (N_15146,N_14375,N_12561);
and U15147 (N_15147,N_14534,N_13683);
nand U15148 (N_15148,N_13617,N_13129);
and U15149 (N_15149,N_11609,N_14954);
and U15150 (N_15150,N_11839,N_13473);
nor U15151 (N_15151,N_14449,N_10439);
nand U15152 (N_15152,N_12661,N_14755);
nor U15153 (N_15153,N_13751,N_14611);
nor U15154 (N_15154,N_10980,N_10370);
and U15155 (N_15155,N_10424,N_12359);
nand U15156 (N_15156,N_14396,N_10948);
nor U15157 (N_15157,N_11444,N_11224);
and U15158 (N_15158,N_11225,N_14531);
nor U15159 (N_15159,N_11879,N_11766);
or U15160 (N_15160,N_14327,N_14485);
and U15161 (N_15161,N_12829,N_13427);
nor U15162 (N_15162,N_14566,N_13942);
nor U15163 (N_15163,N_13113,N_14609);
nor U15164 (N_15164,N_10286,N_14604);
or U15165 (N_15165,N_10796,N_10691);
or U15166 (N_15166,N_11004,N_13480);
or U15167 (N_15167,N_13490,N_13122);
and U15168 (N_15168,N_13900,N_12238);
nand U15169 (N_15169,N_14590,N_13030);
and U15170 (N_15170,N_10372,N_13347);
nor U15171 (N_15171,N_11739,N_13886);
nor U15172 (N_15172,N_10793,N_10709);
or U15173 (N_15173,N_13951,N_10159);
and U15174 (N_15174,N_12677,N_14622);
nor U15175 (N_15175,N_11966,N_12126);
xor U15176 (N_15176,N_10231,N_11077);
or U15177 (N_15177,N_10678,N_11116);
xor U15178 (N_15178,N_14491,N_14877);
nor U15179 (N_15179,N_12557,N_10572);
or U15180 (N_15180,N_12726,N_14808);
and U15181 (N_15181,N_11339,N_12371);
nor U15182 (N_15182,N_10098,N_13548);
nor U15183 (N_15183,N_12612,N_14781);
or U15184 (N_15184,N_10956,N_14388);
or U15185 (N_15185,N_13529,N_10933);
or U15186 (N_15186,N_13196,N_13532);
and U15187 (N_15187,N_11460,N_11448);
nand U15188 (N_15188,N_13094,N_14626);
or U15189 (N_15189,N_14010,N_11294);
or U15190 (N_15190,N_12349,N_13776);
nor U15191 (N_15191,N_10593,N_13669);
or U15192 (N_15192,N_13706,N_14438);
nand U15193 (N_15193,N_14551,N_14526);
nand U15194 (N_15194,N_12985,N_13790);
nand U15195 (N_15195,N_11384,N_14648);
nor U15196 (N_15196,N_14624,N_12942);
nor U15197 (N_15197,N_13395,N_12960);
nand U15198 (N_15198,N_11603,N_12303);
xnor U15199 (N_15199,N_13883,N_10506);
nor U15200 (N_15200,N_11084,N_12013);
and U15201 (N_15201,N_14173,N_13381);
nor U15202 (N_15202,N_11740,N_10351);
or U15203 (N_15203,N_12971,N_13324);
and U15204 (N_15204,N_12408,N_14656);
and U15205 (N_15205,N_14822,N_12733);
nand U15206 (N_15206,N_14736,N_10407);
and U15207 (N_15207,N_14380,N_12354);
or U15208 (N_15208,N_13530,N_14577);
and U15209 (N_15209,N_13736,N_10258);
nand U15210 (N_15210,N_13821,N_11172);
nor U15211 (N_15211,N_11887,N_14362);
and U15212 (N_15212,N_13008,N_14540);
and U15213 (N_15213,N_10251,N_12654);
nor U15214 (N_15214,N_13575,N_12553);
and U15215 (N_15215,N_12360,N_12921);
nor U15216 (N_15216,N_11539,N_10784);
nor U15217 (N_15217,N_13267,N_11223);
and U15218 (N_15218,N_12920,N_12207);
nand U15219 (N_15219,N_10838,N_13235);
or U15220 (N_15220,N_12054,N_12946);
or U15221 (N_15221,N_14206,N_12652);
nand U15222 (N_15222,N_10574,N_14965);
or U15223 (N_15223,N_10339,N_11174);
or U15224 (N_15224,N_14299,N_12687);
nor U15225 (N_15225,N_14576,N_12846);
nor U15226 (N_15226,N_12155,N_11368);
and U15227 (N_15227,N_11397,N_10026);
nor U15228 (N_15228,N_13555,N_14831);
and U15229 (N_15229,N_14586,N_12897);
nand U15230 (N_15230,N_11562,N_10900);
and U15231 (N_15231,N_12742,N_11506);
nor U15232 (N_15232,N_14970,N_13981);
or U15233 (N_15233,N_11695,N_14653);
nor U15234 (N_15234,N_12369,N_12773);
nor U15235 (N_15235,N_14915,N_14415);
nand U15236 (N_15236,N_12051,N_10474);
nor U15237 (N_15237,N_13364,N_13626);
and U15238 (N_15238,N_14291,N_13774);
and U15239 (N_15239,N_10324,N_12175);
and U15240 (N_15240,N_13588,N_14373);
nor U15241 (N_15241,N_10477,N_13693);
nor U15242 (N_15242,N_11934,N_14497);
nor U15243 (N_15243,N_14649,N_10420);
nand U15244 (N_15244,N_10299,N_13881);
and U15245 (N_15245,N_11098,N_11616);
nor U15246 (N_15246,N_10955,N_12965);
nor U15247 (N_15247,N_10632,N_14058);
or U15248 (N_15248,N_12110,N_12728);
or U15249 (N_15249,N_11509,N_13013);
nand U15250 (N_15250,N_11193,N_14441);
nand U15251 (N_15251,N_12464,N_13054);
or U15252 (N_15252,N_10813,N_11551);
nand U15253 (N_15253,N_11295,N_10832);
nor U15254 (N_15254,N_12864,N_10057);
or U15255 (N_15255,N_13458,N_10880);
and U15256 (N_15256,N_14465,N_14588);
nor U15257 (N_15257,N_14002,N_10139);
nor U15258 (N_15258,N_10280,N_10571);
or U15259 (N_15259,N_10353,N_11813);
nand U15260 (N_15260,N_11108,N_14717);
nand U15261 (N_15261,N_10894,N_14353);
nor U15262 (N_15262,N_14255,N_11302);
or U15263 (N_15263,N_12415,N_12090);
nand U15264 (N_15264,N_13800,N_12673);
nor U15265 (N_15265,N_10913,N_13224);
nand U15266 (N_15266,N_13190,N_11082);
nand U15267 (N_15267,N_14592,N_13405);
nor U15268 (N_15268,N_11537,N_13780);
or U15269 (N_15269,N_13741,N_12005);
xnor U15270 (N_15270,N_13937,N_12658);
nor U15271 (N_15271,N_10826,N_13412);
and U15272 (N_15272,N_10570,N_14399);
nand U15273 (N_15273,N_12746,N_10889);
or U15274 (N_15274,N_10175,N_12160);
and U15275 (N_15275,N_11841,N_12329);
and U15276 (N_15276,N_10846,N_13646);
nand U15277 (N_15277,N_11112,N_10465);
or U15278 (N_15278,N_12637,N_13558);
and U15279 (N_15279,N_13365,N_10937);
or U15280 (N_15280,N_12707,N_14574);
nor U15281 (N_15281,N_12964,N_14405);
and U15282 (N_15282,N_12438,N_12824);
and U15283 (N_15283,N_10421,N_13147);
nor U15284 (N_15284,N_12681,N_13421);
nand U15285 (N_15285,N_10549,N_10247);
nand U15286 (N_15286,N_11528,N_11162);
and U15287 (N_15287,N_10695,N_13783);
nor U15288 (N_15288,N_12657,N_13023);
or U15289 (N_15289,N_14940,N_13359);
and U15290 (N_15290,N_11949,N_13615);
nor U15291 (N_15291,N_11171,N_13944);
nand U15292 (N_15292,N_13566,N_11214);
or U15293 (N_15293,N_11386,N_14557);
and U15294 (N_15294,N_14471,N_11820);
and U15295 (N_15295,N_11724,N_13545);
nor U15296 (N_15296,N_14138,N_14135);
and U15297 (N_15297,N_13371,N_12593);
nor U15298 (N_15298,N_10278,N_11794);
or U15299 (N_15299,N_10330,N_13229);
nor U15300 (N_15300,N_10189,N_11204);
nor U15301 (N_15301,N_10654,N_12665);
and U15302 (N_15302,N_12844,N_13465);
and U15303 (N_15303,N_10845,N_13144);
nand U15304 (N_15304,N_14231,N_14893);
nor U15305 (N_15305,N_13020,N_12491);
and U15306 (N_15306,N_13809,N_10769);
nand U15307 (N_15307,N_14844,N_12406);
or U15308 (N_15308,N_14128,N_10959);
nand U15309 (N_15309,N_12075,N_12104);
and U15310 (N_15310,N_10403,N_10469);
and U15311 (N_15311,N_13346,N_14018);
or U15312 (N_15312,N_13258,N_13428);
and U15313 (N_15313,N_11598,N_14579);
or U15314 (N_15314,N_14536,N_12865);
nor U15315 (N_15315,N_13358,N_13404);
and U15316 (N_15316,N_10261,N_11130);
and U15317 (N_15317,N_10780,N_13813);
nor U15318 (N_15318,N_10906,N_13453);
or U15319 (N_15319,N_12888,N_14172);
or U15320 (N_15320,N_14752,N_14003);
and U15321 (N_15321,N_12301,N_13043);
or U15322 (N_15322,N_10461,N_12487);
and U15323 (N_15323,N_12918,N_11308);
or U15324 (N_15324,N_11986,N_13521);
nand U15325 (N_15325,N_12385,N_14164);
and U15326 (N_15326,N_12237,N_13618);
nor U15327 (N_15327,N_11585,N_14317);
and U15328 (N_15328,N_10360,N_12061);
nor U15329 (N_15329,N_14771,N_12591);
nand U15330 (N_15330,N_12571,N_11495);
nand U15331 (N_15331,N_10563,N_14807);
nand U15332 (N_15332,N_12396,N_12202);
nor U15333 (N_15333,N_13477,N_11305);
nor U15334 (N_15334,N_10272,N_13895);
and U15335 (N_15335,N_13005,N_14553);
nand U15336 (N_15336,N_14004,N_11645);
nor U15337 (N_15337,N_11040,N_14275);
or U15338 (N_15338,N_10011,N_10984);
nand U15339 (N_15339,N_12906,N_13578);
and U15340 (N_15340,N_12993,N_14148);
or U15341 (N_15341,N_13954,N_13183);
nor U15342 (N_15342,N_12697,N_12927);
and U15343 (N_15343,N_10199,N_10336);
and U15344 (N_15344,N_11775,N_13910);
nor U15345 (N_15345,N_11189,N_13165);
and U15346 (N_15346,N_13389,N_13659);
and U15347 (N_15347,N_10789,N_12086);
nand U15348 (N_15348,N_11090,N_12527);
nor U15349 (N_15349,N_12326,N_11242);
and U15350 (N_15350,N_12530,N_10783);
and U15351 (N_15351,N_12919,N_14938);
nor U15352 (N_15352,N_10497,N_10655);
or U15353 (N_15353,N_11178,N_14113);
or U15354 (N_15354,N_12148,N_10652);
and U15355 (N_15355,N_10679,N_13928);
nand U15356 (N_15356,N_11252,N_11100);
and U15357 (N_15357,N_11930,N_14778);
nand U15358 (N_15358,N_11009,N_13785);
nor U15359 (N_15359,N_12603,N_13251);
or U15360 (N_15360,N_11882,N_14160);
or U15361 (N_15361,N_12869,N_14767);
nand U15362 (N_15362,N_13022,N_14139);
and U15363 (N_15363,N_11001,N_10504);
nand U15364 (N_15364,N_12089,N_14919);
nand U15365 (N_15365,N_13505,N_11892);
and U15366 (N_15366,N_14763,N_13816);
or U15367 (N_15367,N_10473,N_14756);
or U15368 (N_15368,N_12395,N_10920);
or U15369 (N_15369,N_12070,N_11203);
nand U15370 (N_15370,N_12445,N_10172);
and U15371 (N_15371,N_12573,N_11610);
nor U15372 (N_15372,N_14639,N_13402);
nand U15373 (N_15373,N_14634,N_13670);
nor U15374 (N_15374,N_11029,N_11309);
and U15375 (N_15375,N_12857,N_10438);
or U15376 (N_15376,N_12414,N_13668);
and U15377 (N_15377,N_14424,N_10737);
or U15378 (N_15378,N_12125,N_11976);
nand U15379 (N_15379,N_10283,N_14957);
and U15380 (N_15380,N_11039,N_14105);
nand U15381 (N_15381,N_13246,N_10233);
and U15382 (N_15382,N_10773,N_13423);
nor U15383 (N_15383,N_14030,N_13250);
nor U15384 (N_15384,N_13090,N_12295);
nor U15385 (N_15385,N_11455,N_12248);
nor U15386 (N_15386,N_10914,N_11088);
and U15387 (N_15387,N_12336,N_14633);
and U15388 (N_15388,N_12345,N_14750);
nor U15389 (N_15389,N_12288,N_13637);
or U15390 (N_15390,N_11725,N_14406);
and U15391 (N_15391,N_11848,N_14731);
and U15392 (N_15392,N_11964,N_13085);
nand U15393 (N_15393,N_11391,N_12625);
xor U15394 (N_15394,N_12499,N_11519);
or U15395 (N_15395,N_14647,N_13330);
nor U15396 (N_15396,N_12623,N_14197);
nand U15397 (N_15397,N_13853,N_10823);
and U15398 (N_15398,N_11952,N_12362);
or U15399 (N_15399,N_14762,N_10540);
and U15400 (N_15400,N_13854,N_10434);
or U15401 (N_15401,N_11123,N_14072);
or U15402 (N_15402,N_14470,N_13759);
nor U15403 (N_15403,N_13304,N_10896);
and U15404 (N_15404,N_12390,N_11333);
nor U15405 (N_15405,N_13155,N_10781);
nand U15406 (N_15406,N_11315,N_13851);
and U15407 (N_15407,N_10618,N_11960);
or U15408 (N_15408,N_10756,N_10790);
nor U15409 (N_15409,N_11299,N_14720);
or U15410 (N_15410,N_10966,N_13784);
and U15411 (N_15411,N_13537,N_10706);
nand U15412 (N_15412,N_13517,N_10964);
and U15413 (N_15413,N_11671,N_14532);
or U15414 (N_15414,N_13417,N_12451);
and U15415 (N_15415,N_13604,N_11941);
nor U15416 (N_15416,N_12700,N_10073);
nand U15417 (N_15417,N_11497,N_10911);
or U15418 (N_15418,N_12091,N_10816);
or U15419 (N_15419,N_10198,N_13060);
and U15420 (N_15420,N_11301,N_11626);
nor U15421 (N_15421,N_13117,N_12239);
or U15422 (N_15422,N_12568,N_10917);
nor U15423 (N_15423,N_11997,N_12113);
and U15424 (N_15424,N_11845,N_10295);
or U15425 (N_15425,N_10942,N_11742);
or U15426 (N_15426,N_11982,N_13439);
nor U15427 (N_15427,N_12520,N_11971);
and U15428 (N_15428,N_14802,N_11066);
or U15429 (N_15429,N_13674,N_10552);
nor U15430 (N_15430,N_12796,N_13950);
nor U15431 (N_15431,N_12738,N_11121);
nand U15432 (N_15432,N_11991,N_11468);
nand U15433 (N_15433,N_11896,N_12114);
nand U15434 (N_15434,N_13745,N_13848);
and U15435 (N_15435,N_12862,N_13265);
and U15436 (N_15436,N_13058,N_14365);
nand U15437 (N_15437,N_11659,N_11692);
nor U15438 (N_15438,N_10381,N_10114);
nand U15439 (N_15439,N_11017,N_12800);
nand U15440 (N_15440,N_13167,N_13711);
nand U15441 (N_15441,N_13924,N_14316);
nand U15442 (N_15442,N_13727,N_14530);
nor U15443 (N_15443,N_11898,N_12409);
nor U15444 (N_15444,N_10772,N_13689);
and U15445 (N_15445,N_11332,N_10634);
nand U15446 (N_15446,N_10944,N_11450);
nand U15447 (N_15447,N_14378,N_12249);
nor U15448 (N_15448,N_12884,N_11360);
and U15449 (N_15449,N_12496,N_10758);
or U15450 (N_15450,N_14056,N_13519);
nor U15451 (N_15451,N_12073,N_14149);
and U15452 (N_15452,N_10413,N_13287);
or U15453 (N_15453,N_11325,N_12852);
or U15454 (N_15454,N_12639,N_10788);
nor U15455 (N_15455,N_10850,N_14243);
and U15456 (N_15456,N_11366,N_14971);
and U15457 (N_15457,N_12968,N_14951);
and U15458 (N_15458,N_13255,N_12656);
or U15459 (N_15459,N_14501,N_10794);
nand U15460 (N_15460,N_12162,N_11910);
and U15461 (N_15461,N_13808,N_12552);
nand U15462 (N_15462,N_12660,N_11097);
nor U15463 (N_15463,N_13091,N_10455);
or U15464 (N_15464,N_12894,N_11618);
or U15465 (N_15465,N_10364,N_14675);
nor U15466 (N_15466,N_12837,N_13915);
or U15467 (N_15467,N_12741,N_13598);
nand U15468 (N_15468,N_10106,N_14772);
and U15469 (N_15469,N_14573,N_11018);
or U15470 (N_15470,N_12327,N_11587);
nand U15471 (N_15471,N_10119,N_10677);
and U15472 (N_15472,N_10032,N_11087);
nand U15473 (N_15473,N_14224,N_12318);
nor U15474 (N_15474,N_14753,N_12401);
and U15475 (N_15475,N_10458,N_10260);
and U15476 (N_15476,N_12472,N_14064);
and U15477 (N_15477,N_14201,N_10156);
nor U15478 (N_15478,N_10386,N_13581);
or U15479 (N_15479,N_11220,N_13590);
nand U15480 (N_15480,N_13798,N_14937);
nor U15481 (N_15481,N_11142,N_11005);
nor U15482 (N_15482,N_14575,N_12886);
and U15483 (N_15483,N_11246,N_14458);
nor U15484 (N_15484,N_11258,N_13956);
nand U15485 (N_15485,N_12133,N_13918);
and U15486 (N_15486,N_10141,N_10837);
nand U15487 (N_15487,N_12426,N_13237);
and U15488 (N_15488,N_13709,N_10414);
or U15489 (N_15489,N_12232,N_11691);
nand U15490 (N_15490,N_10624,N_11769);
nand U15491 (N_15491,N_11160,N_14725);
and U15492 (N_15492,N_12165,N_11103);
nor U15493 (N_15493,N_12743,N_13350);
and U15494 (N_15494,N_12860,N_13969);
or U15495 (N_15495,N_12122,N_11852);
nor U15496 (N_15496,N_13471,N_13778);
nand U15497 (N_15497,N_12605,N_13651);
nor U15498 (N_15498,N_13791,N_10935);
and U15499 (N_15499,N_13343,N_13045);
or U15500 (N_15500,N_13753,N_13510);
and U15501 (N_15501,N_12947,N_12180);
nor U15502 (N_15502,N_13622,N_13717);
nor U15503 (N_15503,N_13180,N_11086);
and U15504 (N_15504,N_11422,N_11744);
and U15505 (N_15505,N_12779,N_12430);
nor U15506 (N_15506,N_13616,N_12234);
and U15507 (N_15507,N_12466,N_12097);
nor U15508 (N_15508,N_14706,N_12159);
or U15509 (N_15509,N_14223,N_11552);
and U15510 (N_15510,N_14301,N_14827);
and U15511 (N_15511,N_10193,N_12285);
nand U15512 (N_15512,N_14507,N_11916);
xnor U15513 (N_15513,N_11890,N_12412);
and U15514 (N_15514,N_14888,N_13682);
and U15515 (N_15515,N_14815,N_14236);
or U15516 (N_15516,N_14986,N_14100);
or U15517 (N_15517,N_13499,N_13936);
nor U15518 (N_15518,N_12889,N_12631);
and U15519 (N_15519,N_10603,N_13974);
and U15520 (N_15520,N_10205,N_13002);
nor U15521 (N_15521,N_13264,N_11735);
nand U15522 (N_15522,N_13082,N_14266);
nor U15523 (N_15523,N_10901,N_10858);
nand U15524 (N_15524,N_10861,N_12554);
nand U15525 (N_15525,N_11905,N_10777);
or U15526 (N_15526,N_13017,N_11625);
or U15527 (N_15527,N_13803,N_10241);
nor U15528 (N_15528,N_13802,N_11822);
and U15529 (N_15529,N_14422,N_14533);
or U15530 (N_15530,N_13740,N_14537);
nor U15531 (N_15531,N_13688,N_12289);
and U15532 (N_15532,N_14384,N_14228);
or U15533 (N_15533,N_10994,N_11939);
or U15534 (N_15534,N_14329,N_13312);
and U15535 (N_15535,N_12210,N_14229);
nand U15536 (N_15536,N_12930,N_11853);
or U15537 (N_15537,N_14182,N_11458);
or U15538 (N_15538,N_13478,N_11791);
or U15539 (N_15539,N_13975,N_12006);
nand U15540 (N_15540,N_14187,N_13432);
nand U15541 (N_15541,N_11232,N_12476);
and U15542 (N_15542,N_13686,N_10206);
and U15543 (N_15543,N_14712,N_14645);
or U15544 (N_15544,N_13414,N_11738);
and U15545 (N_15545,N_11421,N_13691);
and U15546 (N_15546,N_11061,N_11440);
nand U15547 (N_15547,N_10870,N_12556);
nand U15548 (N_15548,N_14091,N_10037);
and U15549 (N_15549,N_14605,N_11606);
nand U15550 (N_15550,N_13551,N_11727);
nand U15551 (N_15551,N_14456,N_12152);
or U15552 (N_15552,N_11762,N_10396);
nor U15553 (N_15553,N_14459,N_11837);
and U15554 (N_15554,N_11072,N_12138);
or U15555 (N_15555,N_12515,N_13037);
and U15556 (N_15556,N_12391,N_11772);
or U15557 (N_15557,N_14437,N_12014);
nand U15558 (N_15558,N_10819,N_12141);
and U15559 (N_15559,N_13109,N_10453);
and U15560 (N_15560,N_13282,N_10389);
or U15561 (N_15561,N_10704,N_11131);
nand U15562 (N_15562,N_13495,N_11286);
and U15563 (N_15563,N_11502,N_11247);
or U15564 (N_15564,N_14315,N_12891);
nand U15565 (N_15565,N_12205,N_14142);
and U15566 (N_15566,N_12381,N_12002);
nand U15567 (N_15567,N_13624,N_10498);
and U15568 (N_15568,N_10713,N_12222);
or U15569 (N_15569,N_12291,N_11437);
or U15570 (N_15570,N_13133,N_12216);
nand U15571 (N_15571,N_12335,N_14811);
or U15572 (N_15572,N_14219,N_11657);
or U15573 (N_15573,N_10003,N_11687);
and U15574 (N_15574,N_14220,N_11254);
or U15575 (N_15575,N_11633,N_14235);
and U15576 (N_15576,N_14212,N_13823);
nor U15577 (N_15577,N_12638,N_12227);
nand U15578 (N_15578,N_10016,N_12281);
nand U15579 (N_15579,N_10085,N_10312);
nand U15580 (N_15580,N_13917,N_14366);
and U15581 (N_15581,N_12775,N_11936);
and U15582 (N_15582,N_13757,N_13567);
nor U15583 (N_15583,N_13019,N_10539);
or U15584 (N_15584,N_13143,N_11900);
or U15585 (N_15585,N_12382,N_14710);
nand U15586 (N_15586,N_12598,N_11875);
nand U15587 (N_15587,N_12941,N_14925);
or U15588 (N_15588,N_11191,N_10764);
nor U15589 (N_15589,N_11581,N_13696);
nand U15590 (N_15590,N_10785,N_10173);
and U15591 (N_15591,N_13205,N_10072);
nor U15592 (N_15592,N_12525,N_12776);
or U15593 (N_15593,N_13723,N_11327);
nor U15594 (N_15594,N_13374,N_11876);
nor U15595 (N_15595,N_13665,N_12766);
nor U15596 (N_15596,N_12340,N_11222);
nor U15597 (N_15597,N_13986,N_12333);
and U15598 (N_15598,N_10612,N_14766);
nor U15599 (N_15599,N_13361,N_13443);
nor U15600 (N_15600,N_14014,N_12176);
and U15601 (N_15601,N_10502,N_14897);
and U15602 (N_15602,N_13072,N_10101);
and U15603 (N_15603,N_14157,N_13511);
nand U15604 (N_15604,N_11185,N_10532);
or U15605 (N_15605,N_10686,N_14933);
nor U15606 (N_15606,N_11467,N_14892);
or U15607 (N_15607,N_12795,N_14383);
and U15608 (N_15608,N_13430,N_13597);
and U15609 (N_15609,N_10811,N_12763);
nor U15610 (N_15610,N_10064,N_13396);
and U15611 (N_15611,N_14005,N_13300);
or U15612 (N_15612,N_13187,N_12449);
or U15613 (N_15613,N_14518,N_11781);
or U15614 (N_15614,N_12737,N_11475);
and U15615 (N_15615,N_10800,N_13763);
nand U15616 (N_15616,N_10883,N_12046);
nand U15617 (N_15617,N_11394,N_11076);
nor U15618 (N_15618,N_13627,N_11867);
nand U15619 (N_15619,N_11545,N_13171);
nor U15620 (N_15620,N_12200,N_13606);
or U15621 (N_15621,N_13123,N_11752);
nand U15622 (N_15622,N_14661,N_14085);
and U15623 (N_15623,N_14425,N_11092);
and U15624 (N_15624,N_12047,N_10213);
nor U15625 (N_15625,N_13259,N_13509);
xor U15626 (N_15626,N_14423,N_11465);
nor U15627 (N_15627,N_12422,N_14601);
nor U15628 (N_15628,N_13857,N_14020);
nand U15629 (N_15629,N_14809,N_11860);
or U15630 (N_15630,N_14793,N_13996);
or U15631 (N_15631,N_14896,N_12350);
nand U15632 (N_15632,N_13284,N_13283);
nor U15633 (N_15633,N_14025,N_13656);
and U15634 (N_15634,N_10134,N_14848);
and U15635 (N_15635,N_11260,N_10776);
and U15636 (N_15636,N_13363,N_14071);
or U15637 (N_15637,N_12690,N_10442);
nand U15638 (N_15638,N_12375,N_10609);
and U15639 (N_15639,N_13609,N_13595);
and U15640 (N_15640,N_13625,N_10248);
or U15641 (N_15641,N_14073,N_10534);
or U15642 (N_15642,N_13351,N_13049);
or U15643 (N_15643,N_12826,N_12720);
nand U15644 (N_15644,N_14398,N_12261);
nor U15645 (N_15645,N_11003,N_13847);
xnor U15646 (N_15646,N_14394,N_13087);
nor U15647 (N_15647,N_13501,N_10436);
and U15648 (N_15648,N_10292,N_12425);
and U15649 (N_15649,N_14079,N_14411);
or U15650 (N_15650,N_10354,N_11899);
nand U15651 (N_15651,N_12565,N_11357);
nand U15652 (N_15652,N_11402,N_12128);
or U15653 (N_15653,N_10126,N_11054);
and U15654 (N_15654,N_10086,N_14854);
or U15655 (N_15655,N_13572,N_11190);
nand U15656 (N_15656,N_14562,N_12505);
and U15657 (N_15657,N_12224,N_13564);
or U15658 (N_15658,N_10194,N_10629);
nor U15659 (N_15659,N_12192,N_11601);
or U15660 (N_15660,N_11496,N_14615);
or U15661 (N_15661,N_13372,N_12049);
or U15662 (N_15662,N_10435,N_12590);
and U15663 (N_15663,N_11215,N_11317);
nand U15664 (N_15664,N_13661,N_13279);
nand U15665 (N_15665,N_14814,N_14075);
and U15666 (N_15666,N_13882,N_11165);
nor U15667 (N_15667,N_10009,N_12948);
nor U15668 (N_15668,N_10830,N_14882);
and U15669 (N_15669,N_10475,N_12555);
nor U15670 (N_15670,N_10950,N_14863);
nor U15671 (N_15671,N_14618,N_10856);
and U15672 (N_15672,N_10171,N_11874);
and U15673 (N_15673,N_12686,N_12924);
nand U15674 (N_15674,N_13079,N_14042);
or U15675 (N_15675,N_11356,N_12617);
nor U15676 (N_15676,N_14932,N_10307);
nand U15677 (N_15677,N_14321,N_10521);
and U15678 (N_15678,N_11851,N_11776);
or U15679 (N_15679,N_12870,N_11136);
or U15680 (N_15680,N_12167,N_10462);
nand U15681 (N_15681,N_14688,N_13337);
nand U15682 (N_15682,N_13767,N_11372);
nand U15683 (N_15683,N_11320,N_11216);
or U15684 (N_15684,N_11617,N_12950);
nor U15685 (N_15685,N_12154,N_11833);
nand U15686 (N_15686,N_13905,N_13083);
xnor U15687 (N_15687,N_12821,N_13313);
nand U15688 (N_15688,N_13871,N_14141);
nor U15689 (N_15689,N_14635,N_12095);
nor U15690 (N_15690,N_13793,N_11685);
or U15691 (N_15691,N_12981,N_10237);
and U15692 (N_15692,N_12030,N_10940);
or U15693 (N_15693,N_10298,N_13931);
nor U15694 (N_15694,N_10638,N_10149);
nand U15695 (N_15695,N_10426,N_11487);
nor U15696 (N_15696,N_14845,N_12050);
nand U15697 (N_15697,N_13967,N_10518);
and U15698 (N_15698,N_10042,N_11654);
nor U15699 (N_15699,N_10708,N_13185);
and U15700 (N_15700,N_13150,N_11125);
nor U15701 (N_15701,N_10760,N_10945);
or U15702 (N_15702,N_12121,N_10033);
nor U15703 (N_15703,N_13873,N_11346);
nand U15704 (N_15704,N_12419,N_12302);
or U15705 (N_15705,N_13101,N_10730);
and U15706 (N_15706,N_12446,N_14782);
or U15707 (N_15707,N_10118,N_13787);
nand U15708 (N_15708,N_14820,N_13483);
or U15709 (N_15709,N_14351,N_10581);
or U15710 (N_15710,N_10694,N_14221);
nor U15711 (N_15711,N_10422,N_14457);
nand U15712 (N_15712,N_11326,N_14047);
nor U15713 (N_15713,N_13940,N_14926);
nand U15714 (N_15714,N_13340,N_14281);
and U15715 (N_15715,N_10239,N_11520);
or U15716 (N_15716,N_14700,N_12209);
and U15717 (N_15717,N_14446,N_14427);
or U15718 (N_15718,N_13535,N_13218);
or U15719 (N_15719,N_10641,N_13406);
and U15720 (N_15720,N_10265,N_14326);
or U15721 (N_15721,N_12084,N_11266);
nand U15722 (N_15722,N_12691,N_11243);
or U15723 (N_15723,N_13426,N_13479);
nor U15724 (N_15724,N_10484,N_14026);
and U15725 (N_15725,N_14024,N_11147);
or U15726 (N_15726,N_13845,N_11211);
and U15727 (N_15727,N_11408,N_11033);
nand U15728 (N_15728,N_14883,N_13737);
nor U15729 (N_15729,N_13557,N_13916);
or U15730 (N_15730,N_10281,N_14905);
nor U15731 (N_15731,N_12018,N_12348);
and U15732 (N_15732,N_13368,N_11237);
nand U15733 (N_15733,N_12062,N_14702);
nor U15734 (N_15734,N_13010,N_10878);
nand U15735 (N_15735,N_10733,N_11998);
nand U15736 (N_15736,N_13390,N_13935);
nor U15737 (N_15737,N_11307,N_10727);
nand U15738 (N_15738,N_12298,N_13052);
nor U15739 (N_15739,N_12969,N_10061);
nand U15740 (N_15740,N_14869,N_11790);
nor U15741 (N_15741,N_11296,N_14217);
and U15742 (N_15742,N_13339,N_12468);
nand U15743 (N_15743,N_12024,N_12789);
and U15744 (N_15744,N_11358,N_10428);
nor U15745 (N_15745,N_13097,N_14770);
and U15746 (N_15746,N_14078,N_10931);
nand U15747 (N_15747,N_13526,N_14697);
or U15748 (N_15748,N_11137,N_10221);
nor U15749 (N_15749,N_14650,N_12984);
or U15750 (N_15750,N_12830,N_14641);
nor U15751 (N_15751,N_11909,N_11541);
xnor U15752 (N_15752,N_11710,N_14463);
nand U15753 (N_15753,N_14156,N_14527);
nor U15754 (N_15754,N_14946,N_11032);
and U15755 (N_15755,N_12975,N_11277);
nand U15756 (N_15756,N_11133,N_13862);
nand U15757 (N_15757,N_10334,N_13614);
and U15758 (N_15758,N_11012,N_12799);
and U15759 (N_15759,N_10992,N_11170);
nand U15760 (N_15760,N_14245,N_10667);
and U15761 (N_15761,N_10416,N_10608);
nand U15762 (N_15762,N_13574,N_12320);
or U15763 (N_15763,N_14296,N_14227);
nor U15764 (N_15764,N_14548,N_14895);
or U15765 (N_15765,N_10160,N_11180);
and U15766 (N_15766,N_10749,N_13481);
or U15767 (N_15767,N_11996,N_10855);
nor U15768 (N_15768,N_10957,N_14070);
nor U15769 (N_15769,N_11293,N_12936);
xor U15770 (N_15770,N_12734,N_14311);
and U15771 (N_15771,N_14549,N_14867);
nor U15772 (N_15772,N_13398,N_13534);
and U15773 (N_15773,N_12866,N_11800);
and U15774 (N_15774,N_11793,N_12702);
nand U15775 (N_15775,N_11127,N_11488);
and U15776 (N_15776,N_12600,N_10492);
and U15777 (N_15777,N_11990,N_10423);
and U15778 (N_15778,N_14364,N_12416);
nand U15779 (N_15779,N_14797,N_11605);
and U15780 (N_15780,N_11331,N_12581);
and U15781 (N_15781,N_12998,N_11415);
and U15782 (N_15782,N_10325,N_13213);
nand U15783 (N_15783,N_11268,N_13994);
nor U15784 (N_15784,N_12580,N_14027);
or U15785 (N_15785,N_13685,N_10580);
and U15786 (N_15786,N_10125,N_14041);
or U15787 (N_15787,N_11643,N_13207);
nand U15788 (N_15788,N_14593,N_13493);
nand U15789 (N_15789,N_13584,N_14455);
and U15790 (N_15790,N_13518,N_13498);
xnor U15791 (N_15791,N_10328,N_12267);
nor U15792 (N_15792,N_12902,N_13742);
nor U15793 (N_15793,N_11396,N_11802);
nor U15794 (N_15794,N_11132,N_13680);
and U15795 (N_15795,N_12319,N_12300);
nand U15796 (N_15796,N_10488,N_10881);
nor U15797 (N_15797,N_13531,N_10511);
or U15798 (N_15798,N_11536,N_11778);
nor U15799 (N_15799,N_14692,N_10135);
and U15800 (N_15800,N_13130,N_14642);
nand U15801 (N_15801,N_14324,N_12762);
xor U15802 (N_15802,N_11938,N_14890);
nor U15803 (N_15803,N_13675,N_12490);
nand U15804 (N_15804,N_11508,N_10680);
or U15805 (N_15805,N_11071,N_10770);
or U15806 (N_15806,N_10553,N_13474);
nand U15807 (N_15807,N_11197,N_13170);
nand U15808 (N_15808,N_13344,N_12613);
and U15809 (N_15809,N_10196,N_10561);
nand U15810 (N_15810,N_13464,N_12954);
nor U15811 (N_15811,N_14962,N_13933);
or U15812 (N_15812,N_14040,N_14453);
nand U15813 (N_15813,N_14719,N_10522);
or U15814 (N_15814,N_12098,N_11674);
or U15815 (N_15815,N_12945,N_11267);
xnor U15816 (N_15816,N_11377,N_12041);
and U15817 (N_15817,N_11281,N_10002);
and U15818 (N_15818,N_14564,N_10088);
nand U15819 (N_15819,N_12297,N_12169);
and U15820 (N_15820,N_14265,N_11345);
nor U15821 (N_15821,N_13826,N_12076);
nor U15822 (N_15822,N_14840,N_12276);
nor U15823 (N_15823,N_10587,N_11324);
or U15824 (N_15824,N_14341,N_11022);
nor U15825 (N_15825,N_10388,N_14994);
or U15826 (N_15826,N_10229,N_11383);
nand U15827 (N_15827,N_14256,N_12454);
or U15828 (N_15828,N_10082,N_12646);
nand U15829 (N_15829,N_13219,N_13111);
and U15830 (N_15830,N_11798,N_13568);
nor U15831 (N_15831,N_11849,N_13141);
and U15832 (N_15832,N_11694,N_13177);
or U15833 (N_15833,N_13869,N_13592);
or U15834 (N_15834,N_10663,N_12398);
nand U15835 (N_15835,N_13416,N_13429);
nand U15836 (N_15836,N_14330,N_10755);
nand U15837 (N_15837,N_10812,N_11576);
nor U15838 (N_15838,N_14818,N_14261);
and U15839 (N_15839,N_14825,N_10866);
or U15840 (N_15840,N_10547,N_13858);
and U15841 (N_15841,N_10023,N_11779);
nor U15842 (N_15842,N_11970,N_10107);
or U15843 (N_15843,N_10771,N_12995);
and U15844 (N_15844,N_13275,N_13647);
nor U15845 (N_15845,N_11175,N_12861);
or U15846 (N_15846,N_11613,N_13599);
and U15847 (N_15847,N_10512,N_12182);
nor U15848 (N_15848,N_13121,N_10373);
and U15849 (N_15849,N_10376,N_13542);
or U15850 (N_15850,N_14595,N_10347);
nand U15851 (N_15851,N_11291,N_12713);
or U15852 (N_15852,N_14308,N_12193);
nand U15853 (N_15853,N_12099,N_11414);
or U15854 (N_15854,N_12976,N_14912);
or U15855 (N_15855,N_11571,N_12712);
nor U15856 (N_15856,N_13692,N_13174);
nand U15857 (N_15857,N_13249,N_12827);
nor U15858 (N_15858,N_13725,N_14451);
or U15859 (N_15859,N_14120,N_12616);
and U15860 (N_15860,N_13909,N_12170);
and U15861 (N_15861,N_14000,N_14603);
and U15862 (N_15862,N_12640,N_13385);
nand U15863 (N_15863,N_13710,N_10517);
and U15864 (N_15864,N_14043,N_14240);
or U15865 (N_15865,N_11269,N_14961);
and U15866 (N_15866,N_13547,N_10659);
or U15867 (N_15867,N_13811,N_14859);
nand U15868 (N_15868,N_13088,N_13262);
nand U15869 (N_15869,N_11289,N_11328);
nor U15870 (N_15870,N_14183,N_11079);
nor U15871 (N_15871,N_12740,N_12279);
nand U15872 (N_15872,N_14066,N_14117);
or U15873 (N_15873,N_13874,N_10545);
nor U15874 (N_15874,N_14244,N_11621);
nor U15875 (N_15875,N_12265,N_12206);
nand U15876 (N_15876,N_10100,N_10322);
nand U15877 (N_15877,N_11051,N_13322);
nor U15878 (N_15878,N_12410,N_11866);
nor U15879 (N_15879,N_11361,N_14664);
or U15880 (N_15880,N_14337,N_12236);
or U15881 (N_15881,N_12518,N_12380);
and U15882 (N_15882,N_10702,N_14478);
nor U15883 (N_15883,N_11231,N_14958);
nor U15884 (N_15884,N_10015,N_13999);
or U15885 (N_15885,N_12818,N_10728);
nor U15886 (N_15886,N_13527,N_11917);
and U15887 (N_15887,N_14407,N_12633);
or U15888 (N_15888,N_13952,N_14776);
nor U15889 (N_15889,N_10946,N_10633);
and U15890 (N_15890,N_14200,N_11572);
nor U15891 (N_15891,N_14979,N_12484);
or U15892 (N_15892,N_10912,N_14924);
nand U15893 (N_15893,N_13482,N_13484);
and U15894 (N_15894,N_12788,N_10501);
or U15895 (N_15895,N_14977,N_11922);
and U15896 (N_15896,N_11764,N_12501);
nor U15897 (N_15897,N_11436,N_12247);
nor U15898 (N_15898,N_14137,N_14715);
and U15899 (N_15899,N_10909,N_13028);
nor U15900 (N_15900,N_10797,N_11693);
or U15901 (N_15901,N_12842,N_14230);
nand U15902 (N_15902,N_12080,N_13770);
or U15903 (N_15903,N_11698,N_10035);
nand U15904 (N_15904,N_13314,N_12716);
nand U15905 (N_15905,N_11196,N_13708);
nor U15906 (N_15906,N_12641,N_14196);
nand U15907 (N_15907,N_12688,N_14880);
and U15908 (N_15908,N_14598,N_13446);
nor U15909 (N_15909,N_11696,N_10161);
or U15910 (N_15910,N_10097,N_12246);
and U15911 (N_15911,N_11835,N_13294);
and U15912 (N_15912,N_10323,N_13160);
and U15913 (N_15913,N_11016,N_10232);
nand U15914 (N_15914,N_14060,N_13731);
nand U15915 (N_15915,N_14335,N_13835);
nor U15916 (N_15916,N_14722,N_12465);
or U15917 (N_15917,N_14812,N_13162);
and U15918 (N_15918,N_10808,N_10165);
nor U15919 (N_15919,N_12280,N_10362);
nand U15920 (N_15920,N_11709,N_12745);
nand U15921 (N_15921,N_10123,N_11785);
nor U15922 (N_15922,N_12653,N_12388);
nand U15923 (N_15923,N_12118,N_12153);
and U15924 (N_15924,N_11256,N_14805);
nand U15925 (N_15925,N_12082,N_13619);
xor U15926 (N_15926,N_12231,N_13653);
nor U15927 (N_15927,N_14444,N_11043);
nand U15928 (N_15928,N_12915,N_10672);
or U15929 (N_15929,N_13644,N_13842);
nor U15930 (N_15930,N_11953,N_11002);
nand U15931 (N_15931,N_10411,N_13032);
nor U15932 (N_15932,N_13961,N_12758);
or U15933 (N_15933,N_12088,N_14738);
nor U15934 (N_15934,N_13342,N_13514);
and U15935 (N_15935,N_14097,N_12334);
nand U15936 (N_15936,N_10535,N_13260);
nand U15937 (N_15937,N_11903,N_11885);
and U15938 (N_15938,N_10108,N_10871);
nor U15939 (N_15939,N_10939,N_14127);
nor U15940 (N_15940,N_11729,N_12540);
and U15941 (N_15941,N_14008,N_10863);
and U15942 (N_15942,N_13291,N_12913);
nand U15943 (N_15943,N_14668,N_10683);
and U15944 (N_15944,N_12611,N_14269);
or U15945 (N_15945,N_13523,N_11059);
nand U15946 (N_15946,N_11803,N_14279);
nand U15947 (N_15947,N_12719,N_11730);
nor U15948 (N_15948,N_11322,N_13269);
nand U15949 (N_15949,N_10710,N_11809);
nor U15950 (N_15950,N_10207,N_13536);
and U15951 (N_15951,N_10711,N_14701);
and U15952 (N_15952,N_10853,N_10297);
or U15953 (N_15953,N_10869,N_14711);
nand U15954 (N_15954,N_11884,N_12718);
or U15955 (N_15955,N_13463,N_14631);
nor U15956 (N_15956,N_13943,N_12724);
or U15957 (N_15957,N_13806,N_13115);
and U15958 (N_15958,N_11008,N_14462);
nor U15959 (N_15959,N_11166,N_12373);
nand U15960 (N_15960,N_13290,N_10962);
and U15961 (N_15961,N_11321,N_11110);
or U15962 (N_15962,N_12037,N_12447);
nor U15963 (N_15963,N_13818,N_12696);
nor U15964 (N_15964,N_10689,N_14663);
nor U15965 (N_15965,N_12177,N_10500);
or U15966 (N_15966,N_13642,N_10153);
nand U15967 (N_15967,N_12701,N_12308);
or U15968 (N_15968,N_12757,N_10244);
and U15969 (N_15969,N_11094,N_12240);
nand U15970 (N_15970,N_13601,N_13698);
or U15971 (N_15971,N_13201,N_10440);
nand U15972 (N_15972,N_10300,N_10145);
and U15973 (N_15973,N_10131,N_13315);
nand U15974 (N_15974,N_13435,N_11430);
nor U15975 (N_15975,N_10988,N_10342);
or U15976 (N_15976,N_14798,N_12878);
nor U15977 (N_15977,N_11962,N_12218);
or U15978 (N_15978,N_11099,N_13839);
nor U15979 (N_15979,N_11846,N_13234);
nor U15980 (N_15980,N_13701,N_14567);
nand U15981 (N_15981,N_12052,N_13880);
nor U15982 (N_15982,N_13833,N_11983);
nand U15983 (N_15983,N_12199,N_11575);
xor U15984 (N_15984,N_12683,N_13026);
and U15985 (N_15985,N_12443,N_11492);
or U15986 (N_15986,N_12032,N_13247);
nor U15987 (N_15987,N_10147,N_14943);
or U15988 (N_15988,N_11273,N_14861);
or U15989 (N_15989,N_14214,N_11122);
and U15990 (N_15990,N_10658,N_14918);
or U15991 (N_15991,N_12321,N_12831);
or U15992 (N_15992,N_13894,N_11515);
and U15993 (N_15993,N_12574,N_14426);
or U15994 (N_15994,N_10786,N_14777);
nand U15995 (N_15995,N_14847,N_11682);
and U15996 (N_15996,N_11221,N_13041);
or U15997 (N_15997,N_12871,N_12475);
and U15998 (N_15998,N_10916,N_11089);
and U15999 (N_15999,N_12925,N_14684);
or U16000 (N_16000,N_13775,N_11723);
nand U16001 (N_16001,N_11750,N_10600);
nand U16002 (N_16002,N_10304,N_13303);
and U16003 (N_16003,N_10675,N_12548);
or U16004 (N_16004,N_11491,N_10595);
nand U16005 (N_16005,N_13103,N_10012);
and U16006 (N_16006,N_13795,N_11034);
or U16007 (N_16007,N_13074,N_12450);
nor U16008 (N_16008,N_13843,N_12692);
nor U16009 (N_16009,N_10671,N_11823);
nor U16010 (N_16010,N_12197,N_11746);
or U16011 (N_16011,N_12817,N_10903);
or U16012 (N_16012,N_10577,N_13230);
and U16013 (N_16013,N_12706,N_14114);
and U16014 (N_16014,N_13503,N_10885);
nor U16015 (N_16015,N_12079,N_14927);
or U16016 (N_16016,N_10441,N_13724);
and U16017 (N_16017,N_10622,N_14644);
and U16018 (N_16018,N_11010,N_11338);
nand U16019 (N_16019,N_11257,N_13056);
nor U16020 (N_16020,N_10187,N_13718);
nor U16021 (N_16021,N_11169,N_13437);
nor U16022 (N_16022,N_13878,N_14813);
nand U16023 (N_16023,N_10401,N_13594);
or U16024 (N_16024,N_14741,N_10765);
nand U16025 (N_16025,N_11556,N_12174);
and U16026 (N_16026,N_11985,N_12599);
nand U16027 (N_16027,N_13442,N_14570);
nor U16028 (N_16028,N_13127,N_14665);
nor U16029 (N_16029,N_11665,N_11407);
and U16030 (N_16030,N_14474,N_12150);
nand U16031 (N_16031,N_11913,N_14552);
nor U16032 (N_16032,N_14352,N_11999);
or U16033 (N_16033,N_14188,N_10739);
nor U16034 (N_16034,N_14044,N_14758);
and U16035 (N_16035,N_11920,N_10262);
nor U16036 (N_16036,N_14166,N_13671);
nor U16037 (N_16037,N_10294,N_10208);
nand U16038 (N_16038,N_14338,N_13722);
and U16039 (N_16039,N_12053,N_10938);
and U16040 (N_16040,N_13009,N_10907);
or U16041 (N_16041,N_11213,N_14354);
and U16042 (N_16042,N_10398,N_11801);
or U16043 (N_16043,N_14369,N_13139);
and U16044 (N_16044,N_11479,N_10974);
and U16045 (N_16045,N_14232,N_12020);
nor U16046 (N_16046,N_10817,N_12235);
nor U16047 (N_16047,N_10223,N_12256);
nand U16048 (N_16048,N_14511,N_12698);
nand U16049 (N_16049,N_10093,N_10296);
nand U16050 (N_16050,N_11661,N_11313);
and U16051 (N_16051,N_10647,N_10698);
nand U16052 (N_16052,N_13765,N_13387);
or U16053 (N_16053,N_10775,N_13204);
or U16054 (N_16054,N_11511,N_14864);
nor U16055 (N_16055,N_14484,N_10188);
or U16056 (N_16056,N_13946,N_13664);
nor U16057 (N_16057,N_10519,N_14659);
nor U16058 (N_16058,N_14830,N_10017);
and U16059 (N_16059,N_10742,N_11512);
nor U16060 (N_16060,N_11955,N_10782);
nand U16061 (N_16061,N_12467,N_11474);
nand U16062 (N_16062,N_10140,N_13163);
nand U16063 (N_16063,N_12078,N_14159);
or U16064 (N_16064,N_11423,N_14328);
nand U16065 (N_16065,N_13989,N_11399);
and U16066 (N_16066,N_14443,N_10390);
or U16067 (N_16067,N_12999,N_11865);
or U16068 (N_16068,N_12178,N_13104);
nand U16069 (N_16069,N_10065,N_12689);
or U16070 (N_16070,N_12312,N_12471);
or U16071 (N_16071,N_10951,N_14023);
and U16072 (N_16072,N_14363,N_10495);
nor U16073 (N_16073,N_12517,N_13216);
and U16074 (N_16074,N_10872,N_13161);
nand U16075 (N_16075,N_10841,N_14528);
nor U16076 (N_16076,N_10092,N_11093);
or U16077 (N_16077,N_12498,N_13062);
and U16078 (N_16078,N_11412,N_13308);
or U16079 (N_16079,N_10650,N_10997);
nand U16080 (N_16080,N_10558,N_14673);
nor U16081 (N_16081,N_11834,N_12973);
nor U16082 (N_16082,N_14403,N_13288);
nand U16083 (N_16083,N_11179,N_10266);
and U16084 (N_16084,N_12510,N_12131);
and U16085 (N_16085,N_14824,N_11514);
and U16086 (N_16086,N_12044,N_13470);
and U16087 (N_16087,N_12780,N_11429);
or U16088 (N_16088,N_14773,N_12022);
nand U16089 (N_16089,N_11967,N_14346);
nand U16090 (N_16090,N_10310,N_11804);
nor U16091 (N_16091,N_10452,N_11770);
or U16092 (N_16092,N_14799,N_12033);
or U16093 (N_16093,N_12767,N_14572);
and U16094 (N_16094,N_14504,N_11102);
or U16095 (N_16095,N_11278,N_12010);
nand U16096 (N_16096,N_14262,N_11788);
nand U16097 (N_16097,N_10991,N_11622);
and U16098 (N_16098,N_10005,N_13189);
nand U16099 (N_16099,N_14794,N_13561);
or U16100 (N_16100,N_11636,N_11201);
or U16101 (N_16101,N_11897,N_12494);
and U16102 (N_16102,N_14395,N_14239);
and U16103 (N_16103,N_13679,N_13252);
nand U16104 (N_16104,N_11639,N_13863);
or U16105 (N_16105,N_10104,N_11248);
nand U16106 (N_16106,N_12662,N_10170);
nand U16107 (N_16107,N_11554,N_14432);
and U16108 (N_16108,N_13522,N_12626);
nor U16109 (N_16109,N_10556,N_12987);
and U16110 (N_16110,N_12228,N_14628);
nor U16111 (N_16111,N_11550,N_13865);
nor U16112 (N_16112,N_11516,N_13050);
nand U16113 (N_16113,N_14342,N_12317);
and U16114 (N_16114,N_12634,N_10692);
or U16115 (N_16115,N_13911,N_13243);
and U16116 (N_16116,N_10983,N_12481);
and U16117 (N_16117,N_10833,N_10516);
nand U16118 (N_16118,N_14136,N_12157);
and U16119 (N_16119,N_11205,N_11925);
nand U16120 (N_16120,N_12896,N_14774);
and U16121 (N_16121,N_14929,N_14500);
or U16122 (N_16122,N_10227,N_14356);
nor U16123 (N_16123,N_13166,N_13012);
or U16124 (N_16124,N_12252,N_14129);
nand U16125 (N_16125,N_14723,N_12083);
nand U16126 (N_16126,N_13197,N_14257);
nand U16127 (N_16127,N_12566,N_12650);
and U16128 (N_16128,N_14760,N_14996);
and U16129 (N_16129,N_13948,N_12394);
nor U16130 (N_16130,N_11927,N_13070);
and U16131 (N_16131,N_10457,N_12093);
nor U16132 (N_16132,N_12843,N_14810);
nand U16133 (N_16133,N_14826,N_10890);
and U16134 (N_16134,N_14022,N_14714);
or U16135 (N_16135,N_10700,N_13345);
nand U16136 (N_16136,N_12695,N_14123);
or U16137 (N_16137,N_12156,N_12072);
nand U16138 (N_16138,N_13508,N_10494);
and U16139 (N_16139,N_14133,N_13292);
nand U16140 (N_16140,N_14886,N_11631);
or U16141 (N_16141,N_10277,N_13241);
nor U16142 (N_16142,N_12310,N_11279);
or U16143 (N_16143,N_10929,N_14401);
or U16144 (N_16144,N_12777,N_13006);
nor U16145 (N_16145,N_11038,N_14332);
or U16146 (N_16146,N_13684,N_12341);
nand U16147 (N_16147,N_12783,N_13929);
nand U16148 (N_16148,N_10392,N_13356);
xor U16149 (N_16149,N_14305,N_12480);
nand U16150 (N_16150,N_11164,N_11113);
nand U16151 (N_16151,N_13084,N_14630);
and U16152 (N_16152,N_12579,N_10467);
and U16153 (N_16153,N_14016,N_14303);
nand U16154 (N_16154,N_12802,N_10287);
nor U16155 (N_16155,N_10067,N_13634);
nand U16156 (N_16156,N_10925,N_11138);
or U16157 (N_16157,N_11259,N_12361);
xor U16158 (N_16158,N_10449,N_13812);
nand U16159 (N_16159,N_14726,N_12511);
nand U16160 (N_16160,N_13239,N_13159);
and U16161 (N_16161,N_13657,N_12161);
and U16162 (N_16162,N_12001,N_10714);
nor U16163 (N_16163,N_10562,N_13301);
or U16164 (N_16164,N_13034,N_12368);
xnor U16165 (N_16165,N_11153,N_12060);
nor U16166 (N_16166,N_11815,N_13131);
or U16167 (N_16167,N_13295,N_10024);
and U16168 (N_16168,N_13504,N_11375);
and U16169 (N_16169,N_10174,N_10152);
and U16170 (N_16170,N_11392,N_12048);
xor U16171 (N_16171,N_14355,N_14241);
nor U16172 (N_16172,N_12262,N_12606);
or U16173 (N_16173,N_11395,N_10579);
and U16174 (N_16174,N_14737,N_11975);
nor U16175 (N_16175,N_11830,N_14218);
nor U16176 (N_16176,N_11647,N_14242);
nor U16177 (N_16177,N_14414,N_13102);
and U16178 (N_16178,N_12833,N_13154);
or U16179 (N_16179,N_11124,N_13733);
or U16180 (N_16180,N_10062,N_11843);
and U16181 (N_16181,N_12595,N_10243);
nand U16182 (N_16182,N_10745,N_14655);
nand U16183 (N_16183,N_12711,N_10169);
nand U16184 (N_16184,N_11173,N_10410);
nor U16185 (N_16185,N_11493,N_12989);
nor U16186 (N_16186,N_13240,N_14473);
and U16187 (N_16187,N_11888,N_11359);
nor U16188 (N_16188,N_10217,N_11842);
nor U16189 (N_16189,N_10987,N_10696);
or U16190 (N_16190,N_13538,N_11297);
nand U16191 (N_16191,N_12710,N_12432);
nor U16192 (N_16192,N_14209,N_14907);
nor U16193 (N_16193,N_10590,N_13593);
and U16194 (N_16194,N_12991,N_14503);
nor U16195 (N_16195,N_12594,N_11045);
nand U16196 (N_16196,N_10990,N_13990);
nor U16197 (N_16197,N_13318,N_14469);
nand U16198 (N_16198,N_13231,N_13015);
nor U16199 (N_16199,N_10201,N_11957);
nand U16200 (N_16200,N_11947,N_14089);
nor U16201 (N_16201,N_11206,N_11371);
nand U16202 (N_16202,N_13063,N_10471);
and U16203 (N_16203,N_11114,N_11642);
and U16204 (N_16204,N_14600,N_10610);
and U16205 (N_16205,N_12739,N_11376);
nor U16206 (N_16206,N_10326,N_14082);
nor U16207 (N_16207,N_14872,N_10079);
or U16208 (N_16208,N_13591,N_13902);
nor U16209 (N_16209,N_13051,N_11409);
nand U16210 (N_16210,N_12727,N_10554);
or U16211 (N_16211,N_10605,N_11859);
nand U16212 (N_16212,N_14181,N_10192);
xor U16213 (N_16213,N_14963,N_14658);
xor U16214 (N_16214,N_14178,N_11500);
or U16215 (N_16215,N_14703,N_14063);
nand U16216 (N_16216,N_10001,N_10214);
nor U16217 (N_16217,N_10332,N_11350);
or U16218 (N_16218,N_12436,N_10155);
and U16219 (N_16219,N_13904,N_14400);
and U16220 (N_16220,N_11672,N_11342);
or U16221 (N_16221,N_12264,N_10377);
and U16222 (N_16222,N_13678,N_13824);
or U16223 (N_16223,N_11229,N_13829);
nand U16224 (N_16224,N_14666,N_14237);
or U16225 (N_16225,N_13641,N_13515);
and U16226 (N_16226,N_10829,N_12761);
nand U16227 (N_16227,N_12828,N_10639);
nor U16228 (N_16228,N_14162,N_13496);
nor U16229 (N_16229,N_10820,N_10365);
nand U16230 (N_16230,N_13738,N_13232);
nor U16231 (N_16231,N_13541,N_10008);
or U16232 (N_16232,N_14865,N_13947);
nand U16233 (N_16233,N_14966,N_13156);
and U16234 (N_16234,N_12108,N_14821);
nand U16235 (N_16235,N_14109,N_11080);
and U16236 (N_16236,N_12721,N_13794);
nor U16237 (N_16237,N_13086,N_12952);
and U16238 (N_16238,N_11810,N_12735);
or U16239 (N_16239,N_14514,N_14729);
or U16240 (N_16240,N_14785,N_10415);
or U16241 (N_16241,N_14467,N_13587);
or U16242 (N_16242,N_10493,N_12023);
nor U16243 (N_16243,N_11619,N_12263);
or U16244 (N_16244,N_12458,N_10824);
or U16245 (N_16245,N_11540,N_14998);
nor U16246 (N_16246,N_13899,N_10224);
nor U16247 (N_16247,N_14360,N_11827);
or U16248 (N_16248,N_14490,N_12676);
and U16249 (N_16249,N_10757,N_14862);
nor U16250 (N_16250,N_10039,N_12251);
or U16251 (N_16251,N_13906,N_12841);
nand U16252 (N_16252,N_11535,N_11245);
nand U16253 (N_16253,N_14594,N_10491);
or U16254 (N_16254,N_10601,N_10766);
and U16255 (N_16255,N_14153,N_13452);
and U16256 (N_16256,N_12164,N_10981);
nand U16257 (N_16257,N_14512,N_10483);
and U16258 (N_16258,N_13468,N_13388);
nand U16259 (N_16259,N_11819,N_14554);
nor U16260 (N_16260,N_12972,N_10318);
and U16261 (N_16261,N_11035,N_11593);
and U16262 (N_16262,N_13838,N_11668);
nor U16263 (N_16263,N_14390,N_13921);
nand U16264 (N_16264,N_11447,N_14286);
nor U16265 (N_16265,N_13585,N_14984);
nand U16266 (N_16266,N_13837,N_10831);
and U16267 (N_16267,N_12931,N_14191);
nor U16268 (N_16268,N_14541,N_12506);
or U16269 (N_16269,N_10291,N_10747);
nand U16270 (N_16270,N_10450,N_11689);
or U16271 (N_16271,N_14061,N_11736);
or U16272 (N_16272,N_14150,N_13004);
nor U16273 (N_16273,N_10922,N_14636);
nor U16274 (N_16274,N_11664,N_11690);
nor U16275 (N_16275,N_10930,N_10010);
nor U16276 (N_16276,N_10752,N_14868);
and U16277 (N_16277,N_10703,N_14331);
and U16278 (N_16278,N_11706,N_14995);
nand U16279 (N_16279,N_13348,N_13971);
nor U16280 (N_16280,N_12725,N_13335);
nand U16281 (N_16281,N_12723,N_12453);
nand U16282 (N_16282,N_13376,N_12142);
nor U16283 (N_16283,N_12124,N_14344);
and U16284 (N_16284,N_14679,N_11195);
and U16285 (N_16285,N_11027,N_12507);
nor U16286 (N_16286,N_13107,N_10670);
nor U16287 (N_16287,N_10975,N_11298);
nand U16288 (N_16288,N_11640,N_11861);
nor U16289 (N_16289,N_11352,N_14515);
nand U16290 (N_16290,N_13891,N_14053);
nor U16291 (N_16291,N_12299,N_13145);
nor U16292 (N_16292,N_14387,N_10557);
nor U16293 (N_16293,N_10805,N_14747);
or U16294 (N_16294,N_11483,N_12455);
or U16295 (N_16295,N_13338,N_11836);
or U16296 (N_16296,N_10795,N_11091);
or U16297 (N_16297,N_13633,N_12970);
or U16298 (N_16298,N_11290,N_10606);
nor U16299 (N_16299,N_14629,N_10734);
nand U16300 (N_16300,N_12963,N_12417);
and U16301 (N_16301,N_10409,N_12293);
nand U16302 (N_16302,N_11319,N_12383);
and U16303 (N_16303,N_10753,N_10614);
nor U16304 (N_16304,N_11006,N_10367);
nand U16305 (N_16305,N_10443,N_12069);
nand U16306 (N_16306,N_14952,N_11380);
and U16307 (N_16307,N_13705,N_12188);
nand U16308 (N_16308,N_13970,N_14372);
and U16309 (N_16309,N_13221,N_13277);
and U16310 (N_16310,N_13920,N_10971);
and U16311 (N_16311,N_10113,N_11057);
and U16312 (N_16312,N_12541,N_14522);
or U16313 (N_16313,N_14621,N_14580);
nor U16314 (N_16314,N_13544,N_13353);
nand U16315 (N_16315,N_14294,N_14452);
nand U16316 (N_16316,N_14483,N_10958);
or U16317 (N_16317,N_10303,N_11111);
nand U16318 (N_16318,N_11449,N_12628);
or U16319 (N_16319,N_11561,N_12352);
and U16320 (N_16320,N_14982,N_12338);
or U16321 (N_16321,N_11594,N_12521);
nor U16322 (N_16322,N_13093,N_11053);
and U16323 (N_16323,N_14358,N_10122);
or U16324 (N_16324,N_12904,N_10051);
and U16325 (N_16325,N_11518,N_10701);
and U16326 (N_16326,N_14899,N_13257);
xnor U16327 (N_16327,N_10978,N_12890);
or U16328 (N_16328,N_12708,N_13089);
or U16329 (N_16329,N_12774,N_13704);
nor U16330 (N_16330,N_11335,N_13077);
nor U16331 (N_16331,N_13153,N_14608);
nor U16332 (N_16332,N_12233,N_11159);
and U16333 (N_16333,N_11484,N_12961);
and U16334 (N_16334,N_11343,N_13867);
or U16335 (N_16335,N_11940,N_11943);
and U16336 (N_16336,N_12460,N_12250);
or U16337 (N_16337,N_14171,N_11662);
nand U16338 (N_16338,N_12143,N_13203);
nor U16339 (N_16339,N_10857,N_11774);
and U16340 (N_16340,N_11937,N_14122);
nand U16341 (N_16341,N_14439,N_11824);
or U16342 (N_16342,N_10676,N_14314);
nand U16343 (N_16343,N_11292,N_10528);
nand U16344 (N_16344,N_13877,N_14103);
or U16345 (N_16345,N_13801,N_10496);
nand U16346 (N_16346,N_11431,N_13797);
nor U16347 (N_16347,N_13407,N_10982);
and U16348 (N_16348,N_14045,N_10544);
and U16349 (N_16349,N_12994,N_12379);
or U16350 (N_16350,N_12100,N_10660);
nor U16351 (N_16351,N_13434,N_11150);
or U16352 (N_16352,N_10616,N_12437);
and U16353 (N_16353,N_14377,N_13700);
nor U16354 (N_16354,N_14662,N_10619);
nand U16355 (N_16355,N_10076,N_12672);
and U16356 (N_16356,N_11981,N_14558);
nand U16357 (N_16357,N_11863,N_14460);
and U16358 (N_16358,N_11538,N_11466);
and U16359 (N_16359,N_10892,N_12539);
nor U16360 (N_16360,N_10615,N_14578);
or U16361 (N_16361,N_11272,N_10099);
and U16362 (N_16362,N_12106,N_12254);
or U16363 (N_16363,N_11184,N_13068);
nand U16364 (N_16364,N_10732,N_11818);
nand U16365 (N_16365,N_10274,N_14280);
nor U16366 (N_16366,N_14493,N_13730);
and U16367 (N_16367,N_10058,N_13645);
nor U16368 (N_16368,N_14691,N_10048);
and U16369 (N_16369,N_12448,N_10949);
or U16370 (N_16370,N_10059,N_13573);
nand U16371 (N_16371,N_12895,N_13173);
and U16372 (N_16372,N_14479,N_14461);
nand U16373 (N_16373,N_14302,N_12029);
nor U16374 (N_16374,N_10589,N_10673);
nand U16375 (N_16375,N_14051,N_10427);
nand U16376 (N_16376,N_12940,N_13583);
or U16377 (N_16377,N_11807,N_10529);
or U16378 (N_16378,N_14881,N_14385);
nand U16379 (N_16379,N_13998,N_13934);
and U16380 (N_16380,N_14253,N_10162);
and U16381 (N_16381,N_10447,N_10004);
nor U16382 (N_16382,N_14735,N_14121);
nand U16383 (N_16383,N_10041,N_11638);
nand U16384 (N_16384,N_12066,N_13146);
nor U16385 (N_16385,N_13263,N_12856);
nand U16386 (N_16386,N_11526,N_12839);
and U16387 (N_16387,N_11634,N_11312);
or U16388 (N_16388,N_13138,N_10095);
xnor U16389 (N_16389,N_12027,N_10275);
nor U16390 (N_16390,N_11945,N_13922);
nor U16391 (N_16391,N_14203,N_10886);
xor U16392 (N_16392,N_14757,N_10740);
or U16393 (N_16393,N_13329,N_12358);
or U16394 (N_16394,N_12201,N_14289);
and U16395 (N_16395,N_12572,N_12705);
nor U16396 (N_16396,N_10664,N_12367);
nand U16397 (N_16397,N_14350,N_14625);
nor U16398 (N_16398,N_13636,N_14683);
nand U16399 (N_16399,N_11713,N_13827);
nor U16400 (N_16400,N_11688,N_13849);
nand U16401 (N_16401,N_12374,N_12274);
or U16402 (N_16402,N_11513,N_13000);
or U16403 (N_16403,N_14107,N_13184);
nor U16404 (N_16404,N_14431,N_10166);
and U16405 (N_16405,N_10523,N_11489);
or U16406 (N_16406,N_13516,N_14263);
or U16407 (N_16407,N_13226,N_13716);
nor U16408 (N_16408,N_13248,N_14972);
or U16409 (N_16409,N_13119,N_13297);
or U16410 (N_16410,N_12532,N_14769);
and U16411 (N_16411,N_10568,N_11367);
and U16412 (N_16412,N_13786,N_10060);
or U16413 (N_16413,N_11832,N_14442);
nor U16414 (N_16414,N_10363,N_10329);
and U16415 (N_16415,N_12194,N_11199);
nand U16416 (N_16416,N_13949,N_14989);
nor U16417 (N_16417,N_12642,N_11919);
and U16418 (N_16418,N_13175,N_11993);
and U16419 (N_16419,N_13885,N_12771);
and U16420 (N_16420,N_10094,N_14627);
nand U16421 (N_16421,N_11306,N_13756);
or U16422 (N_16422,N_14151,N_12257);
or U16423 (N_16423,N_11574,N_11135);
and U16424 (N_16424,N_12004,N_14846);
or U16425 (N_16425,N_11980,N_11037);
or U16426 (N_16426,N_13425,N_10385);
or U16427 (N_16427,N_12615,N_12386);
nand U16428 (N_16428,N_12549,N_14285);
and U16429 (N_16429,N_13053,N_11419);
or U16430 (N_16430,N_11207,N_14152);
nor U16431 (N_16431,N_13977,N_13469);
nand U16432 (N_16432,N_14476,N_11425);
or U16433 (N_16433,N_13341,N_10382);
nand U16434 (N_16434,N_12754,N_10693);
nand U16435 (N_16435,N_12957,N_10117);
nand U16436 (N_16436,N_11811,N_13702);
and U16437 (N_16437,N_12463,N_10091);
or U16438 (N_16438,N_12473,N_13714);
or U16439 (N_16439,N_11577,N_14494);
nand U16440 (N_16440,N_10531,N_11741);
nand U16441 (N_16441,N_12399,N_12551);
nand U16442 (N_16442,N_11989,N_13152);
or U16443 (N_16443,N_13289,N_12223);
nor U16444 (N_16444,N_13782,N_14513);
or U16445 (N_16445,N_13305,N_13655);
nand U16446 (N_16446,N_14146,N_11632);
or U16447 (N_16447,N_11628,N_12909);
nor U16448 (N_16448,N_12901,N_13409);
and U16449 (N_16449,N_14238,N_12619);
or U16450 (N_16450,N_14038,N_14304);
and U16451 (N_16451,N_11974,N_13400);
or U16452 (N_16452,N_14613,N_10560);
nand U16453 (N_16453,N_13440,N_14999);
xor U16454 (N_16454,N_10842,N_13941);
nand U16455 (N_16455,N_12704,N_14361);
or U16456 (N_16456,N_13098,N_13320);
and U16457 (N_16457,N_13273,N_12260);
and U16458 (N_16458,N_11062,N_13772);
nand U16459 (N_16459,N_14674,N_12042);
nand U16460 (N_16460,N_13607,N_10314);
or U16461 (N_16461,N_14694,N_10311);
nor U16462 (N_16462,N_11288,N_14800);
or U16463 (N_16463,N_11705,N_11969);
nand U16464 (N_16464,N_10406,N_12195);
nor U16465 (N_16465,N_14913,N_11314);
or U16466 (N_16466,N_11208,N_13377);
and U16467 (N_16467,N_12123,N_14509);
nand U16468 (N_16468,N_10726,N_10627);
or U16469 (N_16469,N_13846,N_12868);
nand U16470 (N_16470,N_11773,N_14816);
and U16471 (N_16471,N_14857,N_14836);
and U16472 (N_16472,N_12709,N_10514);
nand U16473 (N_16473,N_12608,N_10116);
nor U16474 (N_16474,N_11401,N_11915);
or U16475 (N_16475,N_13461,N_11390);
nor U16476 (N_16476,N_10030,N_10029);
and U16477 (N_16477,N_12872,N_13168);
nand U16478 (N_16478,N_10464,N_12191);
or U16479 (N_16479,N_10315,N_11950);
nand U16480 (N_16480,N_10668,N_14764);
nor U16481 (N_16481,N_10055,N_14950);
nor U16482 (N_16482,N_10379,N_14900);
nor U16483 (N_16483,N_12129,N_12275);
nor U16484 (N_16484,N_13276,N_13447);
or U16485 (N_16485,N_12116,N_12016);
or U16486 (N_16486,N_11456,N_10976);
nor U16487 (N_16487,N_10509,N_13957);
nor U16488 (N_16488,N_13069,N_11000);
nand U16489 (N_16489,N_14167,N_10290);
and U16490 (N_16490,N_10533,N_14734);
nand U16491 (N_16491,N_10799,N_11649);
nand U16492 (N_16492,N_12832,N_12057);
nor U16493 (N_16493,N_12534,N_13703);
nor U16494 (N_16494,N_14955,N_12136);
nand U16495 (N_16495,N_12715,N_13603);
or U16496 (N_16496,N_14559,N_10238);
nand U16497 (N_16497,N_13553,N_11675);
nor U16498 (N_16498,N_11096,N_13820);
and U16499 (N_16499,N_13065,N_12622);
nor U16500 (N_16500,N_11878,N_12636);
and U16501 (N_16501,N_14607,N_11965);
or U16502 (N_16502,N_12055,N_10898);
and U16503 (N_16503,N_12112,N_12760);
and U16504 (N_16504,N_12411,N_12266);
or U16505 (N_16505,N_12764,N_12887);
nand U16506 (N_16506,N_10718,N_10848);
nor U16507 (N_16507,N_14780,N_12578);
nand U16508 (N_16508,N_11163,N_10341);
nand U16509 (N_16509,N_11381,N_14852);
or U16510 (N_16510,N_10437,N_14784);
or U16511 (N_16511,N_12311,N_12514);
nor U16512 (N_16512,N_10588,N_10986);
or U16513 (N_16513,N_11478,N_11047);
or U16514 (N_16514,N_12874,N_12305);
or U16515 (N_16515,N_10604,N_14765);
and U16516 (N_16516,N_10611,N_14832);
nor U16517 (N_16517,N_10179,N_13191);
or U16518 (N_16518,N_11653,N_11648);
nand U16519 (N_16519,N_13394,N_11826);
nor U16520 (N_16520,N_10761,N_11490);
nand U16521 (N_16521,N_14084,N_14472);
nor U16522 (N_16522,N_13182,N_10284);
or U16523 (N_16523,N_14433,N_12364);
nor U16524 (N_16524,N_12145,N_10736);
or U16525 (N_16525,N_11678,N_13908);
and U16526 (N_16526,N_10066,N_13640);
and U16527 (N_16527,N_11812,N_11720);
and U16528 (N_16528,N_13945,N_10387);
xor U16529 (N_16529,N_10725,N_11891);
or U16530 (N_16530,N_10888,N_10054);
nor U16531 (N_16531,N_10459,N_14939);
nand U16532 (N_16532,N_10383,N_14193);
and U16533 (N_16533,N_10215,N_10743);
nand U16534 (N_16534,N_10182,N_12759);
nor U16535 (N_16535,N_10448,N_12614);
and U16536 (N_16536,N_14612,N_13868);
or U16537 (N_16537,N_12693,N_11684);
and U16538 (N_16538,N_10000,N_14001);
and U16539 (N_16539,N_10302,N_13268);
nand U16540 (N_16540,N_13266,N_14054);
or U16541 (N_16541,N_13889,N_11877);
or U16542 (N_16542,N_11428,N_11544);
nand U16543 (N_16543,N_14696,N_10110);
nand U16544 (N_16544,N_10867,N_12003);
nand U16545 (N_16545,N_12620,N_12937);
nand U16546 (N_16546,N_13095,N_14077);
nor U16547 (N_16547,N_10977,N_10645);
nand U16548 (N_16548,N_11060,N_14581);
nor U16549 (N_16549,N_14088,N_11789);
xnor U16550 (N_16550,N_10628,N_14806);
nor U16551 (N_16551,N_14728,N_14032);
and U16552 (N_16552,N_10006,N_10177);
nor U16553 (N_16553,N_10225,N_13985);
or U16554 (N_16554,N_10337,N_14874);
nand U16555 (N_16555,N_14523,N_12034);
or U16556 (N_16556,N_12287,N_12813);
nor U16557 (N_16557,N_11323,N_14654);
nand U16558 (N_16558,N_13559,N_10384);
nor U16559 (N_16559,N_12400,N_10137);
nand U16560 (N_16560,N_14102,N_11410);
nand U16561 (N_16561,N_14685,N_10210);
nor U16562 (N_16562,N_11912,N_10078);
nand U16563 (N_16563,N_12847,N_11504);
nor U16564 (N_16564,N_12893,N_11024);
and U16565 (N_16565,N_13044,N_14492);
or U16566 (N_16566,N_12990,N_11271);
and U16567 (N_16567,N_11956,N_13764);
and U16568 (N_16568,N_11984,N_11902);
nand U16569 (N_16569,N_10715,N_10536);
or U16570 (N_16570,N_10357,N_11911);
nor U16571 (N_16571,N_12602,N_10395);
nand U16572 (N_16572,N_11463,N_13789);
nor U16573 (N_16573,N_12403,N_14597);
and U16574 (N_16574,N_14368,N_14850);
and U16575 (N_16575,N_13907,N_13076);
nand U16576 (N_16576,N_13913,N_11411);
nand U16577 (N_16577,N_12081,N_11107);
and U16578 (N_16578,N_12092,N_12147);
or U16579 (N_16579,N_13872,N_14234);
nor U16580 (N_16580,N_13120,N_14282);
and U16581 (N_16581,N_10875,N_10129);
and U16582 (N_16582,N_10960,N_13328);
nand U16583 (N_16583,N_14006,N_14293);
nor U16584 (N_16584,N_12558,N_14300);
nor U16585 (N_16585,N_11445,N_14709);
and U16586 (N_16586,N_10164,N_13781);
or U16587 (N_16587,N_14505,N_11336);
nand U16588 (N_16588,N_14017,N_10741);
nand U16589 (N_16589,N_10220,N_12537);
nor U16590 (N_16590,N_12756,N_11155);
nand U16591 (N_16591,N_14619,N_13048);
nor U16592 (N_16592,N_11151,N_13973);
nand U16593 (N_16593,N_13014,N_14225);
and U16594 (N_16594,N_13744,N_10320);
and U16595 (N_16595,N_12019,N_11978);
nand U16596 (N_16596,N_12907,N_12103);
or U16597 (N_16597,N_11567,N_12378);
and U16598 (N_16598,N_14186,N_12085);
nor U16599 (N_16599,N_13768,N_14744);
and U16600 (N_16600,N_12292,N_12938);
nor U16601 (N_16601,N_11304,N_13687);
or U16602 (N_16602,N_14544,N_13420);
nand U16603 (N_16603,N_12324,N_10970);
or U16604 (N_16604,N_12714,N_12139);
nor U16605 (N_16605,N_11751,N_12958);
or U16606 (N_16606,N_12294,N_14276);
and U16607 (N_16607,N_12241,N_12651);
nor U16608 (N_16608,N_13450,N_12217);
and U16609 (N_16609,N_13752,N_12495);
nor U16610 (N_16610,N_12822,N_13628);
nor U16611 (N_16611,N_14391,N_14495);
and U16612 (N_16612,N_11181,N_12026);
nor U16613 (N_16613,N_13293,N_13410);
and U16614 (N_16614,N_11120,N_10127);
nor U16615 (N_16615,N_12282,N_10084);
nand U16616 (N_16616,N_13380,N_12528);
nor U16617 (N_16617,N_11719,N_10635);
nor U16618 (N_16618,N_13841,N_14671);
nor U16619 (N_16619,N_13563,N_12670);
nand U16620 (N_16620,N_14732,N_12967);
or U16621 (N_16621,N_11139,N_11453);
nor U16622 (N_16622,N_12258,N_13178);
nor U16623 (N_16623,N_11049,N_10564);
and U16624 (N_16624,N_10046,N_13834);
nor U16625 (N_16625,N_14849,N_13582);
and U16626 (N_16626,N_11287,N_12245);
and U16627 (N_16627,N_12569,N_11115);
nor U16628 (N_16628,N_11255,N_10852);
nor U16629 (N_16629,N_10651,N_14312);
nor U16630 (N_16630,N_10524,N_11404);
nor U16631 (N_16631,N_13307,N_12007);
and U16632 (N_16632,N_14529,N_14817);
nor U16633 (N_16633,N_14379,N_10625);
and U16634 (N_16634,N_11817,N_13896);
or U16635 (N_16635,N_14297,N_12666);
nor U16636 (N_16636,N_12474,N_11707);
or U16637 (N_16637,N_13209,N_13984);
nor U16638 (N_16638,N_10617,N_11734);
nand U16639 (N_16639,N_14180,N_10818);
nand U16640 (N_16640,N_14093,N_11948);
or U16641 (N_16641,N_13311,N_12898);
and U16642 (N_16642,N_14448,N_10874);
and U16643 (N_16643,N_12225,N_10526);
nor U16644 (N_16644,N_12911,N_13431);
or U16645 (N_16645,N_10063,N_10510);
nor U16646 (N_16646,N_10267,N_11233);
nor U16647 (N_16647,N_12187,N_11608);
nand U16648 (N_16648,N_12736,N_14434);
or U16649 (N_16649,N_12933,N_11056);
and U16650 (N_16650,N_14392,N_12939);
nand U16651 (N_16651,N_11763,N_13939);
or U16652 (N_16652,N_13875,N_12951);
nand U16653 (N_16653,N_10582,N_10999);
or U16654 (N_16654,N_13976,N_12853);
nor U16655 (N_16655,N_11868,N_11579);
nand U16656 (N_16656,N_14270,N_14185);
and U16657 (N_16657,N_11757,N_14652);
or U16658 (N_16658,N_13887,N_13600);
and U16659 (N_16659,N_10486,N_10985);
nand U16660 (N_16660,N_10662,N_13198);
or U16661 (N_16661,N_10053,N_14052);
nand U16662 (N_16662,N_10380,N_10657);
nand U16663 (N_16663,N_11451,N_10585);
and U16664 (N_16664,N_12810,N_10105);
nor U16665 (N_16665,N_10350,N_11933);
and U16666 (N_16666,N_14320,N_14101);
or U16667 (N_16667,N_11660,N_13792);
or U16668 (N_16668,N_12744,N_14155);
nor U16669 (N_16669,N_13962,N_13586);
and U16670 (N_16670,N_11073,N_14428);
nor U16671 (N_16671,N_12526,N_13832);
nand U16672 (N_16672,N_11560,N_12137);
or U16673 (N_16673,N_11726,N_12664);
and U16674 (N_16674,N_12962,N_14420);
and U16675 (N_16675,N_11977,N_14922);
nor U16676 (N_16676,N_11716,N_13067);
and U16677 (N_16677,N_14889,N_12149);
and U16678 (N_16678,N_13373,N_10451);
or U16679 (N_16679,N_14019,N_14546);
and U16680 (N_16680,N_10924,N_14547);
nor U16681 (N_16681,N_13271,N_10697);
or U16682 (N_16682,N_12596,N_14359);
and U16683 (N_16683,N_10918,N_11935);
or U16684 (N_16684,N_14539,N_10197);
nand U16685 (N_16685,N_14521,N_13176);
or U16686 (N_16686,N_11523,N_11250);
and U16687 (N_16687,N_12179,N_13136);
or U16688 (N_16688,N_13596,N_12435);
and U16689 (N_16689,N_11200,N_12959);
nor U16690 (N_16690,N_10391,N_11285);
nand U16691 (N_16691,N_11042,N_11334);
and U16692 (N_16692,N_11607,N_14682);
or U16693 (N_16693,N_14901,N_12377);
and U16694 (N_16694,N_11020,N_10200);
nor U16695 (N_16695,N_11783,N_11251);
and U16696 (N_16696,N_10027,N_12926);
or U16697 (N_16697,N_10269,N_11988);
nand U16698 (N_16698,N_11749,N_14481);
nor U16699 (N_16699,N_11918,N_14318);
nand U16700 (N_16700,N_14252,N_12669);
or U16701 (N_16701,N_10802,N_10807);
nor U16702 (N_16702,N_13799,N_13524);
nor U16703 (N_16703,N_14357,N_13472);
nand U16704 (N_16704,N_11480,N_14858);
and U16705 (N_16705,N_10744,N_12542);
nand U16706 (N_16706,N_10333,N_13316);
and U16707 (N_16707,N_13489,N_11722);
nor U16708 (N_16708,N_10253,N_13520);
nand U16709 (N_16709,N_11129,N_10049);
or U16710 (N_16710,N_10317,N_11889);
and U16711 (N_16711,N_10576,N_14177);
and U16712 (N_16712,N_11354,N_14602);
nor U16713 (N_16713,N_10040,N_14370);
nor U16714 (N_16714,N_12365,N_13932);
and U16715 (N_16715,N_10862,N_11149);
nor U16716 (N_16716,N_13078,N_14502);
nand U16717 (N_16717,N_12166,N_14823);
and U16718 (N_16718,N_14796,N_10932);
or U16719 (N_16719,N_12226,N_13850);
nor U16720 (N_16720,N_14997,N_11441);
or U16721 (N_16721,N_11973,N_14065);
or U16722 (N_16722,N_13334,N_10887);
or U16723 (N_16723,N_10735,N_11187);
and U16724 (N_16724,N_10259,N_10613);
nand U16725 (N_16725,N_12908,N_14258);
and U16726 (N_16726,N_13543,N_14928);
or U16727 (N_16727,N_12444,N_10584);
and U16728 (N_16728,N_13217,N_11686);
nor U16729 (N_16729,N_12028,N_11235);
and U16730 (N_16730,N_11680,N_14960);
nand U16731 (N_16731,N_14418,N_14339);
or U16732 (N_16732,N_13064,N_10344);
nor U16733 (N_16733,N_13445,N_10178);
and U16734 (N_16734,N_14569,N_14873);
nor U16735 (N_16735,N_13721,N_10282);
or U16736 (N_16736,N_10778,N_14184);
and U16737 (N_16737,N_12597,N_11758);
and U16738 (N_16738,N_14374,N_11753);
nand U16739 (N_16739,N_11472,N_11534);
and U16740 (N_16740,N_10998,N_12790);
xor U16741 (N_16741,N_11081,N_12355);
nor U16742 (N_16742,N_12560,N_10602);
nor U16743 (N_16743,N_14404,N_10393);
nand U16744 (N_16744,N_10148,N_13128);
and U16745 (N_16745,N_11021,N_10219);
nor U16746 (N_16746,N_13357,N_10124);
or U16747 (N_16747,N_11611,N_12801);
nand U16748 (N_16748,N_11477,N_13610);
or U16749 (N_16749,N_12621,N_10397);
or U16750 (N_16750,N_14048,N_10366);
and U16751 (N_16751,N_12679,N_13719);
nor U16752 (N_16752,N_12064,N_14875);
nor U16753 (N_16753,N_12943,N_12781);
nor U16754 (N_16754,N_14969,N_12461);
nand U16755 (N_16755,N_11406,N_11134);
or U16756 (N_16756,N_14525,N_13424);
or U16757 (N_16757,N_14985,N_11067);
nand U16758 (N_16758,N_13158,N_13983);
or U16759 (N_16759,N_14435,N_14205);
or U16760 (N_16760,N_10358,N_12879);
nor U16761 (N_16761,N_12722,N_11063);
nand U16762 (N_16762,N_13169,N_12575);
and U16763 (N_16763,N_11031,N_14386);
nor U16764 (N_16764,N_11434,N_10102);
nand U16765 (N_16765,N_13467,N_11028);
nor U16766 (N_16766,N_14693,N_11074);
or U16767 (N_16767,N_10273,N_10120);
or U16768 (N_16768,N_14413,N_14246);
and U16769 (N_16769,N_13914,N_13893);
and U16770 (N_16770,N_11030,N_14591);
xnor U16771 (N_16771,N_12570,N_14081);
nor U16772 (N_16772,N_11656,N_12198);
nand U16773 (N_16773,N_13525,N_13677);
and U16774 (N_16774,N_13762,N_10167);
nand U16775 (N_16775,N_12798,N_12863);
and U16776 (N_16776,N_11711,N_11767);
or U16777 (N_16777,N_14902,N_14450);
nand U16778 (N_16778,N_13033,N_14916);
or U16779 (N_16779,N_11721,N_10729);
nand U16780 (N_16780,N_10460,N_10661);
nor U16781 (N_16781,N_13796,N_12130);
or U16782 (N_16782,N_12949,N_11582);
xor U16783 (N_16783,N_13658,N_11473);
nand U16784 (N_16784,N_12431,N_10212);
or U16785 (N_16785,N_12880,N_11921);
nor U16786 (N_16786,N_12659,N_10319);
nand U16787 (N_16787,N_10368,N_11677);
nor U16788 (N_16788,N_11310,N_10112);
nand U16789 (N_16789,N_14011,N_12751);
nor U16790 (N_16790,N_14283,N_11923);
or U16791 (N_16791,N_13927,N_11101);
nand U16792 (N_16792,N_11942,N_14981);
and U16793 (N_16793,N_11873,N_12820);
or U16794 (N_16794,N_13643,N_13608);
nor U16795 (N_16795,N_10252,N_14112);
nor U16796 (N_16796,N_11814,N_13100);
xnor U16797 (N_16797,N_10682,N_14519);
or U16798 (N_16798,N_13336,N_12424);
nor U16799 (N_16799,N_11944,N_11731);
xnor U16800 (N_16800,N_13879,N_14941);
or U16801 (N_16801,N_14990,N_12021);
or U16802 (N_16802,N_13466,N_10133);
nand U16803 (N_16803,N_12101,N_13897);
nand U16804 (N_16804,N_13393,N_11737);
nor U16805 (N_16805,N_12087,N_13815);
or U16806 (N_16806,N_14730,N_11078);
or U16807 (N_16807,N_13747,N_12273);
nor U16808 (N_16808,N_13728,N_14934);
and U16809 (N_16809,N_14617,N_10973);
nor U16810 (N_16810,N_10952,N_11655);
nand U16811 (N_16811,N_10417,N_10013);
nand U16812 (N_16812,N_12283,N_14190);
nor U16813 (N_16813,N_14640,N_11239);
nand U16814 (N_16814,N_11557,N_11443);
and U16815 (N_16815,N_13613,N_10111);
nand U16816 (N_16816,N_12284,N_10598);
or U16817 (N_16817,N_12259,N_13379);
nand U16818 (N_16818,N_14389,N_11143);
and U16819 (N_16819,N_13707,N_13805);
and U16820 (N_16820,N_10724,N_12485);
and U16821 (N_16821,N_12171,N_13533);
and U16822 (N_16822,N_13760,N_12855);
nand U16823 (N_16823,N_11457,N_14740);
or U16824 (N_16824,N_11699,N_11624);
nor U16825 (N_16825,N_12500,N_11869);
nor U16826 (N_16826,N_11808,N_11227);
or U16827 (N_16827,N_12421,N_11126);
nor U16828 (N_16828,N_10768,N_12434);
nand U16829 (N_16829,N_11300,N_13080);
nand U16830 (N_16830,N_11946,N_10876);
nand U16831 (N_16831,N_10943,N_12457);
xor U16832 (N_16832,N_12337,N_13106);
nor U16833 (N_16833,N_13988,N_11588);
nand U16834 (N_16834,N_10185,N_11228);
and U16835 (N_16835,N_14292,N_11177);
or U16836 (N_16836,N_10136,N_11929);
nor U16837 (N_16837,N_11284,N_11424);
or U16838 (N_16838,N_14894,N_14207);
nand U16839 (N_16839,N_12583,N_14248);
nand U16840 (N_16840,N_14254,N_10767);
xnor U16841 (N_16841,N_12914,N_12242);
or U16842 (N_16842,N_10926,N_10034);
and U16843 (N_16843,N_11525,N_10074);
nor U16844 (N_16844,N_11183,N_14677);
nand U16845 (N_16845,N_12803,N_13310);
nor U16846 (N_16846,N_13360,N_14599);
nand U16847 (N_16847,N_13349,N_14175);
nand U16848 (N_16848,N_10505,N_10378);
and U16849 (N_16849,N_12848,N_13454);
nand U16850 (N_16850,N_10748,N_10226);
nor U16851 (N_16851,N_11584,N_13663);
or U16852 (N_16852,N_12823,N_13383);
nand U16853 (N_16853,N_14542,N_13638);
nor U16854 (N_16854,N_11681,N_14968);
nand U16855 (N_16855,N_13580,N_11370);
nor U16856 (N_16856,N_14745,N_10965);
nand U16857 (N_16857,N_14672,N_11908);
or U16858 (N_16858,N_10597,N_12978);
nor U16859 (N_16859,N_12674,N_11620);
and U16860 (N_16860,N_11276,N_13278);
nor U16861 (N_16861,N_11119,N_13836);
nor U16862 (N_16862,N_10538,N_14216);
and U16863 (N_16863,N_11382,N_11666);
nand U16864 (N_16864,N_14068,N_11786);
nor U16865 (N_16865,N_14334,N_14215);
or U16866 (N_16866,N_12035,N_14208);
or U16867 (N_16867,N_13926,N_13302);
and U16868 (N_16868,N_10222,N_10050);
nor U16869 (N_16869,N_11510,N_13179);
or U16870 (N_16870,N_14707,N_10482);
or U16871 (N_16871,N_10375,N_10476);
nand U16872 (N_16872,N_10941,N_12859);
or U16873 (N_16873,N_11754,N_10089);
or U16874 (N_16874,N_12427,N_11527);
nand U16875 (N_16875,N_12797,N_12272);
nand U16876 (N_16876,N_13898,N_10340);
nand U16877 (N_16877,N_11627,N_11044);
and U16878 (N_16878,N_13272,N_11442);
nor U16879 (N_16879,N_10936,N_12618);
nor U16880 (N_16880,N_12439,N_12546);
or U16881 (N_16881,N_11795,N_13367);
and U16882 (N_16882,N_14409,N_13750);
or U16883 (N_16883,N_12643,N_10543);
nor U16884 (N_16884,N_10839,N_12211);
nand U16885 (N_16885,N_13274,N_13142);
nor U16886 (N_16886,N_12784,N_14930);
or U16887 (N_16887,N_14313,N_10720);
nand U16888 (N_16888,N_10821,N_11629);
and U16889 (N_16889,N_13860,N_13755);
nor U16890 (N_16890,N_13475,N_12519);
and U16891 (N_16891,N_12440,N_13326);
and U16892 (N_16892,N_11501,N_11670);
or U16893 (N_16893,N_14606,N_11283);
nor U16894 (N_16894,N_14498,N_12508);
nor U16895 (N_16895,N_14154,N_10508);
and U16896 (N_16896,N_11280,N_14983);
and U16897 (N_16897,N_12039,N_12645);
and U16898 (N_16898,N_13319,N_14343);
and U16899 (N_16899,N_13589,N_12544);
nand U16900 (N_16900,N_13864,N_10463);
or U16901 (N_16901,N_14098,N_13370);
and U16902 (N_16902,N_14035,N_12576);
nand U16903 (N_16903,N_11240,N_11379);
nand U16904 (N_16904,N_14430,N_13930);
and U16905 (N_16905,N_11128,N_13667);
or U16906 (N_16906,N_13192,N_13754);
and U16907 (N_16907,N_10644,N_11932);
nand U16908 (N_16908,N_11486,N_12699);
or U16909 (N_16909,N_10665,N_14708);
or U16910 (N_16910,N_13552,N_11883);
nor U16911 (N_16911,N_14973,N_13492);
xor U16912 (N_16912,N_14953,N_12503);
nand U16913 (N_16913,N_10068,N_11316);
nand U16914 (N_16914,N_12684,N_10908);
nand U16915 (N_16915,N_11555,N_10513);
and U16916 (N_16916,N_10181,N_14165);
nor U16917 (N_16917,N_14555,N_12854);
or U16918 (N_16918,N_14417,N_14543);
or U16919 (N_16919,N_13306,N_14716);
nor U16920 (N_16920,N_12357,N_13233);
nand U16921 (N_16921,N_10195,N_14689);
nand U16922 (N_16922,N_10321,N_11747);
nor U16923 (N_16923,N_13712,N_10190);
nor U16924 (N_16924,N_10352,N_10705);
and U16925 (N_16925,N_11469,N_14419);
nand U16926 (N_16926,N_11748,N_11673);
nor U16927 (N_16927,N_10707,N_14779);
or U16928 (N_16928,N_12296,N_11630);
and U16929 (N_16929,N_14751,N_10873);
and U16930 (N_16930,N_12974,N_12748);
or U16931 (N_16931,N_10028,N_12627);
nand U16932 (N_16932,N_11236,N_10142);
and U16933 (N_16933,N_12892,N_11209);
nand U16934 (N_16934,N_10240,N_13253);
nand U16935 (N_16935,N_12144,N_12229);
nand U16936 (N_16936,N_13125,N_12325);
or U16937 (N_16937,N_13457,N_12562);
or U16938 (N_16938,N_11590,N_12732);
nor U16939 (N_16939,N_10546,N_13401);
or U16940 (N_16940,N_13476,N_12531);
nand U16941 (N_16941,N_13021,N_14743);
nor U16942 (N_16942,N_14247,N_11275);
xor U16943 (N_16943,N_11265,N_10485);
nand U16944 (N_16944,N_12215,N_10419);
or U16945 (N_16945,N_13748,N_14408);
nand U16946 (N_16946,N_13375,N_11531);
or U16947 (N_16947,N_11348,N_14911);
and U16948 (N_16948,N_11586,N_11599);
nor U16949 (N_16949,N_14277,N_11194);
nand U16950 (N_16950,N_13118,N_10405);
xor U16951 (N_16951,N_10573,N_11700);
nand U16952 (N_16952,N_10257,N_10834);
and U16953 (N_16953,N_12212,N_10763);
nor U16954 (N_16954,N_13673,N_10993);
and U16955 (N_16955,N_12392,N_12717);
xnor U16956 (N_16956,N_12146,N_14792);
nor U16957 (N_16957,N_13285,N_12220);
nor U16958 (N_16958,N_11787,N_13193);
xor U16959 (N_16959,N_13135,N_11417);
or U16960 (N_16960,N_14021,N_11393);
nor U16961 (N_16961,N_14713,N_11530);
nand U16962 (N_16962,N_10762,N_14298);
nor U16963 (N_16963,N_12270,N_11176);
or U16964 (N_16964,N_12168,N_12512);
nand U16965 (N_16965,N_11373,N_12462);
nand U16966 (N_16966,N_11145,N_10327);
and U16967 (N_16967,N_11641,N_13132);
and U16968 (N_16968,N_10128,N_11182);
or U16969 (N_16969,N_14211,N_13486);
or U16970 (N_16970,N_10996,N_10083);
nor U16971 (N_16971,N_14076,N_12836);
or U16972 (N_16972,N_11140,N_10968);
nand U16973 (N_16973,N_10216,N_14310);
nand U16974 (N_16974,N_12059,N_14140);
nor U16975 (N_16975,N_12351,N_11644);
or U16976 (N_16976,N_13148,N_13979);
nor U16977 (N_16977,N_10910,N_13124);
nor U16978 (N_16978,N_14055,N_14454);
or U16979 (N_16979,N_11026,N_11505);
nand U16980 (N_16980,N_12917,N_11427);
or U16981 (N_16981,N_11340,N_14106);
or U16982 (N_16982,N_14168,N_10902);
or U16983 (N_16983,N_14959,N_11604);
and U16984 (N_16984,N_10995,N_12647);
or U16985 (N_16985,N_10176,N_10254);
or U16986 (N_16986,N_12109,N_12181);
nor U16987 (N_16987,N_14724,N_14643);
nor U16988 (N_16988,N_14993,N_13681);
and U16989 (N_16989,N_14189,N_13323);
and U16990 (N_16990,N_12000,N_10804);
and U16991 (N_16991,N_10596,N_10865);
nor U16992 (N_16992,N_10249,N_14876);
nor U16993 (N_16993,N_11188,N_14841);
or U16994 (N_16994,N_10530,N_14143);
or U16995 (N_16995,N_10637,N_10731);
nor U16996 (N_16996,N_10860,N_12588);
nor U16997 (N_16997,N_10138,N_12755);
and U16998 (N_16998,N_13735,N_10309);
and U16999 (N_16999,N_10348,N_12983);
or U17000 (N_17000,N_11580,N_13296);
and U17001 (N_17001,N_10953,N_14170);
nor U17002 (N_17002,N_11755,N_12344);
or U17003 (N_17003,N_12479,N_14520);
or U17004 (N_17004,N_11718,N_14271);
nor U17005 (N_17005,N_10293,N_13332);
and U17006 (N_17006,N_10399,N_11583);
xnor U17007 (N_17007,N_12648,N_10480);
or U17008 (N_17008,N_11347,N_12538);
nand U17009 (N_17009,N_11398,N_14410);
and U17010 (N_17010,N_11146,N_10631);
or U17011 (N_17011,N_12135,N_12815);
and U17012 (N_17012,N_12134,N_14870);
nand U17013 (N_17013,N_13560,N_13140);
nor U17014 (N_17014,N_13225,N_14695);
nand U17015 (N_17015,N_11979,N_10681);
and U17016 (N_17016,N_13362,N_13746);
xnor U17017 (N_17017,N_14879,N_12497);
nor U17018 (N_17018,N_14260,N_10798);
or U17019 (N_17019,N_12214,N_10429);
nor U17020 (N_17020,N_11844,N_13912);
nor U17021 (N_17021,N_10271,N_10750);
xnor U17022 (N_17022,N_10454,N_14956);
nor U17023 (N_17023,N_12017,N_13690);
and U17024 (N_17024,N_14108,N_12009);
or U17025 (N_17025,N_12339,N_14348);
nand U17026 (N_17026,N_12253,N_11023);
nor U17027 (N_17027,N_14837,N_11014);
nand U17028 (N_17028,N_14447,N_10234);
and U17029 (N_17029,N_11792,N_13321);
or U17030 (N_17030,N_14412,N_10331);
nor U17031 (N_17031,N_10815,N_10242);
or U17032 (N_17032,N_14878,N_12807);
nand U17033 (N_17033,N_12486,N_12127);
nor U17034 (N_17034,N_12304,N_10090);
and U17035 (N_17035,N_14834,N_14903);
and U17036 (N_17036,N_11547,N_12730);
and U17037 (N_17037,N_11961,N_14116);
or U17038 (N_17038,N_14871,N_14637);
and U17039 (N_17039,N_11646,N_10646);
nor U17040 (N_17040,N_12025,N_12230);
and U17041 (N_17041,N_11717,N_12667);
nand U17042 (N_17042,N_11470,N_10043);
nand U17043 (N_17043,N_13734,N_13652);
nand U17044 (N_17044,N_10180,N_11829);
and U17045 (N_17045,N_14842,N_12547);
nor U17046 (N_17046,N_14062,N_11459);
or U17047 (N_17047,N_13378,N_11388);
nor U17048 (N_17048,N_14920,N_11141);
nor U17049 (N_17049,N_14596,N_14421);
and U17050 (N_17050,N_11564,N_13413);
nor U17051 (N_17051,N_13333,N_14268);
or U17052 (N_17052,N_10891,N_14669);
and U17053 (N_17053,N_12885,N_10643);
nor U17054 (N_17054,N_12731,N_14987);
nand U17055 (N_17055,N_10921,N_10264);
nand U17056 (N_17056,N_10038,N_14851);
or U17057 (N_17057,N_10343,N_10031);
nor U17058 (N_17058,N_11405,N_13408);
nor U17059 (N_17059,N_13761,N_12632);
nor U17060 (N_17060,N_13938,N_13729);
and U17061 (N_17061,N_14278,N_13042);
nand U17062 (N_17062,N_12749,N_14944);
nor U17063 (N_17063,N_11048,N_12316);
nand U17064 (N_17064,N_14436,N_14923);
nor U17065 (N_17065,N_14274,N_14147);
and U17066 (N_17066,N_13605,N_12785);
nor U17067 (N_17067,N_14632,N_10835);
nand U17068 (N_17068,N_11840,N_13485);
nand U17069 (N_17069,N_13958,N_12812);
nand U17070 (N_17070,N_11362,N_12934);
nand U17071 (N_17071,N_12932,N_10425);
nand U17072 (N_17072,N_14306,N_11784);
and U17073 (N_17073,N_14584,N_14761);
nor U17074 (N_17074,N_10404,N_10445);
nor U17075 (N_17075,N_14949,N_10355);
and U17076 (N_17076,N_13739,N_11733);
nor U17077 (N_17077,N_10897,N_13831);
nand U17078 (N_17078,N_10479,N_14891);
and U17079 (N_17079,N_12184,N_14964);
nand U17080 (N_17080,N_14132,N_10313);
and U17081 (N_17081,N_10621,N_11635);
or U17082 (N_17082,N_14267,N_10507);
or U17083 (N_17083,N_13569,N_11901);
and U17084 (N_17084,N_12899,N_14839);
or U17085 (N_17085,N_11870,N_12065);
and U17086 (N_17086,N_11517,N_14466);
and U17087 (N_17087,N_12286,N_11144);
and U17088 (N_17088,N_12172,N_10263);
nand U17089 (N_17089,N_10989,N_12808);
nand U17090 (N_17090,N_10810,N_13038);
nor U17091 (N_17091,N_12393,N_14975);
and U17092 (N_17092,N_13206,N_13096);
nand U17093 (N_17093,N_12271,N_10555);
and U17094 (N_17094,N_11064,N_10905);
nand U17095 (N_17095,N_10923,N_12753);
or U17096 (N_17096,N_14074,N_12346);
nor U17097 (N_17097,N_10607,N_10044);
nand U17098 (N_17098,N_12805,N_10636);
or U17099 (N_17099,N_11521,N_12208);
or U17100 (N_17100,N_12592,N_13055);
nor U17101 (N_17101,N_13960,N_12814);
or U17102 (N_17102,N_11701,N_10979);
nand U17103 (N_17103,N_11337,N_12876);
nor U17104 (N_17104,N_10515,N_14496);
or U17105 (N_17105,N_11365,N_12982);
nand U17106 (N_17106,N_14887,N_11070);
or U17107 (N_17107,N_14345,N_10859);
or U17108 (N_17108,N_12663,N_10487);
nor U17109 (N_17109,N_10121,N_11847);
and U17110 (N_17110,N_11036,N_12997);
and U17111 (N_17111,N_14090,N_11330);
and U17112 (N_17112,N_12011,N_11566);
nand U17113 (N_17113,N_14718,N_10096);
nor U17114 (N_17114,N_10490,N_10620);
nand U17115 (N_17115,N_12384,N_11471);
nand U17116 (N_17116,N_13556,N_14033);
or U17117 (N_17117,N_11446,N_14482);
nor U17118 (N_17118,N_14194,N_14838);
or U17119 (N_17119,N_13222,N_10209);
nor U17120 (N_17120,N_11972,N_11563);
and U17121 (N_17121,N_13254,N_14092);
nor U17122 (N_17122,N_12535,N_13788);
nand U17123 (N_17123,N_12269,N_10814);
and U17124 (N_17124,N_14110,N_14036);
or U17125 (N_17125,N_13392,N_13978);
nand U17126 (N_17126,N_14853,N_10077);
and U17127 (N_17127,N_12366,N_14333);
nor U17128 (N_17128,N_14325,N_14914);
nor U17129 (N_17129,N_12986,N_12433);
and U17130 (N_17130,N_11241,N_14251);
nor U17131 (N_17131,N_10809,N_14125);
nand U17132 (N_17132,N_13195,N_13919);
nor U17133 (N_17133,N_10235,N_10884);
and U17134 (N_17134,N_10211,N_11872);
or U17135 (N_17135,N_12867,N_13758);
or U17136 (N_17136,N_13713,N_10191);
nor U17137 (N_17137,N_11522,N_10787);
nor U17138 (N_17138,N_11075,N_14163);
or U17139 (N_17139,N_10472,N_13840);
and U17140 (N_17140,N_14080,N_10288);
nor U17141 (N_17141,N_11679,N_10394);
nand U17142 (N_17142,N_14524,N_10684);
or U17143 (N_17143,N_11954,N_14843);
nand U17144 (N_17144,N_10565,N_13355);
and U17145 (N_17145,N_14249,N_13411);
nand U17146 (N_17146,N_10007,N_10712);
nor U17147 (N_17147,N_10432,N_12278);
nand U17148 (N_17148,N_12809,N_14921);
nor U17149 (N_17149,N_10751,N_11568);
and U17150 (N_17150,N_12787,N_11303);
and U17151 (N_17151,N_13959,N_13027);
nand U17152 (N_17152,N_10361,N_11652);
and U17153 (N_17153,N_13071,N_14508);
nor U17154 (N_17154,N_12782,N_12067);
nand U17155 (N_17155,N_12356,N_12120);
nand U17156 (N_17156,N_13126,N_10338);
and U17157 (N_17157,N_14489,N_10446);
nor U17158 (N_17158,N_14319,N_10285);
or U17159 (N_17159,N_10154,N_11959);
and U17160 (N_17160,N_13966,N_14213);
and U17161 (N_17161,N_12903,N_10246);
nand U17162 (N_17162,N_11481,N_13016);
and U17163 (N_17163,N_13110,N_10301);
and U17164 (N_17164,N_11881,N_13861);
nor U17165 (N_17165,N_11387,N_10070);
nor U17166 (N_17166,N_14202,N_14340);
nor U17167 (N_17167,N_10346,N_10575);
nand U17168 (N_17168,N_13317,N_14988);
or U17169 (N_17169,N_11202,N_12420);
nand U17170 (N_17170,N_12882,N_12441);
and U17171 (N_17171,N_14176,N_12190);
and U17172 (N_17172,N_10433,N_12482);
and U17173 (N_17173,N_12342,N_14264);
nand U17174 (N_17174,N_12770,N_14646);
and U17175 (N_17175,N_10109,N_10014);
nor U17176 (N_17176,N_14746,N_14801);
or U17177 (N_17177,N_12586,N_12905);
nor U17178 (N_17178,N_13134,N_11828);
nand U17179 (N_17179,N_12811,N_10412);
nand U17180 (N_17180,N_10836,N_13632);
or U17181 (N_17181,N_14980,N_13639);
nand U17182 (N_17182,N_13066,N_11238);
nand U17183 (N_17183,N_13612,N_14974);
nor U17184 (N_17184,N_11226,N_12405);
and U17185 (N_17185,N_13397,N_14616);
nor U17186 (N_17186,N_11148,N_12469);
or U17187 (N_17187,N_14535,N_12792);
or U17188 (N_17188,N_11589,N_12900);
or U17189 (N_17189,N_11856,N_12330);
and U17190 (N_17190,N_12012,N_10045);
and U17191 (N_17191,N_12834,N_14126);
nor U17192 (N_17192,N_12816,N_10803);
or U17193 (N_17193,N_13623,N_13172);
nor U17194 (N_17194,N_11895,N_13546);
or U17195 (N_17195,N_11858,N_10828);
nor U17196 (N_17196,N_14307,N_14585);
and U17197 (N_17197,N_14676,N_11623);
and U17198 (N_17198,N_12604,N_13965);
or U17199 (N_17199,N_11158,N_10685);
nand U17200 (N_17200,N_14118,N_13031);
nor U17201 (N_17201,N_13270,N_12402);
xor U17202 (N_17202,N_13576,N_10204);
nand U17203 (N_17203,N_10087,N_14195);
nand U17204 (N_17204,N_12550,N_14651);
and U17205 (N_17205,N_14828,N_11542);
nor U17206 (N_17206,N_12630,N_12477);
and U17207 (N_17207,N_14829,N_12644);
nor U17208 (N_17208,N_14866,N_12107);
nand U17209 (N_17209,N_12255,N_13075);
and U17210 (N_17210,N_12516,N_14226);
or U17211 (N_17211,N_12068,N_11085);
or U17212 (N_17212,N_14382,N_14272);
nand U17213 (N_17213,N_11400,N_12524);
or U17214 (N_17214,N_13018,N_12649);
nand U17215 (N_17215,N_10130,N_11703);
nand U17216 (N_17216,N_12313,N_12008);
and U17217 (N_17217,N_11058,N_13200);
nand U17218 (N_17218,N_10230,N_13188);
and U17219 (N_17219,N_10688,N_10103);
nor U17220 (N_17220,N_12980,N_10899);
or U17221 (N_17221,N_12347,N_13220);
or U17222 (N_17222,N_13888,N_14819);
or U17223 (N_17223,N_12306,N_14657);
or U17224 (N_17224,N_13506,N_14884);
or U17225 (N_17225,N_11069,N_10047);
and U17226 (N_17226,N_11524,N_12835);
and U17227 (N_17227,N_12456,N_12750);
nand U17228 (N_17228,N_11926,N_12332);
or U17229 (N_17229,N_12315,N_10020);
and U17230 (N_17230,N_13819,N_14680);
nor U17231 (N_17231,N_10418,N_11476);
or U17232 (N_17232,N_11992,N_12459);
and U17233 (N_17233,N_12675,N_14568);
nand U17234 (N_17234,N_14704,N_13715);
or U17235 (N_17235,N_13953,N_10056);
nor U17236 (N_17236,N_11558,N_11068);
or U17237 (N_17237,N_12094,N_12429);
and U17238 (N_17238,N_11161,N_10719);
and U17239 (N_17239,N_12389,N_11452);
nand U17240 (N_17240,N_12629,N_12912);
or U17241 (N_17241,N_10052,N_12682);
nor U17242 (N_17242,N_11658,N_12509);
nand U17243 (N_17243,N_10470,N_11152);
nor U17244 (N_17244,N_13565,N_11854);
nand U17245 (N_17245,N_10854,N_11041);
and U17246 (N_17246,N_11831,N_14610);
or U17247 (N_17247,N_12765,N_13227);
and U17248 (N_17248,N_11083,N_12105);
nand U17249 (N_17249,N_10847,N_10481);
nand U17250 (N_17250,N_12196,N_14288);
and U17251 (N_17251,N_13766,N_14192);
nand U17252 (N_17252,N_10018,N_11329);
and U17253 (N_17253,N_12015,N_14158);
and U17254 (N_17254,N_13777,N_14445);
and U17255 (N_17255,N_10466,N_11771);
or U17256 (N_17256,N_13817,N_13112);
and U17257 (N_17257,N_10791,N_10542);
nor U17258 (N_17258,N_14623,N_10268);
and U17259 (N_17259,N_10256,N_13866);
nor U17260 (N_17260,N_13852,N_12966);
nor U17261 (N_17261,N_12151,N_12806);
nand U17262 (N_17262,N_12522,N_11548);
and U17263 (N_17263,N_11894,N_12038);
or U17264 (N_17264,N_12470,N_12585);
and U17265 (N_17265,N_12323,N_14748);
or U17266 (N_17266,N_12173,N_11219);
and U17267 (N_17267,N_13699,N_10566);
or U17268 (N_17268,N_13987,N_14130);
and U17269 (N_17269,N_10567,N_13261);
and U17270 (N_17270,N_11614,N_13025);
nand U17271 (N_17271,N_12314,N_13386);
and U17272 (N_17272,N_14115,N_13577);
and U17273 (N_17273,N_10825,N_10157);
nor U17274 (N_17274,N_11862,N_11573);
nand U17275 (N_17275,N_13855,N_12668);
or U17276 (N_17276,N_11270,N_13743);
or U17277 (N_17277,N_12678,N_10184);
nor U17278 (N_17278,N_14131,N_12768);
nor U17279 (N_17279,N_13980,N_11262);
and U17280 (N_17280,N_12988,N_13242);
and U17281 (N_17281,N_13807,N_12277);
nand U17282 (N_17282,N_12413,N_10036);
and U17283 (N_17283,N_14582,N_11796);
nor U17284 (N_17284,N_14034,N_14510);
nor U17285 (N_17285,N_13441,N_14860);
nor U17286 (N_17286,N_13007,N_12533);
and U17287 (N_17287,N_14678,N_14161);
nand U17288 (N_17288,N_13562,N_12442);
and U17289 (N_17289,N_13157,N_11765);
nand U17290 (N_17290,N_11782,N_14323);
nand U17291 (N_17291,N_10774,N_11353);
nand U17292 (N_17292,N_14039,N_11261);
or U17293 (N_17293,N_12610,N_14791);
nor U17294 (N_17294,N_14087,N_10132);
nor U17295 (N_17295,N_10550,N_14429);
and U17296 (N_17296,N_10822,N_10236);
nor U17297 (N_17297,N_14487,N_11050);
and U17298 (N_17298,N_11433,N_10592);
and U17299 (N_17299,N_14145,N_13061);
and U17300 (N_17300,N_14759,N_14909);
nand U17301 (N_17301,N_10895,N_11217);
nor U17302 (N_17302,N_11838,N_10025);
nand U17303 (N_17303,N_13194,N_11253);
nand U17304 (N_17304,N_11244,N_11951);
nor U17305 (N_17305,N_10599,N_10586);
and U17306 (N_17306,N_13040,N_13186);
or U17307 (N_17307,N_11364,N_12221);
or U17308 (N_17308,N_11464,N_11702);
and U17309 (N_17309,N_12322,N_10022);
nand U17310 (N_17310,N_10754,N_12204);
or U17311 (N_17311,N_11413,N_14468);
and U17312 (N_17312,N_12929,N_14111);
nor U17313 (N_17313,N_14788,N_11777);
nand U17314 (N_17314,N_11439,N_14376);
or U17315 (N_17315,N_12840,N_14393);
and U17316 (N_17316,N_13354,N_10759);
or U17317 (N_17317,N_11928,N_12849);
nand U17318 (N_17318,N_12858,N_13352);
or U17319 (N_17319,N_10746,N_13539);
nand U17320 (N_17320,N_10868,N_12353);
nand U17321 (N_17321,N_14199,N_11106);
nor U17322 (N_17322,N_13149,N_14480);
and U17323 (N_17323,N_11344,N_14754);
or U17324 (N_17324,N_11712,N_11499);
nor U17325 (N_17325,N_13828,N_13540);
nand U17326 (N_17326,N_12219,N_11546);
nor U17327 (N_17327,N_14347,N_11569);
nor U17328 (N_17328,N_12545,N_11602);
or U17329 (N_17329,N_10687,N_14367);
and U17330 (N_17330,N_12058,N_13448);
or U17331 (N_17331,N_12397,N_14336);
or U17332 (N_17332,N_12307,N_14475);
and U17333 (N_17333,N_13982,N_11192);
or U17334 (N_17334,N_13629,N_10541);
nor U17335 (N_17335,N_13238,N_13870);
nor U17336 (N_17336,N_14029,N_10674);
or U17337 (N_17337,N_13073,N_14057);
and U17338 (N_17338,N_14936,N_14402);
or U17339 (N_17339,N_12577,N_11864);
nand U17340 (N_17340,N_13164,N_12680);
or U17341 (N_17341,N_14009,N_11212);
or U17342 (N_17342,N_14885,N_13436);
nand U17343 (N_17343,N_13844,N_13964);
nor U17344 (N_17344,N_13732,N_11274);
and U17345 (N_17345,N_11667,N_14295);
nand U17346 (N_17346,N_13092,N_13630);
nor U17347 (N_17347,N_14739,N_10075);
and U17348 (N_17348,N_13047,N_14833);
nor U17349 (N_17349,N_12953,N_10371);
or U17350 (N_17350,N_14775,N_12031);
or U17351 (N_17351,N_10359,N_11095);
nor U17352 (N_17352,N_13528,N_11349);
and U17353 (N_17353,N_10255,N_11186);
nand U17354 (N_17354,N_11821,N_11311);
nand U17355 (N_17355,N_14705,N_13666);
and U17356 (N_17356,N_12786,N_10559);
and U17357 (N_17357,N_14690,N_11669);
nand U17358 (N_17358,N_10402,N_12244);
or U17359 (N_17359,N_13923,N_11756);
or U17360 (N_17360,N_11637,N_11533);
nor U17361 (N_17361,N_11850,N_10228);
nor U17362 (N_17362,N_10648,N_14486);
and U17363 (N_17363,N_13649,N_14992);
and U17364 (N_17364,N_13024,N_10915);
nor U17365 (N_17365,N_14174,N_14687);
and U17366 (N_17366,N_14855,N_10849);
nand U17367 (N_17367,N_11507,N_11704);
and U17368 (N_17368,N_14667,N_12074);
and U17369 (N_17369,N_10893,N_11351);
nor U17370 (N_17370,N_10630,N_12056);
and U17371 (N_17371,N_14733,N_10069);
nor U17372 (N_17372,N_10864,N_13036);
or U17373 (N_17373,N_11715,N_12752);
and U17374 (N_17374,N_12624,N_14083);
nand U17375 (N_17375,N_14976,N_14095);
or U17376 (N_17376,N_10851,N_12873);
or U17377 (N_17377,N_11595,N_11592);
and U17378 (N_17378,N_10144,N_13438);
nor U17379 (N_17379,N_12563,N_14086);
or U17380 (N_17380,N_13057,N_10843);
or U17381 (N_17381,N_10844,N_10904);
or U17382 (N_17382,N_13631,N_14440);
nand U17383 (N_17383,N_11168,N_11105);
nor U17384 (N_17384,N_10369,N_11714);
or U17385 (N_17385,N_14028,N_13925);
and U17386 (N_17386,N_14942,N_10019);
and U17387 (N_17387,N_13620,N_11600);
nand U17388 (N_17388,N_10143,N_13081);
nor U17389 (N_17389,N_11282,N_14727);
and U17390 (N_17390,N_14947,N_10270);
nand U17391 (N_17391,N_14790,N_10527);
nand U17392 (N_17392,N_12478,N_10722);
nand U17393 (N_17393,N_10081,N_11157);
nor U17394 (N_17394,N_10021,N_14620);
or U17395 (N_17395,N_11218,N_12493);
and U17396 (N_17396,N_12529,N_13955);
or U17397 (N_17397,N_14488,N_11745);
xor U17398 (N_17398,N_10456,N_13494);
nand U17399 (N_17399,N_11385,N_11650);
nand U17400 (N_17400,N_12778,N_10669);
or U17401 (N_17401,N_12492,N_11318);
nand U17402 (N_17402,N_12115,N_11857);
nand U17403 (N_17403,N_13654,N_14935);
or U17404 (N_17404,N_11435,N_13550);
nand U17405 (N_17405,N_10158,N_14660);
or U17406 (N_17406,N_11432,N_13433);
nand U17407 (N_17407,N_12916,N_14037);
nand U17408 (N_17408,N_10335,N_10478);
nand U17409 (N_17409,N_13181,N_10349);
and U17410 (N_17410,N_13892,N_10947);
and U17411 (N_17411,N_13995,N_12036);
or U17412 (N_17412,N_11007,N_14795);
nor U17413 (N_17413,N_10183,N_10827);
nor U17414 (N_17414,N_10967,N_11871);
and U17415 (N_17415,N_14031,N_13650);
nand U17416 (N_17416,N_14783,N_14906);
and U17417 (N_17417,N_14134,N_11019);
or U17418 (N_17418,N_12096,N_13549);
nor U17419 (N_17419,N_12996,N_11013);
and U17420 (N_17420,N_13215,N_13228);
or U17421 (N_17421,N_13236,N_11893);
nand U17422 (N_17422,N_12387,N_12851);
or U17423 (N_17423,N_12935,N_10927);
xor U17424 (N_17424,N_12825,N_13223);
nand U17425 (N_17425,N_14013,N_12483);
or U17426 (N_17426,N_10203,N_14560);
or U17427 (N_17427,N_11855,N_13214);
or U17428 (N_17428,N_10723,N_14681);
or U17429 (N_17429,N_13676,N_12328);
and U17430 (N_17430,N_11494,N_12077);
nand U17431 (N_17431,N_14517,N_12309);
nand U17432 (N_17432,N_10716,N_12343);
nor U17433 (N_17433,N_10345,N_13773);
and U17434 (N_17434,N_13487,N_14222);
or U17435 (N_17435,N_13502,N_12607);
nor U17436 (N_17436,N_11651,N_14908);
nor U17437 (N_17437,N_13403,N_11263);
or U17438 (N_17438,N_14059,N_14198);
or U17439 (N_17439,N_11249,N_14545);
nor U17440 (N_17440,N_14322,N_12747);
or U17441 (N_17441,N_13963,N_14967);
nand U17442 (N_17442,N_12418,N_12043);
and U17443 (N_17443,N_10537,N_11761);
and U17444 (N_17444,N_11760,N_14917);
nand U17445 (N_17445,N_13992,N_12213);
nand U17446 (N_17446,N_12489,N_13579);
or U17447 (N_17447,N_13003,N_14898);
or U17448 (N_17448,N_12370,N_13460);
nand U17449 (N_17449,N_11403,N_11987);
nand U17450 (N_17450,N_12979,N_14284);
nand U17451 (N_17451,N_12655,N_13830);
and U17452 (N_17452,N_12564,N_11886);
nand U17453 (N_17453,N_10499,N_12423);
and U17454 (N_17454,N_12587,N_10721);
nor U17455 (N_17455,N_13822,N_13571);
and U17456 (N_17456,N_13997,N_11825);
nand U17457 (N_17457,N_14789,N_13859);
and U17458 (N_17458,N_14749,N_11015);
or U17459 (N_17459,N_11438,N_10218);
or U17460 (N_17460,N_12268,N_14686);
or U17461 (N_17461,N_12132,N_11995);
and U17462 (N_17462,N_13993,N_14904);
and U17463 (N_17463,N_11799,N_12922);
nor U17464 (N_17464,N_10186,N_13694);
and U17465 (N_17465,N_13001,N_13418);
or U17466 (N_17466,N_11596,N_13059);
nand U17467 (N_17467,N_11104,N_14670);
nand U17468 (N_17468,N_14233,N_14587);
or U17469 (N_17469,N_10801,N_12910);
or U17470 (N_17470,N_10245,N_11994);
nand U17471 (N_17471,N_14477,N_14049);
or U17472 (N_17472,N_12838,N_14506);
and U17473 (N_17473,N_13570,N_13972);
nand U17474 (N_17474,N_13991,N_13415);
and U17475 (N_17475,N_10649,N_13212);
nand U17476 (N_17476,N_11549,N_13771);
nand U17477 (N_17477,N_11805,N_10306);
nand U17478 (N_17478,N_11485,N_10163);
nand U17479 (N_17479,N_13298,N_13621);
nand U17480 (N_17480,N_14991,N_13554);
or U17481 (N_17481,N_13046,N_14499);
and U17482 (N_17482,N_10666,N_11046);
nor U17483 (N_17483,N_12363,N_13901);
nand U17484 (N_17484,N_14948,N_12063);
nor U17485 (N_17485,N_14179,N_12111);
or U17486 (N_17486,N_10699,N_12502);
nand U17487 (N_17487,N_12769,N_13968);
or U17488 (N_17488,N_13105,N_10146);
or U17489 (N_17489,N_10168,N_10640);
and U17490 (N_17490,N_14169,N_10840);
nor U17491 (N_17491,N_13391,N_12685);
nor U17492 (N_17492,N_12040,N_13726);
nor U17493 (N_17493,N_11264,N_11968);
and U17494 (N_17494,N_12589,N_14397);
nand U17495 (N_17495,N_13099,N_13108);
nor U17496 (N_17496,N_13491,N_14046);
nor U17497 (N_17497,N_11880,N_14094);
nor U17498 (N_17498,N_14144,N_12158);
nor U17499 (N_17499,N_10879,N_12536);
and U17500 (N_17500,N_10379,N_11705);
and U17501 (N_17501,N_14824,N_10567);
and U17502 (N_17502,N_13389,N_10379);
and U17503 (N_17503,N_11595,N_13093);
nand U17504 (N_17504,N_10899,N_14702);
nand U17505 (N_17505,N_12694,N_10848);
nand U17506 (N_17506,N_12932,N_10519);
nand U17507 (N_17507,N_13681,N_14550);
and U17508 (N_17508,N_14300,N_12448);
or U17509 (N_17509,N_10734,N_12544);
nand U17510 (N_17510,N_14342,N_13291);
nand U17511 (N_17511,N_12342,N_12317);
and U17512 (N_17512,N_11368,N_10382);
and U17513 (N_17513,N_12862,N_13759);
nand U17514 (N_17514,N_10091,N_11113);
nor U17515 (N_17515,N_11625,N_14557);
and U17516 (N_17516,N_13506,N_14506);
nand U17517 (N_17517,N_11619,N_10115);
and U17518 (N_17518,N_14026,N_11296);
nand U17519 (N_17519,N_11151,N_10022);
nor U17520 (N_17520,N_12174,N_12132);
and U17521 (N_17521,N_14695,N_11644);
and U17522 (N_17522,N_12538,N_11272);
nand U17523 (N_17523,N_13923,N_13554);
or U17524 (N_17524,N_14366,N_13775);
or U17525 (N_17525,N_12438,N_11078);
or U17526 (N_17526,N_13434,N_10832);
nor U17527 (N_17527,N_12908,N_13149);
and U17528 (N_17528,N_11015,N_11960);
nor U17529 (N_17529,N_12136,N_13695);
and U17530 (N_17530,N_11764,N_11213);
nand U17531 (N_17531,N_10922,N_10003);
or U17532 (N_17532,N_11064,N_10061);
and U17533 (N_17533,N_14951,N_12901);
nand U17534 (N_17534,N_12683,N_11081);
and U17535 (N_17535,N_10910,N_14130);
nand U17536 (N_17536,N_13649,N_13674);
nand U17537 (N_17537,N_14775,N_14624);
or U17538 (N_17538,N_13038,N_11274);
nor U17539 (N_17539,N_10708,N_13141);
and U17540 (N_17540,N_12552,N_10230);
nor U17541 (N_17541,N_14758,N_14189);
nor U17542 (N_17542,N_14937,N_10176);
nand U17543 (N_17543,N_13764,N_12487);
or U17544 (N_17544,N_14901,N_10396);
and U17545 (N_17545,N_14002,N_12996);
or U17546 (N_17546,N_11359,N_14089);
nor U17547 (N_17547,N_12831,N_14908);
or U17548 (N_17548,N_11648,N_14771);
nor U17549 (N_17549,N_12327,N_14625);
and U17550 (N_17550,N_13026,N_14512);
or U17551 (N_17551,N_10925,N_11253);
nand U17552 (N_17552,N_13074,N_12588);
or U17553 (N_17553,N_13609,N_12160);
nor U17554 (N_17554,N_14264,N_12081);
and U17555 (N_17555,N_12168,N_10601);
nand U17556 (N_17556,N_12916,N_11057);
or U17557 (N_17557,N_14894,N_12367);
nand U17558 (N_17558,N_12363,N_13354);
or U17559 (N_17559,N_11351,N_11200);
xor U17560 (N_17560,N_13880,N_13546);
nor U17561 (N_17561,N_10226,N_13110);
nor U17562 (N_17562,N_14756,N_13768);
nor U17563 (N_17563,N_10632,N_10176);
or U17564 (N_17564,N_13936,N_14864);
nand U17565 (N_17565,N_12142,N_11148);
nor U17566 (N_17566,N_12203,N_10584);
and U17567 (N_17567,N_12870,N_13225);
and U17568 (N_17568,N_11722,N_14329);
and U17569 (N_17569,N_12945,N_13751);
and U17570 (N_17570,N_13174,N_11149);
and U17571 (N_17571,N_12740,N_12473);
nor U17572 (N_17572,N_13581,N_10142);
nor U17573 (N_17573,N_14966,N_10445);
and U17574 (N_17574,N_10342,N_12848);
nand U17575 (N_17575,N_14734,N_14309);
and U17576 (N_17576,N_14063,N_12230);
and U17577 (N_17577,N_11144,N_12688);
or U17578 (N_17578,N_10138,N_11229);
or U17579 (N_17579,N_14846,N_13594);
nor U17580 (N_17580,N_11446,N_10590);
and U17581 (N_17581,N_12040,N_10583);
or U17582 (N_17582,N_10107,N_11306);
nand U17583 (N_17583,N_12263,N_11103);
nor U17584 (N_17584,N_12141,N_12596);
nor U17585 (N_17585,N_11127,N_14671);
nand U17586 (N_17586,N_14630,N_10341);
and U17587 (N_17587,N_14707,N_12702);
nand U17588 (N_17588,N_14490,N_10414);
and U17589 (N_17589,N_11208,N_13524);
nor U17590 (N_17590,N_14565,N_13548);
nand U17591 (N_17591,N_14339,N_12584);
nand U17592 (N_17592,N_11901,N_10919);
and U17593 (N_17593,N_10670,N_11581);
nand U17594 (N_17594,N_13349,N_12002);
or U17595 (N_17595,N_11978,N_13533);
nand U17596 (N_17596,N_13841,N_11196);
xnor U17597 (N_17597,N_10528,N_10749);
or U17598 (N_17598,N_14788,N_10115);
nor U17599 (N_17599,N_14194,N_14895);
and U17600 (N_17600,N_13599,N_14001);
nor U17601 (N_17601,N_14921,N_10817);
nor U17602 (N_17602,N_11486,N_13936);
nand U17603 (N_17603,N_12721,N_12185);
nand U17604 (N_17604,N_13877,N_11632);
and U17605 (N_17605,N_12800,N_11365);
and U17606 (N_17606,N_13822,N_14019);
and U17607 (N_17607,N_13608,N_13536);
or U17608 (N_17608,N_11178,N_13984);
or U17609 (N_17609,N_14513,N_13586);
nand U17610 (N_17610,N_12953,N_12058);
nor U17611 (N_17611,N_13649,N_13770);
nor U17612 (N_17612,N_11687,N_10888);
nor U17613 (N_17613,N_10757,N_11027);
nor U17614 (N_17614,N_13545,N_14203);
or U17615 (N_17615,N_10859,N_13949);
or U17616 (N_17616,N_13657,N_14374);
and U17617 (N_17617,N_12376,N_12932);
and U17618 (N_17618,N_14247,N_10245);
and U17619 (N_17619,N_10276,N_13803);
nor U17620 (N_17620,N_11628,N_13876);
nand U17621 (N_17621,N_12287,N_13769);
nor U17622 (N_17622,N_12192,N_12141);
or U17623 (N_17623,N_14143,N_14482);
nor U17624 (N_17624,N_13979,N_10547);
nand U17625 (N_17625,N_13597,N_13087);
or U17626 (N_17626,N_10065,N_10810);
and U17627 (N_17627,N_13670,N_10748);
nand U17628 (N_17628,N_10290,N_13261);
or U17629 (N_17629,N_13560,N_13267);
nor U17630 (N_17630,N_10625,N_10484);
nor U17631 (N_17631,N_11417,N_10743);
xor U17632 (N_17632,N_12031,N_12380);
nor U17633 (N_17633,N_11325,N_14513);
or U17634 (N_17634,N_10052,N_12445);
or U17635 (N_17635,N_12344,N_11539);
or U17636 (N_17636,N_10055,N_13392);
nor U17637 (N_17637,N_12381,N_11635);
or U17638 (N_17638,N_11971,N_11455);
nor U17639 (N_17639,N_11930,N_14308);
nand U17640 (N_17640,N_10978,N_12390);
or U17641 (N_17641,N_14020,N_11238);
nor U17642 (N_17642,N_14895,N_13334);
nor U17643 (N_17643,N_14562,N_14358);
nand U17644 (N_17644,N_12901,N_14918);
nand U17645 (N_17645,N_11602,N_12843);
nand U17646 (N_17646,N_11309,N_12643);
and U17647 (N_17647,N_12847,N_12647);
or U17648 (N_17648,N_11096,N_12613);
and U17649 (N_17649,N_13421,N_14154);
nand U17650 (N_17650,N_13608,N_11469);
nor U17651 (N_17651,N_11274,N_12293);
nor U17652 (N_17652,N_11348,N_10663);
nand U17653 (N_17653,N_11384,N_12310);
and U17654 (N_17654,N_11422,N_14368);
nand U17655 (N_17655,N_10366,N_11440);
or U17656 (N_17656,N_11798,N_14337);
and U17657 (N_17657,N_12045,N_10603);
and U17658 (N_17658,N_11782,N_10049);
nand U17659 (N_17659,N_12709,N_11568);
or U17660 (N_17660,N_11638,N_13091);
nor U17661 (N_17661,N_11270,N_11565);
and U17662 (N_17662,N_12241,N_10817);
and U17663 (N_17663,N_10966,N_11307);
and U17664 (N_17664,N_14280,N_12041);
and U17665 (N_17665,N_12105,N_12924);
or U17666 (N_17666,N_12766,N_14066);
or U17667 (N_17667,N_12986,N_11584);
nand U17668 (N_17668,N_13965,N_12492);
and U17669 (N_17669,N_11999,N_14081);
nor U17670 (N_17670,N_12360,N_14575);
nand U17671 (N_17671,N_13108,N_12816);
or U17672 (N_17672,N_13758,N_10494);
nor U17673 (N_17673,N_12559,N_14930);
and U17674 (N_17674,N_11703,N_10229);
nor U17675 (N_17675,N_11129,N_11460);
or U17676 (N_17676,N_14638,N_12972);
and U17677 (N_17677,N_11305,N_13142);
nor U17678 (N_17678,N_11092,N_12228);
nand U17679 (N_17679,N_11695,N_11240);
nor U17680 (N_17680,N_12354,N_11121);
or U17681 (N_17681,N_12548,N_11017);
nor U17682 (N_17682,N_14488,N_12548);
or U17683 (N_17683,N_10900,N_14186);
or U17684 (N_17684,N_10755,N_14276);
nor U17685 (N_17685,N_13956,N_11090);
or U17686 (N_17686,N_14135,N_11825);
nor U17687 (N_17687,N_12670,N_12166);
nand U17688 (N_17688,N_12243,N_12325);
and U17689 (N_17689,N_12703,N_10590);
nand U17690 (N_17690,N_13247,N_11772);
nand U17691 (N_17691,N_13293,N_12789);
nor U17692 (N_17692,N_13097,N_14590);
nand U17693 (N_17693,N_11717,N_10647);
and U17694 (N_17694,N_10783,N_12763);
or U17695 (N_17695,N_10197,N_13766);
or U17696 (N_17696,N_11657,N_10604);
and U17697 (N_17697,N_10060,N_12383);
and U17698 (N_17698,N_12584,N_13696);
nor U17699 (N_17699,N_12181,N_10812);
nor U17700 (N_17700,N_12442,N_14019);
nand U17701 (N_17701,N_13469,N_10285);
or U17702 (N_17702,N_10808,N_13055);
and U17703 (N_17703,N_13915,N_12702);
or U17704 (N_17704,N_10387,N_10640);
nand U17705 (N_17705,N_14818,N_13873);
nor U17706 (N_17706,N_14931,N_10577);
and U17707 (N_17707,N_13527,N_11654);
nor U17708 (N_17708,N_12793,N_10721);
nand U17709 (N_17709,N_11787,N_10112);
nand U17710 (N_17710,N_13803,N_12699);
or U17711 (N_17711,N_14023,N_13791);
nand U17712 (N_17712,N_12695,N_12570);
nand U17713 (N_17713,N_11415,N_12022);
nor U17714 (N_17714,N_11817,N_12375);
and U17715 (N_17715,N_12420,N_11754);
and U17716 (N_17716,N_12877,N_10833);
nand U17717 (N_17717,N_11339,N_14458);
nor U17718 (N_17718,N_11905,N_10261);
nand U17719 (N_17719,N_12769,N_14833);
or U17720 (N_17720,N_13872,N_13218);
or U17721 (N_17721,N_12280,N_11739);
or U17722 (N_17722,N_12119,N_12115);
and U17723 (N_17723,N_12124,N_13221);
and U17724 (N_17724,N_13844,N_14914);
or U17725 (N_17725,N_10025,N_13786);
and U17726 (N_17726,N_13258,N_12552);
nor U17727 (N_17727,N_12693,N_11169);
and U17728 (N_17728,N_11862,N_10018);
nand U17729 (N_17729,N_13001,N_13688);
nor U17730 (N_17730,N_11066,N_13108);
or U17731 (N_17731,N_12052,N_13439);
or U17732 (N_17732,N_10159,N_10430);
and U17733 (N_17733,N_13448,N_12587);
and U17734 (N_17734,N_11399,N_10094);
or U17735 (N_17735,N_12585,N_14812);
nand U17736 (N_17736,N_10802,N_12081);
and U17737 (N_17737,N_12088,N_11214);
nor U17738 (N_17738,N_13538,N_10883);
or U17739 (N_17739,N_11839,N_11638);
and U17740 (N_17740,N_10150,N_13326);
nor U17741 (N_17741,N_14207,N_12009);
and U17742 (N_17742,N_14068,N_10773);
and U17743 (N_17743,N_10032,N_14757);
and U17744 (N_17744,N_12187,N_12542);
and U17745 (N_17745,N_10683,N_10463);
nor U17746 (N_17746,N_11241,N_13550);
nor U17747 (N_17747,N_11434,N_11679);
nor U17748 (N_17748,N_11049,N_14389);
nand U17749 (N_17749,N_10402,N_12730);
nor U17750 (N_17750,N_11564,N_14402);
nand U17751 (N_17751,N_11590,N_12528);
nor U17752 (N_17752,N_12601,N_12062);
and U17753 (N_17753,N_11009,N_14602);
nor U17754 (N_17754,N_12137,N_12627);
and U17755 (N_17755,N_11587,N_11197);
nand U17756 (N_17756,N_12861,N_11661);
or U17757 (N_17757,N_14484,N_14524);
and U17758 (N_17758,N_13446,N_10089);
or U17759 (N_17759,N_13390,N_13117);
or U17760 (N_17760,N_13786,N_11273);
nor U17761 (N_17761,N_13703,N_11269);
or U17762 (N_17762,N_10479,N_12770);
and U17763 (N_17763,N_14872,N_10134);
nor U17764 (N_17764,N_14054,N_10451);
nor U17765 (N_17765,N_12810,N_14361);
nand U17766 (N_17766,N_14853,N_13844);
nor U17767 (N_17767,N_13925,N_11819);
or U17768 (N_17768,N_13519,N_14552);
nor U17769 (N_17769,N_12050,N_13080);
and U17770 (N_17770,N_12036,N_11008);
nand U17771 (N_17771,N_13005,N_12750);
or U17772 (N_17772,N_13642,N_14481);
nor U17773 (N_17773,N_12725,N_13360);
and U17774 (N_17774,N_12938,N_11294);
xnor U17775 (N_17775,N_13864,N_12034);
nor U17776 (N_17776,N_11364,N_13502);
or U17777 (N_17777,N_10544,N_11307);
or U17778 (N_17778,N_10699,N_13851);
or U17779 (N_17779,N_14192,N_13904);
nand U17780 (N_17780,N_12401,N_11120);
and U17781 (N_17781,N_14124,N_10859);
and U17782 (N_17782,N_13643,N_10744);
nand U17783 (N_17783,N_12634,N_10108);
and U17784 (N_17784,N_12037,N_12184);
nor U17785 (N_17785,N_12220,N_10508);
nor U17786 (N_17786,N_10636,N_13882);
nand U17787 (N_17787,N_12012,N_10754);
xnor U17788 (N_17788,N_11149,N_10009);
or U17789 (N_17789,N_10254,N_13691);
xnor U17790 (N_17790,N_10330,N_14660);
nand U17791 (N_17791,N_13855,N_13480);
or U17792 (N_17792,N_14157,N_11253);
nor U17793 (N_17793,N_13420,N_13749);
nor U17794 (N_17794,N_13674,N_14866);
and U17795 (N_17795,N_14261,N_10248);
nor U17796 (N_17796,N_13475,N_10607);
or U17797 (N_17797,N_12669,N_11848);
nor U17798 (N_17798,N_13512,N_11819);
and U17799 (N_17799,N_11898,N_14248);
and U17800 (N_17800,N_10790,N_10368);
or U17801 (N_17801,N_10313,N_10004);
nor U17802 (N_17802,N_10785,N_11961);
and U17803 (N_17803,N_11253,N_10364);
or U17804 (N_17804,N_10360,N_14571);
nand U17805 (N_17805,N_10255,N_14137);
and U17806 (N_17806,N_11881,N_14807);
nand U17807 (N_17807,N_14340,N_12637);
or U17808 (N_17808,N_12975,N_10589);
or U17809 (N_17809,N_10352,N_12312);
nand U17810 (N_17810,N_14380,N_14117);
nand U17811 (N_17811,N_14154,N_10670);
nand U17812 (N_17812,N_10716,N_10307);
nor U17813 (N_17813,N_12588,N_13783);
nand U17814 (N_17814,N_13330,N_12750);
or U17815 (N_17815,N_11426,N_13192);
nand U17816 (N_17816,N_12370,N_10662);
and U17817 (N_17817,N_10705,N_13464);
or U17818 (N_17818,N_11037,N_12267);
nor U17819 (N_17819,N_11653,N_12947);
nand U17820 (N_17820,N_12063,N_13118);
nand U17821 (N_17821,N_10764,N_10139);
nand U17822 (N_17822,N_14215,N_14728);
and U17823 (N_17823,N_11386,N_10681);
nand U17824 (N_17824,N_10671,N_11195);
or U17825 (N_17825,N_14712,N_10357);
nor U17826 (N_17826,N_10622,N_13512);
nor U17827 (N_17827,N_11812,N_12933);
nor U17828 (N_17828,N_11559,N_14810);
nor U17829 (N_17829,N_12817,N_13787);
nor U17830 (N_17830,N_12289,N_14598);
nand U17831 (N_17831,N_14558,N_10050);
nor U17832 (N_17832,N_10533,N_13712);
nor U17833 (N_17833,N_14321,N_13240);
nand U17834 (N_17834,N_12562,N_13858);
nor U17835 (N_17835,N_14403,N_11963);
or U17836 (N_17836,N_14274,N_13471);
nand U17837 (N_17837,N_14672,N_12580);
or U17838 (N_17838,N_12305,N_14466);
and U17839 (N_17839,N_10387,N_10482);
nand U17840 (N_17840,N_11008,N_14967);
and U17841 (N_17841,N_10376,N_14536);
or U17842 (N_17842,N_13731,N_13366);
and U17843 (N_17843,N_11697,N_10726);
and U17844 (N_17844,N_11194,N_12666);
nor U17845 (N_17845,N_13101,N_11768);
nand U17846 (N_17846,N_12764,N_10652);
or U17847 (N_17847,N_11148,N_11696);
nor U17848 (N_17848,N_11461,N_13013);
or U17849 (N_17849,N_10280,N_11905);
and U17850 (N_17850,N_10375,N_11595);
or U17851 (N_17851,N_11298,N_12170);
or U17852 (N_17852,N_12597,N_10407);
and U17853 (N_17853,N_14461,N_11882);
and U17854 (N_17854,N_11223,N_12995);
or U17855 (N_17855,N_12725,N_11110);
or U17856 (N_17856,N_13389,N_11391);
and U17857 (N_17857,N_13050,N_14195);
nand U17858 (N_17858,N_12208,N_11174);
nand U17859 (N_17859,N_10993,N_10479);
or U17860 (N_17860,N_14110,N_13872);
nand U17861 (N_17861,N_11076,N_11545);
or U17862 (N_17862,N_12332,N_12542);
xor U17863 (N_17863,N_14030,N_10845);
nor U17864 (N_17864,N_13964,N_13838);
or U17865 (N_17865,N_10342,N_14595);
and U17866 (N_17866,N_13045,N_14969);
nor U17867 (N_17867,N_10631,N_14262);
nor U17868 (N_17868,N_13714,N_14420);
nor U17869 (N_17869,N_11402,N_14945);
and U17870 (N_17870,N_11214,N_13551);
and U17871 (N_17871,N_11424,N_13141);
nand U17872 (N_17872,N_11047,N_13870);
or U17873 (N_17873,N_12232,N_11318);
nor U17874 (N_17874,N_13987,N_11881);
and U17875 (N_17875,N_14694,N_13591);
and U17876 (N_17876,N_11293,N_12351);
nor U17877 (N_17877,N_10176,N_14309);
and U17878 (N_17878,N_14118,N_12061);
nor U17879 (N_17879,N_11355,N_12786);
nand U17880 (N_17880,N_14790,N_11552);
and U17881 (N_17881,N_12776,N_11817);
nand U17882 (N_17882,N_14958,N_11740);
or U17883 (N_17883,N_10784,N_11471);
nand U17884 (N_17884,N_11730,N_13866);
and U17885 (N_17885,N_13271,N_10732);
and U17886 (N_17886,N_14105,N_14797);
or U17887 (N_17887,N_11045,N_12616);
or U17888 (N_17888,N_11264,N_10119);
nor U17889 (N_17889,N_10700,N_12960);
nor U17890 (N_17890,N_13046,N_14004);
nand U17891 (N_17891,N_13465,N_14637);
and U17892 (N_17892,N_12410,N_13554);
nor U17893 (N_17893,N_14672,N_13494);
nor U17894 (N_17894,N_10188,N_11058);
nor U17895 (N_17895,N_14948,N_12014);
nor U17896 (N_17896,N_14465,N_13044);
and U17897 (N_17897,N_14083,N_14502);
nand U17898 (N_17898,N_14727,N_10826);
nor U17899 (N_17899,N_12393,N_14795);
nand U17900 (N_17900,N_12738,N_11421);
or U17901 (N_17901,N_10016,N_12561);
and U17902 (N_17902,N_14121,N_14619);
and U17903 (N_17903,N_13100,N_11070);
nand U17904 (N_17904,N_12611,N_11468);
nand U17905 (N_17905,N_10431,N_12172);
nor U17906 (N_17906,N_11457,N_13147);
or U17907 (N_17907,N_12655,N_14562);
nand U17908 (N_17908,N_14611,N_14719);
and U17909 (N_17909,N_13079,N_11473);
or U17910 (N_17910,N_13275,N_10971);
and U17911 (N_17911,N_12694,N_11428);
nand U17912 (N_17912,N_14593,N_14537);
and U17913 (N_17913,N_13312,N_12624);
and U17914 (N_17914,N_11892,N_14069);
and U17915 (N_17915,N_14756,N_12266);
and U17916 (N_17916,N_14025,N_11963);
nor U17917 (N_17917,N_13054,N_14442);
or U17918 (N_17918,N_14553,N_11283);
and U17919 (N_17919,N_10487,N_14001);
and U17920 (N_17920,N_13231,N_10332);
nor U17921 (N_17921,N_12856,N_13349);
nor U17922 (N_17922,N_12448,N_10562);
or U17923 (N_17923,N_14500,N_11885);
nor U17924 (N_17924,N_10652,N_11328);
or U17925 (N_17925,N_14230,N_14247);
or U17926 (N_17926,N_10983,N_10106);
and U17927 (N_17927,N_10250,N_13006);
and U17928 (N_17928,N_11656,N_11180);
or U17929 (N_17929,N_14486,N_13278);
nor U17930 (N_17930,N_13221,N_14957);
or U17931 (N_17931,N_14279,N_10505);
and U17932 (N_17932,N_12620,N_14423);
nor U17933 (N_17933,N_13571,N_12382);
or U17934 (N_17934,N_10318,N_13475);
nand U17935 (N_17935,N_13738,N_10552);
nand U17936 (N_17936,N_11504,N_12871);
or U17937 (N_17937,N_14143,N_12202);
and U17938 (N_17938,N_13576,N_14993);
nor U17939 (N_17939,N_10918,N_10508);
and U17940 (N_17940,N_10464,N_10056);
or U17941 (N_17941,N_10277,N_10087);
nor U17942 (N_17942,N_13472,N_12748);
nor U17943 (N_17943,N_11352,N_11981);
nand U17944 (N_17944,N_14140,N_13136);
or U17945 (N_17945,N_11389,N_10939);
or U17946 (N_17946,N_13504,N_11497);
and U17947 (N_17947,N_12190,N_12800);
and U17948 (N_17948,N_12636,N_10924);
or U17949 (N_17949,N_11987,N_10001);
and U17950 (N_17950,N_14250,N_14733);
nand U17951 (N_17951,N_13473,N_13844);
and U17952 (N_17952,N_13576,N_10877);
and U17953 (N_17953,N_13295,N_13158);
and U17954 (N_17954,N_14784,N_11494);
and U17955 (N_17955,N_14791,N_13729);
or U17956 (N_17956,N_12681,N_10635);
or U17957 (N_17957,N_12237,N_13762);
and U17958 (N_17958,N_12841,N_14082);
or U17959 (N_17959,N_10958,N_12117);
and U17960 (N_17960,N_11255,N_13491);
and U17961 (N_17961,N_14740,N_12672);
nand U17962 (N_17962,N_11162,N_11462);
and U17963 (N_17963,N_10232,N_14356);
nand U17964 (N_17964,N_10702,N_12626);
or U17965 (N_17965,N_13941,N_10656);
or U17966 (N_17966,N_13786,N_11370);
nor U17967 (N_17967,N_11522,N_13710);
nand U17968 (N_17968,N_10120,N_10335);
nor U17969 (N_17969,N_14918,N_10048);
nand U17970 (N_17970,N_14027,N_14823);
and U17971 (N_17971,N_13063,N_10307);
or U17972 (N_17972,N_11367,N_11406);
and U17973 (N_17973,N_10376,N_13011);
and U17974 (N_17974,N_12284,N_14364);
nor U17975 (N_17975,N_12763,N_12851);
or U17976 (N_17976,N_14717,N_13458);
nand U17977 (N_17977,N_10370,N_11074);
nand U17978 (N_17978,N_10472,N_12212);
and U17979 (N_17979,N_11251,N_13878);
or U17980 (N_17980,N_11072,N_11287);
nor U17981 (N_17981,N_10697,N_11936);
nand U17982 (N_17982,N_14941,N_13617);
and U17983 (N_17983,N_10812,N_12920);
nor U17984 (N_17984,N_13918,N_14774);
nor U17985 (N_17985,N_13915,N_10162);
nand U17986 (N_17986,N_14695,N_11313);
nand U17987 (N_17987,N_14327,N_10255);
and U17988 (N_17988,N_10301,N_12550);
nor U17989 (N_17989,N_13016,N_10334);
and U17990 (N_17990,N_14133,N_14975);
and U17991 (N_17991,N_11190,N_13299);
nand U17992 (N_17992,N_14598,N_12295);
or U17993 (N_17993,N_11793,N_13295);
and U17994 (N_17994,N_13724,N_10364);
or U17995 (N_17995,N_12052,N_10113);
nand U17996 (N_17996,N_10369,N_10879);
and U17997 (N_17997,N_13323,N_13590);
nor U17998 (N_17998,N_14888,N_12450);
or U17999 (N_17999,N_10936,N_14139);
or U18000 (N_18000,N_14450,N_13683);
or U18001 (N_18001,N_13635,N_13875);
or U18002 (N_18002,N_12727,N_10101);
nor U18003 (N_18003,N_12424,N_11666);
nand U18004 (N_18004,N_13750,N_12681);
and U18005 (N_18005,N_11684,N_13489);
or U18006 (N_18006,N_14680,N_13570);
or U18007 (N_18007,N_12307,N_13227);
nand U18008 (N_18008,N_12361,N_13654);
and U18009 (N_18009,N_10373,N_14105);
nand U18010 (N_18010,N_13009,N_13643);
or U18011 (N_18011,N_14244,N_13805);
nand U18012 (N_18012,N_13058,N_10592);
nand U18013 (N_18013,N_12947,N_12597);
or U18014 (N_18014,N_13362,N_11032);
and U18015 (N_18015,N_13283,N_13986);
nor U18016 (N_18016,N_10095,N_13459);
nor U18017 (N_18017,N_12313,N_10337);
nand U18018 (N_18018,N_12679,N_12529);
nor U18019 (N_18019,N_10403,N_12967);
or U18020 (N_18020,N_13928,N_11643);
and U18021 (N_18021,N_12748,N_12597);
nor U18022 (N_18022,N_14877,N_14240);
and U18023 (N_18023,N_10480,N_13131);
nor U18024 (N_18024,N_11911,N_10073);
and U18025 (N_18025,N_10368,N_10421);
or U18026 (N_18026,N_11512,N_14854);
nand U18027 (N_18027,N_13549,N_11864);
nor U18028 (N_18028,N_13857,N_14321);
or U18029 (N_18029,N_13342,N_13232);
or U18030 (N_18030,N_13007,N_11328);
nand U18031 (N_18031,N_14683,N_14573);
nand U18032 (N_18032,N_12588,N_11783);
or U18033 (N_18033,N_12957,N_10631);
nand U18034 (N_18034,N_11226,N_11591);
or U18035 (N_18035,N_13956,N_11854);
and U18036 (N_18036,N_11129,N_14817);
nand U18037 (N_18037,N_12287,N_10141);
or U18038 (N_18038,N_11080,N_13293);
nand U18039 (N_18039,N_14804,N_14088);
or U18040 (N_18040,N_11521,N_12269);
or U18041 (N_18041,N_13286,N_14068);
or U18042 (N_18042,N_11725,N_10202);
or U18043 (N_18043,N_11117,N_10873);
or U18044 (N_18044,N_13572,N_13752);
nand U18045 (N_18045,N_11922,N_13023);
and U18046 (N_18046,N_13108,N_12716);
or U18047 (N_18047,N_10387,N_14196);
xnor U18048 (N_18048,N_11443,N_14681);
and U18049 (N_18049,N_14079,N_13024);
nor U18050 (N_18050,N_12756,N_13247);
or U18051 (N_18051,N_10347,N_12054);
nand U18052 (N_18052,N_10495,N_13311);
nor U18053 (N_18053,N_13720,N_12697);
or U18054 (N_18054,N_10608,N_12108);
and U18055 (N_18055,N_12612,N_11702);
nand U18056 (N_18056,N_13039,N_14342);
and U18057 (N_18057,N_12815,N_10494);
nand U18058 (N_18058,N_11313,N_13360);
and U18059 (N_18059,N_14740,N_12128);
or U18060 (N_18060,N_13296,N_12790);
nand U18061 (N_18061,N_12752,N_14421);
nand U18062 (N_18062,N_12777,N_11237);
or U18063 (N_18063,N_12526,N_13744);
nor U18064 (N_18064,N_14428,N_14262);
or U18065 (N_18065,N_10209,N_12670);
and U18066 (N_18066,N_14336,N_13423);
and U18067 (N_18067,N_12529,N_11640);
or U18068 (N_18068,N_10150,N_12676);
nand U18069 (N_18069,N_12603,N_12639);
or U18070 (N_18070,N_11457,N_14115);
and U18071 (N_18071,N_11324,N_10477);
or U18072 (N_18072,N_12549,N_11160);
nand U18073 (N_18073,N_14621,N_12603);
or U18074 (N_18074,N_10441,N_13223);
or U18075 (N_18075,N_13594,N_11467);
or U18076 (N_18076,N_14804,N_12053);
and U18077 (N_18077,N_13575,N_11208);
and U18078 (N_18078,N_13790,N_13170);
nand U18079 (N_18079,N_12489,N_14667);
and U18080 (N_18080,N_11521,N_13574);
nor U18081 (N_18081,N_13751,N_14930);
or U18082 (N_18082,N_13912,N_10100);
nor U18083 (N_18083,N_13770,N_10925);
or U18084 (N_18084,N_14763,N_11983);
nor U18085 (N_18085,N_14263,N_11575);
or U18086 (N_18086,N_13780,N_12028);
and U18087 (N_18087,N_10249,N_12005);
nand U18088 (N_18088,N_13459,N_12352);
nor U18089 (N_18089,N_14830,N_14735);
or U18090 (N_18090,N_11450,N_11599);
nand U18091 (N_18091,N_11463,N_10249);
xor U18092 (N_18092,N_12810,N_11694);
nand U18093 (N_18093,N_12842,N_14528);
and U18094 (N_18094,N_10793,N_14654);
nor U18095 (N_18095,N_10470,N_13120);
nand U18096 (N_18096,N_11975,N_12710);
xor U18097 (N_18097,N_13238,N_13043);
nor U18098 (N_18098,N_12688,N_13713);
or U18099 (N_18099,N_14602,N_11746);
nor U18100 (N_18100,N_13520,N_11735);
nand U18101 (N_18101,N_14115,N_12368);
and U18102 (N_18102,N_10686,N_11150);
nor U18103 (N_18103,N_13207,N_13714);
and U18104 (N_18104,N_10537,N_13158);
nor U18105 (N_18105,N_10436,N_13788);
and U18106 (N_18106,N_10623,N_10657);
nand U18107 (N_18107,N_10662,N_11891);
xnor U18108 (N_18108,N_13850,N_12785);
and U18109 (N_18109,N_12925,N_13033);
and U18110 (N_18110,N_11273,N_13605);
or U18111 (N_18111,N_14584,N_12773);
and U18112 (N_18112,N_13152,N_13482);
nand U18113 (N_18113,N_11299,N_10870);
nor U18114 (N_18114,N_11405,N_12108);
nand U18115 (N_18115,N_11336,N_11378);
or U18116 (N_18116,N_13663,N_12454);
nand U18117 (N_18117,N_10459,N_12892);
and U18118 (N_18118,N_12440,N_13123);
nand U18119 (N_18119,N_12331,N_14377);
or U18120 (N_18120,N_10764,N_14407);
nor U18121 (N_18121,N_12723,N_11478);
nor U18122 (N_18122,N_13682,N_10867);
or U18123 (N_18123,N_13727,N_10981);
nand U18124 (N_18124,N_10800,N_12550);
or U18125 (N_18125,N_11177,N_11278);
nor U18126 (N_18126,N_14173,N_11362);
nor U18127 (N_18127,N_14894,N_11524);
nor U18128 (N_18128,N_12651,N_14977);
nor U18129 (N_18129,N_11147,N_12098);
and U18130 (N_18130,N_13493,N_10678);
nand U18131 (N_18131,N_11730,N_12954);
or U18132 (N_18132,N_13796,N_13026);
nand U18133 (N_18133,N_11893,N_12973);
nand U18134 (N_18134,N_13619,N_10907);
nand U18135 (N_18135,N_11959,N_10045);
or U18136 (N_18136,N_14490,N_12386);
nand U18137 (N_18137,N_12261,N_10524);
nand U18138 (N_18138,N_12774,N_10886);
nand U18139 (N_18139,N_13805,N_11588);
nand U18140 (N_18140,N_13555,N_10976);
and U18141 (N_18141,N_12632,N_12199);
and U18142 (N_18142,N_11555,N_10967);
nor U18143 (N_18143,N_11698,N_13484);
nor U18144 (N_18144,N_14785,N_14786);
nand U18145 (N_18145,N_10214,N_13395);
nand U18146 (N_18146,N_12983,N_13884);
or U18147 (N_18147,N_10272,N_12761);
or U18148 (N_18148,N_11010,N_14291);
nor U18149 (N_18149,N_12593,N_12983);
or U18150 (N_18150,N_10455,N_12217);
and U18151 (N_18151,N_14258,N_12955);
and U18152 (N_18152,N_11431,N_10864);
nand U18153 (N_18153,N_14402,N_11038);
nor U18154 (N_18154,N_12750,N_12816);
nand U18155 (N_18155,N_14129,N_14470);
nand U18156 (N_18156,N_13757,N_10761);
xnor U18157 (N_18157,N_14613,N_13966);
nand U18158 (N_18158,N_12448,N_13535);
or U18159 (N_18159,N_11189,N_10542);
and U18160 (N_18160,N_13169,N_14423);
and U18161 (N_18161,N_13329,N_12794);
or U18162 (N_18162,N_10134,N_11604);
or U18163 (N_18163,N_14115,N_10026);
or U18164 (N_18164,N_10786,N_13061);
nor U18165 (N_18165,N_14458,N_10542);
nor U18166 (N_18166,N_13886,N_14448);
nor U18167 (N_18167,N_12633,N_13595);
nor U18168 (N_18168,N_10427,N_13565);
or U18169 (N_18169,N_14248,N_11765);
or U18170 (N_18170,N_12751,N_13805);
nor U18171 (N_18171,N_11423,N_13041);
nor U18172 (N_18172,N_13334,N_14344);
and U18173 (N_18173,N_10788,N_12192);
and U18174 (N_18174,N_14216,N_11647);
and U18175 (N_18175,N_11943,N_11261);
nand U18176 (N_18176,N_10502,N_13973);
nor U18177 (N_18177,N_10755,N_12244);
or U18178 (N_18178,N_12727,N_13448);
and U18179 (N_18179,N_10943,N_12942);
nor U18180 (N_18180,N_13799,N_10294);
and U18181 (N_18181,N_14221,N_14514);
nor U18182 (N_18182,N_10470,N_10575);
and U18183 (N_18183,N_14660,N_14265);
nor U18184 (N_18184,N_10439,N_10875);
or U18185 (N_18185,N_14981,N_12039);
and U18186 (N_18186,N_13738,N_12919);
or U18187 (N_18187,N_11999,N_12239);
or U18188 (N_18188,N_14828,N_11409);
nand U18189 (N_18189,N_10212,N_12873);
and U18190 (N_18190,N_14438,N_13864);
and U18191 (N_18191,N_10340,N_14212);
xor U18192 (N_18192,N_10641,N_13816);
and U18193 (N_18193,N_11562,N_11592);
nor U18194 (N_18194,N_11999,N_12916);
and U18195 (N_18195,N_14963,N_12483);
nand U18196 (N_18196,N_13929,N_12529);
or U18197 (N_18197,N_12895,N_12649);
or U18198 (N_18198,N_14276,N_11816);
nand U18199 (N_18199,N_12411,N_12786);
nand U18200 (N_18200,N_11382,N_10714);
nand U18201 (N_18201,N_13679,N_10092);
or U18202 (N_18202,N_10761,N_11234);
nand U18203 (N_18203,N_14082,N_11001);
or U18204 (N_18204,N_10637,N_14893);
nand U18205 (N_18205,N_11275,N_11729);
nor U18206 (N_18206,N_11544,N_12754);
nor U18207 (N_18207,N_12603,N_12792);
nor U18208 (N_18208,N_14895,N_13860);
nor U18209 (N_18209,N_13491,N_11185);
nand U18210 (N_18210,N_10482,N_13396);
nor U18211 (N_18211,N_14316,N_11155);
nand U18212 (N_18212,N_13327,N_12004);
nor U18213 (N_18213,N_12528,N_10530);
nor U18214 (N_18214,N_14538,N_14594);
or U18215 (N_18215,N_11714,N_10142);
and U18216 (N_18216,N_10673,N_11593);
nor U18217 (N_18217,N_10683,N_12705);
and U18218 (N_18218,N_12925,N_14797);
or U18219 (N_18219,N_11843,N_13739);
or U18220 (N_18220,N_12166,N_14209);
and U18221 (N_18221,N_11386,N_14849);
and U18222 (N_18222,N_10775,N_11709);
and U18223 (N_18223,N_12678,N_11585);
or U18224 (N_18224,N_10746,N_12338);
nand U18225 (N_18225,N_10020,N_14433);
or U18226 (N_18226,N_10172,N_11701);
nand U18227 (N_18227,N_11957,N_14764);
nand U18228 (N_18228,N_11246,N_11755);
nor U18229 (N_18229,N_14460,N_12319);
nor U18230 (N_18230,N_13238,N_14209);
or U18231 (N_18231,N_12892,N_13643);
or U18232 (N_18232,N_13440,N_13631);
nor U18233 (N_18233,N_11688,N_10939);
or U18234 (N_18234,N_13120,N_10724);
or U18235 (N_18235,N_10316,N_14719);
or U18236 (N_18236,N_11666,N_12484);
or U18237 (N_18237,N_12870,N_12209);
nor U18238 (N_18238,N_13888,N_13313);
or U18239 (N_18239,N_10567,N_14424);
or U18240 (N_18240,N_11500,N_10685);
and U18241 (N_18241,N_14620,N_13256);
or U18242 (N_18242,N_10234,N_10230);
nand U18243 (N_18243,N_14251,N_11851);
and U18244 (N_18244,N_10187,N_12799);
nand U18245 (N_18245,N_10360,N_11965);
nand U18246 (N_18246,N_11483,N_13071);
nand U18247 (N_18247,N_14156,N_13049);
and U18248 (N_18248,N_13186,N_11296);
and U18249 (N_18249,N_12062,N_14135);
nor U18250 (N_18250,N_11430,N_11306);
nor U18251 (N_18251,N_14476,N_14119);
nor U18252 (N_18252,N_14830,N_13277);
or U18253 (N_18253,N_14295,N_12552);
nand U18254 (N_18254,N_12348,N_13087);
and U18255 (N_18255,N_12834,N_11630);
or U18256 (N_18256,N_11187,N_14716);
and U18257 (N_18257,N_10138,N_12970);
and U18258 (N_18258,N_14534,N_10988);
nor U18259 (N_18259,N_11549,N_13571);
nand U18260 (N_18260,N_11294,N_13344);
or U18261 (N_18261,N_14794,N_13813);
or U18262 (N_18262,N_13677,N_13017);
and U18263 (N_18263,N_13276,N_13807);
nand U18264 (N_18264,N_12073,N_13486);
or U18265 (N_18265,N_11636,N_13986);
and U18266 (N_18266,N_13248,N_12897);
and U18267 (N_18267,N_10905,N_12433);
nor U18268 (N_18268,N_14940,N_11652);
or U18269 (N_18269,N_14475,N_13508);
nor U18270 (N_18270,N_14688,N_13249);
nor U18271 (N_18271,N_13908,N_12660);
nor U18272 (N_18272,N_12986,N_12566);
nand U18273 (N_18273,N_11990,N_11007);
nor U18274 (N_18274,N_10739,N_10955);
nor U18275 (N_18275,N_12039,N_11705);
nor U18276 (N_18276,N_11929,N_14004);
and U18277 (N_18277,N_14232,N_12293);
or U18278 (N_18278,N_14534,N_11959);
nand U18279 (N_18279,N_14871,N_10990);
or U18280 (N_18280,N_14182,N_14395);
nand U18281 (N_18281,N_11259,N_12738);
or U18282 (N_18282,N_12836,N_10854);
nor U18283 (N_18283,N_14098,N_11661);
nor U18284 (N_18284,N_13943,N_10798);
nor U18285 (N_18285,N_11362,N_10029);
and U18286 (N_18286,N_12116,N_10450);
or U18287 (N_18287,N_11415,N_14088);
nand U18288 (N_18288,N_12055,N_10454);
nand U18289 (N_18289,N_11040,N_12573);
and U18290 (N_18290,N_10747,N_14078);
or U18291 (N_18291,N_14122,N_11701);
and U18292 (N_18292,N_10961,N_13992);
nand U18293 (N_18293,N_13004,N_10932);
or U18294 (N_18294,N_10653,N_12558);
nand U18295 (N_18295,N_13024,N_11140);
and U18296 (N_18296,N_14869,N_14506);
and U18297 (N_18297,N_14973,N_11587);
or U18298 (N_18298,N_12320,N_12860);
or U18299 (N_18299,N_10492,N_10646);
or U18300 (N_18300,N_13778,N_11507);
nand U18301 (N_18301,N_10771,N_10441);
or U18302 (N_18302,N_11752,N_14057);
nand U18303 (N_18303,N_14942,N_13778);
or U18304 (N_18304,N_12341,N_12239);
nor U18305 (N_18305,N_12727,N_13514);
and U18306 (N_18306,N_10541,N_12451);
or U18307 (N_18307,N_11665,N_11422);
or U18308 (N_18308,N_14990,N_10640);
and U18309 (N_18309,N_12394,N_11588);
and U18310 (N_18310,N_14041,N_14356);
nor U18311 (N_18311,N_10684,N_13426);
nor U18312 (N_18312,N_14513,N_14846);
and U18313 (N_18313,N_11463,N_12389);
nand U18314 (N_18314,N_11660,N_12115);
nand U18315 (N_18315,N_13544,N_11230);
xor U18316 (N_18316,N_14277,N_10294);
nor U18317 (N_18317,N_10717,N_12882);
and U18318 (N_18318,N_12708,N_13187);
and U18319 (N_18319,N_12375,N_14394);
nand U18320 (N_18320,N_13946,N_11151);
or U18321 (N_18321,N_11900,N_12673);
and U18322 (N_18322,N_12214,N_11673);
nand U18323 (N_18323,N_10172,N_14911);
or U18324 (N_18324,N_10159,N_10576);
nor U18325 (N_18325,N_10525,N_12489);
nor U18326 (N_18326,N_10204,N_13174);
and U18327 (N_18327,N_10354,N_10346);
nand U18328 (N_18328,N_14526,N_14159);
and U18329 (N_18329,N_11552,N_14902);
nor U18330 (N_18330,N_12044,N_12841);
nand U18331 (N_18331,N_12363,N_13880);
and U18332 (N_18332,N_14621,N_10940);
and U18333 (N_18333,N_11963,N_12946);
or U18334 (N_18334,N_10090,N_12828);
and U18335 (N_18335,N_13104,N_14075);
nand U18336 (N_18336,N_13741,N_11536);
or U18337 (N_18337,N_14943,N_13416);
and U18338 (N_18338,N_14296,N_13441);
nand U18339 (N_18339,N_10589,N_10536);
xnor U18340 (N_18340,N_13677,N_14434);
or U18341 (N_18341,N_12043,N_12305);
nor U18342 (N_18342,N_13830,N_12927);
and U18343 (N_18343,N_13903,N_10631);
nor U18344 (N_18344,N_12350,N_13035);
or U18345 (N_18345,N_13364,N_12756);
nand U18346 (N_18346,N_14185,N_10064);
and U18347 (N_18347,N_13271,N_13238);
and U18348 (N_18348,N_12436,N_11137);
and U18349 (N_18349,N_11695,N_13381);
nand U18350 (N_18350,N_10140,N_10529);
nor U18351 (N_18351,N_11664,N_13483);
or U18352 (N_18352,N_11626,N_11821);
and U18353 (N_18353,N_13850,N_11860);
or U18354 (N_18354,N_11080,N_14174);
nor U18355 (N_18355,N_11761,N_12964);
or U18356 (N_18356,N_12321,N_12288);
nor U18357 (N_18357,N_13731,N_14143);
nor U18358 (N_18358,N_13552,N_10413);
and U18359 (N_18359,N_12962,N_11326);
nor U18360 (N_18360,N_10515,N_13380);
or U18361 (N_18361,N_11929,N_14659);
or U18362 (N_18362,N_10529,N_12007);
nor U18363 (N_18363,N_11911,N_13913);
nand U18364 (N_18364,N_13774,N_10594);
nand U18365 (N_18365,N_14820,N_14791);
and U18366 (N_18366,N_11771,N_10581);
xor U18367 (N_18367,N_11521,N_14374);
nand U18368 (N_18368,N_12970,N_13891);
nand U18369 (N_18369,N_10938,N_11538);
nor U18370 (N_18370,N_13065,N_12157);
nor U18371 (N_18371,N_14238,N_11648);
and U18372 (N_18372,N_13718,N_13287);
or U18373 (N_18373,N_14892,N_10735);
nand U18374 (N_18374,N_12646,N_13541);
or U18375 (N_18375,N_14514,N_10127);
nand U18376 (N_18376,N_10426,N_13793);
nor U18377 (N_18377,N_14586,N_11908);
nand U18378 (N_18378,N_14058,N_14874);
and U18379 (N_18379,N_11314,N_10892);
or U18380 (N_18380,N_12420,N_10380);
and U18381 (N_18381,N_13486,N_14129);
nor U18382 (N_18382,N_14927,N_12700);
nor U18383 (N_18383,N_10737,N_14957);
and U18384 (N_18384,N_12335,N_10846);
nand U18385 (N_18385,N_12658,N_11073);
and U18386 (N_18386,N_10330,N_14705);
or U18387 (N_18387,N_14205,N_14793);
nor U18388 (N_18388,N_11518,N_10304);
or U18389 (N_18389,N_13753,N_10129);
and U18390 (N_18390,N_13445,N_11593);
xor U18391 (N_18391,N_14341,N_13783);
and U18392 (N_18392,N_14048,N_14422);
and U18393 (N_18393,N_10336,N_10560);
nor U18394 (N_18394,N_13981,N_13312);
or U18395 (N_18395,N_10249,N_14650);
or U18396 (N_18396,N_10242,N_14752);
or U18397 (N_18397,N_12902,N_11366);
or U18398 (N_18398,N_11261,N_12091);
or U18399 (N_18399,N_12733,N_13935);
and U18400 (N_18400,N_12509,N_12340);
or U18401 (N_18401,N_11219,N_10125);
nor U18402 (N_18402,N_12517,N_12130);
nand U18403 (N_18403,N_13765,N_13577);
and U18404 (N_18404,N_13055,N_10110);
nor U18405 (N_18405,N_14595,N_11776);
and U18406 (N_18406,N_11695,N_11066);
nand U18407 (N_18407,N_11758,N_11926);
xor U18408 (N_18408,N_10424,N_14521);
or U18409 (N_18409,N_13307,N_11770);
and U18410 (N_18410,N_13333,N_12908);
nand U18411 (N_18411,N_14092,N_12511);
nor U18412 (N_18412,N_14147,N_10294);
nand U18413 (N_18413,N_11449,N_13959);
or U18414 (N_18414,N_11714,N_13265);
and U18415 (N_18415,N_14647,N_10093);
and U18416 (N_18416,N_10348,N_10418);
nand U18417 (N_18417,N_13270,N_11793);
or U18418 (N_18418,N_10046,N_10037);
and U18419 (N_18419,N_12318,N_10826);
nand U18420 (N_18420,N_10257,N_11517);
nand U18421 (N_18421,N_13914,N_12014);
and U18422 (N_18422,N_10409,N_14395);
or U18423 (N_18423,N_12520,N_13191);
nor U18424 (N_18424,N_10123,N_14320);
nand U18425 (N_18425,N_13301,N_11551);
nand U18426 (N_18426,N_13265,N_13598);
or U18427 (N_18427,N_14463,N_11891);
and U18428 (N_18428,N_14292,N_11959);
or U18429 (N_18429,N_13628,N_13253);
or U18430 (N_18430,N_13830,N_13549);
or U18431 (N_18431,N_10745,N_11920);
or U18432 (N_18432,N_11552,N_11217);
nor U18433 (N_18433,N_11314,N_12005);
and U18434 (N_18434,N_12653,N_11979);
or U18435 (N_18435,N_12086,N_14517);
nand U18436 (N_18436,N_11435,N_11123);
nand U18437 (N_18437,N_10221,N_11630);
nand U18438 (N_18438,N_14203,N_13508);
nor U18439 (N_18439,N_14131,N_11844);
or U18440 (N_18440,N_13473,N_14116);
or U18441 (N_18441,N_14596,N_12894);
nand U18442 (N_18442,N_11745,N_11410);
or U18443 (N_18443,N_11910,N_11688);
or U18444 (N_18444,N_14740,N_13929);
or U18445 (N_18445,N_10691,N_14887);
nand U18446 (N_18446,N_14477,N_12330);
or U18447 (N_18447,N_13545,N_14277);
nor U18448 (N_18448,N_13964,N_10517);
nand U18449 (N_18449,N_13417,N_11660);
xor U18450 (N_18450,N_10689,N_13828);
nor U18451 (N_18451,N_10271,N_11966);
nor U18452 (N_18452,N_14688,N_13512);
or U18453 (N_18453,N_14936,N_14750);
xnor U18454 (N_18454,N_12843,N_10987);
nor U18455 (N_18455,N_10350,N_12730);
and U18456 (N_18456,N_10649,N_11370);
nand U18457 (N_18457,N_13225,N_11137);
and U18458 (N_18458,N_12565,N_14660);
nand U18459 (N_18459,N_10450,N_13411);
and U18460 (N_18460,N_14323,N_12398);
or U18461 (N_18461,N_11042,N_10755);
or U18462 (N_18462,N_10244,N_13771);
or U18463 (N_18463,N_12450,N_12100);
nor U18464 (N_18464,N_14329,N_14237);
nor U18465 (N_18465,N_12387,N_11919);
nor U18466 (N_18466,N_11055,N_10578);
or U18467 (N_18467,N_14965,N_13471);
or U18468 (N_18468,N_10235,N_13098);
nor U18469 (N_18469,N_12999,N_11801);
xor U18470 (N_18470,N_10158,N_14989);
or U18471 (N_18471,N_10464,N_13968);
or U18472 (N_18472,N_14355,N_14731);
and U18473 (N_18473,N_14913,N_10107);
nand U18474 (N_18474,N_10244,N_14360);
and U18475 (N_18475,N_12433,N_13131);
nor U18476 (N_18476,N_14112,N_13716);
or U18477 (N_18477,N_13223,N_10981);
nand U18478 (N_18478,N_12483,N_11987);
and U18479 (N_18479,N_12198,N_12654);
or U18480 (N_18480,N_12871,N_13387);
nor U18481 (N_18481,N_12740,N_13467);
nand U18482 (N_18482,N_14909,N_14833);
nand U18483 (N_18483,N_14474,N_12213);
and U18484 (N_18484,N_13808,N_12566);
or U18485 (N_18485,N_13630,N_13316);
or U18486 (N_18486,N_10175,N_12158);
nand U18487 (N_18487,N_10637,N_11004);
nand U18488 (N_18488,N_14344,N_13265);
nand U18489 (N_18489,N_12286,N_10259);
and U18490 (N_18490,N_14537,N_10611);
nor U18491 (N_18491,N_13301,N_12211);
nand U18492 (N_18492,N_12413,N_10802);
nand U18493 (N_18493,N_14214,N_13291);
nor U18494 (N_18494,N_10239,N_14382);
and U18495 (N_18495,N_14110,N_12681);
or U18496 (N_18496,N_12551,N_12963);
or U18497 (N_18497,N_14871,N_11722);
or U18498 (N_18498,N_12847,N_14351);
nor U18499 (N_18499,N_14936,N_11496);
and U18500 (N_18500,N_13324,N_12409);
nand U18501 (N_18501,N_13400,N_10020);
and U18502 (N_18502,N_13842,N_10160);
nor U18503 (N_18503,N_13874,N_11201);
and U18504 (N_18504,N_14113,N_13718);
nor U18505 (N_18505,N_10620,N_13019);
and U18506 (N_18506,N_11399,N_11324);
or U18507 (N_18507,N_12601,N_13811);
and U18508 (N_18508,N_10179,N_12912);
nand U18509 (N_18509,N_14146,N_12985);
or U18510 (N_18510,N_11263,N_10766);
nor U18511 (N_18511,N_12826,N_13198);
or U18512 (N_18512,N_10424,N_10620);
nand U18513 (N_18513,N_11039,N_10110);
and U18514 (N_18514,N_10639,N_14564);
nor U18515 (N_18515,N_12816,N_11406);
nor U18516 (N_18516,N_14576,N_14955);
or U18517 (N_18517,N_14065,N_14927);
and U18518 (N_18518,N_12559,N_13968);
and U18519 (N_18519,N_12355,N_11080);
nor U18520 (N_18520,N_13931,N_10943);
or U18521 (N_18521,N_10358,N_10923);
and U18522 (N_18522,N_13283,N_14388);
and U18523 (N_18523,N_14238,N_13660);
or U18524 (N_18524,N_14701,N_12719);
or U18525 (N_18525,N_14095,N_13014);
and U18526 (N_18526,N_14406,N_12547);
and U18527 (N_18527,N_11606,N_10467);
nand U18528 (N_18528,N_14869,N_11177);
nor U18529 (N_18529,N_13775,N_10911);
nor U18530 (N_18530,N_12317,N_10263);
nand U18531 (N_18531,N_14191,N_12256);
or U18532 (N_18532,N_12091,N_10254);
or U18533 (N_18533,N_14671,N_10315);
and U18534 (N_18534,N_14764,N_11555);
or U18535 (N_18535,N_11375,N_14832);
and U18536 (N_18536,N_13143,N_10355);
or U18537 (N_18537,N_12347,N_14049);
or U18538 (N_18538,N_14837,N_12428);
or U18539 (N_18539,N_10248,N_11263);
nand U18540 (N_18540,N_14206,N_10648);
nand U18541 (N_18541,N_12660,N_11363);
and U18542 (N_18542,N_11204,N_11020);
or U18543 (N_18543,N_11468,N_12668);
nand U18544 (N_18544,N_11506,N_10967);
and U18545 (N_18545,N_10285,N_11537);
nand U18546 (N_18546,N_12968,N_10171);
nor U18547 (N_18547,N_11645,N_14626);
and U18548 (N_18548,N_12145,N_10262);
nand U18549 (N_18549,N_11235,N_13767);
or U18550 (N_18550,N_12520,N_10480);
nand U18551 (N_18551,N_10605,N_12156);
nand U18552 (N_18552,N_13788,N_10037);
or U18553 (N_18553,N_10993,N_14898);
and U18554 (N_18554,N_14456,N_13431);
nand U18555 (N_18555,N_12592,N_12840);
and U18556 (N_18556,N_12079,N_14425);
and U18557 (N_18557,N_13097,N_11319);
nand U18558 (N_18558,N_10769,N_10970);
nand U18559 (N_18559,N_11815,N_13077);
nand U18560 (N_18560,N_12189,N_12378);
nand U18561 (N_18561,N_10539,N_11308);
or U18562 (N_18562,N_10212,N_12633);
or U18563 (N_18563,N_10907,N_11002);
nor U18564 (N_18564,N_12640,N_12231);
or U18565 (N_18565,N_13057,N_14406);
nand U18566 (N_18566,N_10909,N_13280);
or U18567 (N_18567,N_14467,N_14367);
nor U18568 (N_18568,N_12587,N_14740);
or U18569 (N_18569,N_13148,N_14797);
and U18570 (N_18570,N_12411,N_13564);
nor U18571 (N_18571,N_14009,N_12749);
nand U18572 (N_18572,N_13955,N_11527);
and U18573 (N_18573,N_14701,N_11163);
nand U18574 (N_18574,N_11300,N_11988);
and U18575 (N_18575,N_13732,N_14194);
nor U18576 (N_18576,N_12359,N_14252);
or U18577 (N_18577,N_12887,N_10135);
nor U18578 (N_18578,N_14206,N_14682);
and U18579 (N_18579,N_10058,N_11708);
or U18580 (N_18580,N_14930,N_13498);
nand U18581 (N_18581,N_10771,N_13627);
or U18582 (N_18582,N_11009,N_14299);
and U18583 (N_18583,N_14788,N_12483);
nand U18584 (N_18584,N_13641,N_11681);
or U18585 (N_18585,N_10530,N_12941);
and U18586 (N_18586,N_10642,N_11564);
nand U18587 (N_18587,N_11224,N_10446);
and U18588 (N_18588,N_14819,N_14606);
or U18589 (N_18589,N_10162,N_10545);
or U18590 (N_18590,N_11905,N_12397);
nand U18591 (N_18591,N_12116,N_10911);
nand U18592 (N_18592,N_10299,N_13585);
and U18593 (N_18593,N_14041,N_10495);
nand U18594 (N_18594,N_13603,N_12455);
nand U18595 (N_18595,N_10605,N_12157);
nand U18596 (N_18596,N_12246,N_10021);
nand U18597 (N_18597,N_12061,N_10171);
and U18598 (N_18598,N_10731,N_10638);
nand U18599 (N_18599,N_12681,N_10445);
nand U18600 (N_18600,N_14300,N_12781);
or U18601 (N_18601,N_14244,N_10220);
nor U18602 (N_18602,N_11243,N_13120);
and U18603 (N_18603,N_14665,N_14013);
or U18604 (N_18604,N_11756,N_14949);
or U18605 (N_18605,N_10644,N_10143);
and U18606 (N_18606,N_12830,N_11505);
or U18607 (N_18607,N_11328,N_13363);
nor U18608 (N_18608,N_10129,N_12641);
or U18609 (N_18609,N_10465,N_13820);
and U18610 (N_18610,N_12838,N_12434);
nor U18611 (N_18611,N_12578,N_13381);
or U18612 (N_18612,N_13837,N_10421);
nor U18613 (N_18613,N_12734,N_12263);
and U18614 (N_18614,N_11433,N_13056);
nor U18615 (N_18615,N_14027,N_14391);
and U18616 (N_18616,N_13308,N_12801);
or U18617 (N_18617,N_14599,N_12568);
and U18618 (N_18618,N_11242,N_12999);
or U18619 (N_18619,N_12033,N_11555);
nand U18620 (N_18620,N_11729,N_11323);
nor U18621 (N_18621,N_12704,N_10301);
nand U18622 (N_18622,N_11593,N_11560);
nor U18623 (N_18623,N_13524,N_13963);
and U18624 (N_18624,N_14491,N_12380);
nor U18625 (N_18625,N_12653,N_14570);
nand U18626 (N_18626,N_11456,N_10851);
or U18627 (N_18627,N_13963,N_12852);
nor U18628 (N_18628,N_10590,N_14892);
and U18629 (N_18629,N_13950,N_12216);
and U18630 (N_18630,N_13342,N_10661);
nor U18631 (N_18631,N_11712,N_11626);
nand U18632 (N_18632,N_14804,N_14260);
nand U18633 (N_18633,N_10702,N_12480);
nand U18634 (N_18634,N_11960,N_13328);
nor U18635 (N_18635,N_10381,N_13627);
and U18636 (N_18636,N_14928,N_11786);
nand U18637 (N_18637,N_10162,N_13680);
and U18638 (N_18638,N_11266,N_10506);
and U18639 (N_18639,N_14654,N_13808);
nand U18640 (N_18640,N_10676,N_10723);
and U18641 (N_18641,N_11812,N_10190);
nor U18642 (N_18642,N_12974,N_11724);
or U18643 (N_18643,N_10256,N_10598);
xor U18644 (N_18644,N_12074,N_11833);
nor U18645 (N_18645,N_14989,N_13147);
nor U18646 (N_18646,N_10189,N_11327);
nand U18647 (N_18647,N_14017,N_14755);
or U18648 (N_18648,N_10899,N_12105);
or U18649 (N_18649,N_13532,N_10418);
and U18650 (N_18650,N_13983,N_13343);
and U18651 (N_18651,N_10407,N_14589);
nand U18652 (N_18652,N_14646,N_13292);
and U18653 (N_18653,N_12513,N_13890);
and U18654 (N_18654,N_14513,N_14778);
or U18655 (N_18655,N_11655,N_11257);
nor U18656 (N_18656,N_11322,N_10877);
and U18657 (N_18657,N_10775,N_10159);
or U18658 (N_18658,N_14018,N_11770);
and U18659 (N_18659,N_14842,N_11921);
nor U18660 (N_18660,N_14485,N_14657);
or U18661 (N_18661,N_13051,N_10260);
nor U18662 (N_18662,N_10611,N_14231);
and U18663 (N_18663,N_13318,N_12640);
nand U18664 (N_18664,N_12241,N_12140);
and U18665 (N_18665,N_12284,N_14414);
nand U18666 (N_18666,N_10525,N_12756);
nand U18667 (N_18667,N_11393,N_14963);
and U18668 (N_18668,N_13979,N_11606);
or U18669 (N_18669,N_12496,N_12523);
nand U18670 (N_18670,N_11524,N_11410);
or U18671 (N_18671,N_12142,N_10432);
nor U18672 (N_18672,N_11843,N_11344);
and U18673 (N_18673,N_12404,N_12139);
and U18674 (N_18674,N_11699,N_13150);
or U18675 (N_18675,N_14810,N_12882);
nand U18676 (N_18676,N_13261,N_11651);
nand U18677 (N_18677,N_10769,N_12463);
nor U18678 (N_18678,N_10273,N_10781);
or U18679 (N_18679,N_12453,N_14885);
nor U18680 (N_18680,N_14849,N_11916);
and U18681 (N_18681,N_10466,N_13849);
or U18682 (N_18682,N_14899,N_11623);
nor U18683 (N_18683,N_11399,N_13471);
and U18684 (N_18684,N_11836,N_12658);
and U18685 (N_18685,N_13445,N_12124);
or U18686 (N_18686,N_14430,N_10955);
or U18687 (N_18687,N_12841,N_10188);
nand U18688 (N_18688,N_10395,N_12663);
or U18689 (N_18689,N_10569,N_12815);
nand U18690 (N_18690,N_13306,N_12143);
nor U18691 (N_18691,N_11342,N_11780);
nand U18692 (N_18692,N_13783,N_12608);
nand U18693 (N_18693,N_12063,N_13614);
or U18694 (N_18694,N_10658,N_12572);
and U18695 (N_18695,N_11638,N_13670);
or U18696 (N_18696,N_11524,N_12310);
and U18697 (N_18697,N_14040,N_12544);
and U18698 (N_18698,N_10937,N_11421);
and U18699 (N_18699,N_14589,N_11912);
or U18700 (N_18700,N_11116,N_10771);
and U18701 (N_18701,N_12504,N_12885);
or U18702 (N_18702,N_14645,N_13744);
nor U18703 (N_18703,N_11441,N_12890);
nor U18704 (N_18704,N_13462,N_13935);
nor U18705 (N_18705,N_12831,N_11530);
and U18706 (N_18706,N_12218,N_14456);
or U18707 (N_18707,N_10125,N_12450);
nand U18708 (N_18708,N_11446,N_12900);
nor U18709 (N_18709,N_14155,N_12308);
and U18710 (N_18710,N_11149,N_11797);
and U18711 (N_18711,N_10119,N_11599);
or U18712 (N_18712,N_14274,N_13759);
nand U18713 (N_18713,N_11088,N_10694);
nor U18714 (N_18714,N_14630,N_11353);
nor U18715 (N_18715,N_10951,N_13306);
and U18716 (N_18716,N_13939,N_12635);
or U18717 (N_18717,N_12819,N_11366);
or U18718 (N_18718,N_14606,N_12247);
and U18719 (N_18719,N_10177,N_10228);
and U18720 (N_18720,N_10564,N_10535);
and U18721 (N_18721,N_10333,N_12368);
nor U18722 (N_18722,N_10705,N_10076);
or U18723 (N_18723,N_10334,N_12563);
and U18724 (N_18724,N_13246,N_12722);
or U18725 (N_18725,N_11936,N_10616);
and U18726 (N_18726,N_11126,N_13574);
or U18727 (N_18727,N_14242,N_11219);
and U18728 (N_18728,N_14939,N_14046);
nand U18729 (N_18729,N_13630,N_11209);
nand U18730 (N_18730,N_10134,N_11625);
and U18731 (N_18731,N_11910,N_13777);
nand U18732 (N_18732,N_14063,N_11786);
nand U18733 (N_18733,N_13336,N_11011);
nor U18734 (N_18734,N_14799,N_13789);
and U18735 (N_18735,N_11523,N_12151);
and U18736 (N_18736,N_10641,N_10909);
or U18737 (N_18737,N_12797,N_10924);
nand U18738 (N_18738,N_14727,N_12867);
and U18739 (N_18739,N_11605,N_14994);
nand U18740 (N_18740,N_13581,N_14884);
and U18741 (N_18741,N_14932,N_12009);
nand U18742 (N_18742,N_13739,N_14997);
and U18743 (N_18743,N_10376,N_12638);
nor U18744 (N_18744,N_14104,N_10714);
nand U18745 (N_18745,N_11984,N_14099);
or U18746 (N_18746,N_12430,N_12089);
and U18747 (N_18747,N_13531,N_14802);
nor U18748 (N_18748,N_12384,N_11260);
and U18749 (N_18749,N_14359,N_12898);
nor U18750 (N_18750,N_11998,N_10307);
nor U18751 (N_18751,N_14611,N_12443);
nor U18752 (N_18752,N_14464,N_11211);
and U18753 (N_18753,N_11267,N_11730);
nand U18754 (N_18754,N_14293,N_11696);
or U18755 (N_18755,N_13448,N_10020);
nor U18756 (N_18756,N_10680,N_11318);
xor U18757 (N_18757,N_13595,N_13618);
and U18758 (N_18758,N_12926,N_11787);
nand U18759 (N_18759,N_14257,N_11511);
and U18760 (N_18760,N_11913,N_11416);
or U18761 (N_18761,N_10171,N_14773);
and U18762 (N_18762,N_14336,N_14445);
nand U18763 (N_18763,N_10138,N_14454);
or U18764 (N_18764,N_14446,N_13018);
and U18765 (N_18765,N_14509,N_10535);
nand U18766 (N_18766,N_13371,N_10838);
nand U18767 (N_18767,N_12969,N_13254);
or U18768 (N_18768,N_13741,N_10292);
and U18769 (N_18769,N_13990,N_11319);
or U18770 (N_18770,N_13991,N_10347);
or U18771 (N_18771,N_12696,N_10317);
and U18772 (N_18772,N_10866,N_14472);
and U18773 (N_18773,N_14357,N_10875);
nor U18774 (N_18774,N_11055,N_13151);
or U18775 (N_18775,N_13478,N_12780);
or U18776 (N_18776,N_12829,N_11445);
xnor U18777 (N_18777,N_11445,N_10008);
nand U18778 (N_18778,N_12972,N_11119);
or U18779 (N_18779,N_14808,N_13914);
or U18780 (N_18780,N_11293,N_12136);
nand U18781 (N_18781,N_14607,N_12771);
and U18782 (N_18782,N_14240,N_13376);
nand U18783 (N_18783,N_13359,N_13822);
nand U18784 (N_18784,N_11046,N_14958);
or U18785 (N_18785,N_10149,N_13090);
nor U18786 (N_18786,N_13718,N_10747);
nand U18787 (N_18787,N_14700,N_14303);
or U18788 (N_18788,N_10198,N_13754);
or U18789 (N_18789,N_14112,N_11575);
or U18790 (N_18790,N_11888,N_14200);
nor U18791 (N_18791,N_13389,N_10559);
and U18792 (N_18792,N_12692,N_11448);
nand U18793 (N_18793,N_10459,N_13184);
or U18794 (N_18794,N_10418,N_10314);
or U18795 (N_18795,N_10400,N_11272);
nor U18796 (N_18796,N_11327,N_12899);
nor U18797 (N_18797,N_14148,N_11383);
nand U18798 (N_18798,N_12509,N_10889);
nand U18799 (N_18799,N_10860,N_14336);
nor U18800 (N_18800,N_13370,N_12470);
or U18801 (N_18801,N_10051,N_13294);
and U18802 (N_18802,N_12973,N_11592);
or U18803 (N_18803,N_11179,N_13744);
nand U18804 (N_18804,N_13068,N_13414);
nor U18805 (N_18805,N_10952,N_12798);
and U18806 (N_18806,N_10310,N_11821);
and U18807 (N_18807,N_14627,N_10478);
nor U18808 (N_18808,N_14714,N_12118);
or U18809 (N_18809,N_11431,N_14860);
nand U18810 (N_18810,N_13687,N_13228);
nand U18811 (N_18811,N_14037,N_10966);
and U18812 (N_18812,N_12608,N_10419);
nor U18813 (N_18813,N_11265,N_13227);
and U18814 (N_18814,N_14253,N_14836);
nand U18815 (N_18815,N_11525,N_10687);
or U18816 (N_18816,N_14039,N_14287);
nor U18817 (N_18817,N_14293,N_10410);
and U18818 (N_18818,N_10448,N_12769);
or U18819 (N_18819,N_11345,N_12284);
nor U18820 (N_18820,N_12864,N_13441);
or U18821 (N_18821,N_12736,N_14302);
or U18822 (N_18822,N_12926,N_12412);
nand U18823 (N_18823,N_13977,N_14886);
and U18824 (N_18824,N_11257,N_11089);
nor U18825 (N_18825,N_12055,N_13699);
or U18826 (N_18826,N_14934,N_14072);
nor U18827 (N_18827,N_14876,N_14422);
nor U18828 (N_18828,N_14447,N_12083);
nor U18829 (N_18829,N_11413,N_12912);
nand U18830 (N_18830,N_13804,N_14906);
nor U18831 (N_18831,N_11830,N_14566);
nor U18832 (N_18832,N_13249,N_10546);
nand U18833 (N_18833,N_10646,N_11924);
and U18834 (N_18834,N_11791,N_12083);
nand U18835 (N_18835,N_14065,N_12496);
nor U18836 (N_18836,N_13967,N_12835);
nor U18837 (N_18837,N_10921,N_11579);
and U18838 (N_18838,N_14788,N_14919);
or U18839 (N_18839,N_14578,N_11393);
and U18840 (N_18840,N_10265,N_13940);
nor U18841 (N_18841,N_10639,N_11107);
and U18842 (N_18842,N_14605,N_12209);
nor U18843 (N_18843,N_12026,N_14939);
nor U18844 (N_18844,N_13328,N_13418);
or U18845 (N_18845,N_12780,N_13598);
nor U18846 (N_18846,N_14165,N_12016);
and U18847 (N_18847,N_12320,N_10044);
and U18848 (N_18848,N_10549,N_11164);
or U18849 (N_18849,N_10744,N_12302);
nand U18850 (N_18850,N_13531,N_12293);
nand U18851 (N_18851,N_10776,N_14259);
and U18852 (N_18852,N_12244,N_14379);
and U18853 (N_18853,N_10110,N_12665);
and U18854 (N_18854,N_12392,N_11096);
nand U18855 (N_18855,N_11222,N_10871);
nand U18856 (N_18856,N_12983,N_12413);
or U18857 (N_18857,N_10710,N_13580);
or U18858 (N_18858,N_12236,N_11266);
and U18859 (N_18859,N_11315,N_14607);
nor U18860 (N_18860,N_10851,N_11503);
nor U18861 (N_18861,N_13882,N_10959);
xnor U18862 (N_18862,N_12603,N_13258);
xnor U18863 (N_18863,N_12616,N_14021);
nand U18864 (N_18864,N_13622,N_10338);
or U18865 (N_18865,N_14585,N_11910);
nand U18866 (N_18866,N_11006,N_10957);
nand U18867 (N_18867,N_11129,N_11469);
nand U18868 (N_18868,N_13659,N_10327);
and U18869 (N_18869,N_14874,N_14417);
nor U18870 (N_18870,N_11278,N_13724);
nor U18871 (N_18871,N_12286,N_14168);
and U18872 (N_18872,N_14180,N_14480);
nor U18873 (N_18873,N_13362,N_10943);
nor U18874 (N_18874,N_13430,N_13132);
nor U18875 (N_18875,N_12568,N_12606);
xnor U18876 (N_18876,N_14029,N_11434);
and U18877 (N_18877,N_12866,N_10176);
nand U18878 (N_18878,N_13856,N_13748);
nor U18879 (N_18879,N_13439,N_12874);
nor U18880 (N_18880,N_10603,N_11173);
nand U18881 (N_18881,N_10617,N_12663);
nor U18882 (N_18882,N_14112,N_13037);
and U18883 (N_18883,N_10751,N_10144);
or U18884 (N_18884,N_10695,N_14731);
nor U18885 (N_18885,N_11128,N_13358);
and U18886 (N_18886,N_14515,N_12524);
or U18887 (N_18887,N_11961,N_12524);
and U18888 (N_18888,N_13093,N_14908);
or U18889 (N_18889,N_13737,N_13754);
or U18890 (N_18890,N_12023,N_12427);
or U18891 (N_18891,N_13321,N_14476);
or U18892 (N_18892,N_11446,N_14652);
nand U18893 (N_18893,N_11154,N_14369);
and U18894 (N_18894,N_11235,N_11660);
and U18895 (N_18895,N_14909,N_12685);
nor U18896 (N_18896,N_11134,N_11607);
and U18897 (N_18897,N_11379,N_12772);
or U18898 (N_18898,N_14337,N_13126);
and U18899 (N_18899,N_12144,N_10167);
nand U18900 (N_18900,N_12134,N_14915);
nor U18901 (N_18901,N_10695,N_11275);
and U18902 (N_18902,N_11454,N_13404);
and U18903 (N_18903,N_12038,N_14650);
and U18904 (N_18904,N_12057,N_13911);
or U18905 (N_18905,N_14590,N_13500);
nor U18906 (N_18906,N_13582,N_11217);
nor U18907 (N_18907,N_10080,N_11173);
and U18908 (N_18908,N_14634,N_12422);
and U18909 (N_18909,N_11570,N_14138);
nor U18910 (N_18910,N_12837,N_14928);
and U18911 (N_18911,N_11553,N_13532);
or U18912 (N_18912,N_13025,N_10664);
or U18913 (N_18913,N_13952,N_10912);
and U18914 (N_18914,N_14441,N_14987);
nand U18915 (N_18915,N_13023,N_14270);
or U18916 (N_18916,N_13893,N_10015);
and U18917 (N_18917,N_10359,N_10263);
and U18918 (N_18918,N_12170,N_11955);
and U18919 (N_18919,N_13382,N_10118);
nor U18920 (N_18920,N_13568,N_10925);
and U18921 (N_18921,N_11829,N_10326);
or U18922 (N_18922,N_10156,N_14708);
and U18923 (N_18923,N_10893,N_11108);
and U18924 (N_18924,N_12650,N_14497);
or U18925 (N_18925,N_11375,N_11845);
and U18926 (N_18926,N_11761,N_11379);
nand U18927 (N_18927,N_10245,N_14998);
xnor U18928 (N_18928,N_14511,N_14026);
or U18929 (N_18929,N_11129,N_12610);
nand U18930 (N_18930,N_10348,N_13375);
nor U18931 (N_18931,N_14118,N_11809);
or U18932 (N_18932,N_10643,N_11459);
nor U18933 (N_18933,N_11332,N_14611);
nor U18934 (N_18934,N_14106,N_12705);
or U18935 (N_18935,N_11061,N_13988);
or U18936 (N_18936,N_10591,N_10658);
or U18937 (N_18937,N_10884,N_12155);
nand U18938 (N_18938,N_12085,N_12644);
or U18939 (N_18939,N_13198,N_10387);
and U18940 (N_18940,N_10623,N_13461);
nor U18941 (N_18941,N_10236,N_13390);
nand U18942 (N_18942,N_13564,N_13220);
nand U18943 (N_18943,N_12700,N_14068);
nor U18944 (N_18944,N_12834,N_13863);
and U18945 (N_18945,N_12968,N_10667);
nor U18946 (N_18946,N_10870,N_14361);
or U18947 (N_18947,N_11659,N_13210);
and U18948 (N_18948,N_10817,N_11887);
nand U18949 (N_18949,N_14832,N_12766);
nand U18950 (N_18950,N_10815,N_12149);
or U18951 (N_18951,N_13092,N_13571);
nor U18952 (N_18952,N_12461,N_12422);
nor U18953 (N_18953,N_13909,N_13361);
or U18954 (N_18954,N_13868,N_14669);
or U18955 (N_18955,N_13879,N_10267);
nor U18956 (N_18956,N_10460,N_13873);
and U18957 (N_18957,N_11115,N_12986);
nor U18958 (N_18958,N_14838,N_12634);
nand U18959 (N_18959,N_13015,N_10782);
or U18960 (N_18960,N_14420,N_12966);
or U18961 (N_18961,N_12465,N_13850);
nor U18962 (N_18962,N_11546,N_10523);
nand U18963 (N_18963,N_12497,N_13748);
xnor U18964 (N_18964,N_12199,N_11850);
and U18965 (N_18965,N_13600,N_12594);
or U18966 (N_18966,N_12006,N_13444);
nor U18967 (N_18967,N_10175,N_13029);
and U18968 (N_18968,N_10739,N_14488);
or U18969 (N_18969,N_13820,N_11954);
or U18970 (N_18970,N_10526,N_13703);
and U18971 (N_18971,N_11780,N_12863);
nand U18972 (N_18972,N_14357,N_14358);
or U18973 (N_18973,N_11775,N_12861);
or U18974 (N_18974,N_11712,N_12990);
nor U18975 (N_18975,N_10914,N_13871);
and U18976 (N_18976,N_14076,N_14187);
or U18977 (N_18977,N_12959,N_14505);
nor U18978 (N_18978,N_10682,N_10585);
nand U18979 (N_18979,N_11317,N_10386);
or U18980 (N_18980,N_12785,N_10801);
nand U18981 (N_18981,N_12503,N_11304);
nor U18982 (N_18982,N_14798,N_10228);
nand U18983 (N_18983,N_14886,N_12577);
or U18984 (N_18984,N_10536,N_10856);
and U18985 (N_18985,N_10626,N_11582);
nand U18986 (N_18986,N_11032,N_10909);
and U18987 (N_18987,N_13380,N_14143);
or U18988 (N_18988,N_10507,N_13135);
and U18989 (N_18989,N_11086,N_12578);
and U18990 (N_18990,N_11065,N_13967);
nand U18991 (N_18991,N_11861,N_10331);
and U18992 (N_18992,N_10080,N_10166);
and U18993 (N_18993,N_11241,N_11859);
nor U18994 (N_18994,N_14382,N_11155);
or U18995 (N_18995,N_11730,N_13496);
and U18996 (N_18996,N_10388,N_12320);
and U18997 (N_18997,N_11003,N_10779);
or U18998 (N_18998,N_11621,N_13625);
or U18999 (N_18999,N_12874,N_12065);
nor U19000 (N_19000,N_11159,N_11375);
xnor U19001 (N_19001,N_13733,N_11397);
and U19002 (N_19002,N_13385,N_10869);
nor U19003 (N_19003,N_12073,N_10978);
or U19004 (N_19004,N_10298,N_10290);
and U19005 (N_19005,N_10112,N_12731);
nor U19006 (N_19006,N_12554,N_13424);
nand U19007 (N_19007,N_13502,N_12751);
nor U19008 (N_19008,N_12090,N_13097);
nor U19009 (N_19009,N_13447,N_13227);
or U19010 (N_19010,N_12357,N_13869);
and U19011 (N_19011,N_11278,N_12247);
or U19012 (N_19012,N_12765,N_10876);
or U19013 (N_19013,N_14049,N_14792);
nor U19014 (N_19014,N_13936,N_14051);
or U19015 (N_19015,N_11309,N_14704);
or U19016 (N_19016,N_14716,N_12280);
nor U19017 (N_19017,N_12176,N_14896);
nor U19018 (N_19018,N_13501,N_13273);
and U19019 (N_19019,N_10811,N_12820);
or U19020 (N_19020,N_14820,N_10527);
or U19021 (N_19021,N_10901,N_11358);
and U19022 (N_19022,N_11799,N_14446);
nand U19023 (N_19023,N_10149,N_10524);
nor U19024 (N_19024,N_11779,N_13804);
nor U19025 (N_19025,N_10076,N_14645);
and U19026 (N_19026,N_10137,N_11694);
nor U19027 (N_19027,N_11868,N_11429);
and U19028 (N_19028,N_13051,N_14371);
and U19029 (N_19029,N_10942,N_10630);
or U19030 (N_19030,N_12834,N_14943);
or U19031 (N_19031,N_11730,N_14162);
nand U19032 (N_19032,N_14037,N_12644);
and U19033 (N_19033,N_14084,N_12140);
and U19034 (N_19034,N_12991,N_10947);
or U19035 (N_19035,N_13321,N_12942);
nor U19036 (N_19036,N_12218,N_11650);
or U19037 (N_19037,N_13907,N_14695);
and U19038 (N_19038,N_10266,N_13472);
nand U19039 (N_19039,N_10370,N_13794);
nor U19040 (N_19040,N_11864,N_11782);
or U19041 (N_19041,N_10358,N_14775);
nor U19042 (N_19042,N_11652,N_10877);
nor U19043 (N_19043,N_12032,N_14518);
or U19044 (N_19044,N_14045,N_12359);
nand U19045 (N_19045,N_12307,N_13664);
xor U19046 (N_19046,N_12350,N_13697);
and U19047 (N_19047,N_14408,N_10337);
and U19048 (N_19048,N_10752,N_10793);
nand U19049 (N_19049,N_12939,N_13021);
and U19050 (N_19050,N_11435,N_11061);
nand U19051 (N_19051,N_10657,N_12898);
nand U19052 (N_19052,N_10564,N_10187);
nand U19053 (N_19053,N_11168,N_12981);
xor U19054 (N_19054,N_12707,N_11112);
or U19055 (N_19055,N_12548,N_13801);
or U19056 (N_19056,N_13679,N_10993);
nand U19057 (N_19057,N_11984,N_11891);
nor U19058 (N_19058,N_13018,N_10063);
or U19059 (N_19059,N_13148,N_13053);
or U19060 (N_19060,N_10481,N_11676);
nor U19061 (N_19061,N_11945,N_14878);
and U19062 (N_19062,N_14882,N_11011);
nand U19063 (N_19063,N_13877,N_14092);
nor U19064 (N_19064,N_13948,N_13474);
and U19065 (N_19065,N_11824,N_11835);
or U19066 (N_19066,N_10232,N_12960);
or U19067 (N_19067,N_12375,N_14465);
nor U19068 (N_19068,N_10622,N_10379);
or U19069 (N_19069,N_12706,N_12136);
nor U19070 (N_19070,N_14653,N_13560);
or U19071 (N_19071,N_11625,N_12072);
and U19072 (N_19072,N_14807,N_12836);
and U19073 (N_19073,N_13238,N_14433);
nor U19074 (N_19074,N_10053,N_12401);
nor U19075 (N_19075,N_13957,N_10165);
or U19076 (N_19076,N_13120,N_11592);
and U19077 (N_19077,N_12790,N_13046);
nand U19078 (N_19078,N_10521,N_11520);
nor U19079 (N_19079,N_14657,N_12305);
nand U19080 (N_19080,N_11522,N_12508);
and U19081 (N_19081,N_13730,N_14158);
or U19082 (N_19082,N_14723,N_12531);
nor U19083 (N_19083,N_14217,N_11201);
and U19084 (N_19084,N_11783,N_13931);
nor U19085 (N_19085,N_10154,N_14438);
nor U19086 (N_19086,N_12482,N_13947);
nand U19087 (N_19087,N_12646,N_14631);
and U19088 (N_19088,N_13762,N_14310);
nand U19089 (N_19089,N_10646,N_10990);
nor U19090 (N_19090,N_11407,N_14702);
nand U19091 (N_19091,N_10536,N_13034);
nor U19092 (N_19092,N_10612,N_11939);
and U19093 (N_19093,N_13966,N_10632);
nand U19094 (N_19094,N_14266,N_14879);
nor U19095 (N_19095,N_10664,N_14152);
or U19096 (N_19096,N_12849,N_12799);
nand U19097 (N_19097,N_10395,N_12967);
and U19098 (N_19098,N_11184,N_13361);
or U19099 (N_19099,N_11077,N_10030);
nand U19100 (N_19100,N_10459,N_11771);
or U19101 (N_19101,N_10201,N_11199);
or U19102 (N_19102,N_14648,N_14095);
nor U19103 (N_19103,N_14291,N_13237);
and U19104 (N_19104,N_10276,N_12396);
nor U19105 (N_19105,N_14490,N_13582);
or U19106 (N_19106,N_13325,N_11086);
xnor U19107 (N_19107,N_13971,N_11714);
and U19108 (N_19108,N_14966,N_12917);
or U19109 (N_19109,N_13785,N_11748);
nor U19110 (N_19110,N_11463,N_12530);
nand U19111 (N_19111,N_13119,N_12046);
and U19112 (N_19112,N_14505,N_13061);
nand U19113 (N_19113,N_11579,N_11823);
nor U19114 (N_19114,N_13361,N_13826);
or U19115 (N_19115,N_10806,N_12362);
nand U19116 (N_19116,N_14305,N_10565);
or U19117 (N_19117,N_12945,N_13510);
and U19118 (N_19118,N_13508,N_10426);
and U19119 (N_19119,N_14674,N_14576);
nand U19120 (N_19120,N_11940,N_10031);
and U19121 (N_19121,N_10853,N_13048);
or U19122 (N_19122,N_11713,N_11323);
nand U19123 (N_19123,N_14839,N_14899);
and U19124 (N_19124,N_12839,N_11511);
and U19125 (N_19125,N_13238,N_14620);
or U19126 (N_19126,N_14190,N_13634);
and U19127 (N_19127,N_10155,N_10667);
or U19128 (N_19128,N_11813,N_10157);
nor U19129 (N_19129,N_14600,N_11259);
nand U19130 (N_19130,N_14723,N_11110);
or U19131 (N_19131,N_12259,N_11625);
nor U19132 (N_19132,N_12507,N_11714);
nor U19133 (N_19133,N_12414,N_12729);
and U19134 (N_19134,N_12674,N_13175);
or U19135 (N_19135,N_12077,N_10985);
nor U19136 (N_19136,N_10101,N_14198);
nand U19137 (N_19137,N_12685,N_14669);
nand U19138 (N_19138,N_13186,N_10782);
nor U19139 (N_19139,N_10126,N_14875);
nor U19140 (N_19140,N_13340,N_10983);
nor U19141 (N_19141,N_13216,N_13964);
or U19142 (N_19142,N_12859,N_11623);
and U19143 (N_19143,N_13539,N_14964);
nand U19144 (N_19144,N_10834,N_13448);
nor U19145 (N_19145,N_10640,N_14399);
nor U19146 (N_19146,N_14156,N_11003);
nand U19147 (N_19147,N_12621,N_11790);
nor U19148 (N_19148,N_13829,N_14749);
nor U19149 (N_19149,N_11520,N_12047);
or U19150 (N_19150,N_14315,N_12594);
or U19151 (N_19151,N_10125,N_10983);
nor U19152 (N_19152,N_12807,N_11685);
nor U19153 (N_19153,N_11991,N_13396);
nor U19154 (N_19154,N_13899,N_13220);
and U19155 (N_19155,N_10140,N_10571);
or U19156 (N_19156,N_10543,N_14364);
and U19157 (N_19157,N_11151,N_10942);
or U19158 (N_19158,N_13080,N_12657);
and U19159 (N_19159,N_10495,N_10514);
nor U19160 (N_19160,N_14414,N_13070);
nor U19161 (N_19161,N_10142,N_13020);
nor U19162 (N_19162,N_13884,N_14099);
or U19163 (N_19163,N_14306,N_12416);
nand U19164 (N_19164,N_13376,N_11054);
or U19165 (N_19165,N_12460,N_11442);
nand U19166 (N_19166,N_12238,N_14079);
nand U19167 (N_19167,N_10034,N_13273);
and U19168 (N_19168,N_13830,N_13903);
nand U19169 (N_19169,N_13185,N_12384);
or U19170 (N_19170,N_13252,N_10174);
nand U19171 (N_19171,N_14161,N_12621);
or U19172 (N_19172,N_14588,N_12196);
nor U19173 (N_19173,N_13231,N_14871);
or U19174 (N_19174,N_10327,N_12781);
and U19175 (N_19175,N_12478,N_14644);
nor U19176 (N_19176,N_11449,N_12759);
nor U19177 (N_19177,N_14447,N_13864);
nor U19178 (N_19178,N_14157,N_11370);
or U19179 (N_19179,N_14440,N_10475);
nor U19180 (N_19180,N_14956,N_10828);
and U19181 (N_19181,N_12704,N_14766);
or U19182 (N_19182,N_11970,N_12874);
and U19183 (N_19183,N_14612,N_13748);
and U19184 (N_19184,N_10414,N_12512);
or U19185 (N_19185,N_11930,N_13709);
nand U19186 (N_19186,N_14390,N_10226);
nand U19187 (N_19187,N_11765,N_12945);
nand U19188 (N_19188,N_14838,N_10043);
or U19189 (N_19189,N_13440,N_11867);
and U19190 (N_19190,N_12848,N_10316);
nor U19191 (N_19191,N_11202,N_14289);
nor U19192 (N_19192,N_13141,N_11173);
or U19193 (N_19193,N_14756,N_11884);
and U19194 (N_19194,N_12360,N_11200);
and U19195 (N_19195,N_11599,N_13524);
nor U19196 (N_19196,N_13814,N_10013);
or U19197 (N_19197,N_14600,N_11079);
nand U19198 (N_19198,N_11836,N_11908);
or U19199 (N_19199,N_14156,N_11008);
nor U19200 (N_19200,N_12294,N_10951);
nor U19201 (N_19201,N_14284,N_12221);
or U19202 (N_19202,N_10465,N_14392);
nor U19203 (N_19203,N_12933,N_10015);
and U19204 (N_19204,N_13750,N_14912);
or U19205 (N_19205,N_13409,N_11271);
and U19206 (N_19206,N_10007,N_11310);
and U19207 (N_19207,N_10703,N_14304);
or U19208 (N_19208,N_12782,N_14151);
nand U19209 (N_19209,N_11390,N_13334);
nand U19210 (N_19210,N_12071,N_10528);
nor U19211 (N_19211,N_12001,N_10018);
or U19212 (N_19212,N_13461,N_10139);
nand U19213 (N_19213,N_11613,N_11980);
nor U19214 (N_19214,N_12290,N_13852);
or U19215 (N_19215,N_10894,N_12951);
nor U19216 (N_19216,N_12341,N_14393);
nand U19217 (N_19217,N_11290,N_11348);
or U19218 (N_19218,N_12380,N_12305);
nand U19219 (N_19219,N_10264,N_11897);
and U19220 (N_19220,N_12986,N_10905);
nand U19221 (N_19221,N_14109,N_14246);
and U19222 (N_19222,N_12173,N_13775);
nor U19223 (N_19223,N_12721,N_11504);
nand U19224 (N_19224,N_11804,N_10984);
nand U19225 (N_19225,N_11498,N_10121);
nand U19226 (N_19226,N_11181,N_13686);
nand U19227 (N_19227,N_11747,N_11312);
or U19228 (N_19228,N_14824,N_13313);
nand U19229 (N_19229,N_13944,N_10694);
nor U19230 (N_19230,N_11884,N_12932);
nor U19231 (N_19231,N_13948,N_12836);
nand U19232 (N_19232,N_11633,N_12896);
nor U19233 (N_19233,N_12038,N_11322);
or U19234 (N_19234,N_11372,N_12410);
nor U19235 (N_19235,N_14986,N_12680);
or U19236 (N_19236,N_11617,N_10366);
and U19237 (N_19237,N_12607,N_10172);
and U19238 (N_19238,N_11140,N_11747);
nor U19239 (N_19239,N_11075,N_11974);
nor U19240 (N_19240,N_10740,N_10630);
and U19241 (N_19241,N_12791,N_13434);
nor U19242 (N_19242,N_13386,N_12155);
nand U19243 (N_19243,N_10639,N_14322);
nand U19244 (N_19244,N_14239,N_11302);
and U19245 (N_19245,N_14060,N_14775);
nand U19246 (N_19246,N_11451,N_14959);
nor U19247 (N_19247,N_14817,N_14096);
nand U19248 (N_19248,N_12052,N_11437);
or U19249 (N_19249,N_13892,N_11086);
nor U19250 (N_19250,N_14166,N_10667);
nand U19251 (N_19251,N_11361,N_11384);
nand U19252 (N_19252,N_10157,N_14798);
and U19253 (N_19253,N_13007,N_10900);
and U19254 (N_19254,N_13709,N_10122);
nor U19255 (N_19255,N_11717,N_11059);
or U19256 (N_19256,N_12468,N_13476);
and U19257 (N_19257,N_12266,N_11495);
and U19258 (N_19258,N_13788,N_10814);
nor U19259 (N_19259,N_11211,N_13927);
nor U19260 (N_19260,N_14270,N_13782);
nand U19261 (N_19261,N_12054,N_14550);
and U19262 (N_19262,N_14234,N_13735);
and U19263 (N_19263,N_11782,N_13564);
and U19264 (N_19264,N_12045,N_13907);
and U19265 (N_19265,N_13145,N_12755);
nor U19266 (N_19266,N_13953,N_12511);
and U19267 (N_19267,N_13881,N_12901);
and U19268 (N_19268,N_12933,N_11680);
nand U19269 (N_19269,N_12860,N_13020);
or U19270 (N_19270,N_13154,N_11257);
and U19271 (N_19271,N_13513,N_13137);
nor U19272 (N_19272,N_13719,N_10539);
nand U19273 (N_19273,N_11762,N_13083);
and U19274 (N_19274,N_11427,N_11289);
or U19275 (N_19275,N_10381,N_10930);
and U19276 (N_19276,N_11609,N_13573);
or U19277 (N_19277,N_12721,N_12754);
and U19278 (N_19278,N_14856,N_10738);
nor U19279 (N_19279,N_11226,N_10475);
or U19280 (N_19280,N_11380,N_14162);
nand U19281 (N_19281,N_14090,N_13763);
nor U19282 (N_19282,N_10760,N_12694);
and U19283 (N_19283,N_12448,N_10950);
nand U19284 (N_19284,N_14617,N_11227);
nand U19285 (N_19285,N_11947,N_12772);
nor U19286 (N_19286,N_12509,N_14473);
and U19287 (N_19287,N_12016,N_13360);
nor U19288 (N_19288,N_13766,N_11974);
nor U19289 (N_19289,N_13575,N_13537);
or U19290 (N_19290,N_12376,N_11197);
or U19291 (N_19291,N_13242,N_11494);
or U19292 (N_19292,N_14329,N_12036);
or U19293 (N_19293,N_12273,N_14793);
or U19294 (N_19294,N_12385,N_11380);
or U19295 (N_19295,N_10240,N_14812);
nor U19296 (N_19296,N_10080,N_11185);
or U19297 (N_19297,N_12872,N_11872);
and U19298 (N_19298,N_11600,N_10682);
nor U19299 (N_19299,N_12001,N_13787);
or U19300 (N_19300,N_13473,N_11924);
nor U19301 (N_19301,N_13289,N_11667);
nand U19302 (N_19302,N_10109,N_11765);
nand U19303 (N_19303,N_13337,N_11741);
or U19304 (N_19304,N_13146,N_10926);
nand U19305 (N_19305,N_11359,N_11141);
nand U19306 (N_19306,N_13254,N_14542);
nand U19307 (N_19307,N_14129,N_14207);
nand U19308 (N_19308,N_10980,N_10581);
and U19309 (N_19309,N_10237,N_11290);
nor U19310 (N_19310,N_13830,N_10740);
and U19311 (N_19311,N_13313,N_14041);
and U19312 (N_19312,N_11240,N_10635);
nand U19313 (N_19313,N_12802,N_13434);
and U19314 (N_19314,N_14506,N_10001);
nor U19315 (N_19315,N_12430,N_10254);
nand U19316 (N_19316,N_12846,N_14340);
nor U19317 (N_19317,N_13498,N_11260);
nor U19318 (N_19318,N_12418,N_13253);
nor U19319 (N_19319,N_13161,N_10513);
nand U19320 (N_19320,N_13032,N_13025);
nor U19321 (N_19321,N_11449,N_14969);
nand U19322 (N_19322,N_10774,N_12609);
or U19323 (N_19323,N_11966,N_11169);
and U19324 (N_19324,N_13061,N_12430);
or U19325 (N_19325,N_11795,N_12634);
nor U19326 (N_19326,N_13573,N_14493);
nand U19327 (N_19327,N_14738,N_12159);
nor U19328 (N_19328,N_10698,N_10930);
or U19329 (N_19329,N_12912,N_12879);
nand U19330 (N_19330,N_11333,N_11820);
or U19331 (N_19331,N_10693,N_10012);
and U19332 (N_19332,N_11954,N_12084);
or U19333 (N_19333,N_12457,N_14088);
nor U19334 (N_19334,N_12216,N_14898);
nand U19335 (N_19335,N_11214,N_14536);
and U19336 (N_19336,N_10791,N_10090);
or U19337 (N_19337,N_14640,N_11521);
and U19338 (N_19338,N_12804,N_12851);
nand U19339 (N_19339,N_14796,N_14228);
nor U19340 (N_19340,N_14910,N_12325);
or U19341 (N_19341,N_14553,N_14899);
nor U19342 (N_19342,N_12930,N_14688);
nor U19343 (N_19343,N_14441,N_11383);
and U19344 (N_19344,N_14357,N_14680);
nor U19345 (N_19345,N_13314,N_14576);
or U19346 (N_19346,N_11180,N_10747);
nand U19347 (N_19347,N_10011,N_14508);
xnor U19348 (N_19348,N_11058,N_14544);
xor U19349 (N_19349,N_12540,N_14263);
or U19350 (N_19350,N_13800,N_14515);
or U19351 (N_19351,N_12985,N_14355);
or U19352 (N_19352,N_13222,N_13406);
and U19353 (N_19353,N_14006,N_13193);
nor U19354 (N_19354,N_12161,N_13130);
nor U19355 (N_19355,N_11572,N_11539);
nand U19356 (N_19356,N_14999,N_12856);
xor U19357 (N_19357,N_12037,N_10450);
or U19358 (N_19358,N_12626,N_10288);
nand U19359 (N_19359,N_10488,N_11175);
and U19360 (N_19360,N_10267,N_14982);
nor U19361 (N_19361,N_10701,N_12179);
nand U19362 (N_19362,N_10107,N_10016);
nor U19363 (N_19363,N_14359,N_14733);
or U19364 (N_19364,N_10940,N_14977);
nand U19365 (N_19365,N_13912,N_14121);
nor U19366 (N_19366,N_11856,N_14271);
or U19367 (N_19367,N_14540,N_13338);
or U19368 (N_19368,N_11555,N_11729);
nor U19369 (N_19369,N_10188,N_11603);
nand U19370 (N_19370,N_10569,N_12241);
and U19371 (N_19371,N_12833,N_12343);
nand U19372 (N_19372,N_13304,N_12401);
nor U19373 (N_19373,N_11509,N_10317);
and U19374 (N_19374,N_10038,N_14203);
and U19375 (N_19375,N_13698,N_10658);
or U19376 (N_19376,N_13800,N_10963);
nor U19377 (N_19377,N_12766,N_14070);
or U19378 (N_19378,N_11065,N_14215);
or U19379 (N_19379,N_12969,N_11807);
and U19380 (N_19380,N_11863,N_11580);
and U19381 (N_19381,N_12471,N_11334);
xnor U19382 (N_19382,N_13606,N_13648);
or U19383 (N_19383,N_12973,N_11230);
and U19384 (N_19384,N_14222,N_12083);
nor U19385 (N_19385,N_13712,N_12457);
and U19386 (N_19386,N_12730,N_10191);
nand U19387 (N_19387,N_14709,N_11534);
nand U19388 (N_19388,N_10929,N_11446);
and U19389 (N_19389,N_11398,N_14140);
or U19390 (N_19390,N_12078,N_12761);
or U19391 (N_19391,N_11137,N_12314);
and U19392 (N_19392,N_12104,N_14231);
and U19393 (N_19393,N_10332,N_14194);
or U19394 (N_19394,N_10168,N_12636);
or U19395 (N_19395,N_13584,N_11861);
nor U19396 (N_19396,N_11463,N_13912);
and U19397 (N_19397,N_10668,N_14414);
nand U19398 (N_19398,N_13535,N_12319);
and U19399 (N_19399,N_12064,N_12986);
and U19400 (N_19400,N_13026,N_12217);
and U19401 (N_19401,N_12237,N_10613);
nand U19402 (N_19402,N_10036,N_14015);
nor U19403 (N_19403,N_11376,N_14009);
and U19404 (N_19404,N_11272,N_11880);
nor U19405 (N_19405,N_10870,N_12381);
or U19406 (N_19406,N_10562,N_12663);
nand U19407 (N_19407,N_13495,N_14521);
or U19408 (N_19408,N_10876,N_11612);
or U19409 (N_19409,N_14911,N_12784);
and U19410 (N_19410,N_14208,N_12162);
nor U19411 (N_19411,N_10366,N_14452);
nand U19412 (N_19412,N_14392,N_12474);
nor U19413 (N_19413,N_11942,N_11683);
and U19414 (N_19414,N_10157,N_12083);
or U19415 (N_19415,N_13845,N_12233);
or U19416 (N_19416,N_13969,N_14201);
nor U19417 (N_19417,N_14220,N_14059);
or U19418 (N_19418,N_11330,N_13829);
nor U19419 (N_19419,N_14237,N_10509);
or U19420 (N_19420,N_13200,N_13098);
and U19421 (N_19421,N_14768,N_13352);
nor U19422 (N_19422,N_13601,N_11578);
nand U19423 (N_19423,N_10825,N_13589);
nand U19424 (N_19424,N_10883,N_14534);
nor U19425 (N_19425,N_12279,N_10934);
or U19426 (N_19426,N_10652,N_11918);
or U19427 (N_19427,N_13958,N_11368);
and U19428 (N_19428,N_14829,N_14914);
xor U19429 (N_19429,N_10689,N_11189);
nand U19430 (N_19430,N_12367,N_12977);
nor U19431 (N_19431,N_14804,N_14587);
nand U19432 (N_19432,N_12586,N_11178);
and U19433 (N_19433,N_13621,N_13231);
nor U19434 (N_19434,N_13960,N_14099);
and U19435 (N_19435,N_10614,N_13305);
and U19436 (N_19436,N_14586,N_11723);
and U19437 (N_19437,N_14736,N_13372);
or U19438 (N_19438,N_14354,N_11490);
nand U19439 (N_19439,N_12704,N_10612);
and U19440 (N_19440,N_12003,N_13707);
nand U19441 (N_19441,N_14382,N_11630);
nand U19442 (N_19442,N_12863,N_12919);
nor U19443 (N_19443,N_13637,N_13514);
nor U19444 (N_19444,N_13414,N_14368);
or U19445 (N_19445,N_12219,N_10117);
nand U19446 (N_19446,N_13473,N_13539);
nand U19447 (N_19447,N_13692,N_10692);
nand U19448 (N_19448,N_14298,N_12306);
xor U19449 (N_19449,N_12763,N_11270);
and U19450 (N_19450,N_10298,N_10470);
and U19451 (N_19451,N_10587,N_12796);
or U19452 (N_19452,N_11608,N_13410);
nand U19453 (N_19453,N_12395,N_10981);
or U19454 (N_19454,N_13485,N_11961);
nor U19455 (N_19455,N_13251,N_11800);
or U19456 (N_19456,N_10169,N_14763);
nor U19457 (N_19457,N_13290,N_13092);
nor U19458 (N_19458,N_10767,N_14170);
and U19459 (N_19459,N_13826,N_11233);
nor U19460 (N_19460,N_13513,N_13200);
nand U19461 (N_19461,N_13718,N_14619);
nand U19462 (N_19462,N_14698,N_14522);
nand U19463 (N_19463,N_13579,N_14873);
or U19464 (N_19464,N_14317,N_12678);
and U19465 (N_19465,N_12782,N_10594);
xor U19466 (N_19466,N_14552,N_14596);
or U19467 (N_19467,N_10688,N_14094);
or U19468 (N_19468,N_11646,N_13307);
or U19469 (N_19469,N_14233,N_11849);
nand U19470 (N_19470,N_10212,N_12567);
nor U19471 (N_19471,N_14609,N_12007);
nand U19472 (N_19472,N_10817,N_13098);
nor U19473 (N_19473,N_11160,N_10199);
xor U19474 (N_19474,N_12891,N_10728);
and U19475 (N_19475,N_11894,N_10332);
nand U19476 (N_19476,N_13378,N_10099);
nor U19477 (N_19477,N_14614,N_10112);
and U19478 (N_19478,N_14963,N_11425);
nand U19479 (N_19479,N_13563,N_13501);
nand U19480 (N_19480,N_12210,N_11396);
and U19481 (N_19481,N_13792,N_13666);
nand U19482 (N_19482,N_14267,N_14912);
or U19483 (N_19483,N_14043,N_11771);
or U19484 (N_19484,N_13563,N_12207);
or U19485 (N_19485,N_12954,N_13285);
nand U19486 (N_19486,N_10666,N_12435);
or U19487 (N_19487,N_13064,N_11147);
and U19488 (N_19488,N_12498,N_12819);
nand U19489 (N_19489,N_12700,N_12535);
or U19490 (N_19490,N_13571,N_12519);
and U19491 (N_19491,N_12372,N_11729);
nor U19492 (N_19492,N_13164,N_13187);
xor U19493 (N_19493,N_14163,N_14727);
nand U19494 (N_19494,N_14689,N_12276);
and U19495 (N_19495,N_11784,N_12211);
or U19496 (N_19496,N_13137,N_14381);
nand U19497 (N_19497,N_12047,N_13650);
nand U19498 (N_19498,N_12936,N_13078);
nand U19499 (N_19499,N_13827,N_11904);
or U19500 (N_19500,N_13486,N_11536);
nor U19501 (N_19501,N_14499,N_12437);
nand U19502 (N_19502,N_12987,N_11723);
nor U19503 (N_19503,N_12529,N_11413);
nor U19504 (N_19504,N_10677,N_13094);
nand U19505 (N_19505,N_14938,N_12446);
or U19506 (N_19506,N_10715,N_14312);
and U19507 (N_19507,N_10627,N_12059);
nor U19508 (N_19508,N_13357,N_13082);
and U19509 (N_19509,N_10638,N_13203);
and U19510 (N_19510,N_12739,N_13034);
nand U19511 (N_19511,N_10487,N_13857);
or U19512 (N_19512,N_12086,N_12356);
and U19513 (N_19513,N_12350,N_10039);
nand U19514 (N_19514,N_10441,N_10493);
nand U19515 (N_19515,N_13483,N_11140);
nor U19516 (N_19516,N_11376,N_13971);
nand U19517 (N_19517,N_13892,N_10621);
nor U19518 (N_19518,N_10583,N_12730);
and U19519 (N_19519,N_13601,N_12315);
nand U19520 (N_19520,N_11005,N_12514);
nor U19521 (N_19521,N_13629,N_12944);
and U19522 (N_19522,N_14065,N_13830);
and U19523 (N_19523,N_13491,N_11582);
nor U19524 (N_19524,N_11273,N_12762);
nor U19525 (N_19525,N_12465,N_10751);
or U19526 (N_19526,N_14663,N_14207);
nand U19527 (N_19527,N_14682,N_11628);
nor U19528 (N_19528,N_11095,N_11867);
nand U19529 (N_19529,N_13721,N_11812);
and U19530 (N_19530,N_14391,N_12484);
nand U19531 (N_19531,N_12664,N_11154);
or U19532 (N_19532,N_13555,N_14037);
nand U19533 (N_19533,N_10943,N_12953);
nor U19534 (N_19534,N_11533,N_12524);
and U19535 (N_19535,N_11557,N_12810);
nand U19536 (N_19536,N_11714,N_13948);
nor U19537 (N_19537,N_10604,N_14592);
and U19538 (N_19538,N_14220,N_14281);
and U19539 (N_19539,N_14303,N_13473);
and U19540 (N_19540,N_11535,N_11721);
or U19541 (N_19541,N_10033,N_12939);
or U19542 (N_19542,N_11452,N_11483);
nand U19543 (N_19543,N_10689,N_10405);
or U19544 (N_19544,N_12170,N_12770);
or U19545 (N_19545,N_11538,N_10082);
or U19546 (N_19546,N_13386,N_13476);
and U19547 (N_19547,N_13604,N_11617);
and U19548 (N_19548,N_12659,N_13206);
or U19549 (N_19549,N_11210,N_12960);
and U19550 (N_19550,N_12854,N_14946);
and U19551 (N_19551,N_10369,N_11572);
nand U19552 (N_19552,N_10907,N_11001);
and U19553 (N_19553,N_10713,N_12452);
and U19554 (N_19554,N_13444,N_10064);
nand U19555 (N_19555,N_10596,N_10071);
and U19556 (N_19556,N_12080,N_13460);
nor U19557 (N_19557,N_11761,N_10522);
nor U19558 (N_19558,N_11380,N_10959);
or U19559 (N_19559,N_11362,N_11315);
nand U19560 (N_19560,N_11431,N_14178);
or U19561 (N_19561,N_11803,N_13164);
nor U19562 (N_19562,N_10666,N_11910);
nor U19563 (N_19563,N_10228,N_11470);
nand U19564 (N_19564,N_11212,N_13674);
nand U19565 (N_19565,N_13447,N_13695);
or U19566 (N_19566,N_14834,N_13919);
or U19567 (N_19567,N_10421,N_13447);
nor U19568 (N_19568,N_11903,N_11837);
and U19569 (N_19569,N_11772,N_10021);
and U19570 (N_19570,N_12719,N_11550);
or U19571 (N_19571,N_10002,N_14743);
nor U19572 (N_19572,N_11015,N_14339);
nor U19573 (N_19573,N_14658,N_10810);
nand U19574 (N_19574,N_14387,N_12287);
or U19575 (N_19575,N_12480,N_13713);
and U19576 (N_19576,N_14061,N_11509);
nand U19577 (N_19577,N_11641,N_12199);
xor U19578 (N_19578,N_13301,N_12209);
or U19579 (N_19579,N_13285,N_12029);
and U19580 (N_19580,N_10093,N_12983);
nand U19581 (N_19581,N_11029,N_12098);
and U19582 (N_19582,N_14682,N_14976);
and U19583 (N_19583,N_14479,N_14221);
nand U19584 (N_19584,N_11484,N_14314);
or U19585 (N_19585,N_10169,N_14210);
nor U19586 (N_19586,N_13603,N_11969);
nand U19587 (N_19587,N_12683,N_12424);
nand U19588 (N_19588,N_11109,N_12696);
nand U19589 (N_19589,N_14535,N_12781);
or U19590 (N_19590,N_11256,N_13279);
or U19591 (N_19591,N_13658,N_12342);
nor U19592 (N_19592,N_14808,N_12963);
nand U19593 (N_19593,N_11568,N_10659);
nor U19594 (N_19594,N_11949,N_13040);
and U19595 (N_19595,N_12434,N_10703);
nor U19596 (N_19596,N_10037,N_12578);
nor U19597 (N_19597,N_12149,N_14583);
or U19598 (N_19598,N_11143,N_14801);
nand U19599 (N_19599,N_12429,N_11166);
or U19600 (N_19600,N_13527,N_12282);
and U19601 (N_19601,N_14827,N_14059);
nor U19602 (N_19602,N_10056,N_14642);
and U19603 (N_19603,N_13128,N_12402);
nand U19604 (N_19604,N_13471,N_10821);
and U19605 (N_19605,N_10371,N_13957);
nand U19606 (N_19606,N_10067,N_13366);
nor U19607 (N_19607,N_10055,N_10615);
nand U19608 (N_19608,N_13573,N_14024);
and U19609 (N_19609,N_12238,N_10932);
nand U19610 (N_19610,N_14184,N_11655);
nor U19611 (N_19611,N_14091,N_13816);
nor U19612 (N_19612,N_13893,N_13925);
nand U19613 (N_19613,N_11841,N_13240);
or U19614 (N_19614,N_12734,N_12516);
nor U19615 (N_19615,N_14700,N_12698);
nand U19616 (N_19616,N_12995,N_14281);
or U19617 (N_19617,N_12173,N_10116);
or U19618 (N_19618,N_10330,N_11880);
nor U19619 (N_19619,N_10392,N_12744);
and U19620 (N_19620,N_12232,N_13137);
nor U19621 (N_19621,N_14165,N_14836);
or U19622 (N_19622,N_13230,N_10927);
xor U19623 (N_19623,N_11251,N_13639);
nor U19624 (N_19624,N_14970,N_13492);
nand U19625 (N_19625,N_12709,N_13655);
nor U19626 (N_19626,N_14503,N_11804);
and U19627 (N_19627,N_13036,N_12381);
and U19628 (N_19628,N_14963,N_12970);
and U19629 (N_19629,N_14495,N_12787);
nand U19630 (N_19630,N_13558,N_12305);
nor U19631 (N_19631,N_11377,N_14601);
and U19632 (N_19632,N_12625,N_13603);
nor U19633 (N_19633,N_11342,N_13887);
or U19634 (N_19634,N_12619,N_11213);
xor U19635 (N_19635,N_12488,N_12401);
nand U19636 (N_19636,N_13249,N_11675);
nor U19637 (N_19637,N_11468,N_13170);
nand U19638 (N_19638,N_10714,N_13628);
nor U19639 (N_19639,N_14803,N_11449);
nor U19640 (N_19640,N_14820,N_11515);
and U19641 (N_19641,N_13933,N_14520);
or U19642 (N_19642,N_13959,N_13574);
and U19643 (N_19643,N_11626,N_11047);
nand U19644 (N_19644,N_13050,N_13629);
and U19645 (N_19645,N_10284,N_12555);
nor U19646 (N_19646,N_12616,N_13206);
or U19647 (N_19647,N_11478,N_14729);
nand U19648 (N_19648,N_13203,N_14089);
and U19649 (N_19649,N_12569,N_11774);
or U19650 (N_19650,N_14329,N_10709);
and U19651 (N_19651,N_11942,N_14504);
nor U19652 (N_19652,N_10038,N_11705);
nor U19653 (N_19653,N_13332,N_12654);
nor U19654 (N_19654,N_10986,N_14187);
nand U19655 (N_19655,N_12280,N_11443);
nor U19656 (N_19656,N_12550,N_12959);
or U19657 (N_19657,N_13338,N_11571);
or U19658 (N_19658,N_13170,N_13979);
and U19659 (N_19659,N_10728,N_10819);
nand U19660 (N_19660,N_12291,N_12119);
and U19661 (N_19661,N_14733,N_11615);
and U19662 (N_19662,N_11979,N_11265);
nor U19663 (N_19663,N_12677,N_11364);
nor U19664 (N_19664,N_12074,N_10568);
or U19665 (N_19665,N_12745,N_10380);
and U19666 (N_19666,N_11223,N_10359);
nor U19667 (N_19667,N_12186,N_10833);
nand U19668 (N_19668,N_14100,N_14107);
and U19669 (N_19669,N_14380,N_11083);
or U19670 (N_19670,N_14722,N_10379);
nor U19671 (N_19671,N_14883,N_12260);
and U19672 (N_19672,N_11768,N_11733);
nor U19673 (N_19673,N_14661,N_14053);
and U19674 (N_19674,N_14330,N_14608);
nor U19675 (N_19675,N_14844,N_12136);
nand U19676 (N_19676,N_12276,N_10821);
nor U19677 (N_19677,N_13731,N_12555);
or U19678 (N_19678,N_11752,N_13443);
and U19679 (N_19679,N_12141,N_12069);
or U19680 (N_19680,N_10980,N_10412);
nor U19681 (N_19681,N_10154,N_10854);
nor U19682 (N_19682,N_14515,N_14224);
nor U19683 (N_19683,N_10635,N_12253);
or U19684 (N_19684,N_10548,N_12007);
nand U19685 (N_19685,N_11459,N_10942);
nor U19686 (N_19686,N_10850,N_13030);
and U19687 (N_19687,N_13760,N_10062);
and U19688 (N_19688,N_14401,N_12354);
and U19689 (N_19689,N_12692,N_11659);
and U19690 (N_19690,N_14115,N_12769);
or U19691 (N_19691,N_14627,N_13669);
nor U19692 (N_19692,N_11690,N_10908);
or U19693 (N_19693,N_11547,N_14947);
or U19694 (N_19694,N_13778,N_12733);
and U19695 (N_19695,N_11464,N_14611);
nor U19696 (N_19696,N_14799,N_10457);
or U19697 (N_19697,N_12411,N_12340);
nor U19698 (N_19698,N_14451,N_12105);
or U19699 (N_19699,N_13567,N_11606);
or U19700 (N_19700,N_10185,N_13131);
or U19701 (N_19701,N_12716,N_12131);
nor U19702 (N_19702,N_14432,N_10673);
nand U19703 (N_19703,N_12600,N_10257);
and U19704 (N_19704,N_12497,N_10754);
and U19705 (N_19705,N_10966,N_14632);
xor U19706 (N_19706,N_12274,N_13947);
and U19707 (N_19707,N_11712,N_12531);
and U19708 (N_19708,N_11032,N_13053);
nand U19709 (N_19709,N_10202,N_14917);
nor U19710 (N_19710,N_12051,N_11263);
and U19711 (N_19711,N_12075,N_14659);
nand U19712 (N_19712,N_10457,N_11982);
and U19713 (N_19713,N_11934,N_11763);
nand U19714 (N_19714,N_12370,N_13518);
and U19715 (N_19715,N_10864,N_14027);
and U19716 (N_19716,N_11120,N_13782);
or U19717 (N_19717,N_13720,N_14113);
and U19718 (N_19718,N_12370,N_11625);
and U19719 (N_19719,N_13550,N_12876);
or U19720 (N_19720,N_12115,N_12202);
and U19721 (N_19721,N_13010,N_12493);
nand U19722 (N_19722,N_10324,N_14929);
and U19723 (N_19723,N_10365,N_12875);
nor U19724 (N_19724,N_13489,N_11791);
and U19725 (N_19725,N_10039,N_13648);
and U19726 (N_19726,N_14365,N_10263);
or U19727 (N_19727,N_12446,N_12501);
or U19728 (N_19728,N_10828,N_14827);
nor U19729 (N_19729,N_10892,N_11630);
or U19730 (N_19730,N_14230,N_10295);
and U19731 (N_19731,N_14668,N_12526);
and U19732 (N_19732,N_13762,N_12791);
nand U19733 (N_19733,N_10979,N_10894);
nand U19734 (N_19734,N_14329,N_11213);
nand U19735 (N_19735,N_11188,N_10515);
nor U19736 (N_19736,N_14981,N_13634);
and U19737 (N_19737,N_12151,N_14743);
and U19738 (N_19738,N_10069,N_14291);
nor U19739 (N_19739,N_14651,N_10986);
or U19740 (N_19740,N_14840,N_14117);
and U19741 (N_19741,N_10575,N_13385);
or U19742 (N_19742,N_10558,N_11535);
and U19743 (N_19743,N_12388,N_13688);
nor U19744 (N_19744,N_14388,N_14223);
xnor U19745 (N_19745,N_12976,N_12989);
or U19746 (N_19746,N_12781,N_14711);
or U19747 (N_19747,N_11524,N_13364);
or U19748 (N_19748,N_12810,N_10280);
and U19749 (N_19749,N_10235,N_10841);
and U19750 (N_19750,N_14990,N_13411);
and U19751 (N_19751,N_10926,N_14424);
nand U19752 (N_19752,N_11074,N_12265);
or U19753 (N_19753,N_12049,N_12468);
nor U19754 (N_19754,N_11503,N_10931);
and U19755 (N_19755,N_10067,N_13159);
or U19756 (N_19756,N_11396,N_11983);
xnor U19757 (N_19757,N_12226,N_14664);
nor U19758 (N_19758,N_14546,N_11511);
nor U19759 (N_19759,N_12029,N_10884);
nand U19760 (N_19760,N_12054,N_14753);
or U19761 (N_19761,N_10553,N_12689);
or U19762 (N_19762,N_10015,N_10004);
nand U19763 (N_19763,N_10558,N_12658);
and U19764 (N_19764,N_14741,N_11444);
or U19765 (N_19765,N_11447,N_12775);
nor U19766 (N_19766,N_12647,N_11296);
nand U19767 (N_19767,N_10146,N_10369);
nand U19768 (N_19768,N_13557,N_14782);
or U19769 (N_19769,N_13072,N_11397);
or U19770 (N_19770,N_10894,N_13064);
nor U19771 (N_19771,N_14355,N_13249);
and U19772 (N_19772,N_13695,N_12752);
and U19773 (N_19773,N_12400,N_10698);
nor U19774 (N_19774,N_11540,N_10158);
nor U19775 (N_19775,N_13789,N_14570);
nand U19776 (N_19776,N_11849,N_11086);
or U19777 (N_19777,N_10242,N_12781);
nand U19778 (N_19778,N_10898,N_14388);
or U19779 (N_19779,N_13694,N_13195);
nor U19780 (N_19780,N_13953,N_12128);
nor U19781 (N_19781,N_10002,N_12104);
nor U19782 (N_19782,N_11577,N_11822);
or U19783 (N_19783,N_13961,N_11232);
and U19784 (N_19784,N_10306,N_13868);
nand U19785 (N_19785,N_10422,N_14776);
nor U19786 (N_19786,N_13789,N_14387);
and U19787 (N_19787,N_14125,N_13925);
nor U19788 (N_19788,N_11466,N_11082);
or U19789 (N_19789,N_13271,N_14657);
and U19790 (N_19790,N_14677,N_13491);
nor U19791 (N_19791,N_11023,N_10532);
nor U19792 (N_19792,N_11881,N_14278);
or U19793 (N_19793,N_14240,N_14506);
or U19794 (N_19794,N_12557,N_13157);
nor U19795 (N_19795,N_11521,N_14305);
nand U19796 (N_19796,N_14684,N_11584);
or U19797 (N_19797,N_14684,N_12127);
nand U19798 (N_19798,N_12991,N_13040);
nand U19799 (N_19799,N_12482,N_11702);
nand U19800 (N_19800,N_13733,N_12773);
nor U19801 (N_19801,N_11932,N_13434);
and U19802 (N_19802,N_14839,N_13667);
or U19803 (N_19803,N_10593,N_14661);
or U19804 (N_19804,N_10014,N_13708);
or U19805 (N_19805,N_13661,N_14648);
or U19806 (N_19806,N_10994,N_12357);
nor U19807 (N_19807,N_11292,N_13092);
and U19808 (N_19808,N_13250,N_14440);
or U19809 (N_19809,N_13566,N_12530);
nand U19810 (N_19810,N_10558,N_10378);
nor U19811 (N_19811,N_12061,N_11864);
or U19812 (N_19812,N_13310,N_13357);
or U19813 (N_19813,N_14220,N_10658);
nor U19814 (N_19814,N_14048,N_12532);
nand U19815 (N_19815,N_12586,N_13763);
and U19816 (N_19816,N_10161,N_12090);
xnor U19817 (N_19817,N_13640,N_10539);
nor U19818 (N_19818,N_11845,N_10318);
nand U19819 (N_19819,N_11546,N_10442);
nand U19820 (N_19820,N_11743,N_13587);
nor U19821 (N_19821,N_13757,N_12311);
or U19822 (N_19822,N_13629,N_13182);
nor U19823 (N_19823,N_13425,N_12246);
nand U19824 (N_19824,N_11875,N_10943);
nand U19825 (N_19825,N_10203,N_12515);
or U19826 (N_19826,N_13299,N_14033);
and U19827 (N_19827,N_11384,N_10704);
and U19828 (N_19828,N_12467,N_10934);
nand U19829 (N_19829,N_11820,N_10699);
or U19830 (N_19830,N_12682,N_11804);
and U19831 (N_19831,N_10565,N_11722);
nor U19832 (N_19832,N_12739,N_14891);
and U19833 (N_19833,N_14665,N_10964);
nand U19834 (N_19834,N_13769,N_12475);
or U19835 (N_19835,N_10479,N_14253);
nor U19836 (N_19836,N_11578,N_10160);
and U19837 (N_19837,N_10624,N_12260);
nand U19838 (N_19838,N_11280,N_12151);
nor U19839 (N_19839,N_10677,N_14133);
or U19840 (N_19840,N_13480,N_11016);
nor U19841 (N_19841,N_12274,N_10437);
nor U19842 (N_19842,N_12451,N_12302);
nor U19843 (N_19843,N_13305,N_10207);
nor U19844 (N_19844,N_13367,N_14342);
or U19845 (N_19845,N_14324,N_10124);
nor U19846 (N_19846,N_10793,N_11844);
or U19847 (N_19847,N_11566,N_12980);
nor U19848 (N_19848,N_14324,N_11914);
nand U19849 (N_19849,N_12253,N_10448);
nor U19850 (N_19850,N_14616,N_11438);
or U19851 (N_19851,N_14332,N_10664);
nor U19852 (N_19852,N_10560,N_14041);
or U19853 (N_19853,N_12360,N_14617);
or U19854 (N_19854,N_10418,N_13271);
nor U19855 (N_19855,N_11103,N_11967);
and U19856 (N_19856,N_13231,N_13369);
or U19857 (N_19857,N_13845,N_10479);
nand U19858 (N_19858,N_10694,N_11394);
nand U19859 (N_19859,N_10244,N_12986);
nor U19860 (N_19860,N_11212,N_14839);
or U19861 (N_19861,N_11006,N_13163);
nand U19862 (N_19862,N_12238,N_12543);
nor U19863 (N_19863,N_14281,N_14157);
and U19864 (N_19864,N_14518,N_10664);
and U19865 (N_19865,N_12771,N_11344);
nor U19866 (N_19866,N_10031,N_13917);
or U19867 (N_19867,N_11545,N_14941);
and U19868 (N_19868,N_14988,N_11541);
or U19869 (N_19869,N_10319,N_10885);
nor U19870 (N_19870,N_12186,N_11006);
nand U19871 (N_19871,N_10885,N_11722);
nand U19872 (N_19872,N_14531,N_10948);
or U19873 (N_19873,N_10388,N_10191);
or U19874 (N_19874,N_11745,N_14639);
or U19875 (N_19875,N_10900,N_11276);
nor U19876 (N_19876,N_14090,N_10675);
nor U19877 (N_19877,N_14240,N_13783);
nor U19878 (N_19878,N_11169,N_14989);
and U19879 (N_19879,N_10847,N_14818);
and U19880 (N_19880,N_14233,N_13088);
and U19881 (N_19881,N_10558,N_14367);
nand U19882 (N_19882,N_12456,N_13037);
or U19883 (N_19883,N_13876,N_10643);
nor U19884 (N_19884,N_10173,N_11688);
nand U19885 (N_19885,N_13251,N_14383);
and U19886 (N_19886,N_13990,N_10984);
nor U19887 (N_19887,N_13088,N_12293);
xor U19888 (N_19888,N_11239,N_11545);
or U19889 (N_19889,N_14431,N_12363);
nand U19890 (N_19890,N_12427,N_14003);
nor U19891 (N_19891,N_14613,N_12010);
nor U19892 (N_19892,N_13161,N_14153);
or U19893 (N_19893,N_12188,N_10364);
or U19894 (N_19894,N_13165,N_10746);
or U19895 (N_19895,N_13703,N_13641);
or U19896 (N_19896,N_12194,N_11563);
nand U19897 (N_19897,N_13551,N_12108);
and U19898 (N_19898,N_12314,N_11016);
nor U19899 (N_19899,N_14434,N_14841);
nor U19900 (N_19900,N_12645,N_13344);
nand U19901 (N_19901,N_12172,N_11942);
nand U19902 (N_19902,N_11470,N_10713);
or U19903 (N_19903,N_12874,N_11283);
nand U19904 (N_19904,N_11353,N_14529);
nor U19905 (N_19905,N_13331,N_10966);
and U19906 (N_19906,N_13388,N_13484);
nor U19907 (N_19907,N_14643,N_13823);
and U19908 (N_19908,N_12591,N_14027);
nand U19909 (N_19909,N_10552,N_10943);
and U19910 (N_19910,N_14101,N_14215);
nor U19911 (N_19911,N_14194,N_10582);
nand U19912 (N_19912,N_11676,N_10647);
or U19913 (N_19913,N_10366,N_14466);
and U19914 (N_19914,N_10259,N_13815);
and U19915 (N_19915,N_14427,N_12542);
nand U19916 (N_19916,N_10621,N_10037);
nor U19917 (N_19917,N_14865,N_12099);
or U19918 (N_19918,N_13295,N_11982);
and U19919 (N_19919,N_14283,N_12117);
and U19920 (N_19920,N_14067,N_10328);
nand U19921 (N_19921,N_11283,N_13112);
and U19922 (N_19922,N_11775,N_14050);
and U19923 (N_19923,N_13271,N_10897);
nand U19924 (N_19924,N_10849,N_11805);
and U19925 (N_19925,N_11475,N_11895);
nor U19926 (N_19926,N_13869,N_14973);
nand U19927 (N_19927,N_10842,N_11596);
or U19928 (N_19928,N_14333,N_14683);
and U19929 (N_19929,N_10282,N_14762);
or U19930 (N_19930,N_14034,N_11832);
xor U19931 (N_19931,N_14120,N_10548);
nand U19932 (N_19932,N_13171,N_13534);
nand U19933 (N_19933,N_13214,N_13835);
or U19934 (N_19934,N_11115,N_10624);
or U19935 (N_19935,N_10836,N_13586);
nand U19936 (N_19936,N_14923,N_11354);
nor U19937 (N_19937,N_13858,N_11163);
or U19938 (N_19938,N_10755,N_14422);
nand U19939 (N_19939,N_10217,N_11649);
and U19940 (N_19940,N_10329,N_11302);
and U19941 (N_19941,N_13537,N_10835);
and U19942 (N_19942,N_14466,N_11613);
nor U19943 (N_19943,N_13408,N_10888);
nor U19944 (N_19944,N_13465,N_13455);
nor U19945 (N_19945,N_12125,N_13444);
nand U19946 (N_19946,N_12719,N_13133);
and U19947 (N_19947,N_13116,N_12328);
nand U19948 (N_19948,N_14822,N_12902);
nor U19949 (N_19949,N_12389,N_11827);
xnor U19950 (N_19950,N_11531,N_12237);
nand U19951 (N_19951,N_11622,N_11202);
nor U19952 (N_19952,N_12705,N_11327);
nor U19953 (N_19953,N_14108,N_11153);
and U19954 (N_19954,N_10353,N_11639);
or U19955 (N_19955,N_10394,N_14956);
nor U19956 (N_19956,N_13845,N_13897);
nor U19957 (N_19957,N_12277,N_11138);
nor U19958 (N_19958,N_11398,N_12146);
and U19959 (N_19959,N_10997,N_10631);
or U19960 (N_19960,N_12823,N_10768);
or U19961 (N_19961,N_10410,N_13010);
nor U19962 (N_19962,N_10547,N_14895);
nor U19963 (N_19963,N_13912,N_11540);
and U19964 (N_19964,N_11957,N_14226);
nand U19965 (N_19965,N_13932,N_14081);
or U19966 (N_19966,N_11334,N_14776);
and U19967 (N_19967,N_13661,N_10191);
or U19968 (N_19968,N_14515,N_13439);
nand U19969 (N_19969,N_10215,N_11414);
xor U19970 (N_19970,N_11371,N_10653);
nand U19971 (N_19971,N_12582,N_11332);
nor U19972 (N_19972,N_11164,N_14835);
nor U19973 (N_19973,N_14118,N_13052);
and U19974 (N_19974,N_12297,N_10723);
or U19975 (N_19975,N_13512,N_11864);
and U19976 (N_19976,N_14823,N_11466);
and U19977 (N_19977,N_10528,N_10257);
nand U19978 (N_19978,N_11633,N_12707);
or U19979 (N_19979,N_12426,N_14460);
nand U19980 (N_19980,N_14247,N_12871);
nor U19981 (N_19981,N_10785,N_10957);
and U19982 (N_19982,N_14219,N_11076);
nand U19983 (N_19983,N_11586,N_12174);
nand U19984 (N_19984,N_12641,N_14718);
nand U19985 (N_19985,N_14561,N_10702);
nor U19986 (N_19986,N_13825,N_14278);
and U19987 (N_19987,N_12355,N_14005);
or U19988 (N_19988,N_11641,N_11957);
nand U19989 (N_19989,N_10341,N_13772);
or U19990 (N_19990,N_11905,N_10412);
or U19991 (N_19991,N_12818,N_10254);
and U19992 (N_19992,N_11303,N_13689);
nand U19993 (N_19993,N_14604,N_13419);
nand U19994 (N_19994,N_10976,N_13320);
and U19995 (N_19995,N_12462,N_14617);
and U19996 (N_19996,N_12067,N_13308);
nor U19997 (N_19997,N_11501,N_11002);
xor U19998 (N_19998,N_10547,N_12209);
or U19999 (N_19999,N_11881,N_13038);
and UO_0 (O_0,N_16166,N_19547);
or UO_1 (O_1,N_17411,N_18438);
nor UO_2 (O_2,N_15113,N_16686);
nand UO_3 (O_3,N_19853,N_19552);
xor UO_4 (O_4,N_16910,N_19063);
nand UO_5 (O_5,N_17407,N_15410);
nor UO_6 (O_6,N_17768,N_19215);
nor UO_7 (O_7,N_19868,N_18663);
nand UO_8 (O_8,N_19869,N_15609);
or UO_9 (O_9,N_17646,N_17020);
nor UO_10 (O_10,N_16491,N_15623);
and UO_11 (O_11,N_19298,N_15455);
or UO_12 (O_12,N_16704,N_18932);
or UO_13 (O_13,N_15786,N_19747);
or UO_14 (O_14,N_16307,N_19536);
nor UO_15 (O_15,N_17729,N_15327);
nor UO_16 (O_16,N_16474,N_16794);
and UO_17 (O_17,N_18300,N_18521);
or UO_18 (O_18,N_17555,N_18775);
nor UO_19 (O_19,N_18449,N_15453);
or UO_20 (O_20,N_16104,N_18713);
and UO_21 (O_21,N_16636,N_19583);
nor UO_22 (O_22,N_15395,N_15776);
nor UO_23 (O_23,N_19566,N_19144);
and UO_24 (O_24,N_15350,N_15583);
xnor UO_25 (O_25,N_17224,N_15662);
nand UO_26 (O_26,N_16162,N_15529);
and UO_27 (O_27,N_15899,N_19703);
and UO_28 (O_28,N_18804,N_18689);
and UO_29 (O_29,N_16368,N_17711);
nand UO_30 (O_30,N_19730,N_18532);
and UO_31 (O_31,N_19326,N_17082);
or UO_32 (O_32,N_15325,N_19778);
nor UO_33 (O_33,N_17541,N_18361);
nor UO_34 (O_34,N_16378,N_17064);
nor UO_35 (O_35,N_19361,N_18295);
nand UO_36 (O_36,N_17168,N_19151);
nand UO_37 (O_37,N_16080,N_15942);
nand UO_38 (O_38,N_16717,N_15827);
or UO_39 (O_39,N_17655,N_19192);
and UO_40 (O_40,N_15600,N_19345);
and UO_41 (O_41,N_15199,N_19862);
nand UO_42 (O_42,N_18040,N_18916);
nand UO_43 (O_43,N_17393,N_16493);
and UO_44 (O_44,N_17521,N_19113);
nand UO_45 (O_45,N_17138,N_19591);
or UO_46 (O_46,N_17727,N_19055);
nand UO_47 (O_47,N_18480,N_16906);
nand UO_48 (O_48,N_18027,N_17880);
and UO_49 (O_49,N_16055,N_16659);
and UO_50 (O_50,N_17098,N_19158);
and UO_51 (O_51,N_15062,N_18264);
nor UO_52 (O_52,N_19341,N_16592);
or UO_53 (O_53,N_17472,N_15808);
nand UO_54 (O_54,N_19756,N_19116);
or UO_55 (O_55,N_16469,N_18060);
or UO_56 (O_56,N_16459,N_19305);
nor UO_57 (O_57,N_16830,N_18929);
and UO_58 (O_58,N_17735,N_18848);
and UO_59 (O_59,N_16963,N_15139);
or UO_60 (O_60,N_15613,N_19638);
nor UO_61 (O_61,N_19431,N_18974);
and UO_62 (O_62,N_15332,N_17657);
or UO_63 (O_63,N_16739,N_16457);
nand UO_64 (O_64,N_18716,N_19425);
and UO_65 (O_65,N_16311,N_18789);
nand UO_66 (O_66,N_18165,N_19445);
nand UO_67 (O_67,N_17066,N_17603);
nor UO_68 (O_68,N_18181,N_18741);
or UO_69 (O_69,N_19359,N_19805);
nand UO_70 (O_70,N_18423,N_16173);
nor UO_71 (O_71,N_18428,N_15790);
xor UO_72 (O_72,N_17918,N_15418);
and UO_73 (O_73,N_19844,N_18055);
and UO_74 (O_74,N_17590,N_15391);
nor UO_75 (O_75,N_19319,N_19370);
and UO_76 (O_76,N_19247,N_16816);
and UO_77 (O_77,N_17654,N_16178);
xnor UO_78 (O_78,N_19426,N_18962);
and UO_79 (O_79,N_19164,N_17278);
nor UO_80 (O_80,N_16635,N_19487);
or UO_81 (O_81,N_17562,N_16207);
and UO_82 (O_82,N_16411,N_17758);
and UO_83 (O_83,N_16612,N_17357);
nor UO_84 (O_84,N_17706,N_17034);
nor UO_85 (O_85,N_17995,N_15310);
or UO_86 (O_86,N_16786,N_16965);
nand UO_87 (O_87,N_19238,N_18418);
nand UO_88 (O_88,N_19069,N_16001);
and UO_89 (O_89,N_15510,N_17999);
or UO_90 (O_90,N_19452,N_19236);
or UO_91 (O_91,N_17799,N_16541);
or UO_92 (O_92,N_19795,N_15078);
nand UO_93 (O_93,N_15338,N_16784);
nand UO_94 (O_94,N_16589,N_18651);
nor UO_95 (O_95,N_15145,N_19524);
nand UO_96 (O_96,N_17238,N_16980);
nand UO_97 (O_97,N_16390,N_19360);
xor UO_98 (O_98,N_15784,N_17186);
nor UO_99 (O_99,N_15799,N_16579);
nand UO_100 (O_100,N_19727,N_18864);
nor UO_101 (O_101,N_17163,N_16985);
and UO_102 (O_102,N_17612,N_15427);
nor UO_103 (O_103,N_18095,N_19941);
and UO_104 (O_104,N_15307,N_19136);
nor UO_105 (O_105,N_17302,N_15457);
or UO_106 (O_106,N_18129,N_16680);
or UO_107 (O_107,N_19447,N_19306);
and UO_108 (O_108,N_19088,N_17488);
nand UO_109 (O_109,N_15762,N_17376);
and UO_110 (O_110,N_16931,N_19507);
and UO_111 (O_111,N_19157,N_17973);
nand UO_112 (O_112,N_17964,N_18260);
nor UO_113 (O_113,N_18149,N_18851);
nor UO_114 (O_114,N_15598,N_17901);
and UO_115 (O_115,N_16891,N_15421);
nor UO_116 (O_116,N_15685,N_17150);
and UO_117 (O_117,N_18448,N_19397);
nand UO_118 (O_118,N_16409,N_16553);
and UO_119 (O_119,N_18364,N_15659);
or UO_120 (O_120,N_15910,N_18037);
nand UO_121 (O_121,N_18429,N_18865);
nand UO_122 (O_122,N_16687,N_15582);
nor UO_123 (O_123,N_16530,N_15702);
nand UO_124 (O_124,N_17526,N_17038);
or UO_125 (O_125,N_16498,N_17392);
and UO_126 (O_126,N_18955,N_16093);
or UO_127 (O_127,N_17041,N_19621);
nand UO_128 (O_128,N_17568,N_17923);
and UO_129 (O_129,N_19465,N_19186);
nor UO_130 (O_130,N_15365,N_18119);
and UO_131 (O_131,N_19526,N_17297);
or UO_132 (O_132,N_19123,N_16467);
nor UO_133 (O_133,N_18661,N_16196);
nand UO_134 (O_134,N_19746,N_16572);
nand UO_135 (O_135,N_16747,N_18273);
nand UO_136 (O_136,N_15937,N_18600);
and UO_137 (O_137,N_18893,N_18868);
nor UO_138 (O_138,N_18805,N_19409);
nor UO_139 (O_139,N_18297,N_18696);
or UO_140 (O_140,N_15324,N_19633);
nand UO_141 (O_141,N_18291,N_17725);
and UO_142 (O_142,N_19437,N_15846);
or UO_143 (O_143,N_15349,N_17881);
and UO_144 (O_144,N_15096,N_17193);
and UO_145 (O_145,N_17106,N_16430);
nand UO_146 (O_146,N_15905,N_19578);
or UO_147 (O_147,N_15259,N_18801);
nor UO_148 (O_148,N_18183,N_15483);
and UO_149 (O_149,N_15406,N_19841);
nor UO_150 (O_150,N_19467,N_17253);
nand UO_151 (O_151,N_19916,N_19943);
nand UO_152 (O_152,N_15233,N_15791);
nor UO_153 (O_153,N_19147,N_19567);
and UO_154 (O_154,N_18985,N_15943);
and UO_155 (O_155,N_19394,N_16061);
or UO_156 (O_156,N_18509,N_19721);
and UO_157 (O_157,N_15147,N_16298);
nand UO_158 (O_158,N_18502,N_18909);
and UO_159 (O_159,N_17810,N_15748);
nand UO_160 (O_160,N_15229,N_16256);
nand UO_161 (O_161,N_18201,N_15652);
nand UO_162 (O_162,N_16124,N_16586);
and UO_163 (O_163,N_17484,N_18826);
nor UO_164 (O_164,N_16797,N_15480);
xor UO_165 (O_165,N_18778,N_16342);
or UO_166 (O_166,N_18312,N_17862);
or UO_167 (O_167,N_17434,N_16277);
nor UO_168 (O_168,N_19608,N_17769);
nand UO_169 (O_169,N_15212,N_18798);
nor UO_170 (O_170,N_18918,N_17860);
xnor UO_171 (O_171,N_16836,N_17653);
or UO_172 (O_172,N_16594,N_18795);
and UO_173 (O_173,N_17592,N_17231);
or UO_174 (O_174,N_19269,N_19648);
nand UO_175 (O_175,N_18623,N_16242);
nand UO_176 (O_176,N_15741,N_19275);
nand UO_177 (O_177,N_19863,N_18535);
or UO_178 (O_178,N_17752,N_16289);
and UO_179 (O_179,N_19971,N_15719);
or UO_180 (O_180,N_18359,N_18103);
and UO_181 (O_181,N_19404,N_15572);
or UO_182 (O_182,N_18966,N_19838);
and UO_183 (O_183,N_15697,N_17931);
nand UO_184 (O_184,N_15639,N_17126);
and UO_185 (O_185,N_19111,N_16027);
nand UO_186 (O_186,N_15731,N_17446);
and UO_187 (O_187,N_18155,N_15594);
or UO_188 (O_188,N_16969,N_15793);
or UO_189 (O_189,N_18088,N_19294);
and UO_190 (O_190,N_17382,N_17520);
and UO_191 (O_191,N_19806,N_19324);
nand UO_192 (O_192,N_16622,N_16642);
nand UO_193 (O_193,N_16275,N_15909);
and UO_194 (O_194,N_16873,N_16559);
nand UO_195 (O_195,N_18999,N_16833);
nor UO_196 (O_196,N_16004,N_19557);
and UO_197 (O_197,N_15772,N_17258);
and UO_198 (O_198,N_19135,N_16326);
or UO_199 (O_199,N_15571,N_19995);
nor UO_200 (O_200,N_18907,N_19832);
or UO_201 (O_201,N_15006,N_16258);
and UO_202 (O_202,N_19541,N_15530);
nand UO_203 (O_203,N_15400,N_16267);
or UO_204 (O_204,N_15182,N_18350);
nor UO_205 (O_205,N_17989,N_19796);
and UO_206 (O_206,N_15975,N_16092);
nand UO_207 (O_207,N_17889,N_16658);
nor UO_208 (O_208,N_16600,N_17427);
nand UO_209 (O_209,N_16738,N_18882);
and UO_210 (O_210,N_16375,N_19745);
and UO_211 (O_211,N_15711,N_16395);
or UO_212 (O_212,N_17605,N_17268);
nand UO_213 (O_213,N_16231,N_19016);
nand UO_214 (O_214,N_16823,N_16380);
or UO_215 (O_215,N_18011,N_16304);
or UO_216 (O_216,N_15901,N_17295);
and UO_217 (O_217,N_18812,N_16981);
and UO_218 (O_218,N_18874,N_15911);
nor UO_219 (O_219,N_18348,N_18883);
and UO_220 (O_220,N_16736,N_15932);
and UO_221 (O_221,N_18041,N_16504);
nand UO_222 (O_222,N_16517,N_15879);
nand UO_223 (O_223,N_17948,N_15190);
nor UO_224 (O_224,N_19092,N_17777);
or UO_225 (O_225,N_15517,N_15626);
nor UO_226 (O_226,N_16677,N_16584);
nand UO_227 (O_227,N_16805,N_18067);
nand UO_228 (O_228,N_18970,N_19615);
or UO_229 (O_229,N_15557,N_16879);
or UO_230 (O_230,N_15895,N_15402);
and UO_231 (O_231,N_17188,N_19898);
nand UO_232 (O_232,N_17191,N_16616);
nand UO_233 (O_233,N_16502,N_19423);
or UO_234 (O_234,N_15274,N_16526);
or UO_235 (O_235,N_17543,N_18527);
and UO_236 (O_236,N_17452,N_16463);
nand UO_237 (O_237,N_17629,N_19099);
or UO_238 (O_238,N_18425,N_16669);
nor UO_239 (O_239,N_15467,N_16652);
nor UO_240 (O_240,N_16189,N_17548);
nor UO_241 (O_241,N_15912,N_17828);
nand UO_242 (O_242,N_17131,N_19885);
nand UO_243 (O_243,N_17534,N_19555);
nand UO_244 (O_244,N_18272,N_19701);
or UO_245 (O_245,N_16799,N_16132);
nor UO_246 (O_246,N_15746,N_19379);
or UO_247 (O_247,N_18357,N_16832);
nor UO_248 (O_248,N_15247,N_16661);
nor UO_249 (O_249,N_17703,N_16031);
nand UO_250 (O_250,N_17116,N_19436);
or UO_251 (O_251,N_17609,N_19282);
and UO_252 (O_252,N_16351,N_15605);
and UO_253 (O_253,N_17213,N_15488);
and UO_254 (O_254,N_19666,N_17378);
or UO_255 (O_255,N_15969,N_19751);
and UO_256 (O_256,N_17481,N_15944);
or UO_257 (O_257,N_17697,N_16251);
and UO_258 (O_258,N_19441,N_16676);
nor UO_259 (O_259,N_15713,N_15665);
and UO_260 (O_260,N_17121,N_16970);
or UO_261 (O_261,N_17440,N_19308);
nor UO_262 (O_262,N_19708,N_19657);
and UO_263 (O_263,N_16088,N_18518);
nor UO_264 (O_264,N_15952,N_18306);
xor UO_265 (O_265,N_17432,N_15110);
or UO_266 (O_266,N_17466,N_18915);
or UO_267 (O_267,N_17028,N_19312);
nand UO_268 (O_268,N_17770,N_19910);
xnor UO_269 (O_269,N_16455,N_15164);
nor UO_270 (O_270,N_16942,N_17486);
nand UO_271 (O_271,N_19685,N_15232);
or UO_272 (O_272,N_18588,N_17111);
or UO_273 (O_273,N_18235,N_15503);
nor UO_274 (O_274,N_16780,N_16647);
and UO_275 (O_275,N_15106,N_19558);
nor UO_276 (O_276,N_18757,N_17934);
nor UO_277 (O_277,N_15832,N_18845);
nand UO_278 (O_278,N_19152,N_15282);
nand UO_279 (O_279,N_18758,N_18712);
nand UO_280 (O_280,N_17153,N_16141);
or UO_281 (O_281,N_18597,N_19758);
nor UO_282 (O_282,N_18808,N_18369);
nand UO_283 (O_283,N_17981,N_17281);
and UO_284 (O_284,N_18629,N_19223);
nor UO_285 (O_285,N_16102,N_17864);
nor UO_286 (O_286,N_16255,N_17456);
or UO_287 (O_287,N_15997,N_19737);
nand UO_288 (O_288,N_18049,N_18979);
nand UO_289 (O_289,N_15250,N_16608);
and UO_290 (O_290,N_15159,N_19733);
nand UO_291 (O_291,N_19768,N_18025);
nand UO_292 (O_292,N_19378,N_16766);
and UO_293 (O_293,N_17001,N_15957);
and UO_294 (O_294,N_15722,N_18069);
or UO_295 (O_295,N_19040,N_17873);
and UO_296 (O_296,N_15558,N_16048);
nand UO_297 (O_297,N_18931,N_19546);
nor UO_298 (O_298,N_18515,N_19707);
or UO_299 (O_299,N_17699,N_16744);
or UO_300 (O_300,N_18786,N_16439);
and UO_301 (O_301,N_15223,N_17046);
nor UO_302 (O_302,N_16807,N_17899);
nand UO_303 (O_303,N_18086,N_16683);
nand UO_304 (O_304,N_16388,N_17927);
nand UO_305 (O_305,N_17817,N_16904);
and UO_306 (O_306,N_16427,N_17941);
nand UO_307 (O_307,N_16713,N_17365);
nor UO_308 (O_308,N_17876,N_16456);
nand UO_309 (O_309,N_18329,N_17475);
nor UO_310 (O_310,N_18380,N_17350);
nor UO_311 (O_311,N_17444,N_19814);
nor UO_312 (O_312,N_17494,N_19024);
nor UO_313 (O_313,N_16915,N_16544);
nor UO_314 (O_314,N_19229,N_19492);
or UO_315 (O_315,N_16224,N_17318);
and UO_316 (O_316,N_16522,N_15825);
nand UO_317 (O_317,N_15220,N_19387);
and UO_318 (O_318,N_17803,N_19280);
and UO_319 (O_319,N_15214,N_15743);
and UO_320 (O_320,N_18140,N_19328);
and UO_321 (O_321,N_18124,N_18332);
and UO_322 (O_322,N_15656,N_16776);
nor UO_323 (O_323,N_15297,N_17317);
nand UO_324 (O_324,N_16695,N_15404);
or UO_325 (O_325,N_17401,N_15148);
nor UO_326 (O_326,N_15570,N_19077);
and UO_327 (O_327,N_17537,N_15576);
and UO_328 (O_328,N_18701,N_18494);
and UO_329 (O_329,N_19692,N_18136);
nand UO_330 (O_330,N_18114,N_16999);
or UO_331 (O_331,N_17819,N_19327);
nand UO_332 (O_332,N_18836,N_16337);
nand UO_333 (O_333,N_15411,N_19653);
and UO_334 (O_334,N_19984,N_17890);
and UO_335 (O_335,N_17584,N_15999);
nor UO_336 (O_336,N_19278,N_19766);
or UO_337 (O_337,N_17276,N_18283);
or UO_338 (O_338,N_16049,N_17099);
nor UO_339 (O_339,N_19046,N_18605);
nor UO_340 (O_340,N_18464,N_17264);
nand UO_341 (O_341,N_17691,N_16007);
or UO_342 (O_342,N_18679,N_18520);
nor UO_343 (O_343,N_16334,N_19289);
and UO_344 (O_344,N_17512,N_17969);
or UO_345 (O_345,N_16485,N_18206);
or UO_346 (O_346,N_18310,N_16905);
or UO_347 (O_347,N_19942,N_17485);
or UO_348 (O_348,N_15841,N_15122);
xor UO_349 (O_349,N_17137,N_15837);
nor UO_350 (O_350,N_19400,N_19073);
nand UO_351 (O_351,N_16546,N_15794);
and UO_352 (O_352,N_19550,N_17420);
nand UO_353 (O_353,N_18031,N_19401);
and UO_354 (O_354,N_19089,N_16606);
and UO_355 (O_355,N_16309,N_19994);
nand UO_356 (O_356,N_15188,N_15244);
nor UO_357 (O_357,N_17059,N_19866);
nand UO_358 (O_358,N_19070,N_17510);
nor UO_359 (O_359,N_18569,N_19717);
nor UO_360 (O_360,N_17966,N_15986);
or UO_361 (O_361,N_19230,N_17073);
nand UO_362 (O_362,N_19117,N_19127);
or UO_363 (O_363,N_19835,N_18723);
and UO_364 (O_364,N_15029,N_15820);
nor UO_365 (O_365,N_17967,N_16703);
or UO_366 (O_366,N_16169,N_19281);
nor UO_367 (O_367,N_19977,N_18993);
nand UO_368 (O_368,N_16281,N_19163);
nand UO_369 (O_369,N_15392,N_16129);
nand UO_370 (O_370,N_18514,N_18557);
and UO_371 (O_371,N_15484,N_16547);
or UO_372 (O_372,N_18245,N_17049);
nand UO_373 (O_373,N_19334,N_15017);
nor UO_374 (O_374,N_16926,N_19990);
or UO_375 (O_375,N_17690,N_18138);
and UO_376 (O_376,N_15305,N_15448);
or UO_377 (O_377,N_15777,N_19783);
and UO_378 (O_378,N_18596,N_19313);
nor UO_379 (O_379,N_16042,N_17391);
or UO_380 (O_380,N_19318,N_19697);
nand UO_381 (O_381,N_17070,N_16580);
and UO_382 (O_382,N_15668,N_19877);
and UO_383 (O_383,N_18160,N_18615);
nor UO_384 (O_384,N_18400,N_16480);
and UO_385 (O_385,N_16097,N_19859);
or UO_386 (O_386,N_16690,N_18715);
nor UO_387 (O_387,N_15230,N_17042);
and UO_388 (O_388,N_15556,N_15355);
or UO_389 (O_389,N_18392,N_18358);
or UO_390 (O_390,N_16220,N_17418);
or UO_391 (O_391,N_16699,N_15298);
nand UO_392 (O_392,N_17566,N_19932);
or UO_393 (O_393,N_19671,N_19159);
nor UO_394 (O_394,N_15924,N_15028);
or UO_395 (O_395,N_17728,N_15553);
nor UO_396 (O_396,N_19097,N_17623);
or UO_397 (O_397,N_18875,N_18328);
nor UO_398 (O_398,N_18134,N_18780);
or UO_399 (O_399,N_17771,N_15989);
xnor UO_400 (O_400,N_19054,N_16868);
or UO_401 (O_401,N_15261,N_18132);
and UO_402 (O_402,N_19890,N_19944);
or UO_403 (O_403,N_19191,N_19085);
nand UO_404 (O_404,N_16556,N_19606);
nor UO_405 (O_405,N_16855,N_18495);
or UO_406 (O_406,N_17004,N_18809);
or UO_407 (O_407,N_18531,N_15885);
and UO_408 (O_408,N_19966,N_15979);
and UO_409 (O_409,N_17416,N_18612);
and UO_410 (O_410,N_16361,N_16651);
and UO_411 (O_411,N_19307,N_15495);
nor UO_412 (O_412,N_15803,N_19687);
nor UO_413 (O_413,N_19056,N_19095);
nand UO_414 (O_414,N_17007,N_18579);
and UO_415 (O_415,N_17821,N_17256);
nand UO_416 (O_416,N_19891,N_19443);
nor UO_417 (O_417,N_17710,N_19794);
nor UO_418 (O_418,N_19938,N_16641);
or UO_419 (O_419,N_19224,N_19494);
nor UO_420 (O_420,N_16436,N_19393);
or UO_421 (O_421,N_17354,N_15785);
nor UO_422 (O_422,N_19004,N_18378);
nor UO_423 (O_423,N_15688,N_19875);
or UO_424 (O_424,N_16692,N_16279);
nor UO_425 (O_425,N_15730,N_17305);
and UO_426 (O_426,N_16373,N_18517);
nand UO_427 (O_427,N_18642,N_16585);
and UO_428 (O_428,N_19876,N_16733);
nor UO_429 (O_429,N_17800,N_18263);
nor UO_430 (O_430,N_18156,N_16866);
or UO_431 (O_431,N_19048,N_16561);
and UO_432 (O_432,N_19676,N_19624);
nand UO_433 (O_433,N_18036,N_18513);
and UO_434 (O_434,N_17749,N_18824);
and UO_435 (O_435,N_19052,N_19979);
nor UO_436 (O_436,N_15617,N_17335);
or UO_437 (O_437,N_16523,N_16748);
xor UO_438 (O_438,N_16240,N_16629);
nor UO_439 (O_439,N_18933,N_18912);
nand UO_440 (O_440,N_19248,N_18048);
nor UO_441 (O_441,N_19964,N_18353);
or UO_442 (O_442,N_15379,N_19051);
nand UO_443 (O_443,N_18923,N_19476);
xor UO_444 (O_444,N_19170,N_19471);
and UO_445 (O_445,N_18213,N_15544);
nand UO_446 (O_446,N_17707,N_16993);
and UO_447 (O_447,N_15269,N_16443);
nand UO_448 (O_448,N_19346,N_17892);
or UO_449 (O_449,N_19517,N_19842);
nor UO_450 (O_450,N_17573,N_16109);
or UO_451 (O_451,N_19865,N_19497);
nand UO_452 (O_452,N_16858,N_19510);
nand UO_453 (O_453,N_17117,N_16893);
nand UO_454 (O_454,N_17569,N_15692);
and UO_455 (O_455,N_16028,N_18954);
or UO_456 (O_456,N_15460,N_18895);
or UO_457 (O_457,N_16192,N_16844);
nand UO_458 (O_458,N_16136,N_19506);
nor UO_459 (O_459,N_17961,N_17339);
nor UO_460 (O_460,N_17787,N_17398);
xnor UO_461 (O_461,N_16884,N_17785);
and UO_462 (O_462,N_16849,N_18507);
and UO_463 (O_463,N_19682,N_18549);
and UO_464 (O_464,N_15340,N_16764);
or UO_465 (O_465,N_17262,N_16322);
or UO_466 (O_466,N_15360,N_18718);
and UO_467 (O_467,N_17904,N_17721);
or UO_468 (O_468,N_18068,N_16214);
nand UO_469 (O_469,N_18344,N_19171);
and UO_470 (O_470,N_15792,N_16671);
xor UO_471 (O_471,N_16678,N_16698);
or UO_472 (O_472,N_19086,N_17000);
and UO_473 (O_473,N_15388,N_17146);
nor UO_474 (O_474,N_16313,N_15088);
nand UO_475 (O_475,N_19119,N_18382);
nand UO_476 (O_476,N_16073,N_17499);
or UO_477 (O_477,N_15610,N_19669);
and UO_478 (O_478,N_18568,N_19002);
and UO_479 (O_479,N_19679,N_18232);
and UO_480 (O_480,N_17811,N_15728);
and UO_481 (O_481,N_15318,N_16822);
and UO_482 (O_482,N_19927,N_19991);
or UO_483 (O_483,N_18243,N_18111);
nand UO_484 (O_484,N_17489,N_19490);
or UO_485 (O_485,N_19972,N_18373);
and UO_486 (O_486,N_18877,N_18253);
and UO_487 (O_487,N_15002,N_18844);
or UO_488 (O_488,N_15704,N_19839);
and UO_489 (O_489,N_16348,N_18855);
nor UO_490 (O_490,N_19083,N_15959);
or UO_491 (O_491,N_16759,N_16315);
and UO_492 (O_492,N_17080,N_15373);
and UO_493 (O_493,N_19775,N_18242);
nor UO_494 (O_494,N_19543,N_18115);
nand UO_495 (O_495,N_17282,N_15289);
or UO_496 (O_496,N_16106,N_16529);
or UO_497 (O_497,N_18409,N_17985);
and UO_498 (O_498,N_17279,N_18950);
nand UO_499 (O_499,N_19285,N_15204);
and UO_500 (O_500,N_18788,N_18469);
and UO_501 (O_501,N_16892,N_16164);
and UO_502 (O_502,N_17958,N_17898);
nand UO_503 (O_503,N_16997,N_17836);
nand UO_504 (O_504,N_16755,N_15773);
nor UO_505 (O_505,N_18305,N_17567);
nand UO_506 (O_506,N_19478,N_19268);
nand UO_507 (O_507,N_16190,N_19535);
and UO_508 (O_508,N_18179,N_18389);
nor UO_509 (O_509,N_18178,N_18898);
nand UO_510 (O_510,N_18450,N_19712);
nor UO_511 (O_511,N_19415,N_17523);
nor UO_512 (O_512,N_18952,N_19218);
or UO_513 (O_513,N_17069,N_15775);
nand UO_514 (O_514,N_18412,N_17247);
or UO_515 (O_515,N_17913,N_15971);
nor UO_516 (O_516,N_17953,N_19103);
nand UO_517 (O_517,N_18587,N_16391);
nor UO_518 (O_518,N_19139,N_16146);
and UO_519 (O_519,N_16241,N_18308);
nor UO_520 (O_520,N_17737,N_15314);
nand UO_521 (O_521,N_18168,N_18074);
or UO_522 (O_522,N_16927,N_18639);
or UO_523 (O_523,N_16971,N_18860);
and UO_524 (O_524,N_17225,N_17255);
and UO_525 (O_525,N_18486,N_19603);
and UO_526 (O_526,N_15508,N_15689);
nor UO_527 (O_527,N_19466,N_18983);
nand UO_528 (O_528,N_19260,N_16673);
or UO_529 (O_529,N_17714,N_18583);
nor UO_530 (O_530,N_15137,N_18886);
nor UO_531 (O_531,N_19444,N_19006);
or UO_532 (O_532,N_18393,N_15285);
nand UO_533 (O_533,N_18247,N_18534);
and UO_534 (O_534,N_17181,N_16276);
nor UO_535 (O_535,N_16270,N_15851);
nor UO_536 (O_536,N_15919,N_17431);
and UO_537 (O_537,N_19154,N_15393);
or UO_538 (O_538,N_16047,N_15525);
nor UO_539 (O_539,N_17425,N_15641);
and UO_540 (O_540,N_19323,N_17893);
nand UO_541 (O_541,N_19680,N_16912);
or UO_542 (O_542,N_18098,N_15044);
and UO_543 (O_543,N_18816,N_15705);
nor UO_544 (O_544,N_17700,N_18654);
nand UO_545 (O_545,N_18496,N_16216);
or UO_546 (O_546,N_17878,N_19764);
nand UO_547 (O_547,N_17413,N_18659);
and UO_548 (O_548,N_16053,N_18058);
nor UO_549 (O_549,N_18698,N_15260);
or UO_550 (O_550,N_17935,N_18072);
nor UO_551 (O_551,N_17435,N_19442);
or UO_552 (O_552,N_15519,N_15754);
nor UO_553 (O_553,N_17422,N_17780);
and UO_554 (O_554,N_15160,N_15051);
nor UO_555 (O_555,N_16806,N_18508);
nor UO_556 (O_556,N_19731,N_17433);
nor UO_557 (O_557,N_19166,N_17296);
nand UO_558 (O_558,N_17358,N_17345);
nor UO_559 (O_559,N_19337,N_16247);
nor UO_560 (O_560,N_15643,N_15101);
and UO_561 (O_561,N_17369,N_17778);
or UO_562 (O_562,N_19675,N_16609);
nand UO_563 (O_563,N_16966,N_16705);
and UO_564 (O_564,N_18799,N_16729);
nor UO_565 (O_565,N_17912,N_18504);
and UO_566 (O_566,N_16846,N_17493);
nand UO_567 (O_567,N_17459,N_19508);
nand UO_568 (O_568,N_16860,N_16840);
and UO_569 (O_569,N_19782,N_19340);
and UO_570 (O_570,N_15678,N_18398);
or UO_571 (O_571,N_15071,N_17610);
nand UO_572 (O_572,N_18200,N_17009);
and UO_573 (O_573,N_18564,N_19216);
nand UO_574 (O_574,N_16598,N_15118);
nand UO_575 (O_575,N_18943,N_15804);
and UO_576 (O_576,N_15990,N_15577);
or UO_577 (O_577,N_17204,N_16153);
nor UO_578 (O_578,N_19840,N_18045);
and UO_579 (O_579,N_18207,N_15520);
or UO_580 (O_580,N_15601,N_19061);
or UO_581 (O_581,N_15625,N_17457);
and UO_582 (O_582,N_18237,N_16901);
nor UO_583 (O_583,N_16573,N_16885);
and UO_584 (O_584,N_17845,N_17909);
or UO_585 (O_585,N_16071,N_17443);
or UO_586 (O_586,N_18194,N_16437);
or UO_587 (O_587,N_18014,N_16948);
and UO_588 (O_588,N_17381,N_15302);
or UO_589 (O_589,N_15584,N_18511);
nand UO_590 (O_590,N_15432,N_18797);
or UO_591 (O_591,N_17788,N_17652);
or UO_592 (O_592,N_16872,N_15345);
nand UO_593 (O_593,N_18727,N_18051);
nor UO_594 (O_594,N_15255,N_15474);
nor UO_595 (O_595,N_17036,N_15413);
xor UO_596 (O_596,N_18989,N_15853);
and UO_597 (O_597,N_15817,N_19475);
nand UO_598 (O_598,N_19735,N_19960);
nor UO_599 (O_599,N_19980,N_18284);
or UO_600 (O_600,N_17096,N_17996);
or UO_601 (O_601,N_19986,N_18184);
nor UO_602 (O_602,N_15714,N_17002);
or UO_603 (O_603,N_15485,N_17060);
nand UO_604 (O_604,N_16672,N_16257);
or UO_605 (O_605,N_17776,N_18337);
nand UO_606 (O_606,N_19187,N_18445);
and UO_607 (O_607,N_16707,N_16896);
nand UO_608 (O_608,N_16096,N_16461);
or UO_609 (O_609,N_18946,N_17414);
and UO_610 (O_610,N_17875,N_15934);
and UO_611 (O_611,N_19582,N_17848);
or UO_612 (O_612,N_16656,N_17688);
nor UO_613 (O_613,N_19226,N_17692);
and UO_614 (O_614,N_15915,N_15862);
nor UO_615 (O_615,N_16613,N_17216);
nor UO_616 (O_616,N_19078,N_15858);
nand UO_617 (O_617,N_18558,N_19043);
or UO_618 (O_618,N_18627,N_19632);
or UO_619 (O_619,N_16590,N_18458);
and UO_620 (O_620,N_16588,N_15593);
nor UO_621 (O_621,N_18085,N_18333);
and UO_622 (O_622,N_15676,N_17091);
nor UO_623 (O_623,N_19532,N_17856);
or UO_624 (O_624,N_19909,N_17016);
nand UO_625 (O_625,N_16711,N_19204);
nor UO_626 (O_626,N_19903,N_18018);
and UO_627 (O_627,N_18763,N_15624);
nand UO_628 (O_628,N_19585,N_17460);
nor UO_629 (O_629,N_18546,N_15541);
nand UO_630 (O_630,N_19371,N_17833);
or UO_631 (O_631,N_15154,N_16472);
or UO_632 (O_632,N_18147,N_18575);
or UO_633 (O_633,N_15589,N_16955);
or UO_634 (O_634,N_18703,N_19419);
and UO_635 (O_635,N_18252,N_16972);
nand UO_636 (O_636,N_17614,N_15100);
or UO_637 (O_637,N_18087,N_16741);
nor UO_638 (O_638,N_16149,N_18803);
or UO_639 (O_639,N_16557,N_16008);
and UO_640 (O_640,N_16398,N_18096);
or UO_641 (O_641,N_15767,N_15980);
nand UO_642 (O_642,N_16655,N_15437);
or UO_643 (O_643,N_18035,N_19185);
or UO_644 (O_644,N_15779,N_15596);
nand UO_645 (O_645,N_18510,N_19065);
nand UO_646 (O_646,N_18743,N_15976);
nor UO_647 (O_647,N_16175,N_19008);
and UO_648 (O_648,N_18814,N_17370);
or UO_649 (O_649,N_16688,N_18318);
nor UO_650 (O_650,N_19589,N_15085);
and UO_651 (O_651,N_17341,N_15333);
nor UO_652 (O_652,N_18128,N_17019);
or UO_653 (O_653,N_16983,N_17634);
or UO_654 (O_654,N_16441,N_15708);
and UO_655 (O_655,N_18614,N_16160);
nor UO_656 (O_656,N_16693,N_15947);
nand UO_657 (O_657,N_18968,N_19970);
nand UO_658 (O_658,N_15751,N_17932);
or UO_659 (O_659,N_19973,N_16552);
nand UO_660 (O_660,N_17371,N_18482);
nor UO_661 (O_661,N_17061,N_15595);
and UO_662 (O_662,N_15192,N_17855);
or UO_663 (O_663,N_19072,N_15802);
or UO_664 (O_664,N_19786,N_17071);
and UO_665 (O_665,N_19828,N_15465);
nor UO_666 (O_666,N_17349,N_17552);
and UO_667 (O_667,N_16660,N_16800);
and UO_668 (O_668,N_15251,N_15732);
nor UO_669 (O_669,N_17822,N_15893);
and UO_670 (O_670,N_17338,N_15926);
xor UO_671 (O_671,N_15518,N_19978);
nor UO_672 (O_672,N_17685,N_19924);
nor UO_673 (O_673,N_19831,N_15037);
and UO_674 (O_674,N_16290,N_19562);
nand UO_675 (O_675,N_15735,N_15439);
or UO_676 (O_676,N_18116,N_15532);
and UO_677 (O_677,N_18641,N_15150);
and UO_678 (O_678,N_17717,N_16254);
or UO_679 (O_679,N_18062,N_17217);
nor UO_680 (O_680,N_15539,N_17503);
nor UO_681 (O_681,N_18073,N_18584);
and UO_682 (O_682,N_15579,N_18082);
nor UO_683 (O_683,N_17447,N_15225);
and UO_684 (O_684,N_19141,N_16791);
and UO_685 (O_685,N_18551,N_19933);
and UO_686 (O_686,N_17943,N_19427);
or UO_687 (O_687,N_17324,N_18221);
nand UO_688 (O_688,N_18754,N_15316);
nand UO_689 (O_689,N_17743,N_16497);
nor UO_690 (O_690,N_16486,N_17619);
nor UO_691 (O_691,N_18066,N_15581);
nor UO_692 (O_692,N_16507,N_16300);
and UO_693 (O_693,N_15671,N_16925);
and UO_694 (O_694,N_19087,N_16731);
nand UO_695 (O_695,N_18131,N_18747);
and UO_696 (O_696,N_16213,N_18374);
or UO_697 (O_697,N_16466,N_17669);
or UO_698 (O_698,N_19231,N_15502);
nor UO_699 (O_699,N_17259,N_15384);
nand UO_700 (O_700,N_17753,N_19022);
and UO_701 (O_701,N_15201,N_19596);
nand UO_702 (O_702,N_16853,N_17911);
or UO_703 (O_703,N_17597,N_18960);
or UO_704 (O_704,N_18061,N_16908);
and UO_705 (O_705,N_17340,N_19005);
and UO_706 (O_706,N_19757,N_19132);
and UO_707 (O_707,N_19283,N_18720);
nand UO_708 (O_708,N_17419,N_15627);
and UO_709 (O_709,N_16899,N_17496);
nand UO_710 (O_710,N_19502,N_15165);
and UO_711 (O_711,N_19489,N_19176);
nor UO_712 (O_712,N_15857,N_19373);
nor UO_713 (O_713,N_17716,N_18793);
nand UO_714 (O_714,N_15554,N_19531);
nand UO_715 (O_715,N_16521,N_15954);
and UO_716 (O_716,N_19014,N_15152);
or UO_717 (O_717,N_17482,N_18800);
nor UO_718 (O_718,N_17219,N_16434);
and UO_719 (O_719,N_19178,N_19009);
nor UO_720 (O_720,N_18143,N_18497);
nand UO_721 (O_721,N_17453,N_16023);
or UO_722 (O_722,N_18280,N_16288);
nand UO_723 (O_723,N_15838,N_18403);
or UO_724 (O_724,N_17198,N_15420);
nand UO_725 (O_725,N_18834,N_16468);
nor UO_726 (O_726,N_16179,N_19619);
or UO_727 (O_727,N_16119,N_18064);
nand UO_728 (O_728,N_19481,N_19713);
or UO_729 (O_729,N_15869,N_19321);
nand UO_730 (O_730,N_19018,N_18281);
nand UO_731 (O_731,N_15115,N_19613);
or UO_732 (O_732,N_17373,N_17172);
nand UO_733 (O_733,N_15072,N_19527);
nor UO_734 (O_734,N_17665,N_15962);
and UO_735 (O_735,N_19982,N_16938);
nand UO_736 (O_736,N_16702,N_15938);
nand UO_737 (O_737,N_16916,N_19650);
nand UO_738 (O_738,N_15009,N_15861);
nand UO_739 (O_739,N_16152,N_17514);
nor UO_740 (O_740,N_18439,N_17008);
and UO_741 (O_741,N_15907,N_16236);
nand UO_742 (O_742,N_15016,N_18488);
nor UO_743 (O_743,N_15864,N_16923);
nor UO_744 (O_744,N_17742,N_19239);
and UO_745 (O_745,N_17424,N_15354);
nand UO_746 (O_746,N_18541,N_17403);
and UO_747 (O_747,N_18560,N_17540);
or UO_748 (O_748,N_19076,N_18170);
and UO_749 (O_749,N_16566,N_18043);
and UO_750 (O_750,N_15965,N_17269);
nor UO_751 (O_751,N_18973,N_16015);
nor UO_752 (O_752,N_19568,N_18891);
and UO_753 (O_753,N_17467,N_15181);
or UO_754 (O_754,N_19417,N_18630);
nor UO_755 (O_755,N_16909,N_15351);
nand UO_756 (O_756,N_16226,N_17250);
or UO_757 (O_757,N_17846,N_16813);
nor UO_758 (O_758,N_19576,N_19407);
nand UO_759 (O_759,N_17115,N_19599);
nor UO_760 (O_760,N_18335,N_15326);
nand UO_761 (O_761,N_16076,N_17355);
and UO_762 (O_762,N_15414,N_17994);
or UO_763 (O_763,N_19872,N_15870);
and UO_764 (O_764,N_19469,N_18745);
nor UO_765 (O_765,N_15972,N_18498);
nand UO_766 (O_766,N_17910,N_17386);
nor UO_767 (O_767,N_16924,N_19064);
or UO_768 (O_768,N_15295,N_15487);
nand UO_769 (O_769,N_17739,N_17574);
nor UO_770 (O_770,N_15135,N_16798);
and UO_771 (O_771,N_17593,N_17468);
nand UO_772 (O_772,N_17903,N_15945);
or UO_773 (O_773,N_15621,N_18857);
or UO_774 (O_774,N_15996,N_16575);
nor UO_775 (O_775,N_16295,N_17965);
nor UO_776 (O_776,N_18724,N_19210);
nor UO_777 (O_777,N_19598,N_18601);
or UO_778 (O_778,N_18404,N_18638);
and UO_779 (O_779,N_19353,N_15366);
nand UO_780 (O_780,N_18216,N_19422);
and UO_781 (O_781,N_17043,N_15399);
nand UO_782 (O_782,N_15313,N_15831);
nand UO_783 (O_783,N_15918,N_18383);
nor UO_784 (O_784,N_16161,N_19227);
nor UO_785 (O_785,N_19219,N_17886);
nor UO_786 (O_786,N_17081,N_19213);
or UO_787 (O_787,N_17549,N_17135);
nand UO_788 (O_788,N_15908,N_16861);
nand UO_789 (O_789,N_15454,N_16903);
or UO_790 (O_790,N_18435,N_19572);
or UO_791 (O_791,N_18674,N_18092);
nand UO_792 (O_792,N_18484,N_18794);
and UO_793 (O_793,N_17119,N_19013);
nor UO_794 (O_794,N_18740,N_15867);
nor UO_795 (O_795,N_16754,N_19240);
nor UO_796 (O_796,N_19800,N_17321);
or UO_797 (O_797,N_15551,N_19259);
nor UO_798 (O_798,N_15334,N_19772);
nor UO_799 (O_799,N_15003,N_16354);
nor UO_800 (O_800,N_16475,N_17143);
and UO_801 (O_801,N_18819,N_16895);
nor UO_802 (O_802,N_19612,N_17963);
nand UO_803 (O_803,N_18381,N_15466);
nor UO_804 (O_804,N_16944,N_17740);
and UO_805 (O_805,N_16087,N_16177);
nor UO_806 (O_806,N_17438,N_16232);
nand UO_807 (O_807,N_18982,N_19739);
nor UO_808 (O_808,N_18776,N_17202);
nor UO_809 (O_809,N_19681,N_19906);
or UO_810 (O_810,N_18193,N_19067);
and UO_811 (O_811,N_15272,N_18762);
or UO_812 (O_812,N_16244,N_17167);
nor UO_813 (O_813,N_16305,N_18924);
xor UO_814 (O_814,N_18516,N_19519);
nor UO_815 (O_815,N_16543,N_18222);
nor UO_816 (O_816,N_19150,N_15184);
nor UO_817 (O_817,N_15645,N_16188);
nor UO_818 (O_818,N_18083,N_15967);
nor UO_819 (O_819,N_19754,N_15469);
nand UO_820 (O_820,N_18090,N_18710);
and UO_821 (O_821,N_19382,N_16492);
and UO_822 (O_822,N_16841,N_16332);
and UO_823 (O_823,N_16157,N_16370);
and UO_824 (O_824,N_19246,N_18406);
and UO_825 (O_825,N_19232,N_19664);
nor UO_826 (O_826,N_16835,N_15674);
or UO_827 (O_827,N_19753,N_16176);
or UO_828 (O_828,N_18603,N_19292);
nand UO_829 (O_829,N_15620,N_16122);
nand UO_830 (O_830,N_16429,N_17554);
or UO_831 (O_831,N_16062,N_16266);
and UO_832 (O_832,N_15215,N_16788);
nand UO_833 (O_833,N_17950,N_18325);
nand UO_834 (O_834,N_18817,N_16292);
and UO_835 (O_835,N_16959,N_17229);
and UO_836 (O_836,N_18863,N_18956);
nor UO_837 (O_837,N_16432,N_18198);
nor UO_838 (O_838,N_18965,N_18624);
and UO_839 (O_839,N_19822,N_17968);
nor UO_840 (O_840,N_15607,N_17397);
or UO_841 (O_841,N_17683,N_17763);
nand UO_842 (O_842,N_17228,N_17977);
or UO_843 (O_843,N_19974,N_17628);
or UO_844 (O_844,N_16939,N_15648);
and UO_845 (O_845,N_15647,N_16320);
nor UO_846 (O_846,N_15927,N_19661);
nand UO_847 (O_847,N_15331,N_16740);
or UO_848 (O_848,N_15057,N_16126);
nand UO_849 (O_849,N_18476,N_18057);
or UO_850 (O_850,N_19569,N_19347);
and UO_851 (O_851,N_17222,N_17576);
or UO_852 (O_852,N_15046,N_16470);
nor UO_853 (O_853,N_16793,N_16331);
and UO_854 (O_854,N_18595,N_16091);
nand UO_855 (O_855,N_16538,N_15068);
nand UO_856 (O_856,N_19655,N_17065);
and UO_857 (O_857,N_18581,N_15178);
or UO_858 (O_858,N_18697,N_16084);
and UO_859 (O_859,N_18012,N_18167);
nor UO_860 (O_860,N_15545,N_19029);
and UO_861 (O_861,N_17077,N_18914);
nand UO_862 (O_862,N_17027,N_19999);
nand UO_863 (O_863,N_18410,N_15111);
or UO_864 (O_864,N_17547,N_17300);
nor UO_865 (O_865,N_16263,N_16448);
or UO_866 (O_866,N_18939,N_18684);
nand UO_867 (O_867,N_18395,N_16719);
nor UO_868 (O_868,N_16995,N_17155);
nor UO_869 (O_869,N_18402,N_18386);
and UO_870 (O_870,N_18655,N_17232);
or UO_871 (O_871,N_15239,N_18530);
or UO_872 (O_872,N_19145,N_18662);
or UO_873 (O_873,N_19594,N_18538);
and UO_874 (O_874,N_15872,N_17023);
and UO_875 (O_875,N_19921,N_18019);
and UO_876 (O_876,N_15567,N_17328);
or UO_877 (O_877,N_15833,N_16262);
or UO_878 (O_878,N_17947,N_17218);
nand UO_879 (O_879,N_16581,N_16783);
nand UO_880 (O_880,N_16419,N_17273);
or UO_881 (O_881,N_18953,N_19434);
or UO_882 (O_882,N_16537,N_16082);
nor UO_883 (O_883,N_19330,N_17448);
nor UO_884 (O_884,N_19670,N_19377);
or UO_885 (O_885,N_19954,N_15758);
or UO_886 (O_886,N_18266,N_18236);
nor UO_887 (O_887,N_16291,N_19937);
nor UO_888 (O_888,N_17748,N_18554);
nor UO_889 (O_889,N_18262,N_19759);
or UO_890 (O_890,N_15372,N_17148);
nor UO_891 (O_891,N_16113,N_17718);
or UO_892 (O_892,N_16476,N_19406);
nand UO_893 (O_893,N_15309,N_18023);
nor UO_894 (O_894,N_16582,N_19477);
nand UO_895 (O_895,N_17601,N_18265);
and UO_896 (O_896,N_17670,N_17618);
and UO_897 (O_897,N_18522,N_18818);
nor UO_898 (O_898,N_18278,N_17157);
or UO_899 (O_899,N_18125,N_16914);
and UO_900 (O_900,N_18223,N_16542);
and UO_901 (O_901,N_15712,N_15022);
or UO_902 (O_902,N_15429,N_18053);
and UO_903 (O_903,N_18971,N_19586);
nand UO_904 (O_904,N_16540,N_17972);
nor UO_905 (O_905,N_16135,N_16587);
or UO_906 (O_906,N_15278,N_18106);
and UO_907 (O_907,N_19118,N_17755);
and UO_908 (O_908,N_15622,N_16945);
nor UO_909 (O_909,N_15049,N_15382);
and UO_910 (O_910,N_18146,N_15168);
nand UO_911 (O_911,N_17177,N_19936);
nand UO_912 (O_912,N_16907,N_19242);
and UO_913 (O_913,N_19639,N_18729);
or UO_914 (O_914,N_15119,N_18345);
and UO_915 (O_915,N_17394,N_18225);
nor UO_916 (O_916,N_16479,N_19925);
nor UO_917 (O_917,N_15425,N_17937);
nor UO_918 (O_918,N_17796,N_18561);
and UO_919 (O_919,N_15315,N_19381);
or UO_920 (O_920,N_16187,N_17417);
nand UO_921 (O_921,N_18153,N_16820);
nand UO_922 (O_922,N_19044,N_16079);
or UO_923 (O_923,N_18761,N_19514);
nand UO_924 (O_924,N_15983,N_17887);
nand UO_925 (O_925,N_19156,N_18781);
or UO_926 (O_926,N_16715,N_15155);
nand UO_927 (O_927,N_16371,N_16743);
nor UO_928 (O_928,N_15105,N_17587);
or UO_929 (O_929,N_19725,N_17471);
nand UO_930 (O_930,N_17643,N_19262);
nor UO_931 (O_931,N_17051,N_15442);
xor UO_932 (O_932,N_18030,N_17089);
nor UO_933 (O_933,N_17841,N_18622);
nor UO_934 (O_934,N_18719,N_17353);
nand UO_935 (O_935,N_18046,N_19380);
nor UO_936 (O_936,N_18327,N_18483);
nor UO_937 (O_937,N_15348,N_16842);
nand UO_938 (O_938,N_15117,N_18802);
and UO_939 (O_939,N_15968,N_18901);
and UO_940 (O_940,N_15174,N_19516);
nor UO_941 (O_941,N_15319,N_15863);
nand UO_942 (O_942,N_19276,N_18997);
nor UO_943 (O_943,N_18958,N_17134);
nor UO_944 (O_944,N_16593,N_17733);
nor UO_945 (O_945,N_19565,N_18753);
or UO_946 (O_946,N_15745,N_17491);
and UO_947 (O_947,N_19511,N_17530);
nand UO_948 (O_948,N_15279,N_19854);
or UO_949 (O_949,N_16534,N_17867);
nand UO_950 (O_950,N_19367,N_17189);
or UO_951 (O_951,N_18726,N_17630);
nor UO_952 (O_952,N_15524,N_17842);
nor UO_953 (O_953,N_16674,N_16296);
nand UO_954 (O_954,N_16838,N_18499);
and UO_955 (O_955,N_15196,N_15536);
xor UO_956 (O_956,N_18244,N_15555);
nand UO_957 (O_957,N_19030,N_18241);
nor UO_958 (O_958,N_15292,N_17854);
nor UO_959 (O_959,N_19011,N_16211);
nor UO_960 (O_960,N_19858,N_15195);
nor UO_961 (O_961,N_16610,N_17578);
nand UO_962 (O_962,N_19130,N_15194);
nor UO_963 (O_963,N_19935,N_16170);
or UO_964 (O_964,N_18363,N_15854);
or UO_965 (O_965,N_16385,N_15890);
and UO_966 (O_966,N_18573,N_15638);
or UO_967 (O_967,N_19365,N_18054);
nand UO_968 (O_968,N_16710,N_19904);
nor UO_969 (O_969,N_17102,N_17542);
nor UO_970 (O_970,N_18694,N_17781);
nor UO_971 (O_971,N_19211,N_15038);
and UO_972 (O_972,N_16935,N_19287);
nor UO_973 (O_973,N_18120,N_19221);
or UO_974 (O_974,N_17334,N_19174);
and UO_975 (O_975,N_15368,N_15061);
and UO_976 (O_976,N_15866,N_19690);
or UO_977 (O_977,N_18311,N_17532);
nand UO_978 (O_978,N_19723,N_17185);
or UO_979 (O_979,N_19143,N_15881);
nand UO_980 (O_980,N_16396,N_19522);
or UO_981 (O_981,N_19563,N_19233);
or UO_982 (O_982,N_19787,N_19432);
nand UO_983 (O_983,N_15953,N_16444);
and UO_984 (O_984,N_19368,N_15739);
nor UO_985 (O_985,N_15920,N_18309);
and UO_986 (O_986,N_18417,N_16115);
nand UO_987 (O_987,N_18220,N_16140);
and UO_988 (O_988,N_15830,N_16870);
nor UO_989 (O_989,N_16977,N_18420);
nand UO_990 (O_990,N_19556,N_17006);
nor UO_991 (O_991,N_19513,N_19709);
and UO_992 (O_992,N_17037,N_19564);
and UO_993 (O_993,N_19581,N_19495);
and UO_994 (O_994,N_17458,N_18003);
and UO_995 (O_995,N_16417,N_18556);
nor UO_996 (O_996,N_16013,N_16054);
and UO_997 (O_997,N_16689,N_19039);
nand UO_998 (O_998,N_16583,N_15288);
nand UO_999 (O_999,N_16036,N_19631);
nand UO_1000 (O_1000,N_17109,N_15163);
nand UO_1001 (O_1001,N_18267,N_19684);
and UO_1002 (O_1002,N_17936,N_18782);
and UO_1003 (O_1003,N_19561,N_17975);
nor UO_1004 (O_1004,N_15205,N_17242);
nand UO_1005 (O_1005,N_18394,N_18742);
or UO_1006 (O_1006,N_17760,N_15898);
nor UO_1007 (O_1007,N_15219,N_16804);
nor UO_1008 (O_1008,N_15347,N_18806);
nand UO_1009 (O_1009,N_17056,N_18407);
and UO_1010 (O_1010,N_16329,N_16996);
nand UO_1011 (O_1011,N_16982,N_17764);
or UO_1012 (O_1012,N_18842,N_15795);
and UO_1013 (O_1013,N_19208,N_15560);
or UO_1014 (O_1014,N_17621,N_15224);
and UO_1015 (O_1015,N_18969,N_19483);
or UO_1016 (O_1016,N_15814,N_19104);
nand UO_1017 (O_1017,N_15724,N_17745);
and UO_1018 (O_1018,N_17531,N_19920);
nor UO_1019 (O_1019,N_16025,N_17551);
or UO_1020 (O_1020,N_16338,N_17680);
and UO_1021 (O_1021,N_19433,N_19694);
nand UO_1022 (O_1022,N_15761,N_16828);
or UO_1023 (O_1023,N_19332,N_18552);
or UO_1024 (O_1024,N_19716,N_19620);
and UO_1025 (O_1025,N_17283,N_15960);
nand UO_1026 (O_1026,N_19983,N_19702);
and UO_1027 (O_1027,N_15357,N_18360);
nor UO_1028 (O_1028,N_18613,N_15112);
nor UO_1029 (O_1029,N_16449,N_19989);
or UO_1030 (O_1030,N_19500,N_19349);
nor UO_1031 (O_1031,N_19658,N_18565);
nor UO_1032 (O_1032,N_18843,N_17715);
nand UO_1033 (O_1033,N_17497,N_15501);
and UO_1034 (O_1034,N_17852,N_19012);
nor UO_1035 (O_1035,N_15422,N_19931);
nor UO_1036 (O_1036,N_17779,N_16075);
and UO_1037 (O_1037,N_15537,N_16215);
and UO_1038 (O_1038,N_16795,N_19461);
nor UO_1039 (O_1039,N_16052,N_15813);
nand UO_1040 (O_1040,N_17118,N_18104);
nand UO_1041 (O_1041,N_16219,N_17075);
xor UO_1042 (O_1042,N_18859,N_18533);
nor UO_1043 (O_1043,N_17426,N_18927);
nand UO_1044 (O_1044,N_16897,N_15902);
nand UO_1045 (O_1045,N_17127,N_18239);
nand UO_1046 (O_1046,N_15042,N_18229);
nor UO_1047 (O_1047,N_16663,N_17789);
or UO_1048 (O_1048,N_19303,N_15974);
or UO_1049 (O_1049,N_17123,N_17270);
and UO_1050 (O_1050,N_19900,N_17129);
nor UO_1051 (O_1051,N_15829,N_16720);
and UO_1052 (O_1052,N_19254,N_17599);
nor UO_1053 (O_1053,N_15878,N_18135);
nand UO_1054 (O_1054,N_15516,N_17738);
or UO_1055 (O_1055,N_17348,N_17477);
and UO_1056 (O_1056,N_17645,N_19245);
and UO_1057 (O_1057,N_18375,N_19034);
or UO_1058 (O_1058,N_19637,N_16278);
nand UO_1059 (O_1059,N_15426,N_19781);
nand UO_1060 (O_1060,N_18044,N_16026);
or UO_1061 (O_1061,N_15103,N_16051);
xor UO_1062 (O_1062,N_17107,N_17402);
nor UO_1063 (O_1063,N_18945,N_19474);
nor UO_1064 (O_1064,N_18598,N_16953);
nor UO_1065 (O_1065,N_18021,N_15521);
and UO_1066 (O_1066,N_16230,N_18777);
nand UO_1067 (O_1067,N_17439,N_18107);
or UO_1068 (O_1068,N_15415,N_18203);
xor UO_1069 (O_1069,N_16888,N_15547);
nor UO_1070 (O_1070,N_16625,N_16509);
nor UO_1071 (O_1071,N_16060,N_15120);
and UO_1072 (O_1072,N_16854,N_15008);
nand UO_1073 (O_1073,N_17145,N_17616);
or UO_1074 (O_1074,N_19214,N_17396);
and UO_1075 (O_1075,N_15151,N_16050);
or UO_1076 (O_1076,N_16330,N_17906);
nor UO_1077 (O_1077,N_15409,N_18405);
nor UO_1078 (O_1078,N_18065,N_18268);
nor UO_1079 (O_1079,N_16346,N_17529);
or UO_1080 (O_1080,N_18150,N_19291);
nor UO_1081 (O_1081,N_15873,N_19082);
nand UO_1082 (O_1082,N_15896,N_18994);
nand UO_1083 (O_1083,N_18084,N_18750);
nor UO_1084 (O_1084,N_16967,N_15686);
nor UO_1085 (O_1085,N_18577,N_17293);
nand UO_1086 (O_1086,N_16975,N_17175);
nor UO_1087 (O_1087,N_18004,N_15376);
or UO_1088 (O_1088,N_18526,N_17088);
and UO_1089 (O_1089,N_16002,N_18991);
and UO_1090 (O_1090,N_19705,N_16011);
or UO_1091 (O_1091,N_18441,N_18224);
nor UO_1092 (O_1092,N_19521,N_19266);
nand UO_1093 (O_1093,N_16628,N_18177);
nor UO_1094 (O_1094,N_19929,N_18653);
nand UO_1095 (O_1095,N_16364,N_17084);
or UO_1096 (O_1096,N_19886,N_18371);
or UO_1097 (O_1097,N_15236,N_16482);
nor UO_1098 (O_1098,N_15789,N_18537);
nor UO_1099 (O_1099,N_15591,N_19930);
or UO_1100 (O_1100,N_15369,N_17641);
nand UO_1101 (O_1101,N_17988,N_17806);
or UO_1102 (O_1102,N_19271,N_19129);
or UO_1103 (O_1103,N_19484,N_15173);
nor UO_1104 (O_1104,N_15303,N_18609);
nand UO_1105 (O_1105,N_16118,N_17765);
nand UO_1106 (O_1106,N_17589,N_19873);
nor UO_1107 (O_1107,N_15496,N_15102);
nand UO_1108 (O_1108,N_17583,N_17580);
or UO_1109 (O_1109,N_17430,N_17063);
nor UO_1110 (O_1110,N_16763,N_15056);
nor UO_1111 (O_1111,N_16000,N_16607);
nor UO_1112 (O_1112,N_18465,N_19908);
nand UO_1113 (O_1113,N_19953,N_17139);
nand UO_1114 (O_1114,N_16183,N_19647);
nor UO_1115 (O_1115,N_19602,N_18699);
and UO_1116 (O_1116,N_19992,N_15543);
or UO_1117 (O_1117,N_15082,N_15073);
nand UO_1118 (O_1118,N_17871,N_15491);
and UO_1119 (O_1119,N_19320,N_18478);
nor UO_1120 (O_1120,N_15852,N_17201);
and UO_1121 (O_1121,N_15015,N_18959);
or UO_1122 (O_1122,N_19315,N_16894);
and UO_1123 (O_1123,N_16405,N_18139);
and UO_1124 (O_1124,N_16412,N_17791);
and UO_1125 (O_1125,N_17518,N_15218);
and UO_1126 (O_1126,N_16640,N_16818);
nor UO_1127 (O_1127,N_16936,N_16171);
nor UO_1128 (O_1128,N_17389,N_19945);
and UO_1129 (O_1129,N_18941,N_19955);
or UO_1130 (O_1130,N_16886,N_19975);
and UO_1131 (O_1131,N_17775,N_16591);
nor UO_1132 (O_1132,N_17974,N_17220);
nor UO_1133 (O_1133,N_17850,N_18990);
nand UO_1134 (O_1134,N_18858,N_17195);
nor UO_1135 (O_1135,N_18454,N_15489);
and UO_1136 (O_1136,N_18547,N_16081);
and UO_1137 (O_1137,N_18489,N_16555);
and UO_1138 (O_1138,N_19212,N_17363);
nand UO_1139 (O_1139,N_18572,N_19042);
and UO_1140 (O_1140,N_15079,N_18543);
and UO_1141 (O_1141,N_19317,N_16269);
and UO_1142 (O_1142,N_17029,N_15398);
xnor UO_1143 (O_1143,N_15107,N_16774);
nor UO_1144 (O_1144,N_16937,N_16511);
and UO_1145 (O_1145,N_16536,N_15461);
and UO_1146 (O_1146,N_15097,N_18890);
nand UO_1147 (O_1147,N_18610,N_17068);
xor UO_1148 (O_1148,N_19454,N_19311);
nand UO_1149 (O_1149,N_17461,N_15588);
and UO_1150 (O_1150,N_17647,N_19691);
and UO_1151 (O_1151,N_15245,N_15655);
or UO_1152 (O_1152,N_19133,N_17375);
or UO_1153 (O_1153,N_15197,N_15162);
nor UO_1154 (O_1154,N_18320,N_16750);
or UO_1155 (O_1155,N_18042,N_16782);
or UO_1156 (O_1156,N_18118,N_15361);
nand UO_1157 (O_1157,N_19408,N_18322);
and UO_1158 (O_1158,N_15629,N_15311);
nand UO_1159 (O_1159,N_18706,N_17940);
and UO_1160 (O_1160,N_16991,N_15463);
nor UO_1161 (O_1161,N_17897,N_17604);
and UO_1162 (O_1162,N_16488,N_19142);
nand UO_1163 (O_1163,N_17544,N_15175);
and UO_1164 (O_1164,N_16238,N_17527);
or UO_1165 (O_1165,N_15252,N_17380);
nor UO_1166 (O_1166,N_16044,N_17839);
nor UO_1167 (O_1167,N_15301,N_15221);
nor UO_1168 (O_1168,N_16034,N_15531);
or UO_1169 (O_1169,N_17100,N_18677);
nor UO_1170 (O_1170,N_19610,N_16558);
nor UO_1171 (O_1171,N_19463,N_16623);
or UO_1172 (O_1172,N_15683,N_18424);
nor UO_1173 (O_1173,N_17325,N_15694);
nand UO_1174 (O_1174,N_18578,N_15913);
nand UO_1175 (O_1175,N_15198,N_15755);
or UO_1176 (O_1176,N_17464,N_19860);
or UO_1177 (O_1177,N_16549,N_19704);
nor UO_1178 (O_1178,N_15424,N_18434);
nand UO_1179 (O_1179,N_17658,N_16984);
nor UO_1180 (O_1180,N_15619,N_15013);
and UO_1181 (O_1181,N_15742,N_15492);
nand UO_1182 (O_1182,N_17344,N_18813);
nand UO_1183 (O_1183,N_17644,N_15287);
nor UO_1184 (O_1184,N_16340,N_18774);
nand UO_1185 (O_1185,N_17640,N_19288);
nand UO_1186 (O_1186,N_16154,N_16762);
nand UO_1187 (O_1187,N_16303,N_18619);
nand UO_1188 (O_1188,N_19388,N_19194);
and UO_1189 (O_1189,N_17272,N_16657);
and UO_1190 (O_1190,N_18089,N_15430);
and UO_1191 (O_1191,N_16245,N_19809);
nand UO_1192 (O_1192,N_17946,N_19060);
nand UO_1193 (O_1193,N_18354,N_16630);
nor UO_1194 (O_1194,N_17178,N_17992);
nor UO_1195 (O_1195,N_16142,N_17939);
nor UO_1196 (O_1196,N_16721,N_17200);
xor UO_1197 (O_1197,N_15440,N_16650);
or UO_1198 (O_1198,N_16195,N_19180);
nand UO_1199 (O_1199,N_18251,N_18372);
and UO_1200 (O_1200,N_18647,N_15805);
nor UO_1201 (O_1201,N_16527,N_17895);
nor UO_1202 (O_1202,N_18676,N_16706);
and UO_1203 (O_1203,N_17267,N_18833);
xnor UO_1204 (O_1204,N_19688,N_16775);
nor UO_1205 (O_1205,N_19348,N_16360);
xor UO_1206 (O_1206,N_19115,N_15126);
nand UO_1207 (O_1207,N_15925,N_17241);
nor UO_1208 (O_1208,N_17136,N_17708);
or UO_1209 (O_1209,N_19846,N_19830);
or UO_1210 (O_1210,N_15535,N_19241);
nand UO_1211 (O_1211,N_17786,N_18702);
nor UO_1212 (O_1212,N_16070,N_17400);
or UO_1213 (O_1213,N_17022,N_15928);
and UO_1214 (O_1214,N_19126,N_18664);
nor UO_1215 (O_1215,N_19902,N_18938);
nor UO_1216 (O_1216,N_16667,N_16550);
or UO_1217 (O_1217,N_16843,N_17945);
or UO_1218 (O_1218,N_15262,N_15651);
and UO_1219 (O_1219,N_19617,N_19148);
and UO_1220 (O_1220,N_15256,N_17347);
or UO_1221 (O_1221,N_16911,N_19389);
nor UO_1222 (O_1222,N_17271,N_17933);
and UO_1223 (O_1223,N_17501,N_15590);
nand UO_1224 (O_1224,N_19000,N_19878);
or UO_1225 (O_1225,N_15880,N_16335);
or UO_1226 (O_1226,N_18524,N_15606);
xor UO_1227 (O_1227,N_19549,N_18078);
nand UO_1228 (O_1228,N_15158,N_17659);
or UO_1229 (O_1229,N_16384,N_17450);
nor UO_1230 (O_1230,N_17311,N_16185);
nor UO_1231 (O_1231,N_16745,N_15946);
nor UO_1232 (O_1232,N_17579,N_15363);
nand UO_1233 (O_1233,N_18259,N_16282);
nand UO_1234 (O_1234,N_16859,N_15138);
nand UO_1235 (O_1235,N_18390,N_19821);
nor UO_1236 (O_1236,N_15133,N_15385);
nor UO_1237 (O_1237,N_15611,N_15657);
and UO_1238 (O_1238,N_17825,N_16108);
and UO_1239 (O_1239,N_17571,N_19058);
and UO_1240 (O_1240,N_16454,N_17681);
nor UO_1241 (O_1241,N_16570,N_19273);
nand UO_1242 (O_1242,N_15023,N_16085);
and UO_1243 (O_1243,N_16345,N_17675);
nor UO_1244 (O_1244,N_19996,N_19744);
xnor UO_1245 (O_1245,N_16321,N_17802);
nor UO_1246 (O_1246,N_17761,N_17563);
nor UO_1247 (O_1247,N_18453,N_17783);
nor UO_1248 (O_1248,N_16229,N_17248);
nand UO_1249 (O_1249,N_18519,N_15308);
and UO_1250 (O_1250,N_17199,N_16974);
nand UO_1251 (O_1251,N_17978,N_17823);
nand UO_1252 (O_1252,N_18755,N_16626);
or UO_1253 (O_1253,N_19265,N_19217);
nand UO_1254 (O_1254,N_19468,N_15527);
nor UO_1255 (O_1255,N_15083,N_19396);
or UO_1256 (O_1256,N_18349,N_18657);
and UO_1257 (O_1257,N_18334,N_17528);
and UO_1258 (O_1258,N_17684,N_19094);
or UO_1259 (O_1259,N_16199,N_15211);
nand UO_1260 (O_1260,N_19528,N_15660);
nand UO_1261 (O_1261,N_18852,N_17774);
or UO_1262 (O_1262,N_17539,N_15780);
nand UO_1263 (O_1263,N_15322,N_18151);
nand UO_1264 (O_1264,N_18276,N_15136);
or UO_1265 (O_1265,N_17596,N_19161);
or UO_1266 (O_1266,N_16250,N_15296);
or UO_1267 (O_1267,N_18287,N_19643);
or UO_1268 (O_1268,N_15018,N_19673);
or UO_1269 (O_1269,N_18866,N_17180);
nor UO_1270 (O_1270,N_16066,N_17724);
or UO_1271 (O_1271,N_18302,N_15931);
nand UO_1272 (O_1272,N_15010,N_15749);
or UO_1273 (O_1273,N_19997,N_18274);
nor UO_1274 (O_1274,N_15364,N_18505);
and UO_1275 (O_1275,N_17352,N_17902);
and UO_1276 (O_1276,N_16212,N_19825);
nand UO_1277 (O_1277,N_19355,N_17309);
nor UO_1278 (O_1278,N_15226,N_19405);
nand UO_1279 (O_1279,N_17798,N_15876);
nor UO_1280 (O_1280,N_15707,N_18112);
and UO_1281 (O_1281,N_15993,N_19662);
nor UO_1282 (O_1282,N_19001,N_17678);
nor UO_1283 (O_1283,N_18940,N_18964);
nand UO_1284 (O_1284,N_15756,N_16318);
nand UO_1285 (O_1285,N_15757,N_18695);
nand UO_1286 (O_1286,N_16058,N_18673);
xnor UO_1287 (O_1287,N_15695,N_19272);
nor UO_1288 (O_1288,N_16852,N_19493);
or UO_1289 (O_1289,N_18002,N_18512);
nor UO_1290 (O_1290,N_19743,N_16059);
and UO_1291 (O_1291,N_16976,N_17951);
nor UO_1292 (O_1292,N_18296,N_17104);
and UO_1293 (O_1293,N_17679,N_17288);
and UO_1294 (O_1294,N_15810,N_19137);
nand UO_1295 (O_1295,N_16812,N_15916);
and UO_1296 (O_1296,N_17290,N_15121);
and UO_1297 (O_1297,N_16821,N_17021);
nor UO_1298 (O_1298,N_18385,N_15575);
nor UO_1299 (O_1299,N_17600,N_18637);
or UO_1300 (O_1300,N_17627,N_16451);
and UO_1301 (O_1301,N_17917,N_18539);
nor UO_1302 (O_1302,N_19125,N_16851);
nand UO_1303 (O_1303,N_18231,N_19491);
or UO_1304 (O_1304,N_15249,N_18342);
nor UO_1305 (O_1305,N_17428,N_19850);
or UO_1306 (O_1306,N_15434,N_17035);
nor UO_1307 (O_1307,N_18182,N_17207);
nand UO_1308 (O_1308,N_16605,N_17695);
or UO_1309 (O_1309,N_18986,N_17025);
and UO_1310 (O_1310,N_15090,N_16929);
nand UO_1311 (O_1311,N_15966,N_16103);
nand UO_1312 (O_1312,N_15995,N_18604);
nor UO_1313 (O_1313,N_15618,N_15464);
nand UO_1314 (O_1314,N_16771,N_15877);
nor UO_1315 (O_1315,N_17956,N_16235);
and UO_1316 (O_1316,N_15736,N_17149);
or UO_1317 (O_1317,N_19091,N_17712);
or UO_1318 (O_1318,N_18079,N_17190);
xnor UO_1319 (O_1319,N_16520,N_17495);
nor UO_1320 (O_1320,N_16484,N_17709);
and UO_1321 (O_1321,N_15950,N_17896);
or UO_1322 (O_1322,N_19263,N_15935);
nand UO_1323 (O_1323,N_15428,N_18876);
nor UO_1324 (O_1324,N_15089,N_15958);
or UO_1325 (O_1325,N_18075,N_19429);
and UO_1326 (O_1326,N_16601,N_15330);
nand UO_1327 (O_1327,N_15189,N_18947);
or UO_1328 (O_1328,N_19856,N_15471);
nor UO_1329 (O_1329,N_16827,N_15077);
nor UO_1330 (O_1330,N_19375,N_16078);
and UO_1331 (O_1331,N_15098,N_15499);
or UO_1332 (O_1332,N_18784,N_18158);
nor UO_1333 (O_1333,N_16045,N_15923);
nand UO_1334 (O_1334,N_16131,N_17885);
or UO_1335 (O_1335,N_19819,N_15691);
nor UO_1336 (O_1336,N_18102,N_15865);
or UO_1337 (O_1337,N_19106,N_18765);
nor UO_1338 (O_1338,N_18026,N_16727);
nor UO_1339 (O_1339,N_16943,N_19096);
and UO_1340 (O_1340,N_19488,N_19153);
and UO_1341 (O_1341,N_19719,N_16510);
and UO_1342 (O_1342,N_17615,N_15533);
nor UO_1343 (O_1343,N_16902,N_19225);
and UO_1344 (O_1344,N_15886,N_17804);
or UO_1345 (O_1345,N_18157,N_17991);
or UO_1346 (O_1346,N_19110,N_17280);
nor UO_1347 (O_1347,N_16890,N_16453);
and UO_1348 (O_1348,N_15149,N_17611);
or UO_1349 (O_1349,N_18721,N_17164);
and UO_1350 (O_1350,N_15490,N_17602);
and UO_1351 (O_1351,N_17490,N_18148);
nor UO_1352 (O_1352,N_15011,N_18491);
or UO_1353 (O_1353,N_17166,N_18101);
nor UO_1354 (O_1354,N_19722,N_16643);
nor UO_1355 (O_1355,N_18911,N_15240);
and UO_1356 (O_1356,N_18341,N_16777);
nand UO_1357 (O_1357,N_19776,N_18109);
nor UO_1358 (O_1358,N_15701,N_19738);
nor UO_1359 (O_1359,N_17319,N_15276);
and UO_1360 (O_1360,N_16714,N_15721);
or UO_1361 (O_1361,N_16578,N_19587);
or UO_1362 (O_1362,N_18432,N_19742);
or UO_1363 (O_1363,N_16301,N_19031);
nor UO_1364 (O_1364,N_16392,N_17984);
and UO_1365 (O_1365,N_15371,N_18871);
nand UO_1366 (O_1366,N_16620,N_15988);
nor UO_1367 (O_1367,N_16228,N_18033);
or UO_1368 (O_1368,N_17313,N_16317);
or UO_1369 (O_1369,N_15844,N_15889);
nor UO_1370 (O_1370,N_15468,N_19577);
nand UO_1371 (O_1371,N_18288,N_19179);
nor UO_1372 (O_1372,N_18304,N_19122);
nand UO_1373 (O_1373,N_19845,N_17374);
or UO_1374 (O_1374,N_16148,N_18477);
and UO_1375 (O_1375,N_17767,N_16406);
nor UO_1376 (O_1376,N_15628,N_19811);
nand UO_1377 (O_1377,N_16681,N_15690);
nor UO_1378 (O_1378,N_17863,N_18691);
nand UO_1379 (O_1379,N_17884,N_15446);
nand UO_1380 (O_1380,N_19537,N_16014);
and UO_1381 (O_1381,N_17916,N_16206);
nand UO_1382 (O_1382,N_15700,N_16947);
nor UO_1383 (O_1383,N_17631,N_16770);
or UO_1384 (O_1384,N_16865,N_18028);
or UO_1385 (O_1385,N_18900,N_17617);
nor UO_1386 (O_1386,N_17197,N_19907);
or UO_1387 (O_1387,N_16941,N_16365);
or UO_1388 (O_1388,N_18426,N_18559);
nand UO_1389 (O_1389,N_18854,N_19264);
nor UO_1390 (O_1390,N_15027,N_18746);
and UO_1391 (O_1391,N_16952,N_15328);
nand UO_1392 (O_1392,N_18725,N_15124);
nor UO_1393 (O_1393,N_19503,N_19080);
and UO_1394 (O_1394,N_15550,N_19108);
nand UO_1395 (O_1395,N_19826,N_19182);
and UO_1396 (O_1396,N_16127,N_19748);
xor UO_1397 (O_1397,N_17686,N_15747);
nand UO_1398 (O_1398,N_16531,N_18669);
nor UO_1399 (O_1399,N_15566,N_15542);
or UO_1400 (O_1400,N_16875,N_18034);
nor UO_1401 (O_1401,N_15515,N_17929);
nor UO_1402 (O_1402,N_17263,N_17650);
nand UO_1403 (O_1403,N_17090,N_17831);
or UO_1404 (O_1404,N_15951,N_17663);
or UO_1405 (O_1405,N_19504,N_17237);
or UO_1406 (O_1406,N_16128,N_19659);
and UO_1407 (O_1407,N_19696,N_16874);
nand UO_1408 (O_1408,N_15370,N_15897);
or UO_1409 (O_1409,N_17747,N_18847);
nand UO_1410 (O_1410,N_15494,N_17266);
or UO_1411 (O_1411,N_18708,N_18161);
nand UO_1412 (O_1412,N_19861,N_17030);
nand UO_1413 (O_1413,N_15447,N_16856);
nor UO_1414 (O_1414,N_19874,N_17792);
or UO_1415 (O_1415,N_15380,N_18925);
or UO_1416 (O_1416,N_16299,N_16261);
nor UO_1417 (O_1417,N_19523,N_19277);
and UO_1418 (O_1418,N_19530,N_16069);
xor UO_1419 (O_1419,N_19812,N_18123);
nor UO_1420 (O_1420,N_16210,N_15505);
nand UO_1421 (O_1421,N_17003,N_16615);
nand UO_1422 (O_1422,N_16381,N_19399);
nor UO_1423 (O_1423,N_18831,N_19790);
and UO_1424 (O_1424,N_16359,N_18832);
nand UO_1425 (O_1425,N_17455,N_15054);
or UO_1426 (O_1426,N_15892,N_17245);
and UO_1427 (O_1427,N_15836,N_15180);
nand UO_1428 (O_1428,N_15698,N_15177);
or UO_1429 (O_1429,N_15764,N_17812);
and UO_1430 (O_1430,N_19062,N_15578);
nand UO_1431 (O_1431,N_15081,N_18121);
or UO_1432 (O_1432,N_18667,N_15763);
and UO_1433 (O_1433,N_19720,N_16325);
nand UO_1434 (O_1434,N_19482,N_18362);
nor UO_1435 (O_1435,N_19988,N_18644);
and UO_1436 (O_1436,N_18714,N_17986);
nor UO_1437 (O_1437,N_19749,N_18256);
or UO_1438 (O_1438,N_15036,N_17942);
or UO_1439 (O_1439,N_17094,N_16111);
and UO_1440 (O_1440,N_15770,N_18100);
or UO_1441 (O_1441,N_15933,N_16144);
nor UO_1442 (O_1442,N_15356,N_15973);
and UO_1443 (O_1443,N_17504,N_18289);
nand UO_1444 (O_1444,N_19168,N_16116);
or UO_1445 (O_1445,N_17469,N_17331);
nand UO_1446 (O_1446,N_15273,N_18175);
and UO_1447 (O_1447,N_19881,N_19762);
nor UO_1448 (O_1448,N_16043,N_15573);
nand UO_1449 (O_1449,N_17169,N_19799);
nand UO_1450 (O_1450,N_16064,N_19993);
nand UO_1451 (O_1451,N_19580,N_15585);
and UO_1452 (O_1452,N_19848,N_19374);
or UO_1453 (O_1453,N_15458,N_15074);
and UO_1454 (O_1454,N_15504,N_17323);
and UO_1455 (O_1455,N_18271,N_16500);
nor UO_1456 (O_1456,N_15840,N_17437);
or UO_1457 (O_1457,N_15268,N_15681);
nand UO_1458 (O_1458,N_15649,N_15684);
and UO_1459 (O_1459,N_17868,N_16041);
nor UO_1460 (O_1460,N_17083,N_15336);
or UO_1461 (O_1461,N_19533,N_15842);
nand UO_1462 (O_1462,N_19948,N_16209);
nor UO_1463 (O_1463,N_19544,N_15848);
and UO_1464 (O_1464,N_17257,N_16143);
nand UO_1465 (O_1465,N_17795,N_19660);
nor UO_1466 (O_1466,N_17128,N_17516);
nor UO_1467 (O_1467,N_17642,N_18897);
nor UO_1468 (O_1468,N_19071,N_18270);
or UO_1469 (O_1469,N_16100,N_15141);
nor UO_1470 (O_1470,N_18617,N_19625);
and UO_1471 (O_1471,N_19829,N_16599);
and UO_1472 (O_1472,N_17938,N_15765);
nand UO_1473 (O_1473,N_17782,N_19571);
and UO_1474 (O_1474,N_16701,N_18314);
or UO_1475 (O_1475,N_17234,N_19736);
nor UO_1476 (O_1476,N_19411,N_17572);
nor UO_1477 (O_1477,N_18738,N_19257);
nand UO_1478 (O_1478,N_17722,N_18347);
nor UO_1479 (O_1479,N_19732,N_15506);
nor UO_1480 (O_1480,N_16336,N_15682);
or UO_1481 (O_1481,N_15007,N_15725);
and UO_1482 (O_1482,N_16627,N_15191);
nor UO_1483 (O_1483,N_17814,N_15548);
and UO_1484 (O_1484,N_17441,N_18422);
or UO_1485 (O_1485,N_19279,N_17078);
nor UO_1486 (O_1486,N_15703,N_18173);
or UO_1487 (O_1487,N_18978,N_19107);
nand UO_1488 (O_1488,N_19033,N_18493);
and UO_1489 (O_1489,N_15816,N_18254);
nand UO_1490 (O_1490,N_16826,N_19627);
nand UO_1491 (O_1491,N_15940,N_19770);
nand UO_1492 (O_1492,N_16362,N_19817);
nor UO_1493 (O_1493,N_18077,N_16961);
or UO_1494 (O_1494,N_15045,N_19366);
and UO_1495 (O_1495,N_18462,N_16353);
nor UO_1496 (O_1496,N_18709,N_18397);
nor UO_1497 (O_1497,N_19777,N_15445);
nand UO_1498 (O_1498,N_17877,N_18269);
nand UO_1499 (O_1499,N_19149,N_16919);
and UO_1500 (O_1500,N_19121,N_19959);
nor UO_1501 (O_1501,N_17463,N_19912);
nand UO_1502 (O_1502,N_16205,N_15766);
nand UO_1503 (O_1503,N_18440,N_15835);
nor UO_1504 (O_1504,N_15482,N_18456);
nand UO_1505 (O_1505,N_15709,N_19237);
nand UO_1506 (O_1506,N_17672,N_16067);
nor UO_1507 (O_1507,N_15994,N_17498);
nor UO_1508 (O_1508,N_18899,N_18117);
and UO_1509 (O_1509,N_15956,N_16501);
nor UO_1510 (O_1510,N_16645,N_19922);
nor UO_1511 (O_1511,N_16708,N_17508);
and UO_1512 (O_1512,N_15964,N_17492);
or UO_1513 (O_1513,N_19820,N_19798);
nor UO_1514 (O_1514,N_16077,N_18772);
and UO_1515 (O_1515,N_19823,N_15227);
nand UO_1516 (O_1516,N_18704,N_19300);
or UO_1517 (O_1517,N_16560,N_16287);
nand UO_1518 (O_1518,N_17320,N_18340);
nor UO_1519 (O_1519,N_15981,N_17635);
nand UO_1520 (O_1520,N_15063,N_17756);
or UO_1521 (O_1521,N_18052,N_17105);
or UO_1522 (O_1522,N_18460,N_19803);
nor UO_1523 (O_1523,N_19788,N_15984);
or UO_1524 (O_1524,N_16294,N_16618);
nor UO_1525 (O_1525,N_18176,N_19172);
or UO_1526 (O_1526,N_15963,N_19169);
nor UO_1527 (O_1527,N_16847,N_17556);
and UO_1528 (O_1528,N_16415,N_16158);
nand UO_1529 (O_1529,N_18199,N_16756);
nand UO_1530 (O_1530,N_19950,N_17536);
and UO_1531 (O_1531,N_16234,N_16962);
or UO_1532 (O_1532,N_17694,N_16181);
or UO_1533 (O_1533,N_16496,N_17159);
nand UO_1534 (O_1534,N_18872,N_18734);
and UO_1535 (O_1535,N_19195,N_15726);
nor UO_1536 (O_1536,N_16595,N_18166);
or UO_1537 (O_1537,N_16839,N_18748);
nand UO_1538 (O_1538,N_18944,N_15323);
and UO_1539 (O_1539,N_19098,N_17205);
nor UO_1540 (O_1540,N_17194,N_15210);
or UO_1541 (O_1541,N_15826,N_18862);
nand UO_1542 (O_1542,N_19416,N_15035);
and UO_1543 (O_1543,N_19545,N_18607);
nor UO_1544 (O_1544,N_18692,N_16960);
nand UO_1545 (O_1545,N_17113,N_16864);
xnor UO_1546 (O_1546,N_17560,N_18022);
or UO_1547 (O_1547,N_19815,N_19414);
or UO_1548 (O_1548,N_19209,N_15511);
and UO_1549 (O_1549,N_16464,N_19667);
or UO_1550 (O_1550,N_19985,N_19343);
nand UO_1551 (O_1551,N_15661,N_16987);
nor UO_1552 (O_1552,N_16525,N_17979);
xor UO_1553 (O_1553,N_19724,N_18205);
nand UO_1554 (O_1554,N_16803,N_18841);
nand UO_1555 (O_1555,N_19892,N_19882);
or UO_1556 (O_1556,N_15476,N_15024);
or UO_1557 (O_1557,N_19718,N_19947);
nand UO_1558 (O_1558,N_17192,N_19622);
nor UO_1559 (O_1559,N_18961,N_19027);
or UO_1560 (O_1560,N_19852,N_18792);
and UO_1561 (O_1561,N_16086,N_16223);
or UO_1562 (O_1562,N_17607,N_16450);
nand UO_1563 (O_1563,N_16567,N_17292);
or UO_1564 (O_1564,N_17844,N_19189);
and UO_1565 (O_1565,N_17114,N_19961);
or UO_1566 (O_1566,N_17757,N_16917);
and UO_1567 (O_1567,N_16401,N_19325);
xnor UO_1568 (O_1568,N_19700,N_18285);
and UO_1569 (O_1569,N_18501,N_19515);
or UO_1570 (O_1570,N_18540,N_15254);
and UO_1571 (O_1571,N_18821,N_18632);
nand UO_1572 (O_1572,N_17809,N_15187);
and UO_1573 (O_1573,N_17588,N_16410);
and UO_1574 (O_1574,N_17894,N_18717);
and UO_1575 (O_1575,N_19940,N_16758);
nor UO_1576 (O_1576,N_19804,N_15109);
or UO_1577 (O_1577,N_16694,N_18926);
nand UO_1578 (O_1578,N_18110,N_17924);
and UO_1579 (O_1579,N_18980,N_16159);
and UO_1580 (O_1580,N_16495,N_15043);
nor UO_1581 (O_1581,N_15636,N_15095);
or UO_1582 (O_1582,N_18550,N_16633);
nor UO_1583 (O_1583,N_19100,N_15290);
nand UO_1584 (O_1584,N_16539,N_16068);
nand UO_1585 (O_1585,N_18553,N_19420);
nor UO_1586 (O_1586,N_16447,N_17920);
and UO_1587 (O_1587,N_17816,N_19976);
nor UO_1588 (O_1588,N_17797,N_16099);
and UO_1589 (O_1589,N_15507,N_18670);
nor UO_1590 (O_1590,N_15679,N_17581);
or UO_1591 (O_1591,N_16239,N_17744);
or UO_1592 (O_1592,N_19695,N_18787);
nor UO_1593 (O_1593,N_17687,N_17805);
and UO_1594 (O_1594,N_17062,N_18678);
nand UO_1595 (O_1595,N_18240,N_16848);
or UO_1596 (O_1596,N_19752,N_16404);
or UO_1597 (O_1597,N_19579,N_19915);
or UO_1598 (O_1598,N_16958,N_17696);
nand UO_1599 (O_1599,N_15782,N_18447);
nand UO_1600 (O_1600,N_18261,N_18039);
nor UO_1601 (O_1601,N_17926,N_19299);
or UO_1602 (O_1602,N_16481,N_19460);
nand UO_1603 (O_1603,N_19595,N_17244);
or UO_1604 (O_1604,N_17594,N_18186);
nand UO_1605 (O_1605,N_16037,N_15673);
or UO_1606 (O_1606,N_17336,N_18324);
and UO_1607 (O_1607,N_17275,N_17651);
nand UO_1608 (O_1608,N_19689,N_19023);
nand UO_1609 (O_1609,N_16248,N_17072);
nand UO_1610 (O_1610,N_19827,N_18290);
nand UO_1611 (O_1611,N_15568,N_18764);
or UO_1612 (O_1612,N_15436,N_16568);
and UO_1613 (O_1613,N_18163,N_15497);
and UO_1614 (O_1614,N_18197,N_18785);
nor UO_1615 (O_1615,N_15128,N_15156);
or UO_1616 (O_1616,N_15374,N_18503);
or UO_1617 (O_1617,N_15563,N_15906);
nand UO_1618 (O_1618,N_17773,N_16825);
and UO_1619 (O_1619,N_16857,N_18127);
nand UO_1620 (O_1620,N_17595,N_16869);
nand UO_1621 (O_1621,N_19651,N_18590);
nor UO_1622 (O_1622,N_15818,N_15202);
nand UO_1623 (O_1623,N_18466,N_17883);
or UO_1624 (O_1624,N_18191,N_19656);
nand UO_1625 (O_1625,N_15004,N_16203);
nor UO_1626 (O_1626,N_17470,N_19818);
or UO_1627 (O_1627,N_15512,N_17383);
or UO_1628 (O_1628,N_15281,N_16483);
nor UO_1629 (O_1629,N_15407,N_19244);
nor UO_1630 (O_1630,N_18665,N_18536);
nand UO_1631 (O_1631,N_16394,N_18849);
and UO_1632 (O_1632,N_16402,N_19755);
and UO_1633 (O_1633,N_19350,N_17306);
or UO_1634 (O_1634,N_17980,N_19889);
nor UO_1635 (O_1635,N_19440,N_18152);
nor UO_1636 (O_1636,N_19301,N_16445);
nor UO_1637 (O_1637,N_18299,N_17287);
nand UO_1638 (O_1638,N_19234,N_18660);
or UO_1639 (O_1639,N_17582,N_15666);
nand UO_1640 (O_1640,N_18856,N_18009);
nor UO_1641 (O_1641,N_17226,N_19267);
nor UO_1642 (O_1642,N_15286,N_15053);
nor UO_1643 (O_1643,N_17794,N_19899);
nor UO_1644 (O_1644,N_19573,N_19833);
or UO_1645 (O_1645,N_19354,N_15807);
or UO_1646 (O_1646,N_18545,N_17412);
and UO_1647 (O_1647,N_18379,N_16271);
or UO_1648 (O_1648,N_15675,N_17284);
nand UO_1649 (O_1649,N_15451,N_19486);
nand UO_1650 (O_1650,N_16880,N_18981);
nor UO_1651 (O_1651,N_18910,N_18133);
nor UO_1652 (O_1652,N_17254,N_16121);
nor UO_1653 (O_1653,N_16024,N_16046);
or UO_1654 (O_1654,N_18825,N_16796);
nand UO_1655 (O_1655,N_18212,N_19358);
nand UO_1656 (O_1656,N_15104,N_19250);
nor UO_1657 (O_1657,N_19010,N_16920);
nand UO_1658 (O_1658,N_15284,N_17005);
nand UO_1659 (O_1659,N_15258,N_15144);
and UO_1660 (O_1660,N_17772,N_16900);
and UO_1661 (O_1661,N_19134,N_15161);
or UO_1662 (O_1662,N_17322,N_17613);
nor UO_1663 (O_1663,N_18672,N_18649);
nor UO_1664 (O_1664,N_17962,N_19505);
or UO_1665 (O_1665,N_18292,N_17506);
or UO_1666 (O_1666,N_17361,N_16155);
and UO_1667 (O_1667,N_16624,N_18419);
nand UO_1668 (O_1668,N_16400,N_19761);
or UO_1669 (O_1669,N_17387,N_15552);
nor UO_1670 (O_1670,N_18528,N_19928);
nor UO_1671 (O_1671,N_18414,N_15903);
and UO_1672 (O_1672,N_16621,N_17406);
or UO_1673 (O_1673,N_17561,N_18415);
nand UO_1674 (O_1674,N_18885,N_19114);
or UO_1675 (O_1675,N_18094,N_15941);
or UO_1676 (O_1676,N_18277,N_17057);
and UO_1677 (O_1677,N_19574,N_17330);
nor UO_1678 (O_1678,N_15092,N_16083);
nor UO_1679 (O_1679,N_15300,N_18790);
nand UO_1680 (O_1680,N_17110,N_17676);
or UO_1681 (O_1681,N_15166,N_16597);
nand UO_1682 (O_1682,N_16010,N_18436);
nor UO_1683 (O_1683,N_18063,N_18070);
nor UO_1684 (O_1684,N_15304,N_19025);
or UO_1685 (O_1685,N_16883,N_19124);
nor UO_1686 (O_1686,N_15183,N_18652);
nor UO_1687 (O_1687,N_16614,N_17368);
nand UO_1688 (O_1688,N_17558,N_15592);
or UO_1689 (O_1689,N_19740,N_17095);
or UO_1690 (O_1690,N_17044,N_19418);
or UO_1691 (O_1691,N_16110,N_15114);
nor UO_1692 (O_1692,N_15720,N_18682);
nor UO_1693 (O_1693,N_15523,N_19963);
and UO_1694 (O_1694,N_17928,N_16403);
nor UO_1695 (O_1695,N_19913,N_16150);
nand UO_1696 (O_1696,N_16057,N_17959);
nor UO_1697 (O_1697,N_15213,N_18567);
nand UO_1698 (O_1698,N_17720,N_17285);
nand UO_1699 (O_1699,N_16730,N_18992);
or UO_1700 (O_1700,N_18113,N_17388);
or UO_1701 (O_1701,N_16341,N_15209);
nand UO_1702 (O_1702,N_15768,N_17997);
and UO_1703 (O_1703,N_15346,N_19626);
and UO_1704 (O_1704,N_16979,N_17298);
and UO_1705 (O_1705,N_15753,N_18683);
nor UO_1706 (O_1706,N_17511,N_19131);
nor UO_1707 (O_1707,N_19045,N_18396);
and UO_1708 (O_1708,N_17577,N_16664);
and UO_1709 (O_1709,N_18902,N_19981);
nand UO_1710 (O_1710,N_17174,N_18996);
or UO_1711 (O_1711,N_15176,N_17379);
and UO_1712 (O_1712,N_17915,N_15839);
nor UO_1713 (O_1713,N_19286,N_17024);
nand UO_1714 (O_1714,N_16662,N_17921);
nand UO_1715 (O_1715,N_17517,N_15206);
nand UO_1716 (O_1716,N_16408,N_19855);
nand UO_1717 (O_1717,N_16347,N_17474);
and UO_1718 (O_1718,N_17736,N_18211);
or UO_1719 (O_1719,N_18646,N_15752);
nand UO_1720 (O_1720,N_19386,N_15847);
or UO_1721 (O_1721,N_16413,N_18204);
or UO_1722 (O_1722,N_16548,N_19470);
nor UO_1723 (O_1723,N_19435,N_15033);
nand UO_1724 (O_1724,N_15312,N_18873);
nor UO_1725 (O_1725,N_19339,N_16387);
or UO_1726 (O_1726,N_17211,N_16990);
and UO_1727 (O_1727,N_16260,N_18576);
and UO_1728 (O_1728,N_17832,N_15587);
nor UO_1729 (O_1729,N_19683,N_19220);
nor UO_1730 (O_1730,N_17337,N_16107);
nand UO_1731 (O_1731,N_16090,N_19079);
nor UO_1732 (O_1732,N_19870,N_16801);
and UO_1733 (O_1733,N_19883,N_17130);
and UO_1734 (O_1734,N_16877,N_17865);
nand UO_1735 (O_1735,N_17014,N_17667);
nor UO_1736 (O_1736,N_19352,N_15514);
and UO_1737 (O_1737,N_18356,N_19710);
nand UO_1738 (O_1738,N_19448,N_18751);
nand UO_1739 (O_1739,N_18388,N_18490);
or UO_1740 (O_1740,N_16186,N_15549);
nand UO_1741 (O_1741,N_19773,N_15815);
or UO_1742 (O_1742,N_18853,N_19628);
and UO_1743 (O_1743,N_18126,N_18563);
or UO_1744 (O_1744,N_18257,N_15108);
nand UO_1745 (O_1745,N_16712,N_18130);
nand UO_1746 (O_1746,N_16139,N_18005);
and UO_1747 (O_1747,N_17026,N_19789);
and UO_1748 (O_1748,N_15362,N_17140);
nor UO_1749 (O_1749,N_19037,N_15828);
nand UO_1750 (O_1750,N_17955,N_17970);
or UO_1751 (O_1751,N_16722,N_19258);
nand UO_1752 (O_1752,N_17666,N_15283);
or UO_1753 (O_1753,N_18884,N_18303);
or UO_1754 (O_1754,N_19093,N_19462);
nor UO_1755 (O_1755,N_15076,N_18091);
nor UO_1756 (O_1756,N_16760,N_17639);
nand UO_1757 (O_1757,N_17239,N_17626);
nand UO_1758 (O_1758,N_19203,N_18013);
and UO_1759 (O_1759,N_17120,N_18487);
and UO_1760 (O_1760,N_17971,N_17067);
and UO_1761 (O_1761,N_18967,N_19630);
nand UO_1762 (O_1762,N_18343,N_17372);
and UO_1763 (O_1763,N_16489,N_16988);
or UO_1764 (O_1764,N_15234,N_19310);
or UO_1765 (O_1765,N_17682,N_18452);
nor UO_1766 (O_1766,N_17525,N_15513);
or UO_1767 (O_1767,N_15052,N_17055);
nor UO_1768 (O_1768,N_19338,N_18766);
or UO_1769 (O_1769,N_19021,N_19290);
or UO_1770 (O_1770,N_17196,N_19138);
nor UO_1771 (O_1771,N_15716,N_15978);
or UO_1772 (O_1772,N_16426,N_19036);
and UO_1773 (O_1773,N_17303,N_19015);
nand UO_1774 (O_1774,N_18008,N_18144);
nor UO_1775 (O_1775,N_18731,N_16742);
and UO_1776 (O_1776,N_16367,N_18840);
nor UO_1777 (O_1777,N_15131,N_19026);
nand UO_1778 (O_1778,N_18020,N_16505);
and UO_1779 (O_1779,N_18523,N_18298);
or UO_1780 (O_1780,N_16306,N_16576);
or UO_1781 (O_1781,N_17017,N_19726);
or UO_1782 (O_1782,N_15843,N_19128);
nand UO_1783 (O_1783,N_18093,N_19140);
nand UO_1784 (O_1784,N_18475,N_15481);
nor UO_1785 (O_1785,N_19542,N_18355);
nand UO_1786 (O_1786,N_19686,N_18735);
nor UO_1787 (O_1787,N_15788,N_17086);
xnor UO_1788 (O_1788,N_17746,N_16193);
or UO_1789 (O_1789,N_19534,N_15670);
and UO_1790 (O_1790,N_17565,N_18010);
nand UO_1791 (O_1791,N_17223,N_16414);
nand UO_1792 (O_1792,N_19652,N_17265);
or UO_1793 (O_1793,N_17859,N_18492);
or UO_1794 (O_1794,N_17058,N_18286);
nor UO_1795 (O_1795,N_19047,N_16933);
nor UO_1796 (O_1796,N_17165,N_17045);
nand UO_1797 (O_1797,N_16253,N_17404);
nor UO_1798 (O_1798,N_18602,N_19951);
or UO_1799 (O_1799,N_16324,N_19962);
or UO_1800 (O_1800,N_19741,N_17054);
nor UO_1801 (O_1801,N_17449,N_16222);
nand UO_1802 (O_1802,N_16913,N_15456);
nand UO_1803 (O_1803,N_18169,N_17214);
nor UO_1804 (O_1804,N_15603,N_15806);
or UO_1805 (O_1805,N_17870,N_15479);
nor UO_1806 (O_1806,N_16272,N_19333);
nand UO_1807 (O_1807,N_17606,N_18294);
nor UO_1808 (O_1808,N_16928,N_17869);
nor UO_1809 (O_1809,N_18467,N_18881);
nor UO_1810 (O_1810,N_18029,N_15528);
nand UO_1811 (O_1811,N_17960,N_19539);
nand UO_1812 (O_1812,N_16648,N_16632);
nor UO_1813 (O_1813,N_15216,N_16377);
and UO_1814 (O_1814,N_17664,N_18071);
and UO_1815 (O_1815,N_15091,N_19075);
nand UO_1816 (O_1816,N_18056,N_19457);
xor UO_1817 (O_1817,N_17230,N_15744);
nand UO_1818 (O_1818,N_15075,N_16333);
or UO_1819 (O_1819,N_18346,N_16471);
and UO_1820 (O_1820,N_19918,N_18625);
nor UO_1821 (O_1821,N_18500,N_16246);
nor UO_1822 (O_1822,N_19398,N_19864);
or UO_1823 (O_1823,N_19485,N_18904);
or UO_1824 (O_1824,N_18171,N_15419);
and UO_1825 (O_1825,N_15936,N_18208);
and UO_1826 (O_1826,N_16029,N_16881);
or UO_1827 (O_1827,N_16518,N_18640);
nand UO_1828 (O_1828,N_17170,N_16876);
or UO_1829 (O_1829,N_18995,N_17723);
nor UO_1830 (O_1830,N_15241,N_19392);
or UO_1831 (O_1831,N_15059,N_19304);
and UO_1832 (O_1832,N_17308,N_17957);
nand UO_1833 (O_1833,N_16477,N_16921);
and UO_1834 (O_1834,N_19395,N_16514);
nor UO_1835 (O_1835,N_18773,N_15050);
nor UO_1836 (O_1836,N_16968,N_18275);
nor UO_1837 (O_1837,N_16117,N_18142);
nor UO_1838 (O_1838,N_17133,N_16989);
or UO_1839 (O_1839,N_17487,N_18401);
nor UO_1840 (O_1840,N_16221,N_15640);
and UO_1841 (O_1841,N_15070,N_15696);
nand UO_1842 (O_1842,N_19635,N_15526);
or UO_1843 (O_1843,N_18437,N_16038);
nand UO_1844 (O_1844,N_16182,N_15734);
nand UO_1845 (O_1845,N_15917,N_15658);
and UO_1846 (O_1846,N_15116,N_16862);
nor UO_1847 (O_1847,N_18822,N_15859);
nand UO_1848 (O_1848,N_16753,N_15416);
nor UO_1849 (O_1849,N_19897,N_16545);
nor UO_1850 (O_1850,N_15561,N_15099);
and UO_1851 (O_1851,N_17097,N_19007);
nor UO_1852 (O_1852,N_18839,N_16973);
and UO_1853 (O_1853,N_17364,N_16817);
or UO_1854 (O_1854,N_16012,N_19057);
nor UO_1855 (O_1855,N_15771,N_19923);
or UO_1856 (O_1856,N_16356,N_19017);
nand UO_1857 (O_1857,N_19911,N_17830);
and UO_1858 (O_1858,N_16787,N_17853);
xor UO_1859 (O_1859,N_18472,N_19314);
nor UO_1860 (O_1860,N_19893,N_15341);
nand UO_1861 (O_1861,N_18935,N_17301);
and UO_1862 (O_1862,N_18368,N_17384);
nand UO_1863 (O_1863,N_17954,N_18468);
or UO_1864 (O_1864,N_17050,N_17294);
nor UO_1865 (O_1865,N_16389,N_17545);
and UO_1866 (O_1866,N_15462,N_19479);
nand UO_1867 (O_1867,N_15654,N_16809);
or UO_1868 (O_1868,N_18180,N_18080);
nand UO_1869 (O_1869,N_19050,N_16174);
or UO_1870 (O_1870,N_18431,N_16438);
and UO_1871 (O_1871,N_16735,N_15375);
or UO_1872 (O_1872,N_18367,N_18728);
and UO_1873 (O_1873,N_19184,N_16473);
or UO_1874 (O_1874,N_15271,N_15034);
nor UO_1875 (O_1875,N_15783,N_16940);
nand UO_1876 (O_1876,N_16746,N_15167);
nor UO_1877 (O_1877,N_17343,N_17689);
nor UO_1878 (O_1878,N_19987,N_15412);
or UO_1879 (O_1879,N_15408,N_18707);
and UO_1880 (O_1880,N_15193,N_15026);
or UO_1881 (O_1881,N_18815,N_15860);
nand UO_1882 (O_1882,N_17598,N_15493);
or UO_1883 (O_1883,N_16120,N_15320);
nor UO_1884 (O_1884,N_17879,N_15821);
and UO_1885 (O_1885,N_15359,N_15787);
nand UO_1886 (O_1886,N_16005,N_16339);
and UO_1887 (O_1887,N_16649,N_16089);
xnor UO_1888 (O_1888,N_17208,N_15243);
and UO_1889 (O_1889,N_17829,N_17632);
and UO_1890 (O_1890,N_15604,N_16564);
and UO_1891 (O_1891,N_15868,N_16217);
nand UO_1892 (O_1892,N_16789,N_18255);
nor UO_1893 (O_1893,N_16637,N_18249);
nor UO_1894 (O_1894,N_19934,N_15900);
nor UO_1895 (O_1895,N_15834,N_16105);
and UO_1896 (O_1896,N_17533,N_15280);
nor UO_1897 (O_1897,N_19403,N_15383);
or UO_1898 (O_1898,N_18326,N_16268);
and UO_1899 (O_1899,N_19160,N_16386);
or UO_1900 (O_1900,N_16040,N_18635);
or UO_1901 (O_1901,N_18370,N_19678);
or UO_1902 (O_1902,N_15329,N_16898);
nor UO_1903 (O_1903,N_16724,N_16191);
and UO_1904 (O_1904,N_18331,N_17849);
nor UO_1905 (O_1905,N_15170,N_16638);
and UO_1906 (O_1906,N_17671,N_18620);
nand UO_1907 (O_1907,N_17147,N_17040);
nand UO_1908 (O_1908,N_16293,N_17861);
and UO_1909 (O_1909,N_15025,N_15615);
nand UO_1910 (O_1910,N_18076,N_16130);
nand UO_1911 (O_1911,N_16328,N_16792);
nand UO_1912 (O_1912,N_19364,N_16440);
and UO_1913 (O_1913,N_15299,N_17813);
and UO_1914 (O_1914,N_15635,N_19356);
and UO_1915 (O_1915,N_19243,N_16922);
or UO_1916 (O_1916,N_16726,N_17750);
nor UO_1917 (O_1917,N_16020,N_16571);
nor UO_1918 (O_1918,N_18234,N_18829);
or UO_1919 (O_1919,N_17751,N_16017);
or UO_1920 (O_1920,N_19041,N_18443);
and UO_1921 (O_1921,N_16133,N_16666);
and UO_1922 (O_1922,N_16138,N_19584);
nor UO_1923 (O_1923,N_15005,N_16603);
nor UO_1924 (O_1924,N_16845,N_15608);
nor UO_1925 (O_1925,N_19496,N_19270);
nand UO_1926 (O_1926,N_15058,N_17922);
or UO_1927 (O_1927,N_16019,N_17039);
or UO_1928 (O_1928,N_16265,N_16494);
or UO_1929 (O_1929,N_17622,N_15871);
and UO_1930 (O_1930,N_18015,N_17847);
or UO_1931 (O_1931,N_16200,N_19956);
nand UO_1932 (O_1932,N_15809,N_15699);
or UO_1933 (O_1933,N_19867,N_18122);
or UO_1934 (O_1934,N_16503,N_17660);
or UO_1935 (O_1935,N_18215,N_16956);
and UO_1936 (O_1936,N_15179,N_18681);
and UO_1937 (O_1937,N_15401,N_19249);
or UO_1938 (O_1938,N_17390,N_18756);
and UO_1939 (O_1939,N_18145,N_15337);
or UO_1940 (O_1940,N_17252,N_15564);
nand UO_1941 (O_1941,N_15352,N_19674);
and UO_1942 (O_1942,N_16634,N_16596);
and UO_1943 (O_1943,N_15140,N_16617);
nor UO_1944 (O_1944,N_18230,N_16095);
nor UO_1945 (O_1945,N_19729,N_15888);
or UO_1946 (O_1946,N_18921,N_15001);
nand UO_1947 (O_1947,N_17637,N_15257);
nand UO_1948 (O_1948,N_17212,N_19424);
or UO_1949 (O_1949,N_18987,N_19952);
nor UO_1950 (O_1950,N_18376,N_19464);
and UO_1951 (O_1951,N_16574,N_18700);
and UO_1952 (O_1952,N_17156,N_17261);
nor UO_1953 (O_1953,N_17734,N_16167);
nor UO_1954 (O_1954,N_19834,N_15630);
nand UO_1955 (O_1955,N_18481,N_16302);
and UO_1956 (O_1956,N_15811,N_18195);
or UO_1957 (O_1957,N_19698,N_16949);
nor UO_1958 (O_1958,N_16490,N_16021);
or UO_1959 (O_1959,N_18566,N_17990);
or UO_1960 (O_1960,N_19553,N_19053);
nand UO_1961 (O_1961,N_17291,N_19605);
nor UO_1962 (O_1962,N_19636,N_16423);
nor UO_1963 (O_1963,N_18455,N_19256);
or UO_1964 (O_1964,N_15849,N_15186);
or UO_1965 (O_1965,N_17559,N_16670);
nor UO_1966 (O_1966,N_17976,N_15231);
nor UO_1967 (O_1967,N_16562,N_15069);
and UO_1968 (O_1968,N_17731,N_15631);
nor UO_1969 (O_1969,N_18411,N_16259);
and UO_1970 (O_1970,N_18192,N_15030);
nor UO_1971 (O_1971,N_15774,N_18820);
nor UO_1972 (O_1972,N_16779,N_15130);
and UO_1973 (O_1973,N_18099,N_16465);
nand UO_1974 (O_1974,N_19808,N_19188);
or UO_1975 (O_1975,N_18744,N_19570);
nand UO_1976 (O_1976,N_16237,N_18470);
nor UO_1977 (O_1977,N_19297,N_16992);
and UO_1978 (O_1978,N_15208,N_17993);
nor UO_1979 (O_1979,N_19793,N_18542);
or UO_1980 (O_1980,N_19779,N_15998);
and UO_1981 (O_1981,N_17500,N_18688);
and UO_1982 (O_1982,N_16918,N_15222);
nor UO_1983 (O_1983,N_15796,N_18218);
nand UO_1984 (O_1984,N_19066,N_15146);
or UO_1985 (O_1985,N_16732,N_15738);
and UO_1986 (O_1986,N_16358,N_18032);
nand UO_1987 (O_1987,N_19654,N_18759);
nand UO_1988 (O_1988,N_17144,N_19351);
nand UO_1989 (O_1989,N_19575,N_15441);
nand UO_1990 (O_1990,N_16343,N_17112);
or UO_1991 (O_1991,N_18024,N_19837);
and UO_1992 (O_1992,N_16227,N_18687);
or UO_1993 (O_1993,N_18749,N_16725);
nor UO_1994 (O_1994,N_15246,N_17550);
and UO_1995 (O_1995,N_17638,N_15729);
and UO_1996 (O_1996,N_16785,N_19847);
and UO_1997 (O_1997,N_17674,N_16165);
or UO_1998 (O_1998,N_19824,N_15798);
nor UO_1999 (O_1999,N_18506,N_16319);
and UO_2000 (O_2000,N_18319,N_17649);
nand UO_2001 (O_2001,N_17011,N_16709);
and UO_2002 (O_2002,N_19887,N_18387);
nor UO_2003 (O_2003,N_19274,N_16383);
or UO_2004 (O_2004,N_18016,N_15405);
and UO_2005 (O_2005,N_18739,N_16654);
nand UO_2006 (O_2006,N_15172,N_17874);
xor UO_2007 (O_2007,N_16878,N_17101);
and UO_2008 (O_2008,N_16700,N_16478);
or UO_2009 (O_2009,N_17332,N_19905);
and UO_2010 (O_2010,N_16515,N_15574);
xor UO_2011 (O_2011,N_17888,N_17012);
and UO_2012 (O_2012,N_15397,N_19296);
and UO_2013 (O_2013,N_19384,N_17240);
nor UO_2014 (O_2014,N_17624,N_18047);
nor UO_2015 (O_2015,N_16684,N_19146);
xor UO_2016 (O_2016,N_15065,N_15014);
and UO_2017 (O_2017,N_16930,N_18172);
nand UO_2018 (O_2018,N_19322,N_17210);
nand UO_2019 (O_2019,N_15733,N_19162);
or UO_2020 (O_2020,N_18711,N_19706);
nor UO_2021 (O_2021,N_19693,N_17726);
or UO_2022 (O_2022,N_18618,N_18446);
or UO_2023 (O_2023,N_16349,N_16030);
and UO_2024 (O_2024,N_15634,N_16273);
and UO_2025 (O_2025,N_19843,N_17158);
or UO_2026 (O_2026,N_17415,N_19715);
nand UO_2027 (O_2027,N_16350,N_19173);
and UO_2028 (O_2028,N_17436,N_17891);
and UO_2029 (O_2029,N_17142,N_16691);
and UO_2030 (O_2030,N_16204,N_18594);
nand UO_2031 (O_2031,N_15856,N_18767);
nor UO_2032 (O_2032,N_17307,N_19646);
nand UO_2033 (O_2033,N_16824,N_15443);
and UO_2034 (O_2034,N_18293,N_15642);
nand UO_2035 (O_2035,N_18957,N_16837);
or UO_2036 (O_2036,N_17366,N_16252);
or UO_2037 (O_2037,N_18908,N_15522);
and UO_2038 (O_2038,N_18591,N_17377);
or UO_2039 (O_2039,N_18922,N_18421);
nor UO_2040 (O_2040,N_16035,N_15032);
nand UO_2041 (O_2041,N_18810,N_17108);
or UO_2042 (O_2042,N_17483,N_16168);
nor UO_2043 (O_2043,N_19228,N_19472);
nor UO_2044 (O_2044,N_18869,N_19540);
or UO_2045 (O_2045,N_19665,N_18000);
nand UO_2046 (O_2046,N_16734,N_16487);
nand UO_2047 (O_2047,N_17608,N_16808);
or UO_2048 (O_2048,N_17032,N_19816);
and UO_2049 (O_2049,N_18585,N_17702);
nor UO_2050 (O_2050,N_16769,N_15238);
or UO_2051 (O_2051,N_19601,N_17312);
and UO_2052 (O_2052,N_17784,N_19771);
or UO_2053 (O_2053,N_19801,N_18301);
or UO_2054 (O_2054,N_17408,N_16513);
nand UO_2055 (O_2055,N_19785,N_18459);
nor UO_2056 (O_2056,N_18771,N_16039);
and UO_2057 (O_2057,N_19901,N_16946);
nand UO_2058 (O_2058,N_16425,N_17636);
nand UO_2059 (O_2059,N_19413,N_16094);
and UO_2060 (O_2060,N_16682,N_17557);
and UO_2061 (O_2061,N_15450,N_19588);
and UO_2062 (O_2062,N_17476,N_18544);
nor UO_2063 (O_2063,N_15378,N_18592);
and UO_2064 (O_2064,N_18154,N_19383);
nor UO_2065 (O_2065,N_18187,N_19919);
nand UO_2066 (O_2066,N_15142,N_17838);
nor UO_2067 (O_2067,N_15433,N_15874);
and UO_2068 (O_2068,N_15500,N_18791);
and UO_2069 (O_2069,N_16932,N_19634);
nand UO_2070 (O_2070,N_15080,N_19629);
or UO_2071 (O_2071,N_18948,N_19450);
nand UO_2072 (O_2072,N_15740,N_18658);
and UO_2073 (O_2073,N_17661,N_16646);
and UO_2074 (O_2074,N_15982,N_15977);
and UO_2075 (O_2075,N_15423,N_18919);
nand UO_2076 (O_2076,N_17329,N_15064);
nand UO_2077 (O_2077,N_19412,N_17346);
nand UO_2078 (O_2078,N_18006,N_16757);
or UO_2079 (O_2079,N_19167,N_18894);
nand UO_2080 (O_2080,N_18686,N_17625);
or UO_2081 (O_2081,N_17274,N_17209);
nor UO_2082 (O_2082,N_19520,N_15169);
or UO_2083 (O_2083,N_19120,N_17249);
and UO_2084 (O_2084,N_16274,N_18906);
nand UO_2085 (O_2085,N_18636,N_17570);
and UO_2086 (O_2086,N_15845,N_17154);
or UO_2087 (O_2087,N_16420,N_18896);
nor UO_2088 (O_2088,N_18928,N_17399);
or UO_2089 (O_2089,N_18408,N_19439);
and UO_2090 (O_2090,N_16675,N_18316);
nor UO_2091 (O_2091,N_16243,N_18770);
or UO_2092 (O_2092,N_15153,N_16357);
nor UO_2093 (O_2093,N_16519,N_15438);
and UO_2094 (O_2094,N_16374,N_17151);
and UO_2095 (O_2095,N_16376,N_17141);
nor UO_2096 (O_2096,N_15377,N_15929);
and UO_2097 (O_2097,N_19331,N_18892);
nand UO_2098 (O_2098,N_16032,N_18141);
or UO_2099 (O_2099,N_15185,N_19946);
nor UO_2100 (O_2100,N_17206,N_19538);
nand UO_2101 (O_2101,N_17949,N_15586);
and UO_2102 (O_2102,N_17820,N_19734);
nand UO_2103 (O_2103,N_16114,N_19028);
nor UO_2104 (O_2104,N_17423,N_19181);
or UO_2105 (O_2105,N_15084,N_18279);
and UO_2106 (O_2106,N_15882,N_15387);
nor UO_2107 (O_2107,N_17462,N_19446);
nor UO_2108 (O_2108,N_15321,N_19177);
or UO_2109 (O_2109,N_15569,N_17766);
nand UO_2110 (O_2110,N_18626,N_18671);
nor UO_2111 (O_2111,N_16871,N_15143);
nand UO_2112 (O_2112,N_16577,N_15157);
xnor UO_2113 (O_2113,N_18685,N_15475);
xnor UO_2114 (O_2114,N_17053,N_19068);
and UO_2115 (O_2115,N_18007,N_19344);
nand UO_2116 (O_2116,N_18586,N_15203);
nor UO_2117 (O_2117,N_18248,N_15565);
nor UO_2118 (O_2118,N_15602,N_15663);
and UO_2119 (O_2119,N_18307,N_19480);
nand UO_2120 (O_2120,N_17815,N_18321);
and UO_2121 (O_2121,N_18190,N_15801);
nand UO_2122 (O_2122,N_18648,N_17677);
nor UO_2123 (O_2123,N_19616,N_18769);
nor UO_2124 (O_2124,N_16065,N_19456);
and UO_2125 (O_2125,N_18850,N_15599);
nand UO_2126 (O_2126,N_18313,N_16314);
and UO_2127 (O_2127,N_19175,N_15335);
and UO_2128 (O_2128,N_15417,N_15509);
nand UO_2129 (O_2129,N_19101,N_16508);
nand UO_2130 (O_2130,N_19600,N_19560);
and UO_2131 (O_2131,N_15264,N_17221);
or UO_2132 (O_2132,N_15894,N_16137);
nor UO_2133 (O_2133,N_17818,N_18416);
and UO_2134 (O_2134,N_16768,N_19525);
and UO_2135 (O_2135,N_15930,N_15727);
or UO_2136 (O_2136,N_15478,N_17673);
or UO_2137 (O_2137,N_17047,N_17451);
nor UO_2138 (O_2138,N_17342,N_15883);
nor UO_2139 (O_2139,N_18861,N_17515);
or UO_2140 (O_2140,N_19020,N_16399);
nor UO_2141 (O_2141,N_19711,N_17215);
nand UO_2142 (O_2142,N_18796,N_16312);
nor UO_2143 (O_2143,N_16197,N_17837);
nor UO_2144 (O_2144,N_18384,N_16697);
or UO_2145 (O_2145,N_18174,N_19105);
nor UO_2146 (O_2146,N_17732,N_16285);
nand UO_2147 (O_2147,N_15339,N_19894);
nor UO_2148 (O_2148,N_19645,N_18830);
nand UO_2149 (O_2149,N_18246,N_17033);
and UO_2150 (O_2150,N_15646,N_17052);
nand UO_2151 (O_2151,N_19251,N_18752);
nand UO_2152 (O_2152,N_17473,N_16554);
nor UO_2153 (O_2153,N_17759,N_17693);
nand UO_2154 (O_2154,N_17395,N_17152);
nor UO_2155 (O_2155,N_15797,N_16156);
nand UO_2156 (O_2156,N_18846,N_16009);
nand UO_2157 (O_2157,N_17359,N_15498);
and UO_2158 (O_2158,N_16957,N_18827);
and UO_2159 (O_2159,N_17807,N_19769);
nor UO_2160 (O_2160,N_19797,N_17858);
and UO_2161 (O_2161,N_16184,N_19884);
nand UO_2162 (O_2162,N_15386,N_17668);
nor UO_2163 (O_2163,N_15047,N_19590);
or UO_2164 (O_2164,N_15914,N_16366);
xnor UO_2165 (O_2165,N_17546,N_15473);
or UO_2166 (O_2166,N_15041,N_19207);
and UO_2167 (O_2167,N_17010,N_18870);
and UO_2168 (O_2168,N_19593,N_16951);
or UO_2169 (O_2169,N_15667,N_17246);
nor UO_2170 (O_2170,N_15171,N_19357);
nand UO_2171 (O_2171,N_16125,N_19197);
and UO_2172 (O_2172,N_17299,N_18473);
and UO_2173 (O_2173,N_19618,N_18250);
and UO_2174 (O_2174,N_18779,N_16225);
or UO_2175 (O_2175,N_17173,N_17074);
or UO_2176 (O_2176,N_16372,N_16723);
nor UO_2177 (O_2177,N_17316,N_19458);
or UO_2178 (O_2178,N_15275,N_18555);
nand UO_2179 (O_2179,N_16639,N_19059);
nand UO_2180 (O_2180,N_16551,N_16882);
or UO_2181 (O_2181,N_18936,N_19183);
and UO_2182 (O_2182,N_17522,N_15486);
nor UO_2183 (O_2183,N_19038,N_16850);
nand UO_2184 (O_2184,N_15891,N_17730);
nand UO_2185 (O_2185,N_17790,N_18097);
nand UO_2186 (O_2186,N_17872,N_16810);
xnor UO_2187 (O_2187,N_18479,N_16249);
or UO_2188 (O_2188,N_15127,N_19640);
or UO_2189 (O_2189,N_18975,N_18562);
nand UO_2190 (O_2190,N_15534,N_19498);
or UO_2191 (O_2191,N_16765,N_15093);
or UO_2192 (O_2192,N_17907,N_17356);
and UO_2193 (O_2193,N_15342,N_16016);
and UO_2194 (O_2194,N_15217,N_17713);
and UO_2195 (O_2195,N_16407,N_16264);
nand UO_2196 (O_2196,N_16382,N_16728);
or UO_2197 (O_2197,N_17203,N_16790);
or UO_2198 (O_2198,N_17705,N_17591);
nor UO_2199 (O_2199,N_18365,N_16393);
or UO_2200 (O_2200,N_16499,N_16831);
nand UO_2201 (O_2201,N_17092,N_19255);
nor UO_2202 (O_2202,N_15394,N_17585);
and UO_2203 (O_2203,N_15277,N_17827);
or UO_2204 (O_2204,N_19677,N_15353);
and UO_2205 (O_2205,N_16134,N_17429);
nor UO_2206 (O_2206,N_18525,N_19428);
or UO_2207 (O_2207,N_17648,N_15020);
nand UO_2208 (O_2208,N_18188,N_16308);
and UO_2209 (O_2209,N_18760,N_18463);
nor UO_2210 (O_2210,N_18351,N_16101);
and UO_2211 (O_2211,N_16442,N_16433);
xnor UO_2212 (O_2212,N_19551,N_17227);
and UO_2213 (O_2213,N_16310,N_16773);
and UO_2214 (O_2214,N_17808,N_18722);
nor UO_2215 (O_2215,N_18162,N_18164);
and UO_2216 (O_2216,N_18330,N_19198);
and UO_2217 (O_2217,N_18998,N_19554);
and UO_2218 (O_2218,N_16685,N_15294);
nor UO_2219 (O_2219,N_17310,N_19081);
nand UO_2220 (O_2220,N_15123,N_18838);
or UO_2221 (O_2221,N_15985,N_16355);
nor UO_2222 (O_2222,N_18352,N_19329);
and UO_2223 (O_2223,N_18889,N_19362);
and UO_2224 (O_2224,N_17362,N_18878);
or UO_2225 (O_2225,N_18258,N_16151);
nor UO_2226 (O_2226,N_15000,N_18963);
and UO_2227 (O_2227,N_19293,N_17286);
nand UO_2228 (O_2228,N_18227,N_17405);
nand UO_2229 (O_2229,N_19699,N_18427);
nand UO_2230 (O_2230,N_16535,N_15612);
or UO_2231 (O_2231,N_17289,N_16458);
nand UO_2232 (O_2232,N_19668,N_16145);
nor UO_2233 (O_2233,N_18628,N_19750);
nand UO_2234 (O_2234,N_16323,N_17662);
nand UO_2235 (O_2235,N_16749,N_18977);
nor UO_2236 (O_2236,N_19074,N_18656);
nand UO_2237 (O_2237,N_15823,N_18942);
and UO_2238 (O_2238,N_19385,N_15449);
nand UO_2239 (O_2239,N_18571,N_15134);
nor UO_2240 (O_2240,N_17132,N_17857);
and UO_2241 (O_2241,N_17719,N_17505);
nand UO_2242 (O_2242,N_17260,N_19459);
nor UO_2243 (O_2243,N_15019,N_15710);
nand UO_2244 (O_2244,N_19529,N_15680);
nor UO_2245 (O_2245,N_18879,N_17478);
nor UO_2246 (O_2246,N_19792,N_17704);
nor UO_2247 (O_2247,N_18934,N_19609);
and UO_2248 (O_2248,N_17905,N_19455);
nor UO_2249 (O_2249,N_18650,N_19284);
and UO_2250 (O_2250,N_18485,N_16022);
and UO_2251 (O_2251,N_18391,N_16112);
or UO_2252 (O_2252,N_17983,N_16767);
and UO_2253 (O_2253,N_18690,N_19765);
or UO_2254 (O_2254,N_16867,N_18457);
nor UO_2255 (O_2255,N_16604,N_15669);
and UO_2256 (O_2256,N_19372,N_19949);
nand UO_2257 (O_2257,N_18196,N_15431);
nor UO_2258 (O_2258,N_17235,N_17277);
or UO_2259 (O_2259,N_16829,N_15444);
or UO_2260 (O_2260,N_19206,N_17987);
or UO_2261 (O_2261,N_17840,N_17633);
nor UO_2262 (O_2262,N_18570,N_15961);
or UO_2263 (O_2263,N_18238,N_16180);
and UO_2264 (O_2264,N_16569,N_19604);
nor UO_2265 (O_2265,N_18733,N_17085);
nor UO_2266 (O_2266,N_17179,N_16611);
nand UO_2267 (O_2267,N_15884,N_17367);
nor UO_2268 (O_2268,N_17176,N_15822);
or UO_2269 (O_2269,N_16286,N_19967);
and UO_2270 (O_2270,N_15580,N_16460);
nor UO_2271 (O_2271,N_15291,N_17701);
nand UO_2272 (O_2272,N_15717,N_19672);
nand UO_2273 (O_2273,N_18209,N_19451);
nor UO_2274 (O_2274,N_18693,N_19449);
nand UO_2275 (O_2275,N_18828,N_15633);
nor UO_2276 (O_2276,N_18339,N_18611);
and UO_2277 (O_2277,N_15824,N_18888);
and UO_2278 (O_2278,N_17251,N_16752);
and UO_2279 (O_2279,N_15693,N_19165);
or UO_2280 (O_2280,N_16418,N_15389);
and UO_2281 (O_2281,N_15778,N_16889);
nor UO_2282 (O_2282,N_15470,N_19592);
or UO_2283 (O_2283,N_15293,N_18471);
nor UO_2284 (O_2284,N_15677,N_18081);
nor UO_2285 (O_2285,N_16379,N_19607);
nor UO_2286 (O_2286,N_18837,N_18038);
or UO_2287 (O_2287,N_15819,N_17586);
nor UO_2288 (O_2288,N_15760,N_15228);
nand UO_2289 (O_2289,N_18631,N_15031);
or UO_2290 (O_2290,N_18608,N_19090);
nor UO_2291 (O_2291,N_15132,N_16964);
and UO_2292 (O_2292,N_17124,N_16954);
or UO_2293 (O_2293,N_18668,N_15904);
nor UO_2294 (O_2294,N_18634,N_18580);
and UO_2295 (O_2295,N_18433,N_19499);
nor UO_2296 (O_2296,N_15129,N_15039);
and UO_2297 (O_2297,N_17187,N_15970);
and UO_2298 (O_2298,N_18737,N_18621);
or UO_2299 (O_2299,N_17524,N_15055);
and UO_2300 (O_2300,N_19807,N_16986);
or UO_2301 (O_2301,N_18185,N_19200);
or UO_2302 (O_2302,N_18880,N_17182);
nand UO_2303 (O_2303,N_16284,N_19222);
nor UO_2304 (O_2304,N_19914,N_16352);
nor UO_2305 (O_2305,N_18589,N_18984);
nand UO_2306 (O_2306,N_18582,N_19957);
and UO_2307 (O_2307,N_15367,N_15207);
or UO_2308 (O_2308,N_16018,N_19917);
nor UO_2309 (O_2309,N_19509,N_19896);
or UO_2310 (O_2310,N_19155,N_16978);
nand UO_2311 (O_2311,N_18574,N_19035);
nand UO_2312 (O_2312,N_18317,N_16446);
and UO_2313 (O_2313,N_18210,N_18202);
nor UO_2314 (O_2314,N_15616,N_15812);
and UO_2315 (O_2315,N_19410,N_19871);
nand UO_2316 (O_2316,N_19958,N_19084);
or UO_2317 (O_2317,N_17161,N_15390);
nand UO_2318 (O_2318,N_17442,N_18451);
nand UO_2319 (O_2319,N_19202,N_17834);
nor UO_2320 (O_2320,N_15887,N_15921);
nand UO_2321 (O_2321,N_16280,N_18413);
nand UO_2322 (O_2322,N_16006,N_17160);
and UO_2323 (O_2323,N_17360,N_15087);
and UO_2324 (O_2324,N_18736,N_15381);
nand UO_2325 (O_2325,N_17502,N_19253);
nor UO_2326 (O_2326,N_19714,N_17326);
and UO_2327 (O_2327,N_17826,N_15769);
and UO_2328 (O_2328,N_15759,N_16416);
nand UO_2329 (O_2329,N_16344,N_15875);
or UO_2330 (O_2330,N_19049,N_18219);
and UO_2331 (O_2331,N_18474,N_17513);
or UO_2332 (O_2332,N_19879,N_16644);
nand UO_2333 (O_2333,N_19663,N_19193);
nor UO_2334 (O_2334,N_16201,N_19109);
nor UO_2335 (O_2335,N_17553,N_15021);
and UO_2336 (O_2336,N_18730,N_15750);
or UO_2337 (O_2337,N_19003,N_19252);
or UO_2338 (O_2338,N_19641,N_16819);
nand UO_2339 (O_2339,N_18645,N_18059);
or UO_2340 (O_2340,N_19335,N_18930);
and UO_2341 (O_2341,N_18867,N_15949);
or UO_2342 (O_2342,N_15948,N_18377);
nor UO_2343 (O_2343,N_19261,N_18807);
nand UO_2344 (O_2344,N_15060,N_16123);
or UO_2345 (O_2345,N_15991,N_15266);
or UO_2346 (O_2346,N_19302,N_16033);
and UO_2347 (O_2347,N_16369,N_15650);
nor UO_2348 (O_2348,N_17930,N_17171);
nor UO_2349 (O_2349,N_16887,N_16218);
and UO_2350 (O_2350,N_16363,N_16003);
nor UO_2351 (O_2351,N_15094,N_19512);
nand UO_2352 (O_2352,N_17793,N_19196);
nor UO_2353 (O_2353,N_18606,N_16863);
nor UO_2354 (O_2354,N_15664,N_18823);
or UO_2355 (O_2355,N_18226,N_19316);
nor UO_2356 (O_2356,N_16679,N_16716);
nand UO_2357 (O_2357,N_15067,N_17351);
nand UO_2358 (O_2358,N_16631,N_19518);
or UO_2359 (O_2359,N_19849,N_15086);
xor UO_2360 (O_2360,N_15253,N_15344);
nand UO_2361 (O_2361,N_15358,N_18336);
or UO_2362 (O_2362,N_19774,N_18887);
nand UO_2363 (O_2363,N_19501,N_18705);
and UO_2364 (O_2364,N_16431,N_17479);
or UO_2365 (O_2365,N_18972,N_18643);
and UO_2366 (O_2366,N_15235,N_19295);
nor UO_2367 (O_2367,N_15265,N_19802);
and UO_2368 (O_2368,N_15614,N_18366);
nand UO_2369 (O_2369,N_16198,N_16772);
or UO_2370 (O_2370,N_17122,N_18633);
or UO_2371 (O_2371,N_18599,N_19767);
and UO_2372 (O_2372,N_16814,N_15306);
nor UO_2373 (O_2373,N_15452,N_18949);
and UO_2374 (O_2374,N_18937,N_15477);
or UO_2375 (O_2375,N_17741,N_16063);
nand UO_2376 (O_2376,N_17754,N_18903);
nor UO_2377 (O_2377,N_18430,N_17982);
nand UO_2378 (O_2378,N_19851,N_17184);
nand UO_2379 (O_2379,N_17015,N_16297);
or UO_2380 (O_2380,N_17314,N_18338);
and UO_2381 (O_2381,N_17018,N_15597);
and UO_2382 (O_2382,N_15987,N_16950);
and UO_2383 (O_2383,N_16718,N_17233);
and UO_2384 (O_2384,N_16524,N_15403);
nand UO_2385 (O_2385,N_17103,N_16233);
nor UO_2386 (O_2386,N_17801,N_15562);
and UO_2387 (O_2387,N_17575,N_18189);
or UO_2388 (O_2388,N_16533,N_19205);
and UO_2389 (O_2389,N_18399,N_15200);
or UO_2390 (O_2390,N_18768,N_16072);
and UO_2391 (O_2391,N_19614,N_19939);
nand UO_2392 (O_2392,N_15472,N_15546);
nand UO_2393 (O_2393,N_16751,N_19728);
or UO_2394 (O_2394,N_16435,N_16422);
and UO_2395 (O_2395,N_18217,N_16424);
nand UO_2396 (O_2396,N_15687,N_15066);
nand UO_2397 (O_2397,N_15955,N_18675);
or UO_2398 (O_2398,N_17762,N_17304);
nor UO_2399 (O_2399,N_16994,N_18913);
nor UO_2400 (O_2400,N_19857,N_19032);
and UO_2401 (O_2401,N_18108,N_19391);
nand UO_2402 (O_2402,N_19623,N_19369);
and UO_2403 (O_2403,N_19968,N_16761);
nand UO_2404 (O_2404,N_19336,N_16506);
xor UO_2405 (O_2405,N_17093,N_18917);
and UO_2406 (O_2406,N_19760,N_15435);
or UO_2407 (O_2407,N_15992,N_17409);
nor UO_2408 (O_2408,N_18811,N_16934);
and UO_2409 (O_2409,N_19376,N_15855);
or UO_2410 (O_2410,N_17900,N_18105);
nor UO_2411 (O_2411,N_18616,N_17851);
nand UO_2412 (O_2412,N_16283,N_17925);
or UO_2413 (O_2413,N_16316,N_15263);
nand UO_2414 (O_2414,N_17087,N_15559);
nand UO_2415 (O_2415,N_15317,N_16172);
and UO_2416 (O_2416,N_19199,N_16074);
nand UO_2417 (O_2417,N_16602,N_17465);
and UO_2418 (O_2418,N_15781,N_15723);
and UO_2419 (O_2419,N_18920,N_19969);
and UO_2420 (O_2420,N_15125,N_19965);
and UO_2421 (O_2421,N_18783,N_17162);
xor UO_2422 (O_2422,N_18050,N_18461);
nand UO_2423 (O_2423,N_16665,N_18666);
or UO_2424 (O_2424,N_16194,N_17835);
and UO_2425 (O_2425,N_16998,N_16452);
nand UO_2426 (O_2426,N_17843,N_17315);
or UO_2427 (O_2427,N_19019,N_19836);
or UO_2428 (O_2428,N_17620,N_17445);
or UO_2429 (O_2429,N_17507,N_16619);
and UO_2430 (O_2430,N_18233,N_19895);
nor UO_2431 (O_2431,N_15672,N_19644);
nor UO_2432 (O_2432,N_17824,N_16696);
nand UO_2433 (O_2433,N_19421,N_16098);
nor UO_2434 (O_2434,N_17327,N_15800);
nor UO_2435 (O_2435,N_19998,N_19430);
and UO_2436 (O_2436,N_16428,N_19548);
xnor UO_2437 (O_2437,N_15459,N_15248);
nand UO_2438 (O_2438,N_15939,N_15538);
or UO_2439 (O_2439,N_18548,N_18593);
and UO_2440 (O_2440,N_15922,N_16532);
and UO_2441 (O_2441,N_19810,N_15718);
or UO_2442 (O_2442,N_19390,N_15632);
nor UO_2443 (O_2443,N_16208,N_16811);
nand UO_2444 (O_2444,N_18951,N_17952);
and UO_2445 (O_2445,N_17944,N_18214);
or UO_2446 (O_2446,N_19791,N_15396);
and UO_2447 (O_2447,N_16163,N_18228);
nor UO_2448 (O_2448,N_17013,N_18835);
or UO_2449 (O_2449,N_15644,N_15242);
and UO_2450 (O_2450,N_15737,N_17048);
or UO_2451 (O_2451,N_17076,N_17031);
nand UO_2452 (O_2452,N_18442,N_18323);
nor UO_2453 (O_2453,N_16516,N_16056);
and UO_2454 (O_2454,N_19559,N_19780);
nand UO_2455 (O_2455,N_19363,N_15267);
nor UO_2456 (O_2456,N_17421,N_19112);
and UO_2457 (O_2457,N_19438,N_19880);
nand UO_2458 (O_2458,N_19309,N_19453);
and UO_2459 (O_2459,N_15706,N_17333);
and UO_2460 (O_2460,N_19784,N_19642);
nand UO_2461 (O_2461,N_15637,N_16397);
nor UO_2462 (O_2462,N_17538,N_16834);
nor UO_2463 (O_2463,N_18315,N_18680);
nand UO_2464 (O_2464,N_19102,N_16815);
nand UO_2465 (O_2465,N_15343,N_17454);
nand UO_2466 (O_2466,N_17656,N_19649);
and UO_2467 (O_2467,N_16147,N_16421);
nand UO_2468 (O_2468,N_15270,N_18001);
and UO_2469 (O_2469,N_16565,N_17410);
or UO_2470 (O_2470,N_17535,N_16668);
nand UO_2471 (O_2471,N_16462,N_19402);
nand UO_2472 (O_2472,N_18282,N_17698);
or UO_2473 (O_2473,N_18017,N_16202);
nand UO_2474 (O_2474,N_16653,N_18905);
or UO_2475 (O_2475,N_15040,N_16802);
or UO_2476 (O_2476,N_16781,N_15715);
and UO_2477 (O_2477,N_19888,N_17564);
and UO_2478 (O_2478,N_15012,N_17908);
or UO_2479 (O_2479,N_16327,N_17079);
or UO_2480 (O_2480,N_18529,N_17243);
nand UO_2481 (O_2481,N_16563,N_18137);
and UO_2482 (O_2482,N_17914,N_19201);
and UO_2483 (O_2483,N_17385,N_17998);
or UO_2484 (O_2484,N_18988,N_15237);
and UO_2485 (O_2485,N_18444,N_19190);
nand UO_2486 (O_2486,N_18976,N_19235);
or UO_2487 (O_2487,N_15850,N_18732);
nor UO_2488 (O_2488,N_19926,N_17480);
nand UO_2489 (O_2489,N_17236,N_17125);
or UO_2490 (O_2490,N_16737,N_17509);
nand UO_2491 (O_2491,N_17183,N_19763);
nand UO_2492 (O_2492,N_18159,N_16512);
nand UO_2493 (O_2493,N_19597,N_19813);
and UO_2494 (O_2494,N_15540,N_15653);
or UO_2495 (O_2495,N_17519,N_17882);
or UO_2496 (O_2496,N_16778,N_19342);
nand UO_2497 (O_2497,N_17919,N_19611);
or UO_2498 (O_2498,N_19473,N_15048);
or UO_2499 (O_2499,N_17866,N_16528);
endmodule