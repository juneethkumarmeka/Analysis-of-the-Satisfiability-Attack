module basic_1500_15000_2000_15_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
or U0 (N_0,In_870,In_1465);
nand U1 (N_1,In_1310,In_1436);
nor U2 (N_2,In_430,In_481);
xnor U3 (N_3,In_282,In_1418);
nand U4 (N_4,In_857,In_736);
nand U5 (N_5,In_807,In_921);
and U6 (N_6,In_544,In_815);
and U7 (N_7,In_436,In_1215);
xnor U8 (N_8,In_153,In_535);
nand U9 (N_9,In_1314,In_53);
and U10 (N_10,In_1189,In_1248);
or U11 (N_11,In_1070,In_543);
or U12 (N_12,In_745,In_103);
or U13 (N_13,In_856,In_628);
or U14 (N_14,In_525,In_587);
xor U15 (N_15,In_1055,In_1482);
or U16 (N_16,In_879,In_1207);
or U17 (N_17,In_654,In_424);
nand U18 (N_18,In_1114,In_1083);
or U19 (N_19,In_751,In_970);
xor U20 (N_20,In_271,In_871);
nand U21 (N_21,In_393,In_573);
or U22 (N_22,In_564,In_144);
or U23 (N_23,In_118,In_1021);
nand U24 (N_24,In_1119,In_312);
nor U25 (N_25,In_1341,In_209);
nor U26 (N_26,In_348,In_148);
or U27 (N_27,In_1067,In_1089);
nand U28 (N_28,In_650,In_1249);
or U29 (N_29,In_522,In_1244);
or U30 (N_30,In_1209,In_1264);
nand U31 (N_31,In_826,In_12);
nand U32 (N_32,In_615,In_1356);
nor U33 (N_33,In_937,In_548);
xnor U34 (N_34,In_1198,In_1022);
nor U35 (N_35,In_537,In_991);
and U36 (N_36,In_74,In_1292);
or U37 (N_37,In_61,In_938);
xor U38 (N_38,In_1174,In_128);
xnor U39 (N_39,In_59,In_859);
or U40 (N_40,In_583,In_444);
or U41 (N_41,In_787,In_323);
nor U42 (N_42,In_1102,In_613);
nand U43 (N_43,In_767,In_11);
nor U44 (N_44,In_1284,In_143);
nor U45 (N_45,In_1117,In_136);
and U46 (N_46,In_299,In_1254);
and U47 (N_47,In_646,In_472);
or U48 (N_48,In_1487,In_105);
and U49 (N_49,In_1076,In_772);
or U50 (N_50,In_530,In_754);
nor U51 (N_51,In_1126,In_1006);
or U52 (N_52,In_477,In_675);
and U53 (N_53,In_1407,In_364);
nand U54 (N_54,In_138,In_1016);
and U55 (N_55,In_170,In_208);
xnor U56 (N_56,In_1060,In_630);
nor U57 (N_57,In_894,In_1192);
and U58 (N_58,In_391,In_1494);
or U59 (N_59,In_419,In_178);
nand U60 (N_60,In_332,In_979);
nand U61 (N_61,In_791,In_235);
and U62 (N_62,In_198,In_80);
or U63 (N_63,In_1395,In_1275);
nand U64 (N_64,In_1128,In_949);
nor U65 (N_65,In_577,In_867);
or U66 (N_66,In_1216,In_1047);
xnor U67 (N_67,In_1136,In_90);
and U68 (N_68,In_596,In_129);
or U69 (N_69,In_1251,In_72);
xnor U70 (N_70,In_1200,In_1228);
and U71 (N_71,In_1353,In_1236);
or U72 (N_72,In_1245,In_1059);
xnor U73 (N_73,In_1010,In_950);
and U74 (N_74,In_724,In_329);
xnor U75 (N_75,In_1288,In_1419);
nor U76 (N_76,In_956,In_232);
nand U77 (N_77,In_32,In_292);
or U78 (N_78,In_24,In_172);
or U79 (N_79,In_658,In_540);
nor U80 (N_80,In_1274,In_351);
xnor U81 (N_81,In_199,In_995);
xnor U82 (N_82,In_353,In_397);
and U83 (N_83,In_431,In_343);
nand U84 (N_84,In_226,In_490);
and U85 (N_85,In_1421,In_1417);
or U86 (N_86,In_983,In_774);
nor U87 (N_87,In_114,In_1342);
or U88 (N_88,In_1387,In_340);
xnor U89 (N_89,In_660,In_741);
or U90 (N_90,In_1149,In_810);
and U91 (N_91,In_1298,In_51);
xor U92 (N_92,In_926,In_1365);
or U93 (N_93,In_1110,In_420);
nand U94 (N_94,In_498,In_940);
nor U95 (N_95,In_177,In_268);
nor U96 (N_96,In_714,In_972);
or U97 (N_97,In_84,In_966);
nor U98 (N_98,In_812,In_180);
or U99 (N_99,In_1397,In_87);
xor U100 (N_100,In_273,In_743);
xnor U101 (N_101,In_1170,In_1265);
and U102 (N_102,In_293,In_819);
xnor U103 (N_103,In_527,In_30);
xor U104 (N_104,In_324,In_201);
or U105 (N_105,In_418,In_415);
or U106 (N_106,In_1478,In_524);
nor U107 (N_107,In_895,In_1481);
nand U108 (N_108,In_451,In_1178);
or U109 (N_109,In_285,In_492);
and U110 (N_110,In_697,In_33);
xor U111 (N_111,In_6,In_1252);
or U112 (N_112,In_716,In_375);
nor U113 (N_113,In_1235,In_249);
or U114 (N_114,In_975,In_484);
nor U115 (N_115,In_473,In_592);
nand U116 (N_116,In_486,In_1327);
or U117 (N_117,In_1375,In_779);
nand U118 (N_118,In_1168,In_1144);
nor U119 (N_119,In_1466,In_528);
nand U120 (N_120,In_464,In_1279);
xnor U121 (N_121,In_456,In_1476);
and U122 (N_122,In_1111,In_1156);
xor U123 (N_123,In_997,In_511);
xnor U124 (N_124,In_920,In_1187);
nand U125 (N_125,In_34,In_1374);
xor U126 (N_126,In_770,In_644);
and U127 (N_127,In_680,In_984);
and U128 (N_128,In_1237,In_831);
nand U129 (N_129,In_744,In_1309);
nor U130 (N_130,In_1243,In_1217);
xor U131 (N_131,In_1088,In_1191);
xnor U132 (N_132,In_1295,In_777);
nand U133 (N_133,In_885,In_1062);
or U134 (N_134,In_1372,In_536);
and U135 (N_135,In_883,In_514);
nor U136 (N_136,In_225,In_556);
or U137 (N_137,In_1322,In_572);
xor U138 (N_138,In_1204,In_679);
xor U139 (N_139,In_1091,In_927);
or U140 (N_140,In_862,In_1496);
or U141 (N_141,In_775,In_400);
nand U142 (N_142,In_196,In_319);
and U143 (N_143,In_252,In_1253);
nor U144 (N_144,In_989,In_880);
nor U145 (N_145,In_1474,In_1137);
nand U146 (N_146,In_1151,In_439);
nand U147 (N_147,In_1409,In_645);
nand U148 (N_148,In_303,In_39);
or U149 (N_149,In_1472,In_1316);
nor U150 (N_150,In_460,In_491);
or U151 (N_151,In_179,In_229);
nor U152 (N_152,In_125,In_78);
xor U153 (N_153,In_414,In_1097);
nand U154 (N_154,In_955,In_900);
nor U155 (N_155,In_270,In_427);
and U156 (N_156,In_374,In_843);
and U157 (N_157,In_1090,In_605);
or U158 (N_158,In_974,In_474);
nor U159 (N_159,In_260,In_10);
and U160 (N_160,In_147,In_488);
xor U161 (N_161,In_304,In_476);
nor U162 (N_162,In_1073,In_803);
nand U163 (N_163,In_107,In_619);
xor U164 (N_164,In_447,In_661);
or U165 (N_165,In_1130,In_590);
xnor U166 (N_166,In_865,In_496);
nand U167 (N_167,In_1049,In_575);
nand U168 (N_168,In_1438,In_98);
or U169 (N_169,In_953,In_68);
nor U170 (N_170,In_578,In_585);
or U171 (N_171,In_1003,In_263);
nand U172 (N_172,In_603,In_933);
and U173 (N_173,In_321,In_501);
xor U174 (N_174,In_295,In_1210);
xnor U175 (N_175,In_916,In_789);
nor U176 (N_176,In_1369,In_1159);
nand U177 (N_177,In_727,In_482);
xnor U178 (N_178,In_403,In_63);
or U179 (N_179,In_794,In_570);
and U180 (N_180,In_708,In_64);
or U181 (N_181,In_1414,In_206);
or U182 (N_182,In_834,In_652);
nor U183 (N_183,In_684,In_1183);
xor U184 (N_184,In_217,In_811);
and U185 (N_185,In_1220,In_1424);
or U186 (N_186,In_1093,In_946);
and U187 (N_187,In_919,In_386);
or U188 (N_188,In_942,In_720);
or U189 (N_189,In_888,In_1164);
nor U190 (N_190,In_1429,In_222);
and U191 (N_191,In_185,In_1082);
nand U192 (N_192,In_366,In_835);
and U193 (N_193,In_686,In_598);
and U194 (N_194,In_426,In_1357);
and U195 (N_195,In_1402,In_541);
nand U196 (N_196,In_574,In_157);
nand U197 (N_197,In_1394,In_766);
nor U198 (N_198,In_623,In_240);
or U199 (N_199,In_274,In_696);
xor U200 (N_200,In_1013,In_493);
nor U201 (N_201,In_553,In_459);
and U202 (N_202,In_126,In_1305);
nor U203 (N_203,In_124,In_1413);
nor U204 (N_204,In_765,In_480);
or U205 (N_205,In_1400,In_504);
and U206 (N_206,In_1473,In_134);
or U207 (N_207,In_1162,In_71);
nand U208 (N_208,In_49,In_993);
nor U209 (N_209,In_694,In_930);
and U210 (N_210,In_89,In_308);
nor U211 (N_211,In_1468,In_731);
or U212 (N_212,In_1108,In_1377);
or U213 (N_213,In_17,In_1354);
and U214 (N_214,In_117,In_1329);
and U215 (N_215,In_761,In_1447);
or U216 (N_216,In_1085,In_212);
xor U217 (N_217,In_120,In_318);
and U218 (N_218,In_494,In_711);
or U219 (N_219,In_1036,In_814);
nand U220 (N_220,In_821,In_958);
nand U221 (N_221,In_756,In_101);
nor U222 (N_222,In_1452,In_326);
xor U223 (N_223,In_1226,In_820);
and U224 (N_224,In_816,In_1283);
nand U225 (N_225,In_19,In_505);
nor U226 (N_226,In_901,In_358);
nand U227 (N_227,In_1432,In_1194);
xnor U228 (N_228,In_625,In_710);
nor U229 (N_229,In_740,In_1074);
and U230 (N_230,In_647,In_663);
and U231 (N_231,In_191,In_643);
xor U232 (N_232,In_705,In_726);
xor U233 (N_233,In_1197,In_194);
and U234 (N_234,In_837,In_762);
xnor U235 (N_235,In_428,In_47);
and U236 (N_236,In_357,In_1320);
and U237 (N_237,In_907,In_1332);
xnor U238 (N_238,In_372,In_119);
and U239 (N_239,In_1359,In_932);
xor U240 (N_240,In_665,In_893);
and U241 (N_241,In_432,In_500);
nor U242 (N_242,In_91,In_1449);
and U243 (N_243,In_192,In_1124);
xnor U244 (N_244,In_193,In_320);
nor U245 (N_245,In_813,In_1142);
nor U246 (N_246,In_610,In_227);
nand U247 (N_247,In_1107,In_988);
xnor U248 (N_248,In_655,In_36);
nor U249 (N_249,In_566,In_759);
or U250 (N_250,In_1173,In_873);
xor U251 (N_251,In_1034,In_195);
nand U252 (N_252,In_636,In_54);
xnor U253 (N_253,In_1287,In_1495);
xnor U254 (N_254,In_1380,In_747);
nor U255 (N_255,In_467,In_702);
xnor U256 (N_256,In_450,In_1340);
or U257 (N_257,In_214,In_839);
nand U258 (N_258,In_887,In_700);
xnor U259 (N_259,In_1058,In_341);
xnor U260 (N_260,In_1460,In_335);
xnor U261 (N_261,In_1238,In_1441);
nor U262 (N_262,In_1229,In_586);
nand U263 (N_263,In_855,In_255);
nor U264 (N_264,In_844,In_796);
and U265 (N_265,In_969,In_1161);
xor U266 (N_266,In_1433,In_306);
and U267 (N_267,In_184,In_874);
nor U268 (N_268,In_634,In_1263);
xor U269 (N_269,In_479,In_653);
or U270 (N_270,In_187,In_689);
and U271 (N_271,In_1368,In_186);
xor U272 (N_272,In_13,In_631);
nand U273 (N_273,In_555,In_682);
xor U274 (N_274,In_985,In_437);
nor U275 (N_275,In_1002,In_96);
or U276 (N_276,In_1373,In_0);
xor U277 (N_277,In_521,In_1045);
xnor U278 (N_278,In_1202,In_1445);
nand U279 (N_279,In_111,In_836);
nor U280 (N_280,In_1464,In_388);
nor U281 (N_281,In_1299,In_1146);
or U282 (N_282,In_1041,In_936);
nor U283 (N_283,In_149,In_238);
xnor U284 (N_284,In_830,In_223);
nand U285 (N_285,In_1218,In_1463);
or U286 (N_286,In_863,In_1440);
nor U287 (N_287,In_1431,In_878);
nor U288 (N_288,In_1133,In_558);
or U289 (N_289,In_1348,In_1430);
xnor U290 (N_290,In_159,In_167);
and U291 (N_291,In_452,In_538);
xnor U292 (N_292,In_569,In_175);
or U293 (N_293,In_924,In_1050);
nor U294 (N_294,In_822,In_687);
xor U295 (N_295,In_1427,In_651);
nor U296 (N_296,In_905,In_325);
or U297 (N_297,In_1317,In_1081);
nand U298 (N_298,In_516,In_1150);
or U299 (N_299,In_1345,In_1379);
or U300 (N_300,In_1385,In_337);
xnor U301 (N_301,In_875,In_565);
and U302 (N_302,In_438,In_365);
nor U303 (N_303,In_549,In_445);
xnor U304 (N_304,In_1393,In_846);
nand U305 (N_305,In_487,In_551);
xor U306 (N_306,In_183,In_1223);
and U307 (N_307,In_383,In_417);
and U308 (N_308,In_1297,In_1469);
nor U309 (N_309,In_841,In_469);
nor U310 (N_310,In_899,In_1423);
xor U311 (N_311,In_632,In_1281);
nor U312 (N_312,In_35,In_1257);
or U313 (N_313,In_877,In_600);
and U314 (N_314,In_559,In_161);
or U315 (N_315,In_440,In_1459);
nand U316 (N_316,In_849,In_639);
or U317 (N_317,In_50,In_331);
nor U318 (N_318,In_345,In_1153);
and U319 (N_319,In_1296,In_829);
xor U320 (N_320,In_1484,In_1328);
nor U321 (N_321,In_406,In_664);
and U322 (N_322,In_1205,In_1160);
or U323 (N_323,In_579,In_57);
xnor U324 (N_324,In_404,In_734);
xnor U325 (N_325,In_845,In_1470);
nand U326 (N_326,In_709,In_1405);
xnor U327 (N_327,In_378,In_1408);
and U328 (N_328,In_352,In_1378);
nor U329 (N_329,In_234,In_890);
nand U330 (N_330,In_595,In_264);
nand U331 (N_331,In_1234,In_1096);
or U332 (N_332,In_1017,In_602);
xor U333 (N_333,In_242,In_1009);
nand U334 (N_334,In_676,In_41);
xnor U335 (N_335,In_1129,In_563);
nor U336 (N_336,In_1222,In_1259);
nand U337 (N_337,In_1271,In_823);
xor U338 (N_338,In_801,In_67);
or U339 (N_339,In_77,In_994);
and U340 (N_340,In_739,In_1280);
or U341 (N_341,In_1318,In_470);
and U342 (N_342,In_718,In_95);
nor U343 (N_343,In_560,In_28);
or U344 (N_344,In_221,In_162);
or U345 (N_345,In_635,In_468);
and U346 (N_346,In_478,In_23);
xnor U347 (N_347,In_1208,In_656);
and U348 (N_348,In_373,In_818);
or U349 (N_349,In_735,In_1426);
and U350 (N_350,In_1388,In_156);
nor U351 (N_351,In_550,In_1391);
nor U352 (N_352,In_1044,In_908);
xor U353 (N_353,In_56,In_638);
xnor U354 (N_354,In_1276,In_1132);
or U355 (N_355,In_1258,In_1330);
or U356 (N_356,In_9,In_568);
or U357 (N_357,In_886,In_588);
and U358 (N_358,In_1437,In_922);
or U359 (N_359,In_611,In_852);
xnor U360 (N_360,In_359,In_305);
nor U361 (N_361,In_29,In_864);
nand U362 (N_362,In_690,In_1072);
nor U363 (N_363,In_1489,In_239);
nand U364 (N_364,In_703,In_442);
xnor U365 (N_365,In_941,In_562);
or U366 (N_366,In_1000,In_1435);
xor U367 (N_367,In_65,In_339);
nor U368 (N_368,In_1381,In_346);
or U369 (N_369,In_116,In_1056);
nand U370 (N_370,In_998,In_783);
or U371 (N_371,In_20,In_286);
nand U372 (N_372,In_982,In_1171);
xnor U373 (N_373,In_173,In_868);
nor U374 (N_374,In_301,In_317);
xor U375 (N_375,In_617,In_1319);
and U376 (N_376,In_462,In_706);
and U377 (N_377,In_1214,In_869);
and U378 (N_378,In_992,In_557);
and U379 (N_379,In_1350,In_166);
nand U380 (N_380,In_1383,In_1172);
or U381 (N_381,In_1268,In_792);
nand U382 (N_382,In_1053,In_1446);
xnor U383 (N_383,In_205,In_842);
and U384 (N_384,In_499,In_928);
xor U385 (N_385,In_788,In_1262);
or U386 (N_386,In_968,In_145);
nor U387 (N_387,In_659,In_1454);
xnor U388 (N_388,In_963,In_188);
xnor U389 (N_389,In_354,In_546);
xor U390 (N_390,In_723,In_1344);
nor U391 (N_391,In_405,In_1182);
or U392 (N_392,In_361,In_413);
and U393 (N_393,In_399,In_959);
xnor U394 (N_394,In_1071,In_510);
nand U395 (N_395,In_1231,In_1075);
nand U396 (N_396,In_925,In_902);
nor U397 (N_397,In_817,In_591);
nand U398 (N_398,In_858,In_376);
xor U399 (N_399,In_580,In_1411);
nand U400 (N_400,In_1486,In_475);
nor U401 (N_401,In_93,In_798);
or U402 (N_402,In_931,In_45);
nor U403 (N_403,In_151,In_1416);
nor U404 (N_404,In_624,In_1054);
xor U405 (N_405,In_939,In_552);
and U406 (N_406,In_211,In_246);
nand U407 (N_407,In_506,In_1131);
and U408 (N_408,In_1079,In_333);
nand U409 (N_409,In_601,In_531);
nand U410 (N_410,In_377,In_730);
or U411 (N_411,In_311,In_254);
xor U412 (N_412,In_1382,In_86);
nand U413 (N_413,In_1007,In_692);
xor U414 (N_414,In_69,In_633);
or U415 (N_415,In_100,In_233);
and U416 (N_416,In_1061,In_999);
nor U417 (N_417,In_778,In_1392);
nor U418 (N_418,In_1358,In_1030);
nor U419 (N_419,In_371,In_497);
xor U420 (N_420,In_1488,In_1029);
nor U421 (N_421,In_1015,In_181);
or U422 (N_422,In_547,In_218);
and U423 (N_423,In_1014,In_457);
and U424 (N_424,In_1256,In_1232);
nor U425 (N_425,In_515,In_929);
or U426 (N_426,In_307,In_1415);
nor U427 (N_427,In_122,In_441);
nand U428 (N_428,In_1106,In_197);
or U429 (N_429,In_349,In_1042);
nand U430 (N_430,In_1152,In_1065);
and U431 (N_431,In_1410,In_790);
nor U432 (N_432,In_1035,In_909);
nand U433 (N_433,In_889,In_449);
xor U434 (N_434,In_1193,In_973);
and U435 (N_435,In_313,In_1491);
nor U436 (N_436,In_674,In_620);
nand U437 (N_437,In_1037,In_502);
xor U438 (N_438,In_146,In_1242);
and U439 (N_439,In_315,In_121);
and U440 (N_440,In_1046,In_27);
nor U441 (N_441,In_278,In_1179);
xor U442 (N_442,In_840,In_1139);
and U443 (N_443,In_594,In_668);
nor U444 (N_444,In_3,In_42);
nor U445 (N_445,In_614,In_597);
and U446 (N_446,In_1304,In_1403);
xor U447 (N_447,In_411,In_485);
and U448 (N_448,In_135,In_1290);
or U449 (N_449,In_81,In_1462);
nand U450 (N_450,In_1457,In_1498);
nor U451 (N_451,In_106,In_1138);
xor U452 (N_452,In_1312,In_1005);
nor U453 (N_453,In_1412,In_1346);
and U454 (N_454,In_267,In_768);
or U455 (N_455,In_1499,In_113);
xor U456 (N_456,In_385,In_1118);
and U457 (N_457,In_109,In_673);
or U458 (N_458,In_275,In_280);
or U459 (N_459,In_666,In_137);
xor U460 (N_460,In_1233,In_422);
nor U461 (N_461,In_1227,In_1155);
nor U462 (N_462,In_1326,In_102);
or U463 (N_463,In_806,In_471);
nor U464 (N_464,In_465,In_1051);
or U465 (N_465,In_746,In_769);
nor U466 (N_466,In_934,In_1370);
xnor U467 (N_467,In_75,In_629);
xor U468 (N_468,In_362,In_827);
or U469 (N_469,In_1289,In_104);
or U470 (N_470,In_257,In_1337);
or U471 (N_471,In_21,In_1143);
xnor U472 (N_472,In_31,In_721);
nor U473 (N_473,In_758,In_785);
nor U474 (N_474,In_1147,In_423);
and U475 (N_475,In_1084,In_1175);
nor U476 (N_476,In_848,In_1336);
or U477 (N_477,In_996,In_1425);
and U478 (N_478,In_520,In_350);
or U479 (N_479,In_707,In_1286);
and U480 (N_480,In_284,In_898);
nand U481 (N_481,In_1371,In_621);
xnor U482 (N_482,In_797,In_108);
nor U483 (N_483,In_1184,In_965);
and U484 (N_484,In_854,In_860);
nor U485 (N_485,In_1255,In_576);
or U486 (N_486,In_897,In_512);
xor U487 (N_487,In_626,In_434);
or U488 (N_488,In_1122,In_97);
or U489 (N_489,In_369,In_685);
nand U490 (N_490,In_748,In_435);
and U491 (N_491,In_960,In_545);
nor U492 (N_492,In_1077,In_70);
and U493 (N_493,In_396,In_912);
nor U494 (N_494,In_251,In_322);
and U495 (N_495,In_713,In_1479);
nand U496 (N_496,In_141,In_18);
or U497 (N_497,In_1165,In_1188);
xor U498 (N_498,In_833,In_1109);
nand U499 (N_499,In_1080,In_328);
xor U500 (N_500,In_446,In_1201);
nand U501 (N_501,In_1450,In_824);
nor U502 (N_502,In_776,In_123);
nand U503 (N_503,In_809,In_957);
or U504 (N_504,In_1347,In_1105);
nor U505 (N_505,In_825,In_1361);
nand U506 (N_506,In_189,In_224);
xor U507 (N_507,In_294,In_1390);
xnor U508 (N_508,In_410,In_207);
nand U509 (N_509,In_1461,In_330);
nand U510 (N_510,In_951,In_1483);
nand U511 (N_511,In_944,In_245);
or U512 (N_512,In_142,In_1480);
nor U513 (N_513,In_1351,In_38);
xor U514 (N_514,In_94,In_1451);
xnor U515 (N_515,In_1303,In_533);
and U516 (N_516,In_1324,In_1169);
xnor U517 (N_517,In_1367,In_230);
or U518 (N_518,In_1066,In_1458);
nand U519 (N_519,In_483,In_1266);
nand U520 (N_520,In_971,In_1196);
or U521 (N_521,In_1331,In_561);
and U522 (N_522,In_455,In_99);
or U523 (N_523,In_612,In_1475);
nor U524 (N_524,In_733,In_1052);
xor U525 (N_525,In_298,In_1241);
nand U526 (N_526,In_805,In_1335);
or U527 (N_527,In_1334,In_279);
and U528 (N_528,In_1493,In_755);
nand U529 (N_529,In_642,In_542);
nor U530 (N_530,In_1,In_892);
nand U531 (N_531,In_523,In_964);
or U532 (N_532,In_1167,In_737);
xnor U533 (N_533,In_911,In_1339);
xnor U534 (N_534,In_683,In_1315);
nor U535 (N_535,In_967,In_637);
xor U536 (N_536,In_976,In_37);
nor U537 (N_537,In_616,In_8);
nor U538 (N_538,In_1270,In_204);
nand U539 (N_539,In_904,In_1278);
and U540 (N_540,In_1057,In_712);
or U541 (N_541,In_913,In_1158);
or U542 (N_542,In_750,In_1338);
nand U543 (N_543,In_981,In_421);
or U544 (N_544,In_784,In_1140);
and U545 (N_545,In_25,In_342);
or U546 (N_546,In_231,In_589);
nor U547 (N_547,In_1355,In_398);
xnor U548 (N_548,In_529,In_237);
xnor U549 (N_549,In_677,In_1120);
xor U550 (N_550,In_1376,In_454);
and U551 (N_551,In_236,In_1293);
and U552 (N_552,In_152,In_1272);
xor U553 (N_553,In_200,In_729);
and U554 (N_554,In_1112,In_903);
and U555 (N_555,In_980,In_881);
nor U556 (N_556,In_216,In_1099);
xnor U557 (N_557,In_1420,In_276);
nand U558 (N_558,In_608,In_606);
nand U559 (N_559,In_407,In_52);
xnor U560 (N_560,In_202,In_1211);
and U561 (N_561,In_1343,In_265);
nor U562 (N_562,In_1068,In_978);
xor U563 (N_563,In_567,In_336);
nor U564 (N_564,In_1246,In_593);
xor U565 (N_565,In_882,In_519);
nand U566 (N_566,In_1043,In_281);
xor U567 (N_567,In_158,In_923);
nand U568 (N_568,In_327,In_1026);
and U569 (N_569,In_808,In_914);
xnor U570 (N_570,In_150,In_872);
and U571 (N_571,In_62,In_243);
nand U572 (N_572,In_262,In_1300);
nand U573 (N_573,In_168,In_15);
xnor U574 (N_574,In_392,In_219);
nor U575 (N_575,In_802,In_627);
and U576 (N_576,In_344,In_990);
xor U577 (N_577,In_253,In_356);
nand U578 (N_578,In_1157,In_133);
or U579 (N_579,In_1185,In_1384);
and U580 (N_580,In_334,In_55);
xnor U581 (N_581,In_1177,In_847);
or U582 (N_582,In_213,In_46);
nor U583 (N_583,In_1492,In_1190);
and U584 (N_584,In_1100,In_948);
and U585 (N_585,In_760,In_1247);
nand U586 (N_586,In_1301,In_917);
nor U587 (N_587,In_640,In_382);
xor U588 (N_588,In_935,In_773);
nand U589 (N_589,In_461,In_1443);
or U590 (N_590,In_503,In_604);
nand U591 (N_591,In_657,In_1148);
or U592 (N_592,In_722,In_266);
nor U593 (N_593,In_368,In_429);
or U594 (N_594,In_513,In_691);
and U595 (N_595,In_1069,In_1311);
nand U596 (N_596,In_669,In_408);
nor U597 (N_597,In_16,In_648);
nand U598 (N_598,In_1490,In_1028);
and U599 (N_599,In_1485,In_1455);
and U600 (N_600,In_699,In_943);
nor U601 (N_601,In_1453,In_76);
or U602 (N_602,In_370,In_1428);
or U603 (N_603,In_1442,In_5);
and U604 (N_604,In_670,In_85);
nand U605 (N_605,In_1180,In_1439);
nor U606 (N_606,In_728,In_508);
nand U607 (N_607,In_244,In_310);
xnor U608 (N_608,In_618,In_509);
nor U609 (N_609,In_582,In_517);
xnor U610 (N_610,In_402,In_1040);
or U611 (N_611,In_387,In_495);
or U612 (N_612,In_667,In_1224);
xnor U613 (N_613,In_1023,In_58);
nand U614 (N_614,In_1399,In_876);
or U615 (N_615,In_609,In_977);
and U616 (N_616,In_554,In_804);
nor U617 (N_617,In_367,In_1321);
or U618 (N_618,In_1020,In_247);
xnor U619 (N_619,In_607,In_584);
xnor U620 (N_620,In_40,In_1098);
and U621 (N_621,In_79,In_1033);
xor U622 (N_622,In_1116,In_954);
nor U623 (N_623,In_662,In_165);
or U624 (N_624,In_297,In_381);
or U625 (N_625,In_302,In_1025);
nor U626 (N_626,In_1141,In_210);
xor U627 (N_627,In_127,In_409);
nor U628 (N_628,In_448,In_678);
nand U629 (N_629,In_1444,In_1113);
and U630 (N_630,In_725,In_891);
nand U631 (N_631,In_83,In_1195);
or U632 (N_632,In_1134,In_782);
or U633 (N_633,In_73,In_338);
xor U634 (N_634,In_1024,In_1135);
or U635 (N_635,In_258,In_715);
or U636 (N_636,In_532,In_163);
or U637 (N_637,In_1497,In_681);
or U638 (N_638,In_1230,In_300);
xnor U639 (N_639,In_132,In_1398);
xor U640 (N_640,In_896,In_1095);
xnor U641 (N_641,In_1219,In_1163);
nor U642 (N_642,In_1277,In_793);
nor U643 (N_643,In_1471,In_1012);
and U644 (N_644,In_1250,In_688);
nand U645 (N_645,In_154,In_190);
nor U646 (N_646,In_704,In_463);
nand U647 (N_647,In_795,In_363);
nand U648 (N_648,In_394,In_433);
nor U649 (N_649,In_1467,In_1396);
xor U650 (N_650,In_228,In_1011);
nand U651 (N_651,In_1308,In_701);
nor U652 (N_652,In_82,In_164);
nand U653 (N_653,In_2,In_1213);
nor U654 (N_654,In_732,In_918);
or U655 (N_655,In_261,In_160);
nor U656 (N_656,In_526,In_719);
and U657 (N_657,In_14,In_752);
nor U658 (N_658,In_1282,In_1260);
xor U659 (N_659,In_1078,In_671);
nand U660 (N_660,In_182,In_220);
and U661 (N_661,In_518,In_1103);
nor U662 (N_662,In_1404,In_1306);
nand U663 (N_663,In_1166,In_379);
and U664 (N_664,In_1032,In_1181);
nand U665 (N_665,In_910,In_155);
nor U666 (N_666,In_915,In_853);
nand U667 (N_667,In_48,In_838);
nor U668 (N_668,In_131,In_1092);
nand U669 (N_669,In_466,In_832);
or U670 (N_670,In_1401,In_1406);
and U671 (N_671,In_693,In_1389);
xnor U672 (N_672,In_1038,In_347);
or U673 (N_673,In_1203,In_241);
and U674 (N_674,In_291,In_1176);
or U675 (N_675,In_1261,In_66);
or U676 (N_676,In_389,In_786);
and U677 (N_677,In_453,In_1086);
xor U678 (N_678,In_1212,In_1206);
xnor U679 (N_679,In_1307,In_1448);
nor U680 (N_680,In_169,In_1104);
or U681 (N_681,In_599,In_1115);
nand U682 (N_682,In_1386,In_1267);
xnor U683 (N_683,In_945,In_112);
nand U684 (N_684,In_269,In_507);
and U685 (N_685,In_742,In_1121);
nand U686 (N_686,In_952,In_277);
nand U687 (N_687,In_26,In_753);
nor U688 (N_688,In_649,In_1333);
or U689 (N_689,In_174,In_250);
nor U690 (N_690,In_780,In_256);
or U691 (N_691,In_1199,In_355);
and U692 (N_692,In_1127,In_489);
nand U693 (N_693,In_1349,In_781);
xor U694 (N_694,In_695,In_749);
nor U695 (N_695,In_861,In_1027);
nor U696 (N_696,In_416,In_248);
xor U697 (N_697,In_1001,In_1048);
or U698 (N_698,In_272,In_130);
and U699 (N_699,In_581,In_1008);
or U700 (N_700,In_1018,In_259);
xnor U701 (N_701,In_139,In_986);
nor U702 (N_702,In_1186,In_88);
nor U703 (N_703,In_1154,In_1145);
xnor U704 (N_704,In_757,In_1123);
nand U705 (N_705,In_866,In_1364);
or U706 (N_706,In_140,In_384);
nand U707 (N_707,In_1434,In_962);
xor U708 (N_708,In_800,In_458);
nand U709 (N_709,In_1291,In_1221);
xor U710 (N_710,In_799,In_906);
or U711 (N_711,In_115,In_110);
and U712 (N_712,In_316,In_987);
xor U713 (N_713,In_1477,In_443);
and U714 (N_714,In_1366,In_309);
nand U715 (N_715,In_1360,In_1363);
and U716 (N_716,In_395,In_1269);
xnor U717 (N_717,In_1352,In_176);
and U718 (N_718,In_203,In_1094);
nand U719 (N_719,In_1125,In_296);
xnor U720 (N_720,In_171,In_44);
or U721 (N_721,In_287,In_884);
or U722 (N_722,In_1313,In_390);
nor U723 (N_723,In_1273,In_1240);
nand U724 (N_724,In_828,In_289);
xor U725 (N_725,In_401,In_290);
or U726 (N_726,In_850,In_22);
and U727 (N_727,In_1422,In_764);
or U728 (N_728,In_215,In_288);
nand U729 (N_729,In_571,In_1031);
nand U730 (N_730,In_7,In_60);
xnor U731 (N_731,In_314,In_1323);
xnor U732 (N_732,In_622,In_763);
and U733 (N_733,In_360,In_1064);
and U734 (N_734,In_1004,In_961);
nand U735 (N_735,In_4,In_92);
nand U736 (N_736,In_283,In_1063);
and U737 (N_737,In_1101,In_43);
nor U738 (N_738,In_717,In_1294);
and U739 (N_739,In_380,In_1039);
or U740 (N_740,In_1239,In_771);
nand U741 (N_741,In_1087,In_412);
nand U742 (N_742,In_1456,In_1325);
nand U743 (N_743,In_539,In_1302);
nand U744 (N_744,In_947,In_738);
nand U745 (N_745,In_641,In_1362);
and U746 (N_746,In_1019,In_1285);
nand U747 (N_747,In_534,In_1225);
nor U748 (N_748,In_425,In_672);
nand U749 (N_749,In_698,In_851);
nor U750 (N_750,In_23,In_530);
and U751 (N_751,In_335,In_732);
nand U752 (N_752,In_952,In_1199);
or U753 (N_753,In_311,In_1186);
xnor U754 (N_754,In_1369,In_188);
xor U755 (N_755,In_730,In_1488);
xnor U756 (N_756,In_1078,In_18);
nand U757 (N_757,In_307,In_468);
and U758 (N_758,In_1304,In_193);
nor U759 (N_759,In_880,In_240);
nor U760 (N_760,In_194,In_734);
and U761 (N_761,In_1190,In_1166);
or U762 (N_762,In_1259,In_451);
nand U763 (N_763,In_1139,In_666);
nor U764 (N_764,In_1371,In_776);
and U765 (N_765,In_186,In_398);
nand U766 (N_766,In_1283,In_1352);
and U767 (N_767,In_461,In_1467);
and U768 (N_768,In_1316,In_296);
nor U769 (N_769,In_218,In_951);
xor U770 (N_770,In_566,In_684);
and U771 (N_771,In_1352,In_972);
and U772 (N_772,In_281,In_782);
nand U773 (N_773,In_858,In_228);
and U774 (N_774,In_109,In_1123);
xnor U775 (N_775,In_804,In_543);
and U776 (N_776,In_145,In_922);
xor U777 (N_777,In_196,In_35);
nor U778 (N_778,In_1370,In_346);
xor U779 (N_779,In_1235,In_143);
nor U780 (N_780,In_812,In_240);
and U781 (N_781,In_938,In_1287);
xor U782 (N_782,In_590,In_481);
xnor U783 (N_783,In_781,In_169);
and U784 (N_784,In_853,In_711);
or U785 (N_785,In_728,In_32);
or U786 (N_786,In_394,In_1173);
or U787 (N_787,In_1338,In_1195);
nor U788 (N_788,In_299,In_1440);
or U789 (N_789,In_794,In_503);
and U790 (N_790,In_593,In_366);
xnor U791 (N_791,In_929,In_356);
nor U792 (N_792,In_698,In_1125);
xnor U793 (N_793,In_997,In_959);
or U794 (N_794,In_546,In_1337);
and U795 (N_795,In_1010,In_1182);
nand U796 (N_796,In_1258,In_217);
nor U797 (N_797,In_625,In_1339);
or U798 (N_798,In_391,In_1136);
nor U799 (N_799,In_605,In_1002);
xor U800 (N_800,In_1450,In_1044);
nor U801 (N_801,In_748,In_721);
nor U802 (N_802,In_805,In_936);
nand U803 (N_803,In_496,In_51);
or U804 (N_804,In_409,In_1427);
or U805 (N_805,In_894,In_96);
nand U806 (N_806,In_1271,In_700);
nand U807 (N_807,In_823,In_177);
xnor U808 (N_808,In_1147,In_1016);
nand U809 (N_809,In_376,In_766);
nor U810 (N_810,In_953,In_1223);
nand U811 (N_811,In_795,In_17);
xor U812 (N_812,In_1025,In_532);
nand U813 (N_813,In_814,In_565);
nor U814 (N_814,In_1392,In_1289);
nor U815 (N_815,In_1389,In_517);
or U816 (N_816,In_108,In_955);
and U817 (N_817,In_73,In_215);
nor U818 (N_818,In_387,In_705);
or U819 (N_819,In_140,In_1484);
or U820 (N_820,In_82,In_757);
nor U821 (N_821,In_1371,In_1498);
nand U822 (N_822,In_467,In_673);
nand U823 (N_823,In_996,In_994);
nor U824 (N_824,In_1398,In_837);
or U825 (N_825,In_620,In_884);
nand U826 (N_826,In_1321,In_404);
and U827 (N_827,In_1413,In_1146);
or U828 (N_828,In_13,In_1381);
nand U829 (N_829,In_289,In_313);
nand U830 (N_830,In_163,In_118);
nor U831 (N_831,In_969,In_190);
nor U832 (N_832,In_236,In_5);
nand U833 (N_833,In_1233,In_1333);
and U834 (N_834,In_1301,In_34);
and U835 (N_835,In_1246,In_878);
or U836 (N_836,In_1322,In_944);
nor U837 (N_837,In_322,In_961);
xnor U838 (N_838,In_984,In_112);
or U839 (N_839,In_110,In_354);
xnor U840 (N_840,In_303,In_621);
nand U841 (N_841,In_884,In_589);
xor U842 (N_842,In_883,In_461);
or U843 (N_843,In_866,In_863);
or U844 (N_844,In_295,In_1199);
or U845 (N_845,In_73,In_219);
nor U846 (N_846,In_686,In_1153);
nor U847 (N_847,In_989,In_1236);
nor U848 (N_848,In_1219,In_334);
xnor U849 (N_849,In_1492,In_2);
nand U850 (N_850,In_830,In_792);
xnor U851 (N_851,In_1249,In_1483);
nor U852 (N_852,In_186,In_732);
and U853 (N_853,In_609,In_1380);
nor U854 (N_854,In_710,In_592);
or U855 (N_855,In_472,In_150);
nand U856 (N_856,In_393,In_1107);
xor U857 (N_857,In_681,In_16);
or U858 (N_858,In_876,In_87);
or U859 (N_859,In_1144,In_711);
nor U860 (N_860,In_1283,In_922);
nor U861 (N_861,In_228,In_561);
or U862 (N_862,In_16,In_838);
and U863 (N_863,In_682,In_1104);
and U864 (N_864,In_811,In_242);
or U865 (N_865,In_490,In_870);
xor U866 (N_866,In_1194,In_1076);
and U867 (N_867,In_1151,In_924);
nand U868 (N_868,In_1417,In_1162);
or U869 (N_869,In_1345,In_562);
or U870 (N_870,In_402,In_80);
nor U871 (N_871,In_1180,In_1250);
nand U872 (N_872,In_603,In_1282);
nand U873 (N_873,In_1095,In_1154);
and U874 (N_874,In_113,In_622);
xnor U875 (N_875,In_1273,In_810);
xor U876 (N_876,In_1421,In_1353);
or U877 (N_877,In_409,In_1004);
xor U878 (N_878,In_906,In_143);
and U879 (N_879,In_191,In_649);
xnor U880 (N_880,In_1289,In_1073);
xor U881 (N_881,In_401,In_62);
and U882 (N_882,In_917,In_961);
nor U883 (N_883,In_1320,In_1451);
nand U884 (N_884,In_1401,In_640);
xor U885 (N_885,In_913,In_671);
xnor U886 (N_886,In_283,In_951);
or U887 (N_887,In_1432,In_823);
and U888 (N_888,In_463,In_483);
and U889 (N_889,In_852,In_993);
nor U890 (N_890,In_830,In_876);
nor U891 (N_891,In_263,In_595);
or U892 (N_892,In_68,In_1250);
nand U893 (N_893,In_1100,In_232);
or U894 (N_894,In_1268,In_955);
or U895 (N_895,In_1066,In_795);
and U896 (N_896,In_811,In_898);
and U897 (N_897,In_162,In_899);
nand U898 (N_898,In_926,In_677);
nor U899 (N_899,In_526,In_1280);
nand U900 (N_900,In_1491,In_1109);
xnor U901 (N_901,In_452,In_294);
xnor U902 (N_902,In_1406,In_1493);
or U903 (N_903,In_1096,In_597);
or U904 (N_904,In_1323,In_980);
nor U905 (N_905,In_405,In_248);
nand U906 (N_906,In_1346,In_357);
nor U907 (N_907,In_1282,In_845);
xor U908 (N_908,In_1486,In_59);
nor U909 (N_909,In_501,In_1300);
nor U910 (N_910,In_1004,In_968);
xnor U911 (N_911,In_377,In_1407);
and U912 (N_912,In_800,In_1332);
and U913 (N_913,In_199,In_878);
or U914 (N_914,In_1443,In_286);
nand U915 (N_915,In_722,In_412);
xor U916 (N_916,In_1215,In_245);
nor U917 (N_917,In_602,In_167);
nand U918 (N_918,In_1373,In_268);
nand U919 (N_919,In_232,In_613);
nor U920 (N_920,In_1211,In_972);
and U921 (N_921,In_67,In_1136);
or U922 (N_922,In_1388,In_454);
and U923 (N_923,In_1397,In_781);
or U924 (N_924,In_610,In_262);
nor U925 (N_925,In_1132,In_237);
xnor U926 (N_926,In_1129,In_1416);
and U927 (N_927,In_353,In_1400);
and U928 (N_928,In_27,In_1067);
and U929 (N_929,In_756,In_223);
nand U930 (N_930,In_854,In_722);
xor U931 (N_931,In_1387,In_929);
and U932 (N_932,In_571,In_327);
or U933 (N_933,In_161,In_1422);
or U934 (N_934,In_214,In_1233);
and U935 (N_935,In_131,In_283);
xnor U936 (N_936,In_843,In_238);
and U937 (N_937,In_671,In_30);
nand U938 (N_938,In_291,In_1488);
xor U939 (N_939,In_1102,In_10);
nand U940 (N_940,In_706,In_333);
xnor U941 (N_941,In_697,In_1080);
or U942 (N_942,In_701,In_634);
and U943 (N_943,In_308,In_773);
xor U944 (N_944,In_1487,In_479);
or U945 (N_945,In_947,In_833);
xnor U946 (N_946,In_1288,In_627);
and U947 (N_947,In_693,In_462);
nand U948 (N_948,In_1067,In_438);
nor U949 (N_949,In_907,In_20);
xnor U950 (N_950,In_1350,In_770);
nand U951 (N_951,In_1047,In_162);
xnor U952 (N_952,In_414,In_1103);
and U953 (N_953,In_321,In_190);
and U954 (N_954,In_831,In_640);
or U955 (N_955,In_1177,In_904);
xnor U956 (N_956,In_417,In_1330);
nand U957 (N_957,In_317,In_607);
and U958 (N_958,In_29,In_595);
nor U959 (N_959,In_755,In_634);
or U960 (N_960,In_1265,In_177);
and U961 (N_961,In_514,In_329);
nor U962 (N_962,In_28,In_568);
nor U963 (N_963,In_433,In_796);
or U964 (N_964,In_622,In_227);
xnor U965 (N_965,In_914,In_696);
and U966 (N_966,In_356,In_411);
and U967 (N_967,In_1053,In_119);
xor U968 (N_968,In_69,In_51);
and U969 (N_969,In_249,In_682);
and U970 (N_970,In_1452,In_148);
or U971 (N_971,In_1450,In_1077);
nor U972 (N_972,In_105,In_422);
nor U973 (N_973,In_825,In_444);
xor U974 (N_974,In_1230,In_890);
xnor U975 (N_975,In_721,In_876);
or U976 (N_976,In_445,In_1136);
xor U977 (N_977,In_19,In_721);
or U978 (N_978,In_1228,In_1134);
nand U979 (N_979,In_590,In_810);
xor U980 (N_980,In_870,In_620);
nand U981 (N_981,In_1259,In_1291);
and U982 (N_982,In_307,In_56);
nor U983 (N_983,In_628,In_710);
xor U984 (N_984,In_918,In_257);
nand U985 (N_985,In_793,In_158);
or U986 (N_986,In_416,In_1474);
xor U987 (N_987,In_885,In_387);
or U988 (N_988,In_1334,In_688);
and U989 (N_989,In_1245,In_1460);
nor U990 (N_990,In_401,In_1190);
xnor U991 (N_991,In_348,In_1300);
nand U992 (N_992,In_629,In_1043);
nand U993 (N_993,In_406,In_987);
or U994 (N_994,In_980,In_695);
and U995 (N_995,In_1397,In_1377);
nand U996 (N_996,In_164,In_1278);
nand U997 (N_997,In_1432,In_628);
nand U998 (N_998,In_1213,In_226);
xor U999 (N_999,In_171,In_789);
and U1000 (N_1000,N_817,N_69);
or U1001 (N_1001,N_763,N_172);
nor U1002 (N_1002,N_436,N_542);
or U1003 (N_1003,N_327,N_324);
xor U1004 (N_1004,N_102,N_533);
nand U1005 (N_1005,N_475,N_952);
nor U1006 (N_1006,N_718,N_947);
or U1007 (N_1007,N_413,N_614);
nand U1008 (N_1008,N_841,N_145);
and U1009 (N_1009,N_309,N_688);
nand U1010 (N_1010,N_365,N_676);
nand U1011 (N_1011,N_690,N_976);
or U1012 (N_1012,N_217,N_496);
xor U1013 (N_1013,N_246,N_455);
nand U1014 (N_1014,N_122,N_687);
nor U1015 (N_1015,N_608,N_626);
nand U1016 (N_1016,N_564,N_294);
and U1017 (N_1017,N_173,N_190);
nor U1018 (N_1018,N_636,N_224);
nand U1019 (N_1019,N_158,N_319);
and U1020 (N_1020,N_485,N_747);
nor U1021 (N_1021,N_38,N_908);
nor U1022 (N_1022,N_81,N_663);
xnor U1023 (N_1023,N_573,N_208);
nand U1024 (N_1024,N_646,N_775);
nand U1025 (N_1025,N_195,N_20);
and U1026 (N_1026,N_417,N_376);
xor U1027 (N_1027,N_18,N_925);
or U1028 (N_1028,N_361,N_649);
and U1029 (N_1029,N_207,N_623);
or U1030 (N_1030,N_235,N_883);
or U1031 (N_1031,N_188,N_461);
or U1032 (N_1032,N_368,N_965);
and U1033 (N_1033,N_354,N_738);
nand U1034 (N_1034,N_279,N_333);
xnor U1035 (N_1035,N_423,N_613);
nor U1036 (N_1036,N_722,N_979);
and U1037 (N_1037,N_844,N_535);
or U1038 (N_1038,N_890,N_14);
or U1039 (N_1039,N_742,N_581);
or U1040 (N_1040,N_507,N_897);
and U1041 (N_1041,N_831,N_713);
or U1042 (N_1042,N_112,N_798);
or U1043 (N_1043,N_739,N_487);
nor U1044 (N_1044,N_26,N_702);
nand U1045 (N_1045,N_509,N_949);
nand U1046 (N_1046,N_956,N_910);
nand U1047 (N_1047,N_212,N_165);
xor U1048 (N_1048,N_761,N_539);
xor U1049 (N_1049,N_290,N_27);
nor U1050 (N_1050,N_149,N_306);
nand U1051 (N_1051,N_557,N_650);
or U1052 (N_1052,N_552,N_266);
xnor U1053 (N_1053,N_252,N_443);
or U1054 (N_1054,N_848,N_736);
xnor U1055 (N_1055,N_271,N_83);
nand U1056 (N_1056,N_437,N_971);
and U1057 (N_1057,N_37,N_359);
or U1058 (N_1058,N_384,N_167);
nand U1059 (N_1059,N_84,N_554);
or U1060 (N_1060,N_877,N_866);
nor U1061 (N_1061,N_625,N_972);
or U1062 (N_1062,N_641,N_981);
nor U1063 (N_1063,N_975,N_375);
xnor U1064 (N_1064,N_449,N_8);
nor U1065 (N_1065,N_293,N_757);
or U1066 (N_1066,N_227,N_703);
xor U1067 (N_1067,N_24,N_510);
xnor U1068 (N_1068,N_355,N_568);
or U1069 (N_1069,N_600,N_401);
nor U1070 (N_1070,N_743,N_729);
and U1071 (N_1071,N_469,N_79);
nor U1072 (N_1072,N_707,N_175);
and U1073 (N_1073,N_353,N_576);
xor U1074 (N_1074,N_901,N_503);
xor U1075 (N_1075,N_813,N_345);
or U1076 (N_1076,N_275,N_807);
nand U1077 (N_1077,N_322,N_456);
xor U1078 (N_1078,N_248,N_396);
nand U1079 (N_1079,N_445,N_860);
xor U1080 (N_1080,N_984,N_887);
xnor U1081 (N_1081,N_385,N_500);
and U1082 (N_1082,N_490,N_67);
nand U1083 (N_1083,N_155,N_301);
xnor U1084 (N_1084,N_618,N_42);
xnor U1085 (N_1085,N_616,N_946);
nor U1086 (N_1086,N_95,N_598);
nor U1087 (N_1087,N_519,N_474);
nand U1088 (N_1088,N_243,N_694);
xnor U1089 (N_1089,N_465,N_842);
or U1090 (N_1090,N_256,N_25);
nor U1091 (N_1091,N_96,N_412);
nand U1092 (N_1092,N_745,N_905);
and U1093 (N_1093,N_681,N_282);
nor U1094 (N_1094,N_340,N_34);
and U1095 (N_1095,N_940,N_723);
xor U1096 (N_1096,N_571,N_849);
and U1097 (N_1097,N_124,N_117);
or U1098 (N_1098,N_872,N_0);
nand U1099 (N_1099,N_797,N_236);
nand U1100 (N_1100,N_214,N_788);
or U1101 (N_1101,N_394,N_434);
nor U1102 (N_1102,N_551,N_504);
nand U1103 (N_1103,N_179,N_666);
and U1104 (N_1104,N_657,N_655);
nand U1105 (N_1105,N_262,N_156);
nor U1106 (N_1106,N_746,N_599);
nand U1107 (N_1107,N_229,N_123);
nor U1108 (N_1108,N_7,N_635);
xor U1109 (N_1109,N_430,N_57);
nand U1110 (N_1110,N_103,N_442);
and U1111 (N_1111,N_191,N_289);
nand U1112 (N_1112,N_17,N_467);
nor U1113 (N_1113,N_16,N_39);
xnor U1114 (N_1114,N_731,N_75);
xor U1115 (N_1115,N_748,N_94);
nand U1116 (N_1116,N_665,N_120);
and U1117 (N_1117,N_386,N_48);
xnor U1118 (N_1118,N_900,N_338);
xor U1119 (N_1119,N_292,N_388);
nand U1120 (N_1120,N_357,N_893);
and U1121 (N_1121,N_662,N_822);
or U1122 (N_1122,N_463,N_712);
and U1123 (N_1123,N_591,N_230);
and U1124 (N_1124,N_994,N_477);
xnor U1125 (N_1125,N_128,N_846);
or U1126 (N_1126,N_476,N_774);
xnor U1127 (N_1127,N_41,N_318);
nand U1128 (N_1128,N_464,N_682);
nor U1129 (N_1129,N_261,N_315);
xor U1130 (N_1130,N_483,N_276);
and U1131 (N_1131,N_137,N_643);
or U1132 (N_1132,N_232,N_851);
xor U1133 (N_1133,N_869,N_420);
nor U1134 (N_1134,N_459,N_967);
xor U1135 (N_1135,N_131,N_285);
and U1136 (N_1136,N_544,N_65);
and U1137 (N_1137,N_634,N_482);
nor U1138 (N_1138,N_522,N_478);
and U1139 (N_1139,N_91,N_101);
and U1140 (N_1140,N_527,N_341);
and U1141 (N_1141,N_950,N_21);
or U1142 (N_1142,N_136,N_534);
and U1143 (N_1143,N_892,N_660);
nand U1144 (N_1144,N_356,N_597);
nand U1145 (N_1145,N_624,N_915);
and U1146 (N_1146,N_547,N_785);
and U1147 (N_1147,N_162,N_426);
xor U1148 (N_1148,N_820,N_644);
xor U1149 (N_1149,N_675,N_493);
nand U1150 (N_1150,N_604,N_786);
and U1151 (N_1151,N_78,N_803);
nand U1152 (N_1152,N_639,N_367);
xor U1153 (N_1153,N_76,N_988);
nand U1154 (N_1154,N_708,N_89);
nand U1155 (N_1155,N_451,N_592);
or U1156 (N_1156,N_22,N_907);
xor U1157 (N_1157,N_258,N_815);
nand U1158 (N_1158,N_141,N_425);
xor U1159 (N_1159,N_611,N_855);
xor U1160 (N_1160,N_250,N_222);
and U1161 (N_1161,N_52,N_495);
nand U1162 (N_1162,N_569,N_358);
xnor U1163 (N_1163,N_444,N_404);
nor U1164 (N_1164,N_307,N_741);
or U1165 (N_1165,N_773,N_839);
and U1166 (N_1166,N_66,N_409);
nor U1167 (N_1167,N_335,N_721);
nor U1168 (N_1168,N_51,N_668);
xnor U1169 (N_1169,N_833,N_310);
xor U1170 (N_1170,N_40,N_287);
nand U1171 (N_1171,N_744,N_196);
or U1172 (N_1172,N_316,N_438);
and U1173 (N_1173,N_470,N_919);
and U1174 (N_1174,N_835,N_536);
and U1175 (N_1175,N_371,N_985);
nand U1176 (N_1176,N_628,N_100);
xor U1177 (N_1177,N_15,N_861);
and U1178 (N_1178,N_164,N_342);
xnor U1179 (N_1179,N_126,N_347);
xnor U1180 (N_1180,N_233,N_6);
or U1181 (N_1181,N_151,N_513);
and U1182 (N_1182,N_810,N_381);
nand U1183 (N_1183,N_868,N_274);
xnor U1184 (N_1184,N_181,N_825);
or U1185 (N_1185,N_778,N_362);
nor U1186 (N_1186,N_269,N_560);
or U1187 (N_1187,N_50,N_422);
nor U1188 (N_1188,N_715,N_935);
nand U1189 (N_1189,N_934,N_867);
and U1190 (N_1190,N_29,N_875);
and U1191 (N_1191,N_264,N_938);
nor U1192 (N_1192,N_90,N_305);
or U1193 (N_1193,N_698,N_427);
nor U1194 (N_1194,N_411,N_959);
and U1195 (N_1195,N_121,N_730);
xor U1196 (N_1196,N_771,N_458);
xor U1197 (N_1197,N_171,N_109);
or U1198 (N_1198,N_990,N_588);
or U1199 (N_1199,N_615,N_819);
nand U1200 (N_1200,N_725,N_637);
nor U1201 (N_1201,N_58,N_480);
nor U1202 (N_1202,N_218,N_987);
xnor U1203 (N_1203,N_139,N_799);
or U1204 (N_1204,N_735,N_737);
nand U1205 (N_1205,N_1,N_134);
and U1206 (N_1206,N_941,N_638);
and U1207 (N_1207,N_170,N_159);
and U1208 (N_1208,N_192,N_762);
and U1209 (N_1209,N_399,N_2);
xnor U1210 (N_1210,N_879,N_727);
nand U1211 (N_1211,N_506,N_829);
xor U1212 (N_1212,N_793,N_847);
nor U1213 (N_1213,N_818,N_334);
or U1214 (N_1214,N_537,N_740);
xor U1215 (N_1215,N_268,N_516);
xnor U1216 (N_1216,N_878,N_512);
nand U1217 (N_1217,N_138,N_667);
or U1218 (N_1218,N_583,N_132);
xnor U1219 (N_1219,N_750,N_749);
and U1220 (N_1220,N_704,N_312);
and U1221 (N_1221,N_800,N_369);
and U1222 (N_1222,N_494,N_553);
and U1223 (N_1223,N_161,N_929);
nand U1224 (N_1224,N_699,N_471);
and U1225 (N_1225,N_549,N_216);
xnor U1226 (N_1226,N_157,N_472);
nor U1227 (N_1227,N_199,N_116);
and U1228 (N_1228,N_286,N_784);
or U1229 (N_1229,N_627,N_99);
nand U1230 (N_1230,N_850,N_177);
or U1231 (N_1231,N_291,N_944);
nand U1232 (N_1232,N_297,N_782);
xnor U1233 (N_1233,N_672,N_806);
nand U1234 (N_1234,N_226,N_105);
or U1235 (N_1235,N_811,N_524);
nor U1236 (N_1236,N_882,N_397);
nor U1237 (N_1237,N_523,N_351);
or U1238 (N_1238,N_717,N_669);
and U1239 (N_1239,N_719,N_673);
or U1240 (N_1240,N_864,N_36);
xnor U1241 (N_1241,N_642,N_751);
xnor U1242 (N_1242,N_968,N_783);
nand U1243 (N_1243,N_240,N_317);
or U1244 (N_1244,N_518,N_272);
xor U1245 (N_1245,N_408,N_193);
or U1246 (N_1246,N_70,N_255);
nand U1247 (N_1247,N_969,N_186);
xnor U1248 (N_1248,N_921,N_350);
and U1249 (N_1249,N_726,N_903);
nor U1250 (N_1250,N_395,N_473);
or U1251 (N_1251,N_119,N_380);
xnor U1252 (N_1252,N_978,N_63);
and U1253 (N_1253,N_795,N_400);
or U1254 (N_1254,N_845,N_241);
nor U1255 (N_1255,N_251,N_452);
nor U1256 (N_1256,N_491,N_610);
xor U1257 (N_1257,N_174,N_219);
and U1258 (N_1258,N_541,N_686);
xor U1259 (N_1259,N_538,N_10);
nor U1260 (N_1260,N_753,N_421);
xnor U1261 (N_1261,N_336,N_194);
or U1262 (N_1262,N_223,N_263);
nand U1263 (N_1263,N_801,N_550);
nand U1264 (N_1264,N_270,N_410);
nor U1265 (N_1265,N_234,N_838);
and U1266 (N_1266,N_928,N_528);
nand U1267 (N_1267,N_966,N_593);
nor U1268 (N_1268,N_435,N_574);
nor U1269 (N_1269,N_446,N_937);
or U1270 (N_1270,N_792,N_772);
xor U1271 (N_1271,N_508,N_603);
or U1272 (N_1272,N_346,N_176);
nand U1273 (N_1273,N_706,N_448);
nor U1274 (N_1274,N_160,N_840);
xor U1275 (N_1275,N_652,N_777);
or U1276 (N_1276,N_209,N_479);
or U1277 (N_1277,N_72,N_352);
and U1278 (N_1278,N_439,N_178);
or U1279 (N_1279,N_764,N_142);
xnor U1280 (N_1280,N_697,N_953);
nor U1281 (N_1281,N_364,N_958);
xor U1282 (N_1282,N_814,N_481);
nor U1283 (N_1283,N_278,N_249);
and U1284 (N_1284,N_951,N_517);
nand U1285 (N_1285,N_497,N_244);
nor U1286 (N_1286,N_433,N_787);
xor U1287 (N_1287,N_837,N_909);
and U1288 (N_1288,N_543,N_280);
nand U1289 (N_1289,N_983,N_816);
xnor U1290 (N_1290,N_828,N_680);
or U1291 (N_1291,N_406,N_632);
nor U1292 (N_1292,N_502,N_607);
and U1293 (N_1293,N_54,N_617);
xnor U1294 (N_1294,N_654,N_752);
or U1295 (N_1295,N_257,N_754);
and U1296 (N_1296,N_700,N_225);
nand U1297 (N_1297,N_836,N_586);
xor U1298 (N_1298,N_325,N_572);
nor U1299 (N_1299,N_133,N_961);
and U1300 (N_1300,N_348,N_942);
and U1301 (N_1301,N_295,N_288);
xor U1302 (N_1302,N_415,N_913);
xor U1303 (N_1303,N_281,N_127);
or U1304 (N_1304,N_955,N_716);
or U1305 (N_1305,N_514,N_621);
nor U1306 (N_1306,N_939,N_821);
nor U1307 (N_1307,N_633,N_765);
xor U1308 (N_1308,N_894,N_143);
nor U1309 (N_1309,N_43,N_379);
nand U1310 (N_1310,N_180,N_885);
nor U1311 (N_1311,N_904,N_923);
nor U1312 (N_1312,N_974,N_857);
nor U1313 (N_1313,N_153,N_457);
nand U1314 (N_1314,N_488,N_182);
nor U1315 (N_1315,N_47,N_204);
xor U1316 (N_1316,N_854,N_881);
and U1317 (N_1317,N_239,N_68);
and U1318 (N_1318,N_578,N_656);
nor U1319 (N_1319,N_671,N_484);
nor U1320 (N_1320,N_349,N_498);
nand U1321 (N_1321,N_201,N_677);
nor U1322 (N_1322,N_450,N_189);
and U1323 (N_1323,N_62,N_556);
xnor U1324 (N_1324,N_343,N_429);
xor U1325 (N_1325,N_203,N_372);
and U1326 (N_1326,N_871,N_277);
xnor U1327 (N_1327,N_674,N_303);
xor U1328 (N_1328,N_242,N_834);
or U1329 (N_1329,N_93,N_407);
xnor U1330 (N_1330,N_794,N_943);
nand U1331 (N_1331,N_49,N_403);
xor U1332 (N_1332,N_977,N_374);
and U1333 (N_1333,N_812,N_30);
and U1334 (N_1334,N_525,N_521);
and U1335 (N_1335,N_526,N_602);
or U1336 (N_1336,N_555,N_302);
nor U1337 (N_1337,N_460,N_629);
and U1338 (N_1338,N_640,N_414);
xor U1339 (N_1339,N_922,N_808);
and U1340 (N_1340,N_843,N_389);
nand U1341 (N_1341,N_912,N_960);
and U1342 (N_1342,N_115,N_734);
or U1343 (N_1343,N_997,N_447);
nand U1344 (N_1344,N_859,N_238);
and U1345 (N_1345,N_582,N_418);
and U1346 (N_1346,N_780,N_314);
xor U1347 (N_1347,N_462,N_612);
and U1348 (N_1348,N_331,N_804);
or U1349 (N_1349,N_653,N_659);
or U1350 (N_1350,N_44,N_696);
or U1351 (N_1351,N_758,N_382);
nand U1352 (N_1352,N_530,N_97);
and U1353 (N_1353,N_917,N_805);
or U1354 (N_1354,N_962,N_273);
xor U1355 (N_1355,N_620,N_714);
and U1356 (N_1356,N_931,N_147);
nand U1357 (N_1357,N_323,N_92);
xor U1358 (N_1358,N_996,N_619);
and U1359 (N_1359,N_609,N_670);
xnor U1360 (N_1360,N_701,N_118);
xnor U1361 (N_1361,N_344,N_299);
and U1362 (N_1362,N_695,N_19);
nor U1363 (N_1363,N_11,N_933);
nand U1364 (N_1364,N_895,N_781);
nor U1365 (N_1365,N_954,N_441);
nor U1366 (N_1366,N_211,N_724);
and U1367 (N_1367,N_957,N_28);
and U1368 (N_1368,N_46,N_865);
or U1369 (N_1369,N_107,N_982);
nor U1370 (N_1370,N_532,N_129);
nand U1371 (N_1371,N_98,N_565);
and U1372 (N_1372,N_733,N_71);
nor U1373 (N_1373,N_140,N_924);
or U1374 (N_1374,N_284,N_796);
nand U1375 (N_1375,N_56,N_989);
or U1376 (N_1376,N_31,N_370);
xor U1377 (N_1377,N_265,N_630);
xor U1378 (N_1378,N_253,N_489);
or U1379 (N_1379,N_12,N_705);
xor U1380 (N_1380,N_999,N_776);
nand U1381 (N_1381,N_53,N_454);
or U1382 (N_1382,N_377,N_326);
nor U1383 (N_1383,N_790,N_930);
and U1384 (N_1384,N_566,N_826);
and U1385 (N_1385,N_948,N_899);
and U1386 (N_1386,N_768,N_77);
xor U1387 (N_1387,N_245,N_492);
or U1388 (N_1388,N_631,N_5);
xor U1389 (N_1389,N_330,N_313);
xor U1390 (N_1390,N_584,N_113);
xnor U1391 (N_1391,N_683,N_832);
nand U1392 (N_1392,N_387,N_144);
and U1393 (N_1393,N_74,N_468);
nand U1394 (N_1394,N_995,N_320);
or U1395 (N_1395,N_732,N_185);
xor U1396 (N_1396,N_254,N_183);
or U1397 (N_1397,N_767,N_73);
nor U1398 (N_1398,N_645,N_898);
or U1399 (N_1399,N_321,N_501);
or U1400 (N_1400,N_689,N_827);
nor U1401 (N_1401,N_260,N_486);
nor U1402 (N_1402,N_283,N_114);
and U1403 (N_1403,N_769,N_213);
xnor U1404 (N_1404,N_558,N_390);
and U1405 (N_1405,N_166,N_932);
or U1406 (N_1406,N_154,N_440);
xor U1407 (N_1407,N_601,N_998);
xnor U1408 (N_1408,N_873,N_548);
or U1409 (N_1409,N_964,N_80);
xor U1410 (N_1410,N_383,N_197);
nand U1411 (N_1411,N_300,N_32);
and U1412 (N_1412,N_791,N_963);
nor U1413 (N_1413,N_579,N_85);
xor U1414 (N_1414,N_595,N_45);
xor U1415 (N_1415,N_945,N_587);
xor U1416 (N_1416,N_728,N_824);
xor U1417 (N_1417,N_884,N_130);
and U1418 (N_1418,N_902,N_60);
xor U1419 (N_1419,N_152,N_809);
or U1420 (N_1420,N_594,N_858);
or U1421 (N_1421,N_205,N_59);
nand U1422 (N_1422,N_148,N_973);
nor U1423 (N_1423,N_247,N_515);
nand U1424 (N_1424,N_328,N_756);
or U1425 (N_1425,N_661,N_889);
nand U1426 (N_1426,N_391,N_82);
and U1427 (N_1427,N_927,N_187);
nand U1428 (N_1428,N_914,N_339);
xnor U1429 (N_1429,N_916,N_168);
nand U1430 (N_1430,N_332,N_64);
and U1431 (N_1431,N_789,N_709);
nand U1432 (N_1432,N_135,N_453);
or U1433 (N_1433,N_267,N_311);
nand U1434 (N_1434,N_980,N_685);
and U1435 (N_1435,N_86,N_545);
and U1436 (N_1436,N_590,N_163);
and U1437 (N_1437,N_647,N_9);
nand U1438 (N_1438,N_378,N_499);
or U1439 (N_1439,N_392,N_691);
xor U1440 (N_1440,N_304,N_870);
nor U1441 (N_1441,N_605,N_329);
and U1442 (N_1442,N_876,N_658);
nor U1443 (N_1443,N_760,N_770);
or U1444 (N_1444,N_511,N_228);
xor U1445 (N_1445,N_992,N_398);
nand U1446 (N_1446,N_993,N_169);
and U1447 (N_1447,N_880,N_580);
and U1448 (N_1448,N_431,N_110);
nand U1449 (N_1449,N_4,N_221);
nand U1450 (N_1450,N_33,N_540);
nand U1451 (N_1451,N_679,N_823);
or U1452 (N_1452,N_710,N_852);
xor U1453 (N_1453,N_862,N_184);
nand U1454 (N_1454,N_200,N_678);
xnor U1455 (N_1455,N_202,N_432);
nand U1456 (N_1456,N_886,N_684);
nor U1457 (N_1457,N_428,N_35);
nand U1458 (N_1458,N_802,N_888);
nand U1459 (N_1459,N_651,N_692);
xnor U1460 (N_1460,N_520,N_405);
xor U1461 (N_1461,N_13,N_373);
or U1462 (N_1462,N_970,N_206);
nand U1463 (N_1463,N_363,N_559);
and U1464 (N_1464,N_906,N_986);
nor U1465 (N_1465,N_622,N_55);
nand U1466 (N_1466,N_606,N_237);
nand U1467 (N_1467,N_991,N_360);
nor U1468 (N_1468,N_529,N_575);
xnor U1469 (N_1469,N_402,N_759);
and U1470 (N_1470,N_874,N_23);
nor U1471 (N_1471,N_296,N_926);
xor U1472 (N_1472,N_298,N_570);
nor U1473 (N_1473,N_61,N_466);
xnor U1474 (N_1474,N_891,N_711);
or U1475 (N_1475,N_3,N_863);
xnor U1476 (N_1476,N_416,N_911);
or U1477 (N_1477,N_337,N_88);
nor U1478 (N_1478,N_393,N_720);
or U1479 (N_1479,N_308,N_693);
and U1480 (N_1480,N_111,N_366);
xnor U1481 (N_1481,N_896,N_150);
nor U1482 (N_1482,N_108,N_505);
or U1483 (N_1483,N_830,N_531);
xnor U1484 (N_1484,N_87,N_419);
and U1485 (N_1485,N_210,N_424);
and U1486 (N_1486,N_856,N_220);
nand U1487 (N_1487,N_936,N_125);
nand U1488 (N_1488,N_585,N_104);
or U1489 (N_1489,N_198,N_766);
xor U1490 (N_1490,N_664,N_146);
nor U1491 (N_1491,N_546,N_577);
and U1492 (N_1492,N_853,N_648);
nand U1493 (N_1493,N_231,N_561);
xnor U1494 (N_1494,N_106,N_563);
nand U1495 (N_1495,N_755,N_562);
nor U1496 (N_1496,N_596,N_920);
or U1497 (N_1497,N_215,N_918);
xnor U1498 (N_1498,N_567,N_589);
nor U1499 (N_1499,N_779,N_259);
nand U1500 (N_1500,N_244,N_506);
and U1501 (N_1501,N_300,N_152);
and U1502 (N_1502,N_200,N_394);
or U1503 (N_1503,N_105,N_969);
nor U1504 (N_1504,N_826,N_724);
nor U1505 (N_1505,N_76,N_685);
xnor U1506 (N_1506,N_374,N_835);
xor U1507 (N_1507,N_440,N_455);
nand U1508 (N_1508,N_347,N_417);
or U1509 (N_1509,N_775,N_509);
and U1510 (N_1510,N_445,N_734);
xnor U1511 (N_1511,N_594,N_227);
and U1512 (N_1512,N_462,N_88);
nand U1513 (N_1513,N_257,N_366);
nand U1514 (N_1514,N_601,N_458);
or U1515 (N_1515,N_374,N_610);
and U1516 (N_1516,N_579,N_86);
nor U1517 (N_1517,N_475,N_288);
nor U1518 (N_1518,N_378,N_177);
nand U1519 (N_1519,N_189,N_212);
or U1520 (N_1520,N_164,N_786);
nor U1521 (N_1521,N_687,N_614);
and U1522 (N_1522,N_473,N_9);
nand U1523 (N_1523,N_13,N_198);
nor U1524 (N_1524,N_761,N_326);
nand U1525 (N_1525,N_131,N_636);
and U1526 (N_1526,N_752,N_998);
xnor U1527 (N_1527,N_590,N_774);
nand U1528 (N_1528,N_674,N_242);
and U1529 (N_1529,N_492,N_442);
xor U1530 (N_1530,N_336,N_504);
and U1531 (N_1531,N_961,N_49);
and U1532 (N_1532,N_452,N_96);
xor U1533 (N_1533,N_107,N_862);
xnor U1534 (N_1534,N_742,N_669);
xor U1535 (N_1535,N_103,N_420);
and U1536 (N_1536,N_588,N_815);
nand U1537 (N_1537,N_211,N_577);
or U1538 (N_1538,N_970,N_755);
and U1539 (N_1539,N_558,N_30);
xnor U1540 (N_1540,N_395,N_484);
nor U1541 (N_1541,N_839,N_370);
or U1542 (N_1542,N_319,N_507);
nand U1543 (N_1543,N_537,N_566);
and U1544 (N_1544,N_255,N_186);
or U1545 (N_1545,N_922,N_121);
nand U1546 (N_1546,N_323,N_868);
nor U1547 (N_1547,N_453,N_556);
and U1548 (N_1548,N_485,N_636);
or U1549 (N_1549,N_705,N_637);
nor U1550 (N_1550,N_300,N_25);
or U1551 (N_1551,N_775,N_180);
nor U1552 (N_1552,N_239,N_636);
and U1553 (N_1553,N_852,N_684);
or U1554 (N_1554,N_785,N_385);
xor U1555 (N_1555,N_621,N_110);
nand U1556 (N_1556,N_962,N_29);
nand U1557 (N_1557,N_194,N_916);
or U1558 (N_1558,N_375,N_672);
nand U1559 (N_1559,N_394,N_176);
nand U1560 (N_1560,N_338,N_404);
or U1561 (N_1561,N_725,N_497);
and U1562 (N_1562,N_391,N_328);
xor U1563 (N_1563,N_554,N_101);
nand U1564 (N_1564,N_325,N_208);
nor U1565 (N_1565,N_916,N_637);
xnor U1566 (N_1566,N_314,N_967);
nand U1567 (N_1567,N_878,N_217);
or U1568 (N_1568,N_563,N_636);
nand U1569 (N_1569,N_858,N_882);
xnor U1570 (N_1570,N_784,N_405);
nor U1571 (N_1571,N_697,N_244);
nor U1572 (N_1572,N_970,N_812);
nand U1573 (N_1573,N_934,N_803);
and U1574 (N_1574,N_48,N_677);
and U1575 (N_1575,N_566,N_358);
nand U1576 (N_1576,N_782,N_51);
or U1577 (N_1577,N_29,N_441);
or U1578 (N_1578,N_794,N_724);
nand U1579 (N_1579,N_425,N_909);
or U1580 (N_1580,N_408,N_712);
or U1581 (N_1581,N_66,N_530);
and U1582 (N_1582,N_302,N_898);
or U1583 (N_1583,N_467,N_139);
xnor U1584 (N_1584,N_991,N_751);
and U1585 (N_1585,N_229,N_165);
and U1586 (N_1586,N_193,N_842);
nand U1587 (N_1587,N_818,N_110);
nor U1588 (N_1588,N_77,N_844);
or U1589 (N_1589,N_123,N_463);
nor U1590 (N_1590,N_503,N_564);
xor U1591 (N_1591,N_542,N_526);
nand U1592 (N_1592,N_788,N_783);
nor U1593 (N_1593,N_970,N_321);
and U1594 (N_1594,N_726,N_84);
nand U1595 (N_1595,N_359,N_896);
xor U1596 (N_1596,N_877,N_750);
or U1597 (N_1597,N_990,N_282);
and U1598 (N_1598,N_296,N_999);
xnor U1599 (N_1599,N_555,N_654);
nor U1600 (N_1600,N_52,N_118);
and U1601 (N_1601,N_196,N_979);
xor U1602 (N_1602,N_189,N_166);
nand U1603 (N_1603,N_400,N_664);
and U1604 (N_1604,N_41,N_14);
nor U1605 (N_1605,N_780,N_686);
nand U1606 (N_1606,N_420,N_359);
or U1607 (N_1607,N_904,N_838);
nand U1608 (N_1608,N_868,N_749);
xor U1609 (N_1609,N_563,N_719);
or U1610 (N_1610,N_927,N_218);
or U1611 (N_1611,N_957,N_196);
and U1612 (N_1612,N_132,N_428);
and U1613 (N_1613,N_565,N_594);
and U1614 (N_1614,N_999,N_678);
nor U1615 (N_1615,N_566,N_945);
xnor U1616 (N_1616,N_12,N_414);
xor U1617 (N_1617,N_176,N_429);
nand U1618 (N_1618,N_443,N_932);
nor U1619 (N_1619,N_542,N_753);
and U1620 (N_1620,N_551,N_351);
or U1621 (N_1621,N_687,N_522);
and U1622 (N_1622,N_751,N_834);
xnor U1623 (N_1623,N_174,N_99);
xnor U1624 (N_1624,N_61,N_554);
nor U1625 (N_1625,N_4,N_235);
and U1626 (N_1626,N_338,N_107);
and U1627 (N_1627,N_774,N_318);
and U1628 (N_1628,N_491,N_267);
and U1629 (N_1629,N_950,N_37);
or U1630 (N_1630,N_5,N_779);
nor U1631 (N_1631,N_540,N_611);
nor U1632 (N_1632,N_983,N_26);
nand U1633 (N_1633,N_194,N_816);
or U1634 (N_1634,N_789,N_566);
nor U1635 (N_1635,N_440,N_744);
xnor U1636 (N_1636,N_565,N_199);
or U1637 (N_1637,N_596,N_683);
xnor U1638 (N_1638,N_767,N_442);
and U1639 (N_1639,N_273,N_323);
xor U1640 (N_1640,N_643,N_772);
xnor U1641 (N_1641,N_822,N_243);
nand U1642 (N_1642,N_825,N_905);
nor U1643 (N_1643,N_273,N_765);
or U1644 (N_1644,N_483,N_230);
xnor U1645 (N_1645,N_307,N_929);
nand U1646 (N_1646,N_211,N_984);
xnor U1647 (N_1647,N_580,N_426);
and U1648 (N_1648,N_106,N_843);
nand U1649 (N_1649,N_667,N_781);
and U1650 (N_1650,N_606,N_200);
xnor U1651 (N_1651,N_316,N_346);
nand U1652 (N_1652,N_634,N_201);
xnor U1653 (N_1653,N_465,N_18);
or U1654 (N_1654,N_566,N_205);
or U1655 (N_1655,N_67,N_144);
xnor U1656 (N_1656,N_892,N_624);
nor U1657 (N_1657,N_285,N_639);
xnor U1658 (N_1658,N_32,N_478);
and U1659 (N_1659,N_944,N_757);
and U1660 (N_1660,N_356,N_277);
and U1661 (N_1661,N_318,N_88);
and U1662 (N_1662,N_191,N_667);
xnor U1663 (N_1663,N_470,N_682);
or U1664 (N_1664,N_355,N_750);
nor U1665 (N_1665,N_359,N_582);
and U1666 (N_1666,N_319,N_619);
xnor U1667 (N_1667,N_19,N_198);
or U1668 (N_1668,N_934,N_452);
nand U1669 (N_1669,N_696,N_727);
or U1670 (N_1670,N_327,N_332);
nand U1671 (N_1671,N_198,N_666);
nand U1672 (N_1672,N_598,N_32);
xor U1673 (N_1673,N_801,N_755);
or U1674 (N_1674,N_599,N_365);
xnor U1675 (N_1675,N_618,N_954);
or U1676 (N_1676,N_948,N_16);
xor U1677 (N_1677,N_116,N_129);
or U1678 (N_1678,N_887,N_843);
or U1679 (N_1679,N_968,N_690);
nand U1680 (N_1680,N_621,N_811);
and U1681 (N_1681,N_989,N_878);
and U1682 (N_1682,N_408,N_73);
or U1683 (N_1683,N_419,N_193);
nor U1684 (N_1684,N_316,N_258);
and U1685 (N_1685,N_308,N_463);
nand U1686 (N_1686,N_364,N_761);
nand U1687 (N_1687,N_697,N_545);
and U1688 (N_1688,N_363,N_293);
nor U1689 (N_1689,N_418,N_17);
nand U1690 (N_1690,N_559,N_739);
xnor U1691 (N_1691,N_825,N_724);
nor U1692 (N_1692,N_521,N_822);
or U1693 (N_1693,N_312,N_736);
or U1694 (N_1694,N_409,N_437);
or U1695 (N_1695,N_343,N_909);
nand U1696 (N_1696,N_35,N_442);
and U1697 (N_1697,N_717,N_169);
xor U1698 (N_1698,N_537,N_431);
xor U1699 (N_1699,N_723,N_716);
nand U1700 (N_1700,N_56,N_533);
nand U1701 (N_1701,N_402,N_758);
and U1702 (N_1702,N_516,N_75);
nand U1703 (N_1703,N_394,N_239);
or U1704 (N_1704,N_209,N_323);
nor U1705 (N_1705,N_366,N_835);
nand U1706 (N_1706,N_511,N_503);
nand U1707 (N_1707,N_737,N_548);
nand U1708 (N_1708,N_196,N_76);
and U1709 (N_1709,N_321,N_308);
xor U1710 (N_1710,N_979,N_400);
nand U1711 (N_1711,N_224,N_286);
or U1712 (N_1712,N_109,N_180);
xnor U1713 (N_1713,N_643,N_248);
xnor U1714 (N_1714,N_675,N_200);
nor U1715 (N_1715,N_808,N_249);
xor U1716 (N_1716,N_80,N_763);
and U1717 (N_1717,N_188,N_568);
and U1718 (N_1718,N_435,N_326);
nor U1719 (N_1719,N_686,N_80);
or U1720 (N_1720,N_149,N_553);
or U1721 (N_1721,N_117,N_891);
and U1722 (N_1722,N_431,N_118);
and U1723 (N_1723,N_219,N_911);
or U1724 (N_1724,N_12,N_962);
xnor U1725 (N_1725,N_199,N_693);
xor U1726 (N_1726,N_862,N_460);
and U1727 (N_1727,N_254,N_842);
and U1728 (N_1728,N_163,N_505);
nor U1729 (N_1729,N_427,N_663);
xor U1730 (N_1730,N_727,N_846);
or U1731 (N_1731,N_443,N_717);
xor U1732 (N_1732,N_502,N_255);
nand U1733 (N_1733,N_257,N_913);
nor U1734 (N_1734,N_909,N_490);
nor U1735 (N_1735,N_129,N_96);
nor U1736 (N_1736,N_205,N_295);
and U1737 (N_1737,N_833,N_607);
nand U1738 (N_1738,N_513,N_978);
nand U1739 (N_1739,N_16,N_402);
nor U1740 (N_1740,N_425,N_635);
or U1741 (N_1741,N_886,N_667);
or U1742 (N_1742,N_26,N_96);
or U1743 (N_1743,N_875,N_633);
nor U1744 (N_1744,N_957,N_940);
nor U1745 (N_1745,N_633,N_466);
xnor U1746 (N_1746,N_693,N_15);
nand U1747 (N_1747,N_678,N_728);
or U1748 (N_1748,N_273,N_869);
xnor U1749 (N_1749,N_421,N_438);
nand U1750 (N_1750,N_362,N_564);
and U1751 (N_1751,N_343,N_630);
and U1752 (N_1752,N_239,N_2);
nand U1753 (N_1753,N_497,N_697);
xnor U1754 (N_1754,N_451,N_209);
nand U1755 (N_1755,N_931,N_27);
nor U1756 (N_1756,N_970,N_937);
nor U1757 (N_1757,N_577,N_56);
nand U1758 (N_1758,N_249,N_681);
and U1759 (N_1759,N_20,N_694);
nor U1760 (N_1760,N_647,N_393);
nand U1761 (N_1761,N_431,N_500);
and U1762 (N_1762,N_584,N_709);
nor U1763 (N_1763,N_722,N_450);
and U1764 (N_1764,N_88,N_300);
nor U1765 (N_1765,N_852,N_902);
and U1766 (N_1766,N_484,N_530);
nand U1767 (N_1767,N_506,N_584);
nand U1768 (N_1768,N_378,N_878);
xor U1769 (N_1769,N_978,N_870);
and U1770 (N_1770,N_463,N_726);
or U1771 (N_1771,N_330,N_806);
nand U1772 (N_1772,N_215,N_758);
nand U1773 (N_1773,N_872,N_345);
and U1774 (N_1774,N_792,N_243);
and U1775 (N_1775,N_319,N_372);
nor U1776 (N_1776,N_65,N_899);
nor U1777 (N_1777,N_520,N_165);
nand U1778 (N_1778,N_3,N_894);
or U1779 (N_1779,N_283,N_111);
or U1780 (N_1780,N_404,N_198);
nand U1781 (N_1781,N_34,N_99);
nand U1782 (N_1782,N_989,N_164);
xnor U1783 (N_1783,N_922,N_940);
or U1784 (N_1784,N_27,N_108);
nor U1785 (N_1785,N_286,N_915);
nor U1786 (N_1786,N_114,N_395);
and U1787 (N_1787,N_749,N_788);
and U1788 (N_1788,N_704,N_710);
or U1789 (N_1789,N_177,N_355);
xnor U1790 (N_1790,N_153,N_143);
xor U1791 (N_1791,N_726,N_136);
or U1792 (N_1792,N_306,N_382);
xnor U1793 (N_1793,N_480,N_148);
nand U1794 (N_1794,N_913,N_10);
and U1795 (N_1795,N_72,N_620);
nand U1796 (N_1796,N_960,N_207);
xnor U1797 (N_1797,N_390,N_275);
or U1798 (N_1798,N_907,N_482);
nand U1799 (N_1799,N_304,N_970);
xnor U1800 (N_1800,N_525,N_80);
or U1801 (N_1801,N_21,N_727);
or U1802 (N_1802,N_978,N_922);
nor U1803 (N_1803,N_553,N_890);
xnor U1804 (N_1804,N_105,N_632);
nor U1805 (N_1805,N_256,N_549);
or U1806 (N_1806,N_387,N_247);
xnor U1807 (N_1807,N_581,N_101);
xor U1808 (N_1808,N_347,N_472);
nand U1809 (N_1809,N_643,N_587);
and U1810 (N_1810,N_29,N_822);
nor U1811 (N_1811,N_134,N_76);
or U1812 (N_1812,N_795,N_547);
xor U1813 (N_1813,N_901,N_282);
nand U1814 (N_1814,N_279,N_486);
and U1815 (N_1815,N_595,N_768);
or U1816 (N_1816,N_982,N_823);
xnor U1817 (N_1817,N_498,N_874);
or U1818 (N_1818,N_848,N_561);
xnor U1819 (N_1819,N_370,N_809);
and U1820 (N_1820,N_232,N_754);
and U1821 (N_1821,N_575,N_562);
or U1822 (N_1822,N_501,N_264);
and U1823 (N_1823,N_959,N_694);
xor U1824 (N_1824,N_320,N_400);
xnor U1825 (N_1825,N_582,N_829);
and U1826 (N_1826,N_259,N_798);
nand U1827 (N_1827,N_603,N_979);
nor U1828 (N_1828,N_24,N_204);
nor U1829 (N_1829,N_915,N_648);
and U1830 (N_1830,N_582,N_850);
or U1831 (N_1831,N_210,N_482);
and U1832 (N_1832,N_937,N_849);
xnor U1833 (N_1833,N_328,N_428);
nor U1834 (N_1834,N_245,N_210);
and U1835 (N_1835,N_105,N_663);
and U1836 (N_1836,N_734,N_178);
and U1837 (N_1837,N_383,N_317);
and U1838 (N_1838,N_787,N_712);
or U1839 (N_1839,N_142,N_618);
nand U1840 (N_1840,N_104,N_411);
or U1841 (N_1841,N_188,N_789);
xor U1842 (N_1842,N_845,N_149);
nor U1843 (N_1843,N_920,N_479);
nand U1844 (N_1844,N_478,N_107);
nand U1845 (N_1845,N_219,N_448);
xnor U1846 (N_1846,N_481,N_337);
nand U1847 (N_1847,N_520,N_13);
or U1848 (N_1848,N_991,N_830);
nand U1849 (N_1849,N_137,N_14);
nor U1850 (N_1850,N_31,N_762);
nor U1851 (N_1851,N_0,N_894);
and U1852 (N_1852,N_43,N_176);
nor U1853 (N_1853,N_798,N_176);
and U1854 (N_1854,N_852,N_935);
xnor U1855 (N_1855,N_932,N_364);
or U1856 (N_1856,N_486,N_365);
nand U1857 (N_1857,N_879,N_693);
and U1858 (N_1858,N_87,N_673);
xor U1859 (N_1859,N_897,N_551);
xor U1860 (N_1860,N_106,N_599);
nand U1861 (N_1861,N_813,N_901);
and U1862 (N_1862,N_518,N_279);
nor U1863 (N_1863,N_679,N_796);
xor U1864 (N_1864,N_565,N_253);
or U1865 (N_1865,N_234,N_214);
xor U1866 (N_1866,N_90,N_678);
nor U1867 (N_1867,N_853,N_601);
and U1868 (N_1868,N_8,N_666);
or U1869 (N_1869,N_187,N_91);
or U1870 (N_1870,N_788,N_737);
xnor U1871 (N_1871,N_897,N_164);
xor U1872 (N_1872,N_43,N_120);
or U1873 (N_1873,N_8,N_520);
xor U1874 (N_1874,N_231,N_884);
nand U1875 (N_1875,N_416,N_240);
and U1876 (N_1876,N_49,N_688);
nand U1877 (N_1877,N_753,N_620);
nand U1878 (N_1878,N_88,N_834);
xor U1879 (N_1879,N_392,N_980);
and U1880 (N_1880,N_992,N_210);
or U1881 (N_1881,N_151,N_831);
and U1882 (N_1882,N_699,N_348);
or U1883 (N_1883,N_579,N_967);
and U1884 (N_1884,N_559,N_835);
and U1885 (N_1885,N_186,N_455);
or U1886 (N_1886,N_554,N_249);
nor U1887 (N_1887,N_102,N_52);
or U1888 (N_1888,N_393,N_372);
nand U1889 (N_1889,N_764,N_526);
and U1890 (N_1890,N_952,N_73);
xor U1891 (N_1891,N_124,N_202);
nor U1892 (N_1892,N_530,N_48);
nand U1893 (N_1893,N_944,N_895);
or U1894 (N_1894,N_837,N_724);
xnor U1895 (N_1895,N_992,N_43);
xor U1896 (N_1896,N_597,N_224);
or U1897 (N_1897,N_325,N_903);
or U1898 (N_1898,N_686,N_860);
nor U1899 (N_1899,N_430,N_691);
and U1900 (N_1900,N_564,N_795);
or U1901 (N_1901,N_918,N_895);
nor U1902 (N_1902,N_989,N_582);
nand U1903 (N_1903,N_609,N_838);
and U1904 (N_1904,N_754,N_245);
nand U1905 (N_1905,N_992,N_460);
nor U1906 (N_1906,N_84,N_299);
xor U1907 (N_1907,N_816,N_402);
and U1908 (N_1908,N_602,N_329);
xor U1909 (N_1909,N_127,N_988);
xor U1910 (N_1910,N_330,N_582);
nand U1911 (N_1911,N_288,N_685);
nor U1912 (N_1912,N_406,N_896);
or U1913 (N_1913,N_850,N_316);
nand U1914 (N_1914,N_830,N_150);
nor U1915 (N_1915,N_298,N_705);
xnor U1916 (N_1916,N_582,N_450);
and U1917 (N_1917,N_874,N_956);
nor U1918 (N_1918,N_233,N_930);
nand U1919 (N_1919,N_537,N_956);
nor U1920 (N_1920,N_614,N_225);
xnor U1921 (N_1921,N_82,N_727);
and U1922 (N_1922,N_459,N_468);
or U1923 (N_1923,N_389,N_608);
nor U1924 (N_1924,N_584,N_578);
nor U1925 (N_1925,N_50,N_671);
or U1926 (N_1926,N_906,N_884);
nor U1927 (N_1927,N_240,N_437);
xnor U1928 (N_1928,N_965,N_668);
nor U1929 (N_1929,N_403,N_560);
nor U1930 (N_1930,N_495,N_659);
xnor U1931 (N_1931,N_966,N_990);
nor U1932 (N_1932,N_881,N_157);
or U1933 (N_1933,N_544,N_787);
and U1934 (N_1934,N_503,N_424);
xor U1935 (N_1935,N_273,N_319);
and U1936 (N_1936,N_394,N_64);
or U1937 (N_1937,N_205,N_60);
nand U1938 (N_1938,N_331,N_806);
nand U1939 (N_1939,N_376,N_304);
and U1940 (N_1940,N_207,N_981);
nor U1941 (N_1941,N_431,N_332);
xor U1942 (N_1942,N_598,N_295);
nor U1943 (N_1943,N_80,N_500);
and U1944 (N_1944,N_841,N_998);
nand U1945 (N_1945,N_664,N_191);
or U1946 (N_1946,N_838,N_104);
xnor U1947 (N_1947,N_435,N_959);
or U1948 (N_1948,N_467,N_54);
or U1949 (N_1949,N_328,N_181);
or U1950 (N_1950,N_527,N_815);
and U1951 (N_1951,N_100,N_703);
or U1952 (N_1952,N_63,N_543);
nor U1953 (N_1953,N_394,N_786);
or U1954 (N_1954,N_779,N_98);
xor U1955 (N_1955,N_285,N_602);
or U1956 (N_1956,N_151,N_928);
nand U1957 (N_1957,N_629,N_832);
nor U1958 (N_1958,N_974,N_589);
xor U1959 (N_1959,N_591,N_983);
nand U1960 (N_1960,N_308,N_554);
and U1961 (N_1961,N_538,N_748);
nand U1962 (N_1962,N_688,N_883);
and U1963 (N_1963,N_19,N_554);
or U1964 (N_1964,N_630,N_35);
and U1965 (N_1965,N_643,N_717);
nor U1966 (N_1966,N_564,N_63);
or U1967 (N_1967,N_135,N_38);
nor U1968 (N_1968,N_119,N_956);
nor U1969 (N_1969,N_991,N_747);
and U1970 (N_1970,N_307,N_678);
xor U1971 (N_1971,N_881,N_66);
or U1972 (N_1972,N_91,N_108);
nand U1973 (N_1973,N_576,N_358);
nor U1974 (N_1974,N_305,N_810);
or U1975 (N_1975,N_532,N_415);
xnor U1976 (N_1976,N_28,N_926);
xor U1977 (N_1977,N_272,N_968);
nand U1978 (N_1978,N_31,N_304);
xnor U1979 (N_1979,N_366,N_619);
nor U1980 (N_1980,N_491,N_929);
or U1981 (N_1981,N_673,N_339);
nand U1982 (N_1982,N_190,N_724);
nor U1983 (N_1983,N_495,N_769);
nor U1984 (N_1984,N_251,N_785);
xnor U1985 (N_1985,N_267,N_948);
nor U1986 (N_1986,N_658,N_305);
nand U1987 (N_1987,N_712,N_859);
nand U1988 (N_1988,N_381,N_692);
or U1989 (N_1989,N_141,N_40);
nor U1990 (N_1990,N_383,N_747);
or U1991 (N_1991,N_544,N_470);
nor U1992 (N_1992,N_269,N_768);
and U1993 (N_1993,N_737,N_68);
and U1994 (N_1994,N_265,N_133);
nor U1995 (N_1995,N_894,N_349);
xor U1996 (N_1996,N_839,N_614);
and U1997 (N_1997,N_8,N_647);
or U1998 (N_1998,N_326,N_912);
nor U1999 (N_1999,N_987,N_820);
xor U2000 (N_2000,N_1734,N_1462);
or U2001 (N_2001,N_1416,N_1547);
nand U2002 (N_2002,N_1459,N_1347);
or U2003 (N_2003,N_1889,N_1259);
and U2004 (N_2004,N_1074,N_1905);
xor U2005 (N_2005,N_1831,N_1963);
nand U2006 (N_2006,N_1010,N_1062);
xnor U2007 (N_2007,N_1508,N_1884);
xnor U2008 (N_2008,N_1495,N_1470);
xor U2009 (N_2009,N_1932,N_1761);
or U2010 (N_2010,N_1853,N_1035);
and U2011 (N_2011,N_1634,N_1666);
xnor U2012 (N_2012,N_1450,N_1431);
nand U2013 (N_2013,N_1673,N_1807);
nor U2014 (N_2014,N_1435,N_1935);
nor U2015 (N_2015,N_1391,N_1419);
or U2016 (N_2016,N_1771,N_1927);
or U2017 (N_2017,N_1638,N_1886);
xor U2018 (N_2018,N_1162,N_1251);
nand U2019 (N_2019,N_1876,N_1755);
nor U2020 (N_2020,N_1401,N_1464);
xnor U2021 (N_2021,N_1517,N_1710);
nand U2022 (N_2022,N_1155,N_1285);
nor U2023 (N_2023,N_1213,N_1306);
nand U2024 (N_2024,N_1972,N_1539);
xor U2025 (N_2025,N_1667,N_1240);
or U2026 (N_2026,N_1489,N_1036);
nor U2027 (N_2027,N_1848,N_1530);
nand U2028 (N_2028,N_1990,N_1013);
or U2029 (N_2029,N_1800,N_1523);
nand U2030 (N_2030,N_1438,N_1718);
and U2031 (N_2031,N_1882,N_1366);
xnor U2032 (N_2032,N_1555,N_1049);
or U2033 (N_2033,N_1510,N_1891);
nor U2034 (N_2034,N_1135,N_1146);
nand U2035 (N_2035,N_1015,N_1749);
nor U2036 (N_2036,N_1016,N_1744);
nor U2037 (N_2037,N_1389,N_1448);
and U2038 (N_2038,N_1370,N_1936);
xor U2039 (N_2039,N_1997,N_1287);
nor U2040 (N_2040,N_1014,N_1242);
or U2041 (N_2041,N_1696,N_1962);
nand U2042 (N_2042,N_1823,N_1143);
and U2043 (N_2043,N_1473,N_1437);
xnor U2044 (N_2044,N_1356,N_1982);
nor U2045 (N_2045,N_1186,N_1930);
and U2046 (N_2046,N_1158,N_1989);
nand U2047 (N_2047,N_1501,N_1652);
nor U2048 (N_2048,N_1184,N_1579);
nor U2049 (N_2049,N_1388,N_1960);
xnor U2050 (N_2050,N_1142,N_1782);
nor U2051 (N_2051,N_1797,N_1918);
nor U2052 (N_2052,N_1599,N_1225);
and U2053 (N_2053,N_1502,N_1252);
xor U2054 (N_2054,N_1767,N_1392);
nor U2055 (N_2055,N_1527,N_1828);
nand U2056 (N_2056,N_1360,N_1157);
or U2057 (N_2057,N_1913,N_1613);
nor U2058 (N_2058,N_1938,N_1382);
xor U2059 (N_2059,N_1421,N_1039);
xor U2060 (N_2060,N_1921,N_1808);
xor U2061 (N_2061,N_1358,N_1364);
nor U2062 (N_2062,N_1716,N_1955);
or U2063 (N_2063,N_1603,N_1496);
xor U2064 (N_2064,N_1660,N_1646);
xnor U2065 (N_2065,N_1053,N_1228);
and U2066 (N_2066,N_1139,N_1060);
and U2067 (N_2067,N_1798,N_1407);
nor U2068 (N_2068,N_1304,N_1846);
nor U2069 (N_2069,N_1693,N_1261);
xor U2070 (N_2070,N_1316,N_1885);
and U2071 (N_2071,N_1216,N_1958);
xor U2072 (N_2072,N_1558,N_1959);
and U2073 (N_2073,N_1217,N_1094);
and U2074 (N_2074,N_1293,N_1363);
or U2075 (N_2075,N_1608,N_1441);
or U2076 (N_2076,N_1461,N_1737);
or U2077 (N_2077,N_1103,N_1125);
xnor U2078 (N_2078,N_1170,N_1888);
nand U2079 (N_2079,N_1815,N_1398);
or U2080 (N_2080,N_1832,N_1690);
nand U2081 (N_2081,N_1999,N_1500);
nand U2082 (N_2082,N_1116,N_1159);
xor U2083 (N_2083,N_1107,N_1641);
and U2084 (N_2084,N_1453,N_1611);
nor U2085 (N_2085,N_1499,N_1195);
nand U2086 (N_2086,N_1816,N_1271);
nor U2087 (N_2087,N_1911,N_1210);
nand U2088 (N_2088,N_1393,N_1790);
nor U2089 (N_2089,N_1004,N_1181);
and U2090 (N_2090,N_1903,N_1319);
nand U2091 (N_2091,N_1102,N_1747);
xnor U2092 (N_2092,N_1514,N_1731);
nand U2093 (N_2093,N_1837,N_1680);
or U2094 (N_2094,N_1325,N_1650);
nor U2095 (N_2095,N_1410,N_1354);
and U2096 (N_2096,N_1099,N_1223);
xor U2097 (N_2097,N_1739,N_1144);
nand U2098 (N_2098,N_1402,N_1909);
and U2099 (N_2099,N_1339,N_1804);
or U2100 (N_2100,N_1414,N_1200);
xor U2101 (N_2101,N_1505,N_1332);
nand U2102 (N_2102,N_1824,N_1208);
or U2103 (N_2103,N_1668,N_1374);
xor U2104 (N_2104,N_1260,N_1097);
nand U2105 (N_2105,N_1685,N_1561);
xnor U2106 (N_2106,N_1621,N_1644);
nor U2107 (N_2107,N_1289,N_1156);
or U2108 (N_2108,N_1653,N_1536);
nand U2109 (N_2109,N_1232,N_1408);
nor U2110 (N_2110,N_1780,N_1745);
xnor U2111 (N_2111,N_1413,N_1597);
or U2112 (N_2112,N_1481,N_1753);
nor U2113 (N_2113,N_1236,N_1709);
nor U2114 (N_2114,N_1836,N_1342);
and U2115 (N_2115,N_1017,N_1629);
or U2116 (N_2116,N_1040,N_1104);
xor U2117 (N_2117,N_1073,N_1023);
xor U2118 (N_2118,N_1132,N_1185);
nor U2119 (N_2119,N_1840,N_1406);
nor U2120 (N_2120,N_1434,N_1340);
and U2121 (N_2121,N_1041,N_1020);
nor U2122 (N_2122,N_1814,N_1371);
nor U2123 (N_2123,N_1549,N_1246);
and U2124 (N_2124,N_1276,N_1605);
nand U2125 (N_2125,N_1609,N_1063);
xnor U2126 (N_2126,N_1328,N_1108);
nand U2127 (N_2127,N_1244,N_1861);
xnor U2128 (N_2128,N_1148,N_1830);
and U2129 (N_2129,N_1803,N_1770);
and U2130 (N_2130,N_1738,N_1268);
nor U2131 (N_2131,N_1351,N_1983);
or U2132 (N_2132,N_1720,N_1320);
nand U2133 (N_2133,N_1671,N_1967);
and U2134 (N_2134,N_1839,N_1973);
and U2135 (N_2135,N_1559,N_1065);
nor U2136 (N_2136,N_1458,N_1521);
xor U2137 (N_2137,N_1772,N_1865);
xor U2138 (N_2138,N_1429,N_1851);
xor U2139 (N_2139,N_1949,N_1457);
xor U2140 (N_2140,N_1551,N_1492);
nor U2141 (N_2141,N_1593,N_1266);
and U2142 (N_2142,N_1301,N_1706);
and U2143 (N_2143,N_1858,N_1842);
nand U2144 (N_2144,N_1309,N_1651);
nand U2145 (N_2145,N_1787,N_1532);
and U2146 (N_2146,N_1866,N_1031);
xnor U2147 (N_2147,N_1606,N_1460);
and U2148 (N_2148,N_1415,N_1026);
nand U2149 (N_2149,N_1472,N_1783);
nor U2150 (N_2150,N_1519,N_1980);
xor U2151 (N_2151,N_1996,N_1140);
or U2152 (N_2152,N_1326,N_1984);
or U2153 (N_2153,N_1614,N_1484);
nor U2154 (N_2154,N_1684,N_1698);
and U2155 (N_2155,N_1722,N_1257);
nand U2156 (N_2156,N_1211,N_1528);
nand U2157 (N_2157,N_1488,N_1595);
nand U2158 (N_2158,N_1399,N_1456);
and U2159 (N_2159,N_1096,N_1190);
nand U2160 (N_2160,N_1029,N_1544);
nand U2161 (N_2161,N_1970,N_1265);
and U2162 (N_2162,N_1243,N_1754);
xor U2163 (N_2163,N_1682,N_1471);
xor U2164 (N_2164,N_1656,N_1942);
xor U2165 (N_2165,N_1833,N_1677);
xor U2166 (N_2166,N_1119,N_1292);
or U2167 (N_2167,N_1198,N_1580);
or U2168 (N_2168,N_1288,N_1428);
nand U2169 (N_2169,N_1610,N_1679);
xor U2170 (N_2170,N_1577,N_1929);
nand U2171 (N_2171,N_1589,N_1047);
nand U2172 (N_2172,N_1663,N_1134);
and U2173 (N_2173,N_1333,N_1030);
nor U2174 (N_2174,N_1919,N_1707);
and U2175 (N_2175,N_1160,N_1843);
or U2176 (N_2176,N_1713,N_1486);
xor U2177 (N_2177,N_1516,N_1801);
nand U2178 (N_2178,N_1191,N_1147);
xor U2179 (N_2179,N_1150,N_1893);
and U2180 (N_2180,N_1943,N_1114);
nand U2181 (N_2181,N_1623,N_1655);
xnor U2182 (N_2182,N_1222,N_1057);
nand U2183 (N_2183,N_1620,N_1979);
nand U2184 (N_2184,N_1341,N_1338);
xnor U2185 (N_2185,N_1052,N_1786);
nor U2186 (N_2186,N_1440,N_1986);
or U2187 (N_2187,N_1506,N_1068);
nand U2188 (N_2188,N_1477,N_1249);
and U2189 (N_2189,N_1080,N_1708);
nand U2190 (N_2190,N_1897,N_1977);
nor U2191 (N_2191,N_1400,N_1542);
nor U2192 (N_2192,N_1504,N_1587);
or U2193 (N_2193,N_1088,N_1622);
and U2194 (N_2194,N_1733,N_1083);
nand U2195 (N_2195,N_1604,N_1231);
xor U2196 (N_2196,N_1649,N_1908);
nand U2197 (N_2197,N_1335,N_1695);
or U2198 (N_2198,N_1046,N_1479);
nor U2199 (N_2199,N_1939,N_1238);
and U2200 (N_2200,N_1256,N_1728);
xor U2201 (N_2201,N_1409,N_1571);
and U2202 (N_2202,N_1183,N_1529);
or U2203 (N_2203,N_1957,N_1475);
nor U2204 (N_2204,N_1233,N_1331);
nand U2205 (N_2205,N_1379,N_1618);
nand U2206 (N_2206,N_1284,N_1381);
nand U2207 (N_2207,N_1002,N_1037);
xnor U2208 (N_2208,N_1896,N_1133);
and U2209 (N_2209,N_1491,N_1813);
or U2210 (N_2210,N_1607,N_1018);
and U2211 (N_2211,N_1138,N_1785);
xor U2212 (N_2212,N_1601,N_1303);
nand U2213 (N_2213,N_1974,N_1359);
nor U2214 (N_2214,N_1697,N_1075);
nor U2215 (N_2215,N_1164,N_1550);
or U2216 (N_2216,N_1054,N_1206);
xor U2217 (N_2217,N_1845,N_1255);
or U2218 (N_2218,N_1291,N_1890);
or U2219 (N_2219,N_1205,N_1556);
nand U2220 (N_2220,N_1446,N_1533);
nor U2221 (N_2221,N_1567,N_1071);
nand U2222 (N_2222,N_1688,N_1854);
and U2223 (N_2223,N_1793,N_1920);
nor U2224 (N_2224,N_1910,N_1978);
or U2225 (N_2225,N_1283,N_1730);
and U2226 (N_2226,N_1686,N_1027);
or U2227 (N_2227,N_1177,N_1072);
and U2228 (N_2228,N_1005,N_1277);
nand U2229 (N_2229,N_1365,N_1476);
or U2230 (N_2230,N_1215,N_1353);
nand U2231 (N_2231,N_1070,N_1992);
xor U2232 (N_2232,N_1025,N_1873);
nand U2233 (N_2233,N_1424,N_1384);
nand U2234 (N_2234,N_1534,N_1313);
or U2235 (N_2235,N_1906,N_1724);
nand U2236 (N_2236,N_1821,N_1746);
nand U2237 (N_2237,N_1681,N_1509);
xor U2238 (N_2238,N_1372,N_1971);
or U2239 (N_2239,N_1714,N_1067);
nor U2240 (N_2240,N_1993,N_1221);
nand U2241 (N_2241,N_1498,N_1664);
and U2242 (N_2242,N_1554,N_1180);
nand U2243 (N_2243,N_1480,N_1113);
nand U2244 (N_2244,N_1482,N_1220);
and U2245 (N_2245,N_1760,N_1563);
and U2246 (N_2246,N_1825,N_1254);
xor U2247 (N_2247,N_1058,N_1574);
nor U2248 (N_2248,N_1868,N_1172);
nand U2249 (N_2249,N_1590,N_1762);
nand U2250 (N_2250,N_1581,N_1654);
xnor U2251 (N_2251,N_1166,N_1011);
nor U2252 (N_2252,N_1427,N_1672);
nand U2253 (N_2253,N_1169,N_1087);
or U2254 (N_2254,N_1230,N_1084);
or U2255 (N_2255,N_1628,N_1055);
nor U2256 (N_2256,N_1619,N_1021);
and U2257 (N_2257,N_1545,N_1892);
xnor U2258 (N_2258,N_1615,N_1859);
xnor U2259 (N_2259,N_1658,N_1178);
nor U2260 (N_2260,N_1091,N_1145);
xnor U2261 (N_2261,N_1214,N_1701);
and U2262 (N_2262,N_1578,N_1552);
xnor U2263 (N_2263,N_1076,N_1700);
xnor U2264 (N_2264,N_1447,N_1901);
or U2265 (N_2265,N_1841,N_1451);
nor U2266 (N_2266,N_1759,N_1857);
and U2267 (N_2267,N_1925,N_1361);
nor U2268 (N_2268,N_1442,N_1637);
or U2269 (N_2269,N_1624,N_1860);
or U2270 (N_2270,N_1310,N_1740);
nand U2271 (N_2271,N_1069,N_1727);
nand U2272 (N_2272,N_1455,N_1847);
xor U2273 (N_2273,N_1900,N_1926);
and U2274 (N_2274,N_1369,N_1912);
xor U2275 (N_2275,N_1207,N_1674);
nor U2276 (N_2276,N_1095,N_1121);
xnor U2277 (N_2277,N_1237,N_1297);
and U2278 (N_2278,N_1819,N_1423);
xor U2279 (N_2279,N_1630,N_1570);
xnor U2280 (N_2280,N_1687,N_1602);
nand U2281 (N_2281,N_1917,N_1732);
or U2282 (N_2282,N_1404,N_1849);
or U2283 (N_2283,N_1092,N_1694);
and U2284 (N_2284,N_1817,N_1625);
or U2285 (N_2285,N_1582,N_1497);
or U2286 (N_2286,N_1902,N_1115);
or U2287 (N_2287,N_1743,N_1262);
nor U2288 (N_2288,N_1032,N_1538);
and U2289 (N_2289,N_1736,N_1835);
xnor U2290 (N_2290,N_1112,N_1966);
xor U2291 (N_2291,N_1741,N_1312);
nand U2292 (N_2292,N_1717,N_1417);
nand U2293 (N_2293,N_1875,N_1869);
xor U2294 (N_2294,N_1245,N_1019);
nor U2295 (N_2295,N_1635,N_1171);
xnor U2296 (N_2296,N_1766,N_1418);
nand U2297 (N_2297,N_1305,N_1937);
or U2298 (N_2298,N_1443,N_1203);
or U2299 (N_2299,N_1253,N_1775);
and U2300 (N_2300,N_1077,N_1947);
nand U2301 (N_2301,N_1520,N_1273);
xnor U2302 (N_2302,N_1352,N_1763);
nor U2303 (N_2303,N_1167,N_1518);
or U2304 (N_2304,N_1856,N_1811);
nand U2305 (N_2305,N_1278,N_1553);
nand U2306 (N_2306,N_1362,N_1774);
or U2307 (N_2307,N_1126,N_1566);
nor U2308 (N_2308,N_1838,N_1194);
xnor U2309 (N_2309,N_1511,N_1474);
or U2310 (N_2310,N_1248,N_1662);
and U2311 (N_2311,N_1945,N_1196);
nand U2312 (N_2312,N_1235,N_1323);
and U2313 (N_2313,N_1380,N_1600);
or U2314 (N_2314,N_1794,N_1061);
nor U2315 (N_2315,N_1494,N_1961);
xor U2316 (N_2316,N_1812,N_1944);
xor U2317 (N_2317,N_1874,N_1594);
xnor U2318 (N_2318,N_1466,N_1969);
and U2319 (N_2319,N_1308,N_1994);
xnor U2320 (N_2320,N_1683,N_1209);
and U2321 (N_2321,N_1742,N_1101);
and U2322 (N_2322,N_1617,N_1985);
nand U2323 (N_2323,N_1764,N_1922);
or U2324 (N_2324,N_1390,N_1881);
or U2325 (N_2325,N_1526,N_1591);
xor U2326 (N_2326,N_1368,N_1344);
xor U2327 (N_2327,N_1872,N_1204);
and U2328 (N_2328,N_1569,N_1295);
and U2329 (N_2329,N_1182,N_1954);
or U2330 (N_2330,N_1723,N_1704);
xor U2331 (N_2331,N_1537,N_1968);
nand U2332 (N_2332,N_1468,N_1531);
nor U2333 (N_2333,N_1281,N_1585);
nor U2334 (N_2334,N_1296,N_1051);
or U2335 (N_2335,N_1991,N_1109);
nor U2336 (N_2336,N_1050,N_1128);
xnor U2337 (N_2337,N_1756,N_1899);
xor U2338 (N_2338,N_1124,N_1202);
nor U2339 (N_2339,N_1877,N_1946);
xnor U2340 (N_2340,N_1512,N_1564);
nor U2341 (N_2341,N_1998,N_1174);
nor U2342 (N_2342,N_1090,N_1657);
and U2343 (N_2343,N_1425,N_1726);
and U2344 (N_2344,N_1089,N_1093);
nand U2345 (N_2345,N_1263,N_1175);
xor U2346 (N_2346,N_1465,N_1643);
nor U2347 (N_2347,N_1367,N_1867);
xor U2348 (N_2348,N_1640,N_1689);
nor U2349 (N_2349,N_1226,N_1598);
nor U2350 (N_2350,N_1546,N_1639);
nor U2351 (N_2351,N_1820,N_1279);
or U2352 (N_2352,N_1676,N_1863);
nor U2353 (N_2353,N_1665,N_1192);
or U2354 (N_2354,N_1022,N_1934);
xnor U2355 (N_2355,N_1078,N_1632);
or U2356 (N_2356,N_1227,N_1350);
nand U2357 (N_2357,N_1543,N_1012);
or U2358 (N_2358,N_1118,N_1454);
xnor U2359 (N_2359,N_1082,N_1463);
or U2360 (N_2360,N_1003,N_1397);
xnor U2361 (N_2361,N_1862,N_1924);
xor U2362 (N_2362,N_1294,N_1324);
nand U2363 (N_2363,N_1280,N_1286);
and U2364 (N_2364,N_1168,N_1343);
and U2365 (N_2365,N_1444,N_1928);
nor U2366 (N_2366,N_1137,N_1478);
nor U2367 (N_2367,N_1224,N_1758);
nor U2368 (N_2368,N_1678,N_1420);
and U2369 (N_2369,N_1735,N_1290);
xor U2370 (N_2370,N_1034,N_1247);
or U2371 (N_2371,N_1490,N_1487);
nor U2372 (N_2372,N_1043,N_1059);
xor U2373 (N_2373,N_1631,N_1376);
or U2374 (N_2374,N_1711,N_1321);
or U2375 (N_2375,N_1098,N_1777);
and U2376 (N_2376,N_1907,N_1522);
nand U2377 (N_2377,N_1931,N_1880);
xnor U2378 (N_2378,N_1299,N_1241);
nand U2379 (N_2379,N_1776,N_1513);
nor U2380 (N_2380,N_1894,N_1130);
nor U2381 (N_2381,N_1229,N_1871);
nor U2382 (N_2382,N_1322,N_1525);
nand U2383 (N_2383,N_1179,N_1085);
and U2384 (N_2384,N_1282,N_1565);
and U2385 (N_2385,N_1334,N_1616);
or U2386 (N_2386,N_1933,N_1769);
or U2387 (N_2387,N_1028,N_1818);
xor U2388 (N_2388,N_1412,N_1948);
or U2389 (N_2389,N_1752,N_1000);
nand U2390 (N_2390,N_1395,N_1383);
nor U2391 (N_2391,N_1445,N_1311);
or U2392 (N_2392,N_1850,N_1789);
or U2393 (N_2393,N_1173,N_1914);
xnor U2394 (N_2394,N_1201,N_1802);
xnor U2395 (N_2395,N_1715,N_1879);
or U2396 (N_2396,N_1066,N_1044);
xor U2397 (N_2397,N_1636,N_1779);
nand U2398 (N_2398,N_1795,N_1483);
xor U2399 (N_2399,N_1302,N_1106);
xnor U2400 (N_2400,N_1612,N_1009);
xor U2401 (N_2401,N_1377,N_1267);
nand U2402 (N_2402,N_1557,N_1895);
xor U2403 (N_2403,N_1503,N_1659);
and U2404 (N_2404,N_1127,N_1033);
and U2405 (N_2405,N_1757,N_1864);
nor U2406 (N_2406,N_1583,N_1219);
xor U2407 (N_2407,N_1940,N_1100);
or U2408 (N_2408,N_1189,N_1386);
nand U2409 (N_2409,N_1541,N_1315);
nor U2410 (N_2410,N_1218,N_1535);
nand U2411 (N_2411,N_1791,N_1187);
and U2412 (N_2412,N_1792,N_1799);
or U2413 (N_2413,N_1524,N_1452);
or U2414 (N_2414,N_1300,N_1669);
and U2415 (N_2415,N_1258,N_1729);
nand U2416 (N_2416,N_1136,N_1941);
and U2417 (N_2417,N_1199,N_1576);
and U2418 (N_2418,N_1349,N_1165);
or U2419 (N_2419,N_1560,N_1852);
xor U2420 (N_2420,N_1645,N_1703);
nand U2421 (N_2421,N_1430,N_1348);
nand U2422 (N_2422,N_1675,N_1056);
and U2423 (N_2423,N_1826,N_1827);
or U2424 (N_2424,N_1163,N_1307);
or U2425 (N_2425,N_1433,N_1064);
and U2426 (N_2426,N_1117,N_1568);
nand U2427 (N_2427,N_1887,N_1153);
and U2428 (N_2428,N_1008,N_1336);
nor U2429 (N_2429,N_1272,N_1317);
or U2430 (N_2430,N_1784,N_1952);
xor U2431 (N_2431,N_1314,N_1626);
or U2432 (N_2432,N_1086,N_1212);
and U2433 (N_2433,N_1120,N_1141);
nand U2434 (N_2434,N_1467,N_1976);
or U2435 (N_2435,N_1439,N_1396);
xor U2436 (N_2436,N_1298,N_1956);
and U2437 (N_2437,N_1691,N_1796);
and U2438 (N_2438,N_1330,N_1898);
xnor U2439 (N_2439,N_1152,N_1584);
xnor U2440 (N_2440,N_1250,N_1805);
and U2441 (N_2441,N_1647,N_1904);
nor U2442 (N_2442,N_1436,N_1870);
nand U2443 (N_2443,N_1829,N_1721);
nand U2444 (N_2444,N_1411,N_1329);
xnor U2445 (N_2445,N_1834,N_1001);
xor U2446 (N_2446,N_1234,N_1197);
nor U2447 (N_2447,N_1048,N_1642);
nor U2448 (N_2448,N_1318,N_1995);
xor U2449 (N_2449,N_1122,N_1110);
nor U2450 (N_2450,N_1765,N_1403);
nor U2451 (N_2451,N_1562,N_1916);
or U2452 (N_2452,N_1822,N_1176);
xnor U2453 (N_2453,N_1105,N_1081);
nor U2454 (N_2454,N_1809,N_1485);
nor U2455 (N_2455,N_1469,N_1129);
xor U2456 (N_2456,N_1586,N_1422);
xor U2457 (N_2457,N_1269,N_1964);
xor U2458 (N_2458,N_1337,N_1702);
nand U2459 (N_2459,N_1670,N_1024);
nand U2460 (N_2460,N_1111,N_1855);
xor U2461 (N_2461,N_1042,N_1161);
xor U2462 (N_2462,N_1951,N_1327);
xnor U2463 (N_2463,N_1987,N_1592);
xor U2464 (N_2464,N_1193,N_1394);
or U2465 (N_2465,N_1575,N_1264);
nand U2466 (N_2466,N_1274,N_1275);
nand U2467 (N_2467,N_1633,N_1493);
and U2468 (N_2468,N_1750,N_1540);
or U2469 (N_2469,N_1751,N_1572);
xnor U2470 (N_2470,N_1426,N_1806);
nor U2471 (N_2471,N_1648,N_1965);
nor U2472 (N_2472,N_1953,N_1270);
or U2473 (N_2473,N_1719,N_1507);
and U2474 (N_2474,N_1154,N_1588);
nand U2475 (N_2475,N_1788,N_1405);
or U2476 (N_2476,N_1778,N_1045);
or U2477 (N_2477,N_1844,N_1627);
or U2478 (N_2478,N_1692,N_1006);
nand U2479 (N_2479,N_1123,N_1038);
xnor U2480 (N_2480,N_1883,N_1149);
or U2481 (N_2481,N_1079,N_1007);
nor U2482 (N_2482,N_1573,N_1548);
or U2483 (N_2483,N_1975,N_1748);
and U2484 (N_2484,N_1375,N_1239);
xor U2485 (N_2485,N_1781,N_1432);
or U2486 (N_2486,N_1773,N_1712);
nand U2487 (N_2487,N_1378,N_1515);
xor U2488 (N_2488,N_1449,N_1915);
xor U2489 (N_2489,N_1151,N_1131);
xor U2490 (N_2490,N_1725,N_1596);
nand U2491 (N_2491,N_1878,N_1373);
or U2492 (N_2492,N_1981,N_1387);
nand U2493 (N_2493,N_1661,N_1988);
and U2494 (N_2494,N_1357,N_1768);
and U2495 (N_2495,N_1923,N_1705);
nor U2496 (N_2496,N_1950,N_1699);
nand U2497 (N_2497,N_1810,N_1385);
and U2498 (N_2498,N_1345,N_1346);
xnor U2499 (N_2499,N_1188,N_1355);
and U2500 (N_2500,N_1795,N_1216);
nor U2501 (N_2501,N_1224,N_1836);
nor U2502 (N_2502,N_1746,N_1949);
nand U2503 (N_2503,N_1772,N_1299);
nand U2504 (N_2504,N_1981,N_1223);
or U2505 (N_2505,N_1284,N_1159);
xnor U2506 (N_2506,N_1160,N_1736);
nand U2507 (N_2507,N_1871,N_1490);
nand U2508 (N_2508,N_1907,N_1840);
or U2509 (N_2509,N_1945,N_1589);
or U2510 (N_2510,N_1094,N_1694);
nor U2511 (N_2511,N_1894,N_1356);
nand U2512 (N_2512,N_1570,N_1647);
and U2513 (N_2513,N_1624,N_1569);
and U2514 (N_2514,N_1312,N_1962);
and U2515 (N_2515,N_1121,N_1186);
nor U2516 (N_2516,N_1428,N_1176);
nor U2517 (N_2517,N_1881,N_1857);
xor U2518 (N_2518,N_1309,N_1204);
and U2519 (N_2519,N_1383,N_1482);
nand U2520 (N_2520,N_1410,N_1724);
nand U2521 (N_2521,N_1505,N_1674);
or U2522 (N_2522,N_1672,N_1845);
nor U2523 (N_2523,N_1601,N_1820);
xnor U2524 (N_2524,N_1887,N_1455);
nand U2525 (N_2525,N_1797,N_1968);
nand U2526 (N_2526,N_1604,N_1285);
nor U2527 (N_2527,N_1149,N_1114);
nand U2528 (N_2528,N_1687,N_1592);
nand U2529 (N_2529,N_1365,N_1612);
xor U2530 (N_2530,N_1698,N_1317);
and U2531 (N_2531,N_1777,N_1155);
and U2532 (N_2532,N_1542,N_1556);
nand U2533 (N_2533,N_1633,N_1347);
or U2534 (N_2534,N_1394,N_1376);
xor U2535 (N_2535,N_1775,N_1938);
or U2536 (N_2536,N_1916,N_1724);
or U2537 (N_2537,N_1966,N_1258);
xnor U2538 (N_2538,N_1505,N_1739);
nand U2539 (N_2539,N_1688,N_1134);
nand U2540 (N_2540,N_1768,N_1721);
nor U2541 (N_2541,N_1305,N_1830);
and U2542 (N_2542,N_1115,N_1600);
and U2543 (N_2543,N_1668,N_1531);
xnor U2544 (N_2544,N_1750,N_1841);
and U2545 (N_2545,N_1389,N_1450);
and U2546 (N_2546,N_1424,N_1781);
and U2547 (N_2547,N_1122,N_1739);
or U2548 (N_2548,N_1814,N_1533);
nand U2549 (N_2549,N_1532,N_1200);
nand U2550 (N_2550,N_1678,N_1744);
xor U2551 (N_2551,N_1083,N_1365);
nand U2552 (N_2552,N_1423,N_1814);
and U2553 (N_2553,N_1736,N_1476);
xor U2554 (N_2554,N_1582,N_1409);
xor U2555 (N_2555,N_1117,N_1650);
or U2556 (N_2556,N_1020,N_1514);
or U2557 (N_2557,N_1758,N_1120);
and U2558 (N_2558,N_1385,N_1639);
nor U2559 (N_2559,N_1839,N_1704);
and U2560 (N_2560,N_1445,N_1016);
xnor U2561 (N_2561,N_1015,N_1147);
nor U2562 (N_2562,N_1928,N_1659);
xor U2563 (N_2563,N_1648,N_1360);
nand U2564 (N_2564,N_1758,N_1321);
nand U2565 (N_2565,N_1428,N_1657);
nand U2566 (N_2566,N_1419,N_1062);
and U2567 (N_2567,N_1522,N_1944);
nand U2568 (N_2568,N_1216,N_1279);
xor U2569 (N_2569,N_1395,N_1220);
and U2570 (N_2570,N_1880,N_1381);
or U2571 (N_2571,N_1056,N_1862);
or U2572 (N_2572,N_1146,N_1919);
nand U2573 (N_2573,N_1225,N_1937);
nand U2574 (N_2574,N_1696,N_1150);
nor U2575 (N_2575,N_1245,N_1064);
nor U2576 (N_2576,N_1753,N_1872);
nand U2577 (N_2577,N_1411,N_1081);
or U2578 (N_2578,N_1454,N_1445);
xor U2579 (N_2579,N_1990,N_1451);
and U2580 (N_2580,N_1175,N_1387);
and U2581 (N_2581,N_1064,N_1519);
and U2582 (N_2582,N_1676,N_1682);
nor U2583 (N_2583,N_1866,N_1064);
and U2584 (N_2584,N_1051,N_1819);
xnor U2585 (N_2585,N_1879,N_1236);
nor U2586 (N_2586,N_1547,N_1657);
or U2587 (N_2587,N_1113,N_1586);
nor U2588 (N_2588,N_1901,N_1103);
or U2589 (N_2589,N_1623,N_1611);
nor U2590 (N_2590,N_1841,N_1380);
nand U2591 (N_2591,N_1131,N_1033);
xnor U2592 (N_2592,N_1030,N_1440);
xor U2593 (N_2593,N_1311,N_1705);
xnor U2594 (N_2594,N_1682,N_1297);
and U2595 (N_2595,N_1873,N_1498);
or U2596 (N_2596,N_1141,N_1420);
nand U2597 (N_2597,N_1983,N_1370);
nand U2598 (N_2598,N_1530,N_1589);
nand U2599 (N_2599,N_1724,N_1958);
nand U2600 (N_2600,N_1058,N_1498);
nand U2601 (N_2601,N_1851,N_1741);
nor U2602 (N_2602,N_1564,N_1134);
or U2603 (N_2603,N_1455,N_1080);
nand U2604 (N_2604,N_1438,N_1394);
and U2605 (N_2605,N_1541,N_1838);
and U2606 (N_2606,N_1961,N_1776);
or U2607 (N_2607,N_1637,N_1709);
xor U2608 (N_2608,N_1288,N_1756);
nor U2609 (N_2609,N_1322,N_1464);
xnor U2610 (N_2610,N_1779,N_1991);
or U2611 (N_2611,N_1211,N_1926);
and U2612 (N_2612,N_1951,N_1744);
xnor U2613 (N_2613,N_1538,N_1519);
nand U2614 (N_2614,N_1362,N_1414);
nand U2615 (N_2615,N_1004,N_1550);
and U2616 (N_2616,N_1092,N_1935);
and U2617 (N_2617,N_1687,N_1897);
nand U2618 (N_2618,N_1862,N_1010);
nand U2619 (N_2619,N_1050,N_1977);
nand U2620 (N_2620,N_1230,N_1029);
xor U2621 (N_2621,N_1037,N_1290);
and U2622 (N_2622,N_1753,N_1268);
nor U2623 (N_2623,N_1367,N_1752);
and U2624 (N_2624,N_1574,N_1512);
xor U2625 (N_2625,N_1237,N_1510);
and U2626 (N_2626,N_1011,N_1177);
or U2627 (N_2627,N_1582,N_1863);
xor U2628 (N_2628,N_1118,N_1434);
or U2629 (N_2629,N_1798,N_1907);
or U2630 (N_2630,N_1145,N_1405);
and U2631 (N_2631,N_1570,N_1948);
or U2632 (N_2632,N_1989,N_1322);
nor U2633 (N_2633,N_1205,N_1744);
nand U2634 (N_2634,N_1577,N_1571);
and U2635 (N_2635,N_1106,N_1342);
nor U2636 (N_2636,N_1675,N_1771);
xor U2637 (N_2637,N_1790,N_1243);
and U2638 (N_2638,N_1131,N_1436);
xnor U2639 (N_2639,N_1093,N_1203);
nor U2640 (N_2640,N_1944,N_1765);
nor U2641 (N_2641,N_1847,N_1005);
xnor U2642 (N_2642,N_1515,N_1808);
xnor U2643 (N_2643,N_1180,N_1236);
nand U2644 (N_2644,N_1837,N_1287);
nand U2645 (N_2645,N_1067,N_1710);
nor U2646 (N_2646,N_1496,N_1354);
and U2647 (N_2647,N_1933,N_1242);
and U2648 (N_2648,N_1694,N_1838);
xnor U2649 (N_2649,N_1912,N_1091);
nor U2650 (N_2650,N_1643,N_1281);
xor U2651 (N_2651,N_1165,N_1226);
nor U2652 (N_2652,N_1856,N_1880);
or U2653 (N_2653,N_1510,N_1231);
and U2654 (N_2654,N_1716,N_1755);
nand U2655 (N_2655,N_1620,N_1594);
xnor U2656 (N_2656,N_1209,N_1978);
nor U2657 (N_2657,N_1761,N_1943);
nor U2658 (N_2658,N_1102,N_1626);
nand U2659 (N_2659,N_1695,N_1947);
xnor U2660 (N_2660,N_1938,N_1028);
and U2661 (N_2661,N_1204,N_1593);
xor U2662 (N_2662,N_1087,N_1900);
nor U2663 (N_2663,N_1416,N_1487);
nor U2664 (N_2664,N_1734,N_1635);
xor U2665 (N_2665,N_1828,N_1686);
nand U2666 (N_2666,N_1334,N_1993);
or U2667 (N_2667,N_1134,N_1913);
or U2668 (N_2668,N_1414,N_1111);
nand U2669 (N_2669,N_1727,N_1239);
nor U2670 (N_2670,N_1637,N_1374);
nand U2671 (N_2671,N_1606,N_1995);
nand U2672 (N_2672,N_1701,N_1806);
nor U2673 (N_2673,N_1247,N_1191);
xor U2674 (N_2674,N_1577,N_1999);
nor U2675 (N_2675,N_1409,N_1623);
or U2676 (N_2676,N_1771,N_1932);
xnor U2677 (N_2677,N_1052,N_1563);
nand U2678 (N_2678,N_1301,N_1541);
nor U2679 (N_2679,N_1260,N_1390);
nand U2680 (N_2680,N_1630,N_1018);
and U2681 (N_2681,N_1352,N_1040);
xor U2682 (N_2682,N_1047,N_1368);
nand U2683 (N_2683,N_1383,N_1945);
and U2684 (N_2684,N_1871,N_1590);
nand U2685 (N_2685,N_1371,N_1314);
nor U2686 (N_2686,N_1264,N_1478);
xor U2687 (N_2687,N_1305,N_1884);
and U2688 (N_2688,N_1746,N_1015);
nand U2689 (N_2689,N_1998,N_1270);
or U2690 (N_2690,N_1017,N_1393);
nand U2691 (N_2691,N_1378,N_1933);
or U2692 (N_2692,N_1671,N_1235);
nand U2693 (N_2693,N_1655,N_1469);
nand U2694 (N_2694,N_1232,N_1824);
nand U2695 (N_2695,N_1724,N_1698);
xor U2696 (N_2696,N_1132,N_1719);
nand U2697 (N_2697,N_1646,N_1226);
nand U2698 (N_2698,N_1404,N_1244);
or U2699 (N_2699,N_1784,N_1648);
nand U2700 (N_2700,N_1473,N_1022);
nor U2701 (N_2701,N_1896,N_1836);
nor U2702 (N_2702,N_1432,N_1137);
nand U2703 (N_2703,N_1294,N_1746);
nand U2704 (N_2704,N_1279,N_1916);
or U2705 (N_2705,N_1721,N_1976);
or U2706 (N_2706,N_1767,N_1982);
and U2707 (N_2707,N_1143,N_1627);
or U2708 (N_2708,N_1493,N_1800);
or U2709 (N_2709,N_1758,N_1154);
nor U2710 (N_2710,N_1193,N_1621);
nor U2711 (N_2711,N_1519,N_1918);
and U2712 (N_2712,N_1764,N_1399);
nand U2713 (N_2713,N_1226,N_1788);
xnor U2714 (N_2714,N_1164,N_1101);
nor U2715 (N_2715,N_1601,N_1459);
or U2716 (N_2716,N_1089,N_1347);
and U2717 (N_2717,N_1949,N_1296);
nand U2718 (N_2718,N_1085,N_1013);
xor U2719 (N_2719,N_1982,N_1023);
xnor U2720 (N_2720,N_1129,N_1758);
and U2721 (N_2721,N_1876,N_1135);
nand U2722 (N_2722,N_1056,N_1211);
or U2723 (N_2723,N_1719,N_1743);
nor U2724 (N_2724,N_1892,N_1757);
nand U2725 (N_2725,N_1537,N_1153);
or U2726 (N_2726,N_1297,N_1238);
or U2727 (N_2727,N_1434,N_1834);
or U2728 (N_2728,N_1902,N_1338);
or U2729 (N_2729,N_1453,N_1564);
nor U2730 (N_2730,N_1972,N_1773);
or U2731 (N_2731,N_1355,N_1168);
and U2732 (N_2732,N_1612,N_1520);
or U2733 (N_2733,N_1701,N_1035);
nor U2734 (N_2734,N_1609,N_1101);
or U2735 (N_2735,N_1124,N_1463);
xnor U2736 (N_2736,N_1925,N_1944);
nor U2737 (N_2737,N_1094,N_1027);
or U2738 (N_2738,N_1924,N_1925);
and U2739 (N_2739,N_1548,N_1624);
and U2740 (N_2740,N_1459,N_1819);
nand U2741 (N_2741,N_1758,N_1223);
or U2742 (N_2742,N_1540,N_1475);
nand U2743 (N_2743,N_1686,N_1207);
or U2744 (N_2744,N_1303,N_1029);
nor U2745 (N_2745,N_1881,N_1380);
and U2746 (N_2746,N_1673,N_1761);
xor U2747 (N_2747,N_1143,N_1357);
nand U2748 (N_2748,N_1354,N_1925);
and U2749 (N_2749,N_1141,N_1574);
nand U2750 (N_2750,N_1873,N_1380);
or U2751 (N_2751,N_1565,N_1495);
and U2752 (N_2752,N_1078,N_1267);
xor U2753 (N_2753,N_1177,N_1848);
xnor U2754 (N_2754,N_1107,N_1204);
nand U2755 (N_2755,N_1542,N_1777);
xnor U2756 (N_2756,N_1350,N_1674);
or U2757 (N_2757,N_1098,N_1352);
nand U2758 (N_2758,N_1222,N_1627);
xor U2759 (N_2759,N_1827,N_1039);
nand U2760 (N_2760,N_1763,N_1181);
nand U2761 (N_2761,N_1207,N_1427);
or U2762 (N_2762,N_1692,N_1548);
or U2763 (N_2763,N_1020,N_1957);
nand U2764 (N_2764,N_1466,N_1220);
nor U2765 (N_2765,N_1218,N_1930);
and U2766 (N_2766,N_1161,N_1239);
nor U2767 (N_2767,N_1297,N_1458);
or U2768 (N_2768,N_1864,N_1341);
nor U2769 (N_2769,N_1461,N_1835);
and U2770 (N_2770,N_1301,N_1402);
or U2771 (N_2771,N_1632,N_1017);
or U2772 (N_2772,N_1812,N_1248);
or U2773 (N_2773,N_1515,N_1256);
nor U2774 (N_2774,N_1794,N_1445);
and U2775 (N_2775,N_1752,N_1982);
nor U2776 (N_2776,N_1659,N_1766);
and U2777 (N_2777,N_1965,N_1089);
nor U2778 (N_2778,N_1971,N_1822);
or U2779 (N_2779,N_1029,N_1825);
xnor U2780 (N_2780,N_1356,N_1449);
nand U2781 (N_2781,N_1408,N_1732);
and U2782 (N_2782,N_1569,N_1944);
xnor U2783 (N_2783,N_1579,N_1333);
nor U2784 (N_2784,N_1157,N_1821);
or U2785 (N_2785,N_1462,N_1250);
xnor U2786 (N_2786,N_1593,N_1675);
xnor U2787 (N_2787,N_1750,N_1431);
nor U2788 (N_2788,N_1089,N_1286);
nor U2789 (N_2789,N_1266,N_1753);
nor U2790 (N_2790,N_1685,N_1198);
nor U2791 (N_2791,N_1189,N_1013);
nor U2792 (N_2792,N_1480,N_1908);
nand U2793 (N_2793,N_1863,N_1790);
nand U2794 (N_2794,N_1300,N_1397);
xor U2795 (N_2795,N_1422,N_1143);
nand U2796 (N_2796,N_1692,N_1866);
or U2797 (N_2797,N_1578,N_1425);
xor U2798 (N_2798,N_1035,N_1384);
xor U2799 (N_2799,N_1973,N_1349);
nand U2800 (N_2800,N_1843,N_1520);
nand U2801 (N_2801,N_1410,N_1149);
xor U2802 (N_2802,N_1746,N_1602);
and U2803 (N_2803,N_1277,N_1099);
and U2804 (N_2804,N_1758,N_1623);
or U2805 (N_2805,N_1307,N_1528);
or U2806 (N_2806,N_1981,N_1379);
and U2807 (N_2807,N_1795,N_1993);
xor U2808 (N_2808,N_1431,N_1797);
nand U2809 (N_2809,N_1005,N_1925);
or U2810 (N_2810,N_1463,N_1737);
xor U2811 (N_2811,N_1902,N_1834);
nand U2812 (N_2812,N_1164,N_1228);
nor U2813 (N_2813,N_1967,N_1969);
or U2814 (N_2814,N_1906,N_1974);
nor U2815 (N_2815,N_1305,N_1514);
or U2816 (N_2816,N_1265,N_1611);
or U2817 (N_2817,N_1791,N_1893);
or U2818 (N_2818,N_1534,N_1916);
xnor U2819 (N_2819,N_1078,N_1826);
xor U2820 (N_2820,N_1451,N_1211);
nor U2821 (N_2821,N_1747,N_1064);
nand U2822 (N_2822,N_1967,N_1398);
nand U2823 (N_2823,N_1819,N_1458);
nor U2824 (N_2824,N_1562,N_1302);
xor U2825 (N_2825,N_1719,N_1143);
nor U2826 (N_2826,N_1629,N_1308);
or U2827 (N_2827,N_1885,N_1389);
nor U2828 (N_2828,N_1188,N_1965);
nand U2829 (N_2829,N_1030,N_1899);
nor U2830 (N_2830,N_1583,N_1663);
and U2831 (N_2831,N_1236,N_1100);
nor U2832 (N_2832,N_1035,N_1607);
xor U2833 (N_2833,N_1926,N_1905);
and U2834 (N_2834,N_1670,N_1623);
xnor U2835 (N_2835,N_1403,N_1472);
or U2836 (N_2836,N_1962,N_1201);
nor U2837 (N_2837,N_1893,N_1335);
and U2838 (N_2838,N_1472,N_1134);
xor U2839 (N_2839,N_1976,N_1079);
xor U2840 (N_2840,N_1196,N_1963);
nor U2841 (N_2841,N_1146,N_1581);
or U2842 (N_2842,N_1392,N_1573);
or U2843 (N_2843,N_1324,N_1472);
xnor U2844 (N_2844,N_1896,N_1974);
or U2845 (N_2845,N_1258,N_1424);
nor U2846 (N_2846,N_1774,N_1200);
nor U2847 (N_2847,N_1578,N_1843);
nor U2848 (N_2848,N_1871,N_1309);
nor U2849 (N_2849,N_1825,N_1767);
xnor U2850 (N_2850,N_1705,N_1406);
and U2851 (N_2851,N_1298,N_1924);
or U2852 (N_2852,N_1805,N_1443);
or U2853 (N_2853,N_1664,N_1367);
nand U2854 (N_2854,N_1408,N_1823);
nand U2855 (N_2855,N_1362,N_1829);
or U2856 (N_2856,N_1881,N_1255);
or U2857 (N_2857,N_1958,N_1723);
nand U2858 (N_2858,N_1949,N_1928);
or U2859 (N_2859,N_1320,N_1263);
or U2860 (N_2860,N_1895,N_1147);
nor U2861 (N_2861,N_1378,N_1424);
nand U2862 (N_2862,N_1388,N_1393);
xor U2863 (N_2863,N_1668,N_1728);
xor U2864 (N_2864,N_1265,N_1903);
or U2865 (N_2865,N_1272,N_1391);
and U2866 (N_2866,N_1601,N_1035);
xnor U2867 (N_2867,N_1152,N_1817);
and U2868 (N_2868,N_1746,N_1946);
nand U2869 (N_2869,N_1046,N_1381);
nand U2870 (N_2870,N_1211,N_1537);
or U2871 (N_2871,N_1494,N_1876);
xnor U2872 (N_2872,N_1826,N_1407);
and U2873 (N_2873,N_1536,N_1977);
xnor U2874 (N_2874,N_1107,N_1441);
or U2875 (N_2875,N_1237,N_1978);
and U2876 (N_2876,N_1439,N_1212);
and U2877 (N_2877,N_1237,N_1229);
or U2878 (N_2878,N_1710,N_1632);
nand U2879 (N_2879,N_1617,N_1594);
and U2880 (N_2880,N_1455,N_1138);
nor U2881 (N_2881,N_1046,N_1751);
or U2882 (N_2882,N_1874,N_1506);
nor U2883 (N_2883,N_1259,N_1927);
nand U2884 (N_2884,N_1073,N_1935);
or U2885 (N_2885,N_1987,N_1243);
xor U2886 (N_2886,N_1100,N_1858);
nand U2887 (N_2887,N_1241,N_1746);
and U2888 (N_2888,N_1746,N_1202);
and U2889 (N_2889,N_1906,N_1007);
and U2890 (N_2890,N_1079,N_1994);
nand U2891 (N_2891,N_1837,N_1529);
nand U2892 (N_2892,N_1698,N_1247);
nand U2893 (N_2893,N_1135,N_1405);
xnor U2894 (N_2894,N_1795,N_1298);
nor U2895 (N_2895,N_1806,N_1049);
or U2896 (N_2896,N_1743,N_1687);
nor U2897 (N_2897,N_1892,N_1554);
nand U2898 (N_2898,N_1124,N_1274);
nand U2899 (N_2899,N_1495,N_1742);
and U2900 (N_2900,N_1031,N_1988);
nand U2901 (N_2901,N_1579,N_1446);
xnor U2902 (N_2902,N_1408,N_1020);
xor U2903 (N_2903,N_1797,N_1212);
xnor U2904 (N_2904,N_1351,N_1053);
xor U2905 (N_2905,N_1255,N_1447);
nor U2906 (N_2906,N_1816,N_1560);
xor U2907 (N_2907,N_1284,N_1859);
nor U2908 (N_2908,N_1801,N_1672);
nand U2909 (N_2909,N_1669,N_1751);
nor U2910 (N_2910,N_1186,N_1464);
xnor U2911 (N_2911,N_1641,N_1020);
nand U2912 (N_2912,N_1016,N_1108);
or U2913 (N_2913,N_1225,N_1091);
nor U2914 (N_2914,N_1085,N_1143);
and U2915 (N_2915,N_1626,N_1601);
or U2916 (N_2916,N_1310,N_1231);
and U2917 (N_2917,N_1609,N_1858);
xnor U2918 (N_2918,N_1716,N_1547);
or U2919 (N_2919,N_1171,N_1859);
nor U2920 (N_2920,N_1108,N_1555);
nor U2921 (N_2921,N_1954,N_1607);
or U2922 (N_2922,N_1275,N_1523);
and U2923 (N_2923,N_1729,N_1597);
nor U2924 (N_2924,N_1250,N_1763);
and U2925 (N_2925,N_1772,N_1007);
nor U2926 (N_2926,N_1464,N_1019);
nand U2927 (N_2927,N_1759,N_1527);
nand U2928 (N_2928,N_1055,N_1081);
and U2929 (N_2929,N_1249,N_1696);
nor U2930 (N_2930,N_1460,N_1793);
xnor U2931 (N_2931,N_1726,N_1780);
or U2932 (N_2932,N_1297,N_1356);
xor U2933 (N_2933,N_1739,N_1006);
nand U2934 (N_2934,N_1198,N_1522);
xnor U2935 (N_2935,N_1013,N_1111);
nor U2936 (N_2936,N_1732,N_1715);
nor U2937 (N_2937,N_1043,N_1081);
xnor U2938 (N_2938,N_1093,N_1359);
nand U2939 (N_2939,N_1378,N_1770);
xnor U2940 (N_2940,N_1587,N_1733);
xnor U2941 (N_2941,N_1721,N_1036);
nor U2942 (N_2942,N_1154,N_1670);
nand U2943 (N_2943,N_1438,N_1164);
nand U2944 (N_2944,N_1122,N_1283);
and U2945 (N_2945,N_1825,N_1940);
and U2946 (N_2946,N_1796,N_1826);
nor U2947 (N_2947,N_1696,N_1489);
xor U2948 (N_2948,N_1003,N_1139);
nand U2949 (N_2949,N_1315,N_1241);
xnor U2950 (N_2950,N_1161,N_1177);
nor U2951 (N_2951,N_1705,N_1398);
xnor U2952 (N_2952,N_1671,N_1285);
nor U2953 (N_2953,N_1320,N_1749);
and U2954 (N_2954,N_1843,N_1785);
nor U2955 (N_2955,N_1531,N_1099);
nor U2956 (N_2956,N_1913,N_1170);
xor U2957 (N_2957,N_1024,N_1603);
and U2958 (N_2958,N_1497,N_1638);
or U2959 (N_2959,N_1529,N_1324);
or U2960 (N_2960,N_1744,N_1180);
xnor U2961 (N_2961,N_1564,N_1488);
xor U2962 (N_2962,N_1479,N_1104);
nor U2963 (N_2963,N_1874,N_1338);
xnor U2964 (N_2964,N_1884,N_1387);
nor U2965 (N_2965,N_1482,N_1897);
or U2966 (N_2966,N_1852,N_1467);
nor U2967 (N_2967,N_1544,N_1361);
xnor U2968 (N_2968,N_1707,N_1139);
or U2969 (N_2969,N_1339,N_1560);
and U2970 (N_2970,N_1890,N_1084);
xor U2971 (N_2971,N_1062,N_1164);
xnor U2972 (N_2972,N_1071,N_1970);
nand U2973 (N_2973,N_1655,N_1219);
nor U2974 (N_2974,N_1832,N_1326);
and U2975 (N_2975,N_1311,N_1179);
xor U2976 (N_2976,N_1280,N_1705);
nor U2977 (N_2977,N_1608,N_1906);
xnor U2978 (N_2978,N_1552,N_1278);
and U2979 (N_2979,N_1403,N_1493);
nand U2980 (N_2980,N_1639,N_1967);
and U2981 (N_2981,N_1819,N_1560);
and U2982 (N_2982,N_1191,N_1839);
and U2983 (N_2983,N_1149,N_1353);
and U2984 (N_2984,N_1297,N_1057);
xor U2985 (N_2985,N_1742,N_1114);
and U2986 (N_2986,N_1421,N_1131);
and U2987 (N_2987,N_1326,N_1243);
and U2988 (N_2988,N_1111,N_1316);
nand U2989 (N_2989,N_1220,N_1131);
or U2990 (N_2990,N_1043,N_1945);
and U2991 (N_2991,N_1910,N_1023);
nand U2992 (N_2992,N_1940,N_1801);
xnor U2993 (N_2993,N_1938,N_1657);
xnor U2994 (N_2994,N_1836,N_1079);
nand U2995 (N_2995,N_1878,N_1059);
nand U2996 (N_2996,N_1255,N_1503);
nand U2997 (N_2997,N_1951,N_1477);
and U2998 (N_2998,N_1551,N_1736);
nor U2999 (N_2999,N_1915,N_1370);
xor U3000 (N_3000,N_2914,N_2428);
nand U3001 (N_3001,N_2520,N_2563);
nand U3002 (N_3002,N_2489,N_2098);
nand U3003 (N_3003,N_2132,N_2610);
and U3004 (N_3004,N_2230,N_2949);
nand U3005 (N_3005,N_2095,N_2123);
xor U3006 (N_3006,N_2897,N_2993);
nor U3007 (N_3007,N_2577,N_2127);
and U3008 (N_3008,N_2517,N_2820);
and U3009 (N_3009,N_2937,N_2814);
nand U3010 (N_3010,N_2131,N_2602);
nand U3011 (N_3011,N_2427,N_2142);
nand U3012 (N_3012,N_2621,N_2877);
nor U3013 (N_3013,N_2351,N_2768);
nor U3014 (N_3014,N_2863,N_2958);
nand U3015 (N_3015,N_2025,N_2928);
xor U3016 (N_3016,N_2411,N_2499);
nand U3017 (N_3017,N_2306,N_2181);
xnor U3018 (N_3018,N_2390,N_2216);
xor U3019 (N_3019,N_2367,N_2043);
xnor U3020 (N_3020,N_2195,N_2940);
nand U3021 (N_3021,N_2109,N_2959);
or U3022 (N_3022,N_2705,N_2175);
or U3023 (N_3023,N_2723,N_2388);
or U3024 (N_3024,N_2720,N_2589);
or U3025 (N_3025,N_2373,N_2270);
xnor U3026 (N_3026,N_2240,N_2442);
nand U3027 (N_3027,N_2544,N_2509);
nor U3028 (N_3028,N_2515,N_2709);
or U3029 (N_3029,N_2700,N_2627);
or U3030 (N_3030,N_2867,N_2683);
and U3031 (N_3031,N_2458,N_2795);
and U3032 (N_3032,N_2218,N_2561);
or U3033 (N_3033,N_2271,N_2360);
and U3034 (N_3034,N_2116,N_2465);
and U3035 (N_3035,N_2706,N_2732);
xor U3036 (N_3036,N_2920,N_2617);
nand U3037 (N_3037,N_2840,N_2026);
and U3038 (N_3038,N_2283,N_2259);
nand U3039 (N_3039,N_2649,N_2243);
xor U3040 (N_3040,N_2102,N_2145);
or U3041 (N_3041,N_2072,N_2611);
nor U3042 (N_3042,N_2997,N_2954);
nand U3043 (N_3043,N_2524,N_2299);
xor U3044 (N_3044,N_2454,N_2895);
xor U3045 (N_3045,N_2153,N_2381);
nand U3046 (N_3046,N_2235,N_2823);
nor U3047 (N_3047,N_2595,N_2981);
xnor U3048 (N_3048,N_2481,N_2199);
nand U3049 (N_3049,N_2125,N_2069);
nor U3050 (N_3050,N_2518,N_2001);
or U3051 (N_3051,N_2212,N_2872);
nand U3052 (N_3052,N_2943,N_2900);
and U3053 (N_3053,N_2809,N_2088);
xor U3054 (N_3054,N_2267,N_2780);
or U3055 (N_3055,N_2850,N_2298);
or U3056 (N_3056,N_2277,N_2207);
and U3057 (N_3057,N_2213,N_2331);
nor U3058 (N_3058,N_2639,N_2164);
nor U3059 (N_3059,N_2944,N_2317);
or U3060 (N_3060,N_2321,N_2057);
and U3061 (N_3061,N_2533,N_2078);
xor U3062 (N_3062,N_2491,N_2531);
xor U3063 (N_3063,N_2614,N_2136);
or U3064 (N_3064,N_2676,N_2716);
nand U3065 (N_3065,N_2340,N_2906);
nor U3066 (N_3066,N_2336,N_2786);
xor U3067 (N_3067,N_2041,N_2403);
or U3068 (N_3068,N_2358,N_2324);
and U3069 (N_3069,N_2335,N_2392);
xnor U3070 (N_3070,N_2543,N_2334);
and U3071 (N_3071,N_2387,N_2528);
or U3072 (N_3072,N_2788,N_2751);
nor U3073 (N_3073,N_2580,N_2440);
nor U3074 (N_3074,N_2038,N_2694);
and U3075 (N_3075,N_2276,N_2757);
xnor U3076 (N_3076,N_2049,N_2300);
nor U3077 (N_3077,N_2368,N_2138);
or U3078 (N_3078,N_2452,N_2607);
xor U3079 (N_3079,N_2082,N_2279);
nor U3080 (N_3080,N_2684,N_2460);
nor U3081 (N_3081,N_2477,N_2268);
nor U3082 (N_3082,N_2034,N_2327);
nor U3083 (N_3083,N_2285,N_2999);
nand U3084 (N_3084,N_2922,N_2737);
nand U3085 (N_3085,N_2409,N_2464);
nand U3086 (N_3086,N_2902,N_2446);
and U3087 (N_3087,N_2762,N_2573);
xnor U3088 (N_3088,N_2891,N_2957);
nor U3089 (N_3089,N_2092,N_2721);
or U3090 (N_3090,N_2763,N_2730);
or U3091 (N_3091,N_2115,N_2157);
xnor U3092 (N_3092,N_2070,N_2713);
nand U3093 (N_3093,N_2979,N_2414);
nor U3094 (N_3094,N_2538,N_2167);
or U3095 (N_3095,N_2842,N_2469);
nand U3096 (N_3096,N_2502,N_2576);
and U3097 (N_3097,N_2590,N_2323);
nand U3098 (N_3098,N_2624,N_2238);
and U3099 (N_3099,N_2861,N_2309);
and U3100 (N_3100,N_2080,N_2698);
or U3101 (N_3101,N_2813,N_2779);
nand U3102 (N_3102,N_2598,N_2745);
or U3103 (N_3103,N_2746,N_2626);
nor U3104 (N_3104,N_2508,N_2227);
nand U3105 (N_3105,N_2063,N_2522);
and U3106 (N_3106,N_2680,N_2091);
and U3107 (N_3107,N_2951,N_2586);
nand U3108 (N_3108,N_2056,N_2475);
xnor U3109 (N_3109,N_2945,N_2927);
or U3110 (N_3110,N_2790,N_2090);
or U3111 (N_3111,N_2512,N_2597);
xor U3112 (N_3112,N_2688,N_2225);
nand U3113 (N_3113,N_2148,N_2249);
nor U3114 (N_3114,N_2364,N_2756);
nor U3115 (N_3115,N_2913,N_2420);
and U3116 (N_3116,N_2455,N_2006);
nor U3117 (N_3117,N_2844,N_2206);
or U3118 (N_3118,N_2896,N_2162);
and U3119 (N_3119,N_2176,N_2657);
and U3120 (N_3120,N_2966,N_2605);
nor U3121 (N_3121,N_2124,N_2868);
nand U3122 (N_3122,N_2521,N_2578);
xor U3123 (N_3123,N_2883,N_2690);
xor U3124 (N_3124,N_2401,N_2969);
nor U3125 (N_3125,N_2618,N_2169);
xor U3126 (N_3126,N_2992,N_2998);
and U3127 (N_3127,N_2677,N_2702);
or U3128 (N_3128,N_2479,N_2282);
nor U3129 (N_3129,N_2988,N_2474);
xor U3130 (N_3130,N_2357,N_2847);
nand U3131 (N_3131,N_2168,N_2425);
nand U3132 (N_3132,N_2485,N_2386);
xor U3133 (N_3133,N_2066,N_2105);
or U3134 (N_3134,N_2826,N_2224);
and U3135 (N_3135,N_2260,N_2806);
and U3136 (N_3136,N_2669,N_2223);
or U3137 (N_3137,N_2322,N_2412);
and U3138 (N_3138,N_2472,N_2871);
or U3139 (N_3139,N_2740,N_2585);
nand U3140 (N_3140,N_2160,N_2430);
xor U3141 (N_3141,N_2137,N_2210);
xnor U3142 (N_3142,N_2699,N_2421);
nand U3143 (N_3143,N_2854,N_2909);
and U3144 (N_3144,N_2894,N_2591);
nor U3145 (N_3145,N_2916,N_2356);
xor U3146 (N_3146,N_2444,N_2004);
xor U3147 (N_3147,N_2575,N_2165);
nor U3148 (N_3148,N_2217,N_2667);
xnor U3149 (N_3149,N_2985,N_2478);
or U3150 (N_3150,N_2486,N_2725);
nor U3151 (N_3151,N_2028,N_2560);
and U3152 (N_3152,N_2365,N_2439);
xnor U3153 (N_3153,N_2384,N_2231);
nand U3154 (N_3154,N_2693,N_2250);
nor U3155 (N_3155,N_2892,N_2808);
or U3156 (N_3156,N_2059,N_2058);
nor U3157 (N_3157,N_2641,N_2042);
xnor U3158 (N_3158,N_2845,N_2076);
xnor U3159 (N_3159,N_2822,N_2687);
nor U3160 (N_3160,N_2426,N_2048);
nand U3161 (N_3161,N_2177,N_2121);
or U3162 (N_3162,N_2704,N_2400);
xnor U3163 (N_3163,N_2291,N_2111);
or U3164 (N_3164,N_2143,N_2545);
xnor U3165 (N_3165,N_2749,N_2396);
or U3166 (N_3166,N_2956,N_2960);
or U3167 (N_3167,N_2950,N_2819);
and U3168 (N_3168,N_2482,N_2150);
and U3169 (N_3169,N_2829,N_2461);
nor U3170 (N_3170,N_2976,N_2931);
xor U3171 (N_3171,N_2510,N_2539);
xnor U3172 (N_3172,N_2601,N_2050);
nor U3173 (N_3173,N_2438,N_2659);
and U3174 (N_3174,N_2752,N_2413);
nand U3175 (N_3175,N_2803,N_2064);
xor U3176 (N_3176,N_2933,N_2226);
nand U3177 (N_3177,N_2326,N_2848);
nor U3178 (N_3178,N_2394,N_2180);
nand U3179 (N_3179,N_2009,N_2583);
xor U3180 (N_3180,N_2010,N_2158);
xor U3181 (N_3181,N_2068,N_2441);
and U3182 (N_3182,N_2798,N_2110);
xor U3183 (N_3183,N_2404,N_2348);
or U3184 (N_3184,N_2592,N_2075);
and U3185 (N_3185,N_2535,N_2172);
nor U3186 (N_3186,N_2194,N_2263);
or U3187 (N_3187,N_2293,N_2112);
xor U3188 (N_3188,N_2670,N_2566);
nand U3189 (N_3189,N_2380,N_2946);
and U3190 (N_3190,N_2003,N_2410);
nor U3191 (N_3191,N_2715,N_2081);
and U3192 (N_3192,N_2492,N_2565);
xnor U3193 (N_3193,N_2242,N_2214);
xor U3194 (N_3194,N_2273,N_2769);
or U3195 (N_3195,N_2371,N_2343);
nand U3196 (N_3196,N_2262,N_2569);
and U3197 (N_3197,N_2087,N_2362);
or U3198 (N_3198,N_2532,N_2604);
and U3199 (N_3199,N_2910,N_2040);
or U3200 (N_3200,N_2506,N_2564);
nand U3201 (N_3201,N_2741,N_2289);
xor U3202 (N_3202,N_2328,N_2338);
nand U3203 (N_3203,N_2977,N_2220);
and U3204 (N_3204,N_2366,N_2661);
and U3205 (N_3205,N_2612,N_2278);
nor U3206 (N_3206,N_2800,N_2727);
nand U3207 (N_3207,N_2930,N_2921);
or U3208 (N_3208,N_2529,N_2128);
nor U3209 (N_3209,N_2376,N_2556);
nor U3210 (N_3210,N_2007,N_2253);
xnor U3211 (N_3211,N_2385,N_2325);
nor U3212 (N_3212,N_2834,N_2496);
nor U3213 (N_3213,N_2567,N_2651);
xor U3214 (N_3214,N_2903,N_2682);
and U3215 (N_3215,N_2630,N_2961);
xnor U3216 (N_3216,N_2793,N_2189);
nand U3217 (N_3217,N_2039,N_2196);
xnor U3218 (N_3218,N_2773,N_2789);
xor U3219 (N_3219,N_2830,N_2572);
xor U3220 (N_3220,N_2085,N_2729);
nand U3221 (N_3221,N_2159,N_2519);
nand U3222 (N_3222,N_2369,N_2209);
or U3223 (N_3223,N_2971,N_2615);
nand U3224 (N_3224,N_2352,N_2691);
nand U3225 (N_3225,N_2215,N_2000);
xor U3226 (N_3226,N_2349,N_2660);
and U3227 (N_3227,N_2642,N_2857);
and U3228 (N_3228,N_2925,N_2514);
or U3229 (N_3229,N_2051,N_2097);
or U3230 (N_3230,N_2986,N_2760);
xor U3231 (N_3231,N_2837,N_2962);
xnor U3232 (N_3232,N_2024,N_2938);
xor U3233 (N_3233,N_2133,N_2712);
or U3234 (N_3234,N_2391,N_2758);
or U3235 (N_3235,N_2622,N_2451);
and U3236 (N_3236,N_2689,N_2707);
or U3237 (N_3237,N_2989,N_2272);
nand U3238 (N_3238,N_2785,N_2089);
xnor U3239 (N_3239,N_2077,N_2620);
nand U3240 (N_3240,N_2174,N_2146);
xnor U3241 (N_3241,N_2681,N_2314);
xor U3242 (N_3242,N_2726,N_2295);
xor U3243 (N_3243,N_2201,N_2232);
nor U3244 (N_3244,N_2536,N_2023);
or U3245 (N_3245,N_2054,N_2449);
nor U3246 (N_3246,N_2653,N_2636);
and U3247 (N_3247,N_2257,N_2770);
nor U3248 (N_3248,N_2134,N_2866);
and U3249 (N_3249,N_2841,N_2915);
and U3250 (N_3250,N_2672,N_2632);
nor U3251 (N_3251,N_2487,N_2332);
nand U3252 (N_3252,N_2233,N_2155);
xnor U3253 (N_3253,N_2771,N_2596);
nand U3254 (N_3254,N_2523,N_2047);
nor U3255 (N_3255,N_2178,N_2675);
and U3256 (N_3256,N_2679,N_2484);
or U3257 (N_3257,N_2637,N_2315);
and U3258 (N_3258,N_2045,N_2188);
nand U3259 (N_3259,N_2724,N_2608);
nor U3260 (N_3260,N_2129,N_2970);
nand U3261 (N_3261,N_2084,N_2852);
xnor U3262 (N_3262,N_2965,N_2935);
or U3263 (N_3263,N_2173,N_2817);
and U3264 (N_3264,N_2831,N_2313);
nor U3265 (N_3265,N_2382,N_2031);
or U3266 (N_3266,N_2305,N_2337);
nand U3267 (N_3267,N_2821,N_2296);
and U3268 (N_3268,N_2383,N_2436);
or U3269 (N_3269,N_2053,N_2899);
nand U3270 (N_3270,N_2372,N_2011);
nor U3271 (N_3271,N_2422,N_2511);
xnor U3272 (N_3272,N_2244,N_2967);
and U3273 (N_3273,N_2046,N_2154);
nor U3274 (N_3274,N_2149,N_2804);
and U3275 (N_3275,N_2911,N_2581);
xnor U3276 (N_3276,N_2122,N_2754);
nor U3277 (N_3277,N_2103,N_2942);
xnor U3278 (N_3278,N_2530,N_2333);
xnor U3279 (N_3279,N_2810,N_2002);
xnor U3280 (N_3280,N_2584,N_2666);
and U3281 (N_3281,N_2701,N_2640);
nand U3282 (N_3282,N_2980,N_2397);
nor U3283 (N_3283,N_2638,N_2494);
nor U3284 (N_3284,N_2650,N_2893);
or U3285 (N_3285,N_2166,N_2812);
xor U3286 (N_3286,N_2185,N_2504);
or U3287 (N_3287,N_2493,N_2488);
or U3288 (N_3288,N_2836,N_2549);
nor U3289 (N_3289,N_2934,N_2568);
and U3290 (N_3290,N_2377,N_2443);
nand U3291 (N_3291,N_2792,N_2929);
nor U3292 (N_3292,N_2582,N_2885);
or U3293 (N_3293,N_2525,N_2113);
nor U3294 (N_3294,N_2062,N_2312);
xnor U3295 (N_3295,N_2643,N_2497);
and U3296 (N_3296,N_2304,N_2389);
and U3297 (N_3297,N_2468,N_2717);
nor U3298 (N_3298,N_2748,N_2835);
nand U3299 (N_3299,N_2805,N_2246);
and U3300 (N_3300,N_2731,N_2901);
and U3301 (N_3301,N_2858,N_2658);
nand U3302 (N_3302,N_2987,N_2629);
xnor U3303 (N_3303,N_2086,N_2603);
or U3304 (N_3304,N_2203,N_2471);
and U3305 (N_3305,N_2634,N_2781);
or U3306 (N_3306,N_2761,N_2470);
and U3307 (N_3307,N_2353,N_2251);
and U3308 (N_3308,N_2908,N_2579);
or U3309 (N_3309,N_2875,N_2557);
and U3310 (N_3310,N_2307,N_2375);
nor U3311 (N_3311,N_2912,N_2747);
nand U3312 (N_3312,N_2711,N_2733);
or U3313 (N_3313,N_2065,N_2859);
nand U3314 (N_3314,N_2035,N_2106);
nor U3315 (N_3315,N_2936,N_2738);
and U3316 (N_3316,N_2236,N_2437);
xnor U3317 (N_3317,N_2490,N_2548);
nor U3318 (N_3318,N_2973,N_2483);
nand U3319 (N_3319,N_2184,N_2955);
or U3320 (N_3320,N_2876,N_2542);
or U3321 (N_3321,N_2645,N_2555);
and U3322 (N_3322,N_2884,N_2354);
or U3323 (N_3323,N_2219,N_2551);
nor U3324 (N_3324,N_2600,N_2179);
and U3325 (N_3325,N_2361,N_2797);
nor U3326 (N_3326,N_2824,N_2541);
nand U3327 (N_3327,N_2550,N_2516);
nand U3328 (N_3328,N_2774,N_2553);
and U3329 (N_3329,N_2135,N_2743);
and U3330 (N_3330,N_2265,N_2014);
xor U3331 (N_3331,N_2099,N_2755);
nor U3332 (N_3332,N_2722,N_2764);
and U3333 (N_3333,N_2668,N_2860);
or U3334 (N_3334,N_2290,N_2318);
and U3335 (N_3335,N_2783,N_2952);
or U3336 (N_3336,N_2431,N_2308);
and U3337 (N_3337,N_2182,N_2811);
nor U3338 (N_3338,N_2211,N_2513);
or U3339 (N_3339,N_2017,N_2570);
nand U3340 (N_3340,N_2772,N_2186);
xnor U3341 (N_3341,N_2994,N_2968);
and U3342 (N_3342,N_2644,N_2656);
and U3343 (N_3343,N_2898,N_2562);
nand U3344 (N_3344,N_2280,N_2887);
nand U3345 (N_3345,N_2419,N_2237);
nand U3346 (N_3346,N_2429,N_2345);
nor U3347 (N_3347,N_2163,N_2234);
or U3348 (N_3348,N_2571,N_2021);
nand U3349 (N_3349,N_2923,N_2399);
or U3350 (N_3350,N_2120,N_2873);
or U3351 (N_3351,N_2648,N_2100);
nor U3352 (N_3352,N_2393,N_2245);
nand U3353 (N_3353,N_2558,N_2071);
or U3354 (N_3354,N_2750,N_2073);
nor U3355 (N_3355,N_2126,N_2674);
nor U3356 (N_3356,N_2093,N_2032);
and U3357 (N_3357,N_2222,N_2547);
nand U3358 (N_3358,N_2445,N_2616);
nor U3359 (N_3359,N_2972,N_2316);
xor U3360 (N_3360,N_2171,N_2526);
nor U3361 (N_3361,N_2416,N_2292);
xnor U3362 (N_3362,N_2433,N_2139);
or U3363 (N_3363,N_2654,N_2924);
nand U3364 (N_3364,N_2882,N_2200);
or U3365 (N_3365,N_2108,N_2505);
nand U3366 (N_3366,N_2008,N_2415);
nor U3367 (N_3367,N_2456,N_2374);
xor U3368 (N_3368,N_2030,N_2398);
nor U3369 (N_3369,N_2540,N_2287);
nor U3370 (N_3370,N_2784,N_2839);
and U3371 (N_3371,N_2663,N_2407);
or U3372 (N_3372,N_2864,N_2261);
and U3373 (N_3373,N_2878,N_2061);
xor U3374 (N_3374,N_2818,N_2500);
nand U3375 (N_3375,N_2865,N_2881);
xnor U3376 (N_3376,N_2782,N_2778);
and U3377 (N_3377,N_2984,N_2775);
or U3378 (N_3378,N_2406,N_2350);
and U3379 (N_3379,N_2853,N_2495);
or U3380 (N_3380,N_2631,N_2889);
nor U3381 (N_3381,N_2628,N_2151);
xnor U3382 (N_3382,N_2119,N_2395);
and U3383 (N_3383,N_2594,N_2450);
and U3384 (N_3384,N_2588,N_2708);
nand U3385 (N_3385,N_2802,N_2114);
nand U3386 (N_3386,N_2963,N_2417);
or U3387 (N_3387,N_2948,N_2739);
and U3388 (N_3388,N_2703,N_2828);
nor U3389 (N_3389,N_2258,N_2880);
xnor U3390 (N_3390,N_2247,N_2339);
or U3391 (N_3391,N_2147,N_2501);
nor U3392 (N_3392,N_2953,N_2671);
nor U3393 (N_3393,N_2466,N_2060);
and U3394 (N_3394,N_2917,N_2187);
and U3395 (N_3395,N_2507,N_2275);
nor U3396 (N_3396,N_2083,N_2310);
or U3397 (N_3397,N_2183,N_2801);
xnor U3398 (N_3398,N_2606,N_2130);
xor U3399 (N_3399,N_2728,N_2647);
nor U3400 (N_3400,N_2037,N_2554);
or U3401 (N_3401,N_2996,N_2074);
nor U3402 (N_3402,N_2208,N_2467);
xnor U3403 (N_3403,N_2418,N_2140);
xnor U3404 (N_3404,N_2435,N_2574);
and U3405 (N_3405,N_2052,N_2067);
and U3406 (N_3406,N_2975,N_2964);
or U3407 (N_3407,N_2678,N_2241);
nand U3408 (N_3408,N_2297,N_2855);
nor U3409 (N_3409,N_2978,N_2019);
xnor U3410 (N_3410,N_2619,N_2827);
nand U3411 (N_3411,N_2777,N_2286);
and U3412 (N_3412,N_2117,N_2347);
and U3413 (N_3413,N_2424,N_2005);
nor U3414 (N_3414,N_2613,N_2264);
xnor U3415 (N_3415,N_2794,N_2288);
nand U3416 (N_3416,N_2905,N_2423);
xor U3417 (N_3417,N_2016,N_2799);
nor U3418 (N_3418,N_2281,N_2886);
nor U3419 (N_3419,N_2655,N_2753);
xnor U3420 (N_3420,N_2652,N_2370);
or U3421 (N_3421,N_2869,N_2302);
or U3422 (N_3422,N_2202,N_2319);
nand U3423 (N_3423,N_2995,N_2480);
nand U3424 (N_3424,N_2022,N_2197);
and U3425 (N_3425,N_2825,N_2849);
and U3426 (N_3426,N_2888,N_2686);
nand U3427 (N_3427,N_2719,N_2759);
xnor U3428 (N_3428,N_2974,N_2402);
xnor U3429 (N_3429,N_2646,N_2599);
nor U3430 (N_3430,N_2018,N_2269);
or U3431 (N_3431,N_2363,N_2294);
and U3432 (N_3432,N_2856,N_2587);
nand U3433 (N_3433,N_2807,N_2448);
nand U3434 (N_3434,N_2463,N_2879);
and U3435 (N_3435,N_2862,N_2434);
or U3436 (N_3436,N_2152,N_2685);
nor U3437 (N_3437,N_2537,N_2055);
nor U3438 (N_3438,N_2341,N_2255);
xnor U3439 (N_3439,N_2457,N_2256);
xnor U3440 (N_3440,N_2796,N_2252);
nand U3441 (N_3441,N_2301,N_2890);
nand U3442 (N_3442,N_2593,N_2329);
nor U3443 (N_3443,N_2816,N_2221);
or U3444 (N_3444,N_2776,N_2107);
and U3445 (N_3445,N_2559,N_2462);
xnor U3446 (N_3446,N_2734,N_2714);
and U3447 (N_3447,N_2355,N_2696);
nor U3448 (N_3448,N_2838,N_2346);
or U3449 (N_3449,N_2330,N_2228);
and U3450 (N_3450,N_2718,N_2405);
and U3451 (N_3451,N_2408,N_2204);
or U3452 (N_3452,N_2191,N_2033);
nor U3453 (N_3453,N_2765,N_2919);
xnor U3454 (N_3454,N_2029,N_2190);
nor U3455 (N_3455,N_2344,N_2735);
nand U3456 (N_3456,N_2079,N_2534);
or U3457 (N_3457,N_2015,N_2609);
nor U3458 (N_3458,N_2161,N_2904);
nand U3459 (N_3459,N_2141,N_2266);
nand U3460 (N_3460,N_2284,N_2044);
nor U3461 (N_3461,N_2623,N_2274);
and U3462 (N_3462,N_2459,N_2476);
nor U3463 (N_3463,N_2027,N_2673);
xnor U3464 (N_3464,N_2198,N_2012);
or U3465 (N_3465,N_2094,N_2311);
nand U3466 (N_3466,N_2378,N_2742);
nor U3467 (N_3467,N_2527,N_2303);
nand U3468 (N_3468,N_2744,N_2665);
and U3469 (N_3469,N_2432,N_2787);
nor U3470 (N_3470,N_2503,N_2498);
or U3471 (N_3471,N_2695,N_2020);
and U3472 (N_3472,N_2766,N_2379);
nor U3473 (N_3473,N_2453,N_2447);
and U3474 (N_3474,N_2248,N_2833);
and U3475 (N_3475,N_2947,N_2697);
nor U3476 (N_3476,N_2851,N_2101);
and U3477 (N_3477,N_2767,N_2144);
xnor U3478 (N_3478,N_2552,N_2736);
nand U3479 (N_3479,N_2662,N_2156);
nand U3480 (N_3480,N_2983,N_2832);
or U3481 (N_3481,N_2664,N_2990);
nor U3482 (N_3482,N_2254,N_2846);
nand U3483 (N_3483,N_2635,N_2791);
xor U3484 (N_3484,N_2118,N_2170);
or U3485 (N_3485,N_2633,N_2939);
nand U3486 (N_3486,N_2096,N_2239);
nand U3487 (N_3487,N_2546,N_2473);
xor U3488 (N_3488,N_2192,N_2193);
and U3489 (N_3489,N_2874,N_2815);
nand U3490 (N_3490,N_2710,N_2036);
xor U3491 (N_3491,N_2013,N_2991);
or U3492 (N_3492,N_2692,N_2229);
nand U3493 (N_3493,N_2320,N_2870);
xor U3494 (N_3494,N_2932,N_2342);
xnor U3495 (N_3495,N_2918,N_2941);
and U3496 (N_3496,N_2359,N_2926);
nand U3497 (N_3497,N_2843,N_2982);
xor U3498 (N_3498,N_2104,N_2205);
nand U3499 (N_3499,N_2625,N_2907);
nor U3500 (N_3500,N_2847,N_2927);
nand U3501 (N_3501,N_2916,N_2918);
and U3502 (N_3502,N_2888,N_2085);
or U3503 (N_3503,N_2406,N_2622);
nand U3504 (N_3504,N_2463,N_2565);
xor U3505 (N_3505,N_2840,N_2399);
or U3506 (N_3506,N_2862,N_2385);
xnor U3507 (N_3507,N_2994,N_2551);
or U3508 (N_3508,N_2323,N_2566);
and U3509 (N_3509,N_2438,N_2665);
or U3510 (N_3510,N_2742,N_2226);
nor U3511 (N_3511,N_2130,N_2330);
or U3512 (N_3512,N_2937,N_2217);
and U3513 (N_3513,N_2884,N_2728);
nand U3514 (N_3514,N_2410,N_2661);
and U3515 (N_3515,N_2078,N_2742);
or U3516 (N_3516,N_2614,N_2899);
nor U3517 (N_3517,N_2676,N_2315);
or U3518 (N_3518,N_2430,N_2472);
nand U3519 (N_3519,N_2894,N_2840);
nand U3520 (N_3520,N_2582,N_2995);
xor U3521 (N_3521,N_2767,N_2942);
and U3522 (N_3522,N_2827,N_2580);
and U3523 (N_3523,N_2635,N_2524);
and U3524 (N_3524,N_2975,N_2200);
or U3525 (N_3525,N_2963,N_2603);
and U3526 (N_3526,N_2753,N_2934);
and U3527 (N_3527,N_2317,N_2053);
and U3528 (N_3528,N_2263,N_2167);
or U3529 (N_3529,N_2541,N_2567);
xor U3530 (N_3530,N_2705,N_2294);
nor U3531 (N_3531,N_2604,N_2138);
nand U3532 (N_3532,N_2257,N_2006);
or U3533 (N_3533,N_2526,N_2746);
and U3534 (N_3534,N_2579,N_2173);
nand U3535 (N_3535,N_2519,N_2033);
nor U3536 (N_3536,N_2045,N_2768);
or U3537 (N_3537,N_2960,N_2082);
nand U3538 (N_3538,N_2159,N_2211);
nor U3539 (N_3539,N_2256,N_2314);
or U3540 (N_3540,N_2884,N_2801);
and U3541 (N_3541,N_2038,N_2000);
nor U3542 (N_3542,N_2255,N_2797);
xnor U3543 (N_3543,N_2042,N_2235);
xor U3544 (N_3544,N_2430,N_2532);
and U3545 (N_3545,N_2086,N_2325);
and U3546 (N_3546,N_2925,N_2847);
nor U3547 (N_3547,N_2583,N_2530);
nor U3548 (N_3548,N_2798,N_2794);
nand U3549 (N_3549,N_2799,N_2547);
and U3550 (N_3550,N_2103,N_2505);
xor U3551 (N_3551,N_2059,N_2994);
and U3552 (N_3552,N_2427,N_2099);
and U3553 (N_3553,N_2856,N_2979);
xnor U3554 (N_3554,N_2795,N_2675);
xnor U3555 (N_3555,N_2470,N_2008);
xor U3556 (N_3556,N_2191,N_2669);
and U3557 (N_3557,N_2439,N_2151);
or U3558 (N_3558,N_2724,N_2858);
nand U3559 (N_3559,N_2965,N_2104);
or U3560 (N_3560,N_2472,N_2166);
xnor U3561 (N_3561,N_2425,N_2416);
xnor U3562 (N_3562,N_2017,N_2661);
xor U3563 (N_3563,N_2017,N_2878);
or U3564 (N_3564,N_2376,N_2806);
nand U3565 (N_3565,N_2293,N_2254);
and U3566 (N_3566,N_2619,N_2717);
nor U3567 (N_3567,N_2458,N_2279);
and U3568 (N_3568,N_2581,N_2662);
nor U3569 (N_3569,N_2804,N_2329);
and U3570 (N_3570,N_2447,N_2753);
and U3571 (N_3571,N_2464,N_2097);
nand U3572 (N_3572,N_2650,N_2471);
nand U3573 (N_3573,N_2836,N_2971);
and U3574 (N_3574,N_2804,N_2144);
xor U3575 (N_3575,N_2917,N_2526);
or U3576 (N_3576,N_2910,N_2132);
xor U3577 (N_3577,N_2619,N_2466);
nor U3578 (N_3578,N_2672,N_2498);
or U3579 (N_3579,N_2721,N_2375);
and U3580 (N_3580,N_2942,N_2585);
xnor U3581 (N_3581,N_2115,N_2712);
or U3582 (N_3582,N_2954,N_2992);
nand U3583 (N_3583,N_2848,N_2570);
nor U3584 (N_3584,N_2220,N_2797);
or U3585 (N_3585,N_2760,N_2221);
or U3586 (N_3586,N_2160,N_2476);
nand U3587 (N_3587,N_2612,N_2622);
xor U3588 (N_3588,N_2057,N_2072);
nor U3589 (N_3589,N_2611,N_2526);
nor U3590 (N_3590,N_2080,N_2459);
or U3591 (N_3591,N_2043,N_2622);
xnor U3592 (N_3592,N_2493,N_2022);
nand U3593 (N_3593,N_2197,N_2740);
xor U3594 (N_3594,N_2701,N_2279);
or U3595 (N_3595,N_2779,N_2094);
and U3596 (N_3596,N_2674,N_2786);
nor U3597 (N_3597,N_2542,N_2524);
or U3598 (N_3598,N_2072,N_2012);
xor U3599 (N_3599,N_2765,N_2703);
nor U3600 (N_3600,N_2079,N_2702);
nand U3601 (N_3601,N_2973,N_2411);
xnor U3602 (N_3602,N_2615,N_2595);
and U3603 (N_3603,N_2735,N_2766);
or U3604 (N_3604,N_2159,N_2910);
nand U3605 (N_3605,N_2503,N_2552);
nand U3606 (N_3606,N_2373,N_2909);
xnor U3607 (N_3607,N_2000,N_2370);
nor U3608 (N_3608,N_2471,N_2436);
xnor U3609 (N_3609,N_2105,N_2817);
and U3610 (N_3610,N_2679,N_2393);
nor U3611 (N_3611,N_2327,N_2157);
or U3612 (N_3612,N_2088,N_2938);
or U3613 (N_3613,N_2889,N_2955);
and U3614 (N_3614,N_2290,N_2465);
xnor U3615 (N_3615,N_2354,N_2753);
nor U3616 (N_3616,N_2652,N_2068);
nor U3617 (N_3617,N_2506,N_2207);
nand U3618 (N_3618,N_2065,N_2017);
nor U3619 (N_3619,N_2791,N_2345);
and U3620 (N_3620,N_2303,N_2966);
or U3621 (N_3621,N_2449,N_2896);
and U3622 (N_3622,N_2269,N_2541);
nand U3623 (N_3623,N_2398,N_2496);
or U3624 (N_3624,N_2814,N_2169);
nand U3625 (N_3625,N_2113,N_2480);
nor U3626 (N_3626,N_2693,N_2080);
nand U3627 (N_3627,N_2883,N_2682);
xor U3628 (N_3628,N_2580,N_2257);
or U3629 (N_3629,N_2896,N_2725);
xnor U3630 (N_3630,N_2229,N_2266);
and U3631 (N_3631,N_2662,N_2270);
nor U3632 (N_3632,N_2841,N_2557);
and U3633 (N_3633,N_2170,N_2500);
nor U3634 (N_3634,N_2998,N_2550);
nor U3635 (N_3635,N_2811,N_2227);
and U3636 (N_3636,N_2509,N_2417);
and U3637 (N_3637,N_2368,N_2749);
nand U3638 (N_3638,N_2765,N_2372);
nor U3639 (N_3639,N_2442,N_2046);
nor U3640 (N_3640,N_2121,N_2937);
xnor U3641 (N_3641,N_2936,N_2826);
xnor U3642 (N_3642,N_2318,N_2243);
nor U3643 (N_3643,N_2603,N_2368);
xnor U3644 (N_3644,N_2252,N_2966);
or U3645 (N_3645,N_2104,N_2747);
and U3646 (N_3646,N_2150,N_2527);
and U3647 (N_3647,N_2426,N_2420);
and U3648 (N_3648,N_2683,N_2602);
nand U3649 (N_3649,N_2315,N_2724);
and U3650 (N_3650,N_2234,N_2954);
and U3651 (N_3651,N_2023,N_2659);
or U3652 (N_3652,N_2400,N_2439);
or U3653 (N_3653,N_2024,N_2196);
xnor U3654 (N_3654,N_2446,N_2187);
nand U3655 (N_3655,N_2272,N_2198);
and U3656 (N_3656,N_2632,N_2443);
nand U3657 (N_3657,N_2261,N_2452);
and U3658 (N_3658,N_2910,N_2377);
and U3659 (N_3659,N_2179,N_2194);
nor U3660 (N_3660,N_2016,N_2981);
xor U3661 (N_3661,N_2342,N_2267);
nand U3662 (N_3662,N_2547,N_2010);
and U3663 (N_3663,N_2828,N_2971);
nand U3664 (N_3664,N_2306,N_2652);
nor U3665 (N_3665,N_2961,N_2119);
or U3666 (N_3666,N_2587,N_2706);
or U3667 (N_3667,N_2811,N_2022);
xnor U3668 (N_3668,N_2215,N_2100);
xnor U3669 (N_3669,N_2423,N_2077);
nor U3670 (N_3670,N_2522,N_2303);
and U3671 (N_3671,N_2726,N_2681);
xnor U3672 (N_3672,N_2740,N_2410);
xnor U3673 (N_3673,N_2798,N_2144);
nor U3674 (N_3674,N_2670,N_2001);
nand U3675 (N_3675,N_2206,N_2114);
xnor U3676 (N_3676,N_2582,N_2585);
xnor U3677 (N_3677,N_2898,N_2118);
and U3678 (N_3678,N_2201,N_2008);
nor U3679 (N_3679,N_2347,N_2644);
nand U3680 (N_3680,N_2982,N_2097);
or U3681 (N_3681,N_2503,N_2377);
xor U3682 (N_3682,N_2268,N_2538);
or U3683 (N_3683,N_2621,N_2015);
or U3684 (N_3684,N_2719,N_2560);
nand U3685 (N_3685,N_2785,N_2607);
nor U3686 (N_3686,N_2279,N_2562);
or U3687 (N_3687,N_2157,N_2079);
or U3688 (N_3688,N_2410,N_2357);
nor U3689 (N_3689,N_2890,N_2402);
xor U3690 (N_3690,N_2647,N_2743);
and U3691 (N_3691,N_2016,N_2763);
nor U3692 (N_3692,N_2061,N_2286);
xnor U3693 (N_3693,N_2147,N_2375);
nor U3694 (N_3694,N_2857,N_2115);
xnor U3695 (N_3695,N_2200,N_2585);
xor U3696 (N_3696,N_2303,N_2572);
nor U3697 (N_3697,N_2303,N_2346);
and U3698 (N_3698,N_2631,N_2731);
nor U3699 (N_3699,N_2868,N_2634);
xor U3700 (N_3700,N_2078,N_2859);
and U3701 (N_3701,N_2309,N_2942);
or U3702 (N_3702,N_2959,N_2718);
xnor U3703 (N_3703,N_2461,N_2469);
nand U3704 (N_3704,N_2990,N_2190);
nor U3705 (N_3705,N_2092,N_2787);
or U3706 (N_3706,N_2873,N_2541);
nor U3707 (N_3707,N_2590,N_2196);
xor U3708 (N_3708,N_2259,N_2235);
xnor U3709 (N_3709,N_2531,N_2038);
and U3710 (N_3710,N_2156,N_2062);
and U3711 (N_3711,N_2446,N_2328);
nand U3712 (N_3712,N_2796,N_2683);
nand U3713 (N_3713,N_2435,N_2997);
and U3714 (N_3714,N_2060,N_2710);
and U3715 (N_3715,N_2895,N_2725);
xnor U3716 (N_3716,N_2642,N_2463);
and U3717 (N_3717,N_2323,N_2384);
xnor U3718 (N_3718,N_2076,N_2234);
nand U3719 (N_3719,N_2660,N_2839);
nor U3720 (N_3720,N_2531,N_2413);
or U3721 (N_3721,N_2039,N_2501);
xor U3722 (N_3722,N_2725,N_2939);
xor U3723 (N_3723,N_2084,N_2082);
xnor U3724 (N_3724,N_2579,N_2079);
nor U3725 (N_3725,N_2440,N_2257);
nand U3726 (N_3726,N_2872,N_2674);
nor U3727 (N_3727,N_2425,N_2951);
or U3728 (N_3728,N_2328,N_2132);
nor U3729 (N_3729,N_2151,N_2403);
xnor U3730 (N_3730,N_2159,N_2321);
and U3731 (N_3731,N_2936,N_2917);
nor U3732 (N_3732,N_2325,N_2380);
nor U3733 (N_3733,N_2375,N_2124);
nand U3734 (N_3734,N_2852,N_2118);
xnor U3735 (N_3735,N_2315,N_2395);
xnor U3736 (N_3736,N_2843,N_2767);
or U3737 (N_3737,N_2753,N_2058);
xor U3738 (N_3738,N_2114,N_2558);
or U3739 (N_3739,N_2636,N_2979);
or U3740 (N_3740,N_2970,N_2357);
nand U3741 (N_3741,N_2022,N_2814);
and U3742 (N_3742,N_2281,N_2883);
xor U3743 (N_3743,N_2732,N_2253);
nand U3744 (N_3744,N_2335,N_2882);
or U3745 (N_3745,N_2641,N_2061);
xnor U3746 (N_3746,N_2389,N_2374);
xor U3747 (N_3747,N_2837,N_2118);
xnor U3748 (N_3748,N_2267,N_2969);
nand U3749 (N_3749,N_2442,N_2096);
and U3750 (N_3750,N_2706,N_2040);
nor U3751 (N_3751,N_2398,N_2892);
or U3752 (N_3752,N_2546,N_2815);
nor U3753 (N_3753,N_2004,N_2514);
xor U3754 (N_3754,N_2695,N_2190);
xor U3755 (N_3755,N_2124,N_2465);
nor U3756 (N_3756,N_2715,N_2309);
or U3757 (N_3757,N_2880,N_2554);
nand U3758 (N_3758,N_2933,N_2103);
nand U3759 (N_3759,N_2544,N_2240);
xnor U3760 (N_3760,N_2653,N_2801);
nor U3761 (N_3761,N_2526,N_2290);
nand U3762 (N_3762,N_2251,N_2358);
and U3763 (N_3763,N_2921,N_2396);
and U3764 (N_3764,N_2410,N_2147);
nand U3765 (N_3765,N_2048,N_2711);
xor U3766 (N_3766,N_2235,N_2742);
or U3767 (N_3767,N_2223,N_2437);
nand U3768 (N_3768,N_2177,N_2765);
nor U3769 (N_3769,N_2571,N_2681);
and U3770 (N_3770,N_2079,N_2810);
nand U3771 (N_3771,N_2305,N_2912);
xor U3772 (N_3772,N_2602,N_2012);
nor U3773 (N_3773,N_2136,N_2944);
nor U3774 (N_3774,N_2341,N_2146);
nor U3775 (N_3775,N_2905,N_2684);
nand U3776 (N_3776,N_2819,N_2597);
nor U3777 (N_3777,N_2374,N_2692);
nand U3778 (N_3778,N_2220,N_2407);
and U3779 (N_3779,N_2078,N_2367);
and U3780 (N_3780,N_2425,N_2509);
nand U3781 (N_3781,N_2042,N_2906);
nor U3782 (N_3782,N_2466,N_2200);
and U3783 (N_3783,N_2944,N_2823);
and U3784 (N_3784,N_2957,N_2952);
nor U3785 (N_3785,N_2461,N_2775);
nor U3786 (N_3786,N_2263,N_2945);
nor U3787 (N_3787,N_2094,N_2154);
xor U3788 (N_3788,N_2856,N_2851);
nor U3789 (N_3789,N_2559,N_2584);
nor U3790 (N_3790,N_2442,N_2333);
and U3791 (N_3791,N_2462,N_2059);
and U3792 (N_3792,N_2065,N_2655);
xor U3793 (N_3793,N_2083,N_2229);
xnor U3794 (N_3794,N_2065,N_2380);
or U3795 (N_3795,N_2299,N_2276);
and U3796 (N_3796,N_2674,N_2437);
and U3797 (N_3797,N_2715,N_2816);
nor U3798 (N_3798,N_2837,N_2364);
nand U3799 (N_3799,N_2538,N_2859);
nor U3800 (N_3800,N_2036,N_2174);
or U3801 (N_3801,N_2676,N_2252);
nor U3802 (N_3802,N_2423,N_2032);
and U3803 (N_3803,N_2366,N_2646);
nand U3804 (N_3804,N_2895,N_2472);
or U3805 (N_3805,N_2008,N_2742);
or U3806 (N_3806,N_2244,N_2009);
xor U3807 (N_3807,N_2479,N_2928);
nor U3808 (N_3808,N_2436,N_2587);
or U3809 (N_3809,N_2804,N_2519);
nor U3810 (N_3810,N_2193,N_2117);
xnor U3811 (N_3811,N_2391,N_2700);
nand U3812 (N_3812,N_2937,N_2702);
xor U3813 (N_3813,N_2486,N_2091);
nand U3814 (N_3814,N_2382,N_2044);
and U3815 (N_3815,N_2738,N_2013);
nand U3816 (N_3816,N_2499,N_2903);
xnor U3817 (N_3817,N_2781,N_2201);
xor U3818 (N_3818,N_2890,N_2411);
or U3819 (N_3819,N_2170,N_2081);
or U3820 (N_3820,N_2790,N_2972);
and U3821 (N_3821,N_2713,N_2439);
nand U3822 (N_3822,N_2797,N_2849);
nand U3823 (N_3823,N_2122,N_2247);
or U3824 (N_3824,N_2466,N_2634);
or U3825 (N_3825,N_2570,N_2936);
and U3826 (N_3826,N_2328,N_2313);
xor U3827 (N_3827,N_2209,N_2918);
nand U3828 (N_3828,N_2858,N_2270);
nor U3829 (N_3829,N_2484,N_2780);
xor U3830 (N_3830,N_2637,N_2000);
xor U3831 (N_3831,N_2352,N_2647);
or U3832 (N_3832,N_2377,N_2829);
xnor U3833 (N_3833,N_2650,N_2390);
and U3834 (N_3834,N_2037,N_2129);
nor U3835 (N_3835,N_2658,N_2095);
nor U3836 (N_3836,N_2316,N_2472);
nand U3837 (N_3837,N_2120,N_2967);
and U3838 (N_3838,N_2867,N_2488);
nand U3839 (N_3839,N_2440,N_2970);
or U3840 (N_3840,N_2198,N_2508);
nand U3841 (N_3841,N_2638,N_2405);
nor U3842 (N_3842,N_2588,N_2704);
nor U3843 (N_3843,N_2934,N_2998);
or U3844 (N_3844,N_2014,N_2942);
or U3845 (N_3845,N_2115,N_2847);
xor U3846 (N_3846,N_2937,N_2411);
nor U3847 (N_3847,N_2289,N_2384);
nor U3848 (N_3848,N_2326,N_2420);
xor U3849 (N_3849,N_2284,N_2354);
and U3850 (N_3850,N_2194,N_2810);
xnor U3851 (N_3851,N_2856,N_2928);
or U3852 (N_3852,N_2901,N_2882);
and U3853 (N_3853,N_2141,N_2520);
and U3854 (N_3854,N_2926,N_2259);
nand U3855 (N_3855,N_2315,N_2800);
and U3856 (N_3856,N_2933,N_2081);
xor U3857 (N_3857,N_2111,N_2699);
xnor U3858 (N_3858,N_2679,N_2759);
or U3859 (N_3859,N_2337,N_2645);
or U3860 (N_3860,N_2809,N_2237);
nor U3861 (N_3861,N_2056,N_2374);
nor U3862 (N_3862,N_2022,N_2729);
xor U3863 (N_3863,N_2190,N_2793);
or U3864 (N_3864,N_2519,N_2064);
nand U3865 (N_3865,N_2726,N_2563);
xnor U3866 (N_3866,N_2754,N_2486);
nor U3867 (N_3867,N_2076,N_2378);
nand U3868 (N_3868,N_2154,N_2924);
or U3869 (N_3869,N_2445,N_2712);
or U3870 (N_3870,N_2282,N_2757);
xor U3871 (N_3871,N_2093,N_2061);
and U3872 (N_3872,N_2584,N_2096);
or U3873 (N_3873,N_2936,N_2453);
and U3874 (N_3874,N_2454,N_2778);
nor U3875 (N_3875,N_2482,N_2213);
nor U3876 (N_3876,N_2044,N_2697);
and U3877 (N_3877,N_2542,N_2777);
nor U3878 (N_3878,N_2838,N_2063);
nand U3879 (N_3879,N_2292,N_2714);
nor U3880 (N_3880,N_2978,N_2053);
and U3881 (N_3881,N_2660,N_2074);
or U3882 (N_3882,N_2386,N_2156);
nor U3883 (N_3883,N_2732,N_2826);
nand U3884 (N_3884,N_2928,N_2066);
nor U3885 (N_3885,N_2361,N_2614);
nor U3886 (N_3886,N_2412,N_2615);
and U3887 (N_3887,N_2561,N_2727);
nand U3888 (N_3888,N_2674,N_2695);
xor U3889 (N_3889,N_2498,N_2847);
xor U3890 (N_3890,N_2165,N_2455);
and U3891 (N_3891,N_2527,N_2926);
xor U3892 (N_3892,N_2321,N_2754);
nor U3893 (N_3893,N_2461,N_2204);
xor U3894 (N_3894,N_2314,N_2477);
and U3895 (N_3895,N_2495,N_2933);
xnor U3896 (N_3896,N_2365,N_2452);
nor U3897 (N_3897,N_2953,N_2589);
nand U3898 (N_3898,N_2425,N_2353);
nand U3899 (N_3899,N_2727,N_2390);
nor U3900 (N_3900,N_2068,N_2023);
nand U3901 (N_3901,N_2767,N_2056);
and U3902 (N_3902,N_2009,N_2049);
nor U3903 (N_3903,N_2258,N_2176);
nand U3904 (N_3904,N_2415,N_2327);
nand U3905 (N_3905,N_2847,N_2856);
nor U3906 (N_3906,N_2713,N_2401);
nor U3907 (N_3907,N_2895,N_2752);
nand U3908 (N_3908,N_2015,N_2613);
and U3909 (N_3909,N_2918,N_2777);
nand U3910 (N_3910,N_2298,N_2592);
or U3911 (N_3911,N_2415,N_2998);
nand U3912 (N_3912,N_2773,N_2206);
xnor U3913 (N_3913,N_2791,N_2694);
or U3914 (N_3914,N_2483,N_2081);
xnor U3915 (N_3915,N_2663,N_2878);
xnor U3916 (N_3916,N_2583,N_2738);
and U3917 (N_3917,N_2083,N_2489);
xnor U3918 (N_3918,N_2251,N_2139);
xnor U3919 (N_3919,N_2868,N_2938);
nor U3920 (N_3920,N_2678,N_2083);
nand U3921 (N_3921,N_2105,N_2383);
nor U3922 (N_3922,N_2183,N_2783);
and U3923 (N_3923,N_2733,N_2240);
or U3924 (N_3924,N_2525,N_2348);
xnor U3925 (N_3925,N_2338,N_2384);
xnor U3926 (N_3926,N_2866,N_2432);
or U3927 (N_3927,N_2806,N_2794);
xnor U3928 (N_3928,N_2667,N_2951);
nand U3929 (N_3929,N_2892,N_2890);
nor U3930 (N_3930,N_2761,N_2751);
xor U3931 (N_3931,N_2856,N_2618);
nor U3932 (N_3932,N_2419,N_2379);
or U3933 (N_3933,N_2277,N_2485);
nand U3934 (N_3934,N_2501,N_2706);
xnor U3935 (N_3935,N_2940,N_2893);
or U3936 (N_3936,N_2818,N_2883);
xor U3937 (N_3937,N_2154,N_2637);
or U3938 (N_3938,N_2975,N_2360);
xor U3939 (N_3939,N_2165,N_2549);
xor U3940 (N_3940,N_2061,N_2394);
nor U3941 (N_3941,N_2386,N_2190);
xnor U3942 (N_3942,N_2869,N_2803);
xor U3943 (N_3943,N_2341,N_2102);
xor U3944 (N_3944,N_2890,N_2303);
xor U3945 (N_3945,N_2226,N_2709);
nand U3946 (N_3946,N_2648,N_2187);
or U3947 (N_3947,N_2455,N_2869);
xor U3948 (N_3948,N_2070,N_2792);
xor U3949 (N_3949,N_2318,N_2357);
and U3950 (N_3950,N_2178,N_2622);
or U3951 (N_3951,N_2561,N_2888);
or U3952 (N_3952,N_2217,N_2330);
nand U3953 (N_3953,N_2506,N_2131);
nor U3954 (N_3954,N_2442,N_2351);
and U3955 (N_3955,N_2456,N_2714);
or U3956 (N_3956,N_2644,N_2087);
and U3957 (N_3957,N_2486,N_2095);
nor U3958 (N_3958,N_2126,N_2846);
or U3959 (N_3959,N_2811,N_2518);
xor U3960 (N_3960,N_2132,N_2087);
nand U3961 (N_3961,N_2327,N_2205);
or U3962 (N_3962,N_2879,N_2919);
and U3963 (N_3963,N_2238,N_2747);
and U3964 (N_3964,N_2346,N_2957);
or U3965 (N_3965,N_2835,N_2716);
and U3966 (N_3966,N_2999,N_2853);
nor U3967 (N_3967,N_2036,N_2955);
and U3968 (N_3968,N_2137,N_2099);
xor U3969 (N_3969,N_2946,N_2790);
nor U3970 (N_3970,N_2783,N_2196);
or U3971 (N_3971,N_2650,N_2944);
nor U3972 (N_3972,N_2850,N_2701);
nand U3973 (N_3973,N_2496,N_2481);
nor U3974 (N_3974,N_2732,N_2674);
nor U3975 (N_3975,N_2972,N_2584);
or U3976 (N_3976,N_2445,N_2880);
xor U3977 (N_3977,N_2098,N_2254);
or U3978 (N_3978,N_2046,N_2536);
xnor U3979 (N_3979,N_2667,N_2977);
nand U3980 (N_3980,N_2296,N_2794);
and U3981 (N_3981,N_2798,N_2671);
nand U3982 (N_3982,N_2972,N_2154);
xor U3983 (N_3983,N_2877,N_2571);
or U3984 (N_3984,N_2418,N_2085);
nor U3985 (N_3985,N_2035,N_2050);
xor U3986 (N_3986,N_2064,N_2067);
xnor U3987 (N_3987,N_2376,N_2380);
nor U3988 (N_3988,N_2421,N_2114);
nand U3989 (N_3989,N_2231,N_2820);
nor U3990 (N_3990,N_2406,N_2117);
xor U3991 (N_3991,N_2099,N_2077);
xor U3992 (N_3992,N_2174,N_2556);
and U3993 (N_3993,N_2847,N_2347);
xnor U3994 (N_3994,N_2598,N_2588);
nand U3995 (N_3995,N_2440,N_2023);
and U3996 (N_3996,N_2065,N_2374);
and U3997 (N_3997,N_2783,N_2382);
and U3998 (N_3998,N_2030,N_2494);
xnor U3999 (N_3999,N_2165,N_2209);
nor U4000 (N_4000,N_3778,N_3054);
xor U4001 (N_4001,N_3139,N_3996);
nand U4002 (N_4002,N_3458,N_3107);
and U4003 (N_4003,N_3466,N_3822);
or U4004 (N_4004,N_3309,N_3669);
and U4005 (N_4005,N_3568,N_3471);
nand U4006 (N_4006,N_3888,N_3133);
nor U4007 (N_4007,N_3501,N_3104);
xor U4008 (N_4008,N_3140,N_3649);
nor U4009 (N_4009,N_3493,N_3038);
nand U4010 (N_4010,N_3771,N_3548);
xnor U4011 (N_4011,N_3224,N_3575);
nand U4012 (N_4012,N_3457,N_3535);
and U4013 (N_4013,N_3642,N_3354);
nor U4014 (N_4014,N_3141,N_3363);
and U4015 (N_4015,N_3276,N_3366);
nor U4016 (N_4016,N_3526,N_3823);
nor U4017 (N_4017,N_3444,N_3882);
nand U4018 (N_4018,N_3455,N_3904);
xor U4019 (N_4019,N_3052,N_3867);
or U4020 (N_4020,N_3325,N_3659);
xnor U4021 (N_4021,N_3071,N_3772);
xor U4022 (N_4022,N_3543,N_3099);
and U4023 (N_4023,N_3485,N_3293);
xnor U4024 (N_4024,N_3812,N_3709);
xnor U4025 (N_4025,N_3609,N_3060);
nor U4026 (N_4026,N_3044,N_3370);
nand U4027 (N_4027,N_3808,N_3103);
or U4028 (N_4028,N_3983,N_3136);
and U4029 (N_4029,N_3358,N_3591);
nor U4030 (N_4030,N_3583,N_3617);
xnor U4031 (N_4031,N_3936,N_3502);
xor U4032 (N_4032,N_3341,N_3157);
nor U4033 (N_4033,N_3719,N_3712);
xnor U4034 (N_4034,N_3307,N_3547);
and U4035 (N_4035,N_3885,N_3741);
or U4036 (N_4036,N_3556,N_3210);
and U4037 (N_4037,N_3966,N_3550);
xnor U4038 (N_4038,N_3462,N_3542);
or U4039 (N_4039,N_3045,N_3468);
or U4040 (N_4040,N_3766,N_3449);
nand U4041 (N_4041,N_3877,N_3735);
xor U4042 (N_4042,N_3914,N_3582);
and U4043 (N_4043,N_3807,N_3088);
xor U4044 (N_4044,N_3666,N_3160);
xor U4045 (N_4045,N_3789,N_3129);
nand U4046 (N_4046,N_3952,N_3943);
or U4047 (N_4047,N_3475,N_3379);
xnor U4048 (N_4048,N_3237,N_3990);
xnor U4049 (N_4049,N_3149,N_3090);
nor U4050 (N_4050,N_3767,N_3333);
xor U4051 (N_4051,N_3938,N_3442);
and U4052 (N_4052,N_3674,N_3204);
or U4053 (N_4053,N_3275,N_3962);
nand U4054 (N_4054,N_3544,N_3857);
and U4055 (N_4055,N_3170,N_3280);
xor U4056 (N_4056,N_3273,N_3618);
or U4057 (N_4057,N_3514,N_3029);
or U4058 (N_4058,N_3323,N_3711);
and U4059 (N_4059,N_3540,N_3383);
nor U4060 (N_4060,N_3113,N_3120);
nor U4061 (N_4061,N_3768,N_3218);
and U4062 (N_4062,N_3443,N_3085);
xnor U4063 (N_4063,N_3565,N_3788);
or U4064 (N_4064,N_3253,N_3685);
nand U4065 (N_4065,N_3357,N_3042);
and U4066 (N_4066,N_3942,N_3415);
or U4067 (N_4067,N_3026,N_3108);
and U4068 (N_4068,N_3720,N_3167);
nand U4069 (N_4069,N_3790,N_3626);
nor U4070 (N_4070,N_3787,N_3496);
or U4071 (N_4071,N_3021,N_3269);
or U4072 (N_4072,N_3118,N_3916);
and U4073 (N_4073,N_3033,N_3959);
nor U4074 (N_4074,N_3290,N_3834);
or U4075 (N_4075,N_3409,N_3176);
and U4076 (N_4076,N_3206,N_3827);
and U4077 (N_4077,N_3803,N_3607);
or U4078 (N_4078,N_3375,N_3076);
xor U4079 (N_4079,N_3963,N_3726);
nor U4080 (N_4080,N_3640,N_3081);
and U4081 (N_4081,N_3721,N_3845);
xor U4082 (N_4082,N_3267,N_3500);
nor U4083 (N_4083,N_3739,N_3016);
and U4084 (N_4084,N_3271,N_3737);
nor U4085 (N_4085,N_3738,N_3188);
and U4086 (N_4086,N_3478,N_3852);
xor U4087 (N_4087,N_3880,N_3911);
and U4088 (N_4088,N_3374,N_3153);
xor U4089 (N_4089,N_3154,N_3196);
and U4090 (N_4090,N_3704,N_3968);
xor U4091 (N_4091,N_3036,N_3467);
nand U4092 (N_4092,N_3553,N_3855);
or U4093 (N_4093,N_3481,N_3563);
and U4094 (N_4094,N_3873,N_3993);
nand U4095 (N_4095,N_3477,N_3486);
nor U4096 (N_4096,N_3894,N_3367);
and U4097 (N_4097,N_3921,N_3041);
or U4098 (N_4098,N_3804,N_3930);
nand U4099 (N_4099,N_3532,N_3774);
xnor U4100 (N_4100,N_3384,N_3339);
and U4101 (N_4101,N_3809,N_3117);
nor U4102 (N_4102,N_3075,N_3817);
or U4103 (N_4103,N_3572,N_3260);
nor U4104 (N_4104,N_3385,N_3459);
nor U4105 (N_4105,N_3030,N_3424);
xor U4106 (N_4106,N_3512,N_3746);
xnor U4107 (N_4107,N_3345,N_3687);
nor U4108 (N_4108,N_3628,N_3697);
and U4109 (N_4109,N_3780,N_3320);
xnor U4110 (N_4110,N_3889,N_3351);
and U4111 (N_4111,N_3641,N_3219);
and U4112 (N_4112,N_3982,N_3839);
xnor U4113 (N_4113,N_3994,N_3731);
xnor U4114 (N_4114,N_3348,N_3635);
nor U4115 (N_4115,N_3387,N_3710);
nand U4116 (N_4116,N_3503,N_3592);
nand U4117 (N_4117,N_3820,N_3465);
nor U4118 (N_4118,N_3454,N_3322);
or U4119 (N_4119,N_3944,N_3770);
or U4120 (N_4120,N_3631,N_3180);
nand U4121 (N_4121,N_3082,N_3037);
or U4122 (N_4122,N_3250,N_3364);
or U4123 (N_4123,N_3668,N_3574);
nor U4124 (N_4124,N_3225,N_3950);
nor U4125 (N_4125,N_3492,N_3412);
nor U4126 (N_4126,N_3303,N_3272);
nor U4127 (N_4127,N_3066,N_3907);
nand U4128 (N_4128,N_3425,N_3419);
nor U4129 (N_4129,N_3350,N_3517);
and U4130 (N_4130,N_3274,N_3521);
xnor U4131 (N_4131,N_3048,N_3956);
and U4132 (N_4132,N_3578,N_3017);
and U4133 (N_4133,N_3693,N_3009);
or U4134 (N_4134,N_3651,N_3308);
and U4135 (N_4135,N_3025,N_3988);
nor U4136 (N_4136,N_3059,N_3910);
xnor U4137 (N_4137,N_3106,N_3665);
nor U4138 (N_4138,N_3332,N_3560);
and U4139 (N_4139,N_3155,N_3960);
nor U4140 (N_4140,N_3247,N_3362);
or U4141 (N_4141,N_3476,N_3179);
xnor U4142 (N_4142,N_3433,N_3954);
nor U4143 (N_4143,N_3895,N_3184);
and U4144 (N_4144,N_3143,N_3879);
nor U4145 (N_4145,N_3297,N_3671);
and U4146 (N_4146,N_3035,N_3077);
or U4147 (N_4147,N_3003,N_3020);
nor U4148 (N_4148,N_3619,N_3523);
nor U4149 (N_4149,N_3688,N_3317);
and U4150 (N_4150,N_3000,N_3211);
or U4151 (N_4151,N_3352,N_3304);
and U4152 (N_4152,N_3802,N_3973);
and U4153 (N_4153,N_3326,N_3784);
and U4154 (N_4154,N_3122,N_3277);
or U4155 (N_4155,N_3606,N_3340);
nor U4156 (N_4156,N_3215,N_3980);
nand U4157 (N_4157,N_3216,N_3586);
nor U4158 (N_4158,N_3524,N_3414);
or U4159 (N_4159,N_3441,N_3534);
and U4160 (N_4160,N_3594,N_3469);
or U4161 (N_4161,N_3567,N_3028);
and U4162 (N_4162,N_3185,N_3564);
nor U4163 (N_4163,N_3813,N_3252);
nand U4164 (N_4164,N_3504,N_3010);
xnor U4165 (N_4165,N_3530,N_3762);
xor U4166 (N_4166,N_3418,N_3891);
nor U4167 (N_4167,N_3380,N_3699);
nand U4168 (N_4168,N_3102,N_3101);
nand U4169 (N_4169,N_3207,N_3427);
nand U4170 (N_4170,N_3286,N_3740);
nand U4171 (N_4171,N_3368,N_3310);
and U4172 (N_4172,N_3192,N_3198);
and U4173 (N_4173,N_3301,N_3908);
or U4174 (N_4174,N_3654,N_3109);
nand U4175 (N_4175,N_3437,N_3229);
nand U4176 (N_4176,N_3193,N_3981);
or U4177 (N_4177,N_3545,N_3612);
or U4178 (N_4178,N_3602,N_3440);
xnor U4179 (N_4179,N_3240,N_3506);
nand U4180 (N_4180,N_3546,N_3707);
and U4181 (N_4181,N_3974,N_3743);
nand U4182 (N_4182,N_3821,N_3264);
and U4183 (N_4183,N_3757,N_3878);
or U4184 (N_4184,N_3971,N_3448);
xnor U4185 (N_4185,N_3806,N_3844);
xor U4186 (N_4186,N_3865,N_3292);
and U4187 (N_4187,N_3142,N_3859);
and U4188 (N_4188,N_3828,N_3832);
xor U4189 (N_4189,N_3755,N_3324);
nor U4190 (N_4190,N_3881,N_3678);
xnor U4191 (N_4191,N_3646,N_3800);
nor U4192 (N_4192,N_3723,N_3957);
or U4193 (N_4193,N_3660,N_3152);
and U4194 (N_4194,N_3434,N_3151);
xor U4195 (N_4195,N_3393,N_3634);
nand U4196 (N_4196,N_3920,N_3472);
xnor U4197 (N_4197,N_3148,N_3413);
xor U4198 (N_4198,N_3166,N_3681);
or U4199 (N_4199,N_3793,N_3623);
nor U4200 (N_4200,N_3296,N_3664);
nor U4201 (N_4201,N_3933,N_3169);
xnor U4202 (N_4202,N_3769,N_3861);
or U4203 (N_4203,N_3032,N_3031);
or U4204 (N_4204,N_3639,N_3625);
xor U4205 (N_4205,N_3949,N_3846);
nor U4206 (N_4206,N_3482,N_3124);
or U4207 (N_4207,N_3976,N_3979);
nand U4208 (N_4208,N_3573,N_3168);
nor U4209 (N_4209,N_3062,N_3473);
nand U4210 (N_4210,N_3525,N_3715);
xnor U4211 (N_4211,N_3972,N_3138);
nand U4212 (N_4212,N_3835,N_3826);
xor U4213 (N_4213,N_3554,N_3001);
nand U4214 (N_4214,N_3019,N_3285);
or U4215 (N_4215,N_3328,N_3816);
xor U4216 (N_4216,N_3371,N_3116);
nor U4217 (N_4217,N_3334,N_3128);
nor U4218 (N_4218,N_3670,N_3751);
and U4219 (N_4219,N_3584,N_3024);
xor U4220 (N_4220,N_3801,N_3683);
nand U4221 (N_4221,N_3644,N_3661);
and U4222 (N_4222,N_3552,N_3680);
or U4223 (N_4223,N_3928,N_3756);
nand U4224 (N_4224,N_3825,N_3100);
nor U4225 (N_4225,N_3344,N_3588);
or U4226 (N_4226,N_3396,N_3833);
nand U4227 (N_4227,N_3604,N_3401);
and U4228 (N_4228,N_3335,N_3706);
nor U4229 (N_4229,N_3461,N_3522);
xor U4230 (N_4230,N_3776,N_3794);
xnor U4231 (N_4231,N_3255,N_3397);
nor U4232 (N_4232,N_3287,N_3713);
nor U4233 (N_4233,N_3946,N_3094);
nand U4234 (N_4234,N_3915,N_3410);
and U4235 (N_4235,N_3722,N_3676);
and U4236 (N_4236,N_3773,N_3163);
xor U4237 (N_4237,N_3819,N_3953);
and U4238 (N_4238,N_3093,N_3652);
nor U4239 (N_4239,N_3497,N_3539);
and U4240 (N_4240,N_3241,N_3248);
nor U4241 (N_4241,N_3692,N_3940);
xor U4242 (N_4242,N_3509,N_3931);
nand U4243 (N_4243,N_3551,N_3725);
and U4244 (N_4244,N_3923,N_3511);
nor U4245 (N_4245,N_3361,N_3989);
or U4246 (N_4246,N_3447,N_3898);
nor U4247 (N_4247,N_3172,N_3662);
nor U4248 (N_4248,N_3050,N_3558);
or U4249 (N_4249,N_3871,N_3520);
nor U4250 (N_4250,N_3658,N_3369);
xor U4251 (N_4251,N_3905,N_3200);
or U4252 (N_4252,N_3883,N_3708);
nor U4253 (N_4253,N_3555,N_3964);
and U4254 (N_4254,N_3810,N_3047);
nand U4255 (N_4255,N_3201,N_3236);
and U4256 (N_4256,N_3992,N_3799);
and U4257 (N_4257,N_3505,N_3622);
or U4258 (N_4258,N_3637,N_3251);
xnor U4259 (N_4259,N_3159,N_3795);
nor U4260 (N_4260,N_3013,N_3022);
nor U4261 (N_4261,N_3608,N_3394);
nor U4262 (N_4262,N_3446,N_3156);
xor U4263 (N_4263,N_3747,N_3049);
nor U4264 (N_4264,N_3579,N_3230);
nand U4265 (N_4265,N_3538,N_3400);
nor U4266 (N_4266,N_3599,N_3388);
nand U4267 (N_4267,N_3068,N_3329);
or U4268 (N_4268,N_3998,N_3495);
nand U4269 (N_4269,N_3703,N_3146);
nand U4270 (N_4270,N_3408,N_3638);
nand U4271 (N_4271,N_3158,N_3212);
or U4272 (N_4272,N_3053,N_3696);
xor U4273 (N_4273,N_3450,N_3187);
nor U4274 (N_4274,N_3298,N_3842);
xnor U4275 (N_4275,N_3125,N_3906);
xnor U4276 (N_4276,N_3675,N_3753);
nand U4277 (N_4277,N_3811,N_3541);
and U4278 (N_4278,N_3270,N_3111);
nand U4279 (N_4279,N_3299,N_3006);
nor U4280 (N_4280,N_3605,N_3258);
nand U4281 (N_4281,N_3145,N_3643);
nand U4282 (N_4282,N_3282,N_3074);
xor U4283 (N_4283,N_3590,N_3132);
nor U4284 (N_4284,N_3398,N_3884);
or U4285 (N_4285,N_3407,N_3431);
nor U4286 (N_4286,N_3259,N_3829);
nand U4287 (N_4287,N_3015,N_3672);
xnor U4288 (N_4288,N_3648,N_3005);
xor U4289 (N_4289,N_3222,N_3265);
xnor U4290 (N_4290,N_3797,N_3815);
or U4291 (N_4291,N_3718,N_3239);
nand U4292 (N_4292,N_3745,N_3087);
and U4293 (N_4293,N_3621,N_3389);
or U4294 (N_4294,N_3314,N_3734);
nor U4295 (N_4295,N_3945,N_3947);
nor U4296 (N_4296,N_3261,N_3430);
nand U4297 (N_4297,N_3012,N_3464);
and U4298 (N_4298,N_3585,N_3295);
and U4299 (N_4299,N_3866,N_3232);
nor U4300 (N_4300,N_3321,N_3566);
nand U4301 (N_4301,N_3549,N_3647);
nand U4302 (N_4302,N_3254,N_3694);
or U4303 (N_4303,N_3862,N_3202);
nor U4304 (N_4304,N_3775,N_3995);
nor U4305 (N_4305,N_3890,N_3760);
and U4306 (N_4306,N_3228,N_3856);
nor U4307 (N_4307,N_3864,N_3991);
and U4308 (N_4308,N_3597,N_3900);
and U4309 (N_4309,N_3406,N_3040);
nand U4310 (N_4310,N_3342,N_3353);
nand U4311 (N_4311,N_3186,N_3404);
nand U4312 (N_4312,N_3899,N_3925);
xnor U4313 (N_4313,N_3391,N_3456);
nor U4314 (N_4314,N_3513,N_3436);
xor U4315 (N_4315,N_3263,N_3359);
nand U4316 (N_4316,N_3395,N_3684);
or U4317 (N_4317,N_3836,N_3929);
xor U4318 (N_4318,N_3970,N_3932);
and U4319 (N_4319,N_3119,N_3913);
or U4320 (N_4320,N_3438,N_3014);
or U4321 (N_4321,N_3831,N_3377);
and U4322 (N_4322,N_3390,N_3965);
or U4323 (N_4323,N_3955,N_3347);
xor U4324 (N_4324,N_3249,N_3961);
or U4325 (N_4325,N_3203,N_3231);
and U4326 (N_4326,N_3302,N_3315);
nand U4327 (N_4327,N_3096,N_3453);
or U4328 (N_4328,N_3095,N_3234);
and U4329 (N_4329,N_3601,N_3798);
and U4330 (N_4330,N_3969,N_3986);
xor U4331 (N_4331,N_3902,N_3064);
or U4332 (N_4332,N_3392,N_3183);
or U4333 (N_4333,N_3451,N_3399);
or U4334 (N_4334,N_3758,N_3346);
nor U4335 (N_4335,N_3086,N_3761);
nor U4336 (N_4336,N_3221,N_3279);
or U4337 (N_4337,N_3291,N_3901);
nor U4338 (N_4338,N_3338,N_3130);
xor U4339 (N_4339,N_3978,N_3763);
nand U4340 (N_4340,N_3786,N_3097);
xor U4341 (N_4341,N_3135,N_3645);
xor U4342 (N_4342,N_3791,N_3903);
or U4343 (N_4343,N_3887,N_3750);
nand U4344 (N_4344,N_3581,N_3939);
nand U4345 (N_4345,N_3749,N_3373);
nor U4346 (N_4346,N_3084,N_3875);
and U4347 (N_4347,N_3519,N_3381);
or U4348 (N_4348,N_3349,N_3242);
nand U4349 (N_4349,N_3580,N_3405);
or U4350 (N_4350,N_3445,N_3886);
xor U4351 (N_4351,N_3587,N_3226);
or U4352 (N_4352,N_3008,N_3733);
nor U4353 (N_4353,N_3985,N_3951);
nand U4354 (N_4354,N_3208,N_3860);
or U4355 (N_4355,N_3420,N_3417);
and U4356 (N_4356,N_3796,N_3730);
nand U4357 (N_4357,N_3615,N_3863);
and U4358 (N_4358,N_3067,N_3058);
and U4359 (N_4359,N_3736,N_3209);
nand U4360 (N_4360,N_3174,N_3055);
and U4361 (N_4361,N_3557,N_3386);
nor U4362 (N_4362,N_3571,N_3422);
nand U4363 (N_4363,N_3510,N_3765);
nand U4364 (N_4364,N_3570,N_3474);
nand U4365 (N_4365,N_3779,N_3189);
nor U4366 (N_4366,N_3682,N_3777);
nand U4367 (N_4367,N_3217,N_3892);
nand U4368 (N_4368,N_3653,N_3917);
xnor U4369 (N_4369,N_3098,N_3343);
nor U4370 (N_4370,N_3701,N_3092);
and U4371 (N_4371,N_3613,N_3311);
or U4372 (N_4372,N_3171,N_3691);
nand U4373 (N_4373,N_3841,N_3507);
nand U4374 (N_4374,N_3752,N_3175);
or U4375 (N_4375,N_3294,N_3091);
or U4376 (N_4376,N_3110,N_3256);
nand U4377 (N_4377,N_3213,N_3403);
xnor U4378 (N_4378,N_3754,N_3714);
xor U4379 (N_4379,N_3576,N_3165);
nor U4380 (N_4380,N_3620,N_3365);
xor U4381 (N_4381,N_3056,N_3705);
nor U4382 (N_4382,N_3927,N_3488);
nor U4383 (N_4383,N_3480,N_3673);
xnor U4384 (N_4384,N_3593,N_3876);
or U4385 (N_4385,N_3997,N_3063);
xnor U4386 (N_4386,N_3614,N_3850);
nand U4387 (N_4387,N_3463,N_3849);
or U4388 (N_4388,N_3782,N_3837);
and U4389 (N_4389,N_3518,N_3327);
or U4390 (N_4390,N_3818,N_3896);
nand U4391 (N_4391,N_3499,N_3830);
nor U4392 (N_4392,N_3562,N_3987);
and U4393 (N_4393,N_3561,N_3007);
xnor U4394 (N_4394,N_3610,N_3838);
nand U4395 (N_4395,N_3489,N_3070);
or U4396 (N_4396,N_3624,N_3941);
and U4397 (N_4397,N_3182,N_3046);
or U4398 (N_4398,N_3233,N_3569);
xor U4399 (N_4399,N_3874,N_3123);
and U4400 (N_4400,N_3897,N_3069);
nand U4401 (N_4401,N_3266,N_3078);
xor U4402 (N_4402,N_3851,N_3195);
nand U4403 (N_4403,N_3194,N_3729);
nor U4404 (N_4404,N_3533,N_3732);
nor U4405 (N_4405,N_3843,N_3402);
or U4406 (N_4406,N_3783,N_3278);
and U4407 (N_4407,N_3716,N_3173);
xnor U4408 (N_4408,N_3657,N_3686);
or U4409 (N_4409,N_3268,N_3043);
xor U4410 (N_4410,N_3126,N_3717);
and U4411 (N_4411,N_3958,N_3537);
xnor U4412 (N_4412,N_3616,N_3079);
nand U4413 (N_4413,N_3121,N_3337);
or U4414 (N_4414,N_3912,N_3382);
nand U4415 (N_4415,N_3490,N_3805);
xor U4416 (N_4416,N_3004,N_3629);
nor U4417 (N_4417,N_3319,N_3611);
xor U4418 (N_4418,N_3487,N_3262);
or U4419 (N_4419,N_3948,N_3698);
xnor U4420 (N_4420,N_3460,N_3051);
or U4421 (N_4421,N_3061,N_3330);
or U4422 (N_4422,N_3792,N_3702);
or U4423 (N_4423,N_3870,N_3848);
or U4424 (N_4424,N_3423,N_3967);
and U4425 (N_4425,N_3162,N_3284);
or U4426 (N_4426,N_3426,N_3289);
nand U4427 (N_4427,N_3428,N_3360);
nand U4428 (N_4428,N_3840,N_3689);
or U4429 (N_4429,N_3089,N_3245);
and U4430 (N_4430,N_3536,N_3527);
xor U4431 (N_4431,N_3376,N_3679);
and U4432 (N_4432,N_3529,N_3589);
nand U4433 (N_4433,N_3633,N_3065);
or U4434 (N_4434,N_3144,N_3868);
or U4435 (N_4435,N_3114,N_3937);
xor U4436 (N_4436,N_3356,N_3023);
xnor U4437 (N_4437,N_3854,N_3039);
or U4438 (N_4438,N_3127,N_3600);
nor U4439 (N_4439,N_3115,N_3577);
nor U4440 (N_4440,N_3853,N_3781);
nand U4441 (N_4441,N_3214,N_3238);
nor U4442 (N_4442,N_3372,N_3919);
or U4443 (N_4443,N_3695,N_3824);
or U4444 (N_4444,N_3220,N_3281);
nand U4445 (N_4445,N_3002,N_3313);
or U4446 (N_4446,N_3484,N_3105);
and U4447 (N_4447,N_3677,N_3432);
nor U4448 (N_4448,N_3235,N_3147);
or U4449 (N_4449,N_3667,N_3027);
nand U4450 (N_4450,N_3452,N_3283);
and U4451 (N_4451,N_3177,N_3223);
and U4452 (N_4452,N_3999,N_3243);
and U4453 (N_4453,N_3439,N_3134);
nand U4454 (N_4454,N_3197,N_3416);
and U4455 (N_4455,N_3318,N_3312);
xnor U4456 (N_4456,N_3498,N_3636);
xor U4457 (N_4457,N_3748,N_3650);
or U4458 (N_4458,N_3977,N_3656);
nor U4459 (N_4459,N_3516,N_3057);
and U4460 (N_4460,N_3508,N_3494);
or U4461 (N_4461,N_3435,N_3491);
xor U4462 (N_4462,N_3011,N_3975);
nor U4463 (N_4463,N_3858,N_3018);
nor U4464 (N_4464,N_3814,N_3728);
nor U4465 (N_4465,N_3655,N_3421);
and U4466 (N_4466,N_3515,N_3316);
or U4467 (N_4467,N_3724,N_3083);
or U4468 (N_4468,N_3479,N_3531);
nand U4469 (N_4469,N_3227,N_3411);
and U4470 (N_4470,N_3080,N_3922);
or U4471 (N_4471,N_3300,N_3926);
nand U4472 (N_4472,N_3700,N_3872);
or U4473 (N_4473,N_3331,N_3190);
nor U4474 (N_4474,N_3246,N_3663);
nand U4475 (N_4475,N_3181,N_3759);
xnor U4476 (N_4476,N_3355,N_3305);
nor U4477 (N_4477,N_3984,N_3528);
and U4478 (N_4478,N_3690,N_3598);
nand U4479 (N_4479,N_3630,N_3924);
or U4480 (N_4480,N_3137,N_3191);
xnor U4481 (N_4481,N_3178,N_3131);
nor U4482 (N_4482,N_3199,N_3847);
nor U4483 (N_4483,N_3378,N_3596);
xor U4484 (N_4484,N_3306,N_3918);
nor U4485 (N_4485,N_3257,N_3785);
nor U4486 (N_4486,N_3244,N_3744);
or U4487 (N_4487,N_3934,N_3072);
nor U4488 (N_4488,N_3164,N_3603);
nand U4489 (N_4489,N_3112,N_3161);
or U4490 (N_4490,N_3429,N_3205);
nor U4491 (N_4491,N_3336,N_3627);
nor U4492 (N_4492,N_3483,N_3595);
nor U4493 (N_4493,N_3150,N_3909);
and U4494 (N_4494,N_3764,N_3727);
or U4495 (N_4495,N_3869,N_3034);
and U4496 (N_4496,N_3559,N_3073);
and U4497 (N_4497,N_3470,N_3742);
nand U4498 (N_4498,N_3935,N_3288);
nor U4499 (N_4499,N_3893,N_3632);
nand U4500 (N_4500,N_3603,N_3739);
xnor U4501 (N_4501,N_3032,N_3573);
nand U4502 (N_4502,N_3350,N_3767);
nand U4503 (N_4503,N_3749,N_3919);
or U4504 (N_4504,N_3017,N_3529);
xor U4505 (N_4505,N_3044,N_3212);
nor U4506 (N_4506,N_3639,N_3994);
nor U4507 (N_4507,N_3865,N_3201);
nor U4508 (N_4508,N_3227,N_3165);
xor U4509 (N_4509,N_3764,N_3328);
nor U4510 (N_4510,N_3036,N_3220);
or U4511 (N_4511,N_3380,N_3016);
or U4512 (N_4512,N_3181,N_3908);
xor U4513 (N_4513,N_3054,N_3111);
nor U4514 (N_4514,N_3428,N_3779);
nand U4515 (N_4515,N_3925,N_3397);
xor U4516 (N_4516,N_3227,N_3321);
or U4517 (N_4517,N_3002,N_3511);
nor U4518 (N_4518,N_3173,N_3974);
or U4519 (N_4519,N_3490,N_3730);
nor U4520 (N_4520,N_3401,N_3767);
and U4521 (N_4521,N_3555,N_3523);
xor U4522 (N_4522,N_3373,N_3708);
xor U4523 (N_4523,N_3569,N_3244);
or U4524 (N_4524,N_3237,N_3188);
or U4525 (N_4525,N_3521,N_3817);
or U4526 (N_4526,N_3476,N_3927);
xor U4527 (N_4527,N_3099,N_3519);
xor U4528 (N_4528,N_3496,N_3770);
and U4529 (N_4529,N_3452,N_3915);
nor U4530 (N_4530,N_3341,N_3931);
and U4531 (N_4531,N_3881,N_3113);
nor U4532 (N_4532,N_3183,N_3256);
nor U4533 (N_4533,N_3076,N_3748);
or U4534 (N_4534,N_3436,N_3570);
xnor U4535 (N_4535,N_3864,N_3826);
and U4536 (N_4536,N_3403,N_3729);
and U4537 (N_4537,N_3229,N_3499);
and U4538 (N_4538,N_3276,N_3055);
or U4539 (N_4539,N_3801,N_3587);
or U4540 (N_4540,N_3782,N_3301);
nor U4541 (N_4541,N_3383,N_3833);
xnor U4542 (N_4542,N_3688,N_3055);
xnor U4543 (N_4543,N_3251,N_3451);
or U4544 (N_4544,N_3106,N_3307);
or U4545 (N_4545,N_3049,N_3782);
nand U4546 (N_4546,N_3558,N_3093);
xnor U4547 (N_4547,N_3781,N_3181);
nand U4548 (N_4548,N_3378,N_3303);
nor U4549 (N_4549,N_3004,N_3514);
nand U4550 (N_4550,N_3540,N_3176);
nand U4551 (N_4551,N_3232,N_3698);
nand U4552 (N_4552,N_3775,N_3417);
nor U4553 (N_4553,N_3080,N_3656);
or U4554 (N_4554,N_3627,N_3241);
nand U4555 (N_4555,N_3392,N_3996);
nand U4556 (N_4556,N_3329,N_3056);
and U4557 (N_4557,N_3527,N_3564);
nor U4558 (N_4558,N_3470,N_3494);
xnor U4559 (N_4559,N_3967,N_3977);
xor U4560 (N_4560,N_3952,N_3311);
xnor U4561 (N_4561,N_3252,N_3982);
nor U4562 (N_4562,N_3493,N_3477);
nor U4563 (N_4563,N_3492,N_3850);
or U4564 (N_4564,N_3234,N_3648);
or U4565 (N_4565,N_3849,N_3960);
or U4566 (N_4566,N_3193,N_3870);
or U4567 (N_4567,N_3922,N_3894);
nand U4568 (N_4568,N_3169,N_3253);
nor U4569 (N_4569,N_3535,N_3066);
nand U4570 (N_4570,N_3301,N_3735);
nor U4571 (N_4571,N_3388,N_3034);
nor U4572 (N_4572,N_3267,N_3395);
xor U4573 (N_4573,N_3186,N_3175);
and U4574 (N_4574,N_3345,N_3914);
xor U4575 (N_4575,N_3709,N_3152);
or U4576 (N_4576,N_3991,N_3675);
or U4577 (N_4577,N_3663,N_3722);
or U4578 (N_4578,N_3351,N_3569);
xor U4579 (N_4579,N_3727,N_3927);
or U4580 (N_4580,N_3502,N_3266);
xor U4581 (N_4581,N_3589,N_3948);
nand U4582 (N_4582,N_3957,N_3825);
or U4583 (N_4583,N_3131,N_3779);
xnor U4584 (N_4584,N_3572,N_3484);
xor U4585 (N_4585,N_3238,N_3448);
or U4586 (N_4586,N_3180,N_3218);
or U4587 (N_4587,N_3079,N_3114);
and U4588 (N_4588,N_3841,N_3806);
and U4589 (N_4589,N_3848,N_3422);
nand U4590 (N_4590,N_3273,N_3938);
xnor U4591 (N_4591,N_3451,N_3593);
nor U4592 (N_4592,N_3493,N_3868);
and U4593 (N_4593,N_3749,N_3248);
nor U4594 (N_4594,N_3542,N_3383);
and U4595 (N_4595,N_3179,N_3033);
xnor U4596 (N_4596,N_3130,N_3989);
xor U4597 (N_4597,N_3929,N_3648);
and U4598 (N_4598,N_3610,N_3800);
or U4599 (N_4599,N_3810,N_3397);
xnor U4600 (N_4600,N_3096,N_3290);
and U4601 (N_4601,N_3682,N_3473);
or U4602 (N_4602,N_3401,N_3849);
nor U4603 (N_4603,N_3917,N_3434);
xor U4604 (N_4604,N_3669,N_3379);
or U4605 (N_4605,N_3365,N_3277);
xor U4606 (N_4606,N_3875,N_3768);
xnor U4607 (N_4607,N_3385,N_3890);
nor U4608 (N_4608,N_3052,N_3060);
or U4609 (N_4609,N_3470,N_3684);
or U4610 (N_4610,N_3609,N_3282);
xnor U4611 (N_4611,N_3027,N_3242);
nor U4612 (N_4612,N_3556,N_3833);
nand U4613 (N_4613,N_3836,N_3887);
nand U4614 (N_4614,N_3641,N_3061);
and U4615 (N_4615,N_3461,N_3447);
xor U4616 (N_4616,N_3565,N_3767);
or U4617 (N_4617,N_3560,N_3249);
nand U4618 (N_4618,N_3025,N_3878);
and U4619 (N_4619,N_3546,N_3377);
and U4620 (N_4620,N_3385,N_3816);
and U4621 (N_4621,N_3372,N_3271);
nor U4622 (N_4622,N_3787,N_3892);
nor U4623 (N_4623,N_3437,N_3907);
xor U4624 (N_4624,N_3884,N_3908);
or U4625 (N_4625,N_3213,N_3822);
nor U4626 (N_4626,N_3385,N_3916);
nand U4627 (N_4627,N_3842,N_3643);
nand U4628 (N_4628,N_3095,N_3822);
xnor U4629 (N_4629,N_3139,N_3112);
nor U4630 (N_4630,N_3174,N_3962);
or U4631 (N_4631,N_3004,N_3023);
and U4632 (N_4632,N_3549,N_3544);
and U4633 (N_4633,N_3395,N_3300);
nand U4634 (N_4634,N_3014,N_3391);
nor U4635 (N_4635,N_3123,N_3610);
nand U4636 (N_4636,N_3654,N_3658);
or U4637 (N_4637,N_3320,N_3641);
xnor U4638 (N_4638,N_3587,N_3320);
or U4639 (N_4639,N_3761,N_3226);
nand U4640 (N_4640,N_3077,N_3711);
xnor U4641 (N_4641,N_3033,N_3929);
and U4642 (N_4642,N_3761,N_3069);
nor U4643 (N_4643,N_3550,N_3369);
xor U4644 (N_4644,N_3768,N_3938);
or U4645 (N_4645,N_3649,N_3438);
and U4646 (N_4646,N_3200,N_3806);
nand U4647 (N_4647,N_3610,N_3848);
nor U4648 (N_4648,N_3219,N_3149);
nand U4649 (N_4649,N_3912,N_3567);
nor U4650 (N_4650,N_3426,N_3167);
nand U4651 (N_4651,N_3305,N_3465);
xnor U4652 (N_4652,N_3093,N_3151);
and U4653 (N_4653,N_3497,N_3226);
or U4654 (N_4654,N_3269,N_3751);
nor U4655 (N_4655,N_3297,N_3834);
or U4656 (N_4656,N_3467,N_3184);
nor U4657 (N_4657,N_3953,N_3847);
xor U4658 (N_4658,N_3340,N_3500);
xor U4659 (N_4659,N_3354,N_3600);
and U4660 (N_4660,N_3093,N_3409);
xnor U4661 (N_4661,N_3750,N_3148);
and U4662 (N_4662,N_3431,N_3663);
xor U4663 (N_4663,N_3148,N_3344);
nand U4664 (N_4664,N_3827,N_3452);
nor U4665 (N_4665,N_3471,N_3520);
and U4666 (N_4666,N_3855,N_3265);
or U4667 (N_4667,N_3215,N_3759);
xor U4668 (N_4668,N_3790,N_3697);
or U4669 (N_4669,N_3563,N_3962);
and U4670 (N_4670,N_3438,N_3748);
nor U4671 (N_4671,N_3475,N_3336);
or U4672 (N_4672,N_3323,N_3371);
and U4673 (N_4673,N_3412,N_3185);
xor U4674 (N_4674,N_3675,N_3269);
nand U4675 (N_4675,N_3753,N_3085);
nand U4676 (N_4676,N_3031,N_3816);
nand U4677 (N_4677,N_3698,N_3363);
xnor U4678 (N_4678,N_3888,N_3382);
and U4679 (N_4679,N_3333,N_3072);
and U4680 (N_4680,N_3757,N_3550);
or U4681 (N_4681,N_3931,N_3024);
or U4682 (N_4682,N_3314,N_3445);
nor U4683 (N_4683,N_3776,N_3407);
nor U4684 (N_4684,N_3807,N_3750);
xnor U4685 (N_4685,N_3137,N_3022);
nor U4686 (N_4686,N_3787,N_3012);
nor U4687 (N_4687,N_3110,N_3976);
nor U4688 (N_4688,N_3015,N_3251);
or U4689 (N_4689,N_3586,N_3009);
xnor U4690 (N_4690,N_3933,N_3774);
nand U4691 (N_4691,N_3283,N_3169);
nor U4692 (N_4692,N_3486,N_3356);
and U4693 (N_4693,N_3293,N_3102);
nor U4694 (N_4694,N_3796,N_3045);
xnor U4695 (N_4695,N_3110,N_3736);
and U4696 (N_4696,N_3561,N_3321);
and U4697 (N_4697,N_3037,N_3867);
nor U4698 (N_4698,N_3947,N_3951);
xor U4699 (N_4699,N_3239,N_3490);
nor U4700 (N_4700,N_3626,N_3509);
and U4701 (N_4701,N_3895,N_3009);
xor U4702 (N_4702,N_3271,N_3051);
xor U4703 (N_4703,N_3749,N_3995);
and U4704 (N_4704,N_3416,N_3776);
nand U4705 (N_4705,N_3560,N_3456);
xor U4706 (N_4706,N_3286,N_3847);
or U4707 (N_4707,N_3472,N_3782);
xor U4708 (N_4708,N_3605,N_3692);
or U4709 (N_4709,N_3253,N_3953);
xor U4710 (N_4710,N_3499,N_3700);
or U4711 (N_4711,N_3910,N_3674);
xnor U4712 (N_4712,N_3533,N_3992);
nand U4713 (N_4713,N_3483,N_3308);
nand U4714 (N_4714,N_3288,N_3812);
xor U4715 (N_4715,N_3073,N_3061);
nand U4716 (N_4716,N_3960,N_3150);
or U4717 (N_4717,N_3124,N_3037);
nor U4718 (N_4718,N_3425,N_3938);
or U4719 (N_4719,N_3736,N_3875);
or U4720 (N_4720,N_3416,N_3707);
nand U4721 (N_4721,N_3946,N_3229);
and U4722 (N_4722,N_3184,N_3605);
nor U4723 (N_4723,N_3004,N_3308);
nand U4724 (N_4724,N_3743,N_3668);
nor U4725 (N_4725,N_3562,N_3635);
or U4726 (N_4726,N_3600,N_3629);
xnor U4727 (N_4727,N_3392,N_3469);
or U4728 (N_4728,N_3836,N_3123);
nor U4729 (N_4729,N_3941,N_3315);
and U4730 (N_4730,N_3310,N_3671);
nor U4731 (N_4731,N_3610,N_3377);
nand U4732 (N_4732,N_3666,N_3229);
or U4733 (N_4733,N_3652,N_3110);
and U4734 (N_4734,N_3701,N_3536);
and U4735 (N_4735,N_3379,N_3944);
xor U4736 (N_4736,N_3027,N_3988);
and U4737 (N_4737,N_3000,N_3341);
nor U4738 (N_4738,N_3265,N_3570);
xor U4739 (N_4739,N_3608,N_3178);
nand U4740 (N_4740,N_3138,N_3108);
and U4741 (N_4741,N_3321,N_3415);
and U4742 (N_4742,N_3613,N_3756);
and U4743 (N_4743,N_3730,N_3334);
nor U4744 (N_4744,N_3861,N_3064);
or U4745 (N_4745,N_3502,N_3571);
or U4746 (N_4746,N_3538,N_3895);
xnor U4747 (N_4747,N_3543,N_3822);
nor U4748 (N_4748,N_3258,N_3593);
or U4749 (N_4749,N_3766,N_3821);
xnor U4750 (N_4750,N_3978,N_3756);
or U4751 (N_4751,N_3842,N_3377);
nor U4752 (N_4752,N_3551,N_3752);
nand U4753 (N_4753,N_3164,N_3286);
nor U4754 (N_4754,N_3726,N_3199);
or U4755 (N_4755,N_3507,N_3089);
xnor U4756 (N_4756,N_3285,N_3739);
xor U4757 (N_4757,N_3806,N_3763);
nor U4758 (N_4758,N_3948,N_3317);
or U4759 (N_4759,N_3069,N_3701);
xnor U4760 (N_4760,N_3835,N_3554);
nor U4761 (N_4761,N_3590,N_3330);
nand U4762 (N_4762,N_3913,N_3668);
and U4763 (N_4763,N_3043,N_3430);
or U4764 (N_4764,N_3641,N_3433);
nand U4765 (N_4765,N_3045,N_3429);
nor U4766 (N_4766,N_3062,N_3351);
or U4767 (N_4767,N_3389,N_3846);
nor U4768 (N_4768,N_3494,N_3374);
and U4769 (N_4769,N_3953,N_3568);
or U4770 (N_4770,N_3663,N_3682);
nor U4771 (N_4771,N_3757,N_3408);
nor U4772 (N_4772,N_3828,N_3366);
or U4773 (N_4773,N_3268,N_3320);
or U4774 (N_4774,N_3177,N_3790);
and U4775 (N_4775,N_3352,N_3669);
and U4776 (N_4776,N_3051,N_3205);
or U4777 (N_4777,N_3876,N_3337);
nor U4778 (N_4778,N_3917,N_3389);
or U4779 (N_4779,N_3708,N_3468);
nand U4780 (N_4780,N_3646,N_3568);
and U4781 (N_4781,N_3017,N_3506);
nor U4782 (N_4782,N_3982,N_3630);
and U4783 (N_4783,N_3918,N_3731);
xor U4784 (N_4784,N_3974,N_3431);
nand U4785 (N_4785,N_3546,N_3654);
and U4786 (N_4786,N_3821,N_3379);
and U4787 (N_4787,N_3878,N_3919);
or U4788 (N_4788,N_3602,N_3469);
or U4789 (N_4789,N_3868,N_3628);
xnor U4790 (N_4790,N_3038,N_3098);
nand U4791 (N_4791,N_3045,N_3551);
xnor U4792 (N_4792,N_3249,N_3435);
xor U4793 (N_4793,N_3591,N_3327);
nor U4794 (N_4794,N_3831,N_3628);
and U4795 (N_4795,N_3290,N_3303);
or U4796 (N_4796,N_3562,N_3990);
nand U4797 (N_4797,N_3170,N_3208);
nor U4798 (N_4798,N_3536,N_3401);
and U4799 (N_4799,N_3226,N_3505);
and U4800 (N_4800,N_3482,N_3430);
nor U4801 (N_4801,N_3893,N_3554);
or U4802 (N_4802,N_3855,N_3340);
nor U4803 (N_4803,N_3978,N_3073);
xor U4804 (N_4804,N_3130,N_3982);
xnor U4805 (N_4805,N_3156,N_3919);
nand U4806 (N_4806,N_3860,N_3206);
or U4807 (N_4807,N_3859,N_3467);
or U4808 (N_4808,N_3059,N_3417);
or U4809 (N_4809,N_3806,N_3373);
nor U4810 (N_4810,N_3590,N_3530);
or U4811 (N_4811,N_3596,N_3134);
or U4812 (N_4812,N_3292,N_3250);
and U4813 (N_4813,N_3316,N_3721);
xnor U4814 (N_4814,N_3151,N_3875);
or U4815 (N_4815,N_3137,N_3694);
nor U4816 (N_4816,N_3572,N_3219);
xor U4817 (N_4817,N_3717,N_3847);
xnor U4818 (N_4818,N_3157,N_3131);
and U4819 (N_4819,N_3601,N_3221);
nand U4820 (N_4820,N_3374,N_3475);
xnor U4821 (N_4821,N_3310,N_3892);
nor U4822 (N_4822,N_3138,N_3597);
nand U4823 (N_4823,N_3710,N_3512);
nor U4824 (N_4824,N_3050,N_3020);
nand U4825 (N_4825,N_3149,N_3036);
xor U4826 (N_4826,N_3332,N_3160);
nor U4827 (N_4827,N_3021,N_3116);
and U4828 (N_4828,N_3446,N_3296);
nor U4829 (N_4829,N_3723,N_3347);
nand U4830 (N_4830,N_3025,N_3881);
nor U4831 (N_4831,N_3435,N_3873);
xor U4832 (N_4832,N_3009,N_3665);
nor U4833 (N_4833,N_3127,N_3245);
nand U4834 (N_4834,N_3138,N_3821);
and U4835 (N_4835,N_3669,N_3892);
xnor U4836 (N_4836,N_3539,N_3366);
nor U4837 (N_4837,N_3853,N_3293);
or U4838 (N_4838,N_3064,N_3345);
xnor U4839 (N_4839,N_3615,N_3327);
nor U4840 (N_4840,N_3236,N_3129);
xnor U4841 (N_4841,N_3049,N_3649);
and U4842 (N_4842,N_3067,N_3432);
nand U4843 (N_4843,N_3153,N_3109);
or U4844 (N_4844,N_3850,N_3148);
and U4845 (N_4845,N_3544,N_3744);
nor U4846 (N_4846,N_3929,N_3375);
nand U4847 (N_4847,N_3681,N_3588);
and U4848 (N_4848,N_3132,N_3310);
or U4849 (N_4849,N_3949,N_3481);
nor U4850 (N_4850,N_3879,N_3969);
nand U4851 (N_4851,N_3399,N_3860);
and U4852 (N_4852,N_3245,N_3802);
xor U4853 (N_4853,N_3310,N_3389);
and U4854 (N_4854,N_3724,N_3196);
nor U4855 (N_4855,N_3372,N_3375);
or U4856 (N_4856,N_3570,N_3721);
and U4857 (N_4857,N_3928,N_3651);
nand U4858 (N_4858,N_3696,N_3024);
nand U4859 (N_4859,N_3101,N_3074);
nand U4860 (N_4860,N_3630,N_3116);
or U4861 (N_4861,N_3557,N_3859);
xnor U4862 (N_4862,N_3725,N_3821);
and U4863 (N_4863,N_3496,N_3188);
or U4864 (N_4864,N_3941,N_3349);
nand U4865 (N_4865,N_3000,N_3560);
or U4866 (N_4866,N_3598,N_3232);
xnor U4867 (N_4867,N_3201,N_3991);
xnor U4868 (N_4868,N_3569,N_3728);
xor U4869 (N_4869,N_3688,N_3130);
or U4870 (N_4870,N_3496,N_3762);
xnor U4871 (N_4871,N_3935,N_3638);
or U4872 (N_4872,N_3983,N_3266);
or U4873 (N_4873,N_3794,N_3947);
xor U4874 (N_4874,N_3311,N_3507);
nand U4875 (N_4875,N_3485,N_3084);
nor U4876 (N_4876,N_3468,N_3180);
nor U4877 (N_4877,N_3090,N_3675);
and U4878 (N_4878,N_3770,N_3301);
or U4879 (N_4879,N_3039,N_3538);
and U4880 (N_4880,N_3109,N_3335);
xor U4881 (N_4881,N_3465,N_3730);
nor U4882 (N_4882,N_3621,N_3641);
or U4883 (N_4883,N_3833,N_3423);
nand U4884 (N_4884,N_3525,N_3708);
nand U4885 (N_4885,N_3456,N_3422);
and U4886 (N_4886,N_3251,N_3317);
nor U4887 (N_4887,N_3405,N_3849);
nand U4888 (N_4888,N_3893,N_3053);
or U4889 (N_4889,N_3089,N_3123);
nand U4890 (N_4890,N_3030,N_3437);
and U4891 (N_4891,N_3859,N_3227);
nor U4892 (N_4892,N_3557,N_3188);
or U4893 (N_4893,N_3211,N_3035);
and U4894 (N_4894,N_3665,N_3182);
and U4895 (N_4895,N_3652,N_3510);
nand U4896 (N_4896,N_3569,N_3291);
or U4897 (N_4897,N_3593,N_3847);
nor U4898 (N_4898,N_3509,N_3836);
xor U4899 (N_4899,N_3881,N_3365);
nand U4900 (N_4900,N_3266,N_3836);
xor U4901 (N_4901,N_3804,N_3820);
nor U4902 (N_4902,N_3879,N_3102);
xor U4903 (N_4903,N_3595,N_3364);
xor U4904 (N_4904,N_3428,N_3482);
nor U4905 (N_4905,N_3216,N_3921);
or U4906 (N_4906,N_3471,N_3894);
nand U4907 (N_4907,N_3314,N_3951);
xor U4908 (N_4908,N_3470,N_3053);
nor U4909 (N_4909,N_3951,N_3448);
or U4910 (N_4910,N_3682,N_3513);
nor U4911 (N_4911,N_3197,N_3414);
nand U4912 (N_4912,N_3611,N_3335);
or U4913 (N_4913,N_3889,N_3121);
nand U4914 (N_4914,N_3699,N_3815);
and U4915 (N_4915,N_3300,N_3233);
nor U4916 (N_4916,N_3562,N_3191);
nor U4917 (N_4917,N_3065,N_3995);
xor U4918 (N_4918,N_3933,N_3203);
and U4919 (N_4919,N_3856,N_3273);
or U4920 (N_4920,N_3102,N_3133);
and U4921 (N_4921,N_3694,N_3275);
or U4922 (N_4922,N_3880,N_3246);
nor U4923 (N_4923,N_3309,N_3326);
nor U4924 (N_4924,N_3711,N_3725);
or U4925 (N_4925,N_3922,N_3574);
nor U4926 (N_4926,N_3649,N_3563);
or U4927 (N_4927,N_3211,N_3515);
and U4928 (N_4928,N_3159,N_3305);
and U4929 (N_4929,N_3991,N_3378);
nor U4930 (N_4930,N_3600,N_3744);
xnor U4931 (N_4931,N_3959,N_3669);
nor U4932 (N_4932,N_3594,N_3848);
or U4933 (N_4933,N_3555,N_3832);
nand U4934 (N_4934,N_3602,N_3425);
nor U4935 (N_4935,N_3147,N_3467);
nor U4936 (N_4936,N_3141,N_3137);
xnor U4937 (N_4937,N_3718,N_3597);
nor U4938 (N_4938,N_3355,N_3191);
xnor U4939 (N_4939,N_3340,N_3027);
nand U4940 (N_4940,N_3725,N_3766);
and U4941 (N_4941,N_3127,N_3235);
and U4942 (N_4942,N_3250,N_3695);
nand U4943 (N_4943,N_3219,N_3658);
and U4944 (N_4944,N_3962,N_3338);
nor U4945 (N_4945,N_3042,N_3062);
or U4946 (N_4946,N_3945,N_3633);
nand U4947 (N_4947,N_3067,N_3565);
or U4948 (N_4948,N_3098,N_3804);
xnor U4949 (N_4949,N_3757,N_3381);
nand U4950 (N_4950,N_3727,N_3944);
or U4951 (N_4951,N_3423,N_3926);
and U4952 (N_4952,N_3475,N_3580);
nor U4953 (N_4953,N_3162,N_3878);
nand U4954 (N_4954,N_3614,N_3705);
and U4955 (N_4955,N_3160,N_3509);
and U4956 (N_4956,N_3281,N_3197);
xnor U4957 (N_4957,N_3129,N_3682);
nor U4958 (N_4958,N_3375,N_3912);
and U4959 (N_4959,N_3813,N_3801);
and U4960 (N_4960,N_3987,N_3606);
nor U4961 (N_4961,N_3807,N_3511);
nor U4962 (N_4962,N_3736,N_3019);
xor U4963 (N_4963,N_3387,N_3537);
and U4964 (N_4964,N_3056,N_3195);
nor U4965 (N_4965,N_3076,N_3854);
nor U4966 (N_4966,N_3010,N_3424);
or U4967 (N_4967,N_3577,N_3755);
xnor U4968 (N_4968,N_3797,N_3174);
nor U4969 (N_4969,N_3577,N_3014);
and U4970 (N_4970,N_3343,N_3208);
xnor U4971 (N_4971,N_3072,N_3812);
nand U4972 (N_4972,N_3043,N_3660);
nand U4973 (N_4973,N_3241,N_3402);
xor U4974 (N_4974,N_3686,N_3184);
and U4975 (N_4975,N_3883,N_3699);
nand U4976 (N_4976,N_3634,N_3009);
nor U4977 (N_4977,N_3104,N_3969);
nand U4978 (N_4978,N_3317,N_3151);
nand U4979 (N_4979,N_3688,N_3723);
nand U4980 (N_4980,N_3762,N_3795);
xor U4981 (N_4981,N_3485,N_3011);
and U4982 (N_4982,N_3137,N_3778);
or U4983 (N_4983,N_3673,N_3852);
xnor U4984 (N_4984,N_3142,N_3118);
and U4985 (N_4985,N_3101,N_3813);
and U4986 (N_4986,N_3883,N_3255);
and U4987 (N_4987,N_3997,N_3006);
nor U4988 (N_4988,N_3091,N_3006);
or U4989 (N_4989,N_3982,N_3890);
nand U4990 (N_4990,N_3938,N_3677);
nor U4991 (N_4991,N_3991,N_3340);
nor U4992 (N_4992,N_3425,N_3083);
xnor U4993 (N_4993,N_3645,N_3578);
xor U4994 (N_4994,N_3177,N_3304);
xor U4995 (N_4995,N_3865,N_3993);
nand U4996 (N_4996,N_3500,N_3081);
nand U4997 (N_4997,N_3017,N_3491);
or U4998 (N_4998,N_3390,N_3716);
and U4999 (N_4999,N_3669,N_3544);
or U5000 (N_5000,N_4074,N_4864);
and U5001 (N_5001,N_4839,N_4451);
nor U5002 (N_5002,N_4202,N_4669);
nand U5003 (N_5003,N_4491,N_4267);
xnor U5004 (N_5004,N_4506,N_4969);
xor U5005 (N_5005,N_4510,N_4799);
nor U5006 (N_5006,N_4767,N_4374);
nor U5007 (N_5007,N_4789,N_4077);
nor U5008 (N_5008,N_4948,N_4290);
nand U5009 (N_5009,N_4396,N_4993);
nor U5010 (N_5010,N_4618,N_4414);
nand U5011 (N_5011,N_4141,N_4911);
and U5012 (N_5012,N_4447,N_4349);
nand U5013 (N_5013,N_4521,N_4189);
nand U5014 (N_5014,N_4909,N_4619);
or U5015 (N_5015,N_4338,N_4710);
xor U5016 (N_5016,N_4931,N_4024);
and U5017 (N_5017,N_4539,N_4643);
nor U5018 (N_5018,N_4719,N_4365);
nand U5019 (N_5019,N_4605,N_4484);
or U5020 (N_5020,N_4623,N_4314);
xor U5021 (N_5021,N_4846,N_4638);
xnor U5022 (N_5022,N_4676,N_4677);
xor U5023 (N_5023,N_4187,N_4337);
nor U5024 (N_5024,N_4462,N_4995);
and U5025 (N_5025,N_4952,N_4318);
or U5026 (N_5026,N_4299,N_4340);
nor U5027 (N_5027,N_4031,N_4256);
nor U5028 (N_5028,N_4956,N_4281);
nor U5029 (N_5029,N_4431,N_4656);
nor U5030 (N_5030,N_4511,N_4153);
xnor U5031 (N_5031,N_4670,N_4372);
xor U5032 (N_5032,N_4501,N_4014);
nor U5033 (N_5033,N_4070,N_4645);
nand U5034 (N_5034,N_4901,N_4184);
or U5035 (N_5035,N_4884,N_4761);
nor U5036 (N_5036,N_4019,N_4801);
or U5037 (N_5037,N_4116,N_4962);
nand U5038 (N_5038,N_4742,N_4207);
or U5039 (N_5039,N_4291,N_4311);
nor U5040 (N_5040,N_4143,N_4192);
or U5041 (N_5041,N_4792,N_4992);
nor U5042 (N_5042,N_4756,N_4673);
xnor U5043 (N_5043,N_4403,N_4715);
nand U5044 (N_5044,N_4428,N_4853);
and U5045 (N_5045,N_4978,N_4465);
nand U5046 (N_5046,N_4286,N_4829);
xor U5047 (N_5047,N_4251,N_4629);
xor U5048 (N_5048,N_4781,N_4865);
nand U5049 (N_5049,N_4800,N_4186);
nor U5050 (N_5050,N_4371,N_4814);
or U5051 (N_5051,N_4463,N_4749);
nand U5052 (N_5052,N_4035,N_4613);
nand U5053 (N_5053,N_4602,N_4348);
nand U5054 (N_5054,N_4620,N_4518);
nor U5055 (N_5055,N_4044,N_4214);
nand U5056 (N_5056,N_4998,N_4507);
xnor U5057 (N_5057,N_4907,N_4553);
or U5058 (N_5058,N_4776,N_4085);
and U5059 (N_5059,N_4900,N_4022);
or U5060 (N_5060,N_4101,N_4516);
nand U5061 (N_5061,N_4176,N_4603);
xnor U5062 (N_5062,N_4261,N_4012);
and U5063 (N_5063,N_4276,N_4493);
and U5064 (N_5064,N_4064,N_4357);
and U5065 (N_5065,N_4342,N_4148);
nand U5066 (N_5066,N_4566,N_4432);
nor U5067 (N_5067,N_4633,N_4018);
nand U5068 (N_5068,N_4275,N_4939);
xnor U5069 (N_5069,N_4177,N_4890);
nand U5070 (N_5070,N_4914,N_4960);
or U5071 (N_5071,N_4888,N_4413);
and U5072 (N_5072,N_4058,N_4115);
or U5073 (N_5073,N_4441,N_4168);
nand U5074 (N_5074,N_4504,N_4343);
nand U5075 (N_5075,N_4703,N_4784);
xor U5076 (N_5076,N_4273,N_4555);
nand U5077 (N_5077,N_4351,N_4512);
nand U5078 (N_5078,N_4968,N_4777);
nand U5079 (N_5079,N_4872,N_4097);
nor U5080 (N_5080,N_4034,N_4332);
nor U5081 (N_5081,N_4720,N_4768);
or U5082 (N_5082,N_4363,N_4745);
or U5083 (N_5083,N_4653,N_4098);
nand U5084 (N_5084,N_4461,N_4255);
and U5085 (N_5085,N_4200,N_4798);
nand U5086 (N_5086,N_4127,N_4306);
and U5087 (N_5087,N_4005,N_4717);
or U5088 (N_5088,N_4743,N_4046);
nand U5089 (N_5089,N_4389,N_4878);
nor U5090 (N_5090,N_4201,N_4775);
nor U5091 (N_5091,N_4500,N_4446);
and U5092 (N_5092,N_4236,N_4054);
and U5093 (N_5093,N_4233,N_4402);
and U5094 (N_5094,N_4837,N_4271);
nand U5095 (N_5095,N_4094,N_4631);
xor U5096 (N_5096,N_4686,N_4297);
and U5097 (N_5097,N_4532,N_4434);
or U5098 (N_5098,N_4104,N_4378);
and U5099 (N_5099,N_4688,N_4644);
xnor U5100 (N_5100,N_4660,N_4259);
nand U5101 (N_5101,N_4575,N_4408);
nand U5102 (N_5102,N_4301,N_4657);
xor U5103 (N_5103,N_4833,N_4099);
or U5104 (N_5104,N_4119,N_4066);
or U5105 (N_5105,N_4102,N_4223);
and U5106 (N_5106,N_4515,N_4114);
xor U5107 (N_5107,N_4771,N_4976);
nor U5108 (N_5108,N_4786,N_4088);
xor U5109 (N_5109,N_4812,N_4145);
xnor U5110 (N_5110,N_4885,N_4364);
nand U5111 (N_5111,N_4460,N_4687);
xor U5112 (N_5112,N_4078,N_4272);
xnor U5113 (N_5113,N_4997,N_4591);
or U5114 (N_5114,N_4950,N_4048);
or U5115 (N_5115,N_4758,N_4661);
and U5116 (N_5116,N_4377,N_4154);
nand U5117 (N_5117,N_4095,N_4017);
nor U5118 (N_5118,N_4527,N_4531);
nor U5119 (N_5119,N_4123,N_4152);
xnor U5120 (N_5120,N_4319,N_4409);
or U5121 (N_5121,N_4163,N_4367);
and U5122 (N_5122,N_4448,N_4739);
nand U5123 (N_5123,N_4795,N_4254);
and U5124 (N_5124,N_4140,N_4601);
and U5125 (N_5125,N_4245,N_4215);
nor U5126 (N_5126,N_4160,N_4838);
xnor U5127 (N_5127,N_4390,N_4690);
xor U5128 (N_5128,N_4737,N_4172);
nor U5129 (N_5129,N_4320,N_4821);
or U5130 (N_5130,N_4815,N_4651);
or U5131 (N_5131,N_4898,N_4525);
or U5132 (N_5132,N_4564,N_4877);
nor U5133 (N_5133,N_4309,N_4964);
and U5134 (N_5134,N_4668,N_4196);
nor U5135 (N_5135,N_4667,N_4622);
xnor U5136 (N_5136,N_4604,N_4862);
nand U5137 (N_5137,N_4039,N_4928);
or U5138 (N_5138,N_4716,N_4635);
nand U5139 (N_5139,N_4639,N_4664);
or U5140 (N_5140,N_4930,N_4100);
nand U5141 (N_5141,N_4361,N_4105);
and U5142 (N_5142,N_4130,N_4831);
or U5143 (N_5143,N_4443,N_4356);
or U5144 (N_5144,N_4033,N_4509);
nor U5145 (N_5145,N_4117,N_4004);
nor U5146 (N_5146,N_4963,N_4246);
nand U5147 (N_5147,N_4937,N_4834);
xnor U5148 (N_5148,N_4769,N_4029);
xor U5149 (N_5149,N_4126,N_4355);
and U5150 (N_5150,N_4183,N_4496);
nand U5151 (N_5151,N_4961,N_4763);
or U5152 (N_5152,N_4212,N_4991);
or U5153 (N_5153,N_4455,N_4472);
nand U5154 (N_5154,N_4237,N_4544);
nor U5155 (N_5155,N_4079,N_4996);
and U5156 (N_5156,N_4387,N_4983);
nor U5157 (N_5157,N_4327,N_4707);
nor U5158 (N_5158,N_4628,N_4709);
nand U5159 (N_5159,N_4535,N_4084);
xnor U5160 (N_5160,N_4806,N_4508);
xor U5161 (N_5161,N_4547,N_4832);
or U5162 (N_5162,N_4727,N_4208);
nor U5163 (N_5163,N_4418,N_4436);
or U5164 (N_5164,N_4241,N_4059);
or U5165 (N_5165,N_4173,N_4899);
nor U5166 (N_5166,N_4866,N_4615);
nor U5167 (N_5167,N_4442,N_4551);
or U5168 (N_5168,N_4287,N_4572);
xor U5169 (N_5169,N_4333,N_4445);
nor U5170 (N_5170,N_4411,N_4435);
nand U5171 (N_5171,N_4316,N_4379);
nand U5172 (N_5172,N_4003,N_4166);
or U5173 (N_5173,N_4230,N_4923);
nand U5174 (N_5174,N_4748,N_4701);
nand U5175 (N_5175,N_4897,N_4659);
nand U5176 (N_5176,N_4522,N_4596);
xor U5177 (N_5177,N_4787,N_4439);
nand U5178 (N_5178,N_4308,N_4876);
nand U5179 (N_5179,N_4250,N_4274);
or U5180 (N_5180,N_4556,N_4277);
nand U5181 (N_5181,N_4452,N_4951);
nor U5182 (N_5182,N_4981,N_4910);
nor U5183 (N_5183,N_4144,N_4975);
or U5184 (N_5184,N_4178,N_4430);
xor U5185 (N_5185,N_4157,N_4942);
nor U5186 (N_5186,N_4852,N_4699);
nand U5187 (N_5187,N_4696,N_4695);
or U5188 (N_5188,N_4616,N_4180);
or U5189 (N_5189,N_4811,N_4548);
nand U5190 (N_5190,N_4217,N_4469);
xnor U5191 (N_5191,N_4257,N_4825);
nand U5192 (N_5192,N_4871,N_4886);
and U5193 (N_5193,N_4336,N_4211);
and U5194 (N_5194,N_4822,N_4807);
nor U5195 (N_5195,N_4557,N_4398);
and U5196 (N_5196,N_4826,N_4940);
nand U5197 (N_5197,N_4471,N_4171);
xnor U5198 (N_5198,N_4785,N_4597);
or U5199 (N_5199,N_4027,N_4794);
and U5200 (N_5200,N_4561,N_4934);
nor U5201 (N_5201,N_4827,N_4858);
nor U5202 (N_5202,N_4497,N_4790);
nor U5203 (N_5203,N_4503,N_4570);
and U5204 (N_5204,N_4381,N_4331);
and U5205 (N_5205,N_4824,N_4574);
xor U5206 (N_5206,N_4725,N_4300);
nand U5207 (N_5207,N_4869,N_4793);
nor U5208 (N_5208,N_4219,N_4809);
nor U5209 (N_5209,N_4240,N_4971);
or U5210 (N_5210,N_4694,N_4685);
xnor U5211 (N_5211,N_4652,N_4209);
nand U5212 (N_5212,N_4195,N_4354);
xnor U5213 (N_5213,N_4921,N_4055);
xor U5214 (N_5214,N_4071,N_4175);
and U5215 (N_5215,N_4206,N_4627);
and U5216 (N_5216,N_4713,N_4540);
xnor U5217 (N_5217,N_4086,N_4167);
xor U5218 (N_5218,N_4658,N_4181);
xnor U5219 (N_5219,N_4285,N_4955);
and U5220 (N_5220,N_4642,N_4429);
nand U5221 (N_5221,N_4524,N_4326);
xnor U5222 (N_5222,N_4315,N_4662);
xor U5223 (N_5223,N_4689,N_4947);
nand U5224 (N_5224,N_4056,N_4323);
nand U5225 (N_5225,N_4844,N_4068);
xnor U5226 (N_5226,N_4227,N_4595);
and U5227 (N_5227,N_4334,N_4502);
and U5228 (N_5228,N_4953,N_4624);
xor U5229 (N_5229,N_4693,N_4067);
nand U5230 (N_5230,N_4288,N_4213);
or U5231 (N_5231,N_4358,N_4370);
and U5232 (N_5232,N_4249,N_4751);
and U5233 (N_5233,N_4857,N_4382);
nor U5234 (N_5234,N_4816,N_4530);
xor U5235 (N_5235,N_4120,N_4580);
nor U5236 (N_5236,N_4860,N_4185);
or U5237 (N_5237,N_4646,N_4517);
nand U5238 (N_5238,N_4835,N_4045);
nand U5239 (N_5239,N_4766,N_4736);
nor U5240 (N_5240,N_4782,N_4984);
nand U5241 (N_5241,N_4464,N_4945);
xnor U5242 (N_5242,N_4009,N_4577);
and U5243 (N_5243,N_4573,N_4474);
nand U5244 (N_5244,N_4149,N_4134);
nor U5245 (N_5245,N_4599,N_4704);
or U5246 (N_5246,N_4242,N_4051);
or U5247 (N_5247,N_4922,N_4891);
or U5248 (N_5248,N_4295,N_4558);
nand U5249 (N_5249,N_4234,N_4422);
nor U5250 (N_5250,N_4121,N_4020);
nand U5251 (N_5251,N_4731,N_4567);
or U5252 (N_5252,N_4142,N_4892);
nand U5253 (N_5253,N_4165,N_4889);
nor U5254 (N_5254,N_4093,N_4394);
nand U5255 (N_5255,N_4823,N_4083);
nor U5256 (N_5256,N_4882,N_4714);
nand U5257 (N_5257,N_4526,N_4873);
nand U5258 (N_5258,N_4729,N_4543);
and U5259 (N_5259,N_4855,N_4069);
nand U5260 (N_5260,N_4546,N_4060);
xor U5261 (N_5261,N_4129,N_4158);
or U5262 (N_5262,N_4162,N_4006);
nand U5263 (N_5263,N_4926,N_4279);
or U5264 (N_5264,N_4708,N_4298);
and U5265 (N_5265,N_4265,N_4985);
nand U5266 (N_5266,N_4542,N_4625);
nor U5267 (N_5267,N_4746,N_4593);
nor U5268 (N_5268,N_4682,N_4549);
xnor U5269 (N_5269,N_4994,N_4359);
nor U5270 (N_5270,N_4216,N_4438);
nand U5271 (N_5271,N_4589,N_4513);
or U5272 (N_5272,N_4966,N_4550);
and U5273 (N_5273,N_4845,N_4458);
and U5274 (N_5274,N_4916,N_4170);
xnor U5275 (N_5275,N_4481,N_4150);
nor U5276 (N_5276,N_4151,N_4393);
xnor U5277 (N_5277,N_4959,N_4459);
or U5278 (N_5278,N_4426,N_4606);
and U5279 (N_5279,N_4841,N_4023);
nand U5280 (N_5280,N_4702,N_4637);
xnor U5281 (N_5281,N_4982,N_4405);
xnor U5282 (N_5282,N_4920,N_4747);
nor U5283 (N_5283,N_4388,N_4346);
or U5284 (N_5284,N_4042,N_4002);
nand U5285 (N_5285,N_4808,N_4565);
or U5286 (N_5286,N_4568,N_4541);
nor U5287 (N_5287,N_4712,N_4610);
nand U5288 (N_5288,N_4147,N_4312);
nor U5289 (N_5289,N_4569,N_4609);
nor U5290 (N_5290,N_4278,N_4305);
nand U5291 (N_5291,N_4385,N_4466);
nor U5292 (N_5292,N_4943,N_4819);
or U5293 (N_5293,N_4905,N_4016);
nand U5294 (N_5294,N_4999,N_4182);
or U5295 (N_5295,N_4650,N_4376);
nand U5296 (N_5296,N_4013,N_4025);
and U5297 (N_5297,N_4373,N_4190);
xnor U5298 (N_5298,N_4457,N_4655);
xnor U5299 (N_5299,N_4345,N_4118);
nand U5300 (N_5300,N_4425,N_4681);
xnor U5301 (N_5301,N_4938,N_4954);
nand U5302 (N_5302,N_4562,N_4559);
xnor U5303 (N_5303,N_4738,N_4037);
nor U5304 (N_5304,N_4107,N_4958);
xor U5305 (N_5305,N_4967,N_4444);
and U5306 (N_5306,N_4818,N_4698);
xnor U5307 (N_5307,N_4571,N_4990);
nand U5308 (N_5308,N_4584,N_4988);
nor U5309 (N_5309,N_4483,N_4339);
and U5310 (N_5310,N_4598,N_4590);
and U5311 (N_5311,N_4863,N_4137);
xnor U5312 (N_5312,N_4310,N_4244);
or U5313 (N_5313,N_4529,N_4796);
and U5314 (N_5314,N_4235,N_4062);
or U5315 (N_5315,N_4607,N_4733);
nor U5316 (N_5316,N_4840,N_4392);
xnor U5317 (N_5317,N_4258,N_4700);
xnor U5318 (N_5318,N_4061,N_4049);
or U5319 (N_5319,N_4433,N_4292);
nor U5320 (N_5320,N_4854,N_4893);
nand U5321 (N_5321,N_4269,N_4554);
nor U5322 (N_5322,N_4454,N_4936);
and U5323 (N_5323,N_4280,N_4762);
nand U5324 (N_5324,N_4894,N_4404);
xor U5325 (N_5325,N_4296,N_4247);
nor U5326 (N_5326,N_4155,N_4828);
nand U5327 (N_5327,N_4270,N_4802);
and U5328 (N_5328,N_4397,N_4581);
nand U5329 (N_5329,N_4538,N_4908);
nand U5330 (N_5330,N_4335,N_4552);
nor U5331 (N_5331,N_4805,N_4096);
or U5332 (N_5332,N_4110,N_4919);
nand U5333 (N_5333,N_4132,N_4477);
or U5334 (N_5334,N_4325,N_4427);
nand U5335 (N_5335,N_4011,N_4222);
xor U5336 (N_5336,N_4913,N_4933);
xor U5337 (N_5337,N_4412,N_4220);
nor U5338 (N_5338,N_4671,N_4680);
nor U5339 (N_5339,N_4849,N_4239);
nor U5340 (N_5340,N_4489,N_4475);
and U5341 (N_5341,N_4161,N_4663);
xnor U5342 (N_5342,N_4076,N_4592);
nor U5343 (N_5343,N_4740,N_4935);
or U5344 (N_5344,N_4205,N_4986);
nand U5345 (N_5345,N_4523,N_4401);
xnor U5346 (N_5346,N_4804,N_4410);
xor U5347 (N_5347,N_4294,N_4912);
xor U5348 (N_5348,N_4896,N_4759);
or U5349 (N_5349,N_4082,N_4156);
xnor U5350 (N_5350,N_4199,N_4588);
nor U5351 (N_5351,N_4399,N_4050);
nor U5352 (N_5352,N_4360,N_4440);
nor U5353 (N_5353,N_4494,N_4263);
or U5354 (N_5354,N_4416,N_4586);
nor U5355 (N_5355,N_4253,N_4052);
and U5356 (N_5356,N_4282,N_4437);
nor U5357 (N_5357,N_4957,N_4228);
xor U5358 (N_5358,N_4423,N_4760);
or U5359 (N_5359,N_4772,N_4848);
or U5360 (N_5360,N_4861,N_4090);
or U5361 (N_5361,N_4973,N_4752);
or U5362 (N_5362,N_4053,N_4368);
or U5363 (N_5363,N_4924,N_4868);
nor U5364 (N_5364,N_4534,N_4036);
nand U5365 (N_5365,N_4600,N_4779);
or U5366 (N_5366,N_4634,N_4081);
or U5367 (N_5367,N_4225,N_4879);
xnor U5368 (N_5368,N_4203,N_4103);
and U5369 (N_5369,N_4000,N_4488);
xnor U5370 (N_5370,N_4753,N_4266);
nor U5371 (N_5371,N_4765,N_4473);
nor U5372 (N_5372,N_4684,N_4197);
or U5373 (N_5373,N_4450,N_4136);
nand U5374 (N_5374,N_4386,N_4353);
and U5375 (N_5375,N_4672,N_4917);
xor U5376 (N_5376,N_4362,N_4974);
nand U5377 (N_5377,N_4395,N_4859);
xnor U5378 (N_5378,N_4728,N_4970);
and U5379 (N_5379,N_4722,N_4499);
xnor U5380 (N_5380,N_4467,N_4870);
xor U5381 (N_5381,N_4578,N_4579);
nand U5382 (N_5382,N_4453,N_4867);
nor U5383 (N_5383,N_4730,N_4449);
and U5384 (N_5384,N_4075,N_4063);
or U5385 (N_5385,N_4350,N_4918);
nand U5386 (N_5386,N_4179,N_4065);
or U5387 (N_5387,N_4611,N_4734);
and U5388 (N_5388,N_4721,N_4262);
nand U5389 (N_5389,N_4906,N_4773);
nand U5390 (N_5390,N_4881,N_4480);
xnor U5391 (N_5391,N_4585,N_4987);
or U5392 (N_5392,N_4038,N_4492);
or U5393 (N_5393,N_4293,N_4243);
nand U5394 (N_5394,N_4226,N_4621);
nor U5395 (N_5395,N_4490,N_4109);
or U5396 (N_5396,N_4537,N_4674);
xor U5397 (N_5397,N_4560,N_4304);
nand U5398 (N_5398,N_4417,N_4232);
nand U5399 (N_5399,N_4112,N_4666);
nor U5400 (N_5400,N_4965,N_4008);
and U5401 (N_5401,N_4057,N_4617);
nand U5402 (N_5402,N_4904,N_4007);
xor U5403 (N_5403,N_4697,N_4159);
nand U5404 (N_5404,N_4317,N_4903);
or U5405 (N_5405,N_4757,N_4755);
xor U5406 (N_5406,N_4091,N_4576);
and U5407 (N_5407,N_4384,N_4724);
or U5408 (N_5408,N_4092,N_4977);
nand U5409 (N_5409,N_4648,N_4188);
or U5410 (N_5410,N_4264,N_4420);
and U5411 (N_5411,N_4505,N_4224);
and U5412 (N_5412,N_4321,N_4851);
and U5413 (N_5413,N_4106,N_4347);
or U5414 (N_5414,N_4582,N_4283);
xor U5415 (N_5415,N_4400,N_4783);
nand U5416 (N_5416,N_4972,N_4847);
nand U5417 (N_5417,N_4630,N_4303);
and U5418 (N_5418,N_4989,N_4407);
xor U5419 (N_5419,N_4632,N_4883);
nand U5420 (N_5420,N_4665,N_4640);
nor U5421 (N_5421,N_4260,N_4754);
nor U5422 (N_5422,N_4268,N_4647);
or U5423 (N_5423,N_4626,N_4380);
nor U5424 (N_5424,N_4679,N_4842);
or U5425 (N_5425,N_4850,N_4880);
and U5426 (N_5426,N_4391,N_4415);
or U5427 (N_5427,N_4307,N_4778);
and U5428 (N_5428,N_4583,N_4229);
xnor U5429 (N_5429,N_4041,N_4032);
xor U5430 (N_5430,N_4528,N_4139);
and U5431 (N_5431,N_4612,N_4043);
nor U5432 (N_5432,N_4944,N_4289);
or U5433 (N_5433,N_4636,N_4111);
xnor U5434 (N_5434,N_4198,N_4191);
nor U5435 (N_5435,N_4476,N_4369);
and U5436 (N_5436,N_4741,N_4820);
and U5437 (N_5437,N_4533,N_4485);
xor U5438 (N_5438,N_4675,N_4419);
nor U5439 (N_5439,N_4221,N_4514);
nor U5440 (N_5440,N_4744,N_4813);
nor U5441 (N_5441,N_4113,N_4706);
xor U5442 (N_5442,N_4887,N_4705);
nand U5443 (N_5443,N_4138,N_4536);
and U5444 (N_5444,N_4780,N_4010);
xor U5445 (N_5445,N_4366,N_4193);
nand U5446 (N_5446,N_4545,N_4594);
and U5447 (N_5447,N_4726,N_4238);
nor U5448 (N_5448,N_4949,N_4080);
nor U5449 (N_5449,N_4830,N_4470);
nor U5450 (N_5450,N_4128,N_4895);
or U5451 (N_5451,N_4482,N_4692);
and U5452 (N_5452,N_4204,N_4015);
xnor U5453 (N_5453,N_4302,N_4980);
xnor U5454 (N_5454,N_4764,N_4875);
xnor U5455 (N_5455,N_4468,N_4073);
nor U5456 (N_5456,N_4486,N_4519);
xnor U5457 (N_5457,N_4479,N_4563);
and U5458 (N_5458,N_4711,N_4047);
or U5459 (N_5459,N_4498,N_4788);
xnor U5460 (N_5460,N_4683,N_4169);
nand U5461 (N_5461,N_4735,N_4026);
and U5462 (N_5462,N_4941,N_4135);
nor U5463 (N_5463,N_4108,N_4587);
and U5464 (N_5464,N_4797,N_4125);
nand U5465 (N_5465,N_4352,N_4028);
nand U5466 (N_5466,N_4608,N_4344);
xnor U5467 (N_5467,N_4328,N_4284);
or U5468 (N_5468,N_4836,N_4252);
nand U5469 (N_5469,N_4021,N_4322);
nor U5470 (N_5470,N_4248,N_4614);
xor U5471 (N_5471,N_4691,N_4231);
or U5472 (N_5472,N_4932,N_4146);
xnor U5473 (N_5473,N_4803,N_4649);
xnor U5474 (N_5474,N_4678,N_4495);
or U5475 (N_5475,N_4131,N_4194);
or U5476 (N_5476,N_4929,N_4770);
nor U5477 (N_5477,N_4089,N_4520);
and U5478 (N_5478,N_4383,N_4774);
nand U5479 (N_5479,N_4030,N_4791);
nand U5480 (N_5480,N_4723,N_4925);
or U5481 (N_5481,N_4330,N_4124);
nand U5482 (N_5482,N_4424,N_4641);
and U5483 (N_5483,N_4856,N_4456);
and U5484 (N_5484,N_4927,N_4718);
nand U5485 (N_5485,N_4087,N_4654);
nor U5486 (N_5486,N_4487,N_4001);
nor U5487 (N_5487,N_4329,N_4072);
nand U5488 (N_5488,N_4313,N_4164);
or U5489 (N_5489,N_4122,N_4133);
and U5490 (N_5490,N_4810,N_4915);
xnor U5491 (N_5491,N_4341,N_4874);
nand U5492 (N_5492,N_4040,N_4421);
nand U5493 (N_5493,N_4406,N_4946);
or U5494 (N_5494,N_4218,N_4817);
nand U5495 (N_5495,N_4174,N_4478);
or U5496 (N_5496,N_4324,N_4732);
or U5497 (N_5497,N_4979,N_4843);
or U5498 (N_5498,N_4750,N_4375);
or U5499 (N_5499,N_4902,N_4210);
and U5500 (N_5500,N_4318,N_4186);
nor U5501 (N_5501,N_4468,N_4787);
or U5502 (N_5502,N_4637,N_4397);
nor U5503 (N_5503,N_4079,N_4061);
nand U5504 (N_5504,N_4769,N_4027);
nand U5505 (N_5505,N_4912,N_4545);
xor U5506 (N_5506,N_4304,N_4281);
xnor U5507 (N_5507,N_4134,N_4948);
nand U5508 (N_5508,N_4574,N_4211);
xor U5509 (N_5509,N_4744,N_4778);
xor U5510 (N_5510,N_4347,N_4061);
and U5511 (N_5511,N_4740,N_4881);
nand U5512 (N_5512,N_4573,N_4709);
or U5513 (N_5513,N_4719,N_4355);
nand U5514 (N_5514,N_4304,N_4235);
and U5515 (N_5515,N_4369,N_4536);
nor U5516 (N_5516,N_4104,N_4756);
and U5517 (N_5517,N_4011,N_4604);
and U5518 (N_5518,N_4102,N_4751);
or U5519 (N_5519,N_4039,N_4674);
or U5520 (N_5520,N_4733,N_4164);
xor U5521 (N_5521,N_4194,N_4394);
and U5522 (N_5522,N_4871,N_4181);
nand U5523 (N_5523,N_4437,N_4887);
xnor U5524 (N_5524,N_4606,N_4793);
xor U5525 (N_5525,N_4063,N_4139);
nor U5526 (N_5526,N_4871,N_4684);
nand U5527 (N_5527,N_4835,N_4211);
nand U5528 (N_5528,N_4096,N_4321);
and U5529 (N_5529,N_4416,N_4724);
nor U5530 (N_5530,N_4680,N_4311);
nand U5531 (N_5531,N_4747,N_4523);
nand U5532 (N_5532,N_4761,N_4375);
nor U5533 (N_5533,N_4021,N_4765);
nor U5534 (N_5534,N_4482,N_4309);
xnor U5535 (N_5535,N_4161,N_4014);
xor U5536 (N_5536,N_4298,N_4838);
nor U5537 (N_5537,N_4513,N_4139);
nor U5538 (N_5538,N_4378,N_4128);
and U5539 (N_5539,N_4309,N_4155);
xor U5540 (N_5540,N_4289,N_4279);
xor U5541 (N_5541,N_4950,N_4904);
or U5542 (N_5542,N_4734,N_4865);
nor U5543 (N_5543,N_4921,N_4986);
and U5544 (N_5544,N_4291,N_4406);
nand U5545 (N_5545,N_4682,N_4341);
xnor U5546 (N_5546,N_4353,N_4279);
xnor U5547 (N_5547,N_4969,N_4424);
and U5548 (N_5548,N_4406,N_4188);
or U5549 (N_5549,N_4714,N_4062);
nand U5550 (N_5550,N_4526,N_4397);
nand U5551 (N_5551,N_4215,N_4633);
nand U5552 (N_5552,N_4783,N_4457);
or U5553 (N_5553,N_4396,N_4774);
xnor U5554 (N_5554,N_4163,N_4987);
or U5555 (N_5555,N_4191,N_4109);
or U5556 (N_5556,N_4079,N_4285);
nand U5557 (N_5557,N_4234,N_4131);
or U5558 (N_5558,N_4482,N_4859);
nand U5559 (N_5559,N_4269,N_4726);
nand U5560 (N_5560,N_4524,N_4678);
and U5561 (N_5561,N_4780,N_4917);
and U5562 (N_5562,N_4781,N_4919);
xnor U5563 (N_5563,N_4481,N_4233);
xnor U5564 (N_5564,N_4246,N_4106);
nand U5565 (N_5565,N_4187,N_4815);
xnor U5566 (N_5566,N_4459,N_4223);
nand U5567 (N_5567,N_4768,N_4067);
nor U5568 (N_5568,N_4728,N_4832);
nor U5569 (N_5569,N_4634,N_4682);
or U5570 (N_5570,N_4452,N_4184);
or U5571 (N_5571,N_4140,N_4135);
nand U5572 (N_5572,N_4551,N_4423);
and U5573 (N_5573,N_4455,N_4152);
or U5574 (N_5574,N_4833,N_4282);
or U5575 (N_5575,N_4343,N_4584);
xor U5576 (N_5576,N_4914,N_4700);
or U5577 (N_5577,N_4485,N_4745);
and U5578 (N_5578,N_4942,N_4616);
nand U5579 (N_5579,N_4861,N_4869);
or U5580 (N_5580,N_4105,N_4890);
nor U5581 (N_5581,N_4379,N_4866);
or U5582 (N_5582,N_4381,N_4839);
nand U5583 (N_5583,N_4827,N_4616);
xor U5584 (N_5584,N_4826,N_4995);
nand U5585 (N_5585,N_4549,N_4556);
or U5586 (N_5586,N_4263,N_4159);
and U5587 (N_5587,N_4870,N_4228);
nand U5588 (N_5588,N_4958,N_4117);
xor U5589 (N_5589,N_4646,N_4596);
or U5590 (N_5590,N_4135,N_4093);
xnor U5591 (N_5591,N_4453,N_4107);
nor U5592 (N_5592,N_4670,N_4721);
nand U5593 (N_5593,N_4264,N_4956);
or U5594 (N_5594,N_4235,N_4749);
nand U5595 (N_5595,N_4007,N_4537);
or U5596 (N_5596,N_4137,N_4446);
xor U5597 (N_5597,N_4478,N_4872);
xnor U5598 (N_5598,N_4604,N_4398);
nand U5599 (N_5599,N_4448,N_4998);
xnor U5600 (N_5600,N_4634,N_4685);
nand U5601 (N_5601,N_4165,N_4733);
or U5602 (N_5602,N_4833,N_4246);
or U5603 (N_5603,N_4082,N_4254);
nand U5604 (N_5604,N_4480,N_4631);
nand U5605 (N_5605,N_4753,N_4149);
nor U5606 (N_5606,N_4846,N_4847);
nand U5607 (N_5607,N_4942,N_4387);
nand U5608 (N_5608,N_4099,N_4152);
or U5609 (N_5609,N_4684,N_4378);
nand U5610 (N_5610,N_4231,N_4334);
nor U5611 (N_5611,N_4579,N_4656);
or U5612 (N_5612,N_4280,N_4788);
nand U5613 (N_5613,N_4728,N_4368);
nor U5614 (N_5614,N_4222,N_4423);
and U5615 (N_5615,N_4945,N_4002);
xnor U5616 (N_5616,N_4111,N_4861);
nor U5617 (N_5617,N_4233,N_4867);
nor U5618 (N_5618,N_4690,N_4559);
xnor U5619 (N_5619,N_4328,N_4320);
and U5620 (N_5620,N_4061,N_4699);
and U5621 (N_5621,N_4259,N_4598);
and U5622 (N_5622,N_4045,N_4396);
nand U5623 (N_5623,N_4839,N_4316);
nand U5624 (N_5624,N_4334,N_4513);
and U5625 (N_5625,N_4222,N_4783);
xnor U5626 (N_5626,N_4638,N_4523);
or U5627 (N_5627,N_4254,N_4358);
nor U5628 (N_5628,N_4801,N_4439);
nand U5629 (N_5629,N_4754,N_4076);
nor U5630 (N_5630,N_4499,N_4677);
and U5631 (N_5631,N_4364,N_4103);
xnor U5632 (N_5632,N_4940,N_4387);
and U5633 (N_5633,N_4441,N_4392);
and U5634 (N_5634,N_4787,N_4824);
xnor U5635 (N_5635,N_4671,N_4620);
xor U5636 (N_5636,N_4977,N_4604);
and U5637 (N_5637,N_4930,N_4407);
or U5638 (N_5638,N_4893,N_4947);
and U5639 (N_5639,N_4158,N_4471);
nor U5640 (N_5640,N_4718,N_4845);
nor U5641 (N_5641,N_4484,N_4029);
and U5642 (N_5642,N_4844,N_4922);
nor U5643 (N_5643,N_4568,N_4487);
nor U5644 (N_5644,N_4023,N_4067);
xnor U5645 (N_5645,N_4808,N_4101);
and U5646 (N_5646,N_4196,N_4955);
and U5647 (N_5647,N_4687,N_4225);
nand U5648 (N_5648,N_4746,N_4435);
xor U5649 (N_5649,N_4303,N_4544);
or U5650 (N_5650,N_4178,N_4121);
xor U5651 (N_5651,N_4265,N_4746);
nand U5652 (N_5652,N_4128,N_4380);
nor U5653 (N_5653,N_4486,N_4201);
nor U5654 (N_5654,N_4505,N_4163);
or U5655 (N_5655,N_4426,N_4524);
nand U5656 (N_5656,N_4867,N_4009);
or U5657 (N_5657,N_4789,N_4157);
or U5658 (N_5658,N_4911,N_4040);
nand U5659 (N_5659,N_4188,N_4796);
nor U5660 (N_5660,N_4777,N_4933);
nand U5661 (N_5661,N_4616,N_4595);
nor U5662 (N_5662,N_4943,N_4243);
nor U5663 (N_5663,N_4338,N_4349);
nor U5664 (N_5664,N_4338,N_4732);
or U5665 (N_5665,N_4417,N_4324);
and U5666 (N_5666,N_4233,N_4683);
nor U5667 (N_5667,N_4265,N_4784);
and U5668 (N_5668,N_4548,N_4291);
nor U5669 (N_5669,N_4925,N_4206);
xor U5670 (N_5670,N_4134,N_4727);
or U5671 (N_5671,N_4509,N_4124);
and U5672 (N_5672,N_4786,N_4821);
nor U5673 (N_5673,N_4937,N_4330);
xnor U5674 (N_5674,N_4093,N_4553);
nand U5675 (N_5675,N_4834,N_4582);
nand U5676 (N_5676,N_4703,N_4172);
nand U5677 (N_5677,N_4944,N_4735);
and U5678 (N_5678,N_4679,N_4733);
nand U5679 (N_5679,N_4402,N_4514);
xnor U5680 (N_5680,N_4312,N_4194);
or U5681 (N_5681,N_4127,N_4637);
nor U5682 (N_5682,N_4182,N_4179);
nand U5683 (N_5683,N_4148,N_4255);
and U5684 (N_5684,N_4116,N_4614);
xor U5685 (N_5685,N_4730,N_4988);
and U5686 (N_5686,N_4116,N_4421);
nor U5687 (N_5687,N_4831,N_4256);
and U5688 (N_5688,N_4676,N_4225);
nor U5689 (N_5689,N_4500,N_4025);
xnor U5690 (N_5690,N_4414,N_4228);
and U5691 (N_5691,N_4771,N_4200);
xnor U5692 (N_5692,N_4521,N_4230);
nand U5693 (N_5693,N_4068,N_4360);
xnor U5694 (N_5694,N_4960,N_4228);
nor U5695 (N_5695,N_4178,N_4182);
and U5696 (N_5696,N_4222,N_4767);
nand U5697 (N_5697,N_4322,N_4825);
xnor U5698 (N_5698,N_4574,N_4417);
nand U5699 (N_5699,N_4651,N_4238);
and U5700 (N_5700,N_4853,N_4850);
nand U5701 (N_5701,N_4966,N_4247);
and U5702 (N_5702,N_4962,N_4223);
nand U5703 (N_5703,N_4467,N_4070);
nand U5704 (N_5704,N_4263,N_4287);
nand U5705 (N_5705,N_4413,N_4346);
and U5706 (N_5706,N_4655,N_4915);
nand U5707 (N_5707,N_4129,N_4539);
or U5708 (N_5708,N_4309,N_4369);
nand U5709 (N_5709,N_4405,N_4046);
and U5710 (N_5710,N_4507,N_4509);
nor U5711 (N_5711,N_4052,N_4251);
and U5712 (N_5712,N_4329,N_4008);
nor U5713 (N_5713,N_4860,N_4088);
nor U5714 (N_5714,N_4713,N_4459);
xor U5715 (N_5715,N_4213,N_4717);
nand U5716 (N_5716,N_4121,N_4580);
xnor U5717 (N_5717,N_4968,N_4034);
nor U5718 (N_5718,N_4505,N_4412);
and U5719 (N_5719,N_4805,N_4233);
xnor U5720 (N_5720,N_4210,N_4252);
nand U5721 (N_5721,N_4987,N_4119);
and U5722 (N_5722,N_4258,N_4108);
and U5723 (N_5723,N_4486,N_4939);
and U5724 (N_5724,N_4042,N_4154);
xor U5725 (N_5725,N_4236,N_4657);
nor U5726 (N_5726,N_4877,N_4070);
nand U5727 (N_5727,N_4443,N_4499);
and U5728 (N_5728,N_4317,N_4929);
xor U5729 (N_5729,N_4130,N_4294);
and U5730 (N_5730,N_4086,N_4771);
nand U5731 (N_5731,N_4356,N_4630);
or U5732 (N_5732,N_4515,N_4647);
or U5733 (N_5733,N_4446,N_4262);
or U5734 (N_5734,N_4294,N_4587);
and U5735 (N_5735,N_4324,N_4413);
or U5736 (N_5736,N_4321,N_4050);
and U5737 (N_5737,N_4584,N_4021);
or U5738 (N_5738,N_4080,N_4569);
nand U5739 (N_5739,N_4449,N_4931);
nor U5740 (N_5740,N_4812,N_4390);
or U5741 (N_5741,N_4644,N_4279);
xor U5742 (N_5742,N_4316,N_4600);
nor U5743 (N_5743,N_4558,N_4268);
xnor U5744 (N_5744,N_4785,N_4924);
and U5745 (N_5745,N_4016,N_4208);
and U5746 (N_5746,N_4592,N_4427);
nor U5747 (N_5747,N_4483,N_4259);
or U5748 (N_5748,N_4662,N_4126);
nand U5749 (N_5749,N_4826,N_4948);
nor U5750 (N_5750,N_4201,N_4475);
nor U5751 (N_5751,N_4129,N_4032);
nor U5752 (N_5752,N_4853,N_4771);
nor U5753 (N_5753,N_4670,N_4057);
and U5754 (N_5754,N_4318,N_4945);
nor U5755 (N_5755,N_4295,N_4592);
xnor U5756 (N_5756,N_4805,N_4130);
nor U5757 (N_5757,N_4849,N_4117);
nor U5758 (N_5758,N_4187,N_4117);
nand U5759 (N_5759,N_4163,N_4696);
nand U5760 (N_5760,N_4394,N_4338);
nand U5761 (N_5761,N_4316,N_4752);
and U5762 (N_5762,N_4836,N_4872);
and U5763 (N_5763,N_4360,N_4065);
xor U5764 (N_5764,N_4465,N_4860);
and U5765 (N_5765,N_4324,N_4064);
xor U5766 (N_5766,N_4335,N_4520);
nand U5767 (N_5767,N_4701,N_4382);
xnor U5768 (N_5768,N_4057,N_4855);
or U5769 (N_5769,N_4307,N_4969);
or U5770 (N_5770,N_4170,N_4632);
nor U5771 (N_5771,N_4628,N_4448);
xnor U5772 (N_5772,N_4920,N_4292);
xnor U5773 (N_5773,N_4300,N_4310);
or U5774 (N_5774,N_4395,N_4027);
xnor U5775 (N_5775,N_4848,N_4093);
nor U5776 (N_5776,N_4860,N_4351);
nor U5777 (N_5777,N_4918,N_4158);
nand U5778 (N_5778,N_4067,N_4291);
nand U5779 (N_5779,N_4638,N_4571);
xor U5780 (N_5780,N_4958,N_4623);
xnor U5781 (N_5781,N_4405,N_4619);
and U5782 (N_5782,N_4487,N_4689);
nand U5783 (N_5783,N_4119,N_4574);
and U5784 (N_5784,N_4921,N_4559);
or U5785 (N_5785,N_4782,N_4386);
nor U5786 (N_5786,N_4494,N_4831);
xor U5787 (N_5787,N_4314,N_4788);
nand U5788 (N_5788,N_4933,N_4398);
or U5789 (N_5789,N_4929,N_4839);
nand U5790 (N_5790,N_4497,N_4701);
nand U5791 (N_5791,N_4194,N_4088);
nand U5792 (N_5792,N_4888,N_4070);
xnor U5793 (N_5793,N_4253,N_4248);
nand U5794 (N_5794,N_4717,N_4625);
xor U5795 (N_5795,N_4238,N_4092);
nor U5796 (N_5796,N_4579,N_4945);
nor U5797 (N_5797,N_4786,N_4269);
nand U5798 (N_5798,N_4255,N_4212);
xor U5799 (N_5799,N_4907,N_4523);
nor U5800 (N_5800,N_4325,N_4422);
nor U5801 (N_5801,N_4558,N_4853);
xor U5802 (N_5802,N_4225,N_4510);
and U5803 (N_5803,N_4187,N_4512);
nand U5804 (N_5804,N_4525,N_4355);
xor U5805 (N_5805,N_4837,N_4464);
and U5806 (N_5806,N_4013,N_4113);
xor U5807 (N_5807,N_4274,N_4332);
nor U5808 (N_5808,N_4783,N_4366);
xnor U5809 (N_5809,N_4230,N_4706);
nand U5810 (N_5810,N_4717,N_4344);
nor U5811 (N_5811,N_4903,N_4991);
or U5812 (N_5812,N_4415,N_4876);
or U5813 (N_5813,N_4439,N_4724);
nand U5814 (N_5814,N_4309,N_4811);
and U5815 (N_5815,N_4627,N_4056);
or U5816 (N_5816,N_4665,N_4092);
and U5817 (N_5817,N_4687,N_4192);
or U5818 (N_5818,N_4119,N_4792);
nand U5819 (N_5819,N_4265,N_4425);
nor U5820 (N_5820,N_4180,N_4734);
or U5821 (N_5821,N_4160,N_4107);
or U5822 (N_5822,N_4797,N_4327);
nand U5823 (N_5823,N_4619,N_4955);
xor U5824 (N_5824,N_4783,N_4173);
xnor U5825 (N_5825,N_4321,N_4039);
xor U5826 (N_5826,N_4898,N_4832);
or U5827 (N_5827,N_4167,N_4425);
or U5828 (N_5828,N_4116,N_4484);
and U5829 (N_5829,N_4923,N_4881);
nor U5830 (N_5830,N_4549,N_4871);
or U5831 (N_5831,N_4974,N_4885);
and U5832 (N_5832,N_4952,N_4378);
nand U5833 (N_5833,N_4926,N_4327);
and U5834 (N_5834,N_4937,N_4513);
and U5835 (N_5835,N_4642,N_4876);
nor U5836 (N_5836,N_4527,N_4764);
and U5837 (N_5837,N_4630,N_4747);
and U5838 (N_5838,N_4383,N_4151);
or U5839 (N_5839,N_4122,N_4113);
nor U5840 (N_5840,N_4396,N_4282);
nand U5841 (N_5841,N_4268,N_4786);
xor U5842 (N_5842,N_4873,N_4246);
or U5843 (N_5843,N_4519,N_4866);
nand U5844 (N_5844,N_4914,N_4364);
nor U5845 (N_5845,N_4347,N_4014);
nand U5846 (N_5846,N_4544,N_4503);
or U5847 (N_5847,N_4994,N_4843);
nand U5848 (N_5848,N_4481,N_4421);
and U5849 (N_5849,N_4346,N_4401);
nor U5850 (N_5850,N_4705,N_4900);
xor U5851 (N_5851,N_4139,N_4943);
or U5852 (N_5852,N_4932,N_4807);
or U5853 (N_5853,N_4728,N_4608);
nor U5854 (N_5854,N_4333,N_4349);
and U5855 (N_5855,N_4676,N_4617);
or U5856 (N_5856,N_4393,N_4463);
nand U5857 (N_5857,N_4868,N_4698);
or U5858 (N_5858,N_4932,N_4227);
or U5859 (N_5859,N_4578,N_4254);
xor U5860 (N_5860,N_4273,N_4727);
nand U5861 (N_5861,N_4609,N_4932);
and U5862 (N_5862,N_4474,N_4004);
xor U5863 (N_5863,N_4775,N_4432);
or U5864 (N_5864,N_4863,N_4423);
nand U5865 (N_5865,N_4342,N_4383);
xnor U5866 (N_5866,N_4541,N_4757);
xnor U5867 (N_5867,N_4163,N_4734);
nor U5868 (N_5868,N_4507,N_4495);
nand U5869 (N_5869,N_4904,N_4707);
nand U5870 (N_5870,N_4664,N_4985);
or U5871 (N_5871,N_4634,N_4128);
nand U5872 (N_5872,N_4575,N_4267);
or U5873 (N_5873,N_4257,N_4278);
nor U5874 (N_5874,N_4520,N_4138);
or U5875 (N_5875,N_4345,N_4412);
xnor U5876 (N_5876,N_4535,N_4564);
and U5877 (N_5877,N_4504,N_4937);
xnor U5878 (N_5878,N_4400,N_4880);
xnor U5879 (N_5879,N_4822,N_4065);
and U5880 (N_5880,N_4815,N_4537);
nor U5881 (N_5881,N_4403,N_4676);
xor U5882 (N_5882,N_4020,N_4382);
or U5883 (N_5883,N_4696,N_4203);
nand U5884 (N_5884,N_4146,N_4828);
nand U5885 (N_5885,N_4255,N_4815);
and U5886 (N_5886,N_4229,N_4319);
nand U5887 (N_5887,N_4979,N_4902);
nor U5888 (N_5888,N_4454,N_4486);
or U5889 (N_5889,N_4979,N_4390);
nor U5890 (N_5890,N_4438,N_4902);
nor U5891 (N_5891,N_4689,N_4287);
xnor U5892 (N_5892,N_4098,N_4921);
nand U5893 (N_5893,N_4138,N_4788);
xor U5894 (N_5894,N_4293,N_4218);
and U5895 (N_5895,N_4963,N_4795);
nor U5896 (N_5896,N_4434,N_4769);
and U5897 (N_5897,N_4826,N_4889);
or U5898 (N_5898,N_4320,N_4702);
nand U5899 (N_5899,N_4540,N_4828);
nand U5900 (N_5900,N_4312,N_4062);
or U5901 (N_5901,N_4018,N_4725);
xnor U5902 (N_5902,N_4794,N_4951);
or U5903 (N_5903,N_4841,N_4077);
nand U5904 (N_5904,N_4835,N_4561);
nand U5905 (N_5905,N_4625,N_4211);
nor U5906 (N_5906,N_4406,N_4373);
nor U5907 (N_5907,N_4812,N_4717);
xor U5908 (N_5908,N_4103,N_4647);
nand U5909 (N_5909,N_4595,N_4669);
xor U5910 (N_5910,N_4829,N_4477);
nor U5911 (N_5911,N_4829,N_4097);
xor U5912 (N_5912,N_4179,N_4091);
and U5913 (N_5913,N_4211,N_4395);
nor U5914 (N_5914,N_4871,N_4693);
and U5915 (N_5915,N_4034,N_4189);
or U5916 (N_5916,N_4154,N_4120);
and U5917 (N_5917,N_4251,N_4539);
or U5918 (N_5918,N_4427,N_4231);
and U5919 (N_5919,N_4444,N_4088);
and U5920 (N_5920,N_4297,N_4066);
nor U5921 (N_5921,N_4268,N_4607);
xnor U5922 (N_5922,N_4374,N_4563);
or U5923 (N_5923,N_4985,N_4626);
xor U5924 (N_5924,N_4994,N_4816);
and U5925 (N_5925,N_4573,N_4546);
and U5926 (N_5926,N_4010,N_4267);
xor U5927 (N_5927,N_4029,N_4422);
nand U5928 (N_5928,N_4660,N_4992);
nor U5929 (N_5929,N_4639,N_4822);
nand U5930 (N_5930,N_4346,N_4482);
nor U5931 (N_5931,N_4168,N_4791);
nor U5932 (N_5932,N_4699,N_4825);
nand U5933 (N_5933,N_4235,N_4525);
xor U5934 (N_5934,N_4767,N_4162);
nand U5935 (N_5935,N_4958,N_4027);
and U5936 (N_5936,N_4409,N_4236);
nor U5937 (N_5937,N_4492,N_4771);
and U5938 (N_5938,N_4241,N_4297);
nand U5939 (N_5939,N_4277,N_4827);
or U5940 (N_5940,N_4259,N_4107);
and U5941 (N_5941,N_4003,N_4516);
and U5942 (N_5942,N_4603,N_4026);
xnor U5943 (N_5943,N_4802,N_4215);
xor U5944 (N_5944,N_4080,N_4554);
and U5945 (N_5945,N_4016,N_4465);
nor U5946 (N_5946,N_4121,N_4684);
xnor U5947 (N_5947,N_4591,N_4910);
nor U5948 (N_5948,N_4116,N_4758);
nor U5949 (N_5949,N_4781,N_4577);
and U5950 (N_5950,N_4503,N_4648);
and U5951 (N_5951,N_4602,N_4172);
xnor U5952 (N_5952,N_4301,N_4476);
and U5953 (N_5953,N_4337,N_4527);
and U5954 (N_5954,N_4585,N_4247);
nor U5955 (N_5955,N_4737,N_4897);
nor U5956 (N_5956,N_4232,N_4082);
xor U5957 (N_5957,N_4213,N_4856);
nor U5958 (N_5958,N_4827,N_4313);
and U5959 (N_5959,N_4929,N_4006);
nor U5960 (N_5960,N_4852,N_4385);
or U5961 (N_5961,N_4152,N_4228);
xor U5962 (N_5962,N_4517,N_4806);
and U5963 (N_5963,N_4597,N_4495);
and U5964 (N_5964,N_4941,N_4799);
or U5965 (N_5965,N_4834,N_4616);
nor U5966 (N_5966,N_4510,N_4168);
and U5967 (N_5967,N_4508,N_4316);
and U5968 (N_5968,N_4818,N_4001);
nor U5969 (N_5969,N_4501,N_4502);
nor U5970 (N_5970,N_4229,N_4049);
and U5971 (N_5971,N_4757,N_4918);
nor U5972 (N_5972,N_4832,N_4913);
and U5973 (N_5973,N_4342,N_4576);
and U5974 (N_5974,N_4888,N_4177);
or U5975 (N_5975,N_4526,N_4035);
xnor U5976 (N_5976,N_4162,N_4584);
nor U5977 (N_5977,N_4533,N_4464);
nand U5978 (N_5978,N_4972,N_4279);
or U5979 (N_5979,N_4869,N_4699);
nand U5980 (N_5980,N_4307,N_4632);
or U5981 (N_5981,N_4216,N_4830);
or U5982 (N_5982,N_4092,N_4370);
xnor U5983 (N_5983,N_4957,N_4256);
nor U5984 (N_5984,N_4826,N_4201);
nor U5985 (N_5985,N_4829,N_4884);
and U5986 (N_5986,N_4607,N_4423);
xor U5987 (N_5987,N_4155,N_4116);
xor U5988 (N_5988,N_4190,N_4120);
nand U5989 (N_5989,N_4627,N_4814);
and U5990 (N_5990,N_4660,N_4354);
or U5991 (N_5991,N_4836,N_4785);
and U5992 (N_5992,N_4512,N_4001);
nor U5993 (N_5993,N_4986,N_4217);
nor U5994 (N_5994,N_4662,N_4828);
or U5995 (N_5995,N_4951,N_4932);
xnor U5996 (N_5996,N_4477,N_4399);
and U5997 (N_5997,N_4318,N_4108);
or U5998 (N_5998,N_4866,N_4370);
or U5999 (N_5999,N_4334,N_4309);
and U6000 (N_6000,N_5376,N_5794);
xor U6001 (N_6001,N_5296,N_5931);
or U6002 (N_6002,N_5907,N_5530);
nor U6003 (N_6003,N_5825,N_5326);
and U6004 (N_6004,N_5954,N_5335);
and U6005 (N_6005,N_5166,N_5743);
and U6006 (N_6006,N_5348,N_5320);
and U6007 (N_6007,N_5725,N_5570);
and U6008 (N_6008,N_5845,N_5992);
and U6009 (N_6009,N_5361,N_5585);
or U6010 (N_6010,N_5473,N_5742);
xnor U6011 (N_6011,N_5556,N_5922);
nor U6012 (N_6012,N_5325,N_5112);
nor U6013 (N_6013,N_5155,N_5211);
xor U6014 (N_6014,N_5067,N_5905);
nand U6015 (N_6015,N_5417,N_5766);
or U6016 (N_6016,N_5430,N_5612);
nor U6017 (N_6017,N_5968,N_5105);
xnor U6018 (N_6018,N_5672,N_5757);
nor U6019 (N_6019,N_5765,N_5664);
xor U6020 (N_6020,N_5700,N_5862);
and U6021 (N_6021,N_5269,N_5812);
xor U6022 (N_6022,N_5983,N_5520);
nor U6023 (N_6023,N_5486,N_5649);
xor U6024 (N_6024,N_5314,N_5303);
or U6025 (N_6025,N_5752,N_5493);
nand U6026 (N_6026,N_5912,N_5744);
xor U6027 (N_6027,N_5746,N_5514);
and U6028 (N_6028,N_5178,N_5481);
nand U6029 (N_6029,N_5265,N_5138);
and U6030 (N_6030,N_5604,N_5057);
and U6031 (N_6031,N_5301,N_5893);
nor U6032 (N_6032,N_5411,N_5975);
nand U6033 (N_6033,N_5060,N_5627);
and U6034 (N_6034,N_5892,N_5786);
nor U6035 (N_6035,N_5690,N_5216);
nand U6036 (N_6036,N_5559,N_5891);
xor U6037 (N_6037,N_5973,N_5441);
or U6038 (N_6038,N_5226,N_5637);
xor U6039 (N_6039,N_5307,N_5807);
and U6040 (N_6040,N_5680,N_5151);
or U6041 (N_6041,N_5222,N_5251);
xnor U6042 (N_6042,N_5182,N_5305);
xor U6043 (N_6043,N_5580,N_5568);
nor U6044 (N_6044,N_5756,N_5927);
nor U6045 (N_6045,N_5154,N_5542);
nand U6046 (N_6046,N_5780,N_5404);
or U6047 (N_6047,N_5477,N_5191);
nand U6048 (N_6048,N_5978,N_5260);
or U6049 (N_6049,N_5084,N_5176);
xnor U6050 (N_6050,N_5229,N_5450);
nand U6051 (N_6051,N_5609,N_5037);
or U6052 (N_6052,N_5819,N_5820);
or U6053 (N_6053,N_5491,N_5662);
xnor U6054 (N_6054,N_5099,N_5942);
and U6055 (N_6055,N_5435,N_5209);
and U6056 (N_6056,N_5342,N_5101);
and U6057 (N_6057,N_5340,N_5703);
or U6058 (N_6058,N_5242,N_5088);
nor U6059 (N_6059,N_5377,N_5434);
xor U6060 (N_6060,N_5162,N_5352);
nand U6061 (N_6061,N_5152,N_5076);
nand U6062 (N_6062,N_5599,N_5136);
nor U6063 (N_6063,N_5413,N_5082);
or U6064 (N_6064,N_5180,N_5605);
xor U6065 (N_6065,N_5480,N_5564);
or U6066 (N_6066,N_5402,N_5839);
nand U6067 (N_6067,N_5522,N_5210);
and U6068 (N_6068,N_5939,N_5512);
xor U6069 (N_6069,N_5643,N_5697);
nor U6070 (N_6070,N_5165,N_5333);
xnor U6071 (N_6071,N_5338,N_5691);
nor U6072 (N_6072,N_5050,N_5842);
and U6073 (N_6073,N_5941,N_5550);
nor U6074 (N_6074,N_5295,N_5192);
nor U6075 (N_6075,N_5863,N_5663);
nand U6076 (N_6076,N_5218,N_5231);
nand U6077 (N_6077,N_5114,N_5901);
and U6078 (N_6078,N_5408,N_5317);
and U6079 (N_6079,N_5124,N_5925);
xnor U6080 (N_6080,N_5339,N_5537);
nor U6081 (N_6081,N_5444,N_5039);
or U6082 (N_6082,N_5715,N_5988);
nand U6083 (N_6083,N_5017,N_5647);
xor U6084 (N_6084,N_5056,N_5517);
nand U6085 (N_6085,N_5745,N_5908);
or U6086 (N_6086,N_5967,N_5671);
xnor U6087 (N_6087,N_5618,N_5467);
nor U6088 (N_6088,N_5699,N_5019);
xnor U6089 (N_6089,N_5915,N_5897);
xor U6090 (N_6090,N_5816,N_5916);
xor U6091 (N_6091,N_5658,N_5137);
or U6092 (N_6092,N_5418,N_5737);
nor U6093 (N_6093,N_5379,N_5791);
and U6094 (N_6094,N_5667,N_5634);
or U6095 (N_6095,N_5783,N_5249);
nand U6096 (N_6096,N_5610,N_5072);
nor U6097 (N_6097,N_5372,N_5148);
nor U6098 (N_6098,N_5334,N_5704);
and U6099 (N_6099,N_5494,N_5598);
or U6100 (N_6100,N_5661,N_5507);
xnor U6101 (N_6101,N_5062,N_5886);
and U6102 (N_6102,N_5217,N_5052);
nor U6103 (N_6103,N_5426,N_5692);
and U6104 (N_6104,N_5669,N_5923);
or U6105 (N_6105,N_5346,N_5287);
nand U6106 (N_6106,N_5038,N_5075);
or U6107 (N_6107,N_5852,N_5068);
and U6108 (N_6108,N_5194,N_5563);
and U6109 (N_6109,N_5410,N_5804);
nor U6110 (N_6110,N_5013,N_5471);
and U6111 (N_6111,N_5767,N_5063);
nor U6112 (N_6112,N_5048,N_5469);
nor U6113 (N_6113,N_5183,N_5321);
and U6114 (N_6114,N_5866,N_5518);
or U6115 (N_6115,N_5960,N_5091);
nor U6116 (N_6116,N_5904,N_5523);
nand U6117 (N_6117,N_5382,N_5140);
and U6118 (N_6118,N_5130,N_5965);
and U6119 (N_6119,N_5508,N_5841);
xnor U6120 (N_6120,N_5100,N_5574);
xnor U6121 (N_6121,N_5133,N_5813);
nand U6122 (N_6122,N_5538,N_5531);
xor U6123 (N_6123,N_5738,N_5781);
and U6124 (N_6124,N_5490,N_5318);
nand U6125 (N_6125,N_5511,N_5393);
nor U6126 (N_6126,N_5438,N_5007);
or U6127 (N_6127,N_5289,N_5142);
or U6128 (N_6128,N_5423,N_5840);
nand U6129 (N_6129,N_5844,N_5645);
xnor U6130 (N_6130,N_5732,N_5449);
nor U6131 (N_6131,N_5122,N_5716);
and U6132 (N_6132,N_5364,N_5985);
or U6133 (N_6133,N_5870,N_5392);
or U6134 (N_6134,N_5546,N_5628);
and U6135 (N_6135,N_5115,N_5261);
or U6136 (N_6136,N_5108,N_5758);
xnor U6137 (N_6137,N_5505,N_5003);
nor U6138 (N_6138,N_5278,N_5665);
or U6139 (N_6139,N_5991,N_5555);
or U6140 (N_6140,N_5407,N_5689);
and U6141 (N_6141,N_5833,N_5920);
or U6142 (N_6142,N_5759,N_5624);
nor U6143 (N_6143,N_5044,N_5143);
xnor U6144 (N_6144,N_5219,N_5843);
nand U6145 (N_6145,N_5461,N_5502);
xor U6146 (N_6146,N_5214,N_5323);
nand U6147 (N_6147,N_5932,N_5458);
xnor U6148 (N_6148,N_5189,N_5810);
nand U6149 (N_6149,N_5644,N_5104);
nor U6150 (N_6150,N_5388,N_5808);
and U6151 (N_6151,N_5824,N_5313);
or U6152 (N_6152,N_5846,N_5046);
or U6153 (N_6153,N_5240,N_5969);
or U6154 (N_6154,N_5011,N_5830);
nand U6155 (N_6155,N_5943,N_5077);
xor U6156 (N_6156,N_5371,N_5771);
xor U6157 (N_6157,N_5127,N_5120);
or U6158 (N_6158,N_5509,N_5298);
nor U6159 (N_6159,N_5341,N_5254);
xnor U6160 (N_6160,N_5874,N_5888);
nand U6161 (N_6161,N_5685,N_5113);
nand U6162 (N_6162,N_5970,N_5118);
xnor U6163 (N_6163,N_5020,N_5462);
or U6164 (N_6164,N_5391,N_5974);
or U6165 (N_6165,N_5872,N_5573);
and U6166 (N_6166,N_5638,N_5468);
nor U6167 (N_6167,N_5395,N_5859);
and U6168 (N_6168,N_5709,N_5456);
nand U6169 (N_6169,N_5749,N_5906);
and U6170 (N_6170,N_5607,N_5919);
xnor U6171 (N_6171,N_5253,N_5894);
nor U6172 (N_6172,N_5561,N_5476);
xor U6173 (N_6173,N_5951,N_5398);
and U6174 (N_6174,N_5110,N_5149);
and U6175 (N_6175,N_5995,N_5729);
xor U6176 (N_6176,N_5762,N_5054);
xnor U6177 (N_6177,N_5596,N_5986);
xnor U6178 (N_6178,N_5173,N_5717);
or U6179 (N_6179,N_5448,N_5064);
or U6180 (N_6180,N_5835,N_5656);
xor U6181 (N_6181,N_5768,N_5197);
nand U6182 (N_6182,N_5220,N_5237);
or U6183 (N_6183,N_5267,N_5528);
xnor U6184 (N_6184,N_5792,N_5213);
and U6185 (N_6185,N_5315,N_5740);
nand U6186 (N_6186,N_5292,N_5386);
or U6187 (N_6187,N_5299,N_5982);
nand U6188 (N_6188,N_5940,N_5741);
or U6189 (N_6189,N_5642,N_5529);
nor U6190 (N_6190,N_5666,N_5350);
or U6191 (N_6191,N_5910,N_5146);
nor U6192 (N_6192,N_5713,N_5543);
or U6193 (N_6193,N_5051,N_5484);
and U6194 (N_6194,N_5818,N_5890);
nor U6195 (N_6195,N_5466,N_5557);
and U6196 (N_6196,N_5701,N_5553);
nor U6197 (N_6197,N_5205,N_5772);
and U6198 (N_6198,N_5565,N_5276);
nand U6199 (N_6199,N_5238,N_5728);
and U6200 (N_6200,N_5021,N_5080);
and U6201 (N_6201,N_5111,N_5053);
xnor U6202 (N_6202,N_5310,N_5014);
and U6203 (N_6203,N_5707,N_5345);
xor U6204 (N_6204,N_5533,N_5290);
nand U6205 (N_6205,N_5400,N_5106);
or U6206 (N_6206,N_5588,N_5623);
nand U6207 (N_6207,N_5470,N_5416);
nor U6208 (N_6208,N_5066,N_5447);
or U6209 (N_6209,N_5510,N_5532);
nor U6210 (N_6210,N_5730,N_5720);
or U6211 (N_6211,N_5536,N_5698);
and U6212 (N_6212,N_5002,N_5592);
or U6213 (N_6213,N_5332,N_5990);
and U6214 (N_6214,N_5161,N_5551);
nor U6215 (N_6215,N_5710,N_5004);
nor U6216 (N_6216,N_5353,N_5065);
xor U6217 (N_6217,N_5145,N_5185);
nand U6218 (N_6218,N_5630,N_5571);
and U6219 (N_6219,N_5950,N_5079);
nand U6220 (N_6220,N_5566,N_5527);
nor U6221 (N_6221,N_5903,N_5487);
nand U6222 (N_6222,N_5453,N_5224);
and U6223 (N_6223,N_5232,N_5562);
and U6224 (N_6224,N_5733,N_5651);
and U6225 (N_6225,N_5653,N_5049);
xor U6226 (N_6226,N_5997,N_5776);
and U6227 (N_6227,N_5695,N_5273);
or U6228 (N_6228,N_5736,N_5164);
nand U6229 (N_6229,N_5674,N_5861);
or U6230 (N_6230,N_5591,N_5567);
and U6231 (N_6231,N_5070,N_5575);
nor U6232 (N_6232,N_5519,N_5934);
or U6233 (N_6233,N_5802,N_5918);
or U6234 (N_6234,N_5123,N_5576);
nand U6235 (N_6235,N_5775,N_5614);
and U6236 (N_6236,N_5621,N_5134);
and U6237 (N_6237,N_5899,N_5172);
nor U6238 (N_6238,N_5147,N_5622);
or U6239 (N_6239,N_5581,N_5412);
and U6240 (N_6240,N_5798,N_5929);
nor U6241 (N_6241,N_5141,N_5297);
or U6242 (N_6242,N_5324,N_5181);
or U6243 (N_6243,N_5409,N_5619);
xor U6244 (N_6244,N_5822,N_5001);
xnor U6245 (N_6245,N_5239,N_5443);
or U6246 (N_6246,N_5437,N_5479);
xnor U6247 (N_6247,N_5836,N_5774);
and U6248 (N_6248,N_5357,N_5788);
and U6249 (N_6249,N_5823,N_5590);
nand U6250 (N_6250,N_5109,N_5170);
or U6251 (N_6251,N_5909,N_5980);
and U6252 (N_6252,N_5957,N_5722);
xor U6253 (N_6253,N_5247,N_5262);
nand U6254 (N_6254,N_5702,N_5953);
and U6255 (N_6255,N_5779,N_5959);
and U6256 (N_6256,N_5761,N_5427);
and U6257 (N_6257,N_5648,N_5615);
or U6258 (N_6258,N_5785,N_5998);
nor U6259 (N_6259,N_5964,N_5883);
or U6260 (N_6260,N_5498,N_5368);
and U6261 (N_6261,N_5308,N_5196);
and U6262 (N_6262,N_5103,N_5790);
nand U6263 (N_6263,N_5005,N_5351);
and U6264 (N_6264,N_5572,N_5635);
or U6265 (N_6265,N_5280,N_5652);
nor U6266 (N_6266,N_5577,N_5979);
nor U6267 (N_6267,N_5286,N_5856);
xor U6268 (N_6268,N_5594,N_5433);
nor U6269 (N_6269,N_5865,N_5465);
or U6270 (N_6270,N_5800,N_5281);
xor U6271 (N_6271,N_5735,N_5102);
nand U6272 (N_6272,N_5474,N_5028);
xor U6273 (N_6273,N_5236,N_5935);
nor U6274 (N_6274,N_5694,N_5160);
and U6275 (N_6275,N_5071,N_5270);
xnor U6276 (N_6276,N_5655,N_5031);
and U6277 (N_6277,N_5300,N_5024);
and U6278 (N_6278,N_5367,N_5380);
or U6279 (N_6279,N_5705,N_5129);
or U6280 (N_6280,N_5739,N_5285);
and U6281 (N_6281,N_5159,N_5304);
nand U6282 (N_6282,N_5687,N_5617);
and U6283 (N_6283,N_5864,N_5283);
nand U6284 (N_6284,N_5483,N_5753);
nor U6285 (N_6285,N_5257,N_5036);
nand U6286 (N_6286,N_5711,N_5936);
and U6287 (N_6287,N_5244,N_5464);
xnor U6288 (N_6288,N_5631,N_5677);
nor U6289 (N_6289,N_5552,N_5442);
and U6290 (N_6290,N_5033,N_5764);
nor U6291 (N_6291,N_5933,N_5616);
or U6292 (N_6292,N_5187,N_5534);
nand U6293 (N_6293,N_5311,N_5363);
and U6294 (N_6294,N_5751,N_5045);
nand U6295 (N_6295,N_5022,N_5815);
or U6296 (N_6296,N_5962,N_5008);
and U6297 (N_6297,N_5747,N_5047);
and U6298 (N_6298,N_5009,N_5268);
and U6299 (N_6299,N_5058,N_5993);
or U6300 (N_6300,N_5938,N_5678);
xnor U6301 (N_6301,N_5535,N_5293);
nand U6302 (N_6302,N_5828,N_5659);
or U6303 (N_6303,N_5291,N_5636);
nor U6304 (N_6304,N_5331,N_5989);
xnor U6305 (N_6305,N_5095,N_5349);
or U6306 (N_6306,N_5343,N_5847);
xor U6307 (N_6307,N_5356,N_5354);
or U6308 (N_6308,N_5179,N_5241);
and U6309 (N_6309,N_5586,N_5688);
nand U6310 (N_6310,N_5175,N_5881);
nor U6311 (N_6311,N_5976,N_5849);
or U6312 (N_6312,N_5259,N_5190);
xnor U6313 (N_6313,N_5706,N_5419);
nand U6314 (N_6314,N_5384,N_5611);
or U6315 (N_6315,N_5803,N_5228);
nand U6316 (N_6316,N_5676,N_5225);
and U6317 (N_6317,N_5206,N_5928);
nor U6318 (N_6318,N_5016,N_5158);
xnor U6319 (N_6319,N_5855,N_5539);
and U6320 (N_6320,N_5385,N_5513);
nor U6321 (N_6321,N_5930,N_5059);
xnor U6322 (N_6322,N_5625,N_5917);
and U6323 (N_6323,N_5401,N_5770);
xor U6324 (N_6324,N_5250,N_5337);
nor U6325 (N_6325,N_5000,N_5668);
or U6326 (N_6326,N_5475,N_5926);
and U6327 (N_6327,N_5055,N_5857);
and U6328 (N_6328,N_5504,N_5420);
nor U6329 (N_6329,N_5362,N_5215);
or U6330 (N_6330,N_5421,N_5156);
and U6331 (N_6331,N_5381,N_5827);
xor U6332 (N_6332,N_5873,N_5579);
or U6333 (N_6333,N_5603,N_5389);
nand U6334 (N_6334,N_5784,N_5006);
or U6335 (N_6335,N_5554,N_5355);
nand U6336 (N_6336,N_5424,N_5272);
or U6337 (N_6337,N_5726,N_5131);
xnor U6338 (N_6338,N_5319,N_5963);
and U6339 (N_6339,N_5485,N_5832);
nor U6340 (N_6340,N_5858,N_5797);
nor U6341 (N_6341,N_5724,N_5042);
xor U6342 (N_6342,N_5482,N_5312);
xnor U6343 (N_6343,N_5578,N_5500);
and U6344 (N_6344,N_5583,N_5074);
or U6345 (N_6345,N_5023,N_5026);
nor U6346 (N_6346,N_5330,N_5640);
nor U6347 (N_6347,N_5454,N_5369);
nor U6348 (N_6348,N_5885,N_5034);
xnor U6349 (N_6349,N_5041,N_5693);
nor U6350 (N_6350,N_5921,N_5457);
xor U6351 (N_6351,N_5924,N_5452);
nand U6352 (N_6352,N_5949,N_5460);
nand U6353 (N_6353,N_5271,N_5383);
nor U6354 (N_6354,N_5947,N_5731);
xor U6355 (N_6355,N_5696,N_5675);
xor U6356 (N_6356,N_5795,N_5425);
xnor U6357 (N_6357,N_5834,N_5937);
and U6358 (N_6358,N_5073,N_5135);
nand U6359 (N_6359,N_5087,N_5378);
xor U6360 (N_6360,N_5463,N_5777);
nor U6361 (N_6361,N_5994,N_5360);
nand U6362 (N_6362,N_5948,N_5032);
nor U6363 (N_6363,N_5329,N_5977);
nor U6364 (N_6364,N_5436,N_5098);
nor U6365 (N_6365,N_5203,N_5639);
or U6366 (N_6366,N_5327,N_5681);
xor U6367 (N_6367,N_5025,N_5439);
nand U6368 (N_6368,N_5186,N_5252);
and U6369 (N_6369,N_5868,N_5415);
nor U6370 (N_6370,N_5956,N_5826);
nand U6371 (N_6371,N_5660,N_5399);
nand U6372 (N_6372,N_5769,N_5488);
and U6373 (N_6373,N_5266,N_5174);
nor U6374 (N_6374,N_5778,N_5274);
and U6375 (N_6375,N_5879,N_5854);
nor U6376 (N_6376,N_5914,N_5188);
or U6377 (N_6377,N_5809,N_5589);
xor U6378 (N_6378,N_5601,N_5850);
or U6379 (N_6379,N_5896,N_5650);
xnor U6380 (N_6380,N_5316,N_5344);
xnor U6381 (N_6381,N_5608,N_5157);
and U6382 (N_6382,N_5083,N_5679);
nand U6383 (N_6383,N_5445,N_5010);
nor U6384 (N_6384,N_5012,N_5712);
xnor U6385 (N_6385,N_5035,N_5789);
xor U6386 (N_6386,N_5495,N_5971);
or U6387 (N_6387,N_5366,N_5620);
and U6388 (N_6388,N_5996,N_5204);
and U6389 (N_6389,N_5263,N_5727);
nor U6390 (N_6390,N_5748,N_5397);
and U6391 (N_6391,N_5328,N_5234);
nand U6392 (N_6392,N_5132,N_5375);
xnor U6393 (N_6393,N_5683,N_5208);
xnor U6394 (N_6394,N_5734,N_5869);
nand U6395 (N_6395,N_5946,N_5431);
nand U6396 (N_6396,N_5472,N_5944);
xnor U6397 (N_6397,N_5125,N_5256);
nand U6398 (N_6398,N_5793,N_5606);
nand U6399 (N_6399,N_5848,N_5212);
nand U6400 (N_6400,N_5718,N_5394);
xor U6401 (N_6401,N_5255,N_5284);
xor U6402 (N_6402,N_5373,N_5760);
nor U6403 (N_6403,N_5370,N_5027);
or U6404 (N_6404,N_5322,N_5549);
nor U6405 (N_6405,N_5913,N_5871);
and U6406 (N_6406,N_5200,N_5030);
or U6407 (N_6407,N_5750,N_5089);
nand U6408 (N_6408,N_5558,N_5119);
nor U6409 (N_6409,N_5121,N_5657);
xor U6410 (N_6410,N_5040,N_5096);
nor U6411 (N_6411,N_5086,N_5686);
xor U6412 (N_6412,N_5150,N_5492);
or U6413 (N_6413,N_5169,N_5955);
nor U6414 (N_6414,N_5945,N_5092);
nand U6415 (N_6415,N_5626,N_5721);
or U6416 (N_6416,N_5902,N_5405);
or U6417 (N_6417,N_5544,N_5821);
or U6418 (N_6418,N_5811,N_5754);
nor U6419 (N_6419,N_5199,N_5396);
and U6420 (N_6420,N_5422,N_5503);
nand U6421 (N_6421,N_5202,N_5043);
nor U6422 (N_6422,N_5646,N_5569);
xor U6423 (N_6423,N_5851,N_5525);
and U6424 (N_6424,N_5227,N_5877);
or U6425 (N_6425,N_5094,N_5167);
nand U6426 (N_6426,N_5587,N_5029);
nor U6427 (N_6427,N_5163,N_5889);
nand U6428 (N_6428,N_5526,N_5501);
and U6429 (N_6429,N_5782,N_5277);
nor U6430 (N_6430,N_5288,N_5069);
nand U6431 (N_6431,N_5602,N_5853);
nand U6432 (N_6432,N_5831,N_5516);
nand U6433 (N_6433,N_5548,N_5884);
xnor U6434 (N_6434,N_5440,N_5429);
or U6435 (N_6435,N_5763,N_5670);
xnor U6436 (N_6436,N_5223,N_5673);
nor U6437 (N_6437,N_5867,N_5207);
or U6438 (N_6438,N_5233,N_5193);
and U6439 (N_6439,N_5595,N_5451);
nor U6440 (N_6440,N_5547,N_5177);
nand U6441 (N_6441,N_5090,N_5258);
xnor U6442 (N_6442,N_5506,N_5279);
nor U6443 (N_6443,N_5860,N_5600);
and U6444 (N_6444,N_5358,N_5799);
xnor U6445 (N_6445,N_5984,N_5126);
xor U6446 (N_6446,N_5294,N_5806);
xor U6447 (N_6447,N_5787,N_5117);
or U6448 (N_6448,N_5875,N_5455);
nor U6449 (N_6449,N_5107,N_5838);
nand U6450 (N_6450,N_5153,N_5414);
nand U6451 (N_6451,N_5814,N_5085);
or U6452 (N_6452,N_5374,N_5243);
nand U6453 (N_6453,N_5309,N_5719);
nand U6454 (N_6454,N_5805,N_5952);
or U6455 (N_6455,N_5478,N_5524);
nor U6456 (N_6456,N_5829,N_5235);
nor U6457 (N_6457,N_5097,N_5246);
nand U6458 (N_6458,N_5882,N_5584);
nor U6459 (N_6459,N_5171,N_5496);
xor U6460 (N_6460,N_5497,N_5282);
xnor U6461 (N_6461,N_5972,N_5061);
nor U6462 (N_6462,N_5406,N_5093);
or U6463 (N_6463,N_5302,N_5184);
or U6464 (N_6464,N_5116,N_5545);
xor U6465 (N_6465,N_5347,N_5521);
nand U6466 (N_6466,N_5911,N_5201);
nor U6467 (N_6467,N_5999,N_5876);
nor U6468 (N_6468,N_5078,N_5015);
nand U6469 (N_6469,N_5613,N_5900);
xnor U6470 (N_6470,N_5987,N_5708);
nor U6471 (N_6471,N_5796,N_5817);
or U6472 (N_6472,N_5966,N_5880);
or U6473 (N_6473,N_5515,N_5632);
nor U6474 (N_6474,N_5144,N_5629);
and U6475 (N_6475,N_5593,N_5641);
nand U6476 (N_6476,N_5081,N_5837);
and U6477 (N_6477,N_5723,N_5432);
nor U6478 (N_6478,N_5887,N_5221);
and U6479 (N_6479,N_5958,N_5895);
xor U6480 (N_6480,N_5633,N_5654);
xnor U6481 (N_6481,N_5540,N_5168);
or U6482 (N_6482,N_5560,N_5230);
xor U6483 (N_6483,N_5264,N_5714);
nor U6484 (N_6484,N_5275,N_5245);
xor U6485 (N_6485,N_5582,N_5773);
nand U6486 (N_6486,N_5387,N_5489);
xnor U6487 (N_6487,N_5878,N_5801);
nand U6488 (N_6488,N_5961,N_5446);
xnor U6489 (N_6489,N_5459,N_5195);
nor U6490 (N_6490,N_5198,N_5403);
nor U6491 (N_6491,N_5306,N_5018);
nand U6492 (N_6492,N_5390,N_5248);
nand U6493 (N_6493,N_5755,N_5139);
and U6494 (N_6494,N_5128,N_5541);
and U6495 (N_6495,N_5359,N_5898);
nand U6496 (N_6496,N_5336,N_5597);
nor U6497 (N_6497,N_5981,N_5428);
and U6498 (N_6498,N_5682,N_5499);
and U6499 (N_6499,N_5365,N_5684);
or U6500 (N_6500,N_5910,N_5627);
nor U6501 (N_6501,N_5339,N_5610);
nand U6502 (N_6502,N_5397,N_5240);
or U6503 (N_6503,N_5998,N_5941);
and U6504 (N_6504,N_5002,N_5402);
xor U6505 (N_6505,N_5566,N_5902);
and U6506 (N_6506,N_5945,N_5813);
nor U6507 (N_6507,N_5505,N_5588);
xnor U6508 (N_6508,N_5545,N_5436);
and U6509 (N_6509,N_5597,N_5881);
or U6510 (N_6510,N_5569,N_5649);
nand U6511 (N_6511,N_5413,N_5691);
nand U6512 (N_6512,N_5636,N_5762);
or U6513 (N_6513,N_5881,N_5708);
and U6514 (N_6514,N_5458,N_5432);
and U6515 (N_6515,N_5257,N_5449);
nand U6516 (N_6516,N_5610,N_5526);
nand U6517 (N_6517,N_5613,N_5656);
nand U6518 (N_6518,N_5672,N_5054);
nor U6519 (N_6519,N_5790,N_5756);
nand U6520 (N_6520,N_5126,N_5434);
xnor U6521 (N_6521,N_5882,N_5016);
nor U6522 (N_6522,N_5115,N_5066);
or U6523 (N_6523,N_5278,N_5282);
nor U6524 (N_6524,N_5359,N_5257);
nor U6525 (N_6525,N_5483,N_5115);
xor U6526 (N_6526,N_5080,N_5768);
or U6527 (N_6527,N_5327,N_5706);
nand U6528 (N_6528,N_5216,N_5910);
and U6529 (N_6529,N_5935,N_5450);
nor U6530 (N_6530,N_5426,N_5751);
nor U6531 (N_6531,N_5437,N_5768);
nor U6532 (N_6532,N_5938,N_5897);
nand U6533 (N_6533,N_5422,N_5835);
and U6534 (N_6534,N_5286,N_5161);
nand U6535 (N_6535,N_5594,N_5712);
xnor U6536 (N_6536,N_5576,N_5235);
nand U6537 (N_6537,N_5353,N_5652);
or U6538 (N_6538,N_5448,N_5467);
xor U6539 (N_6539,N_5144,N_5789);
nor U6540 (N_6540,N_5030,N_5528);
nand U6541 (N_6541,N_5960,N_5230);
and U6542 (N_6542,N_5899,N_5780);
and U6543 (N_6543,N_5038,N_5161);
and U6544 (N_6544,N_5318,N_5170);
or U6545 (N_6545,N_5929,N_5309);
nor U6546 (N_6546,N_5150,N_5811);
nor U6547 (N_6547,N_5674,N_5379);
or U6548 (N_6548,N_5450,N_5800);
nor U6549 (N_6549,N_5559,N_5526);
or U6550 (N_6550,N_5723,N_5697);
nand U6551 (N_6551,N_5619,N_5697);
or U6552 (N_6552,N_5426,N_5503);
xnor U6553 (N_6553,N_5351,N_5534);
nor U6554 (N_6554,N_5033,N_5260);
nand U6555 (N_6555,N_5053,N_5864);
nor U6556 (N_6556,N_5788,N_5538);
nor U6557 (N_6557,N_5091,N_5477);
nor U6558 (N_6558,N_5095,N_5944);
nor U6559 (N_6559,N_5505,N_5850);
and U6560 (N_6560,N_5262,N_5711);
nor U6561 (N_6561,N_5446,N_5311);
nand U6562 (N_6562,N_5895,N_5802);
xor U6563 (N_6563,N_5456,N_5873);
and U6564 (N_6564,N_5124,N_5848);
and U6565 (N_6565,N_5632,N_5262);
xor U6566 (N_6566,N_5735,N_5550);
nor U6567 (N_6567,N_5021,N_5413);
or U6568 (N_6568,N_5208,N_5018);
xor U6569 (N_6569,N_5210,N_5062);
nand U6570 (N_6570,N_5194,N_5693);
and U6571 (N_6571,N_5010,N_5116);
and U6572 (N_6572,N_5398,N_5662);
or U6573 (N_6573,N_5864,N_5535);
or U6574 (N_6574,N_5605,N_5774);
xor U6575 (N_6575,N_5106,N_5124);
xor U6576 (N_6576,N_5406,N_5349);
nor U6577 (N_6577,N_5213,N_5953);
and U6578 (N_6578,N_5087,N_5200);
nand U6579 (N_6579,N_5421,N_5010);
and U6580 (N_6580,N_5017,N_5504);
or U6581 (N_6581,N_5508,N_5975);
nand U6582 (N_6582,N_5633,N_5967);
nor U6583 (N_6583,N_5397,N_5166);
or U6584 (N_6584,N_5147,N_5320);
nand U6585 (N_6585,N_5325,N_5491);
nor U6586 (N_6586,N_5888,N_5096);
nor U6587 (N_6587,N_5475,N_5671);
xor U6588 (N_6588,N_5861,N_5791);
xor U6589 (N_6589,N_5018,N_5921);
nor U6590 (N_6590,N_5934,N_5945);
nor U6591 (N_6591,N_5625,N_5530);
xnor U6592 (N_6592,N_5784,N_5729);
and U6593 (N_6593,N_5878,N_5984);
nor U6594 (N_6594,N_5501,N_5828);
nor U6595 (N_6595,N_5308,N_5093);
and U6596 (N_6596,N_5055,N_5006);
or U6597 (N_6597,N_5478,N_5571);
nand U6598 (N_6598,N_5092,N_5302);
xor U6599 (N_6599,N_5365,N_5860);
xnor U6600 (N_6600,N_5471,N_5488);
nor U6601 (N_6601,N_5718,N_5709);
xor U6602 (N_6602,N_5418,N_5605);
nand U6603 (N_6603,N_5613,N_5317);
or U6604 (N_6604,N_5587,N_5107);
nor U6605 (N_6605,N_5985,N_5796);
xnor U6606 (N_6606,N_5354,N_5079);
nand U6607 (N_6607,N_5794,N_5141);
or U6608 (N_6608,N_5906,N_5898);
nand U6609 (N_6609,N_5460,N_5247);
and U6610 (N_6610,N_5809,N_5864);
or U6611 (N_6611,N_5371,N_5155);
and U6612 (N_6612,N_5785,N_5894);
nand U6613 (N_6613,N_5453,N_5802);
xor U6614 (N_6614,N_5956,N_5575);
and U6615 (N_6615,N_5727,N_5696);
xnor U6616 (N_6616,N_5444,N_5050);
nand U6617 (N_6617,N_5103,N_5251);
xor U6618 (N_6618,N_5997,N_5024);
xor U6619 (N_6619,N_5643,N_5763);
and U6620 (N_6620,N_5496,N_5869);
nand U6621 (N_6621,N_5188,N_5576);
or U6622 (N_6622,N_5058,N_5708);
nand U6623 (N_6623,N_5703,N_5721);
nand U6624 (N_6624,N_5742,N_5036);
and U6625 (N_6625,N_5239,N_5554);
nand U6626 (N_6626,N_5728,N_5438);
xnor U6627 (N_6627,N_5986,N_5859);
or U6628 (N_6628,N_5019,N_5263);
xnor U6629 (N_6629,N_5591,N_5437);
and U6630 (N_6630,N_5686,N_5645);
nor U6631 (N_6631,N_5598,N_5764);
nand U6632 (N_6632,N_5208,N_5039);
nand U6633 (N_6633,N_5771,N_5666);
nand U6634 (N_6634,N_5230,N_5320);
nor U6635 (N_6635,N_5439,N_5470);
nor U6636 (N_6636,N_5473,N_5501);
nor U6637 (N_6637,N_5181,N_5983);
and U6638 (N_6638,N_5081,N_5160);
and U6639 (N_6639,N_5496,N_5747);
xor U6640 (N_6640,N_5397,N_5586);
nor U6641 (N_6641,N_5944,N_5626);
xor U6642 (N_6642,N_5572,N_5612);
nand U6643 (N_6643,N_5288,N_5499);
or U6644 (N_6644,N_5955,N_5437);
or U6645 (N_6645,N_5855,N_5109);
nor U6646 (N_6646,N_5453,N_5168);
or U6647 (N_6647,N_5442,N_5993);
and U6648 (N_6648,N_5302,N_5940);
or U6649 (N_6649,N_5014,N_5632);
or U6650 (N_6650,N_5343,N_5636);
nor U6651 (N_6651,N_5298,N_5761);
xnor U6652 (N_6652,N_5404,N_5260);
and U6653 (N_6653,N_5922,N_5848);
or U6654 (N_6654,N_5445,N_5685);
or U6655 (N_6655,N_5086,N_5606);
nand U6656 (N_6656,N_5474,N_5111);
and U6657 (N_6657,N_5508,N_5407);
xnor U6658 (N_6658,N_5879,N_5908);
xor U6659 (N_6659,N_5927,N_5184);
nor U6660 (N_6660,N_5004,N_5276);
and U6661 (N_6661,N_5606,N_5895);
nand U6662 (N_6662,N_5357,N_5839);
and U6663 (N_6663,N_5194,N_5883);
nor U6664 (N_6664,N_5696,N_5560);
or U6665 (N_6665,N_5701,N_5720);
nor U6666 (N_6666,N_5370,N_5877);
and U6667 (N_6667,N_5595,N_5514);
nor U6668 (N_6668,N_5691,N_5951);
or U6669 (N_6669,N_5154,N_5887);
nor U6670 (N_6670,N_5365,N_5818);
nand U6671 (N_6671,N_5399,N_5627);
nor U6672 (N_6672,N_5525,N_5242);
nor U6673 (N_6673,N_5546,N_5089);
nor U6674 (N_6674,N_5810,N_5946);
xor U6675 (N_6675,N_5043,N_5385);
nor U6676 (N_6676,N_5060,N_5820);
nor U6677 (N_6677,N_5846,N_5945);
nor U6678 (N_6678,N_5372,N_5176);
and U6679 (N_6679,N_5006,N_5785);
and U6680 (N_6680,N_5172,N_5472);
and U6681 (N_6681,N_5178,N_5293);
and U6682 (N_6682,N_5348,N_5905);
xnor U6683 (N_6683,N_5676,N_5483);
or U6684 (N_6684,N_5405,N_5272);
or U6685 (N_6685,N_5909,N_5051);
nor U6686 (N_6686,N_5665,N_5532);
xor U6687 (N_6687,N_5824,N_5126);
xnor U6688 (N_6688,N_5522,N_5418);
xor U6689 (N_6689,N_5126,N_5263);
nand U6690 (N_6690,N_5786,N_5686);
nor U6691 (N_6691,N_5335,N_5403);
xor U6692 (N_6692,N_5746,N_5419);
nand U6693 (N_6693,N_5064,N_5194);
and U6694 (N_6694,N_5764,N_5848);
nand U6695 (N_6695,N_5867,N_5364);
or U6696 (N_6696,N_5361,N_5270);
or U6697 (N_6697,N_5857,N_5621);
xnor U6698 (N_6698,N_5285,N_5371);
xor U6699 (N_6699,N_5542,N_5757);
nor U6700 (N_6700,N_5444,N_5955);
nor U6701 (N_6701,N_5846,N_5614);
or U6702 (N_6702,N_5532,N_5575);
or U6703 (N_6703,N_5842,N_5032);
or U6704 (N_6704,N_5411,N_5243);
xor U6705 (N_6705,N_5321,N_5513);
nor U6706 (N_6706,N_5166,N_5292);
xor U6707 (N_6707,N_5212,N_5877);
and U6708 (N_6708,N_5624,N_5298);
xor U6709 (N_6709,N_5709,N_5457);
xnor U6710 (N_6710,N_5241,N_5497);
nand U6711 (N_6711,N_5573,N_5295);
or U6712 (N_6712,N_5639,N_5982);
xor U6713 (N_6713,N_5717,N_5933);
xnor U6714 (N_6714,N_5661,N_5393);
or U6715 (N_6715,N_5341,N_5472);
or U6716 (N_6716,N_5574,N_5042);
nor U6717 (N_6717,N_5679,N_5758);
xor U6718 (N_6718,N_5643,N_5748);
and U6719 (N_6719,N_5159,N_5257);
nand U6720 (N_6720,N_5043,N_5597);
xnor U6721 (N_6721,N_5700,N_5768);
and U6722 (N_6722,N_5416,N_5081);
xnor U6723 (N_6723,N_5806,N_5897);
nor U6724 (N_6724,N_5391,N_5907);
nor U6725 (N_6725,N_5063,N_5753);
nor U6726 (N_6726,N_5408,N_5316);
and U6727 (N_6727,N_5647,N_5606);
and U6728 (N_6728,N_5048,N_5546);
nand U6729 (N_6729,N_5113,N_5039);
and U6730 (N_6730,N_5030,N_5608);
xnor U6731 (N_6731,N_5339,N_5222);
xnor U6732 (N_6732,N_5176,N_5710);
and U6733 (N_6733,N_5256,N_5385);
nand U6734 (N_6734,N_5189,N_5054);
and U6735 (N_6735,N_5654,N_5200);
xnor U6736 (N_6736,N_5020,N_5654);
nor U6737 (N_6737,N_5965,N_5079);
and U6738 (N_6738,N_5904,N_5142);
nor U6739 (N_6739,N_5958,N_5581);
nor U6740 (N_6740,N_5234,N_5373);
xnor U6741 (N_6741,N_5646,N_5960);
nor U6742 (N_6742,N_5420,N_5352);
or U6743 (N_6743,N_5577,N_5194);
nand U6744 (N_6744,N_5636,N_5680);
nand U6745 (N_6745,N_5670,N_5929);
or U6746 (N_6746,N_5361,N_5326);
xnor U6747 (N_6747,N_5496,N_5338);
xnor U6748 (N_6748,N_5773,N_5133);
or U6749 (N_6749,N_5999,N_5624);
nand U6750 (N_6750,N_5803,N_5859);
xnor U6751 (N_6751,N_5789,N_5186);
nand U6752 (N_6752,N_5241,N_5720);
nand U6753 (N_6753,N_5385,N_5574);
or U6754 (N_6754,N_5278,N_5105);
or U6755 (N_6755,N_5847,N_5617);
nand U6756 (N_6756,N_5481,N_5758);
xnor U6757 (N_6757,N_5011,N_5030);
nor U6758 (N_6758,N_5896,N_5252);
or U6759 (N_6759,N_5982,N_5493);
xor U6760 (N_6760,N_5274,N_5546);
and U6761 (N_6761,N_5040,N_5226);
and U6762 (N_6762,N_5560,N_5477);
xor U6763 (N_6763,N_5383,N_5537);
and U6764 (N_6764,N_5686,N_5144);
nor U6765 (N_6765,N_5226,N_5186);
nor U6766 (N_6766,N_5611,N_5733);
or U6767 (N_6767,N_5536,N_5730);
nor U6768 (N_6768,N_5357,N_5170);
or U6769 (N_6769,N_5241,N_5366);
and U6770 (N_6770,N_5286,N_5343);
and U6771 (N_6771,N_5946,N_5392);
and U6772 (N_6772,N_5410,N_5251);
xnor U6773 (N_6773,N_5658,N_5945);
xnor U6774 (N_6774,N_5000,N_5928);
xnor U6775 (N_6775,N_5074,N_5234);
and U6776 (N_6776,N_5919,N_5624);
and U6777 (N_6777,N_5416,N_5084);
or U6778 (N_6778,N_5152,N_5974);
nor U6779 (N_6779,N_5352,N_5981);
nand U6780 (N_6780,N_5007,N_5190);
and U6781 (N_6781,N_5047,N_5201);
xor U6782 (N_6782,N_5658,N_5767);
nand U6783 (N_6783,N_5910,N_5278);
or U6784 (N_6784,N_5903,N_5079);
nand U6785 (N_6785,N_5008,N_5406);
nand U6786 (N_6786,N_5415,N_5843);
or U6787 (N_6787,N_5015,N_5369);
nand U6788 (N_6788,N_5532,N_5942);
or U6789 (N_6789,N_5891,N_5615);
xor U6790 (N_6790,N_5514,N_5601);
nand U6791 (N_6791,N_5441,N_5962);
and U6792 (N_6792,N_5010,N_5912);
or U6793 (N_6793,N_5592,N_5066);
nand U6794 (N_6794,N_5714,N_5050);
or U6795 (N_6795,N_5363,N_5686);
xor U6796 (N_6796,N_5833,N_5281);
xnor U6797 (N_6797,N_5784,N_5534);
xor U6798 (N_6798,N_5788,N_5992);
nand U6799 (N_6799,N_5669,N_5493);
or U6800 (N_6800,N_5954,N_5515);
xnor U6801 (N_6801,N_5740,N_5822);
xnor U6802 (N_6802,N_5626,N_5027);
nand U6803 (N_6803,N_5025,N_5954);
nand U6804 (N_6804,N_5254,N_5304);
nand U6805 (N_6805,N_5642,N_5549);
nor U6806 (N_6806,N_5046,N_5915);
nor U6807 (N_6807,N_5366,N_5182);
nor U6808 (N_6808,N_5266,N_5345);
and U6809 (N_6809,N_5516,N_5501);
and U6810 (N_6810,N_5887,N_5506);
or U6811 (N_6811,N_5765,N_5748);
xor U6812 (N_6812,N_5537,N_5859);
nand U6813 (N_6813,N_5902,N_5449);
nand U6814 (N_6814,N_5059,N_5601);
xor U6815 (N_6815,N_5269,N_5422);
xor U6816 (N_6816,N_5723,N_5829);
and U6817 (N_6817,N_5548,N_5376);
and U6818 (N_6818,N_5383,N_5097);
nand U6819 (N_6819,N_5721,N_5517);
xnor U6820 (N_6820,N_5297,N_5732);
nand U6821 (N_6821,N_5157,N_5127);
nand U6822 (N_6822,N_5485,N_5416);
or U6823 (N_6823,N_5588,N_5708);
nand U6824 (N_6824,N_5204,N_5469);
nor U6825 (N_6825,N_5231,N_5715);
nand U6826 (N_6826,N_5421,N_5079);
nand U6827 (N_6827,N_5057,N_5371);
nor U6828 (N_6828,N_5613,N_5879);
nand U6829 (N_6829,N_5118,N_5457);
and U6830 (N_6830,N_5030,N_5423);
nor U6831 (N_6831,N_5324,N_5313);
nor U6832 (N_6832,N_5615,N_5939);
nand U6833 (N_6833,N_5771,N_5682);
nor U6834 (N_6834,N_5050,N_5525);
nor U6835 (N_6835,N_5501,N_5913);
xor U6836 (N_6836,N_5392,N_5861);
nand U6837 (N_6837,N_5173,N_5653);
nand U6838 (N_6838,N_5958,N_5445);
and U6839 (N_6839,N_5747,N_5536);
nor U6840 (N_6840,N_5137,N_5690);
and U6841 (N_6841,N_5084,N_5288);
xor U6842 (N_6842,N_5906,N_5085);
or U6843 (N_6843,N_5607,N_5680);
nor U6844 (N_6844,N_5224,N_5087);
xor U6845 (N_6845,N_5131,N_5272);
or U6846 (N_6846,N_5102,N_5188);
nor U6847 (N_6847,N_5992,N_5317);
nor U6848 (N_6848,N_5109,N_5422);
or U6849 (N_6849,N_5458,N_5023);
nor U6850 (N_6850,N_5877,N_5307);
nor U6851 (N_6851,N_5203,N_5458);
and U6852 (N_6852,N_5799,N_5453);
and U6853 (N_6853,N_5080,N_5253);
xor U6854 (N_6854,N_5010,N_5308);
nand U6855 (N_6855,N_5791,N_5161);
nand U6856 (N_6856,N_5996,N_5884);
nor U6857 (N_6857,N_5458,N_5148);
nor U6858 (N_6858,N_5316,N_5671);
nor U6859 (N_6859,N_5616,N_5090);
nor U6860 (N_6860,N_5914,N_5169);
xor U6861 (N_6861,N_5516,N_5407);
nor U6862 (N_6862,N_5959,N_5839);
xnor U6863 (N_6863,N_5601,N_5093);
xor U6864 (N_6864,N_5987,N_5903);
and U6865 (N_6865,N_5416,N_5969);
and U6866 (N_6866,N_5405,N_5804);
xor U6867 (N_6867,N_5188,N_5696);
and U6868 (N_6868,N_5059,N_5547);
xor U6869 (N_6869,N_5999,N_5632);
nor U6870 (N_6870,N_5246,N_5499);
nor U6871 (N_6871,N_5324,N_5058);
nor U6872 (N_6872,N_5487,N_5169);
or U6873 (N_6873,N_5196,N_5931);
nand U6874 (N_6874,N_5857,N_5343);
nand U6875 (N_6875,N_5281,N_5899);
nand U6876 (N_6876,N_5365,N_5551);
and U6877 (N_6877,N_5903,N_5230);
nor U6878 (N_6878,N_5783,N_5662);
and U6879 (N_6879,N_5891,N_5621);
nand U6880 (N_6880,N_5098,N_5050);
xnor U6881 (N_6881,N_5050,N_5637);
or U6882 (N_6882,N_5328,N_5651);
nor U6883 (N_6883,N_5144,N_5721);
nand U6884 (N_6884,N_5167,N_5230);
nand U6885 (N_6885,N_5435,N_5084);
nor U6886 (N_6886,N_5099,N_5396);
or U6887 (N_6887,N_5201,N_5654);
and U6888 (N_6888,N_5201,N_5430);
nor U6889 (N_6889,N_5313,N_5391);
nor U6890 (N_6890,N_5864,N_5012);
and U6891 (N_6891,N_5007,N_5813);
nand U6892 (N_6892,N_5413,N_5158);
xnor U6893 (N_6893,N_5775,N_5518);
and U6894 (N_6894,N_5408,N_5870);
xor U6895 (N_6895,N_5999,N_5973);
xor U6896 (N_6896,N_5219,N_5164);
or U6897 (N_6897,N_5280,N_5977);
xnor U6898 (N_6898,N_5672,N_5394);
and U6899 (N_6899,N_5267,N_5325);
nor U6900 (N_6900,N_5977,N_5387);
nand U6901 (N_6901,N_5960,N_5685);
or U6902 (N_6902,N_5306,N_5780);
and U6903 (N_6903,N_5316,N_5932);
and U6904 (N_6904,N_5054,N_5711);
xnor U6905 (N_6905,N_5171,N_5982);
nand U6906 (N_6906,N_5954,N_5072);
or U6907 (N_6907,N_5218,N_5593);
xnor U6908 (N_6908,N_5609,N_5170);
nand U6909 (N_6909,N_5556,N_5190);
xnor U6910 (N_6910,N_5438,N_5037);
or U6911 (N_6911,N_5400,N_5538);
and U6912 (N_6912,N_5547,N_5988);
nor U6913 (N_6913,N_5772,N_5402);
and U6914 (N_6914,N_5088,N_5064);
xor U6915 (N_6915,N_5767,N_5280);
xor U6916 (N_6916,N_5089,N_5666);
nor U6917 (N_6917,N_5342,N_5070);
nand U6918 (N_6918,N_5536,N_5549);
or U6919 (N_6919,N_5402,N_5619);
nor U6920 (N_6920,N_5205,N_5371);
and U6921 (N_6921,N_5717,N_5370);
nand U6922 (N_6922,N_5267,N_5532);
nand U6923 (N_6923,N_5409,N_5481);
nor U6924 (N_6924,N_5794,N_5791);
nor U6925 (N_6925,N_5103,N_5801);
nand U6926 (N_6926,N_5342,N_5231);
and U6927 (N_6927,N_5727,N_5123);
and U6928 (N_6928,N_5784,N_5472);
nor U6929 (N_6929,N_5743,N_5867);
nor U6930 (N_6930,N_5173,N_5098);
nand U6931 (N_6931,N_5755,N_5600);
and U6932 (N_6932,N_5551,N_5512);
and U6933 (N_6933,N_5297,N_5444);
nand U6934 (N_6934,N_5002,N_5564);
nor U6935 (N_6935,N_5615,N_5671);
or U6936 (N_6936,N_5519,N_5544);
or U6937 (N_6937,N_5774,N_5677);
or U6938 (N_6938,N_5111,N_5177);
xor U6939 (N_6939,N_5142,N_5706);
or U6940 (N_6940,N_5609,N_5204);
xor U6941 (N_6941,N_5742,N_5343);
and U6942 (N_6942,N_5936,N_5511);
and U6943 (N_6943,N_5217,N_5419);
and U6944 (N_6944,N_5234,N_5191);
or U6945 (N_6945,N_5185,N_5113);
nand U6946 (N_6946,N_5262,N_5628);
and U6947 (N_6947,N_5050,N_5045);
xor U6948 (N_6948,N_5035,N_5366);
nor U6949 (N_6949,N_5476,N_5468);
or U6950 (N_6950,N_5648,N_5783);
nand U6951 (N_6951,N_5172,N_5368);
and U6952 (N_6952,N_5716,N_5082);
nand U6953 (N_6953,N_5700,N_5299);
or U6954 (N_6954,N_5797,N_5752);
xor U6955 (N_6955,N_5948,N_5568);
nand U6956 (N_6956,N_5370,N_5114);
and U6957 (N_6957,N_5085,N_5012);
and U6958 (N_6958,N_5066,N_5270);
nor U6959 (N_6959,N_5238,N_5576);
and U6960 (N_6960,N_5595,N_5961);
or U6961 (N_6961,N_5478,N_5063);
or U6962 (N_6962,N_5530,N_5874);
and U6963 (N_6963,N_5087,N_5019);
nor U6964 (N_6964,N_5785,N_5885);
or U6965 (N_6965,N_5085,N_5049);
nand U6966 (N_6966,N_5542,N_5445);
nor U6967 (N_6967,N_5976,N_5091);
nand U6968 (N_6968,N_5316,N_5669);
nor U6969 (N_6969,N_5008,N_5110);
nor U6970 (N_6970,N_5214,N_5614);
and U6971 (N_6971,N_5411,N_5604);
or U6972 (N_6972,N_5931,N_5403);
and U6973 (N_6973,N_5059,N_5898);
nor U6974 (N_6974,N_5470,N_5398);
xnor U6975 (N_6975,N_5737,N_5560);
xnor U6976 (N_6976,N_5781,N_5079);
and U6977 (N_6977,N_5026,N_5754);
or U6978 (N_6978,N_5089,N_5998);
nand U6979 (N_6979,N_5818,N_5726);
or U6980 (N_6980,N_5978,N_5221);
nand U6981 (N_6981,N_5866,N_5912);
nand U6982 (N_6982,N_5702,N_5038);
xor U6983 (N_6983,N_5347,N_5354);
and U6984 (N_6984,N_5553,N_5181);
and U6985 (N_6985,N_5051,N_5498);
nand U6986 (N_6986,N_5034,N_5619);
nand U6987 (N_6987,N_5777,N_5950);
or U6988 (N_6988,N_5597,N_5841);
and U6989 (N_6989,N_5417,N_5028);
or U6990 (N_6990,N_5203,N_5992);
nor U6991 (N_6991,N_5464,N_5349);
nand U6992 (N_6992,N_5908,N_5867);
xor U6993 (N_6993,N_5821,N_5685);
nor U6994 (N_6994,N_5925,N_5172);
nand U6995 (N_6995,N_5864,N_5781);
and U6996 (N_6996,N_5260,N_5789);
and U6997 (N_6997,N_5946,N_5614);
nand U6998 (N_6998,N_5102,N_5501);
nand U6999 (N_6999,N_5010,N_5536);
and U7000 (N_7000,N_6497,N_6083);
xor U7001 (N_7001,N_6583,N_6349);
or U7002 (N_7002,N_6652,N_6487);
xor U7003 (N_7003,N_6137,N_6207);
nand U7004 (N_7004,N_6218,N_6432);
nand U7005 (N_7005,N_6150,N_6530);
and U7006 (N_7006,N_6599,N_6928);
nand U7007 (N_7007,N_6976,N_6328);
or U7008 (N_7008,N_6217,N_6366);
xnor U7009 (N_7009,N_6372,N_6859);
or U7010 (N_7010,N_6513,N_6994);
nor U7011 (N_7011,N_6177,N_6194);
and U7012 (N_7012,N_6744,N_6303);
and U7013 (N_7013,N_6427,N_6109);
or U7014 (N_7014,N_6881,N_6913);
nand U7015 (N_7015,N_6105,N_6781);
nor U7016 (N_7016,N_6082,N_6557);
or U7017 (N_7017,N_6382,N_6592);
and U7018 (N_7018,N_6844,N_6935);
nand U7019 (N_7019,N_6156,N_6827);
and U7020 (N_7020,N_6421,N_6993);
and U7021 (N_7021,N_6478,N_6300);
and U7022 (N_7022,N_6727,N_6039);
nor U7023 (N_7023,N_6369,N_6880);
nor U7024 (N_7024,N_6955,N_6970);
and U7025 (N_7025,N_6721,N_6793);
and U7026 (N_7026,N_6264,N_6950);
or U7027 (N_7027,N_6835,N_6940);
xnor U7028 (N_7028,N_6834,N_6905);
xor U7029 (N_7029,N_6732,N_6331);
or U7030 (N_7030,N_6806,N_6135);
and U7031 (N_7031,N_6275,N_6226);
nand U7032 (N_7032,N_6213,N_6127);
or U7033 (N_7033,N_6733,N_6997);
nand U7034 (N_7034,N_6254,N_6613);
nand U7035 (N_7035,N_6036,N_6528);
and U7036 (N_7036,N_6554,N_6716);
nor U7037 (N_7037,N_6021,N_6821);
nand U7038 (N_7038,N_6851,N_6256);
and U7039 (N_7039,N_6942,N_6222);
nand U7040 (N_7040,N_6591,N_6374);
or U7041 (N_7041,N_6739,N_6023);
nor U7042 (N_7042,N_6816,N_6323);
nor U7043 (N_7043,N_6798,N_6964);
nor U7044 (N_7044,N_6279,N_6734);
or U7045 (N_7045,N_6261,N_6885);
xor U7046 (N_7046,N_6989,N_6471);
xnor U7047 (N_7047,N_6790,N_6130);
and U7048 (N_7048,N_6075,N_6878);
xor U7049 (N_7049,N_6166,N_6304);
and U7050 (N_7050,N_6623,N_6079);
or U7051 (N_7051,N_6125,N_6159);
or U7052 (N_7052,N_6854,N_6832);
xor U7053 (N_7053,N_6355,N_6702);
nor U7054 (N_7054,N_6945,N_6937);
nor U7055 (N_7055,N_6123,N_6726);
xor U7056 (N_7056,N_6643,N_6665);
or U7057 (N_7057,N_6017,N_6977);
xnor U7058 (N_7058,N_6552,N_6291);
or U7059 (N_7059,N_6695,N_6181);
and U7060 (N_7060,N_6296,N_6171);
or U7061 (N_7061,N_6801,N_6051);
nand U7062 (N_7062,N_6338,N_6126);
xor U7063 (N_7063,N_6433,N_6388);
nand U7064 (N_7064,N_6979,N_6451);
nand U7065 (N_7065,N_6968,N_6020);
or U7066 (N_7066,N_6621,N_6059);
or U7067 (N_7067,N_6795,N_6563);
xnor U7068 (N_7068,N_6522,N_6353);
or U7069 (N_7069,N_6581,N_6167);
and U7070 (N_7070,N_6229,N_6667);
and U7071 (N_7071,N_6956,N_6546);
nor U7072 (N_7072,N_6352,N_6629);
nor U7073 (N_7073,N_6312,N_6189);
and U7074 (N_7074,N_6660,N_6515);
xnor U7075 (N_7075,N_6722,N_6814);
nand U7076 (N_7076,N_6289,N_6507);
and U7077 (N_7077,N_6327,N_6991);
nor U7078 (N_7078,N_6933,N_6607);
nor U7079 (N_7079,N_6674,N_6639);
nand U7080 (N_7080,N_6415,N_6406);
nand U7081 (N_7081,N_6266,N_6815);
nor U7082 (N_7082,N_6035,N_6092);
nor U7083 (N_7083,N_6953,N_6762);
xor U7084 (N_7084,N_6957,N_6679);
xnor U7085 (N_7085,N_6142,N_6321);
xor U7086 (N_7086,N_6297,N_6740);
and U7087 (N_7087,N_6718,N_6749);
or U7088 (N_7088,N_6817,N_6715);
xor U7089 (N_7089,N_6484,N_6646);
xor U7090 (N_7090,N_6430,N_6984);
nor U7091 (N_7091,N_6265,N_6408);
nand U7092 (N_7092,N_6418,N_6414);
xnor U7093 (N_7093,N_6416,N_6775);
and U7094 (N_7094,N_6398,N_6999);
or U7095 (N_7095,N_6753,N_6360);
nor U7096 (N_7096,N_6225,N_6305);
nand U7097 (N_7097,N_6966,N_6567);
or U7098 (N_7098,N_6308,N_6258);
nand U7099 (N_7099,N_6384,N_6751);
xnor U7100 (N_7100,N_6129,N_6146);
nand U7101 (N_7101,N_6198,N_6253);
nor U7102 (N_7102,N_6524,N_6120);
and U7103 (N_7103,N_6044,N_6435);
nand U7104 (N_7104,N_6713,N_6981);
and U7105 (N_7105,N_6511,N_6315);
or U7106 (N_7106,N_6234,N_6015);
xnor U7107 (N_7107,N_6914,N_6439);
or U7108 (N_7108,N_6124,N_6049);
nand U7109 (N_7109,N_6499,N_6002);
xor U7110 (N_7110,N_6479,N_6918);
xnor U7111 (N_7111,N_6974,N_6717);
and U7112 (N_7112,N_6568,N_6813);
nand U7113 (N_7113,N_6385,N_6888);
nand U7114 (N_7114,N_6894,N_6469);
nor U7115 (N_7115,N_6411,N_6809);
xnor U7116 (N_7116,N_6985,N_6954);
nor U7117 (N_7117,N_6285,N_6086);
or U7118 (N_7118,N_6370,N_6473);
xor U7119 (N_7119,N_6804,N_6377);
nor U7120 (N_7120,N_6910,N_6431);
and U7121 (N_7121,N_6151,N_6058);
nor U7122 (N_7122,N_6040,N_6470);
nand U7123 (N_7123,N_6493,N_6367);
or U7124 (N_7124,N_6555,N_6019);
xor U7125 (N_7125,N_6833,N_6657);
nor U7126 (N_7126,N_6316,N_6066);
or U7127 (N_7127,N_6277,N_6869);
and U7128 (N_7128,N_6201,N_6050);
nand U7129 (N_7129,N_6383,N_6235);
or U7130 (N_7130,N_6375,N_6533);
nand U7131 (N_7131,N_6429,N_6392);
nor U7132 (N_7132,N_6365,N_6683);
xnor U7133 (N_7133,N_6053,N_6962);
nor U7134 (N_7134,N_6593,N_6428);
nor U7135 (N_7135,N_6608,N_6586);
xor U7136 (N_7136,N_6995,N_6455);
or U7137 (N_7137,N_6875,N_6932);
nor U7138 (N_7138,N_6446,N_6299);
nand U7139 (N_7139,N_6708,N_6873);
and U7140 (N_7140,N_6409,N_6938);
or U7141 (N_7141,N_6559,N_6788);
or U7142 (N_7142,N_6787,N_6260);
nand U7143 (N_7143,N_6005,N_6653);
xor U7144 (N_7144,N_6322,N_6892);
nand U7145 (N_7145,N_6617,N_6893);
nor U7146 (N_7146,N_6257,N_6046);
or U7147 (N_7147,N_6014,N_6401);
or U7148 (N_7148,N_6495,N_6846);
nor U7149 (N_7149,N_6441,N_6792);
xnor U7150 (N_7150,N_6776,N_6246);
nand U7151 (N_7151,N_6687,N_6663);
or U7152 (N_7152,N_6149,N_6025);
nand U7153 (N_7153,N_6670,N_6565);
nor U7154 (N_7154,N_6139,N_6063);
nor U7155 (N_7155,N_6114,N_6115);
nor U7156 (N_7156,N_6154,N_6466);
nor U7157 (N_7157,N_6209,N_6627);
nor U7158 (N_7158,N_6424,N_6822);
or U7159 (N_7159,N_6288,N_6272);
nor U7160 (N_7160,N_6969,N_6172);
xor U7161 (N_7161,N_6248,N_6532);
and U7162 (N_7162,N_6378,N_6140);
and U7163 (N_7163,N_6205,N_6029);
or U7164 (N_7164,N_6443,N_6868);
nand U7165 (N_7165,N_6022,N_6024);
nor U7166 (N_7166,N_6199,N_6699);
nand U7167 (N_7167,N_6498,N_6819);
xnor U7168 (N_7168,N_6319,N_6230);
nand U7169 (N_7169,N_6628,N_6697);
nand U7170 (N_7170,N_6179,N_6637);
nand U7171 (N_7171,N_6489,N_6459);
and U7172 (N_7172,N_6197,N_6929);
nor U7173 (N_7173,N_6931,N_6853);
or U7174 (N_7174,N_6756,N_6930);
nand U7175 (N_7175,N_6452,N_6284);
nor U7176 (N_7176,N_6512,N_6476);
xor U7177 (N_7177,N_6803,N_6810);
or U7178 (N_7178,N_6444,N_6601);
nand U7179 (N_7179,N_6061,N_6185);
or U7180 (N_7180,N_6967,N_6691);
or U7181 (N_7181,N_6768,N_6326);
nand U7182 (N_7182,N_6636,N_6820);
or U7183 (N_7183,N_6437,N_6840);
or U7184 (N_7184,N_6763,N_6067);
nor U7185 (N_7185,N_6055,N_6153);
or U7186 (N_7186,N_6774,N_6596);
nor U7187 (N_7187,N_6758,N_6188);
and U7188 (N_7188,N_6348,N_6357);
nor U7189 (N_7189,N_6541,N_6004);
nand U7190 (N_7190,N_6943,N_6417);
xnor U7191 (N_7191,N_6735,N_6915);
xor U7192 (N_7192,N_6706,N_6152);
and U7193 (N_7193,N_6068,N_6693);
nand U7194 (N_7194,N_6602,N_6582);
nor U7195 (N_7195,N_6001,N_6496);
or U7196 (N_7196,N_6381,N_6520);
xor U7197 (N_7197,N_6677,N_6710);
xor U7198 (N_7198,N_6797,N_6219);
nand U7199 (N_7199,N_6924,N_6886);
xnor U7200 (N_7200,N_6902,N_6688);
or U7201 (N_7201,N_6630,N_6842);
and U7202 (N_7202,N_6661,N_6448);
and U7203 (N_7203,N_6397,N_6460);
nor U7204 (N_7204,N_6342,N_6642);
nor U7205 (N_7205,N_6508,N_6765);
nor U7206 (N_7206,N_6645,N_6274);
and U7207 (N_7207,N_6684,N_6088);
nand U7208 (N_7208,N_6477,N_6826);
nand U7209 (N_7209,N_6823,N_6074);
nor U7210 (N_7210,N_6936,N_6671);
nand U7211 (N_7211,N_6566,N_6920);
xnor U7212 (N_7212,N_6690,N_6454);
nor U7213 (N_7213,N_6203,N_6101);
and U7214 (N_7214,N_6594,N_6633);
and U7215 (N_7215,N_6211,N_6604);
or U7216 (N_7216,N_6673,N_6379);
and U7217 (N_7217,N_6099,N_6685);
nand U7218 (N_7218,N_6456,N_6168);
xor U7219 (N_7219,N_6165,N_6413);
nand U7220 (N_7220,N_6490,N_6482);
and U7221 (N_7221,N_6675,N_6286);
nor U7222 (N_7222,N_6784,N_6491);
xor U7223 (N_7223,N_6380,N_6746);
and U7224 (N_7224,N_6231,N_6314);
and U7225 (N_7225,N_6925,N_6526);
xor U7226 (N_7226,N_6098,N_6085);
nand U7227 (N_7227,N_6195,N_6647);
nand U7228 (N_7228,N_6998,N_6527);
nand U7229 (N_7229,N_6811,N_6239);
or U7230 (N_7230,N_6077,N_6073);
or U7231 (N_7231,N_6975,N_6010);
nand U7232 (N_7232,N_6944,N_6777);
nor U7233 (N_7233,N_6148,N_6659);
xor U7234 (N_7234,N_6668,N_6570);
and U7235 (N_7235,N_6605,N_6959);
or U7236 (N_7236,N_6799,N_6503);
nand U7237 (N_7237,N_6650,N_6295);
nand U7238 (N_7238,N_6536,N_6350);
nor U7239 (N_7239,N_6576,N_6064);
xnor U7240 (N_7240,N_6463,N_6506);
and U7241 (N_7241,N_6373,N_6093);
and U7242 (N_7242,N_6542,N_6325);
xnor U7243 (N_7243,N_6584,N_6849);
and U7244 (N_7244,N_6237,N_6707);
xnor U7245 (N_7245,N_6648,N_6644);
nand U7246 (N_7246,N_6324,N_6764);
or U7247 (N_7247,N_6738,N_6026);
nor U7248 (N_7248,N_6119,N_6818);
and U7249 (N_7249,N_6622,N_6157);
or U7250 (N_7250,N_6794,N_6863);
nor U7251 (N_7251,N_6802,N_6233);
nand U7252 (N_7252,N_6951,N_6193);
nor U7253 (N_7253,N_6281,N_6097);
and U7254 (N_7254,N_6133,N_6719);
nand U7255 (N_7255,N_6362,N_6184);
xor U7256 (N_7256,N_6472,N_6867);
xor U7257 (N_7257,N_6094,N_6917);
nor U7258 (N_7258,N_6070,N_6339);
xnor U7259 (N_7259,N_6850,N_6509);
or U7260 (N_7260,N_6882,N_6212);
or U7261 (N_7261,N_6095,N_6462);
nand U7262 (N_7262,N_6041,N_6445);
xnor U7263 (N_7263,N_6042,N_6712);
xnor U7264 (N_7264,N_6830,N_6278);
xnor U7265 (N_7265,N_6603,N_6824);
nand U7266 (N_7266,N_6271,N_6006);
nand U7267 (N_7267,N_6879,N_6761);
or U7268 (N_7268,N_6887,N_6032);
nor U7269 (N_7269,N_6828,N_6676);
and U7270 (N_7270,N_6890,N_6364);
and U7271 (N_7271,N_6048,N_6737);
xor U7272 (N_7272,N_6155,N_6502);
and U7273 (N_7273,N_6494,N_6728);
nor U7274 (N_7274,N_6987,N_6909);
and U7275 (N_7275,N_6293,N_6071);
and U7276 (N_7276,N_6045,N_6216);
nand U7277 (N_7277,N_6919,N_6662);
xor U7278 (N_7278,N_6344,N_6807);
xor U7279 (N_7279,N_6585,N_6600);
nand U7280 (N_7280,N_6741,N_6711);
and U7281 (N_7281,N_6529,N_6837);
nand U7282 (N_7282,N_6615,N_6864);
xnor U7283 (N_7283,N_6680,N_6587);
and U7284 (N_7284,N_6180,N_6825);
nand U7285 (N_7285,N_6488,N_6173);
and U7286 (N_7286,N_6589,N_6333);
or U7287 (N_7287,N_6754,N_6730);
nor U7288 (N_7288,N_6128,N_6301);
xor U7289 (N_7289,N_6877,N_6030);
xnor U7290 (N_7290,N_6899,N_6147);
nor U7291 (N_7291,N_6539,N_6400);
or U7292 (N_7292,N_6263,N_6320);
nor U7293 (N_7293,N_6485,N_6332);
xnor U7294 (N_7294,N_6343,N_6031);
nor U7295 (N_7295,N_6317,N_6723);
and U7296 (N_7296,N_6672,N_6250);
or U7297 (N_7297,N_6860,N_6946);
or U7298 (N_7298,N_6907,N_6089);
nor U7299 (N_7299,N_6525,N_6268);
or U7300 (N_7300,N_6183,N_6390);
xnor U7301 (N_7301,N_6786,N_6874);
xor U7302 (N_7302,N_6556,N_6434);
nor U7303 (N_7303,N_6204,N_6108);
nor U7304 (N_7304,N_6852,N_6341);
xor U7305 (N_7305,N_6076,N_6387);
nand U7306 (N_7306,N_6161,N_6610);
nand U7307 (N_7307,N_6916,N_6939);
nand U7308 (N_7308,N_6992,N_6961);
xor U7309 (N_7309,N_6337,N_6090);
nor U7310 (N_7310,N_6876,N_6122);
nor U7311 (N_7311,N_6871,N_6080);
or U7312 (N_7312,N_6666,N_6612);
xnor U7313 (N_7313,N_6163,N_6412);
nor U7314 (N_7314,N_6043,N_6549);
nor U7315 (N_7315,N_6221,N_6550);
nand U7316 (N_7316,N_6182,N_6904);
or U7317 (N_7317,N_6110,N_6251);
xnor U7318 (N_7318,N_6290,N_6923);
xor U7319 (N_7319,N_6958,N_6096);
and U7320 (N_7320,N_6561,N_6769);
xor U7321 (N_7321,N_6574,N_6689);
nor U7322 (N_7322,N_6145,N_6486);
nand U7323 (N_7323,N_6773,N_6638);
nor U7324 (N_7324,N_6767,N_6404);
or U7325 (N_7325,N_6861,N_6705);
nand U7326 (N_7326,N_6800,N_6116);
nand U7327 (N_7327,N_6696,N_6843);
nand U7328 (N_7328,N_6354,N_6371);
nor U7329 (N_7329,N_6069,N_6169);
and U7330 (N_7330,N_6065,N_6078);
or U7331 (N_7331,N_6008,N_6641);
and U7332 (N_7332,N_6298,N_6011);
nor U7333 (N_7333,N_6597,N_6839);
and U7334 (N_7334,N_6287,N_6252);
nor U7335 (N_7335,N_6208,N_6598);
and U7336 (N_7336,N_6438,N_6698);
or U7337 (N_7337,N_6606,N_6259);
and U7338 (N_7338,N_6947,N_6748);
nor U7339 (N_7339,N_6395,N_6577);
nor U7340 (N_7340,N_6480,N_6033);
xor U7341 (N_7341,N_6483,N_6236);
or U7342 (N_7342,N_6616,N_6573);
xor U7343 (N_7343,N_6847,N_6921);
nor U7344 (N_7344,N_6655,N_6866);
nor U7345 (N_7345,N_6664,N_6791);
xor U7346 (N_7346,N_6162,N_6028);
nor U7347 (N_7347,N_6669,N_6037);
nand U7348 (N_7348,N_6003,N_6276);
and U7349 (N_7349,N_6027,N_6112);
xnor U7350 (N_7350,N_6883,N_6841);
xnor U7351 (N_7351,N_6911,N_6649);
nor U7352 (N_7352,N_6273,N_6562);
nor U7353 (N_7353,N_6747,N_6104);
and U7354 (N_7354,N_6228,N_6922);
and U7355 (N_7355,N_6965,N_6131);
and U7356 (N_7356,N_6619,N_6346);
or U7357 (N_7357,N_6973,N_6521);
nor U7358 (N_7358,N_6531,N_6087);
and U7359 (N_7359,N_6458,N_6564);
or U7360 (N_7360,N_6926,N_6238);
and U7361 (N_7361,N_6419,N_6117);
and U7362 (N_7362,N_6174,N_6245);
xnor U7363 (N_7363,N_6255,N_6505);
nand U7364 (N_7364,N_6215,N_6537);
nand U7365 (N_7365,N_6575,N_6391);
xnor U7366 (N_7366,N_6518,N_6618);
nand U7367 (N_7367,N_6270,N_6190);
nor U7368 (N_7368,N_6113,N_6510);
nand U7369 (N_7369,N_6389,N_6103);
nand U7370 (N_7370,N_6363,N_6934);
xnor U7371 (N_7371,N_6187,N_6329);
or U7372 (N_7372,N_6249,N_6848);
xnor U7373 (N_7373,N_6242,N_6558);
or U7374 (N_7374,N_6340,N_6464);
nand U7375 (N_7375,N_6423,N_6057);
or U7376 (N_7376,N_6681,N_6143);
nand U7377 (N_7377,N_6160,N_6232);
or U7378 (N_7378,N_6560,N_6782);
nor U7379 (N_7379,N_6898,N_6745);
or U7380 (N_7380,N_6426,N_6831);
nor U7381 (N_7381,N_6729,N_6812);
and U7382 (N_7382,N_6492,N_6980);
xnor U7383 (N_7383,N_6703,N_6971);
and U7384 (N_7384,N_6227,N_6358);
or U7385 (N_7385,N_6158,N_6138);
xnor U7386 (N_7386,N_6106,N_6829);
and U7387 (N_7387,N_6241,N_6170);
nor U7388 (N_7388,N_6862,N_6345);
xnor U7389 (N_7389,N_6750,N_6175);
xnor U7390 (N_7390,N_6779,N_6481);
and U7391 (N_7391,N_6052,N_6658);
or U7392 (N_7392,N_6262,N_6440);
and U7393 (N_7393,N_6760,N_6223);
xnor U7394 (N_7394,N_6780,N_6313);
nor U7395 (N_7395,N_6982,N_6724);
xor U7396 (N_7396,N_6118,N_6368);
nand U7397 (N_7397,N_6889,N_6772);
and U7398 (N_7398,N_6538,N_6590);
xnor U7399 (N_7399,N_6062,N_6012);
xor U7400 (N_7400,N_6578,N_6500);
nor U7401 (N_7401,N_6191,N_6694);
nor U7402 (N_7402,N_6900,N_6949);
and U7403 (N_7403,N_6631,N_6176);
nor U7404 (N_7404,N_6196,N_6038);
xnor U7405 (N_7405,N_6422,N_6897);
and U7406 (N_7406,N_6517,N_6865);
nor U7407 (N_7407,N_6941,N_6282);
nor U7408 (N_7408,N_6519,N_6635);
or U7409 (N_7409,N_6091,N_6901);
nor U7410 (N_7410,N_6656,N_6686);
nand U7411 (N_7411,N_6356,N_6056);
xnor U7412 (N_7412,N_6912,N_6283);
xor U7413 (N_7413,N_6571,N_6535);
and U7414 (N_7414,N_6394,N_6475);
or U7415 (N_7415,N_6220,N_6700);
and U7416 (N_7416,N_6678,N_6551);
nand U7417 (N_7417,N_6704,N_6990);
nand U7418 (N_7418,N_6336,N_6202);
nand U7419 (N_7419,N_6224,N_6742);
nor U7420 (N_7420,N_6402,N_6770);
xnor U7421 (N_7421,N_6632,N_6192);
and U7422 (N_7422,N_6620,N_6963);
xnor U7423 (N_7423,N_6359,N_6714);
nor U7424 (N_7424,N_6692,N_6474);
xor U7425 (N_7425,N_6857,N_6436);
and U7426 (N_7426,N_6311,N_6102);
xor U7427 (N_7427,N_6891,N_6872);
xor U7428 (N_7428,N_6569,N_6468);
and U7429 (N_7429,N_6789,N_6624);
xnor U7430 (N_7430,N_6141,N_6200);
nor U7431 (N_7431,N_6420,N_6701);
xor U7432 (N_7432,N_6111,N_6009);
nand U7433 (N_7433,N_6836,N_6461);
nand U7434 (N_7434,N_6785,N_6614);
and U7435 (N_7435,N_6855,N_6292);
and U7436 (N_7436,N_6450,N_6534);
xor U7437 (N_7437,N_6796,N_6178);
nand U7438 (N_7438,N_6410,N_6425);
nor U7439 (N_7439,N_6310,N_6580);
nor U7440 (N_7440,N_6514,N_6838);
nand U7441 (N_7441,N_6743,N_6972);
nand U7442 (N_7442,N_6405,N_6588);
nor U7443 (N_7443,N_6952,N_6752);
and U7444 (N_7444,N_6121,N_6453);
xor U7445 (N_7445,N_6243,N_6280);
or U7446 (N_7446,N_6625,N_6047);
or U7447 (N_7447,N_6054,N_6805);
nand U7448 (N_7448,N_6736,N_6540);
nor U7449 (N_7449,N_6081,N_6547);
nor U7450 (N_7450,N_6783,N_6132);
and U7451 (N_7451,N_6294,N_6579);
and U7452 (N_7452,N_6766,N_6870);
and U7453 (N_7453,N_6609,N_6307);
or U7454 (N_7454,N_6516,N_6978);
nand U7455 (N_7455,N_6757,N_6545);
or U7456 (N_7456,N_6543,N_6611);
or U7457 (N_7457,N_6396,N_6000);
xnor U7458 (N_7458,N_6267,N_6386);
xnor U7459 (N_7459,N_6164,N_6072);
and U7460 (N_7460,N_6501,N_6210);
and U7461 (N_7461,N_6755,N_6351);
and U7462 (N_7462,N_6731,N_6206);
nand U7463 (N_7463,N_6808,N_6908);
xnor U7464 (N_7464,N_6084,N_6640);
or U7465 (N_7465,N_6960,N_6634);
xor U7466 (N_7466,N_6906,N_6759);
or U7467 (N_7467,N_6654,N_6553);
xnor U7468 (N_7468,N_6720,N_6407);
and U7469 (N_7469,N_6983,N_6884);
or U7470 (N_7470,N_6347,N_6626);
or U7471 (N_7471,N_6709,N_6442);
nand U7472 (N_7472,N_6376,N_6100);
and U7473 (N_7473,N_6136,N_6247);
or U7474 (N_7474,N_6034,N_6778);
nor U7475 (N_7475,N_6007,N_6523);
nor U7476 (N_7476,N_6771,N_6996);
nand U7477 (N_7477,N_6651,N_6186);
nand U7478 (N_7478,N_6447,N_6465);
nor U7479 (N_7479,N_6988,N_6335);
nor U7480 (N_7480,N_6449,N_6856);
xnor U7481 (N_7481,N_6504,N_6013);
or U7482 (N_7482,N_6403,N_6309);
and U7483 (N_7483,N_6845,N_6240);
xor U7484 (N_7484,N_6318,N_6927);
nor U7485 (N_7485,N_6858,N_6393);
nand U7486 (N_7486,N_6725,N_6896);
xnor U7487 (N_7487,N_6134,N_6269);
xnor U7488 (N_7488,N_6214,N_6244);
nand U7489 (N_7489,N_6948,N_6334);
xnor U7490 (N_7490,N_6361,N_6016);
nand U7491 (N_7491,N_6548,N_6595);
nand U7492 (N_7492,N_6986,N_6144);
or U7493 (N_7493,N_6895,N_6457);
xnor U7494 (N_7494,N_6060,N_6107);
and U7495 (N_7495,N_6467,N_6682);
xnor U7496 (N_7496,N_6544,N_6903);
or U7497 (N_7497,N_6018,N_6306);
nor U7498 (N_7498,N_6302,N_6399);
or U7499 (N_7499,N_6572,N_6330);
and U7500 (N_7500,N_6491,N_6256);
nor U7501 (N_7501,N_6014,N_6480);
and U7502 (N_7502,N_6657,N_6202);
or U7503 (N_7503,N_6148,N_6930);
nand U7504 (N_7504,N_6249,N_6861);
nor U7505 (N_7505,N_6156,N_6248);
or U7506 (N_7506,N_6252,N_6146);
and U7507 (N_7507,N_6336,N_6206);
and U7508 (N_7508,N_6240,N_6739);
nand U7509 (N_7509,N_6786,N_6955);
xor U7510 (N_7510,N_6667,N_6784);
or U7511 (N_7511,N_6669,N_6359);
and U7512 (N_7512,N_6244,N_6084);
and U7513 (N_7513,N_6122,N_6818);
and U7514 (N_7514,N_6247,N_6691);
nand U7515 (N_7515,N_6378,N_6032);
xnor U7516 (N_7516,N_6193,N_6269);
or U7517 (N_7517,N_6269,N_6381);
nand U7518 (N_7518,N_6347,N_6193);
nand U7519 (N_7519,N_6886,N_6670);
and U7520 (N_7520,N_6231,N_6056);
nand U7521 (N_7521,N_6745,N_6451);
nor U7522 (N_7522,N_6953,N_6576);
or U7523 (N_7523,N_6121,N_6163);
or U7524 (N_7524,N_6779,N_6207);
xnor U7525 (N_7525,N_6990,N_6986);
xnor U7526 (N_7526,N_6651,N_6523);
or U7527 (N_7527,N_6032,N_6475);
xor U7528 (N_7528,N_6680,N_6164);
nor U7529 (N_7529,N_6350,N_6299);
nand U7530 (N_7530,N_6943,N_6567);
or U7531 (N_7531,N_6856,N_6171);
or U7532 (N_7532,N_6736,N_6306);
xnor U7533 (N_7533,N_6713,N_6309);
nor U7534 (N_7534,N_6364,N_6333);
nand U7535 (N_7535,N_6342,N_6271);
or U7536 (N_7536,N_6045,N_6931);
nor U7537 (N_7537,N_6576,N_6057);
nor U7538 (N_7538,N_6731,N_6934);
nor U7539 (N_7539,N_6761,N_6513);
or U7540 (N_7540,N_6428,N_6185);
or U7541 (N_7541,N_6919,N_6513);
and U7542 (N_7542,N_6783,N_6761);
xnor U7543 (N_7543,N_6681,N_6947);
xor U7544 (N_7544,N_6783,N_6338);
nand U7545 (N_7545,N_6290,N_6857);
and U7546 (N_7546,N_6406,N_6655);
nor U7547 (N_7547,N_6726,N_6423);
nor U7548 (N_7548,N_6225,N_6275);
and U7549 (N_7549,N_6220,N_6056);
and U7550 (N_7550,N_6239,N_6056);
nor U7551 (N_7551,N_6907,N_6767);
or U7552 (N_7552,N_6822,N_6537);
and U7553 (N_7553,N_6374,N_6141);
xnor U7554 (N_7554,N_6092,N_6771);
nor U7555 (N_7555,N_6556,N_6892);
nor U7556 (N_7556,N_6824,N_6978);
nand U7557 (N_7557,N_6301,N_6631);
nand U7558 (N_7558,N_6256,N_6325);
xnor U7559 (N_7559,N_6609,N_6874);
and U7560 (N_7560,N_6242,N_6289);
or U7561 (N_7561,N_6186,N_6931);
nor U7562 (N_7562,N_6034,N_6984);
nor U7563 (N_7563,N_6603,N_6367);
and U7564 (N_7564,N_6629,N_6456);
nand U7565 (N_7565,N_6816,N_6695);
nor U7566 (N_7566,N_6900,N_6526);
nor U7567 (N_7567,N_6044,N_6473);
or U7568 (N_7568,N_6220,N_6879);
and U7569 (N_7569,N_6867,N_6699);
xor U7570 (N_7570,N_6996,N_6103);
nor U7571 (N_7571,N_6934,N_6730);
nor U7572 (N_7572,N_6390,N_6156);
or U7573 (N_7573,N_6769,N_6284);
and U7574 (N_7574,N_6396,N_6168);
or U7575 (N_7575,N_6067,N_6131);
nand U7576 (N_7576,N_6305,N_6781);
xnor U7577 (N_7577,N_6047,N_6137);
or U7578 (N_7578,N_6252,N_6434);
nand U7579 (N_7579,N_6366,N_6896);
or U7580 (N_7580,N_6233,N_6133);
and U7581 (N_7581,N_6026,N_6120);
xor U7582 (N_7582,N_6965,N_6247);
xnor U7583 (N_7583,N_6573,N_6750);
nand U7584 (N_7584,N_6101,N_6955);
nand U7585 (N_7585,N_6530,N_6749);
or U7586 (N_7586,N_6051,N_6797);
nand U7587 (N_7587,N_6570,N_6008);
xnor U7588 (N_7588,N_6477,N_6756);
or U7589 (N_7589,N_6782,N_6354);
or U7590 (N_7590,N_6696,N_6950);
xnor U7591 (N_7591,N_6064,N_6633);
or U7592 (N_7592,N_6236,N_6184);
and U7593 (N_7593,N_6432,N_6072);
xnor U7594 (N_7594,N_6255,N_6784);
xnor U7595 (N_7595,N_6264,N_6959);
and U7596 (N_7596,N_6355,N_6704);
xor U7597 (N_7597,N_6588,N_6304);
nand U7598 (N_7598,N_6871,N_6096);
nand U7599 (N_7599,N_6006,N_6654);
xnor U7600 (N_7600,N_6455,N_6028);
nand U7601 (N_7601,N_6610,N_6730);
xor U7602 (N_7602,N_6436,N_6256);
and U7603 (N_7603,N_6069,N_6636);
nor U7604 (N_7604,N_6902,N_6148);
nand U7605 (N_7605,N_6498,N_6038);
nor U7606 (N_7606,N_6777,N_6527);
and U7607 (N_7607,N_6029,N_6899);
and U7608 (N_7608,N_6410,N_6575);
nand U7609 (N_7609,N_6453,N_6906);
or U7610 (N_7610,N_6145,N_6011);
nor U7611 (N_7611,N_6749,N_6068);
and U7612 (N_7612,N_6346,N_6990);
and U7613 (N_7613,N_6317,N_6051);
nand U7614 (N_7614,N_6006,N_6430);
and U7615 (N_7615,N_6888,N_6407);
xor U7616 (N_7616,N_6074,N_6819);
nor U7617 (N_7617,N_6143,N_6776);
xnor U7618 (N_7618,N_6601,N_6592);
xor U7619 (N_7619,N_6633,N_6328);
nor U7620 (N_7620,N_6384,N_6790);
or U7621 (N_7621,N_6313,N_6214);
nand U7622 (N_7622,N_6780,N_6919);
xnor U7623 (N_7623,N_6278,N_6712);
or U7624 (N_7624,N_6587,N_6670);
nor U7625 (N_7625,N_6570,N_6506);
nand U7626 (N_7626,N_6971,N_6854);
nand U7627 (N_7627,N_6159,N_6025);
or U7628 (N_7628,N_6390,N_6658);
nor U7629 (N_7629,N_6500,N_6447);
nor U7630 (N_7630,N_6516,N_6820);
or U7631 (N_7631,N_6359,N_6406);
nand U7632 (N_7632,N_6022,N_6431);
and U7633 (N_7633,N_6786,N_6989);
or U7634 (N_7634,N_6832,N_6789);
or U7635 (N_7635,N_6674,N_6581);
or U7636 (N_7636,N_6552,N_6692);
or U7637 (N_7637,N_6105,N_6248);
nand U7638 (N_7638,N_6226,N_6732);
nor U7639 (N_7639,N_6811,N_6753);
xnor U7640 (N_7640,N_6971,N_6834);
or U7641 (N_7641,N_6445,N_6203);
and U7642 (N_7642,N_6229,N_6354);
or U7643 (N_7643,N_6624,N_6198);
and U7644 (N_7644,N_6489,N_6732);
nor U7645 (N_7645,N_6061,N_6919);
or U7646 (N_7646,N_6645,N_6535);
and U7647 (N_7647,N_6242,N_6992);
and U7648 (N_7648,N_6003,N_6087);
xnor U7649 (N_7649,N_6605,N_6743);
xnor U7650 (N_7650,N_6067,N_6176);
nand U7651 (N_7651,N_6977,N_6479);
nor U7652 (N_7652,N_6748,N_6294);
nand U7653 (N_7653,N_6741,N_6999);
nor U7654 (N_7654,N_6364,N_6372);
nor U7655 (N_7655,N_6358,N_6627);
and U7656 (N_7656,N_6276,N_6312);
xnor U7657 (N_7657,N_6759,N_6490);
nand U7658 (N_7658,N_6634,N_6889);
nor U7659 (N_7659,N_6323,N_6937);
xor U7660 (N_7660,N_6818,N_6194);
nand U7661 (N_7661,N_6141,N_6575);
and U7662 (N_7662,N_6019,N_6979);
xor U7663 (N_7663,N_6690,N_6253);
nor U7664 (N_7664,N_6777,N_6574);
xnor U7665 (N_7665,N_6713,N_6359);
xor U7666 (N_7666,N_6253,N_6754);
nor U7667 (N_7667,N_6067,N_6559);
xor U7668 (N_7668,N_6751,N_6107);
nor U7669 (N_7669,N_6594,N_6194);
or U7670 (N_7670,N_6629,N_6664);
and U7671 (N_7671,N_6779,N_6546);
or U7672 (N_7672,N_6502,N_6134);
nand U7673 (N_7673,N_6647,N_6982);
or U7674 (N_7674,N_6547,N_6833);
or U7675 (N_7675,N_6937,N_6713);
and U7676 (N_7676,N_6572,N_6130);
nand U7677 (N_7677,N_6549,N_6466);
nand U7678 (N_7678,N_6587,N_6949);
xnor U7679 (N_7679,N_6021,N_6956);
or U7680 (N_7680,N_6392,N_6108);
nor U7681 (N_7681,N_6483,N_6033);
nand U7682 (N_7682,N_6399,N_6016);
nor U7683 (N_7683,N_6781,N_6292);
xnor U7684 (N_7684,N_6062,N_6200);
or U7685 (N_7685,N_6031,N_6430);
or U7686 (N_7686,N_6694,N_6095);
nor U7687 (N_7687,N_6868,N_6961);
or U7688 (N_7688,N_6744,N_6252);
or U7689 (N_7689,N_6523,N_6811);
or U7690 (N_7690,N_6633,N_6281);
nor U7691 (N_7691,N_6782,N_6724);
or U7692 (N_7692,N_6560,N_6286);
nor U7693 (N_7693,N_6062,N_6715);
nor U7694 (N_7694,N_6645,N_6417);
nand U7695 (N_7695,N_6207,N_6703);
xor U7696 (N_7696,N_6524,N_6497);
nand U7697 (N_7697,N_6710,N_6183);
nand U7698 (N_7698,N_6570,N_6981);
or U7699 (N_7699,N_6471,N_6633);
and U7700 (N_7700,N_6429,N_6504);
and U7701 (N_7701,N_6276,N_6957);
xor U7702 (N_7702,N_6427,N_6725);
and U7703 (N_7703,N_6489,N_6412);
nor U7704 (N_7704,N_6660,N_6223);
nor U7705 (N_7705,N_6598,N_6761);
or U7706 (N_7706,N_6867,N_6454);
nand U7707 (N_7707,N_6779,N_6086);
and U7708 (N_7708,N_6092,N_6128);
nand U7709 (N_7709,N_6030,N_6748);
nor U7710 (N_7710,N_6525,N_6937);
and U7711 (N_7711,N_6718,N_6434);
and U7712 (N_7712,N_6257,N_6828);
and U7713 (N_7713,N_6117,N_6916);
nor U7714 (N_7714,N_6628,N_6775);
nor U7715 (N_7715,N_6915,N_6302);
nand U7716 (N_7716,N_6176,N_6134);
nor U7717 (N_7717,N_6254,N_6279);
or U7718 (N_7718,N_6605,N_6385);
xor U7719 (N_7719,N_6459,N_6045);
and U7720 (N_7720,N_6677,N_6791);
and U7721 (N_7721,N_6313,N_6122);
or U7722 (N_7722,N_6211,N_6204);
xnor U7723 (N_7723,N_6671,N_6370);
and U7724 (N_7724,N_6954,N_6694);
or U7725 (N_7725,N_6610,N_6746);
or U7726 (N_7726,N_6199,N_6524);
nor U7727 (N_7727,N_6430,N_6082);
or U7728 (N_7728,N_6156,N_6909);
or U7729 (N_7729,N_6158,N_6866);
or U7730 (N_7730,N_6773,N_6137);
xor U7731 (N_7731,N_6926,N_6998);
and U7732 (N_7732,N_6043,N_6577);
nand U7733 (N_7733,N_6999,N_6726);
nor U7734 (N_7734,N_6794,N_6178);
nor U7735 (N_7735,N_6076,N_6791);
nand U7736 (N_7736,N_6358,N_6265);
nand U7737 (N_7737,N_6452,N_6720);
nor U7738 (N_7738,N_6009,N_6584);
xnor U7739 (N_7739,N_6257,N_6233);
or U7740 (N_7740,N_6418,N_6799);
and U7741 (N_7741,N_6755,N_6535);
or U7742 (N_7742,N_6998,N_6465);
xor U7743 (N_7743,N_6156,N_6731);
nor U7744 (N_7744,N_6565,N_6886);
xor U7745 (N_7745,N_6523,N_6210);
xnor U7746 (N_7746,N_6381,N_6879);
xnor U7747 (N_7747,N_6522,N_6570);
and U7748 (N_7748,N_6682,N_6010);
nor U7749 (N_7749,N_6873,N_6206);
or U7750 (N_7750,N_6505,N_6049);
and U7751 (N_7751,N_6824,N_6604);
or U7752 (N_7752,N_6967,N_6245);
nand U7753 (N_7753,N_6414,N_6381);
and U7754 (N_7754,N_6998,N_6135);
or U7755 (N_7755,N_6679,N_6490);
nand U7756 (N_7756,N_6696,N_6036);
nor U7757 (N_7757,N_6594,N_6778);
or U7758 (N_7758,N_6109,N_6381);
or U7759 (N_7759,N_6786,N_6463);
xor U7760 (N_7760,N_6556,N_6180);
xnor U7761 (N_7761,N_6509,N_6797);
or U7762 (N_7762,N_6874,N_6801);
or U7763 (N_7763,N_6827,N_6764);
xor U7764 (N_7764,N_6599,N_6645);
nand U7765 (N_7765,N_6854,N_6630);
nand U7766 (N_7766,N_6356,N_6388);
and U7767 (N_7767,N_6841,N_6597);
and U7768 (N_7768,N_6318,N_6204);
xnor U7769 (N_7769,N_6890,N_6344);
and U7770 (N_7770,N_6640,N_6581);
or U7771 (N_7771,N_6969,N_6898);
nand U7772 (N_7772,N_6933,N_6122);
and U7773 (N_7773,N_6815,N_6200);
nor U7774 (N_7774,N_6287,N_6919);
nor U7775 (N_7775,N_6825,N_6047);
xnor U7776 (N_7776,N_6846,N_6491);
xor U7777 (N_7777,N_6662,N_6428);
nor U7778 (N_7778,N_6021,N_6435);
xnor U7779 (N_7779,N_6833,N_6242);
and U7780 (N_7780,N_6018,N_6560);
nand U7781 (N_7781,N_6603,N_6159);
nand U7782 (N_7782,N_6382,N_6337);
or U7783 (N_7783,N_6323,N_6938);
nor U7784 (N_7784,N_6604,N_6475);
xnor U7785 (N_7785,N_6334,N_6696);
nand U7786 (N_7786,N_6521,N_6032);
nand U7787 (N_7787,N_6238,N_6444);
nor U7788 (N_7788,N_6608,N_6966);
xor U7789 (N_7789,N_6901,N_6906);
and U7790 (N_7790,N_6623,N_6919);
nand U7791 (N_7791,N_6389,N_6680);
xnor U7792 (N_7792,N_6448,N_6515);
xor U7793 (N_7793,N_6166,N_6366);
and U7794 (N_7794,N_6353,N_6127);
xnor U7795 (N_7795,N_6760,N_6651);
nand U7796 (N_7796,N_6048,N_6576);
and U7797 (N_7797,N_6893,N_6095);
nor U7798 (N_7798,N_6612,N_6056);
or U7799 (N_7799,N_6015,N_6660);
xor U7800 (N_7800,N_6385,N_6587);
nor U7801 (N_7801,N_6596,N_6747);
nand U7802 (N_7802,N_6885,N_6110);
and U7803 (N_7803,N_6510,N_6389);
nor U7804 (N_7804,N_6799,N_6356);
nand U7805 (N_7805,N_6926,N_6247);
and U7806 (N_7806,N_6741,N_6833);
xnor U7807 (N_7807,N_6033,N_6323);
nand U7808 (N_7808,N_6122,N_6022);
nand U7809 (N_7809,N_6391,N_6692);
xor U7810 (N_7810,N_6839,N_6350);
xor U7811 (N_7811,N_6498,N_6561);
and U7812 (N_7812,N_6957,N_6429);
nor U7813 (N_7813,N_6533,N_6913);
and U7814 (N_7814,N_6646,N_6980);
nor U7815 (N_7815,N_6926,N_6760);
nor U7816 (N_7816,N_6998,N_6089);
or U7817 (N_7817,N_6533,N_6645);
nand U7818 (N_7818,N_6800,N_6558);
nand U7819 (N_7819,N_6808,N_6374);
nor U7820 (N_7820,N_6727,N_6851);
nand U7821 (N_7821,N_6125,N_6799);
xor U7822 (N_7822,N_6896,N_6985);
nor U7823 (N_7823,N_6395,N_6821);
nand U7824 (N_7824,N_6618,N_6525);
nand U7825 (N_7825,N_6463,N_6780);
nor U7826 (N_7826,N_6190,N_6678);
xor U7827 (N_7827,N_6936,N_6445);
xor U7828 (N_7828,N_6154,N_6387);
and U7829 (N_7829,N_6884,N_6004);
xnor U7830 (N_7830,N_6232,N_6138);
nor U7831 (N_7831,N_6405,N_6350);
and U7832 (N_7832,N_6262,N_6065);
nand U7833 (N_7833,N_6518,N_6719);
xnor U7834 (N_7834,N_6932,N_6409);
or U7835 (N_7835,N_6917,N_6232);
xnor U7836 (N_7836,N_6674,N_6240);
nor U7837 (N_7837,N_6075,N_6208);
and U7838 (N_7838,N_6815,N_6713);
nand U7839 (N_7839,N_6553,N_6799);
nand U7840 (N_7840,N_6489,N_6787);
and U7841 (N_7841,N_6791,N_6883);
and U7842 (N_7842,N_6145,N_6202);
nand U7843 (N_7843,N_6214,N_6352);
nor U7844 (N_7844,N_6385,N_6556);
or U7845 (N_7845,N_6830,N_6532);
xnor U7846 (N_7846,N_6458,N_6355);
nand U7847 (N_7847,N_6918,N_6550);
nor U7848 (N_7848,N_6769,N_6928);
nand U7849 (N_7849,N_6772,N_6263);
and U7850 (N_7850,N_6133,N_6452);
xor U7851 (N_7851,N_6229,N_6907);
nand U7852 (N_7852,N_6217,N_6458);
or U7853 (N_7853,N_6522,N_6652);
nand U7854 (N_7854,N_6775,N_6104);
or U7855 (N_7855,N_6110,N_6263);
xor U7856 (N_7856,N_6011,N_6338);
nand U7857 (N_7857,N_6940,N_6197);
and U7858 (N_7858,N_6152,N_6019);
or U7859 (N_7859,N_6622,N_6707);
nand U7860 (N_7860,N_6058,N_6072);
nor U7861 (N_7861,N_6187,N_6116);
and U7862 (N_7862,N_6877,N_6155);
or U7863 (N_7863,N_6179,N_6696);
xor U7864 (N_7864,N_6525,N_6559);
nand U7865 (N_7865,N_6416,N_6338);
and U7866 (N_7866,N_6345,N_6393);
xnor U7867 (N_7867,N_6463,N_6194);
nand U7868 (N_7868,N_6291,N_6643);
xor U7869 (N_7869,N_6203,N_6618);
nor U7870 (N_7870,N_6302,N_6172);
or U7871 (N_7871,N_6744,N_6472);
xor U7872 (N_7872,N_6083,N_6712);
or U7873 (N_7873,N_6665,N_6190);
and U7874 (N_7874,N_6839,N_6161);
xnor U7875 (N_7875,N_6474,N_6216);
nand U7876 (N_7876,N_6787,N_6847);
nor U7877 (N_7877,N_6317,N_6272);
xor U7878 (N_7878,N_6150,N_6024);
nand U7879 (N_7879,N_6262,N_6102);
xor U7880 (N_7880,N_6346,N_6465);
or U7881 (N_7881,N_6917,N_6748);
nand U7882 (N_7882,N_6101,N_6287);
or U7883 (N_7883,N_6936,N_6625);
xor U7884 (N_7884,N_6589,N_6990);
or U7885 (N_7885,N_6509,N_6414);
and U7886 (N_7886,N_6980,N_6924);
or U7887 (N_7887,N_6165,N_6421);
nand U7888 (N_7888,N_6346,N_6243);
and U7889 (N_7889,N_6389,N_6175);
or U7890 (N_7890,N_6476,N_6980);
xnor U7891 (N_7891,N_6516,N_6539);
or U7892 (N_7892,N_6793,N_6162);
nand U7893 (N_7893,N_6272,N_6273);
xnor U7894 (N_7894,N_6856,N_6759);
or U7895 (N_7895,N_6930,N_6267);
nand U7896 (N_7896,N_6586,N_6522);
or U7897 (N_7897,N_6536,N_6391);
nand U7898 (N_7898,N_6342,N_6545);
xor U7899 (N_7899,N_6690,N_6595);
and U7900 (N_7900,N_6135,N_6759);
nor U7901 (N_7901,N_6362,N_6237);
nor U7902 (N_7902,N_6525,N_6326);
xnor U7903 (N_7903,N_6196,N_6532);
nor U7904 (N_7904,N_6972,N_6103);
nand U7905 (N_7905,N_6803,N_6679);
nand U7906 (N_7906,N_6012,N_6187);
nor U7907 (N_7907,N_6698,N_6617);
xor U7908 (N_7908,N_6363,N_6205);
or U7909 (N_7909,N_6229,N_6736);
or U7910 (N_7910,N_6310,N_6417);
nor U7911 (N_7911,N_6843,N_6423);
xor U7912 (N_7912,N_6280,N_6672);
nand U7913 (N_7913,N_6440,N_6237);
xnor U7914 (N_7914,N_6120,N_6160);
xor U7915 (N_7915,N_6346,N_6411);
nand U7916 (N_7916,N_6208,N_6628);
and U7917 (N_7917,N_6396,N_6149);
nand U7918 (N_7918,N_6781,N_6667);
and U7919 (N_7919,N_6431,N_6729);
or U7920 (N_7920,N_6837,N_6347);
or U7921 (N_7921,N_6405,N_6664);
or U7922 (N_7922,N_6778,N_6135);
nor U7923 (N_7923,N_6232,N_6957);
or U7924 (N_7924,N_6819,N_6524);
nand U7925 (N_7925,N_6726,N_6603);
and U7926 (N_7926,N_6006,N_6351);
xor U7927 (N_7927,N_6263,N_6973);
and U7928 (N_7928,N_6040,N_6641);
or U7929 (N_7929,N_6666,N_6708);
xnor U7930 (N_7930,N_6908,N_6823);
nand U7931 (N_7931,N_6119,N_6597);
nor U7932 (N_7932,N_6142,N_6347);
xnor U7933 (N_7933,N_6186,N_6910);
nor U7934 (N_7934,N_6224,N_6899);
nand U7935 (N_7935,N_6008,N_6305);
or U7936 (N_7936,N_6257,N_6968);
nor U7937 (N_7937,N_6191,N_6976);
nor U7938 (N_7938,N_6422,N_6497);
nor U7939 (N_7939,N_6436,N_6790);
nand U7940 (N_7940,N_6538,N_6987);
nand U7941 (N_7941,N_6738,N_6858);
or U7942 (N_7942,N_6091,N_6423);
xor U7943 (N_7943,N_6064,N_6590);
nor U7944 (N_7944,N_6538,N_6602);
and U7945 (N_7945,N_6325,N_6434);
or U7946 (N_7946,N_6357,N_6028);
nand U7947 (N_7947,N_6498,N_6721);
nand U7948 (N_7948,N_6792,N_6727);
xnor U7949 (N_7949,N_6328,N_6173);
nor U7950 (N_7950,N_6189,N_6833);
nor U7951 (N_7951,N_6322,N_6922);
nand U7952 (N_7952,N_6704,N_6273);
nand U7953 (N_7953,N_6787,N_6980);
nor U7954 (N_7954,N_6285,N_6834);
and U7955 (N_7955,N_6215,N_6308);
or U7956 (N_7956,N_6376,N_6732);
nand U7957 (N_7957,N_6751,N_6822);
nor U7958 (N_7958,N_6732,N_6914);
and U7959 (N_7959,N_6712,N_6050);
or U7960 (N_7960,N_6188,N_6037);
or U7961 (N_7961,N_6390,N_6862);
nor U7962 (N_7962,N_6907,N_6637);
or U7963 (N_7963,N_6536,N_6340);
nand U7964 (N_7964,N_6269,N_6648);
nor U7965 (N_7965,N_6721,N_6973);
or U7966 (N_7966,N_6841,N_6499);
nor U7967 (N_7967,N_6897,N_6162);
xnor U7968 (N_7968,N_6584,N_6607);
or U7969 (N_7969,N_6945,N_6905);
and U7970 (N_7970,N_6519,N_6460);
or U7971 (N_7971,N_6082,N_6425);
and U7972 (N_7972,N_6361,N_6916);
nand U7973 (N_7973,N_6796,N_6098);
xor U7974 (N_7974,N_6884,N_6097);
xor U7975 (N_7975,N_6801,N_6638);
nor U7976 (N_7976,N_6377,N_6437);
nor U7977 (N_7977,N_6694,N_6872);
and U7978 (N_7978,N_6746,N_6392);
and U7979 (N_7979,N_6383,N_6876);
xnor U7980 (N_7980,N_6548,N_6843);
xnor U7981 (N_7981,N_6688,N_6765);
nor U7982 (N_7982,N_6557,N_6866);
xnor U7983 (N_7983,N_6732,N_6972);
nor U7984 (N_7984,N_6913,N_6165);
nor U7985 (N_7985,N_6498,N_6999);
or U7986 (N_7986,N_6670,N_6541);
and U7987 (N_7987,N_6227,N_6760);
or U7988 (N_7988,N_6627,N_6043);
or U7989 (N_7989,N_6186,N_6920);
xnor U7990 (N_7990,N_6647,N_6252);
nor U7991 (N_7991,N_6609,N_6766);
or U7992 (N_7992,N_6769,N_6516);
and U7993 (N_7993,N_6866,N_6520);
xor U7994 (N_7994,N_6703,N_6620);
nor U7995 (N_7995,N_6345,N_6023);
nor U7996 (N_7996,N_6388,N_6012);
nand U7997 (N_7997,N_6013,N_6505);
nand U7998 (N_7998,N_6158,N_6938);
xor U7999 (N_7999,N_6538,N_6082);
nor U8000 (N_8000,N_7966,N_7876);
nand U8001 (N_8001,N_7116,N_7925);
or U8002 (N_8002,N_7172,N_7680);
xnor U8003 (N_8003,N_7366,N_7639);
xor U8004 (N_8004,N_7110,N_7390);
or U8005 (N_8005,N_7891,N_7838);
xor U8006 (N_8006,N_7111,N_7258);
nand U8007 (N_8007,N_7482,N_7570);
and U8008 (N_8008,N_7311,N_7973);
xnor U8009 (N_8009,N_7862,N_7132);
xnor U8010 (N_8010,N_7606,N_7262);
xnor U8011 (N_8011,N_7629,N_7668);
and U8012 (N_8012,N_7193,N_7183);
and U8013 (N_8013,N_7267,N_7125);
and U8014 (N_8014,N_7766,N_7314);
nor U8015 (N_8015,N_7252,N_7104);
nand U8016 (N_8016,N_7481,N_7385);
nand U8017 (N_8017,N_7497,N_7760);
xnor U8018 (N_8018,N_7218,N_7148);
nand U8019 (N_8019,N_7233,N_7012);
xor U8020 (N_8020,N_7277,N_7329);
or U8021 (N_8021,N_7249,N_7100);
nand U8022 (N_8022,N_7750,N_7272);
nand U8023 (N_8023,N_7741,N_7586);
xor U8024 (N_8024,N_7685,N_7503);
and U8025 (N_8025,N_7230,N_7941);
xor U8026 (N_8026,N_7447,N_7227);
nand U8027 (N_8027,N_7664,N_7142);
and U8028 (N_8028,N_7770,N_7328);
xnor U8029 (N_8029,N_7800,N_7571);
nand U8030 (N_8030,N_7032,N_7356);
xor U8031 (N_8031,N_7495,N_7936);
or U8032 (N_8032,N_7200,N_7076);
nand U8033 (N_8033,N_7752,N_7202);
nor U8034 (N_8034,N_7715,N_7030);
nor U8035 (N_8035,N_7265,N_7212);
nand U8036 (N_8036,N_7278,N_7751);
nand U8037 (N_8037,N_7049,N_7374);
nand U8038 (N_8038,N_7687,N_7912);
xnor U8039 (N_8039,N_7705,N_7520);
xnor U8040 (N_8040,N_7960,N_7753);
or U8041 (N_8041,N_7341,N_7194);
nor U8042 (N_8042,N_7562,N_7785);
nand U8043 (N_8043,N_7247,N_7640);
nor U8044 (N_8044,N_7684,N_7820);
or U8045 (N_8045,N_7133,N_7152);
nand U8046 (N_8046,N_7602,N_7072);
nor U8047 (N_8047,N_7694,N_7942);
xnor U8048 (N_8048,N_7608,N_7355);
or U8049 (N_8049,N_7351,N_7555);
or U8050 (N_8050,N_7840,N_7138);
nand U8051 (N_8051,N_7628,N_7733);
xnor U8052 (N_8052,N_7932,N_7810);
or U8053 (N_8053,N_7963,N_7210);
xnor U8054 (N_8054,N_7830,N_7762);
nand U8055 (N_8055,N_7583,N_7509);
and U8056 (N_8056,N_7706,N_7746);
nor U8057 (N_8057,N_7655,N_7739);
and U8058 (N_8058,N_7396,N_7017);
nor U8059 (N_8059,N_7223,N_7834);
nor U8060 (N_8060,N_7057,N_7024);
nand U8061 (N_8061,N_7683,N_7412);
xor U8062 (N_8062,N_7018,N_7471);
nand U8063 (N_8063,N_7397,N_7920);
xor U8064 (N_8064,N_7808,N_7020);
or U8065 (N_8065,N_7547,N_7842);
nand U8066 (N_8066,N_7968,N_7381);
or U8067 (N_8067,N_7224,N_7044);
nand U8068 (N_8068,N_7540,N_7835);
nand U8069 (N_8069,N_7795,N_7059);
xnor U8070 (N_8070,N_7650,N_7423);
nor U8071 (N_8071,N_7198,N_7178);
nor U8072 (N_8072,N_7593,N_7204);
nor U8073 (N_8073,N_7535,N_7675);
xor U8074 (N_8074,N_7690,N_7263);
or U8075 (N_8075,N_7306,N_7500);
xnor U8076 (N_8076,N_7940,N_7274);
xor U8077 (N_8077,N_7275,N_7461);
xor U8078 (N_8078,N_7829,N_7765);
nand U8079 (N_8079,N_7358,N_7873);
xor U8080 (N_8080,N_7354,N_7574);
nor U8081 (N_8081,N_7863,N_7068);
or U8082 (N_8082,N_7435,N_7718);
or U8083 (N_8083,N_7793,N_7735);
and U8084 (N_8084,N_7549,N_7067);
xor U8085 (N_8085,N_7490,N_7162);
or U8086 (N_8086,N_7847,N_7015);
nand U8087 (N_8087,N_7334,N_7157);
and U8088 (N_8088,N_7708,N_7789);
nor U8089 (N_8089,N_7983,N_7081);
or U8090 (N_8090,N_7284,N_7082);
xor U8091 (N_8091,N_7895,N_7253);
xor U8092 (N_8092,N_7324,N_7465);
and U8093 (N_8093,N_7427,N_7295);
or U8094 (N_8094,N_7599,N_7717);
nor U8095 (N_8095,N_7483,N_7980);
xor U8096 (N_8096,N_7310,N_7248);
xnor U8097 (N_8097,N_7908,N_7170);
and U8098 (N_8098,N_7429,N_7995);
nand U8099 (N_8099,N_7950,N_7896);
or U8100 (N_8100,N_7117,N_7518);
nand U8101 (N_8101,N_7696,N_7965);
or U8102 (N_8102,N_7489,N_7097);
and U8103 (N_8103,N_7774,N_7945);
nand U8104 (N_8104,N_7949,N_7446);
or U8105 (N_8105,N_7373,N_7998);
nand U8106 (N_8106,N_7546,N_7644);
xnor U8107 (N_8107,N_7367,N_7177);
and U8108 (N_8108,N_7935,N_7181);
and U8109 (N_8109,N_7804,N_7618);
and U8110 (N_8110,N_7637,N_7330);
xnor U8111 (N_8111,N_7674,N_7442);
xnor U8112 (N_8112,N_7163,N_7221);
or U8113 (N_8113,N_7254,N_7126);
nor U8114 (N_8114,N_7313,N_7841);
or U8115 (N_8115,N_7066,N_7652);
nor U8116 (N_8116,N_7594,N_7927);
nand U8117 (N_8117,N_7409,N_7312);
xor U8118 (N_8118,N_7568,N_7837);
nor U8119 (N_8119,N_7089,N_7440);
xor U8120 (N_8120,N_7947,N_7062);
and U8121 (N_8121,N_7877,N_7276);
nor U8122 (N_8122,N_7058,N_7443);
xnor U8123 (N_8123,N_7332,N_7016);
or U8124 (N_8124,N_7289,N_7772);
nor U8125 (N_8125,N_7523,N_7286);
or U8126 (N_8126,N_7567,N_7937);
or U8127 (N_8127,N_7449,N_7850);
nand U8128 (N_8128,N_7144,N_7827);
nor U8129 (N_8129,N_7080,N_7986);
nor U8130 (N_8130,N_7643,N_7532);
xnor U8131 (N_8131,N_7236,N_7573);
or U8132 (N_8132,N_7971,N_7616);
nor U8133 (N_8133,N_7698,N_7205);
or U8134 (N_8134,N_7472,N_7216);
nand U8135 (N_8135,N_7119,N_7414);
nor U8136 (N_8136,N_7888,N_7638);
nor U8137 (N_8137,N_7634,N_7139);
nor U8138 (N_8138,N_7848,N_7817);
xor U8139 (N_8139,N_7892,N_7333);
or U8140 (N_8140,N_7102,N_7158);
and U8141 (N_8141,N_7768,N_7168);
or U8142 (N_8142,N_7558,N_7539);
and U8143 (N_8143,N_7781,N_7073);
or U8144 (N_8144,N_7240,N_7899);
nand U8145 (N_8145,N_7408,N_7069);
nor U8146 (N_8146,N_7999,N_7667);
xnor U8147 (N_8147,N_7498,N_7331);
or U8148 (N_8148,N_7444,N_7060);
nor U8149 (N_8149,N_7213,N_7607);
and U8150 (N_8150,N_7534,N_7734);
xnor U8151 (N_8151,N_7211,N_7467);
nand U8152 (N_8152,N_7861,N_7775);
xor U8153 (N_8153,N_7515,N_7430);
or U8154 (N_8154,N_7799,N_7384);
xnor U8155 (N_8155,N_7669,N_7419);
or U8156 (N_8156,N_7716,N_7186);
nand U8157 (N_8157,N_7225,N_7123);
nand U8158 (N_8158,N_7093,N_7340);
nand U8159 (N_8159,N_7577,N_7478);
nand U8160 (N_8160,N_7234,N_7411);
or U8161 (N_8161,N_7626,N_7761);
nand U8162 (N_8162,N_7630,N_7933);
or U8163 (N_8163,N_7600,N_7519);
or U8164 (N_8164,N_7953,N_7114);
nand U8165 (N_8165,N_7256,N_7245);
and U8166 (N_8166,N_7801,N_7951);
nor U8167 (N_8167,N_7352,N_7368);
nor U8168 (N_8168,N_7308,N_7543);
and U8169 (N_8169,N_7693,N_7002);
nand U8170 (N_8170,N_7372,N_7359);
nor U8171 (N_8171,N_7703,N_7536);
or U8172 (N_8172,N_7903,N_7271);
nor U8173 (N_8173,N_7450,N_7270);
xnor U8174 (N_8174,N_7242,N_7448);
and U8175 (N_8175,N_7962,N_7038);
nor U8176 (N_8176,N_7956,N_7174);
or U8177 (N_8177,N_7943,N_7764);
xor U8178 (N_8178,N_7851,N_7389);
and U8179 (N_8179,N_7169,N_7156);
or U8180 (N_8180,N_7217,N_7417);
or U8181 (N_8181,N_7106,N_7357);
nor U8182 (N_8182,N_7737,N_7679);
nand U8183 (N_8183,N_7197,N_7074);
nor U8184 (N_8184,N_7228,N_7078);
or U8185 (N_8185,N_7131,N_7985);
and U8186 (N_8186,N_7517,N_7610);
xor U8187 (N_8187,N_7410,N_7376);
nand U8188 (N_8188,N_7363,N_7437);
nor U8189 (N_8189,N_7635,N_7302);
nor U8190 (N_8190,N_7063,N_7548);
nor U8191 (N_8191,N_7917,N_7299);
xnor U8192 (N_8192,N_7296,N_7507);
or U8193 (N_8193,N_7115,N_7147);
nor U8194 (N_8194,N_7743,N_7886);
nand U8195 (N_8195,N_7130,N_7459);
nor U8196 (N_8196,N_7416,N_7480);
or U8197 (N_8197,N_7779,N_7611);
or U8198 (N_8198,N_7484,N_7113);
xor U8199 (N_8199,N_7974,N_7578);
and U8200 (N_8200,N_7151,N_7609);
or U8201 (N_8201,N_7661,N_7619);
or U8202 (N_8202,N_7391,N_7338);
and U8203 (N_8203,N_7499,N_7828);
or U8204 (N_8204,N_7784,N_7707);
nor U8205 (N_8205,N_7836,N_7400);
xnor U8206 (N_8206,N_7127,N_7882);
nand U8207 (N_8207,N_7526,N_7970);
or U8208 (N_8208,N_7524,N_7748);
nor U8209 (N_8209,N_7561,N_7369);
nand U8210 (N_8210,N_7294,N_7179);
nand U8211 (N_8211,N_7161,N_7878);
and U8212 (N_8212,N_7955,N_7273);
xor U8213 (N_8213,N_7788,N_7470);
or U8214 (N_8214,N_7348,N_7996);
and U8215 (N_8215,N_7452,N_7994);
or U8216 (N_8216,N_7572,N_7875);
xnor U8217 (N_8217,N_7129,N_7171);
xnor U8218 (N_8218,N_7720,N_7195);
and U8219 (N_8219,N_7627,N_7670);
nand U8220 (N_8220,N_7822,N_7782);
nand U8221 (N_8221,N_7689,N_7092);
and U8222 (N_8222,N_7426,N_7300);
or U8223 (N_8223,N_7118,N_7624);
and U8224 (N_8224,N_7463,N_7048);
or U8225 (N_8225,N_7033,N_7055);
and U8226 (N_8226,N_7006,N_7292);
nand U8227 (N_8227,N_7736,N_7290);
nor U8228 (N_8228,N_7921,N_7857);
or U8229 (N_8229,N_7466,N_7991);
nor U8230 (N_8230,N_7203,N_7406);
xnor U8231 (N_8231,N_7241,N_7037);
and U8232 (N_8232,N_7166,N_7107);
xor U8233 (N_8233,N_7349,N_7190);
or U8234 (N_8234,N_7283,N_7657);
and U8235 (N_8235,N_7432,N_7553);
xor U8236 (N_8236,N_7375,N_7167);
nor U8237 (N_8237,N_7554,N_7007);
nand U8238 (N_8238,N_7360,N_7528);
nor U8239 (N_8239,N_7053,N_7763);
nor U8240 (N_8240,N_7492,N_7317);
xor U8241 (N_8241,N_7454,N_7721);
nor U8242 (N_8242,N_7339,N_7154);
nand U8243 (N_8243,N_7320,N_7605);
nor U8244 (N_8244,N_7923,N_7196);
xnor U8245 (N_8245,N_7802,N_7336);
xnor U8246 (N_8246,N_7232,N_7914);
nor U8247 (N_8247,N_7948,N_7238);
or U8248 (N_8248,N_7709,N_7281);
xnor U8249 (N_8249,N_7821,N_7860);
nor U8250 (N_8250,N_7034,N_7259);
xnor U8251 (N_8251,N_7464,N_7054);
xor U8252 (N_8252,N_7135,N_7682);
xnor U8253 (N_8253,N_7486,N_7832);
nand U8254 (N_8254,N_7688,N_7910);
or U8255 (N_8255,N_7025,N_7858);
xor U8256 (N_8256,N_7806,N_7846);
nand U8257 (N_8257,N_7362,N_7907);
nor U8258 (N_8258,N_7405,N_7350);
nand U8259 (N_8259,N_7474,N_7323);
and U8260 (N_8260,N_7656,N_7392);
or U8261 (N_8261,N_7428,N_7279);
or U8262 (N_8262,N_7141,N_7394);
xnor U8263 (N_8263,N_7591,N_7601);
or U8264 (N_8264,N_7287,N_7512);
and U8265 (N_8265,N_7964,N_7872);
xor U8266 (N_8266,N_7859,N_7382);
nor U8267 (N_8267,N_7021,N_7590);
xor U8268 (N_8268,N_7431,N_7493);
nor U8269 (N_8269,N_7315,N_7187);
nor U8270 (N_8270,N_7456,N_7757);
and U8271 (N_8271,N_7407,N_7797);
nor U8272 (N_8272,N_7491,N_7645);
and U8273 (N_8273,N_7322,N_7815);
and U8274 (N_8274,N_7701,N_7383);
nand U8275 (N_8275,N_7508,N_7939);
nand U8276 (N_8276,N_7589,N_7958);
or U8277 (N_8277,N_7671,N_7900);
and U8278 (N_8278,N_7103,N_7337);
nand U8279 (N_8279,N_7672,N_7488);
and U8280 (N_8280,N_7377,N_7010);
nand U8281 (N_8281,N_7967,N_7393);
nor U8282 (N_8282,N_7987,N_7421);
nand U8283 (N_8283,N_7565,N_7754);
nor U8284 (N_8284,N_7079,N_7261);
xor U8285 (N_8285,N_7904,N_7959);
and U8286 (N_8286,N_7134,N_7767);
nor U8287 (N_8287,N_7098,N_7468);
or U8288 (N_8288,N_7013,N_7911);
or U8289 (N_8289,N_7087,N_7929);
nand U8290 (N_8290,N_7711,N_7487);
and U8291 (N_8291,N_7982,N_7622);
or U8292 (N_8292,N_7660,N_7327);
and U8293 (N_8293,N_7997,N_7731);
nor U8294 (N_8294,N_7288,N_7649);
or U8295 (N_8295,N_7854,N_7791);
or U8296 (N_8296,N_7365,N_7137);
nor U8297 (N_8297,N_7004,N_7293);
nor U8298 (N_8298,N_7291,N_7977);
nand U8299 (N_8299,N_7344,N_7511);
xnor U8300 (N_8300,N_7798,N_7051);
nor U8301 (N_8301,N_7812,N_7149);
or U8302 (N_8302,N_7124,N_7180);
xnor U8303 (N_8303,N_7208,N_7255);
nor U8304 (N_8304,N_7676,N_7918);
or U8305 (N_8305,N_7475,N_7961);
or U8306 (N_8306,N_7108,N_7266);
xnor U8307 (N_8307,N_7404,N_7109);
and U8308 (N_8308,N_7285,N_7871);
xor U8309 (N_8309,N_7112,N_7691);
xnor U8310 (N_8310,N_7244,N_7260);
nand U8311 (N_8311,N_7813,N_7563);
and U8312 (N_8312,N_7436,N_7192);
nand U8313 (N_8313,N_7831,N_7502);
xnor U8314 (N_8314,N_7335,N_7304);
nand U8315 (N_8315,N_7803,N_7325);
and U8316 (N_8316,N_7595,N_7870);
nor U8317 (N_8317,N_7864,N_7712);
nand U8318 (N_8318,N_7559,N_7919);
and U8319 (N_8319,N_7695,N_7457);
xnor U8320 (N_8320,N_7297,N_7237);
nand U8321 (N_8321,N_7642,N_7727);
and U8322 (N_8322,N_7251,N_7833);
nand U8323 (N_8323,N_7576,N_7105);
xor U8324 (N_8324,N_7207,N_7453);
nor U8325 (N_8325,N_7201,N_7399);
or U8326 (N_8326,N_7071,N_7506);
xnor U8327 (N_8327,N_7867,N_7476);
and U8328 (N_8328,N_7439,N_7975);
or U8329 (N_8329,N_7056,N_7972);
nor U8330 (N_8330,N_7542,N_7040);
xnor U8331 (N_8331,N_7501,N_7379);
nand U8332 (N_8332,N_7773,N_7413);
or U8333 (N_8333,N_7077,N_7922);
or U8334 (N_8334,N_7598,N_7386);
or U8335 (N_8335,N_7807,N_7269);
nand U8336 (N_8336,N_7868,N_7988);
nor U8337 (N_8337,N_7084,N_7301);
nor U8338 (N_8338,N_7726,N_7496);
and U8339 (N_8339,N_7564,N_7879);
xor U8340 (N_8340,N_7027,N_7853);
and U8341 (N_8341,N_7824,N_7028);
or U8342 (N_8342,N_7805,N_7665);
nor U8343 (N_8343,N_7615,N_7525);
or U8344 (N_8344,N_7845,N_7697);
or U8345 (N_8345,N_7155,N_7175);
or U8346 (N_8346,N_7226,N_7710);
nor U8347 (N_8347,N_7176,N_7915);
and U8348 (N_8348,N_7901,N_7632);
nand U8349 (N_8349,N_7597,N_7120);
nor U8350 (N_8350,N_7231,N_7732);
nand U8351 (N_8351,N_7445,N_7825);
or U8352 (N_8352,N_7905,N_7550);
nor U8353 (N_8353,N_7881,N_7462);
nand U8354 (N_8354,N_7658,N_7818);
xnor U8355 (N_8355,N_7094,N_7159);
xor U8356 (N_8356,N_7659,N_7378);
nor U8357 (N_8357,N_7003,N_7346);
nor U8358 (N_8358,N_7849,N_7938);
nor U8359 (N_8359,N_7019,N_7403);
or U8360 (N_8360,N_7722,N_7924);
nor U8361 (N_8361,N_7343,N_7000);
or U8362 (N_8362,N_7326,N_7046);
xnor U8363 (N_8363,N_7008,N_7052);
or U8364 (N_8364,N_7031,N_7099);
nor U8365 (N_8365,N_7724,N_7957);
and U8366 (N_8366,N_7744,N_7814);
xor U8367 (N_8367,N_7855,N_7036);
nand U8368 (N_8368,N_7001,N_7993);
and U8369 (N_8369,N_7264,N_7085);
nor U8370 (N_8370,N_7654,N_7388);
nor U8371 (N_8371,N_7902,N_7662);
nor U8372 (N_8372,N_7954,N_7641);
or U8373 (N_8373,N_7780,N_7364);
or U8374 (N_8374,N_7250,N_7064);
and U8375 (N_8375,N_7422,N_7979);
nor U8376 (N_8376,N_7786,N_7740);
xor U8377 (N_8377,N_7014,N_7566);
and U8378 (N_8378,N_7651,N_7747);
or U8379 (N_8379,N_7096,N_7199);
and U8380 (N_8380,N_7143,N_7719);
and U8381 (N_8381,N_7345,N_7856);
and U8382 (N_8382,N_7581,N_7298);
nor U8383 (N_8383,N_7646,N_7086);
nor U8384 (N_8384,N_7673,N_7229);
nand U8385 (N_8385,N_7700,N_7029);
nor U8386 (N_8386,N_7361,N_7580);
or U8387 (N_8387,N_7603,N_7946);
nor U8388 (N_8388,N_7235,N_7692);
nand U8389 (N_8389,N_7756,N_7926);
nor U8390 (N_8390,N_7887,N_7944);
xor U8391 (N_8391,N_7206,N_7796);
or U8392 (N_8392,N_7434,N_7579);
xnor U8393 (N_8393,N_7022,N_7755);
or U8394 (N_8394,N_7623,N_7494);
and U8395 (N_8395,N_7633,N_7090);
or U8396 (N_8396,N_7425,N_7794);
nand U8397 (N_8397,N_7184,N_7451);
nand U8398 (N_8398,N_7091,N_7749);
nand U8399 (N_8399,N_7189,N_7783);
xnor U8400 (N_8400,N_7560,N_7545);
nor U8401 (N_8401,N_7699,N_7121);
nor U8402 (N_8402,N_7164,N_7898);
xnor U8403 (N_8403,N_7424,N_7792);
nand U8404 (N_8404,N_7584,N_7460);
or U8405 (N_8405,N_7916,N_7844);
nand U8406 (N_8406,N_7575,N_7215);
xor U8407 (N_8407,N_7776,N_7614);
nor U8408 (N_8408,N_7894,N_7023);
and U8409 (N_8409,N_7730,N_7604);
and U8410 (N_8410,N_7398,N_7146);
xnor U8411 (N_8411,N_7913,N_7612);
or U8412 (N_8412,N_7045,N_7047);
nor U8413 (N_8413,N_7569,N_7647);
or U8414 (N_8414,N_7969,N_7625);
or U8415 (N_8415,N_7303,N_7243);
or U8416 (N_8416,N_7485,N_7433);
and U8417 (N_8417,N_7095,N_7582);
nand U8418 (N_8418,N_7257,N_7704);
or U8419 (N_8419,N_7530,N_7050);
or U8420 (N_8420,N_7522,N_7865);
xor U8421 (N_8421,N_7617,N_7771);
or U8422 (N_8422,N_7529,N_7042);
nand U8423 (N_8423,N_7897,N_7702);
and U8424 (N_8424,N_7280,N_7531);
nor U8425 (N_8425,N_7839,N_7819);
and U8426 (N_8426,N_7653,N_7883);
nor U8427 (N_8427,N_7738,N_7631);
nand U8428 (N_8428,N_7636,N_7928);
nor U8429 (N_8429,N_7136,N_7621);
and U8430 (N_8430,N_7347,N_7978);
or U8431 (N_8431,N_7874,N_7185);
xnor U8432 (N_8432,N_7686,N_7477);
and U8433 (N_8433,N_7989,N_7309);
nand U8434 (N_8434,N_7342,N_7976);
nor U8435 (N_8435,N_7930,N_7188);
xor U8436 (N_8436,N_7556,N_7663);
nor U8437 (N_8437,N_7852,N_7745);
xnor U8438 (N_8438,N_7984,N_7319);
nand U8439 (N_8439,N_7909,N_7043);
or U8440 (N_8440,N_7418,N_7811);
xnor U8441 (N_8441,N_7742,N_7415);
xor U8442 (N_8442,N_7214,N_7906);
xor U8443 (N_8443,N_7182,N_7026);
and U8444 (N_8444,N_7714,N_7039);
nand U8445 (N_8445,N_7934,N_7681);
xnor U8446 (N_8446,N_7981,N_7380);
and U8447 (N_8447,N_7401,N_7371);
nor U8448 (N_8448,N_7952,N_7826);
nand U8449 (N_8449,N_7713,N_7521);
and U8450 (N_8450,N_7441,N_7122);
xor U8451 (N_8451,N_7458,N_7551);
xnor U8452 (N_8452,N_7880,N_7843);
xnor U8453 (N_8453,N_7884,N_7552);
and U8454 (N_8454,N_7729,N_7885);
xor U8455 (N_8455,N_7035,N_7469);
or U8456 (N_8456,N_7011,N_7165);
or U8457 (N_8457,N_7239,N_7759);
nand U8458 (N_8458,N_7395,N_7479);
xor U8459 (N_8459,N_7544,N_7889);
nor U8460 (N_8460,N_7220,N_7990);
and U8461 (N_8461,N_7070,N_7769);
nor U8462 (N_8462,N_7402,N_7538);
xor U8463 (N_8463,N_7931,N_7128);
and U8464 (N_8464,N_7787,N_7173);
or U8465 (N_8465,N_7219,N_7140);
nand U8466 (N_8466,N_7101,N_7005);
nor U8467 (N_8467,N_7585,N_7209);
and U8468 (N_8468,N_7678,N_7541);
or U8469 (N_8469,N_7592,N_7307);
or U8470 (N_8470,N_7725,N_7222);
nor U8471 (N_8471,N_7305,N_7083);
nand U8472 (N_8472,N_7648,N_7088);
or U8473 (N_8473,N_7588,N_7516);
or U8474 (N_8474,N_7387,N_7473);
nand U8475 (N_8475,N_7370,N_7510);
nor U8476 (N_8476,N_7150,N_7777);
nand U8477 (N_8477,N_7455,N_7992);
and U8478 (N_8478,N_7268,N_7505);
and U8479 (N_8479,N_7282,N_7318);
xnor U8480 (N_8480,N_7145,N_7758);
or U8481 (N_8481,N_7075,N_7160);
or U8482 (N_8482,N_7041,N_7153);
nor U8483 (N_8483,N_7061,N_7321);
or U8484 (N_8484,N_7866,N_7514);
xor U8485 (N_8485,N_7587,N_7316);
and U8486 (N_8486,N_7728,N_7513);
xor U8487 (N_8487,N_7666,N_7009);
xor U8488 (N_8488,N_7613,N_7869);
nand U8489 (N_8489,N_7533,N_7246);
nor U8490 (N_8490,N_7823,N_7527);
or U8491 (N_8491,N_7809,N_7537);
or U8492 (N_8492,N_7778,N_7191);
xor U8493 (N_8493,N_7504,N_7790);
nor U8494 (N_8494,N_7065,N_7816);
nand U8495 (N_8495,N_7438,N_7677);
xnor U8496 (N_8496,N_7890,N_7353);
nor U8497 (N_8497,N_7596,N_7723);
or U8498 (N_8498,N_7620,N_7893);
nand U8499 (N_8499,N_7557,N_7420);
nor U8500 (N_8500,N_7427,N_7303);
or U8501 (N_8501,N_7097,N_7979);
and U8502 (N_8502,N_7648,N_7534);
or U8503 (N_8503,N_7887,N_7880);
nand U8504 (N_8504,N_7731,N_7551);
and U8505 (N_8505,N_7077,N_7980);
and U8506 (N_8506,N_7382,N_7493);
or U8507 (N_8507,N_7712,N_7783);
nand U8508 (N_8508,N_7478,N_7128);
and U8509 (N_8509,N_7217,N_7064);
nor U8510 (N_8510,N_7745,N_7684);
nand U8511 (N_8511,N_7174,N_7537);
and U8512 (N_8512,N_7456,N_7214);
nor U8513 (N_8513,N_7401,N_7535);
nand U8514 (N_8514,N_7339,N_7871);
or U8515 (N_8515,N_7537,N_7614);
or U8516 (N_8516,N_7545,N_7659);
xnor U8517 (N_8517,N_7381,N_7000);
nand U8518 (N_8518,N_7554,N_7659);
nor U8519 (N_8519,N_7168,N_7825);
nor U8520 (N_8520,N_7329,N_7234);
or U8521 (N_8521,N_7965,N_7827);
or U8522 (N_8522,N_7920,N_7059);
nand U8523 (N_8523,N_7051,N_7116);
nor U8524 (N_8524,N_7383,N_7996);
xor U8525 (N_8525,N_7736,N_7297);
nor U8526 (N_8526,N_7993,N_7326);
xnor U8527 (N_8527,N_7600,N_7243);
nor U8528 (N_8528,N_7717,N_7293);
xnor U8529 (N_8529,N_7709,N_7734);
nor U8530 (N_8530,N_7044,N_7842);
or U8531 (N_8531,N_7080,N_7721);
nand U8532 (N_8532,N_7538,N_7579);
nor U8533 (N_8533,N_7416,N_7362);
nor U8534 (N_8534,N_7621,N_7431);
nand U8535 (N_8535,N_7364,N_7288);
or U8536 (N_8536,N_7390,N_7636);
xor U8537 (N_8537,N_7966,N_7491);
or U8538 (N_8538,N_7526,N_7930);
nand U8539 (N_8539,N_7565,N_7832);
or U8540 (N_8540,N_7392,N_7675);
or U8541 (N_8541,N_7014,N_7234);
nor U8542 (N_8542,N_7412,N_7992);
or U8543 (N_8543,N_7731,N_7209);
and U8544 (N_8544,N_7049,N_7197);
nor U8545 (N_8545,N_7159,N_7956);
and U8546 (N_8546,N_7471,N_7925);
or U8547 (N_8547,N_7020,N_7720);
or U8548 (N_8548,N_7454,N_7443);
xnor U8549 (N_8549,N_7653,N_7122);
or U8550 (N_8550,N_7009,N_7486);
nand U8551 (N_8551,N_7392,N_7571);
nand U8552 (N_8552,N_7413,N_7928);
nand U8553 (N_8553,N_7789,N_7728);
xor U8554 (N_8554,N_7870,N_7140);
or U8555 (N_8555,N_7523,N_7248);
nand U8556 (N_8556,N_7274,N_7115);
nand U8557 (N_8557,N_7531,N_7387);
xnor U8558 (N_8558,N_7692,N_7996);
and U8559 (N_8559,N_7921,N_7183);
and U8560 (N_8560,N_7087,N_7095);
nand U8561 (N_8561,N_7215,N_7803);
nor U8562 (N_8562,N_7828,N_7212);
or U8563 (N_8563,N_7500,N_7415);
or U8564 (N_8564,N_7397,N_7368);
nand U8565 (N_8565,N_7549,N_7665);
and U8566 (N_8566,N_7332,N_7060);
and U8567 (N_8567,N_7358,N_7748);
or U8568 (N_8568,N_7920,N_7211);
or U8569 (N_8569,N_7903,N_7557);
nand U8570 (N_8570,N_7197,N_7040);
and U8571 (N_8571,N_7436,N_7865);
nor U8572 (N_8572,N_7290,N_7472);
nor U8573 (N_8573,N_7189,N_7086);
nand U8574 (N_8574,N_7281,N_7457);
or U8575 (N_8575,N_7938,N_7513);
and U8576 (N_8576,N_7660,N_7754);
xor U8577 (N_8577,N_7034,N_7990);
or U8578 (N_8578,N_7319,N_7863);
and U8579 (N_8579,N_7991,N_7060);
and U8580 (N_8580,N_7134,N_7669);
or U8581 (N_8581,N_7693,N_7725);
nand U8582 (N_8582,N_7233,N_7941);
and U8583 (N_8583,N_7158,N_7681);
nor U8584 (N_8584,N_7116,N_7726);
xor U8585 (N_8585,N_7141,N_7989);
or U8586 (N_8586,N_7408,N_7172);
nor U8587 (N_8587,N_7392,N_7584);
xnor U8588 (N_8588,N_7069,N_7813);
nor U8589 (N_8589,N_7404,N_7224);
xor U8590 (N_8590,N_7447,N_7912);
nand U8591 (N_8591,N_7759,N_7496);
and U8592 (N_8592,N_7319,N_7762);
or U8593 (N_8593,N_7663,N_7040);
nor U8594 (N_8594,N_7176,N_7289);
xor U8595 (N_8595,N_7962,N_7789);
nand U8596 (N_8596,N_7825,N_7068);
nor U8597 (N_8597,N_7313,N_7143);
nor U8598 (N_8598,N_7873,N_7313);
or U8599 (N_8599,N_7350,N_7308);
nor U8600 (N_8600,N_7435,N_7991);
or U8601 (N_8601,N_7967,N_7595);
nand U8602 (N_8602,N_7085,N_7234);
or U8603 (N_8603,N_7715,N_7000);
nand U8604 (N_8604,N_7329,N_7772);
nand U8605 (N_8605,N_7444,N_7482);
nor U8606 (N_8606,N_7146,N_7482);
and U8607 (N_8607,N_7345,N_7515);
xor U8608 (N_8608,N_7776,N_7674);
nor U8609 (N_8609,N_7742,N_7481);
or U8610 (N_8610,N_7091,N_7839);
nand U8611 (N_8611,N_7576,N_7687);
nor U8612 (N_8612,N_7081,N_7321);
nand U8613 (N_8613,N_7592,N_7580);
or U8614 (N_8614,N_7199,N_7832);
nand U8615 (N_8615,N_7407,N_7105);
nor U8616 (N_8616,N_7143,N_7204);
xor U8617 (N_8617,N_7942,N_7283);
nor U8618 (N_8618,N_7329,N_7461);
nand U8619 (N_8619,N_7793,N_7373);
and U8620 (N_8620,N_7813,N_7112);
and U8621 (N_8621,N_7048,N_7455);
or U8622 (N_8622,N_7938,N_7423);
or U8623 (N_8623,N_7262,N_7971);
and U8624 (N_8624,N_7471,N_7558);
or U8625 (N_8625,N_7665,N_7976);
xnor U8626 (N_8626,N_7978,N_7542);
nand U8627 (N_8627,N_7137,N_7851);
or U8628 (N_8628,N_7685,N_7763);
xnor U8629 (N_8629,N_7471,N_7001);
nand U8630 (N_8630,N_7616,N_7658);
or U8631 (N_8631,N_7401,N_7852);
or U8632 (N_8632,N_7297,N_7093);
and U8633 (N_8633,N_7666,N_7369);
or U8634 (N_8634,N_7363,N_7190);
nand U8635 (N_8635,N_7817,N_7130);
nor U8636 (N_8636,N_7092,N_7101);
and U8637 (N_8637,N_7287,N_7756);
and U8638 (N_8638,N_7462,N_7577);
or U8639 (N_8639,N_7846,N_7674);
nor U8640 (N_8640,N_7222,N_7683);
xor U8641 (N_8641,N_7167,N_7901);
xor U8642 (N_8642,N_7069,N_7833);
nand U8643 (N_8643,N_7851,N_7233);
nor U8644 (N_8644,N_7721,N_7619);
nor U8645 (N_8645,N_7665,N_7018);
nor U8646 (N_8646,N_7769,N_7541);
and U8647 (N_8647,N_7898,N_7662);
and U8648 (N_8648,N_7218,N_7294);
nor U8649 (N_8649,N_7171,N_7477);
nor U8650 (N_8650,N_7734,N_7817);
nand U8651 (N_8651,N_7801,N_7605);
xnor U8652 (N_8652,N_7133,N_7597);
or U8653 (N_8653,N_7833,N_7244);
nor U8654 (N_8654,N_7639,N_7966);
nor U8655 (N_8655,N_7542,N_7999);
nand U8656 (N_8656,N_7547,N_7007);
and U8657 (N_8657,N_7899,N_7103);
nor U8658 (N_8658,N_7039,N_7033);
xnor U8659 (N_8659,N_7981,N_7305);
nand U8660 (N_8660,N_7058,N_7553);
nor U8661 (N_8661,N_7095,N_7162);
and U8662 (N_8662,N_7478,N_7008);
or U8663 (N_8663,N_7109,N_7078);
and U8664 (N_8664,N_7420,N_7461);
or U8665 (N_8665,N_7260,N_7096);
nor U8666 (N_8666,N_7361,N_7516);
nand U8667 (N_8667,N_7166,N_7215);
xor U8668 (N_8668,N_7563,N_7280);
and U8669 (N_8669,N_7315,N_7872);
and U8670 (N_8670,N_7473,N_7883);
or U8671 (N_8671,N_7691,N_7849);
nor U8672 (N_8672,N_7221,N_7630);
or U8673 (N_8673,N_7703,N_7632);
nor U8674 (N_8674,N_7836,N_7674);
xor U8675 (N_8675,N_7622,N_7389);
nor U8676 (N_8676,N_7698,N_7508);
or U8677 (N_8677,N_7553,N_7196);
or U8678 (N_8678,N_7595,N_7219);
and U8679 (N_8679,N_7988,N_7395);
nor U8680 (N_8680,N_7743,N_7782);
or U8681 (N_8681,N_7042,N_7248);
and U8682 (N_8682,N_7017,N_7297);
nor U8683 (N_8683,N_7777,N_7036);
xor U8684 (N_8684,N_7901,N_7932);
and U8685 (N_8685,N_7838,N_7794);
nand U8686 (N_8686,N_7952,N_7771);
nand U8687 (N_8687,N_7363,N_7895);
nor U8688 (N_8688,N_7502,N_7866);
nor U8689 (N_8689,N_7692,N_7084);
and U8690 (N_8690,N_7796,N_7483);
or U8691 (N_8691,N_7077,N_7611);
nand U8692 (N_8692,N_7171,N_7616);
nand U8693 (N_8693,N_7117,N_7497);
nand U8694 (N_8694,N_7953,N_7417);
xor U8695 (N_8695,N_7153,N_7168);
or U8696 (N_8696,N_7716,N_7516);
and U8697 (N_8697,N_7383,N_7421);
nand U8698 (N_8698,N_7302,N_7526);
xnor U8699 (N_8699,N_7367,N_7128);
nor U8700 (N_8700,N_7372,N_7288);
nand U8701 (N_8701,N_7247,N_7403);
or U8702 (N_8702,N_7608,N_7941);
and U8703 (N_8703,N_7333,N_7854);
or U8704 (N_8704,N_7291,N_7695);
nand U8705 (N_8705,N_7546,N_7737);
xor U8706 (N_8706,N_7657,N_7768);
nor U8707 (N_8707,N_7207,N_7163);
or U8708 (N_8708,N_7110,N_7796);
or U8709 (N_8709,N_7977,N_7201);
or U8710 (N_8710,N_7600,N_7619);
and U8711 (N_8711,N_7135,N_7902);
xnor U8712 (N_8712,N_7542,N_7415);
nand U8713 (N_8713,N_7296,N_7077);
or U8714 (N_8714,N_7410,N_7603);
nand U8715 (N_8715,N_7071,N_7948);
nor U8716 (N_8716,N_7295,N_7682);
xor U8717 (N_8717,N_7279,N_7103);
xnor U8718 (N_8718,N_7882,N_7707);
xor U8719 (N_8719,N_7267,N_7639);
nor U8720 (N_8720,N_7116,N_7984);
xnor U8721 (N_8721,N_7604,N_7713);
or U8722 (N_8722,N_7381,N_7333);
nor U8723 (N_8723,N_7656,N_7202);
xor U8724 (N_8724,N_7156,N_7802);
or U8725 (N_8725,N_7331,N_7047);
nor U8726 (N_8726,N_7518,N_7013);
or U8727 (N_8727,N_7969,N_7759);
or U8728 (N_8728,N_7582,N_7846);
nor U8729 (N_8729,N_7532,N_7383);
nand U8730 (N_8730,N_7927,N_7600);
xor U8731 (N_8731,N_7605,N_7626);
or U8732 (N_8732,N_7864,N_7054);
xnor U8733 (N_8733,N_7858,N_7694);
or U8734 (N_8734,N_7057,N_7485);
or U8735 (N_8735,N_7085,N_7216);
nor U8736 (N_8736,N_7694,N_7040);
or U8737 (N_8737,N_7088,N_7810);
xor U8738 (N_8738,N_7919,N_7839);
or U8739 (N_8739,N_7923,N_7134);
nand U8740 (N_8740,N_7113,N_7853);
and U8741 (N_8741,N_7499,N_7754);
nor U8742 (N_8742,N_7446,N_7895);
and U8743 (N_8743,N_7616,N_7230);
nand U8744 (N_8744,N_7390,N_7781);
and U8745 (N_8745,N_7547,N_7611);
and U8746 (N_8746,N_7087,N_7216);
nand U8747 (N_8747,N_7693,N_7402);
or U8748 (N_8748,N_7111,N_7301);
xnor U8749 (N_8749,N_7512,N_7887);
and U8750 (N_8750,N_7819,N_7364);
xor U8751 (N_8751,N_7162,N_7414);
xor U8752 (N_8752,N_7814,N_7296);
xnor U8753 (N_8753,N_7698,N_7935);
xor U8754 (N_8754,N_7424,N_7864);
nand U8755 (N_8755,N_7849,N_7038);
nor U8756 (N_8756,N_7565,N_7321);
nand U8757 (N_8757,N_7171,N_7291);
nor U8758 (N_8758,N_7275,N_7560);
nor U8759 (N_8759,N_7803,N_7025);
and U8760 (N_8760,N_7609,N_7671);
and U8761 (N_8761,N_7094,N_7333);
nand U8762 (N_8762,N_7070,N_7228);
or U8763 (N_8763,N_7002,N_7820);
nand U8764 (N_8764,N_7345,N_7844);
nor U8765 (N_8765,N_7368,N_7066);
and U8766 (N_8766,N_7833,N_7035);
nand U8767 (N_8767,N_7551,N_7068);
or U8768 (N_8768,N_7497,N_7784);
and U8769 (N_8769,N_7330,N_7985);
nor U8770 (N_8770,N_7857,N_7272);
or U8771 (N_8771,N_7449,N_7298);
nand U8772 (N_8772,N_7626,N_7935);
nor U8773 (N_8773,N_7840,N_7709);
xnor U8774 (N_8774,N_7864,N_7565);
nor U8775 (N_8775,N_7569,N_7979);
or U8776 (N_8776,N_7493,N_7005);
xnor U8777 (N_8777,N_7460,N_7753);
nand U8778 (N_8778,N_7377,N_7262);
nand U8779 (N_8779,N_7191,N_7634);
or U8780 (N_8780,N_7324,N_7344);
or U8781 (N_8781,N_7969,N_7007);
xnor U8782 (N_8782,N_7252,N_7754);
nand U8783 (N_8783,N_7200,N_7415);
xor U8784 (N_8784,N_7117,N_7866);
nand U8785 (N_8785,N_7716,N_7618);
nor U8786 (N_8786,N_7296,N_7076);
nor U8787 (N_8787,N_7242,N_7512);
nand U8788 (N_8788,N_7052,N_7236);
xnor U8789 (N_8789,N_7690,N_7816);
or U8790 (N_8790,N_7347,N_7441);
or U8791 (N_8791,N_7456,N_7097);
and U8792 (N_8792,N_7104,N_7092);
or U8793 (N_8793,N_7919,N_7335);
or U8794 (N_8794,N_7417,N_7048);
nand U8795 (N_8795,N_7334,N_7261);
and U8796 (N_8796,N_7084,N_7139);
nor U8797 (N_8797,N_7279,N_7997);
or U8798 (N_8798,N_7819,N_7795);
nor U8799 (N_8799,N_7076,N_7443);
nand U8800 (N_8800,N_7045,N_7504);
xnor U8801 (N_8801,N_7153,N_7294);
or U8802 (N_8802,N_7923,N_7583);
nor U8803 (N_8803,N_7804,N_7679);
xor U8804 (N_8804,N_7421,N_7761);
nor U8805 (N_8805,N_7402,N_7941);
nand U8806 (N_8806,N_7267,N_7253);
nor U8807 (N_8807,N_7168,N_7756);
nand U8808 (N_8808,N_7329,N_7526);
or U8809 (N_8809,N_7720,N_7302);
and U8810 (N_8810,N_7346,N_7736);
and U8811 (N_8811,N_7727,N_7368);
and U8812 (N_8812,N_7584,N_7650);
xnor U8813 (N_8813,N_7181,N_7227);
nor U8814 (N_8814,N_7262,N_7160);
nand U8815 (N_8815,N_7887,N_7563);
nor U8816 (N_8816,N_7290,N_7721);
xor U8817 (N_8817,N_7078,N_7877);
xor U8818 (N_8818,N_7552,N_7608);
or U8819 (N_8819,N_7442,N_7881);
nand U8820 (N_8820,N_7521,N_7449);
or U8821 (N_8821,N_7920,N_7931);
or U8822 (N_8822,N_7855,N_7579);
nand U8823 (N_8823,N_7106,N_7658);
nor U8824 (N_8824,N_7205,N_7735);
and U8825 (N_8825,N_7332,N_7018);
nand U8826 (N_8826,N_7461,N_7749);
and U8827 (N_8827,N_7145,N_7940);
and U8828 (N_8828,N_7704,N_7036);
or U8829 (N_8829,N_7015,N_7159);
or U8830 (N_8830,N_7116,N_7793);
nor U8831 (N_8831,N_7517,N_7698);
xor U8832 (N_8832,N_7853,N_7404);
and U8833 (N_8833,N_7907,N_7957);
nand U8834 (N_8834,N_7937,N_7261);
xor U8835 (N_8835,N_7369,N_7818);
xnor U8836 (N_8836,N_7012,N_7462);
or U8837 (N_8837,N_7673,N_7175);
nor U8838 (N_8838,N_7483,N_7293);
or U8839 (N_8839,N_7438,N_7602);
and U8840 (N_8840,N_7779,N_7277);
and U8841 (N_8841,N_7842,N_7550);
nand U8842 (N_8842,N_7066,N_7876);
or U8843 (N_8843,N_7410,N_7331);
or U8844 (N_8844,N_7835,N_7216);
nor U8845 (N_8845,N_7986,N_7745);
and U8846 (N_8846,N_7602,N_7244);
xor U8847 (N_8847,N_7028,N_7945);
nor U8848 (N_8848,N_7011,N_7751);
nand U8849 (N_8849,N_7389,N_7231);
or U8850 (N_8850,N_7083,N_7925);
nand U8851 (N_8851,N_7255,N_7114);
and U8852 (N_8852,N_7522,N_7956);
xor U8853 (N_8853,N_7924,N_7022);
nand U8854 (N_8854,N_7254,N_7428);
nand U8855 (N_8855,N_7315,N_7602);
nand U8856 (N_8856,N_7733,N_7606);
xnor U8857 (N_8857,N_7899,N_7877);
nor U8858 (N_8858,N_7715,N_7410);
or U8859 (N_8859,N_7237,N_7282);
and U8860 (N_8860,N_7009,N_7169);
nor U8861 (N_8861,N_7244,N_7521);
nand U8862 (N_8862,N_7665,N_7168);
or U8863 (N_8863,N_7329,N_7703);
xor U8864 (N_8864,N_7347,N_7704);
or U8865 (N_8865,N_7646,N_7996);
nor U8866 (N_8866,N_7773,N_7359);
or U8867 (N_8867,N_7192,N_7161);
and U8868 (N_8868,N_7293,N_7768);
nand U8869 (N_8869,N_7266,N_7407);
and U8870 (N_8870,N_7660,N_7084);
or U8871 (N_8871,N_7922,N_7133);
nor U8872 (N_8872,N_7956,N_7368);
or U8873 (N_8873,N_7287,N_7215);
nor U8874 (N_8874,N_7531,N_7086);
xnor U8875 (N_8875,N_7416,N_7154);
or U8876 (N_8876,N_7665,N_7704);
nor U8877 (N_8877,N_7868,N_7008);
xor U8878 (N_8878,N_7051,N_7010);
nor U8879 (N_8879,N_7829,N_7861);
nor U8880 (N_8880,N_7454,N_7044);
and U8881 (N_8881,N_7071,N_7419);
and U8882 (N_8882,N_7468,N_7187);
nand U8883 (N_8883,N_7845,N_7787);
nor U8884 (N_8884,N_7285,N_7562);
nor U8885 (N_8885,N_7241,N_7306);
and U8886 (N_8886,N_7650,N_7192);
or U8887 (N_8887,N_7809,N_7876);
nor U8888 (N_8888,N_7710,N_7008);
and U8889 (N_8889,N_7801,N_7950);
xnor U8890 (N_8890,N_7375,N_7966);
or U8891 (N_8891,N_7450,N_7986);
or U8892 (N_8892,N_7676,N_7126);
or U8893 (N_8893,N_7541,N_7868);
nor U8894 (N_8894,N_7049,N_7597);
xnor U8895 (N_8895,N_7979,N_7008);
xnor U8896 (N_8896,N_7509,N_7852);
nor U8897 (N_8897,N_7779,N_7585);
xor U8898 (N_8898,N_7411,N_7907);
and U8899 (N_8899,N_7575,N_7767);
nor U8900 (N_8900,N_7624,N_7004);
nand U8901 (N_8901,N_7937,N_7676);
and U8902 (N_8902,N_7836,N_7212);
nand U8903 (N_8903,N_7601,N_7203);
nor U8904 (N_8904,N_7955,N_7723);
nor U8905 (N_8905,N_7584,N_7246);
nand U8906 (N_8906,N_7919,N_7703);
nand U8907 (N_8907,N_7248,N_7295);
nor U8908 (N_8908,N_7120,N_7059);
or U8909 (N_8909,N_7272,N_7934);
and U8910 (N_8910,N_7273,N_7843);
xnor U8911 (N_8911,N_7811,N_7716);
nand U8912 (N_8912,N_7218,N_7483);
nand U8913 (N_8913,N_7003,N_7076);
xor U8914 (N_8914,N_7931,N_7763);
or U8915 (N_8915,N_7712,N_7808);
xor U8916 (N_8916,N_7451,N_7667);
or U8917 (N_8917,N_7359,N_7329);
nor U8918 (N_8918,N_7128,N_7674);
nand U8919 (N_8919,N_7867,N_7736);
nor U8920 (N_8920,N_7497,N_7214);
nand U8921 (N_8921,N_7433,N_7284);
nand U8922 (N_8922,N_7054,N_7481);
nor U8923 (N_8923,N_7810,N_7839);
and U8924 (N_8924,N_7722,N_7149);
nor U8925 (N_8925,N_7121,N_7802);
or U8926 (N_8926,N_7963,N_7594);
nand U8927 (N_8927,N_7300,N_7288);
nand U8928 (N_8928,N_7633,N_7645);
nor U8929 (N_8929,N_7387,N_7079);
nand U8930 (N_8930,N_7577,N_7109);
nor U8931 (N_8931,N_7991,N_7823);
or U8932 (N_8932,N_7019,N_7959);
nor U8933 (N_8933,N_7502,N_7861);
xnor U8934 (N_8934,N_7717,N_7286);
or U8935 (N_8935,N_7920,N_7409);
or U8936 (N_8936,N_7509,N_7385);
xor U8937 (N_8937,N_7015,N_7452);
and U8938 (N_8938,N_7154,N_7866);
and U8939 (N_8939,N_7410,N_7743);
or U8940 (N_8940,N_7633,N_7141);
nor U8941 (N_8941,N_7464,N_7413);
and U8942 (N_8942,N_7130,N_7295);
or U8943 (N_8943,N_7753,N_7074);
xor U8944 (N_8944,N_7685,N_7519);
or U8945 (N_8945,N_7567,N_7804);
nor U8946 (N_8946,N_7151,N_7968);
xnor U8947 (N_8947,N_7984,N_7178);
nand U8948 (N_8948,N_7938,N_7129);
and U8949 (N_8949,N_7171,N_7118);
nand U8950 (N_8950,N_7981,N_7843);
and U8951 (N_8951,N_7862,N_7697);
and U8952 (N_8952,N_7156,N_7879);
or U8953 (N_8953,N_7720,N_7430);
or U8954 (N_8954,N_7064,N_7952);
and U8955 (N_8955,N_7393,N_7925);
and U8956 (N_8956,N_7125,N_7105);
xnor U8957 (N_8957,N_7259,N_7724);
and U8958 (N_8958,N_7647,N_7025);
xor U8959 (N_8959,N_7723,N_7771);
nor U8960 (N_8960,N_7374,N_7848);
nor U8961 (N_8961,N_7930,N_7443);
nor U8962 (N_8962,N_7694,N_7820);
nor U8963 (N_8963,N_7716,N_7962);
and U8964 (N_8964,N_7026,N_7766);
nand U8965 (N_8965,N_7831,N_7915);
xnor U8966 (N_8966,N_7715,N_7743);
xnor U8967 (N_8967,N_7991,N_7873);
nand U8968 (N_8968,N_7252,N_7982);
nand U8969 (N_8969,N_7335,N_7461);
xnor U8970 (N_8970,N_7464,N_7258);
nor U8971 (N_8971,N_7472,N_7662);
and U8972 (N_8972,N_7354,N_7796);
or U8973 (N_8973,N_7468,N_7425);
and U8974 (N_8974,N_7065,N_7033);
and U8975 (N_8975,N_7267,N_7525);
nand U8976 (N_8976,N_7150,N_7370);
and U8977 (N_8977,N_7763,N_7637);
nand U8978 (N_8978,N_7540,N_7237);
nor U8979 (N_8979,N_7755,N_7563);
nand U8980 (N_8980,N_7415,N_7805);
nor U8981 (N_8981,N_7334,N_7282);
nor U8982 (N_8982,N_7472,N_7407);
and U8983 (N_8983,N_7269,N_7191);
nand U8984 (N_8984,N_7957,N_7196);
nor U8985 (N_8985,N_7603,N_7387);
nand U8986 (N_8986,N_7765,N_7764);
xor U8987 (N_8987,N_7911,N_7137);
nor U8988 (N_8988,N_7363,N_7826);
xnor U8989 (N_8989,N_7357,N_7137);
nor U8990 (N_8990,N_7993,N_7854);
nor U8991 (N_8991,N_7592,N_7710);
xnor U8992 (N_8992,N_7330,N_7392);
or U8993 (N_8993,N_7997,N_7722);
or U8994 (N_8994,N_7767,N_7889);
or U8995 (N_8995,N_7182,N_7614);
or U8996 (N_8996,N_7607,N_7234);
nor U8997 (N_8997,N_7110,N_7373);
and U8998 (N_8998,N_7061,N_7424);
xor U8999 (N_8999,N_7808,N_7397);
and U9000 (N_9000,N_8906,N_8557);
and U9001 (N_9001,N_8545,N_8326);
nand U9002 (N_9002,N_8372,N_8079);
xnor U9003 (N_9003,N_8967,N_8781);
xor U9004 (N_9004,N_8879,N_8133);
xor U9005 (N_9005,N_8756,N_8524);
xnor U9006 (N_9006,N_8089,N_8479);
or U9007 (N_9007,N_8918,N_8937);
or U9008 (N_9008,N_8722,N_8084);
nor U9009 (N_9009,N_8149,N_8527);
xnor U9010 (N_9010,N_8259,N_8220);
xor U9011 (N_9011,N_8564,N_8629);
nand U9012 (N_9012,N_8190,N_8349);
nand U9013 (N_9013,N_8275,N_8968);
xor U9014 (N_9014,N_8934,N_8995);
and U9015 (N_9015,N_8526,N_8869);
nor U9016 (N_9016,N_8344,N_8308);
nand U9017 (N_9017,N_8846,N_8263);
nand U9018 (N_9018,N_8321,N_8228);
nand U9019 (N_9019,N_8902,N_8192);
nor U9020 (N_9020,N_8795,N_8773);
xor U9021 (N_9021,N_8550,N_8333);
or U9022 (N_9022,N_8215,N_8491);
nor U9023 (N_9023,N_8176,N_8168);
or U9024 (N_9024,N_8733,N_8870);
nor U9025 (N_9025,N_8299,N_8067);
nand U9026 (N_9026,N_8681,N_8430);
nand U9027 (N_9027,N_8508,N_8963);
nand U9028 (N_9028,N_8005,N_8535);
and U9029 (N_9029,N_8347,N_8221);
nor U9030 (N_9030,N_8833,N_8266);
nand U9031 (N_9031,N_8831,N_8000);
and U9032 (N_9032,N_8602,N_8893);
or U9033 (N_9033,N_8548,N_8415);
and U9034 (N_9034,N_8287,N_8787);
nand U9035 (N_9035,N_8493,N_8664);
nand U9036 (N_9036,N_8859,N_8576);
nor U9037 (N_9037,N_8990,N_8691);
and U9038 (N_9038,N_8962,N_8026);
and U9039 (N_9039,N_8050,N_8844);
xnor U9040 (N_9040,N_8279,N_8481);
xnor U9041 (N_9041,N_8533,N_8357);
and U9042 (N_9042,N_8606,N_8480);
and U9043 (N_9043,N_8404,N_8815);
nand U9044 (N_9044,N_8579,N_8754);
nand U9045 (N_9045,N_8285,N_8753);
nand U9046 (N_9046,N_8863,N_8181);
nor U9047 (N_9047,N_8763,N_8459);
nand U9048 (N_9048,N_8405,N_8760);
nor U9049 (N_9049,N_8546,N_8441);
xnor U9050 (N_9050,N_8421,N_8179);
nor U9051 (N_9051,N_8074,N_8028);
and U9052 (N_9052,N_8029,N_8495);
and U9053 (N_9053,N_8223,N_8932);
nor U9054 (N_9054,N_8109,N_8626);
and U9055 (N_9055,N_8170,N_8646);
or U9056 (N_9056,N_8057,N_8975);
nand U9057 (N_9057,N_8928,N_8436);
or U9058 (N_9058,N_8832,N_8627);
nor U9059 (N_9059,N_8884,N_8850);
nor U9060 (N_9060,N_8238,N_8213);
nor U9061 (N_9061,N_8999,N_8796);
or U9062 (N_9062,N_8708,N_8729);
nor U9063 (N_9063,N_8858,N_8452);
xnor U9064 (N_9064,N_8689,N_8319);
nor U9065 (N_9065,N_8422,N_8538);
xor U9066 (N_9066,N_8668,N_8229);
nand U9067 (N_9067,N_8560,N_8396);
nand U9068 (N_9068,N_8631,N_8336);
and U9069 (N_9069,N_8061,N_8635);
xor U9070 (N_9070,N_8899,N_8866);
xor U9071 (N_9071,N_8577,N_8439);
or U9072 (N_9072,N_8597,N_8720);
nand U9073 (N_9073,N_8094,N_8182);
nor U9074 (N_9074,N_8009,N_8791);
xnor U9075 (N_9075,N_8512,N_8567);
or U9076 (N_9076,N_8040,N_8240);
nand U9077 (N_9077,N_8301,N_8409);
nor U9078 (N_9078,N_8103,N_8950);
or U9079 (N_9079,N_8854,N_8025);
and U9080 (N_9080,N_8158,N_8628);
and U9081 (N_9081,N_8408,N_8688);
nor U9082 (N_9082,N_8332,N_8751);
nand U9083 (N_9083,N_8713,N_8868);
or U9084 (N_9084,N_8939,N_8563);
or U9085 (N_9085,N_8261,N_8390);
and U9086 (N_9086,N_8216,N_8790);
and U9087 (N_9087,N_8883,N_8978);
nor U9088 (N_9088,N_8352,N_8701);
xor U9089 (N_9089,N_8402,N_8388);
nor U9090 (N_9090,N_8379,N_8852);
xor U9091 (N_9091,N_8268,N_8473);
or U9092 (N_9092,N_8666,N_8324);
and U9093 (N_9093,N_8356,N_8741);
nor U9094 (N_9094,N_8873,N_8813);
nand U9095 (N_9095,N_8260,N_8828);
nor U9096 (N_9096,N_8638,N_8195);
nand U9097 (N_9097,N_8391,N_8021);
nor U9098 (N_9098,N_8594,N_8281);
or U9099 (N_9099,N_8914,N_8426);
and U9100 (N_9100,N_8125,N_8736);
or U9101 (N_9101,N_8194,N_8609);
and U9102 (N_9102,N_8739,N_8387);
and U9103 (N_9103,N_8013,N_8983);
and U9104 (N_9104,N_8106,N_8130);
nor U9105 (N_9105,N_8203,N_8700);
or U9106 (N_9106,N_8414,N_8958);
and U9107 (N_9107,N_8429,N_8143);
nor U9108 (N_9108,N_8399,N_8212);
xnor U9109 (N_9109,N_8857,N_8834);
and U9110 (N_9110,N_8116,N_8816);
xnor U9111 (N_9111,N_8088,N_8601);
or U9112 (N_9112,N_8496,N_8384);
or U9113 (N_9113,N_8059,N_8822);
nor U9114 (N_9114,N_8237,N_8092);
nand U9115 (N_9115,N_8714,N_8592);
nor U9116 (N_9116,N_8742,N_8723);
nor U9117 (N_9117,N_8072,N_8960);
xor U9118 (N_9118,N_8471,N_8435);
nand U9119 (N_9119,N_8389,N_8082);
xor U9120 (N_9120,N_8146,N_8650);
and U9121 (N_9121,N_8175,N_8886);
and U9122 (N_9122,N_8519,N_8805);
nand U9123 (N_9123,N_8393,N_8329);
nor U9124 (N_9124,N_8710,N_8590);
nor U9125 (N_9125,N_8580,N_8537);
and U9126 (N_9126,N_8528,N_8362);
nor U9127 (N_9127,N_8572,N_8808);
xor U9128 (N_9128,N_8171,N_8864);
and U9129 (N_9129,N_8178,N_8358);
nand U9130 (N_9130,N_8929,N_8003);
nor U9131 (N_9131,N_8997,N_8861);
and U9132 (N_9132,N_8525,N_8293);
nand U9133 (N_9133,N_8947,N_8996);
nand U9134 (N_9134,N_8078,N_8989);
or U9135 (N_9135,N_8624,N_8660);
nand U9136 (N_9136,N_8992,N_8322);
xor U9137 (N_9137,N_8411,N_8164);
nand U9138 (N_9138,N_8151,N_8936);
and U9139 (N_9139,N_8539,N_8375);
or U9140 (N_9140,N_8341,N_8090);
and U9141 (N_9141,N_8209,N_8235);
nor U9142 (N_9142,N_8359,N_8063);
nand U9143 (N_9143,N_8381,N_8972);
nand U9144 (N_9144,N_8917,N_8447);
xor U9145 (N_9145,N_8271,N_8921);
xnor U9146 (N_9146,N_8172,N_8353);
xnor U9147 (N_9147,N_8476,N_8284);
xnor U9148 (N_9148,N_8490,N_8591);
xor U9149 (N_9149,N_8184,N_8054);
nor U9150 (N_9150,N_8488,N_8911);
nand U9151 (N_9151,N_8835,N_8186);
nor U9152 (N_9152,N_8219,N_8302);
or U9153 (N_9153,N_8913,N_8135);
xor U9154 (N_9154,N_8363,N_8424);
nand U9155 (N_9155,N_8743,N_8671);
nand U9156 (N_9156,N_8770,N_8113);
xnor U9157 (N_9157,N_8687,N_8839);
and U9158 (N_9158,N_8416,N_8001);
nand U9159 (N_9159,N_8543,N_8717);
or U9160 (N_9160,N_8649,N_8024);
or U9161 (N_9161,N_8725,N_8339);
and U9162 (N_9162,N_8872,N_8300);
xnor U9163 (N_9163,N_8956,N_8320);
nor U9164 (N_9164,N_8498,N_8916);
and U9165 (N_9165,N_8233,N_8019);
nand U9166 (N_9166,N_8286,N_8183);
nor U9167 (N_9167,N_8406,N_8305);
or U9168 (N_9168,N_8241,N_8290);
nand U9169 (N_9169,N_8676,N_8986);
and U9170 (N_9170,N_8607,N_8976);
nor U9171 (N_9171,N_8595,N_8484);
xnor U9172 (N_9172,N_8697,N_8020);
nor U9173 (N_9173,N_8193,N_8295);
xnor U9174 (N_9174,N_8291,N_8786);
and U9175 (N_9175,N_8737,N_8210);
and U9176 (N_9176,N_8513,N_8257);
and U9177 (N_9177,N_8058,N_8923);
xnor U9178 (N_9178,N_8758,N_8069);
or U9179 (N_9179,N_8250,N_8148);
xnor U9180 (N_9180,N_8407,N_8542);
and U9181 (N_9181,N_8675,N_8205);
and U9182 (N_9182,N_8798,N_8244);
or U9183 (N_9183,N_8503,N_8532);
nand U9184 (N_9184,N_8566,N_8711);
nand U9185 (N_9185,N_8905,N_8715);
nor U9186 (N_9186,N_8678,N_8772);
nand U9187 (N_9187,N_8880,N_8618);
and U9188 (N_9188,N_8112,N_8684);
nand U9189 (N_9189,N_8982,N_8892);
nand U9190 (N_9190,N_8392,N_8516);
nand U9191 (N_9191,N_8188,N_8517);
xor U9192 (N_9192,N_8239,N_8276);
nand U9193 (N_9193,N_8598,N_8120);
or U9194 (N_9194,N_8507,N_8129);
or U9195 (N_9195,N_8234,N_8100);
nand U9196 (N_9196,N_8251,N_8316);
or U9197 (N_9197,N_8677,N_8041);
nor U9198 (N_9198,N_8443,N_8199);
nand U9199 (N_9199,N_8957,N_8505);
xor U9200 (N_9200,N_8126,N_8052);
or U9201 (N_9201,N_8101,N_8900);
or U9202 (N_9202,N_8246,N_8462);
or U9203 (N_9203,N_8761,N_8823);
nor U9204 (N_9204,N_8115,N_8282);
nand U9205 (N_9205,N_8111,N_8325);
or U9206 (N_9206,N_8529,N_8465);
nand U9207 (N_9207,N_8682,N_8051);
and U9208 (N_9208,N_8804,N_8327);
nor U9209 (N_9209,N_8719,N_8413);
xor U9210 (N_9210,N_8780,N_8574);
and U9211 (N_9211,N_8838,N_8748);
and U9212 (N_9212,N_8136,N_8127);
and U9213 (N_9213,N_8800,N_8338);
nand U9214 (N_9214,N_8397,N_8346);
xnor U9215 (N_9215,N_8450,N_8487);
nand U9216 (N_9216,N_8478,N_8559);
xnor U9217 (N_9217,N_8885,N_8735);
nand U9218 (N_9218,N_8765,N_8530);
and U9219 (N_9219,N_8056,N_8915);
nor U9220 (N_9220,N_8045,N_8150);
nand U9221 (N_9221,N_8217,N_8904);
nand U9222 (N_9222,N_8940,N_8587);
and U9223 (N_9223,N_8208,N_8762);
nand U9224 (N_9224,N_8144,N_8355);
xnor U9225 (N_9225,N_8202,N_8027);
nor U9226 (N_9226,N_8908,N_8819);
or U9227 (N_9227,N_8901,N_8383);
nand U9228 (N_9228,N_8821,N_8410);
xor U9229 (N_9229,N_8177,N_8740);
and U9230 (N_9230,N_8075,N_8380);
or U9231 (N_9231,N_8836,N_8851);
and U9232 (N_9232,N_8504,N_8242);
and U9233 (N_9233,N_8097,N_8837);
nand U9234 (N_9234,N_8881,N_8412);
xor U9235 (N_9235,N_8469,N_8974);
and U9236 (N_9236,N_8553,N_8042);
or U9237 (N_9237,N_8665,N_8622);
or U9238 (N_9238,N_8738,N_8746);
nand U9239 (N_9239,N_8797,N_8068);
xnor U9240 (N_9240,N_8903,N_8673);
nor U9241 (N_9241,N_8312,N_8254);
and U9242 (N_9242,N_8777,N_8296);
nand U9243 (N_9243,N_8417,N_8946);
nor U9244 (N_9244,N_8653,N_8944);
nand U9245 (N_9245,N_8778,N_8511);
xnor U9246 (N_9246,N_8810,N_8267);
or U9247 (N_9247,N_8897,N_8514);
or U9248 (N_9248,N_8500,N_8599);
or U9249 (N_9249,N_8157,N_8095);
or U9250 (N_9250,N_8247,N_8255);
or U9251 (N_9251,N_8811,N_8752);
and U9252 (N_9252,N_8657,N_8334);
nand U9253 (N_9253,N_8925,N_8658);
nand U9254 (N_9254,N_8343,N_8948);
and U9255 (N_9255,N_8173,N_8464);
nand U9256 (N_9256,N_8812,N_8119);
nand U9257 (N_9257,N_8814,N_8702);
or U9258 (N_9258,N_8224,N_8354);
and U9259 (N_9259,N_8521,N_8612);
xor U9260 (N_9260,N_8776,N_8716);
and U9261 (N_9261,N_8924,N_8970);
and U9262 (N_9262,N_8933,N_8634);
and U9263 (N_9263,N_8782,N_8444);
and U9264 (N_9264,N_8841,N_8039);
nand U9265 (N_9265,N_8878,N_8428);
or U9266 (N_9266,N_8053,N_8656);
xnor U9267 (N_9267,N_8400,N_8034);
nand U9268 (N_9268,N_8745,N_8955);
xor U9269 (N_9269,N_8829,N_8032);
nand U9270 (N_9270,N_8033,N_8686);
and U9271 (N_9271,N_8562,N_8023);
nor U9272 (N_9272,N_8613,N_8558);
xnor U9273 (N_9273,N_8385,N_8573);
and U9274 (N_9274,N_8348,N_8467);
and U9275 (N_9275,N_8792,N_8693);
nand U9276 (N_9276,N_8919,N_8670);
nor U9277 (N_9277,N_8922,N_8337);
and U9278 (N_9278,N_8378,N_8840);
xnor U9279 (N_9279,N_8632,N_8454);
xor U9280 (N_9280,N_8672,N_8249);
xnor U9281 (N_9281,N_8941,N_8489);
nor U9282 (N_9282,N_8340,N_8964);
nand U9283 (N_9283,N_8342,N_8571);
xnor U9284 (N_9284,N_8637,N_8820);
nand U9285 (N_9285,N_8006,N_8108);
nor U9286 (N_9286,N_8098,N_8935);
and U9287 (N_9287,N_8310,N_8757);
nor U9288 (N_9288,N_8138,N_8707);
xor U9289 (N_9289,N_8582,N_8809);
or U9290 (N_9290,N_8002,N_8988);
and U9291 (N_9291,N_8207,N_8588);
nand U9292 (N_9292,N_8446,N_8010);
or U9293 (N_9293,N_8204,N_8482);
xor U9294 (N_9294,N_8584,N_8048);
xor U9295 (N_9295,N_8951,N_8440);
nand U9296 (N_9296,N_8272,N_8449);
nand U9297 (N_9297,N_8008,N_8501);
or U9298 (N_9298,N_8641,N_8642);
nand U9299 (N_9299,N_8142,N_8961);
nor U9300 (N_9300,N_8871,N_8062);
xor U9301 (N_9301,N_8137,N_8920);
or U9302 (N_9302,N_8486,N_8705);
nand U9303 (N_9303,N_8043,N_8382);
and U9304 (N_9304,N_8200,N_8386);
nor U9305 (N_9305,N_8140,N_8724);
nor U9306 (N_9306,N_8377,N_8226);
xnor U9307 (N_9307,N_8522,N_8153);
xor U9308 (N_9308,N_8926,N_8335);
nor U9309 (N_9309,N_8732,N_8654);
nand U9310 (N_9310,N_8853,N_8568);
nor U9311 (N_9311,N_8755,N_8110);
xnor U9312 (N_9312,N_8303,N_8784);
and U9313 (N_9313,N_8160,N_8206);
nand U9314 (N_9314,N_8015,N_8662);
nor U9315 (N_9315,N_8270,N_8827);
xnor U9316 (N_9316,N_8889,N_8448);
nand U9317 (N_9317,N_8734,N_8245);
nand U9318 (N_9318,N_8163,N_8064);
nand U9319 (N_9319,N_8096,N_8065);
and U9320 (N_9320,N_8749,N_8801);
nor U9321 (N_9321,N_8608,N_8842);
nand U9322 (N_9322,N_8086,N_8794);
nor U9323 (N_9323,N_8616,N_8456);
nand U9324 (N_9324,N_8395,N_8690);
nand U9325 (N_9325,N_8818,N_8669);
nand U9326 (N_9326,N_8458,N_8373);
xnor U9327 (N_9327,N_8189,N_8728);
xnor U9328 (N_9328,N_8523,N_8463);
xnor U9329 (N_9329,N_8973,N_8461);
nor U9330 (N_9330,N_8709,N_8766);
and U9331 (N_9331,N_8014,N_8091);
nor U9332 (N_9332,N_8102,N_8663);
xnor U9333 (N_9333,N_8625,N_8230);
and U9334 (N_9334,N_8896,N_8969);
nor U9335 (N_9335,N_8600,N_8018);
nor U9336 (N_9336,N_8977,N_8351);
and U9337 (N_9337,N_8419,N_8265);
or U9338 (N_9338,N_8132,N_8540);
or U9339 (N_9339,N_8161,N_8845);
and U9340 (N_9340,N_8848,N_8617);
xnor U9341 (N_9341,N_8159,N_8423);
xor U9342 (N_9342,N_8603,N_8038);
xnor U9343 (N_9343,N_8147,N_8288);
and U9344 (N_9344,N_8046,N_8965);
xor U9345 (N_9345,N_8593,N_8696);
and U9346 (N_9346,N_8769,N_8644);
nand U9347 (N_9347,N_8518,N_8248);
nor U9348 (N_9348,N_8274,N_8552);
xor U9349 (N_9349,N_8007,N_8698);
nor U9350 (N_9350,N_8912,N_8942);
nor U9351 (N_9351,N_8849,N_8694);
nor U9352 (N_9352,N_8554,N_8575);
nand U9353 (N_9353,N_8368,N_8227);
xnor U9354 (N_9354,N_8107,N_8953);
and U9355 (N_9355,N_8910,N_8768);
and U9356 (N_9356,N_8712,N_8981);
xor U9357 (N_9357,N_8497,N_8704);
and U9358 (N_9358,N_8830,N_8993);
nand U9359 (N_9359,N_8731,N_8509);
xnor U9360 (N_9360,N_8222,N_8536);
or U9361 (N_9361,N_8191,N_8807);
or U9362 (N_9362,N_8647,N_8099);
nor U9363 (N_9363,N_8474,N_8966);
or U9364 (N_9364,N_8451,N_8139);
and U9365 (N_9365,N_8987,N_8547);
or U9366 (N_9366,N_8747,N_8314);
nand U9367 (N_9367,N_8744,N_8198);
xnor U9368 (N_9368,N_8236,N_8971);
xor U9369 (N_9369,N_8699,N_8775);
xor U9370 (N_9370,N_8683,N_8876);
or U9371 (N_9371,N_8468,N_8639);
or U9372 (N_9372,N_8269,N_8252);
nor U9373 (N_9373,N_8292,N_8418);
and U9374 (N_9374,N_8589,N_8306);
and U9375 (N_9375,N_8817,N_8679);
nand U9376 (N_9376,N_8477,N_8196);
nand U9377 (N_9377,N_8201,N_8604);
nand U9378 (N_9378,N_8541,N_8515);
nand U9379 (N_9379,N_8145,N_8605);
nor U9380 (N_9380,N_8979,N_8350);
nand U9381 (N_9381,N_8167,N_8570);
xnor U9382 (N_9382,N_8783,N_8862);
nor U9383 (N_9383,N_8185,N_8485);
nor U9384 (N_9384,N_8596,N_8364);
and U9385 (N_9385,N_8824,N_8083);
or U9386 (N_9386,N_8044,N_8874);
or U9387 (N_9387,N_8492,N_8425);
and U9388 (N_9388,N_8569,N_8499);
and U9389 (N_9389,N_8398,N_8394);
xor U9390 (N_9390,N_8793,N_8531);
nand U9391 (N_9391,N_8453,N_8991);
xor U9392 (N_9392,N_8085,N_8544);
or U9393 (N_9393,N_8225,N_8551);
nand U9394 (N_9394,N_8856,N_8371);
xnor U9395 (N_9395,N_8174,N_8645);
nand U9396 (N_9396,N_8721,N_8894);
or U9397 (N_9397,N_8187,N_8855);
nand U9398 (N_9398,N_8556,N_8081);
nand U9399 (N_9399,N_8370,N_8843);
nand U9400 (N_9400,N_8785,N_8162);
and U9401 (N_9401,N_8433,N_8152);
or U9402 (N_9402,N_8131,N_8938);
xor U9403 (N_9403,N_8360,N_8802);
nand U9404 (N_9404,N_8648,N_8315);
xor U9405 (N_9405,N_8011,N_8374);
and U9406 (N_9406,N_8080,N_8318);
xor U9407 (N_9407,N_8016,N_8888);
and U9408 (N_9408,N_8294,N_8534);
xor U9409 (N_9409,N_8585,N_8431);
nor U9410 (N_9410,N_8949,N_8243);
nor U9411 (N_9411,N_8640,N_8278);
nand U9412 (N_9412,N_8231,N_8909);
or U9413 (N_9413,N_8442,N_8583);
and U9414 (N_9414,N_8718,N_8403);
nand U9415 (N_9415,N_8031,N_8586);
xnor U9416 (N_9416,N_8277,N_8520);
nand U9417 (N_9417,N_8945,N_8166);
or U9418 (N_9418,N_8847,N_8659);
or U9419 (N_9419,N_8105,N_8114);
xnor U9420 (N_9420,N_8361,N_8309);
and U9421 (N_9421,N_8890,N_8012);
nor U9422 (N_9422,N_8117,N_8214);
and U9423 (N_9423,N_8311,N_8943);
or U9424 (N_9424,N_8376,N_8460);
nand U9425 (N_9425,N_8651,N_8262);
or U9426 (N_9426,N_8549,N_8621);
and U9427 (N_9427,N_8211,N_8457);
nor U9428 (N_9428,N_8218,N_8614);
nor U9429 (N_9429,N_8022,N_8197);
xor U9430 (N_9430,N_8472,N_8774);
xnor U9431 (N_9431,N_8049,N_8652);
nor U9432 (N_9432,N_8954,N_8655);
or U9433 (N_9433,N_8298,N_8437);
and U9434 (N_9434,N_8661,N_8331);
or U9435 (N_9435,N_8674,N_8703);
and U9436 (N_9436,N_8093,N_8169);
and U9437 (N_9437,N_8581,N_8017);
and U9438 (N_9438,N_8985,N_8887);
nor U9439 (N_9439,N_8087,N_8667);
nor U9440 (N_9440,N_8789,N_8623);
nand U9441 (N_9441,N_8438,N_8891);
nand U9442 (N_9442,N_8055,N_8004);
nor U9443 (N_9443,N_8779,N_8998);
or U9444 (N_9444,N_8401,N_8898);
and U9445 (N_9445,N_8037,N_8258);
nor U9446 (N_9446,N_8070,N_8121);
xnor U9447 (N_9447,N_8060,N_8633);
nand U9448 (N_9448,N_8502,N_8264);
and U9449 (N_9449,N_8035,N_8141);
or U9450 (N_9450,N_8283,N_8727);
nor U9451 (N_9451,N_8692,N_8289);
or U9452 (N_9452,N_8071,N_8313);
nand U9453 (N_9453,N_8788,N_8565);
xor U9454 (N_9454,N_8952,N_8984);
nor U9455 (N_9455,N_8767,N_8959);
nand U9456 (N_9456,N_8877,N_8104);
or U9457 (N_9457,N_8273,N_8927);
nor U9458 (N_9458,N_8420,N_8445);
and U9459 (N_9459,N_8636,N_8895);
nor U9460 (N_9460,N_8317,N_8134);
nand U9461 (N_9461,N_8304,N_8280);
nor U9462 (N_9462,N_8455,N_8366);
or U9463 (N_9463,N_8860,N_8799);
nor U9464 (N_9464,N_8367,N_8330);
and U9465 (N_9465,N_8726,N_8470);
nand U9466 (N_9466,N_8345,N_8466);
nor U9467 (N_9467,N_8806,N_8610);
or U9468 (N_9468,N_8494,N_8759);
nand U9469 (N_9469,N_8907,N_8826);
and U9470 (N_9470,N_8695,N_8128);
nor U9471 (N_9471,N_8867,N_8369);
and U9472 (N_9472,N_8328,N_8124);
and U9473 (N_9473,N_8077,N_8232);
xnor U9474 (N_9474,N_8155,N_8685);
and U9475 (N_9475,N_8475,N_8620);
nor U9476 (N_9476,N_8076,N_8555);
nor U9477 (N_9477,N_8865,N_8323);
xnor U9478 (N_9478,N_8875,N_8561);
nor U9479 (N_9479,N_8882,N_8066);
xor U9480 (N_9480,N_8483,N_8771);
nor U9481 (N_9481,N_8156,N_8122);
nor U9482 (N_9482,N_8750,N_8803);
xor U9483 (N_9483,N_8427,N_8730);
xnor U9484 (N_9484,N_8510,N_8706);
nor U9485 (N_9485,N_8680,N_8036);
nor U9486 (N_9486,N_8073,N_8030);
xor U9487 (N_9487,N_8118,N_8154);
or U9488 (N_9488,N_8930,N_8578);
or U9489 (N_9489,N_8615,N_8256);
nand U9490 (N_9490,N_8506,N_8931);
nand U9491 (N_9491,N_8434,N_8165);
nand U9492 (N_9492,N_8365,N_8611);
xor U9493 (N_9493,N_8047,N_8994);
nor U9494 (N_9494,N_8253,N_8297);
and U9495 (N_9495,N_8630,N_8980);
or U9496 (N_9496,N_8825,N_8307);
and U9497 (N_9497,N_8432,N_8123);
nor U9498 (N_9498,N_8619,N_8764);
and U9499 (N_9499,N_8180,N_8643);
or U9500 (N_9500,N_8450,N_8077);
xor U9501 (N_9501,N_8287,N_8107);
or U9502 (N_9502,N_8788,N_8681);
or U9503 (N_9503,N_8160,N_8174);
or U9504 (N_9504,N_8700,N_8376);
nand U9505 (N_9505,N_8066,N_8037);
and U9506 (N_9506,N_8389,N_8036);
nand U9507 (N_9507,N_8592,N_8299);
or U9508 (N_9508,N_8966,N_8645);
nand U9509 (N_9509,N_8829,N_8101);
nand U9510 (N_9510,N_8977,N_8241);
or U9511 (N_9511,N_8568,N_8387);
and U9512 (N_9512,N_8138,N_8326);
nor U9513 (N_9513,N_8592,N_8530);
nor U9514 (N_9514,N_8117,N_8523);
and U9515 (N_9515,N_8647,N_8655);
xnor U9516 (N_9516,N_8165,N_8178);
and U9517 (N_9517,N_8921,N_8591);
nor U9518 (N_9518,N_8425,N_8393);
nand U9519 (N_9519,N_8912,N_8699);
and U9520 (N_9520,N_8292,N_8255);
nor U9521 (N_9521,N_8527,N_8055);
nor U9522 (N_9522,N_8222,N_8516);
nor U9523 (N_9523,N_8956,N_8594);
nor U9524 (N_9524,N_8114,N_8277);
and U9525 (N_9525,N_8907,N_8016);
xor U9526 (N_9526,N_8078,N_8064);
xnor U9527 (N_9527,N_8298,N_8694);
or U9528 (N_9528,N_8435,N_8182);
nor U9529 (N_9529,N_8686,N_8383);
or U9530 (N_9530,N_8922,N_8748);
or U9531 (N_9531,N_8815,N_8120);
nor U9532 (N_9532,N_8212,N_8525);
nor U9533 (N_9533,N_8158,N_8607);
nand U9534 (N_9534,N_8152,N_8111);
and U9535 (N_9535,N_8650,N_8469);
xor U9536 (N_9536,N_8311,N_8832);
nor U9537 (N_9537,N_8653,N_8869);
nor U9538 (N_9538,N_8836,N_8936);
nor U9539 (N_9539,N_8089,N_8887);
nand U9540 (N_9540,N_8983,N_8232);
nand U9541 (N_9541,N_8390,N_8975);
and U9542 (N_9542,N_8258,N_8507);
nand U9543 (N_9543,N_8562,N_8216);
and U9544 (N_9544,N_8708,N_8411);
nand U9545 (N_9545,N_8303,N_8380);
nand U9546 (N_9546,N_8145,N_8385);
or U9547 (N_9547,N_8154,N_8678);
nand U9548 (N_9548,N_8814,N_8053);
or U9549 (N_9549,N_8770,N_8539);
nand U9550 (N_9550,N_8997,N_8173);
nand U9551 (N_9551,N_8226,N_8350);
or U9552 (N_9552,N_8149,N_8676);
nand U9553 (N_9553,N_8363,N_8491);
xnor U9554 (N_9554,N_8249,N_8123);
nand U9555 (N_9555,N_8764,N_8202);
xnor U9556 (N_9556,N_8471,N_8433);
nor U9557 (N_9557,N_8083,N_8669);
nor U9558 (N_9558,N_8080,N_8835);
xnor U9559 (N_9559,N_8380,N_8774);
nor U9560 (N_9560,N_8455,N_8631);
xnor U9561 (N_9561,N_8909,N_8680);
nor U9562 (N_9562,N_8632,N_8302);
or U9563 (N_9563,N_8285,N_8929);
xnor U9564 (N_9564,N_8235,N_8584);
nand U9565 (N_9565,N_8380,N_8167);
and U9566 (N_9566,N_8823,N_8208);
and U9567 (N_9567,N_8348,N_8335);
xnor U9568 (N_9568,N_8484,N_8604);
xnor U9569 (N_9569,N_8019,N_8133);
or U9570 (N_9570,N_8469,N_8698);
and U9571 (N_9571,N_8135,N_8246);
nand U9572 (N_9572,N_8436,N_8656);
nor U9573 (N_9573,N_8097,N_8701);
xor U9574 (N_9574,N_8566,N_8347);
nor U9575 (N_9575,N_8826,N_8780);
xor U9576 (N_9576,N_8713,N_8179);
or U9577 (N_9577,N_8660,N_8431);
nor U9578 (N_9578,N_8743,N_8317);
xnor U9579 (N_9579,N_8364,N_8900);
and U9580 (N_9580,N_8817,N_8635);
or U9581 (N_9581,N_8726,N_8178);
nand U9582 (N_9582,N_8411,N_8470);
and U9583 (N_9583,N_8121,N_8456);
nor U9584 (N_9584,N_8921,N_8551);
or U9585 (N_9585,N_8032,N_8841);
nand U9586 (N_9586,N_8461,N_8189);
nor U9587 (N_9587,N_8313,N_8543);
xnor U9588 (N_9588,N_8455,N_8169);
xor U9589 (N_9589,N_8739,N_8176);
nor U9590 (N_9590,N_8937,N_8529);
nor U9591 (N_9591,N_8586,N_8977);
nor U9592 (N_9592,N_8591,N_8239);
and U9593 (N_9593,N_8753,N_8547);
nor U9594 (N_9594,N_8981,N_8413);
nand U9595 (N_9595,N_8622,N_8212);
and U9596 (N_9596,N_8545,N_8919);
nand U9597 (N_9597,N_8182,N_8904);
or U9598 (N_9598,N_8413,N_8203);
or U9599 (N_9599,N_8374,N_8324);
xor U9600 (N_9600,N_8626,N_8270);
xor U9601 (N_9601,N_8894,N_8052);
xnor U9602 (N_9602,N_8477,N_8854);
nor U9603 (N_9603,N_8248,N_8523);
xnor U9604 (N_9604,N_8857,N_8632);
xor U9605 (N_9605,N_8525,N_8843);
nor U9606 (N_9606,N_8268,N_8446);
and U9607 (N_9607,N_8044,N_8184);
nor U9608 (N_9608,N_8530,N_8930);
and U9609 (N_9609,N_8134,N_8900);
nor U9610 (N_9610,N_8048,N_8288);
nand U9611 (N_9611,N_8157,N_8638);
nand U9612 (N_9612,N_8107,N_8709);
or U9613 (N_9613,N_8211,N_8127);
or U9614 (N_9614,N_8576,N_8503);
xor U9615 (N_9615,N_8394,N_8382);
nand U9616 (N_9616,N_8686,N_8917);
nand U9617 (N_9617,N_8562,N_8898);
xor U9618 (N_9618,N_8850,N_8504);
or U9619 (N_9619,N_8467,N_8676);
and U9620 (N_9620,N_8241,N_8749);
nand U9621 (N_9621,N_8490,N_8279);
and U9622 (N_9622,N_8408,N_8111);
and U9623 (N_9623,N_8272,N_8223);
or U9624 (N_9624,N_8745,N_8050);
nor U9625 (N_9625,N_8104,N_8370);
nand U9626 (N_9626,N_8628,N_8274);
and U9627 (N_9627,N_8498,N_8559);
nand U9628 (N_9628,N_8067,N_8141);
nor U9629 (N_9629,N_8878,N_8163);
and U9630 (N_9630,N_8887,N_8880);
and U9631 (N_9631,N_8204,N_8916);
nand U9632 (N_9632,N_8740,N_8440);
nand U9633 (N_9633,N_8988,N_8150);
and U9634 (N_9634,N_8192,N_8960);
or U9635 (N_9635,N_8335,N_8188);
xnor U9636 (N_9636,N_8834,N_8221);
and U9637 (N_9637,N_8650,N_8030);
nand U9638 (N_9638,N_8154,N_8674);
and U9639 (N_9639,N_8568,N_8670);
nand U9640 (N_9640,N_8332,N_8297);
xor U9641 (N_9641,N_8482,N_8491);
xnor U9642 (N_9642,N_8085,N_8371);
and U9643 (N_9643,N_8852,N_8242);
and U9644 (N_9644,N_8013,N_8721);
or U9645 (N_9645,N_8623,N_8681);
nor U9646 (N_9646,N_8248,N_8839);
and U9647 (N_9647,N_8965,N_8161);
xor U9648 (N_9648,N_8848,N_8739);
nand U9649 (N_9649,N_8093,N_8693);
xnor U9650 (N_9650,N_8199,N_8787);
nand U9651 (N_9651,N_8287,N_8455);
xnor U9652 (N_9652,N_8079,N_8176);
or U9653 (N_9653,N_8738,N_8164);
or U9654 (N_9654,N_8010,N_8424);
and U9655 (N_9655,N_8746,N_8942);
or U9656 (N_9656,N_8951,N_8438);
nand U9657 (N_9657,N_8907,N_8468);
xor U9658 (N_9658,N_8803,N_8000);
xnor U9659 (N_9659,N_8438,N_8768);
and U9660 (N_9660,N_8974,N_8441);
and U9661 (N_9661,N_8626,N_8237);
nor U9662 (N_9662,N_8192,N_8304);
nor U9663 (N_9663,N_8228,N_8430);
nand U9664 (N_9664,N_8177,N_8066);
nor U9665 (N_9665,N_8846,N_8880);
nor U9666 (N_9666,N_8382,N_8317);
or U9667 (N_9667,N_8122,N_8292);
nor U9668 (N_9668,N_8596,N_8471);
nand U9669 (N_9669,N_8007,N_8104);
xnor U9670 (N_9670,N_8038,N_8537);
xor U9671 (N_9671,N_8518,N_8071);
and U9672 (N_9672,N_8676,N_8160);
and U9673 (N_9673,N_8818,N_8317);
or U9674 (N_9674,N_8483,N_8440);
or U9675 (N_9675,N_8006,N_8689);
nor U9676 (N_9676,N_8915,N_8946);
nand U9677 (N_9677,N_8875,N_8164);
nand U9678 (N_9678,N_8447,N_8191);
or U9679 (N_9679,N_8348,N_8203);
or U9680 (N_9680,N_8960,N_8184);
nand U9681 (N_9681,N_8509,N_8363);
xor U9682 (N_9682,N_8023,N_8419);
and U9683 (N_9683,N_8282,N_8645);
xnor U9684 (N_9684,N_8634,N_8656);
and U9685 (N_9685,N_8861,N_8334);
nor U9686 (N_9686,N_8751,N_8770);
nand U9687 (N_9687,N_8311,N_8087);
nand U9688 (N_9688,N_8133,N_8034);
xor U9689 (N_9689,N_8864,N_8860);
nand U9690 (N_9690,N_8420,N_8526);
or U9691 (N_9691,N_8169,N_8214);
nand U9692 (N_9692,N_8211,N_8881);
xnor U9693 (N_9693,N_8663,N_8579);
xor U9694 (N_9694,N_8910,N_8044);
nor U9695 (N_9695,N_8618,N_8935);
and U9696 (N_9696,N_8966,N_8125);
or U9697 (N_9697,N_8476,N_8556);
or U9698 (N_9698,N_8566,N_8863);
nor U9699 (N_9699,N_8145,N_8051);
or U9700 (N_9700,N_8491,N_8648);
or U9701 (N_9701,N_8189,N_8270);
xnor U9702 (N_9702,N_8896,N_8082);
nor U9703 (N_9703,N_8583,N_8902);
nand U9704 (N_9704,N_8037,N_8012);
or U9705 (N_9705,N_8658,N_8947);
xnor U9706 (N_9706,N_8238,N_8582);
xnor U9707 (N_9707,N_8099,N_8912);
or U9708 (N_9708,N_8165,N_8514);
and U9709 (N_9709,N_8988,N_8590);
and U9710 (N_9710,N_8238,N_8533);
and U9711 (N_9711,N_8055,N_8662);
or U9712 (N_9712,N_8748,N_8780);
xor U9713 (N_9713,N_8043,N_8645);
and U9714 (N_9714,N_8177,N_8052);
xor U9715 (N_9715,N_8432,N_8908);
and U9716 (N_9716,N_8962,N_8462);
and U9717 (N_9717,N_8221,N_8947);
or U9718 (N_9718,N_8365,N_8030);
or U9719 (N_9719,N_8393,N_8001);
and U9720 (N_9720,N_8651,N_8118);
and U9721 (N_9721,N_8619,N_8626);
nand U9722 (N_9722,N_8152,N_8141);
and U9723 (N_9723,N_8447,N_8500);
nor U9724 (N_9724,N_8040,N_8666);
nand U9725 (N_9725,N_8224,N_8333);
xor U9726 (N_9726,N_8352,N_8384);
or U9727 (N_9727,N_8787,N_8773);
xnor U9728 (N_9728,N_8745,N_8000);
xor U9729 (N_9729,N_8195,N_8122);
nand U9730 (N_9730,N_8580,N_8756);
and U9731 (N_9731,N_8974,N_8093);
nand U9732 (N_9732,N_8099,N_8708);
nor U9733 (N_9733,N_8478,N_8866);
nand U9734 (N_9734,N_8091,N_8312);
nand U9735 (N_9735,N_8523,N_8696);
nand U9736 (N_9736,N_8627,N_8642);
nor U9737 (N_9737,N_8224,N_8736);
xnor U9738 (N_9738,N_8132,N_8117);
nor U9739 (N_9739,N_8841,N_8083);
or U9740 (N_9740,N_8085,N_8770);
nand U9741 (N_9741,N_8689,N_8567);
nand U9742 (N_9742,N_8679,N_8523);
and U9743 (N_9743,N_8396,N_8956);
or U9744 (N_9744,N_8047,N_8170);
or U9745 (N_9745,N_8864,N_8975);
or U9746 (N_9746,N_8546,N_8636);
xor U9747 (N_9747,N_8943,N_8261);
nor U9748 (N_9748,N_8217,N_8012);
nand U9749 (N_9749,N_8901,N_8429);
and U9750 (N_9750,N_8364,N_8385);
xnor U9751 (N_9751,N_8581,N_8092);
xnor U9752 (N_9752,N_8648,N_8336);
and U9753 (N_9753,N_8866,N_8940);
xnor U9754 (N_9754,N_8413,N_8673);
xnor U9755 (N_9755,N_8284,N_8994);
nand U9756 (N_9756,N_8848,N_8025);
nand U9757 (N_9757,N_8468,N_8684);
xnor U9758 (N_9758,N_8612,N_8818);
nand U9759 (N_9759,N_8726,N_8882);
xor U9760 (N_9760,N_8211,N_8234);
or U9761 (N_9761,N_8080,N_8748);
nor U9762 (N_9762,N_8179,N_8587);
nand U9763 (N_9763,N_8865,N_8760);
nand U9764 (N_9764,N_8539,N_8031);
xnor U9765 (N_9765,N_8034,N_8317);
or U9766 (N_9766,N_8470,N_8637);
nand U9767 (N_9767,N_8469,N_8441);
and U9768 (N_9768,N_8594,N_8891);
and U9769 (N_9769,N_8112,N_8760);
xnor U9770 (N_9770,N_8606,N_8461);
or U9771 (N_9771,N_8124,N_8018);
xnor U9772 (N_9772,N_8313,N_8914);
or U9773 (N_9773,N_8913,N_8213);
nor U9774 (N_9774,N_8460,N_8986);
or U9775 (N_9775,N_8561,N_8973);
nand U9776 (N_9776,N_8670,N_8500);
nand U9777 (N_9777,N_8303,N_8542);
nand U9778 (N_9778,N_8685,N_8850);
nor U9779 (N_9779,N_8180,N_8219);
xnor U9780 (N_9780,N_8214,N_8710);
and U9781 (N_9781,N_8333,N_8626);
or U9782 (N_9782,N_8613,N_8639);
and U9783 (N_9783,N_8949,N_8933);
xor U9784 (N_9784,N_8189,N_8384);
or U9785 (N_9785,N_8438,N_8621);
xor U9786 (N_9786,N_8487,N_8972);
or U9787 (N_9787,N_8155,N_8514);
xnor U9788 (N_9788,N_8426,N_8193);
nand U9789 (N_9789,N_8048,N_8213);
nand U9790 (N_9790,N_8890,N_8928);
nor U9791 (N_9791,N_8840,N_8090);
xnor U9792 (N_9792,N_8838,N_8118);
and U9793 (N_9793,N_8250,N_8389);
xor U9794 (N_9794,N_8822,N_8931);
and U9795 (N_9795,N_8093,N_8995);
nand U9796 (N_9796,N_8905,N_8325);
or U9797 (N_9797,N_8291,N_8763);
and U9798 (N_9798,N_8397,N_8940);
and U9799 (N_9799,N_8619,N_8342);
xnor U9800 (N_9800,N_8012,N_8275);
and U9801 (N_9801,N_8357,N_8115);
nand U9802 (N_9802,N_8774,N_8835);
xnor U9803 (N_9803,N_8808,N_8669);
and U9804 (N_9804,N_8757,N_8358);
and U9805 (N_9805,N_8208,N_8400);
or U9806 (N_9806,N_8331,N_8888);
nand U9807 (N_9807,N_8207,N_8201);
xor U9808 (N_9808,N_8784,N_8597);
xor U9809 (N_9809,N_8666,N_8045);
xor U9810 (N_9810,N_8076,N_8545);
nand U9811 (N_9811,N_8648,N_8406);
nand U9812 (N_9812,N_8045,N_8272);
xor U9813 (N_9813,N_8984,N_8722);
or U9814 (N_9814,N_8039,N_8361);
xor U9815 (N_9815,N_8124,N_8633);
xnor U9816 (N_9816,N_8492,N_8136);
nand U9817 (N_9817,N_8062,N_8702);
nand U9818 (N_9818,N_8560,N_8412);
nand U9819 (N_9819,N_8763,N_8450);
or U9820 (N_9820,N_8357,N_8978);
or U9821 (N_9821,N_8387,N_8273);
and U9822 (N_9822,N_8676,N_8010);
and U9823 (N_9823,N_8739,N_8309);
or U9824 (N_9824,N_8678,N_8062);
xor U9825 (N_9825,N_8937,N_8679);
nand U9826 (N_9826,N_8743,N_8365);
and U9827 (N_9827,N_8028,N_8398);
nand U9828 (N_9828,N_8152,N_8320);
and U9829 (N_9829,N_8235,N_8954);
nand U9830 (N_9830,N_8802,N_8695);
xnor U9831 (N_9831,N_8618,N_8658);
xnor U9832 (N_9832,N_8845,N_8843);
xor U9833 (N_9833,N_8950,N_8051);
and U9834 (N_9834,N_8649,N_8186);
and U9835 (N_9835,N_8993,N_8644);
nand U9836 (N_9836,N_8746,N_8078);
or U9837 (N_9837,N_8961,N_8607);
nand U9838 (N_9838,N_8139,N_8400);
nor U9839 (N_9839,N_8968,N_8295);
and U9840 (N_9840,N_8852,N_8716);
xnor U9841 (N_9841,N_8423,N_8366);
xor U9842 (N_9842,N_8230,N_8696);
and U9843 (N_9843,N_8201,N_8435);
and U9844 (N_9844,N_8403,N_8460);
and U9845 (N_9845,N_8143,N_8318);
and U9846 (N_9846,N_8567,N_8591);
or U9847 (N_9847,N_8410,N_8208);
xor U9848 (N_9848,N_8609,N_8797);
or U9849 (N_9849,N_8281,N_8903);
xnor U9850 (N_9850,N_8527,N_8807);
or U9851 (N_9851,N_8973,N_8326);
or U9852 (N_9852,N_8357,N_8858);
nor U9853 (N_9853,N_8163,N_8017);
or U9854 (N_9854,N_8077,N_8458);
or U9855 (N_9855,N_8093,N_8502);
or U9856 (N_9856,N_8580,N_8827);
or U9857 (N_9857,N_8819,N_8740);
nor U9858 (N_9858,N_8724,N_8511);
and U9859 (N_9859,N_8952,N_8576);
xnor U9860 (N_9860,N_8333,N_8122);
and U9861 (N_9861,N_8809,N_8934);
xor U9862 (N_9862,N_8037,N_8845);
xnor U9863 (N_9863,N_8302,N_8845);
and U9864 (N_9864,N_8434,N_8914);
nor U9865 (N_9865,N_8810,N_8967);
nor U9866 (N_9866,N_8300,N_8434);
nor U9867 (N_9867,N_8824,N_8451);
or U9868 (N_9868,N_8562,N_8289);
or U9869 (N_9869,N_8559,N_8529);
nor U9870 (N_9870,N_8586,N_8840);
nor U9871 (N_9871,N_8059,N_8511);
nor U9872 (N_9872,N_8173,N_8565);
nor U9873 (N_9873,N_8853,N_8915);
nand U9874 (N_9874,N_8438,N_8967);
xor U9875 (N_9875,N_8960,N_8880);
xnor U9876 (N_9876,N_8190,N_8408);
and U9877 (N_9877,N_8781,N_8813);
xnor U9878 (N_9878,N_8920,N_8373);
and U9879 (N_9879,N_8919,N_8350);
or U9880 (N_9880,N_8113,N_8615);
or U9881 (N_9881,N_8157,N_8800);
or U9882 (N_9882,N_8795,N_8796);
xnor U9883 (N_9883,N_8372,N_8677);
nor U9884 (N_9884,N_8361,N_8322);
and U9885 (N_9885,N_8127,N_8561);
or U9886 (N_9886,N_8558,N_8837);
or U9887 (N_9887,N_8459,N_8603);
and U9888 (N_9888,N_8488,N_8594);
nor U9889 (N_9889,N_8289,N_8504);
nor U9890 (N_9890,N_8987,N_8068);
xor U9891 (N_9891,N_8148,N_8314);
xnor U9892 (N_9892,N_8785,N_8640);
nor U9893 (N_9893,N_8828,N_8637);
and U9894 (N_9894,N_8258,N_8347);
and U9895 (N_9895,N_8720,N_8050);
xnor U9896 (N_9896,N_8399,N_8208);
nor U9897 (N_9897,N_8825,N_8148);
nand U9898 (N_9898,N_8803,N_8188);
nor U9899 (N_9899,N_8160,N_8916);
and U9900 (N_9900,N_8369,N_8032);
nand U9901 (N_9901,N_8100,N_8072);
and U9902 (N_9902,N_8722,N_8576);
xor U9903 (N_9903,N_8977,N_8537);
or U9904 (N_9904,N_8074,N_8379);
or U9905 (N_9905,N_8535,N_8911);
nand U9906 (N_9906,N_8901,N_8154);
or U9907 (N_9907,N_8650,N_8141);
and U9908 (N_9908,N_8995,N_8475);
xnor U9909 (N_9909,N_8906,N_8585);
and U9910 (N_9910,N_8105,N_8090);
and U9911 (N_9911,N_8589,N_8186);
nor U9912 (N_9912,N_8967,N_8403);
nor U9913 (N_9913,N_8354,N_8130);
or U9914 (N_9914,N_8703,N_8389);
or U9915 (N_9915,N_8302,N_8204);
and U9916 (N_9916,N_8387,N_8964);
nand U9917 (N_9917,N_8578,N_8781);
and U9918 (N_9918,N_8188,N_8653);
or U9919 (N_9919,N_8544,N_8116);
xor U9920 (N_9920,N_8260,N_8800);
and U9921 (N_9921,N_8342,N_8296);
and U9922 (N_9922,N_8435,N_8322);
nor U9923 (N_9923,N_8248,N_8861);
nor U9924 (N_9924,N_8549,N_8229);
nor U9925 (N_9925,N_8637,N_8155);
nand U9926 (N_9926,N_8013,N_8729);
xnor U9927 (N_9927,N_8695,N_8707);
nand U9928 (N_9928,N_8794,N_8106);
and U9929 (N_9929,N_8989,N_8387);
or U9930 (N_9930,N_8562,N_8605);
xor U9931 (N_9931,N_8860,N_8494);
nor U9932 (N_9932,N_8669,N_8382);
xnor U9933 (N_9933,N_8492,N_8616);
xnor U9934 (N_9934,N_8578,N_8011);
xnor U9935 (N_9935,N_8439,N_8632);
or U9936 (N_9936,N_8612,N_8451);
or U9937 (N_9937,N_8854,N_8059);
nand U9938 (N_9938,N_8035,N_8583);
nor U9939 (N_9939,N_8551,N_8370);
or U9940 (N_9940,N_8364,N_8070);
and U9941 (N_9941,N_8420,N_8016);
and U9942 (N_9942,N_8806,N_8887);
or U9943 (N_9943,N_8685,N_8063);
and U9944 (N_9944,N_8651,N_8443);
nor U9945 (N_9945,N_8163,N_8309);
nor U9946 (N_9946,N_8102,N_8431);
nand U9947 (N_9947,N_8700,N_8244);
nand U9948 (N_9948,N_8055,N_8490);
and U9949 (N_9949,N_8625,N_8877);
nor U9950 (N_9950,N_8327,N_8380);
and U9951 (N_9951,N_8416,N_8988);
and U9952 (N_9952,N_8750,N_8522);
xnor U9953 (N_9953,N_8890,N_8055);
nor U9954 (N_9954,N_8512,N_8334);
and U9955 (N_9955,N_8096,N_8572);
xor U9956 (N_9956,N_8586,N_8198);
and U9957 (N_9957,N_8782,N_8479);
and U9958 (N_9958,N_8393,N_8867);
or U9959 (N_9959,N_8174,N_8997);
nor U9960 (N_9960,N_8052,N_8547);
or U9961 (N_9961,N_8042,N_8926);
or U9962 (N_9962,N_8087,N_8419);
nor U9963 (N_9963,N_8543,N_8891);
nand U9964 (N_9964,N_8069,N_8435);
xnor U9965 (N_9965,N_8114,N_8990);
and U9966 (N_9966,N_8189,N_8812);
nand U9967 (N_9967,N_8005,N_8304);
and U9968 (N_9968,N_8837,N_8957);
and U9969 (N_9969,N_8544,N_8806);
xor U9970 (N_9970,N_8299,N_8725);
or U9971 (N_9971,N_8558,N_8595);
xor U9972 (N_9972,N_8907,N_8236);
nor U9973 (N_9973,N_8742,N_8627);
xnor U9974 (N_9974,N_8965,N_8381);
or U9975 (N_9975,N_8695,N_8948);
xor U9976 (N_9976,N_8818,N_8203);
nand U9977 (N_9977,N_8175,N_8074);
nor U9978 (N_9978,N_8780,N_8151);
and U9979 (N_9979,N_8993,N_8252);
nor U9980 (N_9980,N_8193,N_8896);
xnor U9981 (N_9981,N_8271,N_8953);
nor U9982 (N_9982,N_8945,N_8025);
xor U9983 (N_9983,N_8673,N_8607);
xnor U9984 (N_9984,N_8891,N_8537);
and U9985 (N_9985,N_8368,N_8685);
and U9986 (N_9986,N_8971,N_8201);
and U9987 (N_9987,N_8313,N_8537);
nor U9988 (N_9988,N_8586,N_8614);
nor U9989 (N_9989,N_8641,N_8024);
nand U9990 (N_9990,N_8778,N_8008);
or U9991 (N_9991,N_8721,N_8273);
or U9992 (N_9992,N_8405,N_8732);
or U9993 (N_9993,N_8438,N_8962);
nor U9994 (N_9994,N_8216,N_8259);
and U9995 (N_9995,N_8756,N_8983);
xor U9996 (N_9996,N_8351,N_8076);
or U9997 (N_9997,N_8534,N_8779);
nor U9998 (N_9998,N_8410,N_8614);
nand U9999 (N_9999,N_8402,N_8701);
nand U10000 (N_10000,N_9231,N_9165);
and U10001 (N_10001,N_9463,N_9601);
and U10002 (N_10002,N_9209,N_9711);
nor U10003 (N_10003,N_9872,N_9675);
nor U10004 (N_10004,N_9943,N_9327);
or U10005 (N_10005,N_9791,N_9220);
xnor U10006 (N_10006,N_9348,N_9861);
nand U10007 (N_10007,N_9580,N_9741);
and U10008 (N_10008,N_9211,N_9565);
or U10009 (N_10009,N_9730,N_9097);
nand U10010 (N_10010,N_9830,N_9841);
xnor U10011 (N_10011,N_9022,N_9620);
nand U10012 (N_10012,N_9556,N_9956);
or U10013 (N_10013,N_9278,N_9721);
nor U10014 (N_10014,N_9996,N_9469);
nor U10015 (N_10015,N_9948,N_9389);
and U10016 (N_10016,N_9437,N_9552);
xnor U10017 (N_10017,N_9779,N_9099);
and U10018 (N_10018,N_9120,N_9588);
nor U10019 (N_10019,N_9558,N_9973);
nand U10020 (N_10020,N_9893,N_9275);
or U10021 (N_10021,N_9140,N_9570);
nand U10022 (N_10022,N_9160,N_9645);
nand U10023 (N_10023,N_9563,N_9542);
nand U10024 (N_10024,N_9850,N_9131);
or U10025 (N_10025,N_9153,N_9033);
nor U10026 (N_10026,N_9255,N_9221);
nand U10027 (N_10027,N_9486,N_9246);
nand U10028 (N_10028,N_9868,N_9093);
nand U10029 (N_10029,N_9988,N_9931);
nand U10030 (N_10030,N_9627,N_9240);
or U10031 (N_10031,N_9590,N_9933);
nand U10032 (N_10032,N_9470,N_9137);
nand U10033 (N_10033,N_9768,N_9608);
nor U10034 (N_10034,N_9986,N_9226);
nor U10035 (N_10035,N_9669,N_9346);
nand U10036 (N_10036,N_9502,N_9499);
or U10037 (N_10037,N_9998,N_9707);
nor U10038 (N_10038,N_9501,N_9071);
and U10039 (N_10039,N_9800,N_9091);
and U10040 (N_10040,N_9802,N_9966);
nand U10041 (N_10041,N_9717,N_9674);
nand U10042 (N_10042,N_9441,N_9037);
and U10043 (N_10043,N_9155,N_9633);
and U10044 (N_10044,N_9458,N_9798);
xnor U10045 (N_10045,N_9826,N_9701);
and U10046 (N_10046,N_9029,N_9911);
xor U10047 (N_10047,N_9460,N_9951);
xnor U10048 (N_10048,N_9134,N_9766);
and U10049 (N_10049,N_9832,N_9349);
or U10050 (N_10050,N_9239,N_9846);
or U10051 (N_10051,N_9115,N_9173);
nor U10052 (N_10052,N_9159,N_9735);
nand U10053 (N_10053,N_9359,N_9817);
xor U10054 (N_10054,N_9629,N_9733);
or U10055 (N_10055,N_9808,N_9923);
nand U10056 (N_10056,N_9096,N_9285);
nor U10057 (N_10057,N_9320,N_9411);
nand U10058 (N_10058,N_9292,N_9658);
or U10059 (N_10059,N_9856,N_9196);
nor U10060 (N_10060,N_9541,N_9536);
or U10061 (N_10061,N_9754,N_9982);
xor U10062 (N_10062,N_9922,N_9328);
nor U10063 (N_10063,N_9677,N_9077);
or U10064 (N_10064,N_9506,N_9495);
nor U10065 (N_10065,N_9012,N_9807);
xnor U10066 (N_10066,N_9452,N_9414);
and U10067 (N_10067,N_9987,N_9827);
and U10068 (N_10068,N_9522,N_9859);
or U10069 (N_10069,N_9824,N_9573);
or U10070 (N_10070,N_9525,N_9079);
or U10071 (N_10071,N_9537,N_9916);
or U10072 (N_10072,N_9459,N_9069);
and U10073 (N_10073,N_9617,N_9036);
or U10074 (N_10074,N_9533,N_9270);
xnor U10075 (N_10075,N_9141,N_9614);
xnor U10076 (N_10076,N_9528,N_9952);
nand U10077 (N_10077,N_9129,N_9642);
and U10078 (N_10078,N_9118,N_9582);
and U10079 (N_10079,N_9942,N_9600);
or U10080 (N_10080,N_9594,N_9494);
nor U10081 (N_10081,N_9993,N_9087);
or U10082 (N_10082,N_9177,N_9475);
nor U10083 (N_10083,N_9027,N_9377);
xnor U10084 (N_10084,N_9028,N_9063);
nor U10085 (N_10085,N_9716,N_9001);
nor U10086 (N_10086,N_9619,N_9967);
and U10087 (N_10087,N_9186,N_9341);
and U10088 (N_10088,N_9289,N_9198);
nand U10089 (N_10089,N_9078,N_9488);
xnor U10090 (N_10090,N_9946,N_9656);
nand U10091 (N_10091,N_9446,N_9521);
or U10092 (N_10092,N_9920,N_9040);
and U10093 (N_10093,N_9185,N_9139);
nand U10094 (N_10094,N_9516,N_9954);
nand U10095 (N_10095,N_9421,N_9055);
nor U10096 (N_10096,N_9630,N_9272);
and U10097 (N_10097,N_9984,N_9737);
and U10098 (N_10098,N_9613,N_9422);
and U10099 (N_10099,N_9337,N_9105);
or U10100 (N_10100,N_9511,N_9358);
nand U10101 (N_10101,N_9074,N_9941);
or U10102 (N_10102,N_9972,N_9370);
or U10103 (N_10103,N_9783,N_9944);
or U10104 (N_10104,N_9535,N_9273);
or U10105 (N_10105,N_9583,N_9775);
nor U10106 (N_10106,N_9811,N_9968);
nand U10107 (N_10107,N_9336,N_9867);
or U10108 (N_10108,N_9918,N_9661);
xnor U10109 (N_10109,N_9625,N_9064);
xnor U10110 (N_10110,N_9207,N_9695);
xor U10111 (N_10111,N_9568,N_9975);
and U10112 (N_10112,N_9035,N_9863);
and U10113 (N_10113,N_9950,N_9052);
nor U10114 (N_10114,N_9876,N_9329);
nand U10115 (N_10115,N_9393,N_9156);
and U10116 (N_10116,N_9317,N_9248);
and U10117 (N_10117,N_9326,N_9215);
xor U10118 (N_10118,N_9058,N_9383);
nand U10119 (N_10119,N_9472,N_9080);
and U10120 (N_10120,N_9233,N_9151);
xor U10121 (N_10121,N_9133,N_9218);
and U10122 (N_10122,N_9615,N_9531);
xor U10123 (N_10123,N_9126,N_9917);
xor U10124 (N_10124,N_9686,N_9760);
or U10125 (N_10125,N_9764,N_9960);
nor U10126 (N_10126,N_9852,N_9610);
xor U10127 (N_10127,N_9823,N_9748);
and U10128 (N_10128,N_9799,N_9417);
nand U10129 (N_10129,N_9219,N_9050);
xor U10130 (N_10130,N_9713,N_9148);
and U10131 (N_10131,N_9908,N_9031);
or U10132 (N_10132,N_9130,N_9801);
or U10133 (N_10133,N_9976,N_9006);
and U10134 (N_10134,N_9632,N_9862);
nor U10135 (N_10135,N_9789,N_9443);
xnor U10136 (N_10136,N_9263,N_9702);
or U10137 (N_10137,N_9929,N_9427);
or U10138 (N_10138,N_9985,N_9260);
nor U10139 (N_10139,N_9434,N_9896);
or U10140 (N_10140,N_9670,N_9279);
nor U10141 (N_10141,N_9119,N_9201);
or U10142 (N_10142,N_9371,N_9979);
and U10143 (N_10143,N_9212,N_9243);
or U10144 (N_10144,N_9671,N_9401);
xor U10145 (N_10145,N_9145,N_9445);
nor U10146 (N_10146,N_9631,N_9318);
nand U10147 (N_10147,N_9300,N_9236);
nor U10148 (N_10148,N_9049,N_9869);
xor U10149 (N_10149,N_9550,N_9390);
xnor U10150 (N_10150,N_9338,N_9901);
nor U10151 (N_10151,N_9136,N_9291);
and U10152 (N_10152,N_9990,N_9855);
xnor U10153 (N_10153,N_9188,N_9785);
and U10154 (N_10154,N_9725,N_9394);
nand U10155 (N_10155,N_9657,N_9110);
and U10156 (N_10156,N_9415,N_9296);
nor U10157 (N_10157,N_9666,N_9111);
nor U10158 (N_10158,N_9277,N_9391);
or U10159 (N_10159,N_9977,N_9722);
nor U10160 (N_10160,N_9324,N_9771);
xor U10161 (N_10161,N_9780,N_9652);
or U10162 (N_10162,N_9054,N_9308);
and U10163 (N_10163,N_9724,N_9367);
or U10164 (N_10164,N_9903,N_9879);
nand U10165 (N_10165,N_9485,N_9549);
xor U10166 (N_10166,N_9510,N_9624);
nand U10167 (N_10167,N_9758,N_9962);
or U10168 (N_10168,N_9424,N_9727);
or U10169 (N_10169,N_9554,N_9909);
nand U10170 (N_10170,N_9067,N_9526);
nor U10171 (N_10171,N_9072,N_9483);
or U10172 (N_10172,N_9213,N_9761);
and U10173 (N_10173,N_9509,N_9587);
nand U10174 (N_10174,N_9907,N_9312);
xnor U10175 (N_10175,N_9524,N_9860);
nand U10176 (N_10176,N_9679,N_9847);
xor U10177 (N_10177,N_9163,N_9203);
and U10178 (N_10178,N_9643,N_9958);
xnor U10179 (N_10179,N_9599,N_9870);
or U10180 (N_10180,N_9267,N_9407);
nor U10181 (N_10181,N_9913,N_9271);
and U10182 (N_10182,N_9309,N_9405);
nand U10183 (N_10183,N_9892,N_9109);
nand U10184 (N_10184,N_9503,N_9481);
nor U10185 (N_10185,N_9408,N_9915);
xor U10186 (N_10186,N_9476,N_9994);
nand U10187 (N_10187,N_9835,N_9332);
nor U10188 (N_10188,N_9623,N_9086);
and U10189 (N_10189,N_9728,N_9172);
nor U10190 (N_10190,N_9880,N_9821);
nor U10191 (N_10191,N_9238,N_9423);
nor U10192 (N_10192,N_9101,N_9127);
xor U10193 (N_10193,N_9124,N_9607);
xor U10194 (N_10194,N_9303,N_9874);
xor U10195 (N_10195,N_9032,N_9831);
or U10196 (N_10196,N_9106,N_9366);
nand U10197 (N_10197,N_9970,N_9833);
or U10198 (N_10198,N_9378,N_9057);
nand U10199 (N_10199,N_9457,N_9123);
and U10200 (N_10200,N_9878,N_9368);
xnor U10201 (N_10201,N_9492,N_9882);
or U10202 (N_10202,N_9487,N_9819);
and U10203 (N_10203,N_9769,N_9314);
xnor U10204 (N_10204,N_9809,N_9989);
and U10205 (N_10205,N_9949,N_9953);
xnor U10206 (N_10206,N_9822,N_9283);
or U10207 (N_10207,N_9757,N_9429);
nor U10208 (N_10208,N_9781,N_9232);
xor U10209 (N_10209,N_9011,N_9969);
or U10210 (N_10210,N_9190,N_9685);
or U10211 (N_10211,N_9168,N_9744);
xnor U10212 (N_10212,N_9567,N_9584);
nor U10213 (N_10213,N_9256,N_9090);
or U10214 (N_10214,N_9113,N_9650);
and U10215 (N_10215,N_9355,N_9293);
nand U10216 (N_10216,N_9065,N_9450);
nor U10217 (N_10217,N_9651,N_9927);
and U10218 (N_10218,N_9644,N_9191);
or U10219 (N_10219,N_9222,N_9813);
xor U10220 (N_10220,N_9382,N_9726);
and U10221 (N_10221,N_9618,N_9400);
nand U10222 (N_10222,N_9247,N_9265);
nand U10223 (N_10223,N_9540,N_9574);
and U10224 (N_10224,N_9208,N_9519);
xnor U10225 (N_10225,N_9223,N_9350);
and U10226 (N_10226,N_9885,N_9478);
nand U10227 (N_10227,N_9959,N_9444);
nor U10228 (N_10228,N_9076,N_9796);
nor U10229 (N_10229,N_9805,N_9353);
xor U10230 (N_10230,N_9845,N_9362);
or U10231 (N_10231,N_9147,N_9621);
and U10232 (N_10232,N_9965,N_9397);
xor U10233 (N_10233,N_9639,N_9773);
nor U10234 (N_10234,N_9017,N_9683);
xor U10235 (N_10235,N_9392,N_9398);
nor U10236 (N_10236,N_9128,N_9871);
nand U10237 (N_10237,N_9008,N_9112);
nand U10238 (N_10238,N_9684,N_9297);
xnor U10239 (N_10239,N_9810,N_9333);
and U10240 (N_10240,N_9655,N_9244);
nand U10241 (N_10241,N_9047,N_9640);
nor U10242 (N_10242,N_9399,N_9453);
and U10243 (N_10243,N_9396,N_9828);
xor U10244 (N_10244,N_9844,N_9842);
nand U10245 (N_10245,N_9419,N_9418);
xnor U10246 (N_10246,N_9305,N_9138);
xnor U10247 (N_10247,N_9622,N_9498);
nand U10248 (N_10248,N_9276,N_9490);
or U10249 (N_10249,N_9566,N_9334);
or U10250 (N_10250,N_9720,N_9787);
or U10251 (N_10251,N_9774,N_9262);
nand U10252 (N_10252,N_9234,N_9938);
xnor U10253 (N_10253,N_9466,N_9983);
or U10254 (N_10254,N_9663,N_9039);
and U10255 (N_10255,N_9455,N_9322);
or U10256 (N_10256,N_9376,N_9557);
xnor U10257 (N_10257,N_9548,N_9816);
xor U10258 (N_10258,N_9019,N_9315);
xor U10259 (N_10259,N_9932,N_9125);
or U10260 (N_10260,N_9936,N_9529);
nor U10261 (N_10261,N_9009,N_9974);
and U10262 (N_10262,N_9659,N_9225);
xnor U10263 (N_10263,N_9897,N_9092);
nor U10264 (N_10264,N_9611,N_9117);
nand U10265 (N_10265,N_9088,N_9505);
nor U10266 (N_10266,N_9339,N_9189);
nand U10267 (N_10267,N_9082,N_9387);
nor U10268 (N_10268,N_9288,N_9759);
and U10269 (N_10269,N_9280,N_9202);
and U10270 (N_10270,N_9905,N_9045);
nor U10271 (N_10271,N_9325,N_9762);
xnor U10272 (N_10272,N_9053,N_9770);
nand U10273 (N_10273,N_9712,N_9602);
nor U10274 (N_10274,N_9646,N_9157);
nand U10275 (N_10275,N_9734,N_9507);
nand U10276 (N_10276,N_9562,N_9520);
or U10277 (N_10277,N_9016,N_9500);
nor U10278 (N_10278,N_9647,N_9559);
nor U10279 (N_10279,N_9921,N_9089);
nand U10280 (N_10280,N_9797,N_9152);
nand U10281 (N_10281,N_9372,N_9214);
nor U10282 (N_10282,N_9638,N_9068);
and U10283 (N_10283,N_9132,N_9585);
nand U10284 (N_10284,N_9102,N_9820);
nor U10285 (N_10285,N_9178,N_9061);
and U10286 (N_10286,N_9753,N_9561);
xnor U10287 (N_10287,N_9302,N_9484);
nor U10288 (N_10288,N_9204,N_9739);
and U10289 (N_10289,N_9708,N_9402);
nor U10290 (N_10290,N_9480,N_9806);
nor U10291 (N_10291,N_9474,N_9569);
nand U10292 (N_10292,N_9637,N_9409);
xor U10293 (N_10293,N_9307,N_9981);
and U10294 (N_10294,N_9149,N_9678);
nand U10295 (N_10295,N_9731,N_9628);
xor U10296 (N_10296,N_9073,N_9013);
nand U10297 (N_10297,N_9504,N_9877);
nor U10298 (N_10298,N_9210,N_9553);
xor U10299 (N_10299,N_9883,N_9041);
nand U10300 (N_10300,N_9875,N_9829);
nand U10301 (N_10301,N_9146,N_9375);
xnor U10302 (N_10302,N_9200,N_9971);
and U10303 (N_10303,N_9335,N_9992);
or U10304 (N_10304,N_9205,N_9812);
and U10305 (N_10305,N_9606,N_9926);
nand U10306 (N_10306,N_9616,N_9059);
xor U10307 (N_10307,N_9281,N_9538);
nand U10308 (N_10308,N_9866,N_9752);
or U10309 (N_10309,N_9945,N_9085);
nor U10310 (N_10310,N_9530,N_9170);
nand U10311 (N_10311,N_9732,N_9264);
or U10312 (N_10312,N_9319,N_9254);
and U10313 (N_10313,N_9782,N_9161);
nor U10314 (N_10314,N_9104,N_9961);
and U10315 (N_10315,N_9749,N_9406);
nand U10316 (N_10316,N_9473,N_9286);
and U10317 (N_10317,N_9442,N_9311);
or U10318 (N_10318,N_9192,N_9171);
and U10319 (N_10319,N_9023,N_9680);
nand U10320 (N_10320,N_9287,N_9162);
xnor U10321 (N_10321,N_9605,N_9784);
xnor U10322 (N_10322,N_9298,N_9894);
nor U10323 (N_10323,N_9321,N_9589);
nor U10324 (N_10324,N_9745,N_9747);
nor U10325 (N_10325,N_9245,N_9274);
or U10326 (N_10326,N_9268,N_9294);
nor U10327 (N_10327,N_9898,N_9895);
and U10328 (N_10328,N_9636,N_9653);
or U10329 (N_10329,N_9572,N_9266);
nor U10330 (N_10330,N_9062,N_9269);
nor U10331 (N_10331,N_9430,N_9435);
or U10332 (N_10332,N_9888,N_9681);
and U10333 (N_10333,N_9544,N_9925);
nor U10334 (N_10334,N_9697,N_9718);
xor U10335 (N_10335,N_9934,N_9886);
nor U10336 (N_10336,N_9345,N_9000);
or U10337 (N_10337,N_9532,N_9482);
nand U10338 (N_10338,N_9451,N_9386);
and U10339 (N_10339,N_9108,N_9043);
xnor U10340 (N_10340,N_9517,N_9818);
xor U10341 (N_10341,N_9719,N_9042);
nor U10342 (N_10342,N_9682,N_9425);
nand U10343 (N_10343,N_9788,N_9051);
xor U10344 (N_10344,N_9169,N_9249);
xor U10345 (N_10345,N_9676,N_9586);
nand U10346 (N_10346,N_9858,N_9227);
xnor U10347 (N_10347,N_9837,N_9471);
or U10348 (N_10348,N_9374,N_9710);
xnor U10349 (N_10349,N_9497,N_9313);
xnor U10350 (N_10350,N_9662,N_9352);
xor U10351 (N_10351,N_9380,N_9224);
xnor U10352 (N_10352,N_9513,N_9534);
nand U10353 (N_10353,N_9340,N_9344);
nor U10354 (N_10354,N_9593,N_9014);
or U10355 (N_10355,N_9122,N_9449);
and U10356 (N_10356,N_9765,N_9696);
or U10357 (N_10357,N_9384,N_9030);
or U10358 (N_10358,N_9007,N_9515);
nor U10359 (N_10359,N_9714,N_9603);
xor U10360 (N_10360,N_9660,N_9216);
nor U10361 (N_10361,N_9991,N_9121);
xnor U10362 (N_10362,N_9667,N_9709);
nand U10363 (N_10363,N_9595,N_9767);
or U10364 (N_10364,N_9456,N_9034);
xnor U10365 (N_10365,N_9413,N_9436);
and U10366 (N_10366,N_9103,N_9295);
xor U10367 (N_10367,N_9715,N_9323);
and U10368 (N_10368,N_9523,N_9705);
nor U10369 (N_10369,N_9464,N_9454);
or U10370 (N_10370,N_9884,N_9664);
nand U10371 (N_10371,N_9465,N_9546);
nand U10372 (N_10372,N_9839,N_9447);
nor U10373 (N_10373,N_9448,N_9729);
and U10374 (N_10374,N_9235,N_9919);
nor U10375 (N_10375,N_9902,N_9906);
nand U10376 (N_10376,N_9412,N_9410);
nand U10377 (N_10377,N_9539,N_9508);
xnor U10378 (N_10378,N_9564,N_9075);
nand U10379 (N_10379,N_9814,N_9304);
nand U10380 (N_10380,N_9364,N_9776);
and U10381 (N_10381,N_9889,N_9512);
xor U10382 (N_10382,N_9259,N_9258);
xor U10383 (N_10383,N_9598,N_9840);
xnor U10384 (N_10384,N_9107,N_9865);
xor U10385 (N_10385,N_9066,N_9158);
or U10386 (N_10386,N_9021,N_9577);
xnor U10387 (N_10387,N_9851,N_9357);
and U10388 (N_10388,N_9803,N_9070);
nand U10389 (N_10389,N_9467,N_9310);
xnor U10390 (N_10390,N_9648,N_9166);
nand U10391 (N_10391,N_9015,N_9164);
nor U10392 (N_10392,N_9834,N_9230);
nand U10393 (N_10393,N_9228,N_9306);
and U10394 (N_10394,N_9612,N_9257);
and U10395 (N_10395,N_9193,N_9786);
nand U10396 (N_10396,N_9426,N_9253);
xnor U10397 (N_10397,N_9825,N_9928);
nor U10398 (N_10398,N_9356,N_9003);
and U10399 (N_10399,N_9330,N_9116);
and U10400 (N_10400,N_9957,N_9004);
or U10401 (N_10401,N_9252,N_9751);
xnor U10402 (N_10402,N_9777,N_9997);
nor U10403 (N_10403,N_9217,N_9755);
nand U10404 (N_10404,N_9299,N_9388);
nor U10405 (N_10405,N_9242,N_9020);
nand U10406 (N_10406,N_9848,N_9738);
or U10407 (N_10407,N_9044,N_9609);
or U10408 (N_10408,N_9365,N_9995);
and U10409 (N_10409,N_9687,N_9343);
or U10410 (N_10410,N_9914,N_9518);
and U10411 (N_10411,N_9439,N_9433);
nand U10412 (N_10412,N_9964,N_9947);
nor U10413 (N_10413,N_9493,N_9694);
nand U10414 (N_10414,N_9836,N_9545);
nor U10415 (N_10415,N_9527,N_9404);
nand U10416 (N_10416,N_9025,N_9688);
nor U10417 (N_10417,N_9024,N_9369);
nor U10418 (N_10418,N_9199,N_9854);
nand U10419 (N_10419,N_9010,N_9381);
or U10420 (N_10420,N_9700,N_9468);
xnor U10421 (N_10421,N_9999,N_9591);
nor U10422 (N_10422,N_9154,N_9963);
and U10423 (N_10423,N_9910,N_9354);
and U10424 (N_10424,N_9912,N_9691);
xor U10425 (N_10425,N_9795,N_9194);
and U10426 (N_10426,N_9084,N_9261);
and U10427 (N_10427,N_9290,N_9135);
nor U10428 (N_10428,N_9815,N_9100);
nor U10429 (N_10429,N_9668,N_9241);
or U10430 (N_10430,N_9864,N_9881);
nand U10431 (N_10431,N_9432,N_9790);
and U10432 (N_10432,N_9794,N_9150);
xor U10433 (N_10433,N_9690,N_9604);
and U10434 (N_10434,N_9692,N_9385);
and U10435 (N_10435,N_9361,N_9935);
nor U10436 (N_10436,N_9849,N_9060);
nor U10437 (N_10437,N_9176,N_9143);
xnor U10438 (N_10438,N_9547,N_9048);
and U10439 (N_10439,N_9672,N_9181);
nand U10440 (N_10440,N_9635,N_9736);
and U10441 (N_10441,N_9576,N_9543);
xor U10442 (N_10442,N_9250,N_9597);
nand U10443 (N_10443,N_9489,N_9462);
and U10444 (N_10444,N_9750,N_9342);
nand U10445 (N_10445,N_9005,N_9479);
xnor U10446 (N_10446,N_9891,N_9461);
nand U10447 (N_10447,N_9665,N_9699);
and U10448 (N_10448,N_9756,N_9853);
nor U10449 (N_10449,N_9706,N_9793);
or U10450 (N_10450,N_9282,N_9144);
or U10451 (N_10451,N_9187,N_9634);
xor U10452 (N_10452,N_9438,N_9420);
or U10453 (N_10453,N_9184,N_9843);
nor U10454 (N_10454,N_9887,N_9491);
nor U10455 (N_10455,N_9095,N_9673);
xnor U10456 (N_10456,N_9477,N_9174);
nor U10457 (N_10457,N_9002,N_9978);
or U10458 (N_10458,N_9206,N_9596);
xor U10459 (N_10459,N_9804,N_9094);
or U10460 (N_10460,N_9742,N_9743);
nor U10461 (N_10461,N_9571,N_9431);
xnor U10462 (N_10462,N_9083,N_9873);
and U10463 (N_10463,N_9723,N_9496);
nor U10464 (N_10464,N_9980,N_9046);
or U10465 (N_10465,N_9514,N_9195);
and U10466 (N_10466,N_9316,N_9018);
and U10467 (N_10467,N_9180,N_9778);
xnor U10468 (N_10468,N_9363,N_9924);
xor U10469 (N_10469,N_9930,N_9575);
nand U10470 (N_10470,N_9703,N_9581);
or U10471 (N_10471,N_9081,N_9740);
or U10472 (N_10472,N_9939,N_9183);
xnor U10473 (N_10473,N_9693,N_9251);
nand U10474 (N_10474,N_9416,N_9167);
and U10475 (N_10475,N_9763,N_9114);
xnor U10476 (N_10476,N_9237,N_9746);
or U10477 (N_10477,N_9838,N_9229);
xnor U10478 (N_10478,N_9395,N_9179);
nand U10479 (N_10479,N_9440,N_9899);
nand U10480 (N_10480,N_9373,N_9654);
nand U10481 (N_10481,N_9592,N_9284);
nor U10482 (N_10482,N_9857,N_9937);
or U10483 (N_10483,N_9698,N_9772);
nor U10484 (N_10484,N_9641,N_9649);
and U10485 (N_10485,N_9351,N_9331);
and U10486 (N_10486,N_9379,N_9098);
nand U10487 (N_10487,N_9301,N_9360);
xor U10488 (N_10488,N_9428,N_9560);
nor U10489 (N_10489,N_9026,N_9197);
and U10490 (N_10490,N_9182,N_9689);
or U10491 (N_10491,N_9890,N_9900);
nor U10492 (N_10492,N_9056,N_9555);
or U10493 (N_10493,N_9142,N_9038);
or U10494 (N_10494,N_9175,N_9904);
or U10495 (N_10495,N_9792,N_9626);
or U10496 (N_10496,N_9347,N_9579);
and U10497 (N_10497,N_9704,N_9551);
or U10498 (N_10498,N_9578,N_9955);
or U10499 (N_10499,N_9403,N_9940);
and U10500 (N_10500,N_9744,N_9039);
nand U10501 (N_10501,N_9186,N_9004);
nor U10502 (N_10502,N_9525,N_9952);
or U10503 (N_10503,N_9860,N_9856);
nor U10504 (N_10504,N_9466,N_9717);
nor U10505 (N_10505,N_9422,N_9410);
or U10506 (N_10506,N_9372,N_9279);
nor U10507 (N_10507,N_9022,N_9949);
nand U10508 (N_10508,N_9784,N_9369);
or U10509 (N_10509,N_9256,N_9685);
or U10510 (N_10510,N_9317,N_9805);
nand U10511 (N_10511,N_9540,N_9012);
or U10512 (N_10512,N_9641,N_9339);
nor U10513 (N_10513,N_9860,N_9801);
or U10514 (N_10514,N_9048,N_9259);
nor U10515 (N_10515,N_9970,N_9238);
or U10516 (N_10516,N_9268,N_9693);
or U10517 (N_10517,N_9993,N_9418);
or U10518 (N_10518,N_9899,N_9203);
and U10519 (N_10519,N_9770,N_9291);
nand U10520 (N_10520,N_9699,N_9185);
and U10521 (N_10521,N_9537,N_9786);
xor U10522 (N_10522,N_9696,N_9108);
and U10523 (N_10523,N_9771,N_9152);
nor U10524 (N_10524,N_9339,N_9821);
or U10525 (N_10525,N_9009,N_9602);
nand U10526 (N_10526,N_9450,N_9874);
and U10527 (N_10527,N_9543,N_9980);
nand U10528 (N_10528,N_9225,N_9696);
nor U10529 (N_10529,N_9775,N_9339);
and U10530 (N_10530,N_9407,N_9051);
or U10531 (N_10531,N_9214,N_9509);
xor U10532 (N_10532,N_9455,N_9600);
nand U10533 (N_10533,N_9208,N_9720);
xor U10534 (N_10534,N_9346,N_9479);
or U10535 (N_10535,N_9840,N_9184);
nand U10536 (N_10536,N_9178,N_9271);
nand U10537 (N_10537,N_9899,N_9129);
or U10538 (N_10538,N_9498,N_9615);
xnor U10539 (N_10539,N_9197,N_9948);
and U10540 (N_10540,N_9669,N_9788);
or U10541 (N_10541,N_9023,N_9207);
nand U10542 (N_10542,N_9106,N_9105);
xor U10543 (N_10543,N_9383,N_9569);
xnor U10544 (N_10544,N_9409,N_9355);
nand U10545 (N_10545,N_9291,N_9986);
nand U10546 (N_10546,N_9822,N_9414);
or U10547 (N_10547,N_9243,N_9980);
nand U10548 (N_10548,N_9790,N_9462);
xor U10549 (N_10549,N_9781,N_9973);
or U10550 (N_10550,N_9131,N_9341);
or U10551 (N_10551,N_9661,N_9533);
xor U10552 (N_10552,N_9057,N_9179);
xnor U10553 (N_10553,N_9282,N_9604);
nand U10554 (N_10554,N_9251,N_9982);
and U10555 (N_10555,N_9970,N_9228);
xor U10556 (N_10556,N_9385,N_9533);
or U10557 (N_10557,N_9615,N_9823);
nand U10558 (N_10558,N_9722,N_9845);
nand U10559 (N_10559,N_9102,N_9443);
xnor U10560 (N_10560,N_9778,N_9579);
or U10561 (N_10561,N_9117,N_9916);
nand U10562 (N_10562,N_9523,N_9423);
nand U10563 (N_10563,N_9391,N_9928);
or U10564 (N_10564,N_9192,N_9077);
nor U10565 (N_10565,N_9215,N_9727);
nor U10566 (N_10566,N_9568,N_9099);
nand U10567 (N_10567,N_9463,N_9779);
xor U10568 (N_10568,N_9510,N_9020);
nand U10569 (N_10569,N_9901,N_9823);
nor U10570 (N_10570,N_9027,N_9093);
and U10571 (N_10571,N_9964,N_9015);
and U10572 (N_10572,N_9794,N_9871);
or U10573 (N_10573,N_9712,N_9855);
or U10574 (N_10574,N_9456,N_9567);
or U10575 (N_10575,N_9992,N_9327);
and U10576 (N_10576,N_9296,N_9781);
nor U10577 (N_10577,N_9654,N_9785);
nor U10578 (N_10578,N_9086,N_9923);
nand U10579 (N_10579,N_9765,N_9619);
nor U10580 (N_10580,N_9883,N_9192);
nand U10581 (N_10581,N_9282,N_9575);
nand U10582 (N_10582,N_9517,N_9729);
or U10583 (N_10583,N_9116,N_9319);
and U10584 (N_10584,N_9392,N_9533);
and U10585 (N_10585,N_9756,N_9725);
or U10586 (N_10586,N_9803,N_9013);
nand U10587 (N_10587,N_9256,N_9280);
nand U10588 (N_10588,N_9669,N_9656);
nor U10589 (N_10589,N_9326,N_9398);
nor U10590 (N_10590,N_9668,N_9362);
nand U10591 (N_10591,N_9234,N_9931);
and U10592 (N_10592,N_9982,N_9556);
nor U10593 (N_10593,N_9771,N_9890);
or U10594 (N_10594,N_9055,N_9858);
nor U10595 (N_10595,N_9339,N_9315);
nand U10596 (N_10596,N_9445,N_9526);
nor U10597 (N_10597,N_9241,N_9629);
nand U10598 (N_10598,N_9430,N_9687);
xnor U10599 (N_10599,N_9991,N_9065);
and U10600 (N_10600,N_9497,N_9722);
and U10601 (N_10601,N_9901,N_9122);
nor U10602 (N_10602,N_9950,N_9198);
or U10603 (N_10603,N_9595,N_9351);
nand U10604 (N_10604,N_9507,N_9311);
nand U10605 (N_10605,N_9622,N_9735);
and U10606 (N_10606,N_9072,N_9826);
xnor U10607 (N_10607,N_9500,N_9708);
and U10608 (N_10608,N_9783,N_9127);
nand U10609 (N_10609,N_9027,N_9097);
or U10610 (N_10610,N_9251,N_9080);
or U10611 (N_10611,N_9004,N_9392);
and U10612 (N_10612,N_9875,N_9195);
or U10613 (N_10613,N_9582,N_9274);
nor U10614 (N_10614,N_9594,N_9082);
or U10615 (N_10615,N_9967,N_9795);
and U10616 (N_10616,N_9328,N_9659);
nor U10617 (N_10617,N_9886,N_9960);
xor U10618 (N_10618,N_9907,N_9443);
nor U10619 (N_10619,N_9943,N_9743);
or U10620 (N_10620,N_9203,N_9737);
or U10621 (N_10621,N_9570,N_9268);
nor U10622 (N_10622,N_9497,N_9581);
and U10623 (N_10623,N_9707,N_9556);
and U10624 (N_10624,N_9870,N_9037);
or U10625 (N_10625,N_9047,N_9024);
nand U10626 (N_10626,N_9125,N_9867);
xor U10627 (N_10627,N_9000,N_9928);
xnor U10628 (N_10628,N_9529,N_9148);
or U10629 (N_10629,N_9449,N_9512);
nand U10630 (N_10630,N_9354,N_9597);
nor U10631 (N_10631,N_9741,N_9288);
xnor U10632 (N_10632,N_9355,N_9796);
xor U10633 (N_10633,N_9985,N_9978);
and U10634 (N_10634,N_9746,N_9042);
and U10635 (N_10635,N_9773,N_9178);
and U10636 (N_10636,N_9920,N_9687);
or U10637 (N_10637,N_9807,N_9857);
nor U10638 (N_10638,N_9132,N_9058);
nand U10639 (N_10639,N_9244,N_9262);
and U10640 (N_10640,N_9354,N_9615);
or U10641 (N_10641,N_9260,N_9620);
or U10642 (N_10642,N_9836,N_9078);
xnor U10643 (N_10643,N_9621,N_9231);
and U10644 (N_10644,N_9491,N_9145);
or U10645 (N_10645,N_9699,N_9961);
nor U10646 (N_10646,N_9305,N_9404);
xnor U10647 (N_10647,N_9733,N_9703);
or U10648 (N_10648,N_9262,N_9736);
xnor U10649 (N_10649,N_9017,N_9453);
nor U10650 (N_10650,N_9217,N_9647);
xor U10651 (N_10651,N_9767,N_9575);
nand U10652 (N_10652,N_9716,N_9793);
nand U10653 (N_10653,N_9863,N_9197);
nand U10654 (N_10654,N_9535,N_9765);
or U10655 (N_10655,N_9833,N_9763);
and U10656 (N_10656,N_9922,N_9240);
xnor U10657 (N_10657,N_9790,N_9496);
and U10658 (N_10658,N_9409,N_9650);
xnor U10659 (N_10659,N_9723,N_9611);
xor U10660 (N_10660,N_9547,N_9623);
or U10661 (N_10661,N_9671,N_9581);
or U10662 (N_10662,N_9269,N_9625);
and U10663 (N_10663,N_9344,N_9795);
and U10664 (N_10664,N_9565,N_9144);
nand U10665 (N_10665,N_9253,N_9261);
and U10666 (N_10666,N_9589,N_9474);
nor U10667 (N_10667,N_9973,N_9082);
and U10668 (N_10668,N_9794,N_9066);
nor U10669 (N_10669,N_9898,N_9815);
xor U10670 (N_10670,N_9666,N_9125);
or U10671 (N_10671,N_9462,N_9081);
nand U10672 (N_10672,N_9925,N_9756);
or U10673 (N_10673,N_9270,N_9704);
xnor U10674 (N_10674,N_9515,N_9699);
nor U10675 (N_10675,N_9624,N_9430);
nor U10676 (N_10676,N_9458,N_9672);
and U10677 (N_10677,N_9768,N_9368);
nor U10678 (N_10678,N_9821,N_9759);
and U10679 (N_10679,N_9249,N_9013);
nor U10680 (N_10680,N_9064,N_9492);
xnor U10681 (N_10681,N_9955,N_9839);
or U10682 (N_10682,N_9506,N_9211);
and U10683 (N_10683,N_9764,N_9588);
and U10684 (N_10684,N_9833,N_9983);
xor U10685 (N_10685,N_9539,N_9555);
nor U10686 (N_10686,N_9927,N_9214);
xor U10687 (N_10687,N_9328,N_9577);
nor U10688 (N_10688,N_9001,N_9995);
and U10689 (N_10689,N_9561,N_9176);
xor U10690 (N_10690,N_9426,N_9116);
xnor U10691 (N_10691,N_9149,N_9152);
and U10692 (N_10692,N_9611,N_9470);
or U10693 (N_10693,N_9679,N_9886);
nor U10694 (N_10694,N_9815,N_9573);
nor U10695 (N_10695,N_9521,N_9230);
nand U10696 (N_10696,N_9706,N_9300);
xor U10697 (N_10697,N_9180,N_9020);
and U10698 (N_10698,N_9514,N_9229);
and U10699 (N_10699,N_9602,N_9408);
nand U10700 (N_10700,N_9646,N_9180);
and U10701 (N_10701,N_9612,N_9849);
xnor U10702 (N_10702,N_9019,N_9764);
and U10703 (N_10703,N_9182,N_9978);
nand U10704 (N_10704,N_9947,N_9634);
nand U10705 (N_10705,N_9715,N_9502);
xor U10706 (N_10706,N_9406,N_9111);
or U10707 (N_10707,N_9529,N_9789);
xnor U10708 (N_10708,N_9762,N_9607);
and U10709 (N_10709,N_9787,N_9729);
and U10710 (N_10710,N_9527,N_9928);
and U10711 (N_10711,N_9063,N_9178);
nor U10712 (N_10712,N_9091,N_9240);
or U10713 (N_10713,N_9379,N_9564);
nor U10714 (N_10714,N_9822,N_9922);
nor U10715 (N_10715,N_9004,N_9515);
and U10716 (N_10716,N_9270,N_9074);
and U10717 (N_10717,N_9138,N_9850);
or U10718 (N_10718,N_9007,N_9400);
or U10719 (N_10719,N_9441,N_9573);
and U10720 (N_10720,N_9981,N_9555);
or U10721 (N_10721,N_9500,N_9022);
nor U10722 (N_10722,N_9121,N_9787);
nand U10723 (N_10723,N_9565,N_9778);
or U10724 (N_10724,N_9885,N_9025);
nor U10725 (N_10725,N_9636,N_9483);
nand U10726 (N_10726,N_9890,N_9189);
nor U10727 (N_10727,N_9892,N_9637);
or U10728 (N_10728,N_9257,N_9817);
nor U10729 (N_10729,N_9109,N_9917);
or U10730 (N_10730,N_9853,N_9306);
xor U10731 (N_10731,N_9774,N_9856);
xor U10732 (N_10732,N_9059,N_9714);
and U10733 (N_10733,N_9528,N_9215);
and U10734 (N_10734,N_9793,N_9167);
or U10735 (N_10735,N_9544,N_9833);
nand U10736 (N_10736,N_9201,N_9198);
xor U10737 (N_10737,N_9892,N_9979);
nand U10738 (N_10738,N_9397,N_9227);
nand U10739 (N_10739,N_9061,N_9628);
or U10740 (N_10740,N_9859,N_9428);
and U10741 (N_10741,N_9452,N_9053);
and U10742 (N_10742,N_9782,N_9206);
nand U10743 (N_10743,N_9717,N_9239);
nand U10744 (N_10744,N_9407,N_9043);
and U10745 (N_10745,N_9590,N_9817);
nor U10746 (N_10746,N_9242,N_9685);
or U10747 (N_10747,N_9503,N_9142);
and U10748 (N_10748,N_9691,N_9689);
xor U10749 (N_10749,N_9387,N_9038);
nor U10750 (N_10750,N_9545,N_9336);
or U10751 (N_10751,N_9594,N_9166);
nor U10752 (N_10752,N_9568,N_9147);
or U10753 (N_10753,N_9567,N_9449);
and U10754 (N_10754,N_9903,N_9855);
and U10755 (N_10755,N_9970,N_9365);
nor U10756 (N_10756,N_9812,N_9905);
nor U10757 (N_10757,N_9340,N_9805);
nor U10758 (N_10758,N_9621,N_9872);
nand U10759 (N_10759,N_9261,N_9947);
xor U10760 (N_10760,N_9322,N_9789);
xor U10761 (N_10761,N_9803,N_9298);
or U10762 (N_10762,N_9662,N_9155);
nor U10763 (N_10763,N_9580,N_9728);
xor U10764 (N_10764,N_9051,N_9038);
or U10765 (N_10765,N_9881,N_9504);
nor U10766 (N_10766,N_9665,N_9216);
or U10767 (N_10767,N_9800,N_9819);
nor U10768 (N_10768,N_9769,N_9192);
nand U10769 (N_10769,N_9195,N_9094);
xnor U10770 (N_10770,N_9216,N_9137);
or U10771 (N_10771,N_9471,N_9605);
or U10772 (N_10772,N_9765,N_9548);
xnor U10773 (N_10773,N_9581,N_9563);
nor U10774 (N_10774,N_9538,N_9560);
and U10775 (N_10775,N_9565,N_9373);
nor U10776 (N_10776,N_9829,N_9058);
or U10777 (N_10777,N_9092,N_9079);
and U10778 (N_10778,N_9223,N_9573);
xor U10779 (N_10779,N_9280,N_9339);
nand U10780 (N_10780,N_9757,N_9296);
or U10781 (N_10781,N_9796,N_9564);
xor U10782 (N_10782,N_9556,N_9957);
nand U10783 (N_10783,N_9627,N_9160);
xor U10784 (N_10784,N_9335,N_9296);
nand U10785 (N_10785,N_9745,N_9110);
nor U10786 (N_10786,N_9384,N_9792);
and U10787 (N_10787,N_9320,N_9645);
or U10788 (N_10788,N_9616,N_9284);
nand U10789 (N_10789,N_9143,N_9101);
and U10790 (N_10790,N_9533,N_9842);
xnor U10791 (N_10791,N_9779,N_9923);
or U10792 (N_10792,N_9980,N_9880);
nor U10793 (N_10793,N_9012,N_9598);
nor U10794 (N_10794,N_9183,N_9677);
and U10795 (N_10795,N_9192,N_9404);
nor U10796 (N_10796,N_9245,N_9099);
or U10797 (N_10797,N_9351,N_9083);
xor U10798 (N_10798,N_9826,N_9111);
xnor U10799 (N_10799,N_9682,N_9897);
or U10800 (N_10800,N_9454,N_9941);
or U10801 (N_10801,N_9198,N_9879);
nor U10802 (N_10802,N_9950,N_9114);
nor U10803 (N_10803,N_9690,N_9606);
nand U10804 (N_10804,N_9666,N_9652);
and U10805 (N_10805,N_9264,N_9914);
or U10806 (N_10806,N_9056,N_9988);
nand U10807 (N_10807,N_9019,N_9408);
or U10808 (N_10808,N_9950,N_9346);
nor U10809 (N_10809,N_9531,N_9717);
and U10810 (N_10810,N_9363,N_9409);
xor U10811 (N_10811,N_9886,N_9930);
and U10812 (N_10812,N_9127,N_9717);
or U10813 (N_10813,N_9727,N_9783);
xor U10814 (N_10814,N_9067,N_9608);
nand U10815 (N_10815,N_9961,N_9999);
nand U10816 (N_10816,N_9455,N_9679);
nand U10817 (N_10817,N_9611,N_9614);
nand U10818 (N_10818,N_9379,N_9205);
and U10819 (N_10819,N_9905,N_9527);
nand U10820 (N_10820,N_9870,N_9287);
nand U10821 (N_10821,N_9403,N_9299);
or U10822 (N_10822,N_9787,N_9233);
nand U10823 (N_10823,N_9682,N_9806);
nand U10824 (N_10824,N_9450,N_9971);
and U10825 (N_10825,N_9451,N_9101);
nand U10826 (N_10826,N_9782,N_9274);
nor U10827 (N_10827,N_9280,N_9691);
or U10828 (N_10828,N_9247,N_9940);
and U10829 (N_10829,N_9715,N_9858);
nor U10830 (N_10830,N_9728,N_9571);
xor U10831 (N_10831,N_9527,N_9037);
nor U10832 (N_10832,N_9118,N_9970);
and U10833 (N_10833,N_9846,N_9762);
nor U10834 (N_10834,N_9541,N_9037);
nand U10835 (N_10835,N_9307,N_9323);
or U10836 (N_10836,N_9109,N_9423);
nor U10837 (N_10837,N_9350,N_9712);
nor U10838 (N_10838,N_9966,N_9087);
and U10839 (N_10839,N_9502,N_9530);
nor U10840 (N_10840,N_9377,N_9696);
nand U10841 (N_10841,N_9442,N_9193);
xnor U10842 (N_10842,N_9344,N_9965);
or U10843 (N_10843,N_9396,N_9803);
or U10844 (N_10844,N_9310,N_9234);
and U10845 (N_10845,N_9947,N_9244);
or U10846 (N_10846,N_9613,N_9527);
and U10847 (N_10847,N_9895,N_9880);
nor U10848 (N_10848,N_9958,N_9188);
xor U10849 (N_10849,N_9093,N_9412);
xnor U10850 (N_10850,N_9738,N_9504);
xnor U10851 (N_10851,N_9053,N_9599);
or U10852 (N_10852,N_9248,N_9727);
nor U10853 (N_10853,N_9279,N_9269);
xnor U10854 (N_10854,N_9804,N_9058);
nor U10855 (N_10855,N_9700,N_9987);
and U10856 (N_10856,N_9502,N_9238);
nor U10857 (N_10857,N_9168,N_9227);
xnor U10858 (N_10858,N_9461,N_9809);
xnor U10859 (N_10859,N_9407,N_9266);
and U10860 (N_10860,N_9459,N_9181);
xor U10861 (N_10861,N_9929,N_9293);
or U10862 (N_10862,N_9039,N_9507);
nand U10863 (N_10863,N_9279,N_9584);
xnor U10864 (N_10864,N_9352,N_9643);
nand U10865 (N_10865,N_9594,N_9950);
nor U10866 (N_10866,N_9636,N_9481);
or U10867 (N_10867,N_9989,N_9176);
nor U10868 (N_10868,N_9677,N_9460);
or U10869 (N_10869,N_9852,N_9438);
nand U10870 (N_10870,N_9419,N_9351);
nor U10871 (N_10871,N_9100,N_9232);
and U10872 (N_10872,N_9166,N_9852);
and U10873 (N_10873,N_9208,N_9482);
xnor U10874 (N_10874,N_9321,N_9092);
nand U10875 (N_10875,N_9259,N_9008);
nor U10876 (N_10876,N_9329,N_9929);
and U10877 (N_10877,N_9401,N_9611);
or U10878 (N_10878,N_9235,N_9594);
nor U10879 (N_10879,N_9173,N_9714);
nor U10880 (N_10880,N_9245,N_9398);
nor U10881 (N_10881,N_9382,N_9834);
and U10882 (N_10882,N_9824,N_9392);
nand U10883 (N_10883,N_9239,N_9166);
nor U10884 (N_10884,N_9539,N_9836);
or U10885 (N_10885,N_9195,N_9206);
or U10886 (N_10886,N_9229,N_9620);
nand U10887 (N_10887,N_9955,N_9697);
or U10888 (N_10888,N_9360,N_9786);
xor U10889 (N_10889,N_9212,N_9065);
or U10890 (N_10890,N_9635,N_9875);
nand U10891 (N_10891,N_9090,N_9921);
nor U10892 (N_10892,N_9648,N_9903);
or U10893 (N_10893,N_9563,N_9363);
and U10894 (N_10894,N_9101,N_9300);
nor U10895 (N_10895,N_9069,N_9416);
or U10896 (N_10896,N_9621,N_9545);
nand U10897 (N_10897,N_9100,N_9700);
or U10898 (N_10898,N_9800,N_9471);
and U10899 (N_10899,N_9472,N_9519);
or U10900 (N_10900,N_9085,N_9804);
nor U10901 (N_10901,N_9816,N_9014);
or U10902 (N_10902,N_9663,N_9946);
and U10903 (N_10903,N_9035,N_9724);
nand U10904 (N_10904,N_9282,N_9915);
nand U10905 (N_10905,N_9693,N_9033);
nor U10906 (N_10906,N_9678,N_9983);
and U10907 (N_10907,N_9238,N_9357);
and U10908 (N_10908,N_9846,N_9415);
nor U10909 (N_10909,N_9679,N_9386);
xor U10910 (N_10910,N_9176,N_9721);
and U10911 (N_10911,N_9131,N_9413);
nand U10912 (N_10912,N_9733,N_9066);
and U10913 (N_10913,N_9427,N_9129);
and U10914 (N_10914,N_9663,N_9777);
nor U10915 (N_10915,N_9873,N_9865);
xor U10916 (N_10916,N_9885,N_9608);
xor U10917 (N_10917,N_9967,N_9194);
nand U10918 (N_10918,N_9853,N_9576);
xor U10919 (N_10919,N_9481,N_9122);
nor U10920 (N_10920,N_9024,N_9438);
nand U10921 (N_10921,N_9997,N_9827);
or U10922 (N_10922,N_9037,N_9827);
and U10923 (N_10923,N_9323,N_9180);
or U10924 (N_10924,N_9674,N_9533);
or U10925 (N_10925,N_9391,N_9927);
nor U10926 (N_10926,N_9171,N_9915);
or U10927 (N_10927,N_9897,N_9767);
and U10928 (N_10928,N_9107,N_9239);
and U10929 (N_10929,N_9720,N_9607);
nor U10930 (N_10930,N_9482,N_9733);
and U10931 (N_10931,N_9695,N_9895);
xnor U10932 (N_10932,N_9982,N_9736);
nor U10933 (N_10933,N_9743,N_9801);
xnor U10934 (N_10934,N_9702,N_9822);
nor U10935 (N_10935,N_9941,N_9511);
nor U10936 (N_10936,N_9237,N_9944);
and U10937 (N_10937,N_9874,N_9889);
nor U10938 (N_10938,N_9419,N_9945);
or U10939 (N_10939,N_9152,N_9323);
and U10940 (N_10940,N_9749,N_9564);
xnor U10941 (N_10941,N_9165,N_9123);
and U10942 (N_10942,N_9443,N_9126);
xnor U10943 (N_10943,N_9818,N_9012);
nor U10944 (N_10944,N_9662,N_9417);
nand U10945 (N_10945,N_9509,N_9149);
or U10946 (N_10946,N_9460,N_9090);
xor U10947 (N_10947,N_9344,N_9959);
nor U10948 (N_10948,N_9789,N_9877);
nand U10949 (N_10949,N_9710,N_9587);
nand U10950 (N_10950,N_9037,N_9937);
nand U10951 (N_10951,N_9029,N_9239);
nor U10952 (N_10952,N_9004,N_9666);
and U10953 (N_10953,N_9587,N_9781);
nor U10954 (N_10954,N_9419,N_9129);
or U10955 (N_10955,N_9522,N_9293);
and U10956 (N_10956,N_9808,N_9918);
or U10957 (N_10957,N_9774,N_9423);
nor U10958 (N_10958,N_9623,N_9941);
and U10959 (N_10959,N_9823,N_9026);
xor U10960 (N_10960,N_9019,N_9131);
nor U10961 (N_10961,N_9853,N_9630);
nand U10962 (N_10962,N_9174,N_9349);
nand U10963 (N_10963,N_9890,N_9410);
or U10964 (N_10964,N_9451,N_9908);
nand U10965 (N_10965,N_9710,N_9660);
nand U10966 (N_10966,N_9519,N_9754);
nand U10967 (N_10967,N_9458,N_9206);
or U10968 (N_10968,N_9494,N_9802);
xor U10969 (N_10969,N_9229,N_9035);
nor U10970 (N_10970,N_9395,N_9298);
xnor U10971 (N_10971,N_9563,N_9259);
nand U10972 (N_10972,N_9874,N_9206);
or U10973 (N_10973,N_9312,N_9277);
and U10974 (N_10974,N_9495,N_9014);
nand U10975 (N_10975,N_9971,N_9269);
or U10976 (N_10976,N_9489,N_9769);
xnor U10977 (N_10977,N_9114,N_9687);
nand U10978 (N_10978,N_9708,N_9298);
and U10979 (N_10979,N_9786,N_9354);
or U10980 (N_10980,N_9025,N_9314);
and U10981 (N_10981,N_9119,N_9618);
nor U10982 (N_10982,N_9550,N_9799);
nand U10983 (N_10983,N_9015,N_9375);
nor U10984 (N_10984,N_9520,N_9981);
and U10985 (N_10985,N_9199,N_9269);
nand U10986 (N_10986,N_9700,N_9118);
or U10987 (N_10987,N_9538,N_9774);
and U10988 (N_10988,N_9592,N_9833);
nand U10989 (N_10989,N_9402,N_9857);
nand U10990 (N_10990,N_9343,N_9678);
and U10991 (N_10991,N_9609,N_9944);
xor U10992 (N_10992,N_9572,N_9448);
and U10993 (N_10993,N_9086,N_9025);
or U10994 (N_10994,N_9874,N_9305);
or U10995 (N_10995,N_9829,N_9271);
or U10996 (N_10996,N_9255,N_9327);
nand U10997 (N_10997,N_9864,N_9699);
or U10998 (N_10998,N_9087,N_9996);
xnor U10999 (N_10999,N_9155,N_9683);
and U11000 (N_11000,N_10431,N_10256);
and U11001 (N_11001,N_10651,N_10535);
nand U11002 (N_11002,N_10037,N_10747);
xor U11003 (N_11003,N_10975,N_10252);
xor U11004 (N_11004,N_10287,N_10623);
nor U11005 (N_11005,N_10277,N_10600);
nor U11006 (N_11006,N_10095,N_10463);
nor U11007 (N_11007,N_10611,N_10648);
nand U11008 (N_11008,N_10935,N_10384);
nor U11009 (N_11009,N_10634,N_10061);
nand U11010 (N_11010,N_10661,N_10808);
nor U11011 (N_11011,N_10034,N_10388);
nor U11012 (N_11012,N_10212,N_10154);
xnor U11013 (N_11013,N_10862,N_10342);
nor U11014 (N_11014,N_10225,N_10358);
xnor U11015 (N_11015,N_10289,N_10199);
and U11016 (N_11016,N_10314,N_10647);
and U11017 (N_11017,N_10806,N_10950);
xor U11018 (N_11018,N_10231,N_10652);
xor U11019 (N_11019,N_10090,N_10169);
nand U11020 (N_11020,N_10970,N_10695);
nand U11021 (N_11021,N_10297,N_10015);
xnor U11022 (N_11022,N_10163,N_10509);
nand U11023 (N_11023,N_10493,N_10016);
or U11024 (N_11024,N_10189,N_10552);
or U11025 (N_11025,N_10621,N_10781);
nor U11026 (N_11026,N_10292,N_10045);
nand U11027 (N_11027,N_10629,N_10119);
nand U11028 (N_11028,N_10859,N_10641);
and U11029 (N_11029,N_10068,N_10850);
nand U11030 (N_11030,N_10672,N_10805);
xor U11031 (N_11031,N_10481,N_10944);
nand U11032 (N_11032,N_10929,N_10356);
nor U11033 (N_11033,N_10103,N_10098);
nand U11034 (N_11034,N_10601,N_10195);
nand U11035 (N_11035,N_10448,N_10296);
or U11036 (N_11036,N_10395,N_10844);
nand U11037 (N_11037,N_10821,N_10952);
xor U11038 (N_11038,N_10827,N_10876);
xnor U11039 (N_11039,N_10495,N_10976);
or U11040 (N_11040,N_10529,N_10357);
xor U11041 (N_11041,N_10478,N_10345);
nor U11042 (N_11042,N_10698,N_10456);
xnor U11043 (N_11043,N_10108,N_10339);
xor U11044 (N_11044,N_10051,N_10926);
or U11045 (N_11045,N_10590,N_10819);
and U11046 (N_11046,N_10943,N_10525);
nor U11047 (N_11047,N_10288,N_10700);
xnor U11048 (N_11048,N_10500,N_10502);
nor U11049 (N_11049,N_10579,N_10053);
nand U11050 (N_11050,N_10183,N_10749);
xor U11051 (N_11051,N_10304,N_10458);
nand U11052 (N_11052,N_10788,N_10856);
or U11053 (N_11053,N_10804,N_10620);
nor U11054 (N_11054,N_10526,N_10884);
and U11055 (N_11055,N_10278,N_10379);
nand U11056 (N_11056,N_10708,N_10348);
and U11057 (N_11057,N_10073,N_10030);
nand U11058 (N_11058,N_10991,N_10476);
nand U11059 (N_11059,N_10838,N_10835);
nor U11060 (N_11060,N_10956,N_10308);
or U11061 (N_11061,N_10742,N_10176);
nor U11062 (N_11062,N_10168,N_10736);
or U11063 (N_11063,N_10200,N_10043);
xor U11064 (N_11064,N_10038,N_10482);
xor U11065 (N_11065,N_10177,N_10128);
and U11066 (N_11066,N_10100,N_10491);
nand U11067 (N_11067,N_10717,N_10849);
nand U11068 (N_11068,N_10429,N_10414);
xnor U11069 (N_11069,N_10811,N_10673);
nor U11070 (N_11070,N_10837,N_10640);
nor U11071 (N_11071,N_10024,N_10261);
and U11072 (N_11072,N_10487,N_10778);
xor U11073 (N_11073,N_10934,N_10796);
nand U11074 (N_11074,N_10836,N_10910);
or U11075 (N_11075,N_10932,N_10851);
nor U11076 (N_11076,N_10109,N_10550);
or U11077 (N_11077,N_10556,N_10069);
nand U11078 (N_11078,N_10587,N_10421);
xnor U11079 (N_11079,N_10639,N_10813);
nand U11080 (N_11080,N_10219,N_10228);
nand U11081 (N_11081,N_10973,N_10839);
xor U11082 (N_11082,N_10483,N_10179);
nand U11083 (N_11083,N_10178,N_10479);
or U11084 (N_11084,N_10980,N_10968);
xnor U11085 (N_11085,N_10113,N_10000);
xor U11086 (N_11086,N_10824,N_10832);
nand U11087 (N_11087,N_10899,N_10263);
nor U11088 (N_11088,N_10055,N_10086);
and U11089 (N_11089,N_10925,N_10792);
and U11090 (N_11090,N_10675,N_10011);
xor U11091 (N_11091,N_10399,N_10592);
xor U11092 (N_11092,N_10933,N_10918);
nand U11093 (N_11093,N_10696,N_10580);
and U11094 (N_11094,N_10873,N_10951);
or U11095 (N_11095,N_10561,N_10609);
nor U11096 (N_11096,N_10274,N_10092);
and U11097 (N_11097,N_10398,N_10180);
or U11098 (N_11098,N_10924,N_10711);
xnor U11099 (N_11099,N_10149,N_10426);
or U11100 (N_11100,N_10988,N_10901);
or U11101 (N_11101,N_10117,N_10786);
or U11102 (N_11102,N_10834,N_10891);
or U11103 (N_11103,N_10793,N_10449);
nand U11104 (N_11104,N_10267,N_10337);
nand U11105 (N_11105,N_10032,N_10948);
or U11106 (N_11106,N_10567,N_10887);
and U11107 (N_11107,N_10236,N_10983);
and U11108 (N_11108,N_10852,N_10542);
and U11109 (N_11109,N_10381,N_10420);
or U11110 (N_11110,N_10576,N_10725);
xor U11111 (N_11111,N_10662,N_10001);
nand U11112 (N_11112,N_10816,N_10863);
xnor U11113 (N_11113,N_10941,N_10898);
nor U11114 (N_11114,N_10949,N_10018);
or U11115 (N_11115,N_10280,N_10074);
and U11116 (N_11116,N_10057,N_10488);
nand U11117 (N_11117,N_10440,N_10211);
nor U11118 (N_11118,N_10266,N_10779);
xnor U11119 (N_11119,N_10638,N_10966);
and U11120 (N_11120,N_10574,N_10597);
and U11121 (N_11121,N_10503,N_10846);
nand U11122 (N_11122,N_10960,N_10194);
nand U11123 (N_11123,N_10869,N_10294);
nand U11124 (N_11124,N_10689,N_10624);
xor U11125 (N_11125,N_10208,N_10124);
nor U11126 (N_11126,N_10151,N_10114);
xor U11127 (N_11127,N_10247,N_10373);
nor U11128 (N_11128,N_10271,N_10541);
and U11129 (N_11129,N_10222,N_10939);
nor U11130 (N_11130,N_10632,N_10190);
xor U11131 (N_11131,N_10602,N_10082);
xnor U11132 (N_11132,N_10853,N_10413);
and U11133 (N_11133,N_10235,N_10706);
nand U11134 (N_11134,N_10136,N_10870);
or U11135 (N_11135,N_10275,N_10921);
and U11136 (N_11136,N_10106,N_10389);
nor U11137 (N_11137,N_10729,N_10982);
xor U11138 (N_11138,N_10378,N_10671);
or U11139 (N_11139,N_10807,N_10979);
or U11140 (N_11140,N_10336,N_10344);
xor U11141 (N_11141,N_10759,N_10454);
nor U11142 (N_11142,N_10210,N_10115);
or U11143 (N_11143,N_10709,N_10403);
nor U11144 (N_11144,N_10052,N_10062);
nor U11145 (N_11145,N_10505,N_10974);
or U11146 (N_11146,N_10466,N_10627);
and U11147 (N_11147,N_10299,N_10351);
nor U11148 (N_11148,N_10833,N_10202);
and U11149 (N_11149,N_10368,N_10441);
nand U11150 (N_11150,N_10841,N_10260);
xnor U11151 (N_11151,N_10003,N_10452);
xnor U11152 (N_11152,N_10787,N_10059);
xnor U11153 (N_11153,N_10291,N_10654);
or U11154 (N_11154,N_10138,N_10528);
xnor U11155 (N_11155,N_10474,N_10548);
nand U11156 (N_11156,N_10911,N_10460);
and U11157 (N_11157,N_10930,N_10223);
xor U11158 (N_11158,N_10866,N_10945);
and U11159 (N_11159,N_10522,N_10310);
nor U11160 (N_11160,N_10721,N_10005);
and U11161 (N_11161,N_10822,N_10360);
xnor U11162 (N_11162,N_10251,N_10566);
nor U11163 (N_11163,N_10931,N_10328);
or U11164 (N_11164,N_10947,N_10723);
and U11165 (N_11165,N_10126,N_10089);
or U11166 (N_11166,N_10942,N_10048);
xor U11167 (N_11167,N_10265,N_10447);
xor U11168 (N_11168,N_10795,N_10965);
nand U11169 (N_11169,N_10727,N_10442);
nor U11170 (N_11170,N_10175,N_10101);
xnor U11171 (N_11171,N_10380,N_10820);
xnor U11172 (N_11172,N_10083,N_10205);
nand U11173 (N_11173,N_10715,N_10993);
or U11174 (N_11174,N_10570,N_10547);
and U11175 (N_11175,N_10913,N_10171);
and U11176 (N_11176,N_10655,N_10889);
and U11177 (N_11177,N_10847,N_10506);
nor U11178 (N_11178,N_10760,N_10046);
xnor U11179 (N_11179,N_10283,N_10237);
and U11180 (N_11180,N_10519,N_10033);
nand U11181 (N_11181,N_10740,N_10578);
nor U11182 (N_11182,N_10305,N_10318);
nand U11183 (N_11183,N_10707,N_10739);
xnor U11184 (N_11184,N_10042,N_10741);
and U11185 (N_11185,N_10582,N_10025);
nand U11186 (N_11186,N_10686,N_10879);
nand U11187 (N_11187,N_10192,N_10718);
nand U11188 (N_11188,N_10814,N_10354);
and U11189 (N_11189,N_10099,N_10293);
or U11190 (N_11190,N_10860,N_10244);
or U11191 (N_11191,N_10625,N_10303);
and U11192 (N_11192,N_10981,N_10656);
and U11193 (N_11193,N_10613,N_10152);
xor U11194 (N_11194,N_10307,N_10094);
nand U11195 (N_11195,N_10146,N_10990);
xnor U11196 (N_11196,N_10728,N_10087);
nor U11197 (N_11197,N_10664,N_10054);
nand U11198 (N_11198,N_10810,N_10510);
nand U11199 (N_11199,N_10897,N_10070);
or U11200 (N_11200,N_10167,N_10455);
or U11201 (N_11201,N_10894,N_10667);
and U11202 (N_11202,N_10817,N_10184);
nand U11203 (N_11203,N_10226,N_10216);
nand U11204 (N_11204,N_10644,N_10485);
or U11205 (N_11205,N_10010,N_10014);
nand U11206 (N_11206,N_10181,N_10618);
xnor U11207 (N_11207,N_10058,N_10676);
and U11208 (N_11208,N_10703,N_10412);
or U11209 (N_11209,N_10245,N_10464);
nand U11210 (N_11210,N_10912,N_10369);
nand U11211 (N_11211,N_10206,N_10701);
nor U11212 (N_11212,N_10674,N_10524);
xor U11213 (N_11213,N_10290,N_10484);
and U11214 (N_11214,N_10568,N_10188);
xor U11215 (N_11215,N_10300,N_10875);
nor U11216 (N_11216,N_10435,N_10669);
and U11217 (N_11217,N_10699,N_10799);
xnor U11218 (N_11218,N_10955,N_10593);
xnor U11219 (N_11219,N_10645,N_10311);
and U11220 (N_11220,N_10050,N_10868);
and U11221 (N_11221,N_10332,N_10682);
xnor U11222 (N_11222,N_10681,N_10253);
nor U11223 (N_11223,N_10936,N_10122);
nor U11224 (N_11224,N_10325,N_10697);
nand U11225 (N_11225,N_10513,N_10610);
nand U11226 (N_11226,N_10916,N_10159);
xor U11227 (N_11227,N_10688,N_10423);
xor U11228 (N_11228,N_10797,N_10864);
and U11229 (N_11229,N_10782,N_10145);
nor U11230 (N_11230,N_10995,N_10677);
and U11231 (N_11231,N_10013,N_10815);
and U11232 (N_11232,N_10313,N_10858);
nand U11233 (N_11233,N_10143,N_10017);
xnor U11234 (N_11234,N_10480,N_10665);
xor U11235 (N_11235,N_10402,N_10044);
nand U11236 (N_11236,N_10229,N_10374);
xnor U11237 (N_11237,N_10588,N_10599);
and U11238 (N_11238,N_10660,N_10241);
nand U11239 (N_11239,N_10963,N_10893);
nand U11240 (N_11240,N_10872,N_10534);
xor U11241 (N_11241,N_10400,N_10573);
and U11242 (N_11242,N_10996,N_10987);
nor U11243 (N_11243,N_10319,N_10830);
and U11244 (N_11244,N_10238,N_10321);
or U11245 (N_11245,N_10767,N_10475);
nand U11246 (N_11246,N_10954,N_10755);
or U11247 (N_11247,N_10730,N_10465);
or U11248 (N_11248,N_10773,N_10735);
and U11249 (N_11249,N_10022,N_10908);
nor U11250 (N_11250,N_10006,N_10221);
nor U11251 (N_11251,N_10446,N_10978);
or U11252 (N_11252,N_10007,N_10432);
nand U11253 (N_11253,N_10093,N_10826);
nand U11254 (N_11254,N_10603,N_10492);
nor U11255 (N_11255,N_10232,N_10586);
xor U11256 (N_11256,N_10361,N_10085);
and U11257 (N_11257,N_10371,N_10326);
or U11258 (N_11258,N_10433,N_10915);
xor U11259 (N_11259,N_10774,N_10067);
or U11260 (N_11260,N_10196,N_10877);
and U11261 (N_11261,N_10683,N_10763);
xor U11262 (N_11262,N_10035,N_10545);
xnor U11263 (N_11263,N_10331,N_10233);
and U11264 (N_11264,N_10540,N_10418);
and U11265 (N_11265,N_10078,N_10713);
or U11266 (N_11266,N_10129,N_10410);
nand U11267 (N_11267,N_10914,N_10753);
or U11268 (N_11268,N_10633,N_10327);
or U11269 (N_11269,N_10783,N_10091);
nor U11270 (N_11270,N_10992,N_10514);
and U11271 (N_11271,N_10997,N_10445);
or U11272 (N_11272,N_10619,N_10131);
xor U11273 (N_11273,N_10315,N_10594);
nand U11274 (N_11274,N_10752,N_10557);
xnor U11275 (N_11275,N_10121,N_10900);
xor U11276 (N_11276,N_10551,N_10439);
and U11277 (N_11277,N_10306,N_10104);
nor U11278 (N_11278,N_10273,N_10111);
nor U11279 (N_11279,N_10469,N_10857);
nand U11280 (N_11280,N_10262,N_10498);
or U11281 (N_11281,N_10768,N_10546);
and U11282 (N_11282,N_10880,N_10207);
nand U11283 (N_11283,N_10720,N_10972);
or U11284 (N_11284,N_10434,N_10867);
nand U11285 (N_11285,N_10692,N_10854);
nand U11286 (N_11286,N_10964,N_10702);
and U11287 (N_11287,N_10809,N_10130);
and U11288 (N_11288,N_10153,N_10653);
nand U11289 (N_11289,N_10407,N_10563);
xor U11290 (N_11290,N_10451,N_10906);
nor U11291 (N_11291,N_10614,N_10330);
or U11292 (N_11292,N_10516,N_10878);
xnor U11293 (N_11293,N_10575,N_10425);
nor U11294 (N_11294,N_10443,N_10279);
nor U11295 (N_11295,N_10577,N_10512);
xnor U11296 (N_11296,N_10372,N_10203);
nand U11297 (N_11297,N_10604,N_10079);
and U11298 (N_11298,N_10063,N_10888);
and U11299 (N_11299,N_10155,N_10923);
nand U11300 (N_11300,N_10761,N_10029);
nor U11301 (N_11301,N_10218,N_10657);
xnor U11302 (N_11302,N_10554,N_10214);
and U11303 (N_11303,N_10533,N_10081);
nor U11304 (N_11304,N_10714,N_10112);
and U11305 (N_11305,N_10064,N_10269);
nor U11306 (N_11306,N_10937,N_10687);
or U11307 (N_11307,N_10666,N_10543);
nor U11308 (N_11308,N_10558,N_10080);
nand U11309 (N_11309,N_10734,N_10088);
nor U11310 (N_11310,N_10224,N_10562);
nand U11311 (N_11311,N_10612,N_10012);
nor U11312 (N_11312,N_10690,N_10060);
xor U11313 (N_11313,N_10323,N_10270);
nor U11314 (N_11314,N_10871,N_10301);
and U11315 (N_11315,N_10147,N_10023);
nor U11316 (N_11316,N_10071,N_10066);
xnor U11317 (N_11317,N_10705,N_10583);
xnor U11318 (N_11318,N_10608,N_10999);
nand U11319 (N_11319,N_10882,N_10473);
and U11320 (N_11320,N_10077,N_10504);
nand U11321 (N_11321,N_10589,N_10411);
and U11322 (N_11322,N_10401,N_10349);
nor U11323 (N_11323,N_10691,N_10663);
nand U11324 (N_11324,N_10364,N_10377);
and U11325 (N_11325,N_10444,N_10004);
and U11326 (N_11326,N_10668,N_10161);
and U11327 (N_11327,N_10637,N_10107);
nand U11328 (N_11328,N_10282,N_10405);
nand U11329 (N_11329,N_10259,N_10162);
or U11330 (N_11330,N_10333,N_10946);
and U11331 (N_11331,N_10902,N_10748);
nand U11332 (N_11332,N_10750,N_10409);
or U11333 (N_11333,N_10312,N_10538);
nand U11334 (N_11334,N_10967,N_10560);
nor U11335 (N_11335,N_10959,N_10649);
or U11336 (N_11336,N_10234,N_10365);
or U11337 (N_11337,N_10617,N_10422);
nor U11338 (N_11338,N_10084,N_10320);
nor U11339 (N_11339,N_10989,N_10246);
nand U11340 (N_11340,N_10322,N_10470);
or U11341 (N_11341,N_10150,N_10756);
nor U11342 (N_11342,N_10801,N_10555);
xor U11343 (N_11343,N_10896,N_10961);
and U11344 (N_11344,N_10985,N_10744);
or U11345 (N_11345,N_10907,N_10457);
nand U11346 (N_11346,N_10743,N_10704);
nor U11347 (N_11347,N_10164,N_10140);
and U11348 (N_11348,N_10726,N_10284);
nor U11349 (N_11349,N_10105,N_10139);
and U11350 (N_11350,N_10406,N_10678);
xor U11351 (N_11351,N_10340,N_10969);
or U11352 (N_11352,N_10453,N_10367);
and U11353 (N_11353,N_10938,N_10595);
nor U11354 (N_11354,N_10170,N_10928);
xnor U11355 (N_11355,N_10843,N_10775);
nor U11356 (N_11356,N_10515,N_10215);
xor U11357 (N_11357,N_10784,N_10553);
nand U11358 (N_11358,N_10430,N_10459);
and U11359 (N_11359,N_10329,N_10658);
xor U11360 (N_11360,N_10036,N_10772);
nor U11361 (N_11361,N_10239,N_10684);
or U11362 (N_11362,N_10780,N_10518);
and U11363 (N_11363,N_10166,N_10404);
or U11364 (N_11364,N_10040,N_10338);
or U11365 (N_11365,N_10156,N_10628);
or U11366 (N_11366,N_10494,N_10693);
xor U11367 (N_11367,N_10572,N_10376);
xnor U11368 (N_11368,N_10350,N_10471);
nand U11369 (N_11369,N_10142,N_10842);
xor U11370 (N_11370,N_10712,N_10770);
or U11371 (N_11371,N_10776,N_10341);
nor U11372 (N_11372,N_10383,N_10794);
xor U11373 (N_11373,N_10958,N_10679);
nor U11374 (N_11374,N_10895,N_10531);
nor U11375 (N_11375,N_10021,N_10343);
and U11376 (N_11376,N_10905,N_10517);
or U11377 (N_11377,N_10075,N_10118);
nand U11378 (N_11378,N_10606,N_10363);
xnor U11379 (N_11379,N_10771,N_10009);
nand U11380 (N_11380,N_10630,N_10387);
xor U11381 (N_11381,N_10047,N_10392);
and U11382 (N_11382,N_10716,N_10765);
xnor U11383 (N_11383,N_10416,N_10450);
and U11384 (N_11384,N_10636,N_10437);
nand U11385 (N_11385,N_10209,N_10766);
nor U11386 (N_11386,N_10680,N_10722);
and U11387 (N_11387,N_10874,N_10352);
nor U11388 (N_11388,N_10461,N_10317);
nor U11389 (N_11389,N_10883,N_10137);
xnor U11390 (N_11390,N_10120,N_10539);
xor U11391 (N_11391,N_10039,N_10812);
nor U11392 (N_11392,N_10789,N_10255);
and U11393 (N_11393,N_10646,N_10724);
nor U11394 (N_11394,N_10316,N_10710);
or U11395 (N_11395,N_10370,N_10268);
nor U11396 (N_11396,N_10626,N_10994);
nand U11397 (N_11397,N_10160,N_10642);
nor U11398 (N_11398,N_10428,N_10508);
and U11399 (N_11399,N_10382,N_10523);
and U11400 (N_11400,N_10848,N_10840);
or U11401 (N_11401,N_10581,N_10569);
xor U11402 (N_11402,N_10737,N_10845);
nand U11403 (N_11403,N_10396,N_10757);
nor U11404 (N_11404,N_10243,N_10049);
and U11405 (N_11405,N_10468,N_10903);
nand U11406 (N_11406,N_10584,N_10527);
and U11407 (N_11407,N_10616,N_10731);
nor U11408 (N_11408,N_10173,N_10865);
or U11409 (N_11409,N_10591,N_10831);
nor U11410 (N_11410,N_10565,N_10828);
or U11411 (N_11411,N_10719,N_10347);
nor U11412 (N_11412,N_10391,N_10424);
and U11413 (N_11413,N_10385,N_10962);
nor U11414 (N_11414,N_10861,N_10953);
xnor U11415 (N_11415,N_10762,N_10286);
nor U11416 (N_11416,N_10927,N_10746);
nor U11417 (N_11417,N_10355,N_10732);
and U11418 (N_11418,N_10904,N_10031);
or U11419 (N_11419,N_10520,N_10248);
or U11420 (N_11420,N_10986,N_10791);
or U11421 (N_11421,N_10764,N_10123);
nor U11422 (N_11422,N_10258,N_10532);
xor U11423 (N_11423,N_10417,N_10335);
nor U11424 (N_11424,N_10635,N_10818);
and U11425 (N_11425,N_10909,N_10133);
nand U11426 (N_11426,N_10957,N_10298);
or U11427 (N_11427,N_10393,N_10272);
or U11428 (N_11428,N_10511,N_10917);
xnor U11429 (N_11429,N_10020,N_10125);
nand U11430 (N_11430,N_10158,N_10097);
nand U11431 (N_11431,N_10134,N_10738);
and U11432 (N_11432,N_10885,N_10250);
xor U11433 (N_11433,N_10596,N_10019);
xor U11434 (N_11434,N_10501,N_10521);
nand U11435 (N_11435,N_10477,N_10919);
or U11436 (N_11436,N_10920,N_10758);
nor U11437 (N_11437,N_10227,N_10135);
and U11438 (N_11438,N_10220,N_10242);
nor U11439 (N_11439,N_10685,N_10102);
or U11440 (N_11440,N_10467,N_10281);
nand U11441 (N_11441,N_10607,N_10585);
nand U11442 (N_11442,N_10264,N_10198);
nand U11443 (N_11443,N_10174,N_10643);
nand U11444 (N_11444,N_10415,N_10670);
xor U11445 (N_11445,N_10790,N_10886);
or U11446 (N_11446,N_10800,N_10141);
nor U11447 (N_11447,N_10507,N_10733);
and U11448 (N_11448,N_10366,N_10056);
or U11449 (N_11449,N_10375,N_10571);
nand U11450 (N_11450,N_10201,N_10977);
xnor U11451 (N_11451,N_10496,N_10254);
nand U11452 (N_11452,N_10359,N_10922);
xnor U11453 (N_11453,N_10486,N_10823);
or U11454 (N_11454,N_10172,N_10257);
xor U11455 (N_11455,N_10544,N_10998);
xor U11456 (N_11456,N_10605,N_10072);
or U11457 (N_11457,N_10197,N_10390);
xnor U11458 (N_11458,N_10165,N_10204);
or U11459 (N_11459,N_10240,N_10472);
nor U11460 (N_11460,N_10191,N_10362);
xor U11461 (N_11461,N_10096,N_10751);
and U11462 (N_11462,N_10436,N_10427);
nor U11463 (N_11463,N_10419,N_10890);
and U11464 (N_11464,N_10829,N_10694);
or U11465 (N_11465,N_10892,N_10803);
and U11466 (N_11466,N_10881,N_10564);
nor U11467 (N_11467,N_10353,N_10490);
xnor U11468 (N_11468,N_10285,N_10027);
or U11469 (N_11469,N_10041,N_10193);
xnor U11470 (N_11470,N_10230,N_10144);
xnor U11471 (N_11471,N_10530,N_10631);
nor U11472 (N_11472,N_10499,N_10394);
nor U11473 (N_11473,N_10971,N_10346);
and U11474 (N_11474,N_10745,N_10217);
nor U11475 (N_11475,N_10984,N_10802);
and U11476 (N_11476,N_10549,N_10002);
and U11477 (N_11477,N_10132,N_10110);
nand U11478 (N_11478,N_10065,N_10489);
xnor U11479 (N_11479,N_10777,N_10462);
nand U11480 (N_11480,N_10622,N_10324);
nand U11481 (N_11481,N_10769,N_10185);
nor U11482 (N_11482,N_10386,N_10309);
xor U11483 (N_11483,N_10598,N_10559);
and U11484 (N_11484,N_10295,N_10536);
and U11485 (N_11485,N_10213,N_10028);
xor U11486 (N_11486,N_10438,N_10754);
xor U11487 (N_11487,N_10186,N_10249);
and U11488 (N_11488,N_10537,N_10650);
nor U11489 (N_11489,N_10798,N_10825);
or U11490 (N_11490,N_10302,N_10182);
and U11491 (N_11491,N_10148,N_10157);
nand U11492 (N_11492,N_10008,N_10855);
or U11493 (N_11493,N_10785,N_10187);
nand U11494 (N_11494,N_10408,N_10397);
nand U11495 (N_11495,N_10940,N_10615);
or U11496 (N_11496,N_10497,N_10026);
nand U11497 (N_11497,N_10116,N_10076);
nand U11498 (N_11498,N_10127,N_10659);
and U11499 (N_11499,N_10334,N_10276);
or U11500 (N_11500,N_10037,N_10600);
nor U11501 (N_11501,N_10318,N_10974);
nor U11502 (N_11502,N_10501,N_10981);
or U11503 (N_11503,N_10117,N_10003);
and U11504 (N_11504,N_10331,N_10951);
nand U11505 (N_11505,N_10628,N_10670);
nand U11506 (N_11506,N_10947,N_10433);
and U11507 (N_11507,N_10250,N_10208);
nor U11508 (N_11508,N_10889,N_10394);
nand U11509 (N_11509,N_10088,N_10184);
and U11510 (N_11510,N_10522,N_10290);
nor U11511 (N_11511,N_10248,N_10668);
nand U11512 (N_11512,N_10792,N_10456);
xor U11513 (N_11513,N_10742,N_10839);
nor U11514 (N_11514,N_10800,N_10466);
and U11515 (N_11515,N_10871,N_10575);
or U11516 (N_11516,N_10311,N_10619);
xor U11517 (N_11517,N_10697,N_10627);
nand U11518 (N_11518,N_10311,N_10106);
nor U11519 (N_11519,N_10415,N_10442);
xnor U11520 (N_11520,N_10589,N_10744);
and U11521 (N_11521,N_10644,N_10514);
nand U11522 (N_11522,N_10211,N_10477);
and U11523 (N_11523,N_10603,N_10934);
xnor U11524 (N_11524,N_10126,N_10866);
xor U11525 (N_11525,N_10437,N_10774);
nor U11526 (N_11526,N_10479,N_10367);
or U11527 (N_11527,N_10345,N_10849);
nor U11528 (N_11528,N_10567,N_10563);
nor U11529 (N_11529,N_10043,N_10082);
xor U11530 (N_11530,N_10143,N_10106);
or U11531 (N_11531,N_10083,N_10417);
nor U11532 (N_11532,N_10933,N_10376);
and U11533 (N_11533,N_10614,N_10401);
or U11534 (N_11534,N_10106,N_10253);
nand U11535 (N_11535,N_10207,N_10746);
or U11536 (N_11536,N_10936,N_10907);
xor U11537 (N_11537,N_10673,N_10549);
nand U11538 (N_11538,N_10688,N_10768);
xnor U11539 (N_11539,N_10344,N_10708);
nand U11540 (N_11540,N_10279,N_10110);
nor U11541 (N_11541,N_10011,N_10410);
xor U11542 (N_11542,N_10928,N_10162);
and U11543 (N_11543,N_10229,N_10370);
nand U11544 (N_11544,N_10648,N_10335);
xnor U11545 (N_11545,N_10950,N_10126);
nand U11546 (N_11546,N_10306,N_10045);
nand U11547 (N_11547,N_10870,N_10524);
xnor U11548 (N_11548,N_10699,N_10512);
or U11549 (N_11549,N_10471,N_10248);
and U11550 (N_11550,N_10870,N_10634);
and U11551 (N_11551,N_10085,N_10788);
xor U11552 (N_11552,N_10497,N_10893);
nor U11553 (N_11553,N_10344,N_10144);
and U11554 (N_11554,N_10638,N_10521);
nor U11555 (N_11555,N_10221,N_10295);
and U11556 (N_11556,N_10461,N_10580);
xnor U11557 (N_11557,N_10055,N_10453);
and U11558 (N_11558,N_10465,N_10480);
nor U11559 (N_11559,N_10035,N_10393);
xor U11560 (N_11560,N_10004,N_10761);
and U11561 (N_11561,N_10747,N_10297);
nor U11562 (N_11562,N_10458,N_10161);
xor U11563 (N_11563,N_10097,N_10010);
nand U11564 (N_11564,N_10085,N_10509);
xor U11565 (N_11565,N_10620,N_10181);
nor U11566 (N_11566,N_10304,N_10787);
xor U11567 (N_11567,N_10921,N_10943);
or U11568 (N_11568,N_10196,N_10638);
or U11569 (N_11569,N_10839,N_10279);
or U11570 (N_11570,N_10721,N_10209);
nand U11571 (N_11571,N_10187,N_10138);
or U11572 (N_11572,N_10784,N_10418);
nor U11573 (N_11573,N_10544,N_10928);
or U11574 (N_11574,N_10256,N_10022);
nand U11575 (N_11575,N_10973,N_10233);
nand U11576 (N_11576,N_10892,N_10347);
and U11577 (N_11577,N_10995,N_10867);
xnor U11578 (N_11578,N_10601,N_10133);
nor U11579 (N_11579,N_10958,N_10995);
or U11580 (N_11580,N_10310,N_10672);
nor U11581 (N_11581,N_10968,N_10333);
or U11582 (N_11582,N_10215,N_10339);
nand U11583 (N_11583,N_10351,N_10417);
xor U11584 (N_11584,N_10575,N_10226);
nor U11585 (N_11585,N_10426,N_10812);
and U11586 (N_11586,N_10995,N_10019);
and U11587 (N_11587,N_10457,N_10645);
or U11588 (N_11588,N_10517,N_10011);
xnor U11589 (N_11589,N_10766,N_10164);
nor U11590 (N_11590,N_10506,N_10581);
nor U11591 (N_11591,N_10181,N_10716);
nor U11592 (N_11592,N_10284,N_10061);
xnor U11593 (N_11593,N_10063,N_10862);
xnor U11594 (N_11594,N_10257,N_10054);
or U11595 (N_11595,N_10604,N_10369);
nor U11596 (N_11596,N_10991,N_10333);
nand U11597 (N_11597,N_10421,N_10799);
xor U11598 (N_11598,N_10559,N_10483);
nor U11599 (N_11599,N_10754,N_10379);
xnor U11600 (N_11600,N_10038,N_10952);
xnor U11601 (N_11601,N_10384,N_10519);
or U11602 (N_11602,N_10282,N_10098);
and U11603 (N_11603,N_10612,N_10277);
nor U11604 (N_11604,N_10860,N_10726);
nand U11605 (N_11605,N_10475,N_10193);
nand U11606 (N_11606,N_10831,N_10051);
nand U11607 (N_11607,N_10858,N_10982);
xor U11608 (N_11608,N_10595,N_10721);
xor U11609 (N_11609,N_10770,N_10274);
or U11610 (N_11610,N_10342,N_10524);
or U11611 (N_11611,N_10886,N_10309);
nand U11612 (N_11612,N_10304,N_10292);
and U11613 (N_11613,N_10994,N_10410);
nor U11614 (N_11614,N_10879,N_10455);
or U11615 (N_11615,N_10168,N_10181);
xnor U11616 (N_11616,N_10462,N_10693);
or U11617 (N_11617,N_10957,N_10653);
nand U11618 (N_11618,N_10300,N_10636);
nor U11619 (N_11619,N_10189,N_10176);
xnor U11620 (N_11620,N_10551,N_10274);
or U11621 (N_11621,N_10202,N_10528);
nor U11622 (N_11622,N_10046,N_10755);
nor U11623 (N_11623,N_10195,N_10189);
nor U11624 (N_11624,N_10973,N_10920);
nand U11625 (N_11625,N_10164,N_10154);
and U11626 (N_11626,N_10898,N_10093);
xnor U11627 (N_11627,N_10777,N_10004);
nor U11628 (N_11628,N_10229,N_10608);
nand U11629 (N_11629,N_10322,N_10894);
and U11630 (N_11630,N_10423,N_10872);
nor U11631 (N_11631,N_10339,N_10663);
nand U11632 (N_11632,N_10861,N_10800);
xnor U11633 (N_11633,N_10194,N_10400);
xor U11634 (N_11634,N_10953,N_10359);
xor U11635 (N_11635,N_10472,N_10060);
xnor U11636 (N_11636,N_10356,N_10725);
nand U11637 (N_11637,N_10185,N_10286);
nand U11638 (N_11638,N_10750,N_10762);
or U11639 (N_11639,N_10977,N_10726);
nand U11640 (N_11640,N_10740,N_10497);
nor U11641 (N_11641,N_10541,N_10517);
xnor U11642 (N_11642,N_10221,N_10868);
nand U11643 (N_11643,N_10686,N_10354);
nor U11644 (N_11644,N_10788,N_10708);
nor U11645 (N_11645,N_10028,N_10467);
nand U11646 (N_11646,N_10822,N_10932);
or U11647 (N_11647,N_10355,N_10688);
and U11648 (N_11648,N_10561,N_10199);
nand U11649 (N_11649,N_10160,N_10263);
xnor U11650 (N_11650,N_10937,N_10903);
or U11651 (N_11651,N_10098,N_10763);
nor U11652 (N_11652,N_10188,N_10134);
or U11653 (N_11653,N_10262,N_10780);
or U11654 (N_11654,N_10101,N_10696);
and U11655 (N_11655,N_10159,N_10034);
or U11656 (N_11656,N_10161,N_10057);
or U11657 (N_11657,N_10717,N_10289);
nor U11658 (N_11658,N_10850,N_10915);
xor U11659 (N_11659,N_10436,N_10023);
or U11660 (N_11660,N_10349,N_10559);
and U11661 (N_11661,N_10343,N_10947);
nand U11662 (N_11662,N_10530,N_10163);
xor U11663 (N_11663,N_10321,N_10722);
xor U11664 (N_11664,N_10473,N_10344);
xor U11665 (N_11665,N_10126,N_10430);
xnor U11666 (N_11666,N_10425,N_10484);
or U11667 (N_11667,N_10729,N_10873);
and U11668 (N_11668,N_10260,N_10412);
xnor U11669 (N_11669,N_10185,N_10345);
or U11670 (N_11670,N_10030,N_10715);
nor U11671 (N_11671,N_10661,N_10548);
or U11672 (N_11672,N_10498,N_10971);
nand U11673 (N_11673,N_10467,N_10430);
nand U11674 (N_11674,N_10584,N_10482);
nor U11675 (N_11675,N_10480,N_10748);
nor U11676 (N_11676,N_10756,N_10427);
xor U11677 (N_11677,N_10327,N_10565);
nor U11678 (N_11678,N_10879,N_10161);
xnor U11679 (N_11679,N_10145,N_10778);
nor U11680 (N_11680,N_10114,N_10145);
or U11681 (N_11681,N_10451,N_10720);
and U11682 (N_11682,N_10084,N_10453);
xor U11683 (N_11683,N_10653,N_10171);
xor U11684 (N_11684,N_10481,N_10886);
nand U11685 (N_11685,N_10893,N_10143);
or U11686 (N_11686,N_10858,N_10325);
nand U11687 (N_11687,N_10873,N_10616);
and U11688 (N_11688,N_10063,N_10690);
xor U11689 (N_11689,N_10087,N_10231);
nand U11690 (N_11690,N_10194,N_10423);
or U11691 (N_11691,N_10151,N_10327);
xor U11692 (N_11692,N_10251,N_10954);
nand U11693 (N_11693,N_10718,N_10468);
or U11694 (N_11694,N_10032,N_10968);
xor U11695 (N_11695,N_10904,N_10327);
xnor U11696 (N_11696,N_10935,N_10921);
xnor U11697 (N_11697,N_10433,N_10426);
xnor U11698 (N_11698,N_10344,N_10335);
nor U11699 (N_11699,N_10623,N_10425);
and U11700 (N_11700,N_10405,N_10045);
nor U11701 (N_11701,N_10535,N_10221);
nand U11702 (N_11702,N_10274,N_10750);
nor U11703 (N_11703,N_10522,N_10971);
nand U11704 (N_11704,N_10307,N_10861);
or U11705 (N_11705,N_10111,N_10739);
xnor U11706 (N_11706,N_10577,N_10509);
and U11707 (N_11707,N_10371,N_10874);
nand U11708 (N_11708,N_10470,N_10123);
nand U11709 (N_11709,N_10095,N_10937);
nand U11710 (N_11710,N_10240,N_10138);
nor U11711 (N_11711,N_10968,N_10245);
nand U11712 (N_11712,N_10888,N_10225);
or U11713 (N_11713,N_10054,N_10109);
or U11714 (N_11714,N_10983,N_10735);
nor U11715 (N_11715,N_10393,N_10320);
nand U11716 (N_11716,N_10406,N_10378);
xor U11717 (N_11717,N_10511,N_10323);
and U11718 (N_11718,N_10833,N_10954);
and U11719 (N_11719,N_10848,N_10945);
and U11720 (N_11720,N_10017,N_10955);
nor U11721 (N_11721,N_10571,N_10676);
xor U11722 (N_11722,N_10358,N_10429);
nand U11723 (N_11723,N_10624,N_10992);
xor U11724 (N_11724,N_10829,N_10921);
xor U11725 (N_11725,N_10276,N_10630);
nand U11726 (N_11726,N_10593,N_10736);
nand U11727 (N_11727,N_10253,N_10332);
and U11728 (N_11728,N_10805,N_10169);
nor U11729 (N_11729,N_10608,N_10495);
or U11730 (N_11730,N_10713,N_10215);
and U11731 (N_11731,N_10649,N_10910);
nand U11732 (N_11732,N_10348,N_10027);
or U11733 (N_11733,N_10484,N_10006);
nand U11734 (N_11734,N_10008,N_10690);
nor U11735 (N_11735,N_10800,N_10873);
or U11736 (N_11736,N_10108,N_10950);
xnor U11737 (N_11737,N_10960,N_10257);
or U11738 (N_11738,N_10289,N_10389);
nand U11739 (N_11739,N_10269,N_10763);
and U11740 (N_11740,N_10665,N_10591);
or U11741 (N_11741,N_10170,N_10642);
nor U11742 (N_11742,N_10126,N_10104);
or U11743 (N_11743,N_10762,N_10401);
nand U11744 (N_11744,N_10458,N_10986);
nand U11745 (N_11745,N_10014,N_10825);
xnor U11746 (N_11746,N_10130,N_10094);
or U11747 (N_11747,N_10561,N_10296);
nor U11748 (N_11748,N_10248,N_10312);
xnor U11749 (N_11749,N_10052,N_10893);
or U11750 (N_11750,N_10795,N_10873);
nand U11751 (N_11751,N_10347,N_10169);
and U11752 (N_11752,N_10020,N_10024);
nor U11753 (N_11753,N_10745,N_10178);
and U11754 (N_11754,N_10358,N_10413);
xnor U11755 (N_11755,N_10796,N_10538);
or U11756 (N_11756,N_10827,N_10977);
xnor U11757 (N_11757,N_10583,N_10389);
nand U11758 (N_11758,N_10480,N_10894);
and U11759 (N_11759,N_10989,N_10954);
nand U11760 (N_11760,N_10886,N_10681);
nand U11761 (N_11761,N_10045,N_10443);
or U11762 (N_11762,N_10480,N_10504);
nor U11763 (N_11763,N_10836,N_10551);
xor U11764 (N_11764,N_10144,N_10957);
xor U11765 (N_11765,N_10653,N_10978);
nor U11766 (N_11766,N_10479,N_10026);
nor U11767 (N_11767,N_10727,N_10275);
nor U11768 (N_11768,N_10180,N_10298);
or U11769 (N_11769,N_10785,N_10317);
nand U11770 (N_11770,N_10985,N_10125);
xnor U11771 (N_11771,N_10085,N_10540);
xor U11772 (N_11772,N_10381,N_10966);
xnor U11773 (N_11773,N_10220,N_10707);
nor U11774 (N_11774,N_10311,N_10376);
nand U11775 (N_11775,N_10868,N_10445);
or U11776 (N_11776,N_10355,N_10377);
xor U11777 (N_11777,N_10600,N_10462);
and U11778 (N_11778,N_10040,N_10968);
and U11779 (N_11779,N_10650,N_10694);
and U11780 (N_11780,N_10075,N_10202);
xor U11781 (N_11781,N_10623,N_10656);
xor U11782 (N_11782,N_10567,N_10754);
xnor U11783 (N_11783,N_10996,N_10746);
or U11784 (N_11784,N_10705,N_10184);
and U11785 (N_11785,N_10506,N_10573);
nand U11786 (N_11786,N_10224,N_10790);
and U11787 (N_11787,N_10319,N_10117);
nor U11788 (N_11788,N_10271,N_10257);
nor U11789 (N_11789,N_10781,N_10115);
and U11790 (N_11790,N_10186,N_10174);
and U11791 (N_11791,N_10693,N_10595);
nor U11792 (N_11792,N_10760,N_10532);
and U11793 (N_11793,N_10951,N_10206);
xnor U11794 (N_11794,N_10364,N_10079);
or U11795 (N_11795,N_10266,N_10896);
nand U11796 (N_11796,N_10282,N_10352);
or U11797 (N_11797,N_10280,N_10500);
and U11798 (N_11798,N_10999,N_10340);
xnor U11799 (N_11799,N_10732,N_10116);
nand U11800 (N_11800,N_10574,N_10709);
xnor U11801 (N_11801,N_10579,N_10077);
or U11802 (N_11802,N_10394,N_10299);
nor U11803 (N_11803,N_10529,N_10162);
xnor U11804 (N_11804,N_10736,N_10709);
nand U11805 (N_11805,N_10281,N_10225);
and U11806 (N_11806,N_10658,N_10351);
xor U11807 (N_11807,N_10143,N_10300);
xnor U11808 (N_11808,N_10691,N_10348);
nand U11809 (N_11809,N_10456,N_10614);
or U11810 (N_11810,N_10446,N_10011);
nand U11811 (N_11811,N_10090,N_10896);
or U11812 (N_11812,N_10108,N_10426);
xor U11813 (N_11813,N_10277,N_10806);
and U11814 (N_11814,N_10430,N_10150);
and U11815 (N_11815,N_10289,N_10810);
or U11816 (N_11816,N_10344,N_10017);
or U11817 (N_11817,N_10591,N_10662);
xnor U11818 (N_11818,N_10117,N_10525);
and U11819 (N_11819,N_10851,N_10814);
nand U11820 (N_11820,N_10529,N_10174);
nor U11821 (N_11821,N_10807,N_10530);
xor U11822 (N_11822,N_10382,N_10794);
nand U11823 (N_11823,N_10022,N_10674);
or U11824 (N_11824,N_10692,N_10036);
and U11825 (N_11825,N_10168,N_10747);
nand U11826 (N_11826,N_10198,N_10541);
nor U11827 (N_11827,N_10960,N_10735);
nand U11828 (N_11828,N_10079,N_10575);
and U11829 (N_11829,N_10947,N_10129);
nor U11830 (N_11830,N_10397,N_10624);
nand U11831 (N_11831,N_10021,N_10347);
or U11832 (N_11832,N_10767,N_10646);
and U11833 (N_11833,N_10716,N_10666);
xnor U11834 (N_11834,N_10294,N_10645);
or U11835 (N_11835,N_10438,N_10386);
or U11836 (N_11836,N_10580,N_10694);
nor U11837 (N_11837,N_10923,N_10526);
or U11838 (N_11838,N_10126,N_10407);
xor U11839 (N_11839,N_10573,N_10014);
nor U11840 (N_11840,N_10426,N_10353);
xnor U11841 (N_11841,N_10807,N_10390);
nor U11842 (N_11842,N_10186,N_10576);
nand U11843 (N_11843,N_10599,N_10338);
nand U11844 (N_11844,N_10711,N_10745);
nand U11845 (N_11845,N_10575,N_10291);
and U11846 (N_11846,N_10532,N_10865);
xor U11847 (N_11847,N_10271,N_10730);
or U11848 (N_11848,N_10026,N_10747);
nor U11849 (N_11849,N_10358,N_10327);
nand U11850 (N_11850,N_10544,N_10683);
and U11851 (N_11851,N_10540,N_10435);
nor U11852 (N_11852,N_10292,N_10248);
nand U11853 (N_11853,N_10156,N_10527);
or U11854 (N_11854,N_10243,N_10063);
nor U11855 (N_11855,N_10810,N_10340);
and U11856 (N_11856,N_10324,N_10690);
and U11857 (N_11857,N_10062,N_10465);
nor U11858 (N_11858,N_10255,N_10377);
nand U11859 (N_11859,N_10502,N_10887);
or U11860 (N_11860,N_10474,N_10688);
nor U11861 (N_11861,N_10410,N_10968);
or U11862 (N_11862,N_10509,N_10825);
or U11863 (N_11863,N_10355,N_10694);
nor U11864 (N_11864,N_10670,N_10013);
and U11865 (N_11865,N_10616,N_10424);
or U11866 (N_11866,N_10934,N_10564);
xor U11867 (N_11867,N_10021,N_10671);
or U11868 (N_11868,N_10995,N_10285);
xnor U11869 (N_11869,N_10160,N_10202);
xor U11870 (N_11870,N_10388,N_10137);
and U11871 (N_11871,N_10149,N_10620);
nor U11872 (N_11872,N_10011,N_10258);
and U11873 (N_11873,N_10908,N_10795);
or U11874 (N_11874,N_10058,N_10488);
and U11875 (N_11875,N_10960,N_10458);
nand U11876 (N_11876,N_10393,N_10979);
xor U11877 (N_11877,N_10698,N_10018);
or U11878 (N_11878,N_10179,N_10547);
or U11879 (N_11879,N_10083,N_10759);
nand U11880 (N_11880,N_10212,N_10902);
nor U11881 (N_11881,N_10351,N_10743);
or U11882 (N_11882,N_10370,N_10747);
xnor U11883 (N_11883,N_10102,N_10889);
nor U11884 (N_11884,N_10878,N_10141);
xor U11885 (N_11885,N_10485,N_10059);
xor U11886 (N_11886,N_10038,N_10456);
and U11887 (N_11887,N_10863,N_10892);
or U11888 (N_11888,N_10743,N_10931);
and U11889 (N_11889,N_10008,N_10573);
nor U11890 (N_11890,N_10405,N_10680);
and U11891 (N_11891,N_10107,N_10019);
or U11892 (N_11892,N_10942,N_10946);
and U11893 (N_11893,N_10393,N_10940);
or U11894 (N_11894,N_10796,N_10536);
nor U11895 (N_11895,N_10084,N_10893);
xor U11896 (N_11896,N_10287,N_10359);
or U11897 (N_11897,N_10580,N_10316);
and U11898 (N_11898,N_10660,N_10829);
xnor U11899 (N_11899,N_10509,N_10499);
nor U11900 (N_11900,N_10441,N_10127);
nor U11901 (N_11901,N_10442,N_10241);
xnor U11902 (N_11902,N_10936,N_10334);
nand U11903 (N_11903,N_10308,N_10121);
or U11904 (N_11904,N_10612,N_10854);
and U11905 (N_11905,N_10541,N_10697);
nand U11906 (N_11906,N_10711,N_10314);
and U11907 (N_11907,N_10246,N_10440);
and U11908 (N_11908,N_10785,N_10894);
and U11909 (N_11909,N_10179,N_10777);
or U11910 (N_11910,N_10363,N_10144);
and U11911 (N_11911,N_10340,N_10974);
xor U11912 (N_11912,N_10277,N_10629);
xor U11913 (N_11913,N_10071,N_10737);
nor U11914 (N_11914,N_10134,N_10603);
nor U11915 (N_11915,N_10466,N_10975);
xnor U11916 (N_11916,N_10008,N_10753);
xor U11917 (N_11917,N_10409,N_10752);
and U11918 (N_11918,N_10424,N_10164);
and U11919 (N_11919,N_10590,N_10958);
xor U11920 (N_11920,N_10830,N_10507);
nor U11921 (N_11921,N_10245,N_10763);
nor U11922 (N_11922,N_10479,N_10001);
nand U11923 (N_11923,N_10147,N_10551);
nor U11924 (N_11924,N_10715,N_10320);
xnor U11925 (N_11925,N_10069,N_10222);
nand U11926 (N_11926,N_10307,N_10947);
or U11927 (N_11927,N_10305,N_10460);
and U11928 (N_11928,N_10399,N_10326);
xor U11929 (N_11929,N_10820,N_10822);
xor U11930 (N_11930,N_10869,N_10243);
and U11931 (N_11931,N_10452,N_10821);
or U11932 (N_11932,N_10324,N_10559);
nand U11933 (N_11933,N_10440,N_10268);
xor U11934 (N_11934,N_10944,N_10412);
nand U11935 (N_11935,N_10040,N_10203);
nor U11936 (N_11936,N_10709,N_10698);
xnor U11937 (N_11937,N_10692,N_10856);
nor U11938 (N_11938,N_10264,N_10459);
nor U11939 (N_11939,N_10048,N_10730);
xnor U11940 (N_11940,N_10932,N_10623);
nor U11941 (N_11941,N_10483,N_10713);
nand U11942 (N_11942,N_10337,N_10143);
xnor U11943 (N_11943,N_10289,N_10071);
and U11944 (N_11944,N_10572,N_10839);
xnor U11945 (N_11945,N_10026,N_10817);
or U11946 (N_11946,N_10619,N_10120);
and U11947 (N_11947,N_10394,N_10890);
xnor U11948 (N_11948,N_10897,N_10034);
nand U11949 (N_11949,N_10819,N_10745);
and U11950 (N_11950,N_10178,N_10342);
nand U11951 (N_11951,N_10467,N_10595);
xor U11952 (N_11952,N_10704,N_10106);
or U11953 (N_11953,N_10159,N_10119);
or U11954 (N_11954,N_10194,N_10629);
and U11955 (N_11955,N_10031,N_10533);
or U11956 (N_11956,N_10542,N_10782);
nor U11957 (N_11957,N_10383,N_10434);
or U11958 (N_11958,N_10752,N_10118);
and U11959 (N_11959,N_10368,N_10200);
or U11960 (N_11960,N_10529,N_10957);
and U11961 (N_11961,N_10993,N_10972);
nor U11962 (N_11962,N_10299,N_10740);
and U11963 (N_11963,N_10067,N_10579);
and U11964 (N_11964,N_10024,N_10534);
nor U11965 (N_11965,N_10893,N_10871);
nor U11966 (N_11966,N_10964,N_10686);
or U11967 (N_11967,N_10605,N_10640);
or U11968 (N_11968,N_10473,N_10987);
xor U11969 (N_11969,N_10372,N_10494);
and U11970 (N_11970,N_10677,N_10711);
nor U11971 (N_11971,N_10757,N_10335);
xor U11972 (N_11972,N_10230,N_10888);
nor U11973 (N_11973,N_10916,N_10759);
xnor U11974 (N_11974,N_10411,N_10066);
nor U11975 (N_11975,N_10202,N_10558);
nor U11976 (N_11976,N_10341,N_10632);
nor U11977 (N_11977,N_10286,N_10757);
nor U11978 (N_11978,N_10716,N_10075);
nand U11979 (N_11979,N_10279,N_10702);
or U11980 (N_11980,N_10814,N_10395);
xor U11981 (N_11981,N_10029,N_10477);
xnor U11982 (N_11982,N_10896,N_10061);
nand U11983 (N_11983,N_10566,N_10388);
nor U11984 (N_11984,N_10871,N_10603);
nand U11985 (N_11985,N_10360,N_10206);
or U11986 (N_11986,N_10393,N_10382);
nor U11987 (N_11987,N_10079,N_10667);
or U11988 (N_11988,N_10409,N_10882);
nor U11989 (N_11989,N_10115,N_10773);
or U11990 (N_11990,N_10143,N_10931);
nor U11991 (N_11991,N_10559,N_10185);
xnor U11992 (N_11992,N_10603,N_10831);
xor U11993 (N_11993,N_10518,N_10693);
and U11994 (N_11994,N_10557,N_10636);
xnor U11995 (N_11995,N_10638,N_10553);
nor U11996 (N_11996,N_10398,N_10726);
nand U11997 (N_11997,N_10359,N_10745);
and U11998 (N_11998,N_10929,N_10826);
nor U11999 (N_11999,N_10013,N_10693);
xor U12000 (N_12000,N_11875,N_11501);
xor U12001 (N_12001,N_11723,N_11354);
or U12002 (N_12002,N_11164,N_11207);
and U12003 (N_12003,N_11768,N_11303);
nand U12004 (N_12004,N_11361,N_11512);
nand U12005 (N_12005,N_11738,N_11627);
or U12006 (N_12006,N_11706,N_11935);
nand U12007 (N_12007,N_11447,N_11986);
or U12008 (N_12008,N_11269,N_11165);
or U12009 (N_12009,N_11728,N_11541);
xor U12010 (N_12010,N_11286,N_11783);
or U12011 (N_12011,N_11774,N_11691);
xnor U12012 (N_12012,N_11929,N_11277);
or U12013 (N_12013,N_11034,N_11382);
or U12014 (N_12014,N_11786,N_11813);
xor U12015 (N_12015,N_11002,N_11422);
or U12016 (N_12016,N_11588,N_11614);
xor U12017 (N_12017,N_11886,N_11567);
and U12018 (N_12018,N_11654,N_11208);
nor U12019 (N_12019,N_11008,N_11259);
or U12020 (N_12020,N_11298,N_11520);
nand U12021 (N_12021,N_11709,N_11255);
nand U12022 (N_12022,N_11715,N_11579);
nand U12023 (N_12023,N_11630,N_11121);
nor U12024 (N_12024,N_11973,N_11992);
or U12025 (N_12025,N_11885,N_11092);
nor U12026 (N_12026,N_11054,N_11093);
nand U12027 (N_12027,N_11889,N_11392);
xor U12028 (N_12028,N_11249,N_11879);
or U12029 (N_12029,N_11534,N_11735);
and U12030 (N_12030,N_11631,N_11620);
xnor U12031 (N_12031,N_11272,N_11021);
or U12032 (N_12032,N_11946,N_11535);
and U12033 (N_12033,N_11261,N_11496);
nor U12034 (N_12034,N_11058,N_11724);
nor U12035 (N_12035,N_11937,N_11478);
xor U12036 (N_12036,N_11900,N_11116);
nand U12037 (N_12037,N_11721,N_11073);
nand U12038 (N_12038,N_11486,N_11551);
and U12039 (N_12039,N_11677,N_11803);
or U12040 (N_12040,N_11903,N_11055);
xor U12041 (N_12041,N_11802,N_11832);
nor U12042 (N_12042,N_11770,N_11711);
and U12043 (N_12043,N_11598,N_11377);
nand U12044 (N_12044,N_11350,N_11036);
or U12045 (N_12045,N_11862,N_11445);
nand U12046 (N_12046,N_11615,N_11483);
nand U12047 (N_12047,N_11555,N_11290);
nor U12048 (N_12048,N_11751,N_11934);
nor U12049 (N_12049,N_11911,N_11206);
or U12050 (N_12050,N_11909,N_11379);
xor U12051 (N_12051,N_11978,N_11046);
or U12052 (N_12052,N_11572,N_11237);
and U12053 (N_12053,N_11319,N_11893);
nand U12054 (N_12054,N_11729,N_11000);
and U12055 (N_12055,N_11312,N_11841);
xor U12056 (N_12056,N_11926,N_11650);
xor U12057 (N_12057,N_11473,N_11267);
nand U12058 (N_12058,N_11171,N_11367);
and U12059 (N_12059,N_11871,N_11749);
nor U12060 (N_12060,N_11175,N_11405);
xor U12061 (N_12061,N_11632,N_11053);
or U12062 (N_12062,N_11970,N_11480);
xnor U12063 (N_12063,N_11814,N_11087);
and U12064 (N_12064,N_11244,N_11562);
nor U12065 (N_12065,N_11215,N_11993);
xor U12066 (N_12066,N_11605,N_11221);
nand U12067 (N_12067,N_11084,N_11604);
or U12068 (N_12068,N_11157,N_11345);
nand U12069 (N_12069,N_11071,N_11094);
and U12070 (N_12070,N_11219,N_11047);
xor U12071 (N_12071,N_11842,N_11192);
xnor U12072 (N_12072,N_11669,N_11743);
and U12073 (N_12073,N_11883,N_11516);
nor U12074 (N_12074,N_11806,N_11626);
nand U12075 (N_12075,N_11080,N_11460);
or U12076 (N_12076,N_11759,N_11309);
nor U12077 (N_12077,N_11112,N_11590);
and U12078 (N_12078,N_11444,N_11853);
xnor U12079 (N_12079,N_11072,N_11891);
and U12080 (N_12080,N_11180,N_11438);
nor U12081 (N_12081,N_11097,N_11547);
nor U12082 (N_12082,N_11557,N_11141);
nand U12083 (N_12083,N_11417,N_11117);
xor U12084 (N_12084,N_11032,N_11421);
nor U12085 (N_12085,N_11115,N_11293);
xor U12086 (N_12086,N_11147,N_11525);
nand U12087 (N_12087,N_11229,N_11740);
xnor U12088 (N_12088,N_11355,N_11995);
nor U12089 (N_12089,N_11573,N_11754);
nor U12090 (N_12090,N_11936,N_11096);
xnor U12091 (N_12091,N_11051,N_11378);
xor U12092 (N_12092,N_11263,N_11914);
or U12093 (N_12093,N_11888,N_11402);
nand U12094 (N_12094,N_11454,N_11156);
or U12095 (N_12095,N_11228,N_11999);
or U12096 (N_12096,N_11837,N_11872);
and U12097 (N_12097,N_11758,N_11142);
xor U12098 (N_12098,N_11078,N_11281);
or U12099 (N_12099,N_11362,N_11578);
nand U12100 (N_12100,N_11430,N_11288);
nor U12101 (N_12101,N_11082,N_11426);
nor U12102 (N_12102,N_11060,N_11477);
or U12103 (N_12103,N_11482,N_11250);
and U12104 (N_12104,N_11152,N_11506);
nand U12105 (N_12105,N_11118,N_11081);
nand U12106 (N_12106,N_11897,N_11359);
or U12107 (N_12107,N_11710,N_11341);
and U12108 (N_12108,N_11596,N_11302);
and U12109 (N_12109,N_11539,N_11601);
or U12110 (N_12110,N_11540,N_11855);
and U12111 (N_12111,N_11182,N_11083);
nor U12112 (N_12112,N_11067,N_11725);
nand U12113 (N_12113,N_11518,N_11722);
and U12114 (N_12114,N_11038,N_11101);
nand U12115 (N_12115,N_11739,N_11380);
nor U12116 (N_12116,N_11705,N_11857);
nor U12117 (N_12117,N_11876,N_11693);
xor U12118 (N_12118,N_11128,N_11966);
and U12119 (N_12119,N_11890,N_11289);
and U12120 (N_12120,N_11401,N_11481);
xor U12121 (N_12121,N_11386,N_11592);
nand U12122 (N_12122,N_11335,N_11393);
nand U12123 (N_12123,N_11887,N_11780);
nand U12124 (N_12124,N_11894,N_11683);
nand U12125 (N_12125,N_11026,N_11695);
xnor U12126 (N_12126,N_11767,N_11665);
and U12127 (N_12127,N_11205,N_11103);
xnor U12128 (N_12128,N_11273,N_11543);
xnor U12129 (N_12129,N_11874,N_11292);
nand U12130 (N_12130,N_11381,N_11753);
or U12131 (N_12131,N_11530,N_11185);
and U12132 (N_12132,N_11119,N_11079);
nor U12133 (N_12133,N_11960,N_11594);
or U12134 (N_12134,N_11584,N_11406);
nand U12135 (N_12135,N_11622,N_11990);
nand U12136 (N_12136,N_11130,N_11550);
or U12137 (N_12137,N_11351,N_11016);
xor U12138 (N_12138,N_11004,N_11559);
and U12139 (N_12139,N_11574,N_11015);
nand U12140 (N_12140,N_11836,N_11629);
xnor U12141 (N_12141,N_11931,N_11279);
nor U12142 (N_12142,N_11098,N_11689);
nand U12143 (N_12143,N_11659,N_11232);
nor U12144 (N_12144,N_11265,N_11431);
nor U12145 (N_12145,N_11305,N_11007);
nand U12146 (N_12146,N_11258,N_11531);
nor U12147 (N_12147,N_11922,N_11253);
and U12148 (N_12148,N_11191,N_11333);
or U12149 (N_12149,N_11517,N_11176);
nor U12150 (N_12150,N_11927,N_11901);
or U12151 (N_12151,N_11413,N_11808);
nand U12152 (N_12152,N_11339,N_11734);
nor U12153 (N_12153,N_11148,N_11940);
or U12154 (N_12154,N_11399,N_11984);
and U12155 (N_12155,N_11792,N_11200);
nand U12156 (N_12156,N_11979,N_11954);
nor U12157 (N_12157,N_11581,N_11236);
or U12158 (N_12158,N_11301,N_11035);
and U12159 (N_12159,N_11409,N_11190);
and U12160 (N_12160,N_11314,N_11398);
xnor U12161 (N_12161,N_11343,N_11948);
or U12162 (N_12162,N_11595,N_11113);
or U12163 (N_12163,N_11839,N_11254);
and U12164 (N_12164,N_11349,N_11846);
nand U12165 (N_12165,N_11570,N_11070);
or U12166 (N_12166,N_11793,N_11671);
nor U12167 (N_12167,N_11168,N_11921);
nand U12168 (N_12168,N_11681,N_11275);
or U12169 (N_12169,N_11800,N_11025);
and U12170 (N_12170,N_11435,N_11688);
or U12171 (N_12171,N_11987,N_11144);
or U12172 (N_12172,N_11991,N_11684);
xor U12173 (N_12173,N_11642,N_11549);
or U12174 (N_12174,N_11829,N_11737);
nor U12175 (N_12175,N_11226,N_11854);
xnor U12176 (N_12176,N_11100,N_11657);
and U12177 (N_12177,N_11819,N_11612);
or U12178 (N_12178,N_11816,N_11235);
nand U12179 (N_12179,N_11238,N_11155);
xor U12180 (N_12180,N_11143,N_11220);
or U12181 (N_12181,N_11304,N_11068);
and U12182 (N_12182,N_11600,N_11805);
and U12183 (N_12183,N_11717,N_11162);
and U12184 (N_12184,N_11360,N_11436);
and U12185 (N_12185,N_11782,N_11781);
nand U12186 (N_12186,N_11744,N_11641);
nand U12187 (N_12187,N_11005,N_11346);
or U12188 (N_12188,N_11074,N_11713);
nand U12189 (N_12189,N_11509,N_11131);
xnor U12190 (N_12190,N_11432,N_11484);
and U12191 (N_12191,N_11603,N_11407);
nor U12192 (N_12192,N_11280,N_11469);
nor U12193 (N_12193,N_11583,N_11527);
nand U12194 (N_12194,N_11982,N_11702);
xor U12195 (N_12195,N_11917,N_11618);
nor U12196 (N_12196,N_11554,N_11965);
nand U12197 (N_12197,N_11291,N_11459);
and U12198 (N_12198,N_11560,N_11158);
nand U12199 (N_12199,N_11775,N_11045);
or U12200 (N_12200,N_11123,N_11964);
nor U12201 (N_12201,N_11989,N_11619);
xnor U12202 (N_12202,N_11248,N_11499);
or U12203 (N_12203,N_11427,N_11651);
and U12204 (N_12204,N_11497,N_11696);
and U12205 (N_12205,N_11831,N_11344);
and U12206 (N_12206,N_11804,N_11216);
nand U12207 (N_12207,N_11414,N_11838);
or U12208 (N_12208,N_11327,N_11048);
nor U12209 (N_12209,N_11122,N_11400);
xor U12210 (N_12210,N_11988,N_11944);
xor U12211 (N_12211,N_11183,N_11440);
nor U12212 (N_12212,N_11616,N_11779);
xor U12213 (N_12213,N_11593,N_11439);
nor U12214 (N_12214,N_11932,N_11765);
xor U12215 (N_12215,N_11376,N_11546);
nand U12216 (N_12216,N_11500,N_11334);
and U12217 (N_12217,N_11492,N_11633);
xnor U12218 (N_12218,N_11817,N_11680);
or U12219 (N_12219,N_11563,N_11467);
nor U12220 (N_12220,N_11468,N_11542);
or U12221 (N_12221,N_11332,N_11587);
and U12222 (N_12222,N_11336,N_11330);
or U12223 (N_12223,N_11938,N_11848);
and U12224 (N_12224,N_11840,N_11502);
nor U12225 (N_12225,N_11061,N_11971);
xnor U12226 (N_12226,N_11868,N_11154);
xor U12227 (N_12227,N_11858,N_11135);
xnor U12228 (N_12228,N_11247,N_11867);
nand U12229 (N_12229,N_11451,N_11340);
or U12230 (N_12230,N_11692,N_11924);
xnor U12231 (N_12231,N_11714,N_11095);
nor U12232 (N_12232,N_11959,N_11915);
xor U12233 (N_12233,N_11213,N_11251);
nor U12234 (N_12234,N_11752,N_11160);
nand U12235 (N_12235,N_11370,N_11403);
or U12236 (N_12236,N_11283,N_11167);
or U12237 (N_12237,N_11907,N_11690);
nand U12238 (N_12238,N_11150,N_11065);
nand U12239 (N_12239,N_11326,N_11733);
and U12240 (N_12240,N_11028,N_11703);
and U12241 (N_12241,N_11196,N_11151);
nor U12242 (N_12242,N_11834,N_11404);
xor U12243 (N_12243,N_11852,N_11953);
nor U12244 (N_12244,N_11621,N_11504);
and U12245 (N_12245,N_11697,N_11424);
and U12246 (N_12246,N_11957,N_11866);
or U12247 (N_12247,N_11342,N_11088);
nor U12248 (N_12248,N_11225,N_11296);
or U12249 (N_12249,N_11138,N_11371);
nand U12250 (N_12250,N_11287,N_11640);
nand U12251 (N_12251,N_11634,N_11773);
xnor U12252 (N_12252,N_11211,N_11745);
nand U12253 (N_12253,N_11085,N_11129);
and U12254 (N_12254,N_11318,N_11789);
nand U12255 (N_12255,N_11916,N_11170);
or U12256 (N_12256,N_11652,N_11495);
or U12257 (N_12257,N_11408,N_11240);
nand U12258 (N_12258,N_11799,N_11023);
or U12259 (N_12259,N_11218,N_11489);
or U12260 (N_12260,N_11090,N_11163);
nor U12261 (N_12261,N_11297,N_11052);
nor U12262 (N_12262,N_11491,N_11389);
nor U12263 (N_12263,N_11429,N_11599);
nand U12264 (N_12264,N_11976,N_11461);
and U12265 (N_12265,N_11707,N_11464);
nor U12266 (N_12266,N_11294,N_11124);
and U12267 (N_12267,N_11636,N_11214);
and U12268 (N_12268,N_11062,N_11474);
nor U12269 (N_12269,N_11637,N_11257);
xnor U12270 (N_12270,N_11266,N_11794);
and U12271 (N_12271,N_11983,N_11159);
xor U12272 (N_12272,N_11760,N_11647);
nand U12273 (N_12273,N_11284,N_11798);
nand U12274 (N_12274,N_11075,N_11796);
and U12275 (N_12275,N_11653,N_11013);
nor U12276 (N_12276,N_11508,N_11873);
nor U12277 (N_12277,N_11299,N_11086);
and U12278 (N_12278,N_11285,N_11764);
nor U12279 (N_12279,N_11463,N_11544);
xnor U12280 (N_12280,N_11963,N_11968);
xnor U12281 (N_12281,N_11880,N_11201);
or U12282 (N_12282,N_11830,N_11009);
nor U12283 (N_12283,N_11784,N_11177);
nor U12284 (N_12284,N_11383,N_11545);
nor U12285 (N_12285,N_11950,N_11329);
or U12286 (N_12286,N_11981,N_11625);
nor U12287 (N_12287,N_11582,N_11109);
and U12288 (N_12288,N_11278,N_11210);
and U12289 (N_12289,N_11939,N_11996);
nand U12290 (N_12290,N_11041,N_11863);
nor U12291 (N_12291,N_11437,N_11187);
xnor U12292 (N_12292,N_11111,N_11268);
and U12293 (N_12293,N_11611,N_11428);
or U12294 (N_12294,N_11856,N_11698);
nand U12295 (N_12295,N_11747,N_11139);
nand U12296 (N_12296,N_11962,N_11575);
or U12297 (N_12297,N_11423,N_11490);
xnor U12298 (N_12298,N_11977,N_11787);
nor U12299 (N_12299,N_11282,N_11315);
nand U12300 (N_12300,N_11682,N_11374);
nor U12301 (N_12301,N_11452,N_11655);
or U12302 (N_12302,N_11668,N_11186);
and U12303 (N_12303,N_11672,N_11172);
nand U12304 (N_12304,N_11276,N_11676);
and U12305 (N_12305,N_11673,N_11522);
nor U12306 (N_12306,N_11193,N_11687);
xnor U12307 (N_12307,N_11849,N_11912);
or U12308 (N_12308,N_11125,N_11455);
and U12309 (N_12309,N_11757,N_11881);
or U12310 (N_12310,N_11056,N_11373);
xor U12311 (N_12311,N_11179,N_11833);
xnor U12312 (N_12312,N_11997,N_11453);
xnor U12313 (N_12313,N_11864,N_11395);
and U12314 (N_12314,N_11049,N_11391);
nand U12315 (N_12315,N_11951,N_11732);
nand U12316 (N_12316,N_11571,N_11662);
and U12317 (N_12317,N_11017,N_11412);
and U12318 (N_12318,N_11949,N_11772);
nand U12319 (N_12319,N_11624,N_11945);
and U12320 (N_12320,N_11850,N_11843);
xnor U12321 (N_12321,N_11320,N_11030);
nor U12322 (N_12322,N_11791,N_11059);
or U12323 (N_12323,N_11766,N_11233);
nand U12324 (N_12324,N_11140,N_11785);
and U12325 (N_12325,N_11941,N_11569);
xnor U12326 (N_12326,N_11136,N_11755);
nand U12327 (N_12327,N_11602,N_11972);
xor U12328 (N_12328,N_11242,N_11372);
or U12329 (N_12329,N_11899,N_11189);
xnor U12330 (N_12330,N_11942,N_11204);
xnor U12331 (N_12331,N_11010,N_11810);
nor U12332 (N_12332,N_11882,N_11597);
or U12333 (N_12333,N_11558,N_11507);
xnor U12334 (N_12334,N_11515,N_11985);
xor U12335 (N_12335,N_11617,N_11352);
nand U12336 (N_12336,N_11307,N_11011);
nor U12337 (N_12337,N_11040,N_11476);
or U12338 (N_12338,N_11018,N_11149);
nor U12339 (N_12339,N_11521,N_11718);
xor U12340 (N_12340,N_11748,N_11322);
xor U12341 (N_12341,N_11564,N_11252);
and U12342 (N_12342,N_11514,N_11375);
xor U12343 (N_12343,N_11153,N_11526);
nor U12344 (N_12344,N_11245,N_11107);
nor U12345 (N_12345,N_11321,N_11553);
xnor U12346 (N_12346,N_11388,N_11585);
and U12347 (N_12347,N_11146,N_11663);
and U12348 (N_12348,N_11895,N_11456);
or U12349 (N_12349,N_11133,N_11686);
nand U12350 (N_12350,N_11434,N_11699);
nand U12351 (N_12351,N_11064,N_11667);
or U12352 (N_12352,N_11114,N_11566);
and U12353 (N_12353,N_11411,N_11195);
nand U12354 (N_12354,N_11019,N_11106);
xor U12355 (N_12355,N_11828,N_11519);
nand U12356 (N_12356,N_11050,N_11353);
or U12357 (N_12357,N_11712,N_11262);
nand U12358 (N_12358,N_11089,N_11260);
and U12359 (N_12359,N_11369,N_11956);
and U12360 (N_12360,N_11108,N_11586);
xor U12361 (N_12361,N_11664,N_11639);
nand U12362 (N_12362,N_11704,N_11470);
or U12363 (N_12363,N_11536,N_11227);
nand U12364 (N_12364,N_11270,N_11870);
or U12365 (N_12365,N_11356,N_11670);
xor U12366 (N_12366,N_11661,N_11503);
xnor U12367 (N_12367,N_11410,N_11844);
xnor U12368 (N_12368,N_11818,N_11649);
or U12369 (N_12369,N_11811,N_11166);
nand U12370 (N_12370,N_11419,N_11441);
nor U12371 (N_12371,N_11884,N_11488);
nor U12372 (N_12372,N_11325,N_11076);
and U12373 (N_12373,N_11472,N_11824);
nor U12374 (N_12374,N_11826,N_11331);
or U12375 (N_12375,N_11223,N_11920);
or U12376 (N_12376,N_11161,N_11869);
or U12377 (N_12377,N_11556,N_11674);
and U12378 (N_12378,N_11105,N_11433);
or U12379 (N_12379,N_11910,N_11241);
xnor U12380 (N_12380,N_11295,N_11217);
xnor U12381 (N_12381,N_11368,N_11656);
nor U12382 (N_12382,N_11057,N_11308);
and U12383 (N_12383,N_11390,N_11037);
nor U12384 (N_12384,N_11980,N_11835);
xnor U12385 (N_12385,N_11823,N_11385);
and U12386 (N_12386,N_11022,N_11646);
nor U12387 (N_12387,N_11947,N_11033);
or U12388 (N_12388,N_11741,N_11199);
nand U12389 (N_12389,N_11778,N_11892);
nand U12390 (N_12390,N_11537,N_11801);
xnor U12391 (N_12391,N_11077,N_11487);
nand U12392 (N_12392,N_11771,N_11933);
and U12393 (N_12393,N_11243,N_11231);
and U12394 (N_12394,N_11198,N_11418);
or U12395 (N_12395,N_11777,N_11902);
xnor U12396 (N_12396,N_11337,N_11609);
nand U12397 (N_12397,N_11756,N_11638);
nand U12398 (N_12398,N_11449,N_11952);
nand U12399 (N_12399,N_11905,N_11821);
nand U12400 (N_12400,N_11063,N_11316);
xor U12401 (N_12401,N_11031,N_11134);
and U12402 (N_12402,N_11812,N_11099);
nor U12403 (N_12403,N_11091,N_11458);
or U12404 (N_12404,N_11264,N_11324);
nor U12405 (N_12405,N_11648,N_11925);
or U12406 (N_12406,N_11209,N_11448);
or U12407 (N_12407,N_11923,N_11967);
nor U12408 (N_12408,N_11020,N_11027);
nor U12409 (N_12409,N_11790,N_11928);
xnor U12410 (N_12410,N_11736,N_11580);
xnor U12411 (N_12411,N_11918,N_11658);
and U12412 (N_12412,N_11358,N_11202);
or U12413 (N_12413,N_11969,N_11694);
and U12414 (N_12414,N_11003,N_11505);
or U12415 (N_12415,N_11328,N_11174);
and U12416 (N_12416,N_11246,N_11462);
nor U12417 (N_12417,N_11479,N_11865);
nand U12418 (N_12418,N_11761,N_11815);
or U12419 (N_12419,N_11001,N_11538);
and U12420 (N_12420,N_11930,N_11635);
or U12421 (N_12421,N_11137,N_11719);
and U12422 (N_12422,N_11044,N_11708);
or U12423 (N_12423,N_11274,N_11955);
nand U12424 (N_12424,N_11127,N_11446);
nand U12425 (N_12425,N_11606,N_11365);
nor U12426 (N_12426,N_11998,N_11357);
nor U12427 (N_12427,N_11675,N_11797);
xor U12428 (N_12428,N_11443,N_11188);
xnor U12429 (N_12429,N_11102,N_11943);
or U12430 (N_12430,N_11465,N_11120);
nand U12431 (N_12431,N_11577,N_11561);
nor U12432 (N_12432,N_11203,N_11750);
or U12433 (N_12433,N_11679,N_11720);
or U12434 (N_12434,N_11896,N_11742);
and U12435 (N_12435,N_11366,N_11807);
nand U12436 (N_12436,N_11795,N_11110);
xor U12437 (N_12437,N_11104,N_11510);
and U12438 (N_12438,N_11919,N_11532);
and U12439 (N_12439,N_11568,N_11457);
nor U12440 (N_12440,N_11475,N_11394);
and U12441 (N_12441,N_11851,N_11420);
xnor U12442 (N_12442,N_11384,N_11628);
nor U12443 (N_12443,N_11471,N_11822);
xnor U12444 (N_12444,N_11678,N_11877);
nand U12445 (N_12445,N_11184,N_11847);
or U12446 (N_12446,N_11644,N_11511);
and U12447 (N_12447,N_11222,N_11300);
nand U12448 (N_12448,N_11529,N_11913);
nand U12449 (N_12449,N_11126,N_11878);
and U12450 (N_12450,N_11623,N_11169);
nor U12451 (N_12451,N_11666,N_11224);
nand U12452 (N_12452,N_11145,N_11494);
nor U12453 (N_12453,N_11311,N_11898);
and U12454 (N_12454,N_11859,N_11906);
or U12455 (N_12455,N_11425,N_11043);
and U12456 (N_12456,N_11387,N_11994);
and U12457 (N_12457,N_11608,N_11069);
nand U12458 (N_12458,N_11364,N_11528);
nand U12459 (N_12459,N_11014,N_11310);
or U12460 (N_12460,N_11776,N_11396);
nand U12461 (N_12461,N_11042,N_11974);
nand U12462 (N_12462,N_11271,N_11306);
and U12463 (N_12463,N_11416,N_11323);
nand U12464 (N_12464,N_11533,N_11466);
xnor U12465 (N_12465,N_11961,N_11498);
nand U12466 (N_12466,N_11442,N_11727);
nand U12467 (N_12467,N_11450,N_11397);
or U12468 (N_12468,N_11485,N_11006);
xnor U12469 (N_12469,N_11338,N_11716);
or U12470 (N_12470,N_11256,N_11591);
or U12471 (N_12471,N_11513,N_11565);
nand U12472 (N_12472,N_11746,N_11230);
nor U12473 (N_12473,N_11024,N_11039);
xnor U12474 (N_12474,N_11212,N_11763);
or U12475 (N_12475,N_11613,N_11788);
or U12476 (N_12476,N_11769,N_11860);
and U12477 (N_12477,N_11197,N_11347);
or U12478 (N_12478,N_11827,N_11317);
nand U12479 (N_12479,N_11012,N_11194);
nor U12480 (N_12480,N_11975,N_11904);
and U12481 (N_12481,N_11181,N_11548);
nand U12482 (N_12482,N_11820,N_11524);
nor U12483 (N_12483,N_11173,N_11845);
and U12484 (N_12484,N_11660,N_11589);
and U12485 (N_12485,N_11607,N_11731);
xnor U12486 (N_12486,N_11861,N_11825);
nand U12487 (N_12487,N_11239,N_11685);
nand U12488 (N_12488,N_11493,N_11700);
nand U12489 (N_12489,N_11066,N_11730);
xnor U12490 (N_12490,N_11348,N_11234);
nand U12491 (N_12491,N_11363,N_11178);
or U12492 (N_12492,N_11552,N_11132);
and U12493 (N_12493,N_11576,N_11029);
or U12494 (N_12494,N_11701,N_11313);
or U12495 (N_12495,N_11726,N_11523);
nor U12496 (N_12496,N_11645,N_11908);
nor U12497 (N_12497,N_11762,N_11610);
nand U12498 (N_12498,N_11415,N_11643);
xnor U12499 (N_12499,N_11809,N_11958);
or U12500 (N_12500,N_11977,N_11159);
and U12501 (N_12501,N_11773,N_11401);
nor U12502 (N_12502,N_11586,N_11087);
nor U12503 (N_12503,N_11334,N_11337);
xor U12504 (N_12504,N_11987,N_11682);
and U12505 (N_12505,N_11922,N_11464);
nand U12506 (N_12506,N_11422,N_11844);
nand U12507 (N_12507,N_11465,N_11943);
and U12508 (N_12508,N_11442,N_11745);
nand U12509 (N_12509,N_11483,N_11341);
nor U12510 (N_12510,N_11501,N_11021);
nor U12511 (N_12511,N_11173,N_11070);
xnor U12512 (N_12512,N_11936,N_11383);
nand U12513 (N_12513,N_11769,N_11509);
nor U12514 (N_12514,N_11979,N_11451);
nor U12515 (N_12515,N_11522,N_11782);
nand U12516 (N_12516,N_11867,N_11030);
nor U12517 (N_12517,N_11722,N_11032);
nor U12518 (N_12518,N_11455,N_11119);
nand U12519 (N_12519,N_11655,N_11549);
and U12520 (N_12520,N_11829,N_11301);
xor U12521 (N_12521,N_11813,N_11505);
nand U12522 (N_12522,N_11076,N_11760);
nor U12523 (N_12523,N_11379,N_11552);
xor U12524 (N_12524,N_11225,N_11101);
and U12525 (N_12525,N_11898,N_11254);
or U12526 (N_12526,N_11906,N_11827);
and U12527 (N_12527,N_11150,N_11602);
xnor U12528 (N_12528,N_11854,N_11285);
xnor U12529 (N_12529,N_11395,N_11383);
nand U12530 (N_12530,N_11545,N_11927);
nor U12531 (N_12531,N_11707,N_11209);
xor U12532 (N_12532,N_11810,N_11355);
xor U12533 (N_12533,N_11872,N_11907);
and U12534 (N_12534,N_11041,N_11057);
xor U12535 (N_12535,N_11793,N_11706);
or U12536 (N_12536,N_11797,N_11957);
xnor U12537 (N_12537,N_11310,N_11051);
and U12538 (N_12538,N_11583,N_11342);
and U12539 (N_12539,N_11515,N_11911);
nand U12540 (N_12540,N_11390,N_11388);
or U12541 (N_12541,N_11366,N_11013);
and U12542 (N_12542,N_11532,N_11098);
and U12543 (N_12543,N_11130,N_11791);
or U12544 (N_12544,N_11423,N_11391);
nor U12545 (N_12545,N_11645,N_11831);
xnor U12546 (N_12546,N_11852,N_11972);
xor U12547 (N_12547,N_11596,N_11384);
nor U12548 (N_12548,N_11906,N_11064);
and U12549 (N_12549,N_11513,N_11052);
nor U12550 (N_12550,N_11013,N_11217);
and U12551 (N_12551,N_11803,N_11574);
and U12552 (N_12552,N_11873,N_11618);
nand U12553 (N_12553,N_11942,N_11493);
and U12554 (N_12554,N_11345,N_11083);
nand U12555 (N_12555,N_11752,N_11205);
and U12556 (N_12556,N_11340,N_11108);
nor U12557 (N_12557,N_11776,N_11878);
or U12558 (N_12558,N_11422,N_11683);
nand U12559 (N_12559,N_11365,N_11586);
xor U12560 (N_12560,N_11883,N_11704);
and U12561 (N_12561,N_11239,N_11482);
nor U12562 (N_12562,N_11282,N_11679);
xnor U12563 (N_12563,N_11257,N_11738);
and U12564 (N_12564,N_11427,N_11100);
and U12565 (N_12565,N_11070,N_11442);
nand U12566 (N_12566,N_11040,N_11019);
xor U12567 (N_12567,N_11005,N_11831);
or U12568 (N_12568,N_11406,N_11973);
nand U12569 (N_12569,N_11031,N_11300);
nand U12570 (N_12570,N_11216,N_11428);
or U12571 (N_12571,N_11748,N_11131);
xnor U12572 (N_12572,N_11469,N_11368);
and U12573 (N_12573,N_11965,N_11623);
and U12574 (N_12574,N_11931,N_11386);
and U12575 (N_12575,N_11861,N_11605);
xnor U12576 (N_12576,N_11010,N_11200);
nor U12577 (N_12577,N_11075,N_11829);
xor U12578 (N_12578,N_11633,N_11103);
nor U12579 (N_12579,N_11735,N_11903);
and U12580 (N_12580,N_11651,N_11268);
xor U12581 (N_12581,N_11142,N_11440);
xnor U12582 (N_12582,N_11388,N_11764);
or U12583 (N_12583,N_11216,N_11473);
xor U12584 (N_12584,N_11293,N_11831);
or U12585 (N_12585,N_11374,N_11529);
xnor U12586 (N_12586,N_11743,N_11770);
xnor U12587 (N_12587,N_11887,N_11820);
or U12588 (N_12588,N_11749,N_11653);
xor U12589 (N_12589,N_11210,N_11918);
nor U12590 (N_12590,N_11651,N_11198);
xnor U12591 (N_12591,N_11844,N_11353);
or U12592 (N_12592,N_11128,N_11010);
nand U12593 (N_12593,N_11389,N_11999);
and U12594 (N_12594,N_11372,N_11720);
or U12595 (N_12595,N_11068,N_11415);
and U12596 (N_12596,N_11369,N_11295);
nand U12597 (N_12597,N_11022,N_11057);
nand U12598 (N_12598,N_11748,N_11713);
xor U12599 (N_12599,N_11908,N_11168);
and U12600 (N_12600,N_11524,N_11504);
or U12601 (N_12601,N_11150,N_11600);
xor U12602 (N_12602,N_11442,N_11088);
xor U12603 (N_12603,N_11244,N_11656);
nand U12604 (N_12604,N_11673,N_11246);
xor U12605 (N_12605,N_11202,N_11599);
nor U12606 (N_12606,N_11314,N_11219);
and U12607 (N_12607,N_11984,N_11994);
xor U12608 (N_12608,N_11618,N_11751);
or U12609 (N_12609,N_11428,N_11675);
and U12610 (N_12610,N_11560,N_11223);
and U12611 (N_12611,N_11278,N_11492);
nor U12612 (N_12612,N_11335,N_11561);
or U12613 (N_12613,N_11869,N_11218);
nor U12614 (N_12614,N_11652,N_11317);
and U12615 (N_12615,N_11510,N_11205);
xor U12616 (N_12616,N_11852,N_11452);
nand U12617 (N_12617,N_11871,N_11996);
or U12618 (N_12618,N_11329,N_11837);
and U12619 (N_12619,N_11677,N_11087);
and U12620 (N_12620,N_11045,N_11372);
and U12621 (N_12621,N_11503,N_11335);
or U12622 (N_12622,N_11136,N_11787);
xnor U12623 (N_12623,N_11821,N_11959);
nor U12624 (N_12624,N_11661,N_11259);
or U12625 (N_12625,N_11283,N_11124);
and U12626 (N_12626,N_11834,N_11506);
nand U12627 (N_12627,N_11987,N_11367);
nor U12628 (N_12628,N_11999,N_11421);
nand U12629 (N_12629,N_11788,N_11859);
and U12630 (N_12630,N_11351,N_11856);
nand U12631 (N_12631,N_11487,N_11412);
nand U12632 (N_12632,N_11304,N_11973);
nor U12633 (N_12633,N_11044,N_11835);
nand U12634 (N_12634,N_11371,N_11051);
nand U12635 (N_12635,N_11090,N_11213);
nand U12636 (N_12636,N_11336,N_11750);
and U12637 (N_12637,N_11244,N_11975);
nor U12638 (N_12638,N_11234,N_11793);
xor U12639 (N_12639,N_11681,N_11452);
nand U12640 (N_12640,N_11415,N_11801);
and U12641 (N_12641,N_11052,N_11772);
nand U12642 (N_12642,N_11642,N_11240);
nand U12643 (N_12643,N_11876,N_11874);
xor U12644 (N_12644,N_11749,N_11411);
nand U12645 (N_12645,N_11671,N_11080);
and U12646 (N_12646,N_11337,N_11926);
or U12647 (N_12647,N_11501,N_11005);
or U12648 (N_12648,N_11480,N_11684);
nor U12649 (N_12649,N_11654,N_11559);
or U12650 (N_12650,N_11756,N_11814);
nand U12651 (N_12651,N_11970,N_11132);
nor U12652 (N_12652,N_11662,N_11272);
xor U12653 (N_12653,N_11463,N_11842);
xnor U12654 (N_12654,N_11554,N_11250);
and U12655 (N_12655,N_11421,N_11939);
or U12656 (N_12656,N_11542,N_11384);
and U12657 (N_12657,N_11352,N_11144);
nand U12658 (N_12658,N_11366,N_11442);
nor U12659 (N_12659,N_11269,N_11097);
and U12660 (N_12660,N_11930,N_11938);
nor U12661 (N_12661,N_11790,N_11311);
and U12662 (N_12662,N_11816,N_11671);
nand U12663 (N_12663,N_11447,N_11570);
nand U12664 (N_12664,N_11022,N_11806);
nand U12665 (N_12665,N_11669,N_11335);
nor U12666 (N_12666,N_11192,N_11380);
and U12667 (N_12667,N_11799,N_11572);
nor U12668 (N_12668,N_11634,N_11130);
xor U12669 (N_12669,N_11819,N_11970);
and U12670 (N_12670,N_11798,N_11036);
and U12671 (N_12671,N_11501,N_11445);
or U12672 (N_12672,N_11387,N_11774);
and U12673 (N_12673,N_11770,N_11269);
xor U12674 (N_12674,N_11524,N_11938);
and U12675 (N_12675,N_11213,N_11632);
or U12676 (N_12676,N_11745,N_11787);
nand U12677 (N_12677,N_11329,N_11113);
nor U12678 (N_12678,N_11059,N_11273);
nand U12679 (N_12679,N_11334,N_11485);
nand U12680 (N_12680,N_11702,N_11027);
nor U12681 (N_12681,N_11667,N_11035);
or U12682 (N_12682,N_11503,N_11989);
and U12683 (N_12683,N_11381,N_11355);
and U12684 (N_12684,N_11865,N_11896);
and U12685 (N_12685,N_11915,N_11452);
xor U12686 (N_12686,N_11078,N_11487);
nand U12687 (N_12687,N_11135,N_11610);
or U12688 (N_12688,N_11159,N_11575);
and U12689 (N_12689,N_11485,N_11509);
xor U12690 (N_12690,N_11111,N_11447);
nand U12691 (N_12691,N_11391,N_11673);
nor U12692 (N_12692,N_11190,N_11886);
nand U12693 (N_12693,N_11030,N_11300);
nor U12694 (N_12694,N_11450,N_11755);
xor U12695 (N_12695,N_11410,N_11878);
xor U12696 (N_12696,N_11086,N_11825);
xor U12697 (N_12697,N_11455,N_11074);
xor U12698 (N_12698,N_11986,N_11143);
or U12699 (N_12699,N_11101,N_11345);
xor U12700 (N_12700,N_11078,N_11737);
and U12701 (N_12701,N_11198,N_11471);
xor U12702 (N_12702,N_11921,N_11173);
or U12703 (N_12703,N_11050,N_11792);
or U12704 (N_12704,N_11127,N_11869);
nand U12705 (N_12705,N_11691,N_11212);
xnor U12706 (N_12706,N_11321,N_11018);
xnor U12707 (N_12707,N_11834,N_11046);
or U12708 (N_12708,N_11238,N_11200);
or U12709 (N_12709,N_11739,N_11970);
and U12710 (N_12710,N_11345,N_11977);
xnor U12711 (N_12711,N_11065,N_11460);
nand U12712 (N_12712,N_11637,N_11996);
nand U12713 (N_12713,N_11243,N_11029);
nor U12714 (N_12714,N_11258,N_11436);
and U12715 (N_12715,N_11943,N_11804);
and U12716 (N_12716,N_11858,N_11510);
xor U12717 (N_12717,N_11923,N_11312);
nand U12718 (N_12718,N_11608,N_11501);
nor U12719 (N_12719,N_11653,N_11897);
xor U12720 (N_12720,N_11707,N_11900);
nand U12721 (N_12721,N_11832,N_11448);
xor U12722 (N_12722,N_11163,N_11848);
xnor U12723 (N_12723,N_11221,N_11089);
nor U12724 (N_12724,N_11896,N_11603);
and U12725 (N_12725,N_11039,N_11769);
nor U12726 (N_12726,N_11338,N_11829);
and U12727 (N_12727,N_11636,N_11143);
or U12728 (N_12728,N_11556,N_11212);
and U12729 (N_12729,N_11853,N_11711);
or U12730 (N_12730,N_11220,N_11047);
xor U12731 (N_12731,N_11200,N_11192);
nand U12732 (N_12732,N_11339,N_11278);
and U12733 (N_12733,N_11954,N_11173);
nor U12734 (N_12734,N_11421,N_11680);
xor U12735 (N_12735,N_11435,N_11847);
nor U12736 (N_12736,N_11280,N_11543);
or U12737 (N_12737,N_11640,N_11724);
or U12738 (N_12738,N_11310,N_11787);
xor U12739 (N_12739,N_11706,N_11951);
and U12740 (N_12740,N_11874,N_11861);
xor U12741 (N_12741,N_11822,N_11702);
nand U12742 (N_12742,N_11155,N_11956);
nor U12743 (N_12743,N_11669,N_11698);
nand U12744 (N_12744,N_11204,N_11985);
nor U12745 (N_12745,N_11360,N_11965);
xor U12746 (N_12746,N_11315,N_11407);
xnor U12747 (N_12747,N_11581,N_11021);
nand U12748 (N_12748,N_11282,N_11178);
and U12749 (N_12749,N_11984,N_11525);
and U12750 (N_12750,N_11249,N_11192);
or U12751 (N_12751,N_11639,N_11258);
or U12752 (N_12752,N_11213,N_11846);
nor U12753 (N_12753,N_11535,N_11451);
and U12754 (N_12754,N_11490,N_11947);
xnor U12755 (N_12755,N_11666,N_11015);
nor U12756 (N_12756,N_11153,N_11751);
or U12757 (N_12757,N_11870,N_11331);
xnor U12758 (N_12758,N_11075,N_11958);
nand U12759 (N_12759,N_11333,N_11356);
nor U12760 (N_12760,N_11450,N_11642);
nor U12761 (N_12761,N_11086,N_11272);
nor U12762 (N_12762,N_11819,N_11550);
nand U12763 (N_12763,N_11713,N_11782);
xnor U12764 (N_12764,N_11913,N_11034);
xor U12765 (N_12765,N_11224,N_11164);
nand U12766 (N_12766,N_11145,N_11599);
or U12767 (N_12767,N_11153,N_11614);
nor U12768 (N_12768,N_11663,N_11629);
nand U12769 (N_12769,N_11502,N_11569);
nand U12770 (N_12770,N_11883,N_11648);
xnor U12771 (N_12771,N_11214,N_11388);
nand U12772 (N_12772,N_11166,N_11332);
nand U12773 (N_12773,N_11115,N_11737);
xnor U12774 (N_12774,N_11371,N_11960);
or U12775 (N_12775,N_11659,N_11784);
nand U12776 (N_12776,N_11233,N_11214);
nand U12777 (N_12777,N_11105,N_11412);
nor U12778 (N_12778,N_11510,N_11411);
nor U12779 (N_12779,N_11752,N_11147);
or U12780 (N_12780,N_11051,N_11236);
or U12781 (N_12781,N_11508,N_11125);
xor U12782 (N_12782,N_11238,N_11743);
xnor U12783 (N_12783,N_11967,N_11916);
and U12784 (N_12784,N_11903,N_11436);
xnor U12785 (N_12785,N_11148,N_11204);
or U12786 (N_12786,N_11529,N_11587);
xnor U12787 (N_12787,N_11543,N_11071);
and U12788 (N_12788,N_11307,N_11078);
nor U12789 (N_12789,N_11485,N_11712);
nor U12790 (N_12790,N_11863,N_11467);
xor U12791 (N_12791,N_11412,N_11820);
and U12792 (N_12792,N_11088,N_11323);
and U12793 (N_12793,N_11813,N_11927);
or U12794 (N_12794,N_11187,N_11614);
and U12795 (N_12795,N_11203,N_11041);
xnor U12796 (N_12796,N_11458,N_11419);
nor U12797 (N_12797,N_11571,N_11496);
nor U12798 (N_12798,N_11255,N_11824);
xnor U12799 (N_12799,N_11062,N_11119);
nand U12800 (N_12800,N_11031,N_11324);
and U12801 (N_12801,N_11974,N_11440);
xnor U12802 (N_12802,N_11014,N_11008);
nand U12803 (N_12803,N_11008,N_11284);
nor U12804 (N_12804,N_11625,N_11340);
xor U12805 (N_12805,N_11990,N_11679);
and U12806 (N_12806,N_11166,N_11297);
xnor U12807 (N_12807,N_11960,N_11270);
xor U12808 (N_12808,N_11611,N_11232);
nor U12809 (N_12809,N_11950,N_11438);
nor U12810 (N_12810,N_11634,N_11620);
or U12811 (N_12811,N_11264,N_11101);
and U12812 (N_12812,N_11977,N_11722);
and U12813 (N_12813,N_11597,N_11080);
and U12814 (N_12814,N_11591,N_11885);
xor U12815 (N_12815,N_11944,N_11759);
nand U12816 (N_12816,N_11336,N_11210);
or U12817 (N_12817,N_11573,N_11393);
xnor U12818 (N_12818,N_11376,N_11933);
nor U12819 (N_12819,N_11771,N_11797);
nor U12820 (N_12820,N_11754,N_11722);
xor U12821 (N_12821,N_11348,N_11670);
or U12822 (N_12822,N_11196,N_11359);
nand U12823 (N_12823,N_11759,N_11540);
nand U12824 (N_12824,N_11249,N_11630);
nand U12825 (N_12825,N_11075,N_11194);
xor U12826 (N_12826,N_11407,N_11187);
nand U12827 (N_12827,N_11132,N_11162);
xnor U12828 (N_12828,N_11397,N_11053);
or U12829 (N_12829,N_11195,N_11629);
and U12830 (N_12830,N_11635,N_11711);
or U12831 (N_12831,N_11100,N_11005);
and U12832 (N_12832,N_11180,N_11456);
or U12833 (N_12833,N_11945,N_11959);
and U12834 (N_12834,N_11010,N_11209);
nor U12835 (N_12835,N_11887,N_11308);
xnor U12836 (N_12836,N_11167,N_11129);
nand U12837 (N_12837,N_11072,N_11481);
nor U12838 (N_12838,N_11493,N_11397);
nand U12839 (N_12839,N_11491,N_11119);
nor U12840 (N_12840,N_11833,N_11139);
nand U12841 (N_12841,N_11871,N_11302);
or U12842 (N_12842,N_11114,N_11228);
nand U12843 (N_12843,N_11890,N_11782);
and U12844 (N_12844,N_11953,N_11992);
and U12845 (N_12845,N_11392,N_11517);
nor U12846 (N_12846,N_11917,N_11737);
or U12847 (N_12847,N_11407,N_11341);
or U12848 (N_12848,N_11188,N_11239);
xor U12849 (N_12849,N_11430,N_11469);
nor U12850 (N_12850,N_11201,N_11434);
nor U12851 (N_12851,N_11603,N_11573);
and U12852 (N_12852,N_11752,N_11359);
xor U12853 (N_12853,N_11520,N_11829);
or U12854 (N_12854,N_11230,N_11358);
or U12855 (N_12855,N_11788,N_11117);
nand U12856 (N_12856,N_11000,N_11606);
or U12857 (N_12857,N_11399,N_11468);
and U12858 (N_12858,N_11739,N_11381);
nor U12859 (N_12859,N_11334,N_11174);
nand U12860 (N_12860,N_11275,N_11846);
xor U12861 (N_12861,N_11648,N_11123);
nand U12862 (N_12862,N_11855,N_11527);
and U12863 (N_12863,N_11327,N_11413);
nor U12864 (N_12864,N_11228,N_11608);
and U12865 (N_12865,N_11848,N_11144);
and U12866 (N_12866,N_11092,N_11832);
xor U12867 (N_12867,N_11060,N_11224);
and U12868 (N_12868,N_11339,N_11621);
nand U12869 (N_12869,N_11235,N_11472);
nand U12870 (N_12870,N_11011,N_11481);
xnor U12871 (N_12871,N_11844,N_11487);
nand U12872 (N_12872,N_11397,N_11897);
nand U12873 (N_12873,N_11307,N_11029);
and U12874 (N_12874,N_11620,N_11429);
nand U12875 (N_12875,N_11176,N_11162);
xnor U12876 (N_12876,N_11213,N_11004);
nor U12877 (N_12877,N_11360,N_11520);
and U12878 (N_12878,N_11477,N_11090);
or U12879 (N_12879,N_11322,N_11083);
or U12880 (N_12880,N_11393,N_11412);
or U12881 (N_12881,N_11778,N_11195);
nand U12882 (N_12882,N_11962,N_11853);
nor U12883 (N_12883,N_11150,N_11515);
or U12884 (N_12884,N_11414,N_11270);
xnor U12885 (N_12885,N_11959,N_11430);
xnor U12886 (N_12886,N_11029,N_11809);
nor U12887 (N_12887,N_11464,N_11214);
or U12888 (N_12888,N_11336,N_11251);
or U12889 (N_12889,N_11263,N_11533);
nor U12890 (N_12890,N_11763,N_11171);
nor U12891 (N_12891,N_11645,N_11227);
xnor U12892 (N_12892,N_11296,N_11772);
nor U12893 (N_12893,N_11991,N_11876);
or U12894 (N_12894,N_11103,N_11720);
nand U12895 (N_12895,N_11630,N_11174);
or U12896 (N_12896,N_11722,N_11405);
xor U12897 (N_12897,N_11417,N_11215);
nor U12898 (N_12898,N_11917,N_11663);
xor U12899 (N_12899,N_11060,N_11976);
xor U12900 (N_12900,N_11003,N_11254);
or U12901 (N_12901,N_11913,N_11721);
and U12902 (N_12902,N_11795,N_11694);
xor U12903 (N_12903,N_11108,N_11334);
nand U12904 (N_12904,N_11807,N_11973);
or U12905 (N_12905,N_11184,N_11958);
and U12906 (N_12906,N_11589,N_11058);
xor U12907 (N_12907,N_11657,N_11898);
or U12908 (N_12908,N_11291,N_11512);
and U12909 (N_12909,N_11287,N_11920);
xnor U12910 (N_12910,N_11476,N_11285);
nor U12911 (N_12911,N_11157,N_11755);
or U12912 (N_12912,N_11154,N_11338);
nand U12913 (N_12913,N_11305,N_11227);
nor U12914 (N_12914,N_11245,N_11348);
and U12915 (N_12915,N_11375,N_11894);
and U12916 (N_12916,N_11405,N_11154);
and U12917 (N_12917,N_11197,N_11963);
xor U12918 (N_12918,N_11788,N_11390);
nor U12919 (N_12919,N_11693,N_11825);
and U12920 (N_12920,N_11819,N_11999);
nand U12921 (N_12921,N_11005,N_11196);
or U12922 (N_12922,N_11040,N_11394);
xnor U12923 (N_12923,N_11100,N_11620);
or U12924 (N_12924,N_11591,N_11509);
and U12925 (N_12925,N_11013,N_11864);
nand U12926 (N_12926,N_11665,N_11329);
nor U12927 (N_12927,N_11665,N_11387);
xor U12928 (N_12928,N_11763,N_11798);
or U12929 (N_12929,N_11927,N_11331);
nand U12930 (N_12930,N_11758,N_11844);
or U12931 (N_12931,N_11680,N_11386);
xor U12932 (N_12932,N_11201,N_11054);
nand U12933 (N_12933,N_11881,N_11359);
nand U12934 (N_12934,N_11090,N_11069);
xor U12935 (N_12935,N_11324,N_11585);
nand U12936 (N_12936,N_11628,N_11261);
or U12937 (N_12937,N_11896,N_11906);
nand U12938 (N_12938,N_11400,N_11509);
nor U12939 (N_12939,N_11183,N_11985);
nand U12940 (N_12940,N_11695,N_11167);
xnor U12941 (N_12941,N_11120,N_11548);
or U12942 (N_12942,N_11080,N_11006);
nand U12943 (N_12943,N_11582,N_11603);
or U12944 (N_12944,N_11127,N_11464);
xor U12945 (N_12945,N_11250,N_11519);
and U12946 (N_12946,N_11307,N_11536);
nand U12947 (N_12947,N_11284,N_11684);
nor U12948 (N_12948,N_11852,N_11138);
or U12949 (N_12949,N_11643,N_11510);
nand U12950 (N_12950,N_11845,N_11723);
nand U12951 (N_12951,N_11764,N_11027);
and U12952 (N_12952,N_11876,N_11130);
nor U12953 (N_12953,N_11689,N_11758);
xor U12954 (N_12954,N_11108,N_11544);
and U12955 (N_12955,N_11281,N_11143);
and U12956 (N_12956,N_11759,N_11874);
and U12957 (N_12957,N_11054,N_11637);
xor U12958 (N_12958,N_11452,N_11595);
nand U12959 (N_12959,N_11533,N_11109);
and U12960 (N_12960,N_11417,N_11907);
and U12961 (N_12961,N_11933,N_11307);
or U12962 (N_12962,N_11985,N_11688);
nand U12963 (N_12963,N_11769,N_11239);
nor U12964 (N_12964,N_11844,N_11811);
nor U12965 (N_12965,N_11423,N_11150);
and U12966 (N_12966,N_11272,N_11657);
or U12967 (N_12967,N_11304,N_11586);
or U12968 (N_12968,N_11274,N_11114);
or U12969 (N_12969,N_11016,N_11761);
xor U12970 (N_12970,N_11639,N_11813);
and U12971 (N_12971,N_11350,N_11423);
or U12972 (N_12972,N_11417,N_11700);
xor U12973 (N_12973,N_11213,N_11506);
and U12974 (N_12974,N_11264,N_11676);
nand U12975 (N_12975,N_11665,N_11834);
nor U12976 (N_12976,N_11004,N_11152);
nor U12977 (N_12977,N_11651,N_11569);
xor U12978 (N_12978,N_11788,N_11581);
nor U12979 (N_12979,N_11149,N_11171);
or U12980 (N_12980,N_11043,N_11008);
xor U12981 (N_12981,N_11234,N_11948);
nor U12982 (N_12982,N_11190,N_11906);
nand U12983 (N_12983,N_11787,N_11984);
and U12984 (N_12984,N_11587,N_11745);
and U12985 (N_12985,N_11477,N_11275);
nand U12986 (N_12986,N_11136,N_11206);
and U12987 (N_12987,N_11839,N_11087);
nor U12988 (N_12988,N_11648,N_11891);
nand U12989 (N_12989,N_11597,N_11510);
and U12990 (N_12990,N_11239,N_11394);
nor U12991 (N_12991,N_11199,N_11450);
xor U12992 (N_12992,N_11994,N_11086);
and U12993 (N_12993,N_11336,N_11728);
or U12994 (N_12994,N_11169,N_11008);
and U12995 (N_12995,N_11744,N_11329);
and U12996 (N_12996,N_11961,N_11967);
nor U12997 (N_12997,N_11385,N_11072);
and U12998 (N_12998,N_11889,N_11875);
and U12999 (N_12999,N_11029,N_11277);
nor U13000 (N_13000,N_12706,N_12909);
or U13001 (N_13001,N_12774,N_12784);
nor U13002 (N_13002,N_12973,N_12660);
nor U13003 (N_13003,N_12578,N_12567);
or U13004 (N_13004,N_12341,N_12627);
or U13005 (N_13005,N_12086,N_12943);
or U13006 (N_13006,N_12000,N_12599);
or U13007 (N_13007,N_12007,N_12367);
or U13008 (N_13008,N_12139,N_12842);
nand U13009 (N_13009,N_12622,N_12537);
and U13010 (N_13010,N_12179,N_12698);
or U13011 (N_13011,N_12484,N_12661);
and U13012 (N_13012,N_12299,N_12704);
and U13013 (N_13013,N_12041,N_12858);
nor U13014 (N_13014,N_12591,N_12383);
and U13015 (N_13015,N_12992,N_12566);
nor U13016 (N_13016,N_12589,N_12763);
nor U13017 (N_13017,N_12101,N_12662);
nor U13018 (N_13018,N_12320,N_12327);
and U13019 (N_13019,N_12056,N_12946);
nand U13020 (N_13020,N_12441,N_12244);
xor U13021 (N_13021,N_12167,N_12357);
nand U13022 (N_13022,N_12125,N_12918);
nor U13023 (N_13023,N_12982,N_12674);
nor U13024 (N_13024,N_12103,N_12306);
nor U13025 (N_13025,N_12342,N_12733);
or U13026 (N_13026,N_12551,N_12797);
nand U13027 (N_13027,N_12335,N_12488);
or U13028 (N_13028,N_12686,N_12016);
nand U13029 (N_13029,N_12328,N_12980);
nand U13030 (N_13030,N_12334,N_12251);
xnor U13031 (N_13031,N_12318,N_12965);
nor U13032 (N_13032,N_12496,N_12157);
nand U13033 (N_13033,N_12828,N_12431);
xnor U13034 (N_13034,N_12879,N_12501);
xor U13035 (N_13035,N_12750,N_12593);
xnor U13036 (N_13036,N_12022,N_12948);
nor U13037 (N_13037,N_12884,N_12846);
nand U13038 (N_13038,N_12539,N_12647);
nor U13039 (N_13039,N_12655,N_12767);
xor U13040 (N_13040,N_12751,N_12272);
xor U13041 (N_13041,N_12079,N_12527);
nor U13042 (N_13042,N_12074,N_12304);
nand U13043 (N_13043,N_12792,N_12931);
and U13044 (N_13044,N_12678,N_12906);
nor U13045 (N_13045,N_12423,N_12583);
nor U13046 (N_13046,N_12095,N_12407);
xnor U13047 (N_13047,N_12788,N_12021);
nand U13048 (N_13048,N_12302,N_12029);
xor U13049 (N_13049,N_12544,N_12033);
nand U13050 (N_13050,N_12135,N_12082);
and U13051 (N_13051,N_12778,N_12395);
or U13052 (N_13052,N_12497,N_12711);
nand U13053 (N_13053,N_12093,N_12026);
and U13054 (N_13054,N_12668,N_12749);
and U13055 (N_13055,N_12876,N_12229);
or U13056 (N_13056,N_12224,N_12826);
xnor U13057 (N_13057,N_12764,N_12845);
nand U13058 (N_13058,N_12349,N_12143);
and U13059 (N_13059,N_12374,N_12963);
nand U13060 (N_13060,N_12821,N_12449);
xnor U13061 (N_13061,N_12663,N_12574);
nor U13062 (N_13062,N_12008,N_12011);
or U13063 (N_13063,N_12570,N_12832);
or U13064 (N_13064,N_12192,N_12330);
and U13065 (N_13065,N_12260,N_12587);
or U13066 (N_13066,N_12205,N_12837);
and U13067 (N_13067,N_12315,N_12234);
nand U13068 (N_13068,N_12562,N_12576);
nor U13069 (N_13069,N_12927,N_12861);
xnor U13070 (N_13070,N_12178,N_12317);
nand U13071 (N_13071,N_12177,N_12406);
nor U13072 (N_13072,N_12890,N_12631);
nand U13073 (N_13073,N_12579,N_12267);
and U13074 (N_13074,N_12012,N_12250);
or U13075 (N_13075,N_12425,N_12226);
xnor U13076 (N_13076,N_12105,N_12940);
nor U13077 (N_13077,N_12872,N_12671);
nor U13078 (N_13078,N_12947,N_12530);
and U13079 (N_13079,N_12057,N_12731);
nor U13080 (N_13080,N_12380,N_12859);
and U13081 (N_13081,N_12993,N_12922);
xor U13082 (N_13082,N_12572,N_12967);
nand U13083 (N_13083,N_12006,N_12046);
xor U13084 (N_13084,N_12279,N_12217);
xor U13085 (N_13085,N_12734,N_12005);
nand U13086 (N_13086,N_12287,N_12880);
xor U13087 (N_13087,N_12398,N_12408);
and U13088 (N_13088,N_12471,N_12548);
or U13089 (N_13089,N_12636,N_12185);
nor U13090 (N_13090,N_12416,N_12198);
nor U13091 (N_13091,N_12687,N_12116);
xnor U13092 (N_13092,N_12151,N_12144);
or U13093 (N_13093,N_12897,N_12382);
or U13094 (N_13094,N_12856,N_12628);
xor U13095 (N_13095,N_12873,N_12483);
nand U13096 (N_13096,N_12352,N_12819);
and U13097 (N_13097,N_12370,N_12959);
nor U13098 (N_13098,N_12626,N_12487);
and U13099 (N_13099,N_12573,N_12545);
and U13100 (N_13100,N_12417,N_12632);
nand U13101 (N_13101,N_12075,N_12847);
or U13102 (N_13102,N_12600,N_12345);
nand U13103 (N_13103,N_12257,N_12516);
and U13104 (N_13104,N_12585,N_12525);
nand U13105 (N_13105,N_12137,N_12337);
or U13106 (N_13106,N_12189,N_12338);
nor U13107 (N_13107,N_12470,N_12652);
or U13108 (N_13108,N_12605,N_12240);
nor U13109 (N_13109,N_12519,N_12960);
nor U13110 (N_13110,N_12361,N_12493);
xnor U13111 (N_13111,N_12235,N_12929);
xnor U13112 (N_13112,N_12308,N_12386);
xnor U13113 (N_13113,N_12715,N_12122);
nand U13114 (N_13114,N_12688,N_12656);
xnor U13115 (N_13115,N_12590,N_12721);
nor U13116 (N_13116,N_12321,N_12936);
nor U13117 (N_13117,N_12896,N_12957);
nor U13118 (N_13118,N_12363,N_12180);
nand U13119 (N_13119,N_12564,N_12670);
nand U13120 (N_13120,N_12925,N_12916);
nand U13121 (N_13121,N_12709,N_12614);
xnor U13122 (N_13122,N_12791,N_12633);
nor U13123 (N_13123,N_12866,N_12823);
xnor U13124 (N_13124,N_12452,N_12219);
or U13125 (N_13125,N_12696,N_12830);
nor U13126 (N_13126,N_12097,N_12366);
or U13127 (N_13127,N_12263,N_12435);
nor U13128 (N_13128,N_12194,N_12239);
or U13129 (N_13129,N_12804,N_12289);
and U13130 (N_13130,N_12199,N_12119);
and U13131 (N_13131,N_12970,N_12392);
nor U13132 (N_13132,N_12855,N_12448);
xor U13133 (N_13133,N_12816,N_12610);
nor U13134 (N_13134,N_12305,N_12037);
and U13135 (N_13135,N_12789,N_12546);
and U13136 (N_13136,N_12410,N_12404);
and U13137 (N_13137,N_12684,N_12514);
nor U13138 (N_13138,N_12601,N_12252);
nor U13139 (N_13139,N_12988,N_12844);
or U13140 (N_13140,N_12195,N_12466);
nor U13141 (N_13141,N_12039,N_12294);
and U13142 (N_13142,N_12865,N_12874);
or U13143 (N_13143,N_12741,N_12088);
or U13144 (N_13144,N_12048,N_12649);
nand U13145 (N_13145,N_12120,N_12115);
and U13146 (N_13146,N_12813,N_12104);
or U13147 (N_13147,N_12779,N_12635);
nand U13148 (N_13148,N_12498,N_12043);
nor U13149 (N_13149,N_12598,N_12464);
and U13150 (N_13150,N_12910,N_12292);
or U13151 (N_13151,N_12227,N_12723);
nand U13152 (N_13152,N_12463,N_12077);
and U13153 (N_13153,N_12065,N_12140);
nand U13154 (N_13154,N_12754,N_12309);
nand U13155 (N_13155,N_12275,N_12360);
nand U13156 (N_13156,N_12354,N_12486);
xnor U13157 (N_13157,N_12676,N_12860);
nand U13158 (N_13158,N_12637,N_12786);
xnor U13159 (N_13159,N_12414,N_12402);
and U13160 (N_13160,N_12339,N_12439);
xnor U13161 (N_13161,N_12659,N_12164);
and U13162 (N_13162,N_12210,N_12760);
and U13163 (N_13163,N_12976,N_12249);
and U13164 (N_13164,N_12560,N_12454);
xnor U13165 (N_13165,N_12300,N_12166);
nor U13166 (N_13166,N_12350,N_12984);
xnor U13167 (N_13167,N_12556,N_12050);
nand U13168 (N_13168,N_12281,N_12524);
nand U13169 (N_13169,N_12059,N_12076);
xnor U13170 (N_13170,N_12795,N_12549);
nand U13171 (N_13171,N_12301,N_12409);
or U13172 (N_13172,N_12344,N_12325);
and U13173 (N_13173,N_12378,N_12719);
nor U13174 (N_13174,N_12801,N_12520);
nand U13175 (N_13175,N_12231,N_12870);
nand U13176 (N_13176,N_12358,N_12586);
xor U13177 (N_13177,N_12032,N_12747);
nand U13178 (N_13178,N_12228,N_12109);
xor U13179 (N_13179,N_12868,N_12935);
xnor U13180 (N_13180,N_12379,N_12863);
nand U13181 (N_13181,N_12384,N_12616);
or U13182 (N_13182,N_12617,N_12851);
or U13183 (N_13183,N_12434,N_12145);
and U13184 (N_13184,N_12995,N_12031);
nor U13185 (N_13185,N_12468,N_12615);
xnor U13186 (N_13186,N_12500,N_12512);
or U13187 (N_13187,N_12817,N_12974);
nand U13188 (N_13188,N_12359,N_12807);
or U13189 (N_13189,N_12961,N_12611);
and U13190 (N_13190,N_12752,N_12213);
or U13191 (N_13191,N_12665,N_12777);
nor U13192 (N_13192,N_12939,N_12735);
and U13193 (N_13193,N_12171,N_12604);
nor U13194 (N_13194,N_12419,N_12542);
nand U13195 (N_13195,N_12183,N_12700);
and U13196 (N_13196,N_12153,N_12158);
or U13197 (N_13197,N_12504,N_12806);
xnor U13198 (N_13198,N_12442,N_12978);
xnor U13199 (N_13199,N_12081,N_12985);
and U13200 (N_13200,N_12511,N_12803);
nand U13201 (N_13201,N_12117,N_12372);
nor U13202 (N_13202,N_12248,N_12989);
xor U13203 (N_13203,N_12458,N_12550);
xor U13204 (N_13204,N_12852,N_12027);
or U13205 (N_13205,N_12264,N_12477);
nand U13206 (N_13206,N_12757,N_12142);
or U13207 (N_13207,N_12902,N_12800);
nand U13208 (N_13208,N_12373,N_12694);
xnor U13209 (N_13209,N_12203,N_12324);
nor U13210 (N_13210,N_12557,N_12945);
and U13211 (N_13211,N_12403,N_12518);
nor U13212 (N_13212,N_12278,N_12536);
nor U13213 (N_13213,N_12768,N_12618);
nor U13214 (N_13214,N_12653,N_12440);
and U13215 (N_13215,N_12269,N_12717);
nand U13216 (N_13216,N_12206,N_12994);
xor U13217 (N_13217,N_12905,N_12770);
nand U13218 (N_13218,N_12071,N_12232);
xnor U13219 (N_13219,N_12639,N_12907);
xor U13220 (N_13220,N_12729,N_12311);
nor U13221 (N_13221,N_12646,N_12607);
nand U13222 (N_13222,N_12490,N_12133);
xnor U13223 (N_13223,N_12303,N_12332);
nor U13224 (N_13224,N_12951,N_12944);
nor U13225 (N_13225,N_12310,N_12695);
xor U13226 (N_13226,N_12950,N_12351);
nor U13227 (N_13227,N_12675,N_12983);
or U13228 (N_13228,N_12745,N_12161);
xnor U13229 (N_13229,N_12619,N_12201);
xor U13230 (N_13230,N_12038,N_12457);
or U13231 (N_13231,N_12084,N_12934);
nor U13232 (N_13232,N_12193,N_12295);
or U13233 (N_13233,N_12329,N_12450);
nor U13234 (N_13234,N_12644,N_12478);
and U13235 (N_13235,N_12955,N_12273);
nand U13236 (N_13236,N_12322,N_12444);
nand U13237 (N_13237,N_12268,N_12528);
and U13238 (N_13238,N_12815,N_12078);
nor U13239 (N_13239,N_12121,N_12132);
or U13240 (N_13240,N_12538,N_12502);
nor U13241 (N_13241,N_12623,N_12838);
nand U13242 (N_13242,N_12459,N_12010);
or U13243 (N_13243,N_12503,N_12172);
nor U13244 (N_13244,N_12170,N_12356);
nor U13245 (N_13245,N_12176,N_12836);
xor U13246 (N_13246,N_12129,N_12744);
or U13247 (N_13247,N_12689,N_12638);
nand U13248 (N_13248,N_12290,N_12612);
or U13249 (N_13249,N_12389,N_12108);
or U13250 (N_13250,N_12956,N_12952);
nor U13251 (N_13251,N_12932,N_12996);
and U13252 (N_13252,N_12776,N_12505);
and U13253 (N_13253,N_12274,N_12928);
nand U13254 (N_13254,N_12843,N_12377);
xnor U13255 (N_13255,N_12730,N_12679);
nand U13256 (N_13256,N_12283,N_12508);
nor U13257 (N_13257,N_12473,N_12123);
nand U13258 (N_13258,N_12340,N_12424);
nand U13259 (N_13259,N_12368,N_12243);
nand U13260 (N_13260,N_12981,N_12110);
and U13261 (N_13261,N_12141,N_12690);
xnor U13262 (N_13262,N_12810,N_12376);
nor U13263 (N_13263,N_12375,N_12506);
and U13264 (N_13264,N_12885,N_12061);
and U13265 (N_13265,N_12156,N_12181);
xnor U13266 (N_13266,N_12286,N_12085);
and U13267 (N_13267,N_12669,N_12044);
nor U13268 (N_13268,N_12641,N_12480);
nor U13269 (N_13269,N_12924,N_12509);
nor U13270 (N_13270,N_12891,N_12220);
and U13271 (N_13271,N_12024,N_12919);
nand U13272 (N_13272,N_12396,N_12364);
xnor U13273 (N_13273,N_12808,N_12390);
and U13274 (N_13274,N_12881,N_12415);
nor U13275 (N_13275,N_12094,N_12187);
xor U13276 (N_13276,N_12127,N_12042);
nor U13277 (N_13277,N_12580,N_12673);
or U13278 (N_13278,N_12552,N_12047);
xor U13279 (N_13279,N_12840,N_12867);
xnor U13280 (N_13280,N_12758,N_12850);
xnor U13281 (N_13281,N_12738,N_12036);
nand U13282 (N_13282,N_12712,N_12634);
nor U13283 (N_13283,N_12212,N_12908);
nor U13284 (N_13284,N_12451,N_12355);
nand U13285 (N_13285,N_12391,N_12455);
and U13286 (N_13286,N_12812,N_12242);
xnor U13287 (N_13287,N_12233,N_12096);
and U13288 (N_13288,N_12802,N_12857);
or U13289 (N_13289,N_12991,N_12421);
and U13290 (N_13290,N_12559,N_12886);
nor U13291 (N_13291,N_12785,N_12216);
nor U13292 (N_13292,N_12787,N_12058);
or U13293 (N_13293,N_12412,N_12485);
nor U13294 (N_13294,N_12630,N_12186);
nand U13295 (N_13295,N_12561,N_12887);
nor U13296 (N_13296,N_12596,N_12433);
and U13297 (N_13297,N_12159,N_12053);
or U13298 (N_13298,N_12494,N_12878);
nand U13299 (N_13299,N_12667,N_12798);
nand U13300 (N_13300,N_12083,N_12941);
and U13301 (N_13301,N_12405,N_12019);
or U13302 (N_13302,N_12664,N_12237);
or U13303 (N_13303,N_12446,N_12714);
and U13304 (N_13304,N_12262,N_12862);
or U13305 (N_13305,N_12191,N_12298);
and U13306 (N_13306,N_12553,N_12966);
and U13307 (N_13307,N_12765,N_12532);
xor U13308 (N_13308,N_12672,N_12899);
nand U13309 (N_13309,N_12099,N_12426);
nand U13310 (N_13310,N_12657,N_12319);
nand U13311 (N_13311,N_12054,N_12155);
nor U13312 (N_13312,N_12064,N_12825);
and U13313 (N_13313,N_12387,N_12353);
nor U13314 (N_13314,N_12112,N_12102);
and U13315 (N_13315,N_12953,N_12277);
nand U13316 (N_13316,N_12707,N_12015);
and U13317 (N_13317,N_12362,N_12288);
nand U13318 (N_13318,N_12148,N_12197);
nor U13319 (N_13319,N_12221,N_12692);
and U13320 (N_13320,N_12149,N_12903);
nor U13321 (N_13321,N_12128,N_12746);
and U13322 (N_13322,N_12316,N_12312);
nor U13323 (N_13323,N_12642,N_12771);
or U13324 (N_13324,N_12942,N_12581);
nor U13325 (N_13325,N_12418,N_12208);
nand U13326 (N_13326,N_12515,N_12284);
xor U13327 (N_13327,N_12241,N_12002);
nand U13328 (N_13328,N_12877,N_12369);
nor U13329 (N_13329,N_12013,N_12766);
nor U13330 (N_13330,N_12917,N_12540);
xor U13331 (N_13331,N_12914,N_12883);
nand U13332 (N_13332,N_12147,N_12783);
or U13333 (N_13333,N_12113,N_12681);
or U13334 (N_13334,N_12743,N_12713);
xor U13335 (N_13335,N_12892,N_12107);
or U13336 (N_13336,N_12106,N_12429);
nand U13337 (N_13337,N_12018,N_12841);
xor U13338 (N_13338,N_12411,N_12020);
or U13339 (N_13339,N_12276,N_12736);
xor U13340 (N_13340,N_12912,N_12211);
xnor U13341 (N_13341,N_12246,N_12904);
and U13342 (N_13342,N_12092,N_12499);
or U13343 (N_13343,N_12323,N_12901);
nand U13344 (N_13344,N_12975,N_12130);
xnor U13345 (N_13345,N_12629,N_12365);
nand U13346 (N_13346,N_12258,N_12888);
nor U13347 (N_13347,N_12114,N_12979);
nor U13348 (N_13348,N_12162,N_12150);
nor U13349 (N_13349,N_12620,N_12811);
nand U13350 (N_13350,N_12977,N_12467);
or U13351 (N_13351,N_12371,N_12055);
or U13352 (N_13352,N_12245,N_12188);
nand U13353 (N_13353,N_12261,N_12238);
xor U13354 (N_13354,N_12432,N_12571);
nand U13355 (N_13355,N_12526,N_12898);
or U13356 (N_13356,N_12640,N_12069);
or U13357 (N_13357,N_12060,N_12962);
nand U13358 (N_13358,N_12986,N_12954);
nor U13359 (N_13359,N_12650,N_12413);
nand U13360 (N_13360,N_12724,N_12270);
or U13361 (N_13361,N_12937,N_12547);
xor U13362 (N_13362,N_12834,N_12474);
or U13363 (N_13363,N_12326,N_12718);
xor U13364 (N_13364,N_12436,N_12492);
nor U13365 (N_13365,N_12827,N_12430);
or U13366 (N_13366,N_12067,N_12507);
xor U13367 (N_13367,N_12748,N_12009);
or U13368 (N_13368,N_12926,N_12388);
and U13369 (N_13369,N_12759,N_12606);
nor U13370 (N_13370,N_12693,N_12677);
nand U13371 (N_13371,N_12146,N_12160);
xnor U13372 (N_13372,N_12045,N_12182);
nand U13373 (N_13373,N_12100,N_12839);
nand U13374 (N_13374,N_12080,N_12822);
and U13375 (N_13375,N_12438,N_12762);
xor U13376 (N_13376,N_12028,N_12900);
nor U13377 (N_13377,N_12481,N_12462);
and U13378 (N_13378,N_12773,N_12138);
nand U13379 (N_13379,N_12753,N_12790);
or U13380 (N_13380,N_12196,N_12755);
nor U13381 (N_13381,N_12091,N_12666);
xnor U13382 (N_13382,N_12949,N_12603);
xnor U13383 (N_13383,N_12602,N_12535);
and U13384 (N_13384,N_12869,N_12889);
and U13385 (N_13385,N_12111,N_12875);
or U13386 (N_13386,N_12799,N_12814);
xor U13387 (N_13387,N_12399,N_12609);
nor U13388 (N_13388,N_12680,N_12691);
xor U13389 (N_13389,N_12460,N_12445);
and U13390 (N_13390,N_12214,N_12625);
nor U13391 (N_13391,N_12034,N_12207);
or U13392 (N_13392,N_12820,N_12531);
nand U13393 (N_13393,N_12200,N_12254);
and U13394 (N_13394,N_12761,N_12247);
and U13395 (N_13395,N_12654,N_12621);
xnor U13396 (N_13396,N_12482,N_12174);
xnor U13397 (N_13397,N_12597,N_12523);
nor U13398 (N_13398,N_12052,N_12225);
nor U13399 (N_13399,N_12040,N_12282);
nand U13400 (N_13400,N_12645,N_12915);
and U13401 (N_13401,N_12336,N_12202);
or U13402 (N_13402,N_12222,N_12465);
nand U13403 (N_13403,N_12472,N_12168);
xor U13404 (N_13404,N_12204,N_12072);
or U13405 (N_13405,N_12930,N_12397);
xor U13406 (N_13406,N_12933,N_12972);
nor U13407 (N_13407,N_12793,N_12070);
or U13408 (N_13408,N_12479,N_12175);
nor U13409 (N_13409,N_12990,N_12003);
xor U13410 (N_13410,N_12682,N_12999);
xor U13411 (N_13411,N_12595,N_12066);
xnor U13412 (N_13412,N_12969,N_12001);
or U13413 (N_13413,N_12705,N_12521);
or U13414 (N_13414,N_12568,N_12190);
and U13415 (N_13415,N_12090,N_12555);
nand U13416 (N_13416,N_12271,N_12809);
and U13417 (N_13417,N_12259,N_12427);
or U13418 (N_13418,N_12833,N_12911);
xor U13419 (N_13419,N_12702,N_12223);
and U13420 (N_13420,N_12818,N_12920);
xor U13421 (N_13421,N_12307,N_12447);
and U13422 (N_13422,N_12437,N_12737);
and U13423 (N_13423,N_12772,N_12285);
or U13424 (N_13424,N_12265,N_12098);
xor U13425 (N_13425,N_12017,N_12529);
nor U13426 (N_13426,N_12608,N_12893);
or U13427 (N_13427,N_12491,N_12049);
xor U13428 (N_13428,N_12592,N_12255);
nor U13429 (N_13429,N_12805,N_12835);
nor U13430 (N_13430,N_12456,N_12051);
nand U13431 (N_13431,N_12134,N_12333);
nand U13432 (N_13432,N_12683,N_12563);
and U13433 (N_13433,N_12964,N_12968);
nor U13434 (N_13434,N_12215,N_12565);
xnor U13435 (N_13435,N_12781,N_12775);
xor U13436 (N_13436,N_12685,N_12428);
or U13437 (N_13437,N_12004,N_12558);
nand U13438 (N_13438,N_12577,N_12073);
and U13439 (N_13439,N_12400,N_12461);
xor U13440 (N_13440,N_12541,N_12313);
nand U13441 (N_13441,N_12728,N_12184);
nand U13442 (N_13442,N_12296,N_12722);
or U13443 (N_13443,N_12725,N_12780);
xor U13444 (N_13444,N_12293,N_12534);
or U13445 (N_13445,N_12314,N_12513);
nand U13446 (N_13446,N_12697,N_12997);
nand U13447 (N_13447,N_12938,N_12742);
xor U13448 (N_13448,N_12348,N_12126);
nor U13449 (N_13449,N_12124,N_12871);
or U13450 (N_13450,N_12651,N_12297);
nand U13451 (N_13451,N_12726,N_12699);
xor U13452 (N_13452,N_12864,N_12782);
nand U13453 (N_13453,N_12569,N_12266);
or U13454 (N_13454,N_12422,N_12701);
xnor U13455 (N_13455,N_12420,N_12173);
and U13456 (N_13456,N_12643,N_12154);
nor U13457 (N_13457,N_12230,N_12648);
and U13458 (N_13458,N_12543,N_12517);
xor U13459 (N_13459,N_12971,N_12035);
nor U13460 (N_13460,N_12708,N_12913);
nand U13461 (N_13461,N_12469,N_12739);
nand U13462 (N_13462,N_12740,N_12381);
nand U13463 (N_13463,N_12829,N_12089);
nor U13464 (N_13464,N_12152,N_12062);
or U13465 (N_13465,N_12582,N_12769);
xor U13466 (N_13466,N_12331,N_12023);
or U13467 (N_13467,N_12703,N_12236);
nand U13468 (N_13468,N_12958,N_12489);
and U13469 (N_13469,N_12716,N_12554);
nor U13470 (N_13470,N_12824,N_12291);
or U13471 (N_13471,N_12575,N_12253);
or U13472 (N_13472,N_12998,N_12401);
or U13473 (N_13473,N_12475,N_12987);
nand U13474 (N_13474,N_12923,N_12087);
and U13475 (N_13475,N_12209,N_12894);
and U13476 (N_13476,N_12163,N_12895);
nand U13477 (N_13477,N_12063,N_12921);
and U13478 (N_13478,N_12720,N_12594);
or U13479 (N_13479,N_12853,N_12495);
or U13480 (N_13480,N_12014,N_12756);
nand U13481 (N_13481,N_12476,N_12658);
or U13482 (N_13482,N_12510,N_12522);
or U13483 (N_13483,N_12169,N_12533);
and U13484 (N_13484,N_12613,N_12624);
xnor U13485 (N_13485,N_12796,N_12849);
or U13486 (N_13486,N_12394,N_12136);
xnor U13487 (N_13487,N_12831,N_12343);
nor U13488 (N_13488,N_12218,N_12588);
or U13489 (N_13489,N_12131,N_12118);
nor U13490 (N_13490,N_12030,N_12453);
nor U13491 (N_13491,N_12393,N_12794);
or U13492 (N_13492,N_12347,N_12710);
nor U13493 (N_13493,N_12732,N_12882);
or U13494 (N_13494,N_12584,N_12848);
nor U13495 (N_13495,N_12280,N_12443);
and U13496 (N_13496,N_12165,N_12068);
xor U13497 (N_13497,N_12385,N_12854);
nor U13498 (N_13498,N_12025,N_12256);
nor U13499 (N_13499,N_12346,N_12727);
or U13500 (N_13500,N_12767,N_12377);
nand U13501 (N_13501,N_12109,N_12537);
or U13502 (N_13502,N_12250,N_12314);
nand U13503 (N_13503,N_12787,N_12959);
xnor U13504 (N_13504,N_12737,N_12729);
and U13505 (N_13505,N_12729,N_12687);
xor U13506 (N_13506,N_12057,N_12426);
xnor U13507 (N_13507,N_12934,N_12250);
or U13508 (N_13508,N_12735,N_12873);
nand U13509 (N_13509,N_12839,N_12929);
or U13510 (N_13510,N_12062,N_12224);
xor U13511 (N_13511,N_12504,N_12948);
and U13512 (N_13512,N_12113,N_12459);
nand U13513 (N_13513,N_12187,N_12250);
or U13514 (N_13514,N_12159,N_12418);
and U13515 (N_13515,N_12585,N_12322);
or U13516 (N_13516,N_12676,N_12093);
nor U13517 (N_13517,N_12347,N_12940);
nand U13518 (N_13518,N_12552,N_12615);
xor U13519 (N_13519,N_12155,N_12971);
or U13520 (N_13520,N_12257,N_12071);
xor U13521 (N_13521,N_12872,N_12140);
xor U13522 (N_13522,N_12744,N_12727);
and U13523 (N_13523,N_12361,N_12589);
and U13524 (N_13524,N_12467,N_12777);
nor U13525 (N_13525,N_12077,N_12701);
or U13526 (N_13526,N_12098,N_12908);
xnor U13527 (N_13527,N_12163,N_12499);
or U13528 (N_13528,N_12879,N_12797);
xnor U13529 (N_13529,N_12105,N_12175);
or U13530 (N_13530,N_12364,N_12300);
or U13531 (N_13531,N_12127,N_12093);
xnor U13532 (N_13532,N_12081,N_12149);
xor U13533 (N_13533,N_12029,N_12141);
and U13534 (N_13534,N_12125,N_12315);
nor U13535 (N_13535,N_12547,N_12383);
and U13536 (N_13536,N_12172,N_12920);
or U13537 (N_13537,N_12403,N_12342);
xor U13538 (N_13538,N_12203,N_12211);
xnor U13539 (N_13539,N_12914,N_12162);
nand U13540 (N_13540,N_12961,N_12667);
nand U13541 (N_13541,N_12030,N_12245);
nand U13542 (N_13542,N_12626,N_12739);
nor U13543 (N_13543,N_12889,N_12430);
or U13544 (N_13544,N_12770,N_12121);
nand U13545 (N_13545,N_12836,N_12541);
nor U13546 (N_13546,N_12677,N_12901);
nor U13547 (N_13547,N_12826,N_12621);
nor U13548 (N_13548,N_12671,N_12383);
and U13549 (N_13549,N_12333,N_12614);
xor U13550 (N_13550,N_12101,N_12128);
or U13551 (N_13551,N_12115,N_12513);
nor U13552 (N_13552,N_12783,N_12473);
nor U13553 (N_13553,N_12307,N_12840);
or U13554 (N_13554,N_12987,N_12422);
xnor U13555 (N_13555,N_12999,N_12988);
nand U13556 (N_13556,N_12348,N_12489);
nor U13557 (N_13557,N_12122,N_12259);
or U13558 (N_13558,N_12420,N_12775);
and U13559 (N_13559,N_12105,N_12860);
xor U13560 (N_13560,N_12571,N_12799);
nor U13561 (N_13561,N_12786,N_12525);
xor U13562 (N_13562,N_12354,N_12330);
nor U13563 (N_13563,N_12039,N_12195);
nand U13564 (N_13564,N_12985,N_12253);
and U13565 (N_13565,N_12120,N_12283);
nor U13566 (N_13566,N_12024,N_12097);
nand U13567 (N_13567,N_12177,N_12307);
xnor U13568 (N_13568,N_12283,N_12802);
or U13569 (N_13569,N_12010,N_12780);
xor U13570 (N_13570,N_12488,N_12395);
xor U13571 (N_13571,N_12165,N_12296);
or U13572 (N_13572,N_12492,N_12096);
and U13573 (N_13573,N_12909,N_12906);
xor U13574 (N_13574,N_12004,N_12427);
nand U13575 (N_13575,N_12598,N_12551);
nand U13576 (N_13576,N_12565,N_12345);
xnor U13577 (N_13577,N_12985,N_12837);
xnor U13578 (N_13578,N_12397,N_12016);
or U13579 (N_13579,N_12515,N_12226);
or U13580 (N_13580,N_12768,N_12240);
nor U13581 (N_13581,N_12161,N_12239);
or U13582 (N_13582,N_12816,N_12890);
nand U13583 (N_13583,N_12694,N_12600);
or U13584 (N_13584,N_12368,N_12464);
and U13585 (N_13585,N_12804,N_12419);
nand U13586 (N_13586,N_12381,N_12069);
nor U13587 (N_13587,N_12285,N_12572);
xor U13588 (N_13588,N_12243,N_12046);
nand U13589 (N_13589,N_12032,N_12594);
or U13590 (N_13590,N_12767,N_12890);
nor U13591 (N_13591,N_12287,N_12554);
nand U13592 (N_13592,N_12947,N_12528);
nor U13593 (N_13593,N_12587,N_12150);
nand U13594 (N_13594,N_12781,N_12048);
xnor U13595 (N_13595,N_12796,N_12452);
xor U13596 (N_13596,N_12199,N_12650);
xnor U13597 (N_13597,N_12651,N_12534);
or U13598 (N_13598,N_12715,N_12453);
nor U13599 (N_13599,N_12583,N_12614);
nand U13600 (N_13600,N_12497,N_12619);
nor U13601 (N_13601,N_12762,N_12827);
and U13602 (N_13602,N_12513,N_12803);
nor U13603 (N_13603,N_12066,N_12985);
nand U13604 (N_13604,N_12721,N_12127);
xor U13605 (N_13605,N_12201,N_12419);
and U13606 (N_13606,N_12857,N_12009);
nor U13607 (N_13607,N_12424,N_12890);
xor U13608 (N_13608,N_12154,N_12838);
xor U13609 (N_13609,N_12856,N_12022);
xnor U13610 (N_13610,N_12876,N_12115);
xor U13611 (N_13611,N_12648,N_12169);
xor U13612 (N_13612,N_12957,N_12505);
and U13613 (N_13613,N_12076,N_12711);
xor U13614 (N_13614,N_12241,N_12015);
or U13615 (N_13615,N_12708,N_12109);
nand U13616 (N_13616,N_12972,N_12672);
nand U13617 (N_13617,N_12904,N_12175);
and U13618 (N_13618,N_12945,N_12617);
nand U13619 (N_13619,N_12560,N_12992);
or U13620 (N_13620,N_12529,N_12748);
or U13621 (N_13621,N_12057,N_12805);
and U13622 (N_13622,N_12476,N_12509);
nor U13623 (N_13623,N_12487,N_12114);
or U13624 (N_13624,N_12705,N_12632);
nand U13625 (N_13625,N_12225,N_12762);
nor U13626 (N_13626,N_12750,N_12623);
nand U13627 (N_13627,N_12977,N_12055);
nor U13628 (N_13628,N_12140,N_12627);
xor U13629 (N_13629,N_12162,N_12449);
and U13630 (N_13630,N_12864,N_12416);
nand U13631 (N_13631,N_12196,N_12749);
xor U13632 (N_13632,N_12724,N_12702);
or U13633 (N_13633,N_12493,N_12022);
nor U13634 (N_13634,N_12226,N_12575);
and U13635 (N_13635,N_12288,N_12978);
nand U13636 (N_13636,N_12136,N_12779);
nand U13637 (N_13637,N_12612,N_12388);
xnor U13638 (N_13638,N_12562,N_12595);
xnor U13639 (N_13639,N_12937,N_12333);
and U13640 (N_13640,N_12378,N_12307);
xnor U13641 (N_13641,N_12891,N_12082);
nand U13642 (N_13642,N_12117,N_12690);
and U13643 (N_13643,N_12616,N_12925);
nand U13644 (N_13644,N_12384,N_12913);
nor U13645 (N_13645,N_12053,N_12555);
nand U13646 (N_13646,N_12955,N_12304);
nand U13647 (N_13647,N_12349,N_12904);
and U13648 (N_13648,N_12142,N_12680);
and U13649 (N_13649,N_12246,N_12696);
and U13650 (N_13650,N_12219,N_12792);
nor U13651 (N_13651,N_12731,N_12314);
or U13652 (N_13652,N_12941,N_12789);
xnor U13653 (N_13653,N_12505,N_12450);
xnor U13654 (N_13654,N_12009,N_12265);
xor U13655 (N_13655,N_12397,N_12754);
xor U13656 (N_13656,N_12792,N_12503);
xnor U13657 (N_13657,N_12759,N_12936);
or U13658 (N_13658,N_12882,N_12041);
xnor U13659 (N_13659,N_12998,N_12492);
and U13660 (N_13660,N_12449,N_12335);
or U13661 (N_13661,N_12016,N_12021);
nand U13662 (N_13662,N_12076,N_12702);
or U13663 (N_13663,N_12753,N_12914);
or U13664 (N_13664,N_12079,N_12958);
nand U13665 (N_13665,N_12439,N_12763);
xnor U13666 (N_13666,N_12050,N_12797);
or U13667 (N_13667,N_12715,N_12875);
xnor U13668 (N_13668,N_12892,N_12172);
or U13669 (N_13669,N_12585,N_12803);
nor U13670 (N_13670,N_12213,N_12114);
nand U13671 (N_13671,N_12430,N_12413);
and U13672 (N_13672,N_12409,N_12932);
nand U13673 (N_13673,N_12981,N_12220);
or U13674 (N_13674,N_12645,N_12565);
nor U13675 (N_13675,N_12934,N_12579);
or U13676 (N_13676,N_12199,N_12618);
and U13677 (N_13677,N_12286,N_12335);
xor U13678 (N_13678,N_12260,N_12363);
nor U13679 (N_13679,N_12954,N_12898);
and U13680 (N_13680,N_12536,N_12227);
or U13681 (N_13681,N_12551,N_12451);
xnor U13682 (N_13682,N_12744,N_12230);
xor U13683 (N_13683,N_12423,N_12166);
nor U13684 (N_13684,N_12784,N_12198);
xnor U13685 (N_13685,N_12095,N_12428);
nor U13686 (N_13686,N_12840,N_12285);
and U13687 (N_13687,N_12850,N_12207);
xnor U13688 (N_13688,N_12703,N_12024);
or U13689 (N_13689,N_12469,N_12253);
nand U13690 (N_13690,N_12586,N_12415);
nand U13691 (N_13691,N_12961,N_12257);
nand U13692 (N_13692,N_12867,N_12819);
and U13693 (N_13693,N_12998,N_12844);
nor U13694 (N_13694,N_12867,N_12187);
and U13695 (N_13695,N_12198,N_12881);
xor U13696 (N_13696,N_12319,N_12336);
nor U13697 (N_13697,N_12070,N_12230);
nand U13698 (N_13698,N_12339,N_12317);
xor U13699 (N_13699,N_12058,N_12342);
nand U13700 (N_13700,N_12891,N_12321);
or U13701 (N_13701,N_12409,N_12774);
nand U13702 (N_13702,N_12310,N_12951);
and U13703 (N_13703,N_12704,N_12139);
or U13704 (N_13704,N_12728,N_12992);
xnor U13705 (N_13705,N_12947,N_12711);
and U13706 (N_13706,N_12983,N_12766);
xnor U13707 (N_13707,N_12130,N_12911);
xor U13708 (N_13708,N_12019,N_12990);
or U13709 (N_13709,N_12581,N_12477);
or U13710 (N_13710,N_12025,N_12188);
nand U13711 (N_13711,N_12601,N_12171);
xor U13712 (N_13712,N_12713,N_12020);
xor U13713 (N_13713,N_12868,N_12172);
and U13714 (N_13714,N_12564,N_12131);
nand U13715 (N_13715,N_12931,N_12726);
nand U13716 (N_13716,N_12992,N_12231);
xor U13717 (N_13717,N_12469,N_12204);
and U13718 (N_13718,N_12583,N_12797);
or U13719 (N_13719,N_12100,N_12586);
and U13720 (N_13720,N_12645,N_12438);
or U13721 (N_13721,N_12567,N_12383);
xnor U13722 (N_13722,N_12448,N_12946);
and U13723 (N_13723,N_12319,N_12232);
and U13724 (N_13724,N_12316,N_12009);
xnor U13725 (N_13725,N_12853,N_12199);
and U13726 (N_13726,N_12889,N_12739);
nand U13727 (N_13727,N_12517,N_12666);
nor U13728 (N_13728,N_12712,N_12658);
xnor U13729 (N_13729,N_12414,N_12740);
xnor U13730 (N_13730,N_12658,N_12949);
xor U13731 (N_13731,N_12846,N_12106);
and U13732 (N_13732,N_12411,N_12647);
nand U13733 (N_13733,N_12420,N_12344);
or U13734 (N_13734,N_12940,N_12509);
and U13735 (N_13735,N_12680,N_12135);
and U13736 (N_13736,N_12997,N_12747);
xnor U13737 (N_13737,N_12507,N_12647);
xnor U13738 (N_13738,N_12034,N_12940);
nand U13739 (N_13739,N_12366,N_12226);
xnor U13740 (N_13740,N_12556,N_12262);
nand U13741 (N_13741,N_12537,N_12942);
xor U13742 (N_13742,N_12022,N_12968);
and U13743 (N_13743,N_12200,N_12974);
nor U13744 (N_13744,N_12012,N_12840);
and U13745 (N_13745,N_12899,N_12755);
and U13746 (N_13746,N_12238,N_12396);
and U13747 (N_13747,N_12190,N_12597);
and U13748 (N_13748,N_12396,N_12070);
xnor U13749 (N_13749,N_12086,N_12072);
and U13750 (N_13750,N_12733,N_12373);
xor U13751 (N_13751,N_12303,N_12518);
nor U13752 (N_13752,N_12945,N_12714);
nor U13753 (N_13753,N_12805,N_12871);
xnor U13754 (N_13754,N_12274,N_12578);
nand U13755 (N_13755,N_12799,N_12880);
and U13756 (N_13756,N_12256,N_12721);
nor U13757 (N_13757,N_12329,N_12500);
and U13758 (N_13758,N_12435,N_12581);
or U13759 (N_13759,N_12269,N_12913);
and U13760 (N_13760,N_12968,N_12613);
and U13761 (N_13761,N_12348,N_12012);
xnor U13762 (N_13762,N_12024,N_12634);
and U13763 (N_13763,N_12297,N_12684);
nand U13764 (N_13764,N_12388,N_12968);
and U13765 (N_13765,N_12123,N_12102);
xor U13766 (N_13766,N_12031,N_12362);
or U13767 (N_13767,N_12077,N_12335);
or U13768 (N_13768,N_12853,N_12010);
xor U13769 (N_13769,N_12526,N_12755);
xor U13770 (N_13770,N_12492,N_12170);
xor U13771 (N_13771,N_12299,N_12669);
or U13772 (N_13772,N_12585,N_12415);
or U13773 (N_13773,N_12216,N_12125);
xnor U13774 (N_13774,N_12970,N_12789);
or U13775 (N_13775,N_12900,N_12295);
and U13776 (N_13776,N_12212,N_12913);
xnor U13777 (N_13777,N_12789,N_12000);
nor U13778 (N_13778,N_12832,N_12238);
xnor U13779 (N_13779,N_12792,N_12972);
and U13780 (N_13780,N_12538,N_12162);
and U13781 (N_13781,N_12011,N_12228);
nor U13782 (N_13782,N_12893,N_12774);
nor U13783 (N_13783,N_12128,N_12476);
or U13784 (N_13784,N_12687,N_12790);
and U13785 (N_13785,N_12226,N_12701);
or U13786 (N_13786,N_12865,N_12924);
nand U13787 (N_13787,N_12041,N_12047);
xor U13788 (N_13788,N_12572,N_12529);
nand U13789 (N_13789,N_12455,N_12335);
or U13790 (N_13790,N_12220,N_12200);
nand U13791 (N_13791,N_12705,N_12469);
xor U13792 (N_13792,N_12978,N_12715);
nor U13793 (N_13793,N_12985,N_12481);
or U13794 (N_13794,N_12802,N_12161);
xnor U13795 (N_13795,N_12503,N_12057);
or U13796 (N_13796,N_12248,N_12785);
xnor U13797 (N_13797,N_12780,N_12245);
or U13798 (N_13798,N_12587,N_12129);
or U13799 (N_13799,N_12670,N_12038);
xor U13800 (N_13800,N_12241,N_12216);
and U13801 (N_13801,N_12835,N_12636);
nand U13802 (N_13802,N_12751,N_12490);
nand U13803 (N_13803,N_12069,N_12243);
nand U13804 (N_13804,N_12305,N_12682);
or U13805 (N_13805,N_12270,N_12542);
nor U13806 (N_13806,N_12719,N_12221);
xor U13807 (N_13807,N_12434,N_12398);
and U13808 (N_13808,N_12732,N_12966);
nand U13809 (N_13809,N_12768,N_12821);
nand U13810 (N_13810,N_12822,N_12879);
nor U13811 (N_13811,N_12901,N_12907);
nor U13812 (N_13812,N_12283,N_12618);
or U13813 (N_13813,N_12905,N_12346);
nand U13814 (N_13814,N_12665,N_12795);
nand U13815 (N_13815,N_12056,N_12588);
and U13816 (N_13816,N_12573,N_12250);
xor U13817 (N_13817,N_12806,N_12201);
and U13818 (N_13818,N_12487,N_12219);
or U13819 (N_13819,N_12621,N_12949);
nor U13820 (N_13820,N_12865,N_12910);
or U13821 (N_13821,N_12155,N_12127);
nor U13822 (N_13822,N_12232,N_12197);
nand U13823 (N_13823,N_12714,N_12858);
nand U13824 (N_13824,N_12636,N_12642);
or U13825 (N_13825,N_12230,N_12326);
and U13826 (N_13826,N_12060,N_12745);
nor U13827 (N_13827,N_12652,N_12693);
nand U13828 (N_13828,N_12739,N_12088);
nor U13829 (N_13829,N_12669,N_12736);
or U13830 (N_13830,N_12541,N_12710);
or U13831 (N_13831,N_12058,N_12201);
nor U13832 (N_13832,N_12011,N_12640);
and U13833 (N_13833,N_12525,N_12325);
and U13834 (N_13834,N_12780,N_12074);
xnor U13835 (N_13835,N_12256,N_12399);
xor U13836 (N_13836,N_12215,N_12442);
nor U13837 (N_13837,N_12873,N_12766);
nor U13838 (N_13838,N_12925,N_12094);
or U13839 (N_13839,N_12667,N_12819);
nand U13840 (N_13840,N_12215,N_12898);
nor U13841 (N_13841,N_12667,N_12111);
nor U13842 (N_13842,N_12366,N_12919);
or U13843 (N_13843,N_12521,N_12041);
and U13844 (N_13844,N_12841,N_12338);
xnor U13845 (N_13845,N_12401,N_12034);
and U13846 (N_13846,N_12394,N_12828);
nand U13847 (N_13847,N_12224,N_12427);
and U13848 (N_13848,N_12452,N_12877);
or U13849 (N_13849,N_12698,N_12765);
or U13850 (N_13850,N_12278,N_12533);
and U13851 (N_13851,N_12173,N_12914);
xor U13852 (N_13852,N_12188,N_12151);
nor U13853 (N_13853,N_12447,N_12073);
and U13854 (N_13854,N_12596,N_12041);
nand U13855 (N_13855,N_12244,N_12177);
and U13856 (N_13856,N_12571,N_12113);
or U13857 (N_13857,N_12127,N_12708);
or U13858 (N_13858,N_12418,N_12941);
or U13859 (N_13859,N_12916,N_12057);
nor U13860 (N_13860,N_12334,N_12437);
xnor U13861 (N_13861,N_12472,N_12146);
or U13862 (N_13862,N_12438,N_12659);
or U13863 (N_13863,N_12411,N_12167);
or U13864 (N_13864,N_12996,N_12323);
and U13865 (N_13865,N_12144,N_12378);
or U13866 (N_13866,N_12739,N_12903);
and U13867 (N_13867,N_12341,N_12281);
nand U13868 (N_13868,N_12290,N_12911);
nand U13869 (N_13869,N_12646,N_12450);
or U13870 (N_13870,N_12285,N_12924);
and U13871 (N_13871,N_12559,N_12050);
xor U13872 (N_13872,N_12712,N_12209);
nor U13873 (N_13873,N_12582,N_12610);
and U13874 (N_13874,N_12289,N_12120);
or U13875 (N_13875,N_12143,N_12839);
nor U13876 (N_13876,N_12524,N_12737);
nand U13877 (N_13877,N_12116,N_12451);
and U13878 (N_13878,N_12111,N_12022);
xnor U13879 (N_13879,N_12431,N_12188);
or U13880 (N_13880,N_12040,N_12426);
nor U13881 (N_13881,N_12295,N_12747);
and U13882 (N_13882,N_12558,N_12644);
xor U13883 (N_13883,N_12426,N_12258);
or U13884 (N_13884,N_12829,N_12002);
nand U13885 (N_13885,N_12389,N_12544);
and U13886 (N_13886,N_12821,N_12102);
or U13887 (N_13887,N_12790,N_12533);
nand U13888 (N_13888,N_12025,N_12663);
and U13889 (N_13889,N_12453,N_12716);
xor U13890 (N_13890,N_12930,N_12956);
or U13891 (N_13891,N_12826,N_12050);
nand U13892 (N_13892,N_12957,N_12640);
and U13893 (N_13893,N_12714,N_12378);
or U13894 (N_13894,N_12366,N_12247);
xor U13895 (N_13895,N_12105,N_12188);
xnor U13896 (N_13896,N_12516,N_12400);
or U13897 (N_13897,N_12697,N_12879);
nand U13898 (N_13898,N_12602,N_12743);
or U13899 (N_13899,N_12543,N_12844);
or U13900 (N_13900,N_12399,N_12384);
nor U13901 (N_13901,N_12185,N_12087);
nand U13902 (N_13902,N_12364,N_12595);
nor U13903 (N_13903,N_12089,N_12159);
and U13904 (N_13904,N_12872,N_12549);
xor U13905 (N_13905,N_12621,N_12718);
xor U13906 (N_13906,N_12328,N_12158);
and U13907 (N_13907,N_12507,N_12910);
nand U13908 (N_13908,N_12229,N_12134);
or U13909 (N_13909,N_12290,N_12331);
nand U13910 (N_13910,N_12018,N_12825);
nand U13911 (N_13911,N_12300,N_12994);
or U13912 (N_13912,N_12389,N_12353);
and U13913 (N_13913,N_12978,N_12626);
or U13914 (N_13914,N_12928,N_12218);
and U13915 (N_13915,N_12531,N_12292);
nand U13916 (N_13916,N_12482,N_12798);
nor U13917 (N_13917,N_12655,N_12216);
or U13918 (N_13918,N_12820,N_12543);
or U13919 (N_13919,N_12547,N_12251);
or U13920 (N_13920,N_12357,N_12387);
or U13921 (N_13921,N_12958,N_12580);
nand U13922 (N_13922,N_12003,N_12094);
nor U13923 (N_13923,N_12949,N_12014);
or U13924 (N_13924,N_12502,N_12584);
or U13925 (N_13925,N_12309,N_12173);
and U13926 (N_13926,N_12690,N_12866);
nor U13927 (N_13927,N_12272,N_12759);
nor U13928 (N_13928,N_12738,N_12298);
nand U13929 (N_13929,N_12195,N_12349);
or U13930 (N_13930,N_12026,N_12183);
nor U13931 (N_13931,N_12249,N_12309);
nor U13932 (N_13932,N_12840,N_12224);
or U13933 (N_13933,N_12208,N_12967);
and U13934 (N_13934,N_12908,N_12509);
nand U13935 (N_13935,N_12998,N_12982);
and U13936 (N_13936,N_12446,N_12274);
nor U13937 (N_13937,N_12589,N_12935);
nor U13938 (N_13938,N_12614,N_12650);
xor U13939 (N_13939,N_12364,N_12914);
nor U13940 (N_13940,N_12603,N_12863);
nand U13941 (N_13941,N_12720,N_12534);
xor U13942 (N_13942,N_12947,N_12488);
nor U13943 (N_13943,N_12148,N_12377);
nor U13944 (N_13944,N_12986,N_12205);
xnor U13945 (N_13945,N_12477,N_12064);
nor U13946 (N_13946,N_12411,N_12495);
nor U13947 (N_13947,N_12154,N_12585);
xor U13948 (N_13948,N_12260,N_12479);
or U13949 (N_13949,N_12337,N_12779);
or U13950 (N_13950,N_12921,N_12966);
nand U13951 (N_13951,N_12409,N_12436);
nor U13952 (N_13952,N_12637,N_12699);
xnor U13953 (N_13953,N_12660,N_12349);
nor U13954 (N_13954,N_12975,N_12375);
xnor U13955 (N_13955,N_12873,N_12902);
nand U13956 (N_13956,N_12854,N_12706);
and U13957 (N_13957,N_12097,N_12793);
or U13958 (N_13958,N_12015,N_12709);
xor U13959 (N_13959,N_12950,N_12990);
nor U13960 (N_13960,N_12448,N_12366);
nor U13961 (N_13961,N_12334,N_12253);
nand U13962 (N_13962,N_12181,N_12577);
nand U13963 (N_13963,N_12643,N_12720);
and U13964 (N_13964,N_12943,N_12900);
nand U13965 (N_13965,N_12766,N_12447);
nand U13966 (N_13966,N_12532,N_12227);
or U13967 (N_13967,N_12870,N_12529);
and U13968 (N_13968,N_12745,N_12458);
nand U13969 (N_13969,N_12236,N_12870);
and U13970 (N_13970,N_12515,N_12428);
or U13971 (N_13971,N_12009,N_12183);
xnor U13972 (N_13972,N_12527,N_12342);
and U13973 (N_13973,N_12959,N_12487);
xnor U13974 (N_13974,N_12671,N_12754);
and U13975 (N_13975,N_12060,N_12969);
nor U13976 (N_13976,N_12247,N_12081);
or U13977 (N_13977,N_12809,N_12794);
and U13978 (N_13978,N_12131,N_12561);
nor U13979 (N_13979,N_12628,N_12572);
nand U13980 (N_13980,N_12933,N_12642);
nor U13981 (N_13981,N_12068,N_12674);
nor U13982 (N_13982,N_12649,N_12390);
nand U13983 (N_13983,N_12105,N_12334);
or U13984 (N_13984,N_12407,N_12917);
nand U13985 (N_13985,N_12879,N_12937);
nor U13986 (N_13986,N_12026,N_12343);
nand U13987 (N_13987,N_12420,N_12593);
nand U13988 (N_13988,N_12360,N_12143);
xor U13989 (N_13989,N_12886,N_12330);
nor U13990 (N_13990,N_12829,N_12253);
nor U13991 (N_13991,N_12735,N_12053);
xor U13992 (N_13992,N_12388,N_12647);
xnor U13993 (N_13993,N_12232,N_12867);
and U13994 (N_13994,N_12233,N_12564);
or U13995 (N_13995,N_12723,N_12811);
xnor U13996 (N_13996,N_12264,N_12473);
and U13997 (N_13997,N_12777,N_12573);
and U13998 (N_13998,N_12522,N_12034);
and U13999 (N_13999,N_12540,N_12313);
nand U14000 (N_14000,N_13827,N_13832);
nand U14001 (N_14001,N_13410,N_13192);
nand U14002 (N_14002,N_13783,N_13455);
xor U14003 (N_14003,N_13203,N_13684);
or U14004 (N_14004,N_13439,N_13599);
xnor U14005 (N_14005,N_13826,N_13596);
xor U14006 (N_14006,N_13349,N_13677);
and U14007 (N_14007,N_13295,N_13938);
and U14008 (N_14008,N_13634,N_13504);
xor U14009 (N_14009,N_13889,N_13104);
nor U14010 (N_14010,N_13785,N_13760);
nor U14011 (N_14011,N_13285,N_13324);
xor U14012 (N_14012,N_13965,N_13664);
or U14013 (N_14013,N_13071,N_13120);
or U14014 (N_14014,N_13305,N_13655);
nor U14015 (N_14015,N_13541,N_13395);
and U14016 (N_14016,N_13500,N_13091);
nor U14017 (N_14017,N_13121,N_13625);
and U14018 (N_14018,N_13987,N_13834);
or U14019 (N_14019,N_13698,N_13062);
and U14020 (N_14020,N_13372,N_13802);
nand U14021 (N_14021,N_13964,N_13266);
and U14022 (N_14022,N_13034,N_13241);
nor U14023 (N_14023,N_13958,N_13069);
or U14024 (N_14024,N_13301,N_13738);
nor U14025 (N_14025,N_13079,N_13097);
and U14026 (N_14026,N_13982,N_13822);
xnor U14027 (N_14027,N_13323,N_13004);
and U14028 (N_14028,N_13530,N_13752);
and U14029 (N_14029,N_13540,N_13066);
or U14030 (N_14030,N_13138,N_13099);
nand U14031 (N_14031,N_13607,N_13119);
xor U14032 (N_14032,N_13576,N_13011);
or U14033 (N_14033,N_13458,N_13446);
nand U14034 (N_14034,N_13691,N_13812);
xnor U14035 (N_14035,N_13151,N_13952);
nor U14036 (N_14036,N_13989,N_13934);
and U14037 (N_14037,N_13719,N_13311);
nand U14038 (N_14038,N_13152,N_13978);
nor U14039 (N_14039,N_13378,N_13114);
or U14040 (N_14040,N_13058,N_13532);
or U14041 (N_14041,N_13472,N_13307);
and U14042 (N_14042,N_13954,N_13514);
or U14043 (N_14043,N_13581,N_13352);
xor U14044 (N_14044,N_13489,N_13407);
or U14045 (N_14045,N_13523,N_13915);
xor U14046 (N_14046,N_13125,N_13594);
nand U14047 (N_14047,N_13981,N_13588);
xnor U14048 (N_14048,N_13695,N_13375);
nand U14049 (N_14049,N_13267,N_13992);
and U14050 (N_14050,N_13923,N_13354);
nor U14051 (N_14051,N_13927,N_13746);
and U14052 (N_14052,N_13046,N_13436);
nand U14053 (N_14053,N_13328,N_13479);
or U14054 (N_14054,N_13515,N_13419);
or U14055 (N_14055,N_13309,N_13426);
nand U14056 (N_14056,N_13284,N_13363);
or U14057 (N_14057,N_13278,N_13556);
nand U14058 (N_14058,N_13127,N_13142);
xnor U14059 (N_14059,N_13632,N_13757);
nand U14060 (N_14060,N_13068,N_13396);
nor U14061 (N_14061,N_13628,N_13067);
and U14062 (N_14062,N_13296,N_13341);
nor U14063 (N_14063,N_13545,N_13497);
and U14064 (N_14064,N_13254,N_13230);
and U14065 (N_14065,N_13941,N_13379);
or U14066 (N_14066,N_13770,N_13997);
nor U14067 (N_14067,N_13320,N_13245);
or U14068 (N_14068,N_13830,N_13543);
xor U14069 (N_14069,N_13766,N_13031);
xor U14070 (N_14070,N_13551,N_13806);
and U14071 (N_14071,N_13809,N_13158);
or U14072 (N_14072,N_13999,N_13587);
and U14073 (N_14073,N_13200,N_13567);
nand U14074 (N_14074,N_13389,N_13275);
or U14075 (N_14075,N_13351,N_13271);
or U14076 (N_14076,N_13668,N_13956);
or U14077 (N_14077,N_13174,N_13761);
xor U14078 (N_14078,N_13331,N_13998);
or U14079 (N_14079,N_13603,N_13697);
nor U14080 (N_14080,N_13733,N_13844);
and U14081 (N_14081,N_13539,N_13346);
nor U14082 (N_14082,N_13641,N_13926);
nand U14083 (N_14083,N_13913,N_13401);
nor U14084 (N_14084,N_13197,N_13135);
and U14085 (N_14085,N_13525,N_13358);
xor U14086 (N_14086,N_13793,N_13780);
nand U14087 (N_14087,N_13038,N_13442);
nor U14088 (N_14088,N_13018,N_13712);
or U14089 (N_14089,N_13850,N_13888);
or U14090 (N_14090,N_13350,N_13048);
xnor U14091 (N_14091,N_13299,N_13036);
or U14092 (N_14092,N_13165,N_13824);
or U14093 (N_14093,N_13459,N_13434);
nor U14094 (N_14094,N_13220,N_13006);
or U14095 (N_14095,N_13088,N_13409);
xnor U14096 (N_14096,N_13688,N_13858);
and U14097 (N_14097,N_13199,N_13357);
nor U14098 (N_14098,N_13189,N_13518);
and U14099 (N_14099,N_13593,N_13003);
or U14100 (N_14100,N_13529,N_13669);
nand U14101 (N_14101,N_13232,N_13950);
or U14102 (N_14102,N_13920,N_13304);
nand U14103 (N_14103,N_13849,N_13526);
or U14104 (N_14104,N_13654,N_13861);
nand U14105 (N_14105,N_13914,N_13155);
nand U14106 (N_14106,N_13276,N_13162);
nor U14107 (N_14107,N_13799,N_13408);
nand U14108 (N_14108,N_13621,N_13970);
nor U14109 (N_14109,N_13423,N_13393);
xnor U14110 (N_14110,N_13916,N_13743);
nor U14111 (N_14111,N_13933,N_13268);
xor U14112 (N_14112,N_13390,N_13381);
nand U14113 (N_14113,N_13565,N_13671);
and U14114 (N_14114,N_13166,N_13139);
and U14115 (N_14115,N_13601,N_13921);
or U14116 (N_14116,N_13107,N_13869);
xnor U14117 (N_14117,N_13716,N_13623);
nor U14118 (N_14118,N_13430,N_13290);
and U14119 (N_14119,N_13602,N_13486);
xor U14120 (N_14120,N_13385,N_13728);
xor U14121 (N_14121,N_13878,N_13115);
nand U14122 (N_14122,N_13993,N_13772);
nand U14123 (N_14123,N_13735,N_13511);
and U14124 (N_14124,N_13293,N_13510);
nor U14125 (N_14125,N_13703,N_13546);
or U14126 (N_14126,N_13949,N_13150);
or U14127 (N_14127,N_13575,N_13055);
or U14128 (N_14128,N_13624,N_13076);
nor U14129 (N_14129,N_13428,N_13507);
and U14130 (N_14130,N_13364,N_13635);
or U14131 (N_14131,N_13403,N_13481);
and U14132 (N_14132,N_13202,N_13476);
xor U14133 (N_14133,N_13386,N_13231);
and U14134 (N_14134,N_13741,N_13771);
nor U14135 (N_14135,N_13857,N_13347);
nand U14136 (N_14136,N_13219,N_13633);
nor U14137 (N_14137,N_13883,N_13718);
xor U14138 (N_14138,N_13534,N_13140);
nand U14139 (N_14139,N_13056,N_13815);
nand U14140 (N_14140,N_13533,N_13294);
xor U14141 (N_14141,N_13035,N_13249);
and U14142 (N_14142,N_13144,N_13573);
or U14143 (N_14143,N_13255,N_13429);
or U14144 (N_14144,N_13404,N_13397);
nor U14145 (N_14145,N_13637,N_13008);
xor U14146 (N_14146,N_13494,N_13418);
xnor U14147 (N_14147,N_13744,N_13845);
and U14148 (N_14148,N_13180,N_13124);
nor U14149 (N_14149,N_13611,N_13925);
and U14150 (N_14150,N_13779,N_13447);
nand U14151 (N_14151,N_13606,N_13620);
nor U14152 (N_14152,N_13513,N_13000);
nand U14153 (N_14153,N_13387,N_13667);
xor U14154 (N_14154,N_13498,N_13936);
xnor U14155 (N_14155,N_13725,N_13077);
nor U14156 (N_14156,N_13784,N_13880);
or U14157 (N_14157,N_13416,N_13312);
nor U14158 (N_14158,N_13837,N_13558);
and U14159 (N_14159,N_13617,N_13153);
or U14160 (N_14160,N_13417,N_13270);
xor U14161 (N_14161,N_13879,N_13660);
and U14162 (N_14162,N_13638,N_13715);
or U14163 (N_14163,N_13937,N_13570);
nor U14164 (N_14164,N_13610,N_13604);
and U14165 (N_14165,N_13855,N_13973);
and U14166 (N_14166,N_13665,N_13464);
nor U14167 (N_14167,N_13948,N_13911);
or U14168 (N_14168,N_13874,N_13313);
or U14169 (N_14169,N_13361,N_13559);
nor U14170 (N_14170,N_13362,N_13647);
and U14171 (N_14171,N_13683,N_13154);
nor U14172 (N_14172,N_13804,N_13814);
nand U14173 (N_14173,N_13947,N_13616);
xor U14174 (N_14174,N_13078,N_13754);
or U14175 (N_14175,N_13727,N_13359);
nand U14176 (N_14176,N_13173,N_13413);
and U14177 (N_14177,N_13145,N_13467);
or U14178 (N_14178,N_13242,N_13710);
nor U14179 (N_14179,N_13642,N_13908);
or U14180 (N_14180,N_13503,N_13421);
and U14181 (N_14181,N_13485,N_13782);
or U14182 (N_14182,N_13554,N_13005);
nor U14183 (N_14183,N_13663,N_13376);
nor U14184 (N_14184,N_13536,N_13600);
xnor U14185 (N_14185,N_13012,N_13693);
nand U14186 (N_14186,N_13332,N_13383);
xnor U14187 (N_14187,N_13214,N_13685);
or U14188 (N_14188,N_13907,N_13816);
and U14189 (N_14189,N_13994,N_13976);
nand U14190 (N_14190,N_13872,N_13260);
and U14191 (N_14191,N_13890,N_13679);
and U14192 (N_14192,N_13825,N_13469);
and U14193 (N_14193,N_13085,N_13448);
nor U14194 (N_14194,N_13499,N_13807);
and U14195 (N_14195,N_13392,N_13480);
and U14196 (N_14196,N_13918,N_13205);
and U14197 (N_14197,N_13520,N_13509);
xnor U14198 (N_14198,N_13863,N_13083);
and U14199 (N_14199,N_13516,N_13707);
xnor U14200 (N_14200,N_13300,N_13440);
or U14201 (N_14201,N_13778,N_13184);
and U14202 (N_14202,N_13132,N_13412);
or U14203 (N_14203,N_13080,N_13946);
or U14204 (N_14204,N_13527,N_13391);
nor U14205 (N_14205,N_13261,N_13315);
or U14206 (N_14206,N_13985,N_13755);
and U14207 (N_14207,N_13382,N_13325);
nor U14208 (N_14208,N_13488,N_13204);
nor U14209 (N_14209,N_13198,N_13731);
or U14210 (N_14210,N_13027,N_13365);
nor U14211 (N_14211,N_13608,N_13876);
xor U14212 (N_14212,N_13137,N_13473);
nor U14213 (N_14213,N_13052,N_13126);
and U14214 (N_14214,N_13717,N_13156);
nand U14215 (N_14215,N_13690,N_13535);
xor U14216 (N_14216,N_13108,N_13808);
or U14217 (N_14217,N_13096,N_13773);
xnor U14218 (N_14218,N_13269,N_13547);
or U14219 (N_14219,N_13974,N_13291);
xor U14220 (N_14220,N_13327,N_13017);
and U14221 (N_14221,N_13590,N_13569);
and U14222 (N_14222,N_13959,N_13818);
and U14223 (N_14223,N_13692,N_13100);
nand U14224 (N_14224,N_13560,N_13262);
nand U14225 (N_14225,N_13521,N_13118);
xor U14226 (N_14226,N_13578,N_13002);
and U14227 (N_14227,N_13316,N_13902);
xnor U14228 (N_14228,N_13666,N_13229);
nor U14229 (N_14229,N_13045,N_13924);
xnor U14230 (N_14230,N_13615,N_13030);
and U14231 (N_14231,N_13484,N_13433);
and U14232 (N_14232,N_13181,N_13817);
or U14233 (N_14233,N_13028,N_13673);
nand U14234 (N_14234,N_13709,N_13758);
nor U14235 (N_14235,N_13236,N_13061);
nor U14236 (N_14236,N_13722,N_13050);
nand U14237 (N_14237,N_13991,N_13955);
nor U14238 (N_14238,N_13801,N_13435);
xor U14239 (N_14239,N_13847,N_13896);
or U14240 (N_14240,N_13764,N_13649);
nand U14241 (N_14241,N_13839,N_13113);
xor U14242 (N_14242,N_13169,N_13010);
or U14243 (N_14243,N_13742,N_13519);
xor U14244 (N_14244,N_13555,N_13452);
or U14245 (N_14245,N_13706,N_13544);
or U14246 (N_14246,N_13223,N_13828);
nor U14247 (N_14247,N_13714,N_13753);
or U14248 (N_14248,N_13377,N_13583);
and U14249 (N_14249,N_13360,N_13092);
xor U14250 (N_14250,N_13001,N_13552);
nand U14251 (N_14251,N_13314,N_13143);
nand U14252 (N_14252,N_13967,N_13468);
and U14253 (N_14253,N_13033,N_13211);
and U14254 (N_14254,N_13687,N_13968);
nand U14255 (N_14255,N_13463,N_13194);
nand U14256 (N_14256,N_13549,N_13750);
xor U14257 (N_14257,N_13629,N_13636);
or U14258 (N_14258,N_13060,N_13160);
xor U14259 (N_14259,N_13957,N_13209);
nand U14260 (N_14260,N_13877,N_13813);
or U14261 (N_14261,N_13769,N_13905);
or U14262 (N_14262,N_13935,N_13196);
and U14263 (N_14263,N_13420,N_13333);
or U14264 (N_14264,N_13183,N_13644);
or U14265 (N_14265,N_13592,N_13912);
or U14266 (N_14266,N_13550,N_13228);
nand U14267 (N_14267,N_13475,N_13471);
nand U14268 (N_14268,N_13491,N_13356);
nand U14269 (N_14269,N_13944,N_13862);
nand U14270 (N_14270,N_13148,N_13939);
or U14271 (N_14271,N_13910,N_13572);
xnor U14272 (N_14272,N_13415,N_13414);
and U14273 (N_14273,N_13422,N_13568);
and U14274 (N_14274,N_13168,N_13239);
xnor U14275 (N_14275,N_13064,N_13800);
nand U14276 (N_14276,N_13128,N_13431);
and U14277 (N_14277,N_13022,N_13032);
or U14278 (N_14278,N_13882,N_13259);
nor U14279 (N_14279,N_13343,N_13289);
xor U14280 (N_14280,N_13095,N_13508);
or U14281 (N_14281,N_13767,N_13838);
nand U14282 (N_14282,N_13283,N_13645);
xor U14283 (N_14283,N_13675,N_13251);
xnor U14284 (N_14284,N_13371,N_13605);
xor U14285 (N_14285,N_13740,N_13597);
nand U14286 (N_14286,N_13465,N_13334);
or U14287 (N_14287,N_13786,N_13240);
or U14288 (N_14288,N_13235,N_13101);
xor U14289 (N_14289,N_13836,N_13190);
nor U14290 (N_14290,N_13257,N_13394);
nand U14291 (N_14291,N_13894,N_13803);
and U14292 (N_14292,N_13791,N_13049);
xnor U14293 (N_14293,N_13424,N_13213);
xnor U14294 (N_14294,N_13737,N_13795);
xnor U14295 (N_14295,N_13996,N_13306);
or U14296 (N_14296,N_13482,N_13917);
xnor U14297 (N_14297,N_13366,N_13871);
xor U14298 (N_14298,N_13353,N_13007);
xor U14299 (N_14299,N_13072,N_13598);
xnor U14300 (N_14300,N_13098,N_13195);
or U14301 (N_14301,N_13574,N_13167);
nor U14302 (N_14302,N_13265,N_13053);
nand U14303 (N_14303,N_13736,N_13020);
or U14304 (N_14304,N_13584,N_13141);
or U14305 (N_14305,N_13512,N_13810);
or U14306 (N_14306,N_13466,N_13898);
nor U14307 (N_14307,N_13831,N_13739);
xor U14308 (N_14308,N_13759,N_13093);
xnor U14309 (N_14309,N_13747,N_13134);
nand U14310 (N_14310,N_13057,N_13338);
or U14311 (N_14311,N_13713,N_13490);
nor U14312 (N_14312,N_13745,N_13720);
xnor U14313 (N_14313,N_13805,N_13063);
nand U14314 (N_14314,N_13117,N_13963);
xnor U14315 (N_14315,N_13848,N_13402);
nand U14316 (N_14316,N_13942,N_13191);
xor U14317 (N_14317,N_13749,N_13928);
xor U14318 (N_14318,N_13650,N_13164);
nand U14319 (N_14319,N_13852,N_13248);
nand U14320 (N_14320,N_13441,N_13969);
nand U14321 (N_14321,N_13729,N_13321);
or U14322 (N_14322,N_13171,N_13794);
and U14323 (N_14323,N_13614,N_13274);
xor U14324 (N_14324,N_13631,N_13618);
xnor U14325 (N_14325,N_13026,N_13657);
and U14326 (N_14326,N_13225,N_13329);
and U14327 (N_14327,N_13797,N_13406);
and U14328 (N_14328,N_13043,N_13297);
or U14329 (N_14329,N_13264,N_13582);
xnor U14330 (N_14330,N_13129,N_13860);
nand U14331 (N_14331,N_13437,N_13258);
nand U14332 (N_14332,N_13884,N_13317);
and U14333 (N_14333,N_13425,N_13951);
and U14334 (N_14334,N_13345,N_13885);
or U14335 (N_14335,N_13730,N_13843);
or U14336 (N_14336,N_13505,N_13840);
nor U14337 (N_14337,N_13986,N_13961);
and U14338 (N_14338,N_13502,N_13170);
or U14339 (N_14339,N_13252,N_13237);
nand U14340 (N_14340,N_13348,N_13531);
or U14341 (N_14341,N_13227,N_13233);
nor U14342 (N_14342,N_13953,N_13112);
and U14343 (N_14343,N_13013,N_13074);
nor U14344 (N_14344,N_13253,N_13775);
nor U14345 (N_14345,N_13432,N_13875);
or U14346 (N_14346,N_13640,N_13686);
and U14347 (N_14347,N_13157,N_13070);
and U14348 (N_14348,N_13990,N_13103);
xnor U14349 (N_14349,N_13146,N_13374);
xnor U14350 (N_14350,N_13702,N_13286);
and U14351 (N_14351,N_13089,N_13820);
and U14352 (N_14352,N_13024,N_13019);
nand U14353 (N_14353,N_13303,N_13790);
or U14354 (N_14354,N_13319,N_13330);
xor U14355 (N_14355,N_13962,N_13524);
and U14356 (N_14356,N_13528,N_13398);
nand U14357 (N_14357,N_13116,N_13887);
nand U14358 (N_14358,N_13972,N_13930);
nand U14359 (N_14359,N_13111,N_13287);
nand U14360 (N_14360,N_13188,N_13224);
and U14361 (N_14361,N_13210,N_13147);
nand U14362 (N_14362,N_13051,N_13461);
and U14363 (N_14363,N_13851,N_13084);
or U14364 (N_14364,N_13561,N_13277);
or U14365 (N_14365,N_13751,N_13159);
and U14366 (N_14366,N_13798,N_13612);
nor U14367 (N_14367,N_13302,N_13829);
xnor U14368 (N_14368,N_13609,N_13161);
or U14369 (N_14369,N_13444,N_13762);
xor U14370 (N_14370,N_13130,N_13368);
or U14371 (N_14371,N_13622,N_13451);
nand U14372 (N_14372,N_13929,N_13185);
xor U14373 (N_14373,N_13656,N_13842);
and U14374 (N_14374,N_13643,N_13811);
nand U14375 (N_14375,N_13483,N_13589);
or U14376 (N_14376,N_13335,N_13501);
and U14377 (N_14377,N_13651,N_13585);
and U14378 (N_14378,N_13487,N_13859);
or U14379 (N_14379,N_13682,N_13273);
nand U14380 (N_14380,N_13109,N_13975);
xor U14381 (N_14381,N_13591,N_13367);
xnor U14382 (N_14382,N_13774,N_13427);
xor U14383 (N_14383,N_13866,N_13380);
xnor U14384 (N_14384,N_13945,N_13243);
and U14385 (N_14385,N_13659,N_13208);
or U14386 (N_14386,N_13384,N_13517);
nand U14387 (N_14387,N_13014,N_13405);
nor U14388 (N_14388,N_13496,N_13272);
xor U14389 (N_14389,N_13777,N_13370);
xor U14390 (N_14390,N_13648,N_13102);
or U14391 (N_14391,N_13646,N_13222);
nand U14392 (N_14392,N_13279,N_13256);
or U14393 (N_14393,N_13680,N_13699);
or U14394 (N_14394,N_13748,N_13340);
nand U14395 (N_14395,N_13493,N_13041);
nor U14396 (N_14396,N_13653,N_13217);
xnor U14397 (N_14397,N_13661,N_13136);
nor U14398 (N_14398,N_13388,N_13909);
and U14399 (N_14399,N_13971,N_13886);
xnor U14400 (N_14400,N_13563,N_13678);
nand U14401 (N_14401,N_13186,N_13856);
xnor U14402 (N_14402,N_13899,N_13694);
and U14403 (N_14403,N_13023,N_13282);
nor U14404 (N_14404,N_13672,N_13477);
and U14405 (N_14405,N_13221,N_13901);
nor U14406 (N_14406,N_13846,N_13373);
xnor U14407 (N_14407,N_13250,N_13029);
and U14408 (N_14408,N_13670,N_13538);
and U14409 (N_14409,N_13922,N_13630);
or U14410 (N_14410,N_13470,N_13131);
and U14411 (N_14411,N_13411,N_13696);
nor U14412 (N_14412,N_13580,N_13977);
or U14413 (N_14413,N_13579,N_13732);
xnor U14414 (N_14414,N_13586,N_13206);
nand U14415 (N_14415,N_13215,N_13292);
or U14416 (N_14416,N_13537,N_13788);
and U14417 (N_14417,N_13339,N_13548);
or U14418 (N_14418,N_13835,N_13708);
nand U14419 (N_14419,N_13246,N_13149);
and U14420 (N_14420,N_13662,N_13726);
and U14421 (N_14421,N_13787,N_13025);
nor U14422 (N_14422,N_13086,N_13966);
or U14423 (N_14423,N_13867,N_13218);
nor U14424 (N_14424,N_13819,N_13881);
xor U14425 (N_14425,N_13595,N_13841);
nor U14426 (N_14426,N_13322,N_13781);
nor U14427 (N_14427,N_13792,N_13893);
or U14428 (N_14428,N_13821,N_13613);
and U14429 (N_14429,N_13763,N_13979);
nor U14430 (N_14430,N_13895,N_13054);
xnor U14431 (N_14431,N_13919,N_13562);
xor U14432 (N_14432,N_13047,N_13280);
nand U14433 (N_14433,N_13187,N_13075);
nand U14434 (N_14434,N_13336,N_13450);
and U14435 (N_14435,N_13903,N_13021);
nor U14436 (N_14436,N_13234,N_13015);
or U14437 (N_14437,N_13724,N_13897);
or U14438 (N_14438,N_13853,N_13310);
and U14439 (N_14439,N_13619,N_13065);
or U14440 (N_14440,N_13443,N_13756);
and U14441 (N_14441,N_13457,N_13369);
nor U14442 (N_14442,N_13577,N_13522);
nor U14443 (N_14443,N_13564,N_13281);
nor U14444 (N_14444,N_13454,N_13557);
nand U14445 (N_14445,N_13495,N_13073);
nand U14446 (N_14446,N_13399,N_13438);
xor U14447 (N_14447,N_13705,N_13163);
or U14448 (N_14448,N_13960,N_13474);
or U14449 (N_14449,N_13263,N_13326);
nor U14450 (N_14450,N_13639,N_13094);
or U14451 (N_14451,N_13133,N_13040);
nor U14452 (N_14452,N_13833,N_13984);
xnor U14453 (N_14453,N_13226,N_13081);
xnor U14454 (N_14454,N_13122,N_13445);
or U14455 (N_14455,N_13182,N_13865);
and U14456 (N_14456,N_13193,N_13201);
or U14457 (N_14457,N_13566,N_13658);
nand U14458 (N_14458,N_13988,N_13492);
xnor U14459 (N_14459,N_13891,N_13059);
and U14460 (N_14460,N_13980,N_13674);
nor U14461 (N_14461,N_13943,N_13110);
xnor U14462 (N_14462,N_13652,N_13298);
xor U14463 (N_14463,N_13983,N_13087);
or U14464 (N_14464,N_13462,N_13506);
xnor U14465 (N_14465,N_13776,N_13106);
or U14466 (N_14466,N_13932,N_13904);
xnor U14467 (N_14467,N_13288,N_13400);
and U14468 (N_14468,N_13723,N_13123);
and U14469 (N_14469,N_13172,N_13823);
and U14470 (N_14470,N_13870,N_13995);
xor U14471 (N_14471,N_13627,N_13571);
and U14472 (N_14472,N_13626,N_13082);
or U14473 (N_14473,N_13355,N_13768);
or U14474 (N_14474,N_13044,N_13238);
nor U14475 (N_14475,N_13868,N_13892);
and U14476 (N_14476,N_13701,N_13689);
or U14477 (N_14477,N_13676,N_13212);
nand U14478 (N_14478,N_13542,N_13906);
nand U14479 (N_14479,N_13681,N_13765);
nand U14480 (N_14480,N_13175,N_13734);
nand U14481 (N_14481,N_13207,N_13449);
xor U14482 (N_14482,N_13318,N_13721);
nand U14483 (N_14483,N_13009,N_13178);
or U14484 (N_14484,N_13478,N_13700);
or U14485 (N_14485,N_13037,N_13177);
xor U14486 (N_14486,N_13453,N_13342);
or U14487 (N_14487,N_13105,N_13042);
nand U14488 (N_14488,N_13176,N_13244);
nand U14489 (N_14489,N_13016,N_13553);
nor U14490 (N_14490,N_13337,N_13864);
nand U14491 (N_14491,N_13456,N_13344);
nand U14492 (N_14492,N_13796,N_13711);
nand U14493 (N_14493,N_13090,N_13247);
xor U14494 (N_14494,N_13216,N_13900);
nand U14495 (N_14495,N_13179,N_13039);
nor U14496 (N_14496,N_13940,N_13460);
and U14497 (N_14497,N_13308,N_13789);
nand U14498 (N_14498,N_13873,N_13854);
nand U14499 (N_14499,N_13704,N_13931);
or U14500 (N_14500,N_13068,N_13212);
or U14501 (N_14501,N_13814,N_13857);
and U14502 (N_14502,N_13617,N_13896);
nand U14503 (N_14503,N_13233,N_13724);
nor U14504 (N_14504,N_13250,N_13978);
and U14505 (N_14505,N_13670,N_13643);
xnor U14506 (N_14506,N_13447,N_13351);
or U14507 (N_14507,N_13483,N_13968);
or U14508 (N_14508,N_13389,N_13363);
and U14509 (N_14509,N_13482,N_13847);
nor U14510 (N_14510,N_13585,N_13070);
and U14511 (N_14511,N_13567,N_13950);
nor U14512 (N_14512,N_13630,N_13182);
or U14513 (N_14513,N_13335,N_13857);
and U14514 (N_14514,N_13319,N_13471);
nand U14515 (N_14515,N_13844,N_13633);
and U14516 (N_14516,N_13360,N_13452);
nor U14517 (N_14517,N_13650,N_13970);
nor U14518 (N_14518,N_13786,N_13322);
nand U14519 (N_14519,N_13016,N_13414);
and U14520 (N_14520,N_13501,N_13437);
or U14521 (N_14521,N_13953,N_13256);
and U14522 (N_14522,N_13978,N_13800);
or U14523 (N_14523,N_13480,N_13661);
and U14524 (N_14524,N_13890,N_13925);
nor U14525 (N_14525,N_13452,N_13033);
or U14526 (N_14526,N_13044,N_13906);
or U14527 (N_14527,N_13356,N_13823);
and U14528 (N_14528,N_13429,N_13699);
nor U14529 (N_14529,N_13555,N_13117);
or U14530 (N_14530,N_13847,N_13702);
nor U14531 (N_14531,N_13311,N_13155);
and U14532 (N_14532,N_13831,N_13706);
or U14533 (N_14533,N_13004,N_13328);
nor U14534 (N_14534,N_13711,N_13942);
nor U14535 (N_14535,N_13449,N_13080);
nor U14536 (N_14536,N_13240,N_13646);
nand U14537 (N_14537,N_13203,N_13153);
and U14538 (N_14538,N_13662,N_13858);
nor U14539 (N_14539,N_13874,N_13199);
nor U14540 (N_14540,N_13666,N_13378);
nand U14541 (N_14541,N_13896,N_13695);
and U14542 (N_14542,N_13539,N_13833);
nand U14543 (N_14543,N_13227,N_13129);
nor U14544 (N_14544,N_13637,N_13640);
nand U14545 (N_14545,N_13769,N_13672);
and U14546 (N_14546,N_13086,N_13349);
nor U14547 (N_14547,N_13344,N_13320);
xor U14548 (N_14548,N_13621,N_13571);
and U14549 (N_14549,N_13486,N_13607);
and U14550 (N_14550,N_13514,N_13610);
xor U14551 (N_14551,N_13979,N_13203);
nor U14552 (N_14552,N_13455,N_13085);
or U14553 (N_14553,N_13927,N_13515);
and U14554 (N_14554,N_13946,N_13141);
xnor U14555 (N_14555,N_13958,N_13031);
nand U14556 (N_14556,N_13084,N_13378);
xnor U14557 (N_14557,N_13562,N_13028);
or U14558 (N_14558,N_13705,N_13317);
xnor U14559 (N_14559,N_13613,N_13915);
nand U14560 (N_14560,N_13511,N_13521);
nand U14561 (N_14561,N_13289,N_13627);
xnor U14562 (N_14562,N_13982,N_13774);
xnor U14563 (N_14563,N_13374,N_13616);
or U14564 (N_14564,N_13079,N_13565);
nor U14565 (N_14565,N_13355,N_13076);
nand U14566 (N_14566,N_13318,N_13439);
or U14567 (N_14567,N_13011,N_13024);
nand U14568 (N_14568,N_13525,N_13816);
and U14569 (N_14569,N_13202,N_13465);
or U14570 (N_14570,N_13776,N_13061);
xor U14571 (N_14571,N_13526,N_13814);
or U14572 (N_14572,N_13689,N_13706);
xnor U14573 (N_14573,N_13390,N_13677);
or U14574 (N_14574,N_13073,N_13898);
xor U14575 (N_14575,N_13382,N_13807);
xnor U14576 (N_14576,N_13253,N_13991);
or U14577 (N_14577,N_13365,N_13505);
xor U14578 (N_14578,N_13634,N_13426);
and U14579 (N_14579,N_13018,N_13982);
and U14580 (N_14580,N_13565,N_13335);
nor U14581 (N_14581,N_13196,N_13084);
xor U14582 (N_14582,N_13953,N_13117);
nor U14583 (N_14583,N_13038,N_13090);
and U14584 (N_14584,N_13973,N_13515);
nor U14585 (N_14585,N_13944,N_13765);
nor U14586 (N_14586,N_13786,N_13460);
or U14587 (N_14587,N_13331,N_13277);
nor U14588 (N_14588,N_13908,N_13997);
and U14589 (N_14589,N_13405,N_13643);
xor U14590 (N_14590,N_13252,N_13522);
xor U14591 (N_14591,N_13165,N_13491);
nand U14592 (N_14592,N_13998,N_13557);
nor U14593 (N_14593,N_13663,N_13847);
or U14594 (N_14594,N_13418,N_13488);
or U14595 (N_14595,N_13150,N_13083);
or U14596 (N_14596,N_13576,N_13957);
and U14597 (N_14597,N_13883,N_13807);
xor U14598 (N_14598,N_13068,N_13640);
nor U14599 (N_14599,N_13668,N_13021);
and U14600 (N_14600,N_13700,N_13416);
nand U14601 (N_14601,N_13236,N_13904);
or U14602 (N_14602,N_13141,N_13504);
nand U14603 (N_14603,N_13940,N_13897);
xnor U14604 (N_14604,N_13740,N_13088);
and U14605 (N_14605,N_13878,N_13788);
and U14606 (N_14606,N_13771,N_13790);
and U14607 (N_14607,N_13428,N_13040);
and U14608 (N_14608,N_13336,N_13638);
nand U14609 (N_14609,N_13283,N_13694);
nand U14610 (N_14610,N_13066,N_13740);
nand U14611 (N_14611,N_13203,N_13107);
or U14612 (N_14612,N_13549,N_13763);
xnor U14613 (N_14613,N_13421,N_13661);
xnor U14614 (N_14614,N_13198,N_13720);
xnor U14615 (N_14615,N_13183,N_13504);
xnor U14616 (N_14616,N_13330,N_13720);
or U14617 (N_14617,N_13468,N_13743);
xor U14618 (N_14618,N_13410,N_13621);
xor U14619 (N_14619,N_13755,N_13536);
or U14620 (N_14620,N_13553,N_13848);
or U14621 (N_14621,N_13397,N_13818);
nand U14622 (N_14622,N_13318,N_13981);
nand U14623 (N_14623,N_13545,N_13377);
and U14624 (N_14624,N_13827,N_13766);
and U14625 (N_14625,N_13528,N_13482);
or U14626 (N_14626,N_13675,N_13242);
xnor U14627 (N_14627,N_13139,N_13730);
nand U14628 (N_14628,N_13750,N_13552);
or U14629 (N_14629,N_13700,N_13892);
or U14630 (N_14630,N_13866,N_13401);
xnor U14631 (N_14631,N_13364,N_13606);
nand U14632 (N_14632,N_13714,N_13542);
and U14633 (N_14633,N_13441,N_13676);
xor U14634 (N_14634,N_13828,N_13485);
nand U14635 (N_14635,N_13435,N_13060);
nand U14636 (N_14636,N_13882,N_13123);
and U14637 (N_14637,N_13754,N_13504);
or U14638 (N_14638,N_13939,N_13444);
and U14639 (N_14639,N_13539,N_13851);
xnor U14640 (N_14640,N_13653,N_13605);
nand U14641 (N_14641,N_13990,N_13603);
and U14642 (N_14642,N_13715,N_13490);
xnor U14643 (N_14643,N_13569,N_13427);
xnor U14644 (N_14644,N_13847,N_13350);
nor U14645 (N_14645,N_13042,N_13730);
and U14646 (N_14646,N_13003,N_13347);
and U14647 (N_14647,N_13857,N_13513);
xor U14648 (N_14648,N_13039,N_13361);
nor U14649 (N_14649,N_13437,N_13296);
or U14650 (N_14650,N_13463,N_13174);
and U14651 (N_14651,N_13651,N_13966);
nand U14652 (N_14652,N_13323,N_13739);
xor U14653 (N_14653,N_13959,N_13669);
nand U14654 (N_14654,N_13221,N_13751);
or U14655 (N_14655,N_13230,N_13472);
nor U14656 (N_14656,N_13880,N_13587);
or U14657 (N_14657,N_13627,N_13158);
xnor U14658 (N_14658,N_13987,N_13620);
nand U14659 (N_14659,N_13499,N_13909);
xnor U14660 (N_14660,N_13818,N_13322);
or U14661 (N_14661,N_13349,N_13236);
nand U14662 (N_14662,N_13760,N_13551);
and U14663 (N_14663,N_13130,N_13259);
xor U14664 (N_14664,N_13934,N_13118);
nand U14665 (N_14665,N_13176,N_13481);
or U14666 (N_14666,N_13683,N_13369);
nor U14667 (N_14667,N_13327,N_13101);
nand U14668 (N_14668,N_13752,N_13826);
or U14669 (N_14669,N_13843,N_13246);
nor U14670 (N_14670,N_13775,N_13449);
and U14671 (N_14671,N_13505,N_13265);
nor U14672 (N_14672,N_13296,N_13624);
or U14673 (N_14673,N_13192,N_13874);
xor U14674 (N_14674,N_13882,N_13336);
nor U14675 (N_14675,N_13640,N_13551);
nand U14676 (N_14676,N_13954,N_13932);
nor U14677 (N_14677,N_13055,N_13572);
nor U14678 (N_14678,N_13198,N_13341);
nand U14679 (N_14679,N_13973,N_13045);
and U14680 (N_14680,N_13063,N_13610);
and U14681 (N_14681,N_13841,N_13604);
xor U14682 (N_14682,N_13848,N_13118);
xor U14683 (N_14683,N_13972,N_13550);
or U14684 (N_14684,N_13294,N_13778);
or U14685 (N_14685,N_13467,N_13311);
nand U14686 (N_14686,N_13445,N_13036);
nand U14687 (N_14687,N_13283,N_13113);
and U14688 (N_14688,N_13900,N_13162);
and U14689 (N_14689,N_13992,N_13758);
nand U14690 (N_14690,N_13079,N_13246);
and U14691 (N_14691,N_13118,N_13020);
and U14692 (N_14692,N_13988,N_13010);
or U14693 (N_14693,N_13308,N_13084);
xnor U14694 (N_14694,N_13666,N_13642);
nand U14695 (N_14695,N_13080,N_13914);
xor U14696 (N_14696,N_13636,N_13726);
or U14697 (N_14697,N_13668,N_13284);
nor U14698 (N_14698,N_13067,N_13603);
nor U14699 (N_14699,N_13547,N_13579);
or U14700 (N_14700,N_13896,N_13144);
xnor U14701 (N_14701,N_13042,N_13660);
and U14702 (N_14702,N_13377,N_13629);
nand U14703 (N_14703,N_13277,N_13465);
or U14704 (N_14704,N_13262,N_13397);
or U14705 (N_14705,N_13578,N_13594);
or U14706 (N_14706,N_13856,N_13349);
nand U14707 (N_14707,N_13451,N_13656);
nand U14708 (N_14708,N_13831,N_13312);
or U14709 (N_14709,N_13044,N_13918);
xnor U14710 (N_14710,N_13732,N_13199);
and U14711 (N_14711,N_13824,N_13335);
nor U14712 (N_14712,N_13381,N_13440);
nor U14713 (N_14713,N_13745,N_13370);
nor U14714 (N_14714,N_13659,N_13498);
xor U14715 (N_14715,N_13178,N_13583);
nand U14716 (N_14716,N_13403,N_13355);
xor U14717 (N_14717,N_13203,N_13434);
nand U14718 (N_14718,N_13678,N_13370);
nor U14719 (N_14719,N_13910,N_13974);
xor U14720 (N_14720,N_13727,N_13657);
nor U14721 (N_14721,N_13295,N_13695);
and U14722 (N_14722,N_13582,N_13686);
nand U14723 (N_14723,N_13887,N_13149);
xnor U14724 (N_14724,N_13398,N_13854);
nand U14725 (N_14725,N_13620,N_13406);
xnor U14726 (N_14726,N_13109,N_13898);
and U14727 (N_14727,N_13136,N_13168);
nand U14728 (N_14728,N_13392,N_13768);
nand U14729 (N_14729,N_13155,N_13116);
nor U14730 (N_14730,N_13309,N_13759);
nor U14731 (N_14731,N_13475,N_13592);
xnor U14732 (N_14732,N_13369,N_13633);
or U14733 (N_14733,N_13236,N_13277);
xor U14734 (N_14734,N_13661,N_13900);
xnor U14735 (N_14735,N_13964,N_13737);
xor U14736 (N_14736,N_13153,N_13596);
nor U14737 (N_14737,N_13666,N_13905);
nor U14738 (N_14738,N_13390,N_13419);
xnor U14739 (N_14739,N_13576,N_13022);
or U14740 (N_14740,N_13136,N_13560);
or U14741 (N_14741,N_13859,N_13209);
xor U14742 (N_14742,N_13497,N_13367);
or U14743 (N_14743,N_13203,N_13943);
nand U14744 (N_14744,N_13412,N_13566);
nor U14745 (N_14745,N_13847,N_13559);
nand U14746 (N_14746,N_13554,N_13780);
xnor U14747 (N_14747,N_13118,N_13067);
and U14748 (N_14748,N_13864,N_13717);
xnor U14749 (N_14749,N_13915,N_13900);
and U14750 (N_14750,N_13065,N_13908);
and U14751 (N_14751,N_13090,N_13867);
nand U14752 (N_14752,N_13084,N_13183);
xor U14753 (N_14753,N_13807,N_13264);
or U14754 (N_14754,N_13739,N_13883);
nand U14755 (N_14755,N_13120,N_13302);
and U14756 (N_14756,N_13397,N_13335);
nand U14757 (N_14757,N_13822,N_13261);
or U14758 (N_14758,N_13482,N_13427);
xnor U14759 (N_14759,N_13701,N_13288);
and U14760 (N_14760,N_13188,N_13541);
and U14761 (N_14761,N_13755,N_13959);
nor U14762 (N_14762,N_13908,N_13576);
and U14763 (N_14763,N_13855,N_13836);
nor U14764 (N_14764,N_13540,N_13251);
xor U14765 (N_14765,N_13359,N_13350);
nor U14766 (N_14766,N_13120,N_13253);
nor U14767 (N_14767,N_13130,N_13333);
or U14768 (N_14768,N_13207,N_13923);
nand U14769 (N_14769,N_13407,N_13334);
nand U14770 (N_14770,N_13259,N_13712);
xnor U14771 (N_14771,N_13972,N_13075);
nand U14772 (N_14772,N_13892,N_13170);
or U14773 (N_14773,N_13789,N_13497);
nand U14774 (N_14774,N_13886,N_13070);
xnor U14775 (N_14775,N_13424,N_13259);
xnor U14776 (N_14776,N_13196,N_13702);
xnor U14777 (N_14777,N_13964,N_13179);
xnor U14778 (N_14778,N_13700,N_13209);
nand U14779 (N_14779,N_13297,N_13402);
xor U14780 (N_14780,N_13512,N_13505);
nand U14781 (N_14781,N_13011,N_13591);
nor U14782 (N_14782,N_13171,N_13565);
nand U14783 (N_14783,N_13552,N_13077);
nor U14784 (N_14784,N_13359,N_13141);
and U14785 (N_14785,N_13255,N_13912);
xor U14786 (N_14786,N_13898,N_13908);
or U14787 (N_14787,N_13038,N_13256);
xnor U14788 (N_14788,N_13097,N_13978);
xnor U14789 (N_14789,N_13484,N_13771);
and U14790 (N_14790,N_13886,N_13154);
xor U14791 (N_14791,N_13295,N_13613);
xor U14792 (N_14792,N_13636,N_13133);
xnor U14793 (N_14793,N_13085,N_13364);
or U14794 (N_14794,N_13269,N_13668);
and U14795 (N_14795,N_13128,N_13992);
and U14796 (N_14796,N_13959,N_13518);
and U14797 (N_14797,N_13462,N_13980);
nor U14798 (N_14798,N_13008,N_13993);
and U14799 (N_14799,N_13470,N_13862);
and U14800 (N_14800,N_13559,N_13669);
nor U14801 (N_14801,N_13645,N_13184);
nor U14802 (N_14802,N_13722,N_13460);
or U14803 (N_14803,N_13519,N_13365);
and U14804 (N_14804,N_13435,N_13638);
or U14805 (N_14805,N_13725,N_13394);
nor U14806 (N_14806,N_13424,N_13157);
and U14807 (N_14807,N_13800,N_13377);
and U14808 (N_14808,N_13990,N_13096);
or U14809 (N_14809,N_13561,N_13307);
and U14810 (N_14810,N_13462,N_13369);
nand U14811 (N_14811,N_13655,N_13598);
and U14812 (N_14812,N_13040,N_13897);
nor U14813 (N_14813,N_13699,N_13450);
nand U14814 (N_14814,N_13660,N_13428);
nand U14815 (N_14815,N_13342,N_13798);
nand U14816 (N_14816,N_13440,N_13083);
and U14817 (N_14817,N_13298,N_13691);
nor U14818 (N_14818,N_13345,N_13323);
xor U14819 (N_14819,N_13569,N_13731);
and U14820 (N_14820,N_13287,N_13654);
or U14821 (N_14821,N_13552,N_13215);
nand U14822 (N_14822,N_13233,N_13108);
and U14823 (N_14823,N_13930,N_13291);
or U14824 (N_14824,N_13614,N_13782);
nor U14825 (N_14825,N_13789,N_13066);
nand U14826 (N_14826,N_13311,N_13099);
and U14827 (N_14827,N_13295,N_13209);
and U14828 (N_14828,N_13198,N_13296);
nor U14829 (N_14829,N_13617,N_13788);
nand U14830 (N_14830,N_13839,N_13127);
nor U14831 (N_14831,N_13256,N_13268);
and U14832 (N_14832,N_13553,N_13559);
and U14833 (N_14833,N_13384,N_13837);
nand U14834 (N_14834,N_13600,N_13608);
or U14835 (N_14835,N_13971,N_13919);
xor U14836 (N_14836,N_13774,N_13880);
and U14837 (N_14837,N_13823,N_13465);
or U14838 (N_14838,N_13263,N_13367);
xnor U14839 (N_14839,N_13732,N_13656);
nand U14840 (N_14840,N_13663,N_13129);
nand U14841 (N_14841,N_13774,N_13370);
xor U14842 (N_14842,N_13605,N_13910);
nand U14843 (N_14843,N_13045,N_13141);
nand U14844 (N_14844,N_13457,N_13566);
or U14845 (N_14845,N_13084,N_13123);
nand U14846 (N_14846,N_13093,N_13105);
and U14847 (N_14847,N_13692,N_13035);
xor U14848 (N_14848,N_13203,N_13794);
xnor U14849 (N_14849,N_13678,N_13986);
xor U14850 (N_14850,N_13061,N_13071);
xor U14851 (N_14851,N_13894,N_13463);
xor U14852 (N_14852,N_13212,N_13335);
xor U14853 (N_14853,N_13214,N_13182);
and U14854 (N_14854,N_13903,N_13561);
nand U14855 (N_14855,N_13018,N_13279);
nand U14856 (N_14856,N_13486,N_13656);
xor U14857 (N_14857,N_13458,N_13760);
nand U14858 (N_14858,N_13905,N_13913);
and U14859 (N_14859,N_13103,N_13446);
or U14860 (N_14860,N_13732,N_13294);
xor U14861 (N_14861,N_13918,N_13916);
nand U14862 (N_14862,N_13404,N_13984);
and U14863 (N_14863,N_13034,N_13028);
or U14864 (N_14864,N_13719,N_13318);
and U14865 (N_14865,N_13379,N_13266);
nor U14866 (N_14866,N_13681,N_13884);
nor U14867 (N_14867,N_13401,N_13596);
nand U14868 (N_14868,N_13550,N_13284);
nand U14869 (N_14869,N_13795,N_13896);
and U14870 (N_14870,N_13751,N_13599);
and U14871 (N_14871,N_13011,N_13188);
nor U14872 (N_14872,N_13280,N_13764);
xnor U14873 (N_14873,N_13425,N_13064);
xor U14874 (N_14874,N_13522,N_13260);
xor U14875 (N_14875,N_13534,N_13568);
xor U14876 (N_14876,N_13725,N_13162);
nand U14877 (N_14877,N_13330,N_13814);
xnor U14878 (N_14878,N_13739,N_13542);
and U14879 (N_14879,N_13341,N_13071);
xor U14880 (N_14880,N_13208,N_13949);
nand U14881 (N_14881,N_13716,N_13929);
or U14882 (N_14882,N_13650,N_13353);
and U14883 (N_14883,N_13377,N_13353);
nand U14884 (N_14884,N_13678,N_13727);
nor U14885 (N_14885,N_13325,N_13047);
and U14886 (N_14886,N_13744,N_13635);
or U14887 (N_14887,N_13398,N_13383);
nor U14888 (N_14888,N_13725,N_13384);
or U14889 (N_14889,N_13491,N_13933);
nor U14890 (N_14890,N_13334,N_13021);
nor U14891 (N_14891,N_13435,N_13916);
or U14892 (N_14892,N_13513,N_13525);
or U14893 (N_14893,N_13787,N_13823);
nand U14894 (N_14894,N_13075,N_13665);
or U14895 (N_14895,N_13853,N_13057);
xnor U14896 (N_14896,N_13452,N_13927);
and U14897 (N_14897,N_13884,N_13889);
nor U14898 (N_14898,N_13225,N_13681);
nor U14899 (N_14899,N_13960,N_13090);
nor U14900 (N_14900,N_13111,N_13544);
nand U14901 (N_14901,N_13804,N_13198);
nand U14902 (N_14902,N_13092,N_13884);
or U14903 (N_14903,N_13814,N_13139);
nor U14904 (N_14904,N_13554,N_13111);
xnor U14905 (N_14905,N_13545,N_13821);
and U14906 (N_14906,N_13449,N_13521);
nor U14907 (N_14907,N_13397,N_13522);
and U14908 (N_14908,N_13418,N_13682);
or U14909 (N_14909,N_13568,N_13019);
or U14910 (N_14910,N_13999,N_13703);
xnor U14911 (N_14911,N_13192,N_13188);
and U14912 (N_14912,N_13148,N_13073);
xnor U14913 (N_14913,N_13540,N_13760);
nand U14914 (N_14914,N_13196,N_13824);
and U14915 (N_14915,N_13256,N_13168);
and U14916 (N_14916,N_13078,N_13618);
or U14917 (N_14917,N_13236,N_13097);
nor U14918 (N_14918,N_13622,N_13531);
xnor U14919 (N_14919,N_13290,N_13517);
or U14920 (N_14920,N_13580,N_13125);
nor U14921 (N_14921,N_13472,N_13340);
nand U14922 (N_14922,N_13560,N_13880);
xnor U14923 (N_14923,N_13864,N_13939);
nor U14924 (N_14924,N_13433,N_13768);
and U14925 (N_14925,N_13781,N_13180);
nand U14926 (N_14926,N_13702,N_13348);
nor U14927 (N_14927,N_13514,N_13869);
and U14928 (N_14928,N_13061,N_13769);
and U14929 (N_14929,N_13294,N_13156);
and U14930 (N_14930,N_13059,N_13405);
and U14931 (N_14931,N_13261,N_13053);
nand U14932 (N_14932,N_13834,N_13888);
or U14933 (N_14933,N_13211,N_13397);
and U14934 (N_14934,N_13458,N_13620);
xor U14935 (N_14935,N_13243,N_13545);
and U14936 (N_14936,N_13300,N_13095);
nand U14937 (N_14937,N_13047,N_13875);
and U14938 (N_14938,N_13161,N_13349);
nor U14939 (N_14939,N_13028,N_13335);
nor U14940 (N_14940,N_13543,N_13414);
or U14941 (N_14941,N_13251,N_13401);
or U14942 (N_14942,N_13059,N_13193);
nor U14943 (N_14943,N_13454,N_13135);
xnor U14944 (N_14944,N_13505,N_13201);
or U14945 (N_14945,N_13047,N_13485);
nor U14946 (N_14946,N_13277,N_13944);
xnor U14947 (N_14947,N_13968,N_13432);
or U14948 (N_14948,N_13174,N_13705);
nor U14949 (N_14949,N_13200,N_13865);
xnor U14950 (N_14950,N_13231,N_13446);
xor U14951 (N_14951,N_13218,N_13370);
nand U14952 (N_14952,N_13845,N_13746);
or U14953 (N_14953,N_13945,N_13038);
or U14954 (N_14954,N_13459,N_13472);
nor U14955 (N_14955,N_13083,N_13649);
nor U14956 (N_14956,N_13468,N_13174);
nand U14957 (N_14957,N_13197,N_13746);
nor U14958 (N_14958,N_13999,N_13750);
xor U14959 (N_14959,N_13591,N_13532);
or U14960 (N_14960,N_13917,N_13543);
nand U14961 (N_14961,N_13030,N_13883);
nand U14962 (N_14962,N_13729,N_13727);
and U14963 (N_14963,N_13364,N_13218);
xnor U14964 (N_14964,N_13521,N_13235);
xor U14965 (N_14965,N_13811,N_13579);
and U14966 (N_14966,N_13773,N_13278);
and U14967 (N_14967,N_13011,N_13175);
and U14968 (N_14968,N_13812,N_13047);
nand U14969 (N_14969,N_13478,N_13682);
nand U14970 (N_14970,N_13820,N_13487);
nand U14971 (N_14971,N_13116,N_13256);
and U14972 (N_14972,N_13145,N_13867);
nand U14973 (N_14973,N_13595,N_13910);
nand U14974 (N_14974,N_13319,N_13324);
or U14975 (N_14975,N_13924,N_13511);
and U14976 (N_14976,N_13124,N_13788);
and U14977 (N_14977,N_13408,N_13882);
xnor U14978 (N_14978,N_13433,N_13717);
and U14979 (N_14979,N_13587,N_13812);
xor U14980 (N_14980,N_13523,N_13600);
or U14981 (N_14981,N_13498,N_13838);
xor U14982 (N_14982,N_13499,N_13995);
nor U14983 (N_14983,N_13411,N_13885);
nor U14984 (N_14984,N_13854,N_13569);
xnor U14985 (N_14985,N_13178,N_13333);
or U14986 (N_14986,N_13953,N_13137);
and U14987 (N_14987,N_13054,N_13044);
or U14988 (N_14988,N_13709,N_13015);
xnor U14989 (N_14989,N_13006,N_13155);
and U14990 (N_14990,N_13512,N_13117);
and U14991 (N_14991,N_13501,N_13114);
and U14992 (N_14992,N_13073,N_13375);
nand U14993 (N_14993,N_13826,N_13330);
and U14994 (N_14994,N_13386,N_13443);
and U14995 (N_14995,N_13149,N_13761);
nand U14996 (N_14996,N_13212,N_13686);
or U14997 (N_14997,N_13818,N_13891);
nor U14998 (N_14998,N_13400,N_13860);
and U14999 (N_14999,N_13071,N_13818);
xnor UO_0 (O_0,N_14846,N_14528);
xor UO_1 (O_1,N_14086,N_14869);
and UO_2 (O_2,N_14531,N_14926);
xor UO_3 (O_3,N_14737,N_14983);
xnor UO_4 (O_4,N_14703,N_14497);
nor UO_5 (O_5,N_14235,N_14988);
or UO_6 (O_6,N_14655,N_14590);
and UO_7 (O_7,N_14997,N_14393);
or UO_8 (O_8,N_14185,N_14576);
nand UO_9 (O_9,N_14149,N_14602);
and UO_10 (O_10,N_14904,N_14546);
xor UO_11 (O_11,N_14338,N_14770);
or UO_12 (O_12,N_14544,N_14504);
and UO_13 (O_13,N_14698,N_14911);
nor UO_14 (O_14,N_14314,N_14785);
xnor UO_15 (O_15,N_14155,N_14377);
xor UO_16 (O_16,N_14794,N_14351);
xnor UO_17 (O_17,N_14199,N_14230);
and UO_18 (O_18,N_14740,N_14680);
or UO_19 (O_19,N_14500,N_14148);
xor UO_20 (O_20,N_14534,N_14387);
and UO_21 (O_21,N_14746,N_14508);
and UO_22 (O_22,N_14491,N_14592);
or UO_23 (O_23,N_14913,N_14456);
or UO_24 (O_24,N_14815,N_14370);
nand UO_25 (O_25,N_14315,N_14311);
nor UO_26 (O_26,N_14626,N_14608);
nand UO_27 (O_27,N_14567,N_14245);
xor UO_28 (O_28,N_14645,N_14901);
or UO_29 (O_29,N_14925,N_14405);
or UO_30 (O_30,N_14635,N_14458);
nand UO_31 (O_31,N_14298,N_14824);
xnor UO_32 (O_32,N_14417,N_14124);
or UO_33 (O_33,N_14872,N_14734);
nor UO_34 (O_34,N_14397,N_14354);
and UO_35 (O_35,N_14438,N_14960);
xnor UO_36 (O_36,N_14468,N_14836);
and UO_37 (O_37,N_14876,N_14238);
xnor UO_38 (O_38,N_14044,N_14403);
nor UO_39 (O_39,N_14323,N_14220);
and UO_40 (O_40,N_14073,N_14109);
nand UO_41 (O_41,N_14924,N_14956);
nor UO_42 (O_42,N_14411,N_14014);
and UO_43 (O_43,N_14036,N_14946);
nand UO_44 (O_44,N_14176,N_14043);
nor UO_45 (O_45,N_14843,N_14905);
nor UO_46 (O_46,N_14434,N_14198);
xnor UO_47 (O_47,N_14066,N_14413);
nor UO_48 (O_48,N_14473,N_14111);
and UO_49 (O_49,N_14973,N_14143);
or UO_50 (O_50,N_14029,N_14999);
nand UO_51 (O_51,N_14049,N_14871);
xor UO_52 (O_52,N_14979,N_14322);
or UO_53 (O_53,N_14353,N_14263);
xnor UO_54 (O_54,N_14394,N_14117);
and UO_55 (O_55,N_14334,N_14218);
nand UO_56 (O_56,N_14485,N_14395);
xor UO_57 (O_57,N_14229,N_14102);
or UO_58 (O_58,N_14521,N_14051);
or UO_59 (O_59,N_14022,N_14761);
xor UO_60 (O_60,N_14837,N_14250);
or UO_61 (O_61,N_14647,N_14457);
xor UO_62 (O_62,N_14887,N_14669);
nor UO_63 (O_63,N_14064,N_14324);
or UO_64 (O_64,N_14603,N_14551);
or UO_65 (O_65,N_14931,N_14594);
xor UO_66 (O_66,N_14104,N_14278);
and UO_67 (O_67,N_14127,N_14599);
and UO_68 (O_68,N_14577,N_14225);
xor UO_69 (O_69,N_14553,N_14161);
nor UO_70 (O_70,N_14908,N_14628);
xor UO_71 (O_71,N_14652,N_14432);
and UO_72 (O_72,N_14978,N_14646);
nor UO_73 (O_73,N_14184,N_14047);
or UO_74 (O_74,N_14620,N_14749);
xor UO_75 (O_75,N_14723,N_14453);
xnor UO_76 (O_76,N_14526,N_14018);
nand UO_77 (O_77,N_14859,N_14279);
and UO_78 (O_78,N_14063,N_14142);
nor UO_79 (O_79,N_14855,N_14788);
or UO_80 (O_80,N_14344,N_14016);
xor UO_81 (O_81,N_14748,N_14858);
nand UO_82 (O_82,N_14121,N_14820);
nor UO_83 (O_83,N_14671,N_14170);
nor UO_84 (O_84,N_14206,N_14912);
and UO_85 (O_85,N_14296,N_14307);
nor UO_86 (O_86,N_14428,N_14477);
nor UO_87 (O_87,N_14523,N_14829);
or UO_88 (O_88,N_14452,N_14420);
xor UO_89 (O_89,N_14513,N_14834);
or UO_90 (O_90,N_14705,N_14058);
nor UO_91 (O_91,N_14896,N_14284);
nor UO_92 (O_92,N_14079,N_14712);
and UO_93 (O_93,N_14498,N_14759);
nand UO_94 (O_94,N_14255,N_14556);
or UO_95 (O_95,N_14579,N_14103);
xnor UO_96 (O_96,N_14972,N_14765);
nor UO_97 (O_97,N_14164,N_14503);
or UO_98 (O_98,N_14701,N_14747);
and UO_99 (O_99,N_14001,N_14272);
and UO_100 (O_100,N_14548,N_14658);
nand UO_101 (O_101,N_14657,N_14292);
and UO_102 (O_102,N_14024,N_14329);
xor UO_103 (O_103,N_14894,N_14074);
and UO_104 (O_104,N_14787,N_14007);
and UO_105 (O_105,N_14850,N_14482);
nor UO_106 (O_106,N_14437,N_14866);
xor UO_107 (O_107,N_14729,N_14321);
xor UO_108 (O_108,N_14699,N_14550);
nand UO_109 (O_109,N_14260,N_14823);
nor UO_110 (O_110,N_14159,N_14408);
nor UO_111 (O_111,N_14731,N_14118);
and UO_112 (O_112,N_14000,N_14382);
xnor UO_113 (O_113,N_14326,N_14147);
xnor UO_114 (O_114,N_14549,N_14173);
and UO_115 (O_115,N_14727,N_14195);
nor UO_116 (O_116,N_14895,N_14409);
nand UO_117 (O_117,N_14864,N_14474);
nor UO_118 (O_118,N_14089,N_14319);
xnor UO_119 (O_119,N_14793,N_14285);
nand UO_120 (O_120,N_14480,N_14520);
or UO_121 (O_121,N_14939,N_14989);
and UO_122 (O_122,N_14318,N_14750);
nand UO_123 (O_123,N_14542,N_14138);
and UO_124 (O_124,N_14618,N_14339);
and UO_125 (O_125,N_14802,N_14181);
nand UO_126 (O_126,N_14716,N_14336);
nand UO_127 (O_127,N_14714,N_14398);
nor UO_128 (O_128,N_14226,N_14711);
nor UO_129 (O_129,N_14677,N_14707);
or UO_130 (O_130,N_14615,N_14219);
and UO_131 (O_131,N_14153,N_14174);
xnor UO_132 (O_132,N_14154,N_14691);
nor UO_133 (O_133,N_14627,N_14808);
xnor UO_134 (O_134,N_14125,N_14448);
and UO_135 (O_135,N_14958,N_14026);
nor UO_136 (O_136,N_14145,N_14270);
nand UO_137 (O_137,N_14719,N_14665);
or UO_138 (O_138,N_14688,N_14961);
and UO_139 (O_139,N_14650,N_14177);
and UO_140 (O_140,N_14767,N_14123);
nand UO_141 (O_141,N_14916,N_14032);
nand UO_142 (O_142,N_14471,N_14784);
nand UO_143 (O_143,N_14116,N_14854);
nor UO_144 (O_144,N_14466,N_14187);
or UO_145 (O_145,N_14538,N_14903);
nand UO_146 (O_146,N_14130,N_14857);
nand UO_147 (O_147,N_14289,N_14515);
nand UO_148 (O_148,N_14852,N_14088);
nor UO_149 (O_149,N_14302,N_14574);
nor UO_150 (O_150,N_14572,N_14062);
nand UO_151 (O_151,N_14132,N_14190);
nor UO_152 (O_152,N_14333,N_14060);
nand UO_153 (O_153,N_14882,N_14684);
xnor UO_154 (O_154,N_14899,N_14348);
nand UO_155 (O_155,N_14033,N_14668);
nor UO_156 (O_156,N_14672,N_14436);
xnor UO_157 (O_157,N_14945,N_14557);
and UO_158 (O_158,N_14732,N_14922);
and UO_159 (O_159,N_14287,N_14207);
xnor UO_160 (O_160,N_14569,N_14075);
and UO_161 (O_161,N_14414,N_14717);
nor UO_162 (O_162,N_14423,N_14640);
nand UO_163 (O_163,N_14743,N_14976);
nor UO_164 (O_164,N_14885,N_14721);
nor UO_165 (O_165,N_14193,N_14168);
nand UO_166 (O_166,N_14486,N_14992);
or UO_167 (O_167,N_14134,N_14197);
xor UO_168 (O_168,N_14100,N_14256);
nor UO_169 (O_169,N_14402,N_14078);
nand UO_170 (O_170,N_14421,N_14673);
or UO_171 (O_171,N_14930,N_14541);
nor UO_172 (O_172,N_14649,N_14200);
and UO_173 (O_173,N_14383,N_14391);
nand UO_174 (O_174,N_14467,N_14752);
nand UO_175 (O_175,N_14773,N_14779);
and UO_176 (O_176,N_14055,N_14634);
xor UO_177 (O_177,N_14689,N_14380);
and UO_178 (O_178,N_14863,N_14889);
and UO_179 (O_179,N_14275,N_14996);
or UO_180 (O_180,N_14442,N_14416);
nand UO_181 (O_181,N_14360,N_14487);
and UO_182 (O_182,N_14295,N_14212);
nor UO_183 (O_183,N_14347,N_14822);
or UO_184 (O_184,N_14082,N_14617);
nand UO_185 (O_185,N_14087,N_14826);
nand UO_186 (O_186,N_14410,N_14419);
nand UO_187 (O_187,N_14605,N_14372);
xnor UO_188 (O_188,N_14953,N_14936);
xor UO_189 (O_189,N_14265,N_14565);
xnor UO_190 (O_190,N_14994,N_14106);
or UO_191 (O_191,N_14479,N_14084);
and UO_192 (O_192,N_14069,N_14821);
and UO_193 (O_193,N_14811,N_14888);
and UO_194 (O_194,N_14463,N_14097);
and UO_195 (O_195,N_14806,N_14819);
or UO_196 (O_196,N_14827,N_14363);
nand UO_197 (O_197,N_14982,N_14622);
or UO_198 (O_198,N_14596,N_14578);
nand UO_199 (O_199,N_14188,N_14268);
nor UO_200 (O_200,N_14800,N_14529);
xor UO_201 (O_201,N_14968,N_14694);
nand UO_202 (O_202,N_14231,N_14795);
nand UO_203 (O_203,N_14563,N_14425);
xor UO_204 (O_204,N_14552,N_14803);
nor UO_205 (O_205,N_14180,N_14661);
or UO_206 (O_206,N_14755,N_14301);
or UO_207 (O_207,N_14445,N_14909);
nor UO_208 (O_208,N_14637,N_14744);
nand UO_209 (O_209,N_14575,N_14595);
nor UO_210 (O_210,N_14918,N_14129);
xnor UO_211 (O_211,N_14867,N_14758);
and UO_212 (O_212,N_14449,N_14757);
nor UO_213 (O_213,N_14006,N_14274);
nor UO_214 (O_214,N_14067,N_14209);
xor UO_215 (O_215,N_14257,N_14791);
nand UO_216 (O_216,N_14214,N_14966);
xnor UO_217 (O_217,N_14131,N_14775);
and UO_218 (O_218,N_14736,N_14601);
nand UO_219 (O_219,N_14861,N_14283);
and UO_220 (O_220,N_14133,N_14356);
nor UO_221 (O_221,N_14670,N_14878);
and UO_222 (O_222,N_14475,N_14273);
nand UO_223 (O_223,N_14495,N_14633);
nor UO_224 (O_224,N_14790,N_14401);
nor UO_225 (O_225,N_14352,N_14754);
and UO_226 (O_226,N_14678,N_14506);
xnor UO_227 (O_227,N_14585,N_14651);
and UO_228 (O_228,N_14804,N_14952);
and UO_229 (O_229,N_14886,N_14654);
nor UO_230 (O_230,N_14040,N_14305);
or UO_231 (O_231,N_14813,N_14253);
xor UO_232 (O_232,N_14536,N_14934);
xor UO_233 (O_233,N_14955,N_14877);
xor UO_234 (O_234,N_14110,N_14518);
nor UO_235 (O_235,N_14261,N_14848);
and UO_236 (O_236,N_14667,N_14371);
or UO_237 (O_237,N_14091,N_14555);
xnor UO_238 (O_238,N_14929,N_14582);
and UO_239 (O_239,N_14112,N_14581);
and UO_240 (O_240,N_14844,N_14681);
or UO_241 (O_241,N_14019,N_14771);
nor UO_242 (O_242,N_14306,N_14469);
xnor UO_243 (O_243,N_14722,N_14914);
nand UO_244 (O_244,N_14825,N_14208);
xor UO_245 (O_245,N_14012,N_14239);
and UO_246 (O_246,N_14810,N_14171);
nand UO_247 (O_247,N_14932,N_14898);
xnor UO_248 (O_248,N_14362,N_14962);
or UO_249 (O_249,N_14772,N_14817);
and UO_250 (O_250,N_14949,N_14404);
xor UO_251 (O_251,N_14216,N_14881);
and UO_252 (O_252,N_14057,N_14056);
and UO_253 (O_253,N_14986,N_14560);
nor UO_254 (O_254,N_14776,N_14048);
nor UO_255 (O_255,N_14135,N_14604);
nand UO_256 (O_256,N_14527,N_14777);
and UO_257 (O_257,N_14113,N_14830);
nand UO_258 (O_258,N_14258,N_14304);
and UO_259 (O_259,N_14656,N_14325);
and UO_260 (O_260,N_14798,N_14451);
or UO_261 (O_261,N_14248,N_14189);
nor UO_262 (O_262,N_14559,N_14687);
and UO_263 (O_263,N_14612,N_14144);
or UO_264 (O_264,N_14483,N_14856);
and UO_265 (O_265,N_14108,N_14162);
or UO_266 (O_266,N_14316,N_14987);
nor UO_267 (O_267,N_14023,N_14700);
or UO_268 (O_268,N_14537,N_14693);
nor UO_269 (O_269,N_14623,N_14327);
nand UO_270 (O_270,N_14114,N_14037);
and UO_271 (O_271,N_14971,N_14919);
nor UO_272 (O_272,N_14166,N_14061);
nand UO_273 (O_273,N_14464,N_14724);
nand UO_274 (O_274,N_14977,N_14025);
nor UO_275 (O_275,N_14873,N_14241);
and UO_276 (O_276,N_14959,N_14297);
or UO_277 (O_277,N_14799,N_14192);
or UO_278 (O_278,N_14481,N_14774);
and UO_279 (O_279,N_14915,N_14643);
nor UO_280 (O_280,N_14893,N_14963);
nand UO_281 (O_281,N_14429,N_14385);
and UO_282 (O_282,N_14223,N_14492);
and UO_283 (O_283,N_14708,N_14355);
nand UO_284 (O_284,N_14291,N_14373);
nand UO_285 (O_285,N_14710,N_14606);
nor UO_286 (O_286,N_14399,N_14587);
nor UO_287 (O_287,N_14892,N_14476);
nand UO_288 (O_288,N_14686,N_14756);
and UO_289 (O_289,N_14974,N_14860);
and UO_290 (O_290,N_14085,N_14509);
or UO_291 (O_291,N_14030,N_14071);
and UO_292 (O_292,N_14392,N_14342);
nand UO_293 (O_293,N_14041,N_14431);
nor UO_294 (O_294,N_14122,N_14470);
and UO_295 (O_295,N_14598,N_14443);
xor UO_296 (O_296,N_14851,N_14937);
xnor UO_297 (O_297,N_14441,N_14629);
nor UO_298 (O_298,N_14624,N_14046);
nand UO_299 (O_299,N_14516,N_14842);
or UO_300 (O_300,N_14251,N_14638);
or UO_301 (O_301,N_14094,N_14320);
or UO_302 (O_302,N_14675,N_14288);
xor UO_303 (O_303,N_14501,N_14862);
and UO_304 (O_304,N_14357,N_14092);
and UO_305 (O_305,N_14379,N_14293);
nor UO_306 (O_306,N_14910,N_14115);
or UO_307 (O_307,N_14488,N_14940);
and UO_308 (O_308,N_14739,N_14107);
xnor UO_309 (O_309,N_14796,N_14017);
and UO_310 (O_310,N_14349,N_14874);
xnor UO_311 (O_311,N_14807,N_14120);
xnor UO_312 (O_312,N_14610,N_14600);
xnor UO_313 (O_313,N_14942,N_14460);
nor UO_314 (O_314,N_14317,N_14662);
xor UO_315 (O_315,N_14614,N_14158);
and UO_316 (O_316,N_14083,N_14642);
or UO_317 (O_317,N_14227,N_14015);
and UO_318 (O_318,N_14031,N_14512);
and UO_319 (O_319,N_14228,N_14150);
nor UO_320 (O_320,N_14254,N_14493);
or UO_321 (O_321,N_14136,N_14478);
nand UO_322 (O_322,N_14653,N_14462);
xor UO_323 (O_323,N_14616,N_14619);
xnor UO_324 (O_324,N_14897,N_14237);
or UO_325 (O_325,N_14440,N_14780);
nor UO_326 (O_326,N_14718,N_14369);
and UO_327 (O_327,N_14933,N_14591);
or UO_328 (O_328,N_14222,N_14249);
nor UO_329 (O_329,N_14182,N_14126);
nand UO_330 (O_330,N_14702,N_14010);
nor UO_331 (O_331,N_14433,N_14809);
nor UO_332 (O_332,N_14835,N_14981);
xor UO_333 (O_333,N_14993,N_14586);
and UO_334 (O_334,N_14490,N_14735);
or UO_335 (O_335,N_14146,N_14002);
and UO_336 (O_336,N_14359,N_14435);
nor UO_337 (O_337,N_14186,N_14101);
or UO_338 (O_338,N_14879,N_14350);
nor UO_339 (O_339,N_14543,N_14692);
xor UO_340 (O_340,N_14020,N_14196);
nand UO_341 (O_341,N_14525,N_14762);
nor UO_342 (O_342,N_14461,N_14923);
or UO_343 (O_343,N_14011,N_14782);
nor UO_344 (O_344,N_14805,N_14309);
xor UO_345 (O_345,N_14781,N_14831);
xor UO_346 (O_346,N_14883,N_14597);
and UO_347 (O_347,N_14151,N_14328);
nor UO_348 (O_348,N_14259,N_14839);
nor UO_349 (O_349,N_14337,N_14204);
or UO_350 (O_350,N_14105,N_14390);
xnor UO_351 (O_351,N_14816,N_14814);
nor UO_352 (O_352,N_14745,N_14236);
nand UO_353 (O_353,N_14648,N_14096);
or UO_354 (O_354,N_14340,N_14853);
nor UO_355 (O_355,N_14906,N_14489);
xor UO_356 (O_356,N_14191,N_14797);
or UO_357 (O_357,N_14343,N_14008);
or UO_358 (O_358,N_14510,N_14947);
nor UO_359 (O_359,N_14430,N_14169);
or UO_360 (O_360,N_14849,N_14365);
nand UO_361 (O_361,N_14381,N_14917);
nand UO_362 (O_362,N_14611,N_14609);
or UO_363 (O_363,N_14384,N_14639);
and UO_364 (O_364,N_14841,N_14984);
xor UO_365 (O_365,N_14584,N_14003);
and UO_366 (O_366,N_14021,N_14267);
and UO_367 (O_367,N_14928,N_14454);
or UO_368 (O_368,N_14156,N_14980);
or UO_369 (O_369,N_14884,N_14738);
nand UO_370 (O_370,N_14865,N_14530);
and UO_371 (O_371,N_14312,N_14444);
nor UO_372 (O_372,N_14415,N_14346);
nor UO_373 (O_373,N_14558,N_14364);
or UO_374 (O_374,N_14967,N_14580);
or UO_375 (O_375,N_14868,N_14335);
or UO_376 (O_376,N_14472,N_14991);
or UO_377 (O_377,N_14964,N_14484);
nand UO_378 (O_378,N_14554,N_14232);
nor UO_379 (O_379,N_14792,N_14211);
or UO_380 (O_380,N_14139,N_14459);
or UO_381 (O_381,N_14965,N_14564);
or UO_382 (O_382,N_14281,N_14152);
and UO_383 (O_383,N_14300,N_14494);
and UO_384 (O_384,N_14695,N_14539);
nor UO_385 (O_385,N_14213,N_14374);
xnor UO_386 (O_386,N_14004,N_14224);
nand UO_387 (O_387,N_14446,N_14042);
or UO_388 (O_388,N_14367,N_14845);
xnor UO_389 (O_389,N_14280,N_14313);
nand UO_390 (O_390,N_14763,N_14264);
nand UO_391 (O_391,N_14499,N_14998);
or UO_392 (O_392,N_14427,N_14201);
nand UO_393 (O_393,N_14035,N_14660);
or UO_394 (O_394,N_14215,N_14240);
nand UO_395 (O_395,N_14412,N_14666);
xor UO_396 (O_396,N_14517,N_14059);
nor UO_397 (O_397,N_14244,N_14566);
and UO_398 (O_398,N_14080,N_14664);
nor UO_399 (O_399,N_14165,N_14607);
nand UO_400 (O_400,N_14098,N_14386);
nand UO_401 (O_401,N_14262,N_14140);
nand UO_402 (O_402,N_14439,N_14941);
or UO_403 (O_403,N_14065,N_14990);
xor UO_404 (O_404,N_14786,N_14210);
or UO_405 (O_405,N_14345,N_14246);
nand UO_406 (O_406,N_14641,N_14630);
and UO_407 (O_407,N_14540,N_14583);
and UO_408 (O_408,N_14050,N_14632);
or UO_409 (O_409,N_14921,N_14789);
and UO_410 (O_410,N_14715,N_14818);
or UO_411 (O_411,N_14891,N_14948);
or UO_412 (O_412,N_14593,N_14137);
nor UO_413 (O_413,N_14957,N_14400);
xnor UO_414 (O_414,N_14039,N_14706);
xnor UO_415 (O_415,N_14535,N_14674);
nand UO_416 (O_416,N_14613,N_14179);
nor UO_417 (O_417,N_14713,N_14502);
or UO_418 (O_418,N_14450,N_14422);
nand UO_419 (O_419,N_14766,N_14368);
nor UO_420 (O_420,N_14282,N_14571);
nor UO_421 (O_421,N_14072,N_14175);
or UO_422 (O_422,N_14514,N_14507);
xor UO_423 (O_423,N_14833,N_14685);
xnor UO_424 (O_424,N_14778,N_14455);
and UO_425 (O_425,N_14741,N_14663);
or UO_426 (O_426,N_14636,N_14704);
and UO_427 (O_427,N_14880,N_14005);
or UO_428 (O_428,N_14519,N_14054);
nand UO_429 (O_429,N_14217,N_14951);
nand UO_430 (O_430,N_14366,N_14242);
or UO_431 (O_431,N_14970,N_14568);
nand UO_432 (O_432,N_14625,N_14533);
nor UO_433 (O_433,N_14943,N_14682);
nor UO_434 (O_434,N_14095,N_14676);
and UO_435 (O_435,N_14038,N_14768);
or UO_436 (O_436,N_14396,N_14875);
or UO_437 (O_437,N_14985,N_14141);
nand UO_438 (O_438,N_14077,N_14266);
nor UO_439 (O_439,N_14644,N_14028);
and UO_440 (O_440,N_14053,N_14183);
nand UO_441 (O_441,N_14076,N_14303);
nand UO_442 (O_442,N_14832,N_14505);
and UO_443 (O_443,N_14160,N_14332);
nand UO_444 (O_444,N_14099,N_14690);
and UO_445 (O_445,N_14511,N_14969);
or UO_446 (O_446,N_14276,N_14753);
xnor UO_447 (O_447,N_14406,N_14308);
nand UO_448 (O_448,N_14847,N_14760);
xnor UO_449 (O_449,N_14726,N_14203);
and UO_450 (O_450,N_14068,N_14900);
and UO_451 (O_451,N_14358,N_14870);
nor UO_452 (O_452,N_14009,N_14709);
or UO_453 (O_453,N_14330,N_14562);
xnor UO_454 (O_454,N_14388,N_14194);
xor UO_455 (O_455,N_14424,N_14027);
nor UO_456 (O_456,N_14407,N_14221);
nor UO_457 (O_457,N_14045,N_14378);
or UO_458 (O_458,N_14812,N_14840);
nand UO_459 (O_459,N_14172,N_14052);
or UO_460 (O_460,N_14090,N_14728);
or UO_461 (O_461,N_14252,N_14496);
xnor UO_462 (O_462,N_14570,N_14950);
and UO_463 (O_463,N_14720,N_14547);
nor UO_464 (O_464,N_14935,N_14683);
nor UO_465 (O_465,N_14119,N_14081);
nand UO_466 (O_466,N_14679,N_14954);
nor UO_467 (O_467,N_14389,N_14522);
nor UO_468 (O_468,N_14157,N_14167);
nand UO_469 (O_469,N_14975,N_14163);
nand UO_470 (O_470,N_14331,N_14426);
xnor UO_471 (O_471,N_14801,N_14573);
nor UO_472 (O_472,N_14447,N_14532);
nor UO_473 (O_473,N_14233,N_14828);
and UO_474 (O_474,N_14205,N_14178);
xnor UO_475 (O_475,N_14545,N_14269);
and UO_476 (O_476,N_14902,N_14907);
xnor UO_477 (O_477,N_14376,N_14299);
nor UO_478 (O_478,N_14938,N_14271);
xnor UO_479 (O_479,N_14341,N_14310);
or UO_480 (O_480,N_14697,N_14696);
nand UO_481 (O_481,N_14243,N_14769);
xor UO_482 (O_482,N_14128,N_14294);
xnor UO_483 (O_483,N_14277,N_14247);
and UO_484 (O_484,N_14093,N_14286);
or UO_485 (O_485,N_14783,N_14013);
xor UO_486 (O_486,N_14944,N_14631);
nor UO_487 (O_487,N_14659,N_14034);
nand UO_488 (O_488,N_14751,N_14730);
and UO_489 (O_489,N_14234,N_14375);
nor UO_490 (O_490,N_14838,N_14524);
or UO_491 (O_491,N_14588,N_14290);
and UO_492 (O_492,N_14202,N_14927);
nor UO_493 (O_493,N_14995,N_14742);
and UO_494 (O_494,N_14561,N_14070);
nor UO_495 (O_495,N_14890,N_14361);
and UO_496 (O_496,N_14465,N_14621);
xor UO_497 (O_497,N_14418,N_14589);
nand UO_498 (O_498,N_14920,N_14725);
and UO_499 (O_499,N_14733,N_14764);
xor UO_500 (O_500,N_14467,N_14595);
nor UO_501 (O_501,N_14418,N_14331);
nand UO_502 (O_502,N_14161,N_14481);
or UO_503 (O_503,N_14297,N_14917);
nand UO_504 (O_504,N_14742,N_14111);
or UO_505 (O_505,N_14049,N_14545);
nand UO_506 (O_506,N_14345,N_14763);
or UO_507 (O_507,N_14222,N_14073);
xor UO_508 (O_508,N_14147,N_14672);
nor UO_509 (O_509,N_14487,N_14346);
or UO_510 (O_510,N_14555,N_14356);
nand UO_511 (O_511,N_14110,N_14926);
nand UO_512 (O_512,N_14044,N_14948);
or UO_513 (O_513,N_14800,N_14452);
xor UO_514 (O_514,N_14429,N_14986);
xor UO_515 (O_515,N_14260,N_14423);
or UO_516 (O_516,N_14601,N_14009);
nor UO_517 (O_517,N_14837,N_14126);
or UO_518 (O_518,N_14172,N_14123);
and UO_519 (O_519,N_14848,N_14906);
and UO_520 (O_520,N_14732,N_14929);
and UO_521 (O_521,N_14798,N_14336);
nand UO_522 (O_522,N_14135,N_14374);
nor UO_523 (O_523,N_14997,N_14286);
or UO_524 (O_524,N_14506,N_14209);
xor UO_525 (O_525,N_14607,N_14619);
nor UO_526 (O_526,N_14076,N_14986);
xnor UO_527 (O_527,N_14109,N_14071);
xor UO_528 (O_528,N_14384,N_14214);
and UO_529 (O_529,N_14446,N_14708);
or UO_530 (O_530,N_14190,N_14116);
xor UO_531 (O_531,N_14784,N_14664);
nor UO_532 (O_532,N_14424,N_14968);
nor UO_533 (O_533,N_14539,N_14282);
nand UO_534 (O_534,N_14373,N_14008);
xnor UO_535 (O_535,N_14985,N_14348);
xor UO_536 (O_536,N_14166,N_14828);
nand UO_537 (O_537,N_14783,N_14264);
nand UO_538 (O_538,N_14603,N_14420);
xor UO_539 (O_539,N_14893,N_14878);
nor UO_540 (O_540,N_14391,N_14583);
or UO_541 (O_541,N_14589,N_14391);
xor UO_542 (O_542,N_14434,N_14685);
or UO_543 (O_543,N_14385,N_14089);
and UO_544 (O_544,N_14380,N_14056);
and UO_545 (O_545,N_14461,N_14130);
nand UO_546 (O_546,N_14747,N_14913);
xnor UO_547 (O_547,N_14943,N_14326);
or UO_548 (O_548,N_14059,N_14592);
nand UO_549 (O_549,N_14789,N_14911);
xnor UO_550 (O_550,N_14453,N_14433);
xnor UO_551 (O_551,N_14011,N_14439);
and UO_552 (O_552,N_14199,N_14809);
xor UO_553 (O_553,N_14855,N_14660);
xnor UO_554 (O_554,N_14236,N_14984);
and UO_555 (O_555,N_14747,N_14154);
xnor UO_556 (O_556,N_14436,N_14854);
or UO_557 (O_557,N_14324,N_14055);
xor UO_558 (O_558,N_14905,N_14068);
xnor UO_559 (O_559,N_14000,N_14202);
or UO_560 (O_560,N_14104,N_14130);
or UO_561 (O_561,N_14553,N_14746);
xor UO_562 (O_562,N_14366,N_14388);
or UO_563 (O_563,N_14975,N_14230);
or UO_564 (O_564,N_14293,N_14284);
and UO_565 (O_565,N_14381,N_14793);
xor UO_566 (O_566,N_14016,N_14004);
and UO_567 (O_567,N_14158,N_14359);
nor UO_568 (O_568,N_14634,N_14677);
or UO_569 (O_569,N_14358,N_14334);
xnor UO_570 (O_570,N_14840,N_14222);
xor UO_571 (O_571,N_14286,N_14491);
xnor UO_572 (O_572,N_14141,N_14686);
nor UO_573 (O_573,N_14812,N_14517);
xor UO_574 (O_574,N_14152,N_14469);
xor UO_575 (O_575,N_14008,N_14586);
and UO_576 (O_576,N_14615,N_14840);
nand UO_577 (O_577,N_14389,N_14007);
and UO_578 (O_578,N_14879,N_14622);
nor UO_579 (O_579,N_14376,N_14921);
nor UO_580 (O_580,N_14991,N_14301);
nor UO_581 (O_581,N_14274,N_14791);
nand UO_582 (O_582,N_14956,N_14279);
and UO_583 (O_583,N_14152,N_14022);
and UO_584 (O_584,N_14448,N_14323);
nor UO_585 (O_585,N_14781,N_14906);
nand UO_586 (O_586,N_14381,N_14368);
nor UO_587 (O_587,N_14148,N_14730);
nor UO_588 (O_588,N_14911,N_14799);
or UO_589 (O_589,N_14642,N_14413);
and UO_590 (O_590,N_14266,N_14862);
or UO_591 (O_591,N_14595,N_14859);
or UO_592 (O_592,N_14122,N_14705);
and UO_593 (O_593,N_14861,N_14161);
xnor UO_594 (O_594,N_14495,N_14487);
xnor UO_595 (O_595,N_14549,N_14795);
xnor UO_596 (O_596,N_14792,N_14418);
nand UO_597 (O_597,N_14806,N_14392);
and UO_598 (O_598,N_14079,N_14504);
or UO_599 (O_599,N_14449,N_14288);
or UO_600 (O_600,N_14355,N_14249);
nand UO_601 (O_601,N_14424,N_14400);
and UO_602 (O_602,N_14699,N_14152);
nand UO_603 (O_603,N_14199,N_14429);
xnor UO_604 (O_604,N_14894,N_14724);
xor UO_605 (O_605,N_14254,N_14761);
nor UO_606 (O_606,N_14049,N_14025);
nor UO_607 (O_607,N_14094,N_14043);
and UO_608 (O_608,N_14919,N_14236);
xnor UO_609 (O_609,N_14313,N_14500);
or UO_610 (O_610,N_14120,N_14972);
nor UO_611 (O_611,N_14682,N_14021);
xnor UO_612 (O_612,N_14720,N_14662);
xor UO_613 (O_613,N_14256,N_14157);
nor UO_614 (O_614,N_14600,N_14853);
xor UO_615 (O_615,N_14165,N_14450);
or UO_616 (O_616,N_14056,N_14038);
nor UO_617 (O_617,N_14891,N_14523);
nor UO_618 (O_618,N_14454,N_14862);
nand UO_619 (O_619,N_14875,N_14823);
or UO_620 (O_620,N_14349,N_14044);
nor UO_621 (O_621,N_14235,N_14441);
nor UO_622 (O_622,N_14066,N_14776);
or UO_623 (O_623,N_14517,N_14390);
nand UO_624 (O_624,N_14142,N_14575);
nand UO_625 (O_625,N_14285,N_14312);
and UO_626 (O_626,N_14627,N_14764);
xnor UO_627 (O_627,N_14773,N_14495);
or UO_628 (O_628,N_14237,N_14971);
and UO_629 (O_629,N_14764,N_14794);
nand UO_630 (O_630,N_14242,N_14108);
nor UO_631 (O_631,N_14713,N_14369);
xor UO_632 (O_632,N_14623,N_14034);
or UO_633 (O_633,N_14540,N_14298);
nor UO_634 (O_634,N_14362,N_14099);
and UO_635 (O_635,N_14816,N_14684);
and UO_636 (O_636,N_14372,N_14166);
nand UO_637 (O_637,N_14212,N_14005);
nand UO_638 (O_638,N_14394,N_14153);
nor UO_639 (O_639,N_14401,N_14519);
and UO_640 (O_640,N_14542,N_14496);
nand UO_641 (O_641,N_14700,N_14995);
xnor UO_642 (O_642,N_14981,N_14260);
or UO_643 (O_643,N_14655,N_14236);
nor UO_644 (O_644,N_14042,N_14867);
nor UO_645 (O_645,N_14190,N_14083);
nand UO_646 (O_646,N_14842,N_14723);
xnor UO_647 (O_647,N_14749,N_14023);
nand UO_648 (O_648,N_14639,N_14373);
nand UO_649 (O_649,N_14566,N_14856);
xor UO_650 (O_650,N_14641,N_14505);
and UO_651 (O_651,N_14226,N_14698);
nand UO_652 (O_652,N_14783,N_14424);
and UO_653 (O_653,N_14992,N_14913);
and UO_654 (O_654,N_14792,N_14311);
nand UO_655 (O_655,N_14486,N_14380);
nor UO_656 (O_656,N_14948,N_14563);
nor UO_657 (O_657,N_14611,N_14185);
nor UO_658 (O_658,N_14736,N_14585);
or UO_659 (O_659,N_14190,N_14668);
xnor UO_660 (O_660,N_14932,N_14965);
nand UO_661 (O_661,N_14746,N_14035);
and UO_662 (O_662,N_14141,N_14241);
or UO_663 (O_663,N_14024,N_14625);
or UO_664 (O_664,N_14229,N_14967);
and UO_665 (O_665,N_14609,N_14546);
and UO_666 (O_666,N_14305,N_14855);
xor UO_667 (O_667,N_14362,N_14922);
nand UO_668 (O_668,N_14868,N_14608);
nand UO_669 (O_669,N_14381,N_14502);
or UO_670 (O_670,N_14584,N_14539);
xnor UO_671 (O_671,N_14559,N_14656);
and UO_672 (O_672,N_14205,N_14436);
nand UO_673 (O_673,N_14030,N_14913);
xnor UO_674 (O_674,N_14136,N_14958);
xnor UO_675 (O_675,N_14469,N_14874);
xor UO_676 (O_676,N_14885,N_14243);
or UO_677 (O_677,N_14938,N_14431);
nor UO_678 (O_678,N_14763,N_14822);
xnor UO_679 (O_679,N_14919,N_14463);
nor UO_680 (O_680,N_14944,N_14079);
and UO_681 (O_681,N_14470,N_14217);
and UO_682 (O_682,N_14960,N_14187);
xor UO_683 (O_683,N_14431,N_14694);
or UO_684 (O_684,N_14723,N_14477);
and UO_685 (O_685,N_14907,N_14240);
nand UO_686 (O_686,N_14956,N_14192);
nand UO_687 (O_687,N_14528,N_14635);
xor UO_688 (O_688,N_14472,N_14037);
xor UO_689 (O_689,N_14400,N_14192);
and UO_690 (O_690,N_14597,N_14441);
or UO_691 (O_691,N_14181,N_14232);
and UO_692 (O_692,N_14593,N_14419);
or UO_693 (O_693,N_14593,N_14816);
nand UO_694 (O_694,N_14146,N_14196);
xor UO_695 (O_695,N_14892,N_14994);
nand UO_696 (O_696,N_14252,N_14843);
or UO_697 (O_697,N_14721,N_14733);
or UO_698 (O_698,N_14121,N_14955);
and UO_699 (O_699,N_14235,N_14461);
nand UO_700 (O_700,N_14294,N_14758);
or UO_701 (O_701,N_14294,N_14015);
xor UO_702 (O_702,N_14022,N_14275);
nor UO_703 (O_703,N_14197,N_14680);
or UO_704 (O_704,N_14619,N_14068);
xor UO_705 (O_705,N_14053,N_14490);
nor UO_706 (O_706,N_14873,N_14064);
nor UO_707 (O_707,N_14803,N_14254);
xnor UO_708 (O_708,N_14830,N_14844);
or UO_709 (O_709,N_14973,N_14819);
or UO_710 (O_710,N_14323,N_14057);
xor UO_711 (O_711,N_14337,N_14401);
nor UO_712 (O_712,N_14731,N_14440);
or UO_713 (O_713,N_14971,N_14432);
nand UO_714 (O_714,N_14394,N_14912);
or UO_715 (O_715,N_14357,N_14928);
xor UO_716 (O_716,N_14688,N_14455);
or UO_717 (O_717,N_14493,N_14837);
nor UO_718 (O_718,N_14859,N_14519);
or UO_719 (O_719,N_14637,N_14167);
nor UO_720 (O_720,N_14366,N_14890);
nand UO_721 (O_721,N_14458,N_14597);
nor UO_722 (O_722,N_14745,N_14408);
and UO_723 (O_723,N_14643,N_14613);
and UO_724 (O_724,N_14012,N_14102);
nand UO_725 (O_725,N_14609,N_14807);
xnor UO_726 (O_726,N_14303,N_14970);
or UO_727 (O_727,N_14787,N_14308);
xor UO_728 (O_728,N_14346,N_14794);
xnor UO_729 (O_729,N_14974,N_14328);
and UO_730 (O_730,N_14358,N_14142);
xor UO_731 (O_731,N_14599,N_14151);
and UO_732 (O_732,N_14164,N_14887);
nand UO_733 (O_733,N_14381,N_14986);
nor UO_734 (O_734,N_14867,N_14712);
nor UO_735 (O_735,N_14587,N_14117);
nor UO_736 (O_736,N_14786,N_14137);
or UO_737 (O_737,N_14329,N_14542);
nand UO_738 (O_738,N_14726,N_14979);
or UO_739 (O_739,N_14893,N_14097);
nand UO_740 (O_740,N_14366,N_14202);
or UO_741 (O_741,N_14498,N_14519);
and UO_742 (O_742,N_14136,N_14464);
nor UO_743 (O_743,N_14882,N_14850);
xor UO_744 (O_744,N_14451,N_14858);
xnor UO_745 (O_745,N_14803,N_14102);
xnor UO_746 (O_746,N_14298,N_14637);
nor UO_747 (O_747,N_14834,N_14855);
or UO_748 (O_748,N_14111,N_14485);
nand UO_749 (O_749,N_14142,N_14020);
xor UO_750 (O_750,N_14253,N_14606);
and UO_751 (O_751,N_14337,N_14497);
and UO_752 (O_752,N_14487,N_14931);
or UO_753 (O_753,N_14203,N_14784);
nor UO_754 (O_754,N_14794,N_14962);
or UO_755 (O_755,N_14282,N_14900);
or UO_756 (O_756,N_14760,N_14002);
xor UO_757 (O_757,N_14005,N_14967);
xor UO_758 (O_758,N_14146,N_14327);
nor UO_759 (O_759,N_14182,N_14803);
nand UO_760 (O_760,N_14356,N_14343);
xor UO_761 (O_761,N_14424,N_14325);
nor UO_762 (O_762,N_14539,N_14525);
xnor UO_763 (O_763,N_14976,N_14132);
nand UO_764 (O_764,N_14139,N_14664);
nand UO_765 (O_765,N_14349,N_14781);
and UO_766 (O_766,N_14085,N_14781);
xnor UO_767 (O_767,N_14310,N_14012);
xnor UO_768 (O_768,N_14461,N_14249);
and UO_769 (O_769,N_14594,N_14828);
xor UO_770 (O_770,N_14378,N_14256);
nand UO_771 (O_771,N_14771,N_14858);
nand UO_772 (O_772,N_14265,N_14931);
and UO_773 (O_773,N_14070,N_14953);
nor UO_774 (O_774,N_14146,N_14884);
and UO_775 (O_775,N_14643,N_14587);
or UO_776 (O_776,N_14164,N_14069);
nor UO_777 (O_777,N_14903,N_14436);
xor UO_778 (O_778,N_14526,N_14493);
nor UO_779 (O_779,N_14813,N_14720);
and UO_780 (O_780,N_14860,N_14196);
xnor UO_781 (O_781,N_14937,N_14637);
and UO_782 (O_782,N_14007,N_14667);
and UO_783 (O_783,N_14888,N_14137);
and UO_784 (O_784,N_14001,N_14370);
nand UO_785 (O_785,N_14160,N_14511);
nor UO_786 (O_786,N_14759,N_14645);
nor UO_787 (O_787,N_14706,N_14325);
xor UO_788 (O_788,N_14357,N_14177);
xor UO_789 (O_789,N_14549,N_14028);
or UO_790 (O_790,N_14600,N_14142);
xnor UO_791 (O_791,N_14499,N_14819);
or UO_792 (O_792,N_14473,N_14791);
nand UO_793 (O_793,N_14358,N_14630);
nor UO_794 (O_794,N_14367,N_14594);
and UO_795 (O_795,N_14220,N_14142);
nor UO_796 (O_796,N_14058,N_14940);
and UO_797 (O_797,N_14001,N_14398);
xor UO_798 (O_798,N_14550,N_14898);
and UO_799 (O_799,N_14791,N_14134);
nand UO_800 (O_800,N_14156,N_14764);
and UO_801 (O_801,N_14220,N_14692);
nor UO_802 (O_802,N_14426,N_14703);
nand UO_803 (O_803,N_14592,N_14629);
nand UO_804 (O_804,N_14544,N_14803);
nor UO_805 (O_805,N_14001,N_14774);
nor UO_806 (O_806,N_14085,N_14248);
nand UO_807 (O_807,N_14156,N_14921);
nand UO_808 (O_808,N_14231,N_14173);
or UO_809 (O_809,N_14565,N_14800);
and UO_810 (O_810,N_14250,N_14402);
nor UO_811 (O_811,N_14163,N_14646);
and UO_812 (O_812,N_14649,N_14494);
and UO_813 (O_813,N_14621,N_14303);
and UO_814 (O_814,N_14277,N_14419);
or UO_815 (O_815,N_14707,N_14070);
nor UO_816 (O_816,N_14736,N_14176);
nor UO_817 (O_817,N_14427,N_14963);
nor UO_818 (O_818,N_14116,N_14128);
or UO_819 (O_819,N_14941,N_14896);
nand UO_820 (O_820,N_14249,N_14635);
and UO_821 (O_821,N_14092,N_14286);
xor UO_822 (O_822,N_14969,N_14685);
xor UO_823 (O_823,N_14208,N_14109);
nor UO_824 (O_824,N_14325,N_14387);
and UO_825 (O_825,N_14098,N_14192);
nand UO_826 (O_826,N_14252,N_14065);
or UO_827 (O_827,N_14578,N_14192);
or UO_828 (O_828,N_14177,N_14008);
and UO_829 (O_829,N_14664,N_14429);
nor UO_830 (O_830,N_14727,N_14685);
nor UO_831 (O_831,N_14908,N_14380);
xor UO_832 (O_832,N_14176,N_14778);
xor UO_833 (O_833,N_14872,N_14504);
nand UO_834 (O_834,N_14067,N_14235);
nand UO_835 (O_835,N_14477,N_14256);
or UO_836 (O_836,N_14781,N_14463);
and UO_837 (O_837,N_14015,N_14899);
nand UO_838 (O_838,N_14208,N_14643);
nand UO_839 (O_839,N_14346,N_14867);
or UO_840 (O_840,N_14683,N_14317);
nor UO_841 (O_841,N_14686,N_14916);
xor UO_842 (O_842,N_14288,N_14907);
nor UO_843 (O_843,N_14073,N_14216);
nor UO_844 (O_844,N_14815,N_14293);
and UO_845 (O_845,N_14400,N_14574);
nand UO_846 (O_846,N_14047,N_14898);
xor UO_847 (O_847,N_14681,N_14472);
nand UO_848 (O_848,N_14697,N_14561);
xnor UO_849 (O_849,N_14249,N_14712);
nor UO_850 (O_850,N_14553,N_14463);
and UO_851 (O_851,N_14657,N_14648);
nand UO_852 (O_852,N_14293,N_14383);
xnor UO_853 (O_853,N_14349,N_14208);
and UO_854 (O_854,N_14461,N_14365);
or UO_855 (O_855,N_14595,N_14707);
nand UO_856 (O_856,N_14820,N_14754);
nor UO_857 (O_857,N_14396,N_14937);
nor UO_858 (O_858,N_14171,N_14816);
xor UO_859 (O_859,N_14986,N_14033);
or UO_860 (O_860,N_14752,N_14965);
and UO_861 (O_861,N_14975,N_14137);
nor UO_862 (O_862,N_14292,N_14523);
xnor UO_863 (O_863,N_14545,N_14839);
nand UO_864 (O_864,N_14361,N_14224);
and UO_865 (O_865,N_14647,N_14935);
or UO_866 (O_866,N_14338,N_14668);
and UO_867 (O_867,N_14583,N_14767);
xnor UO_868 (O_868,N_14665,N_14395);
xor UO_869 (O_869,N_14485,N_14551);
xnor UO_870 (O_870,N_14912,N_14004);
and UO_871 (O_871,N_14218,N_14835);
xnor UO_872 (O_872,N_14398,N_14000);
nand UO_873 (O_873,N_14295,N_14043);
nand UO_874 (O_874,N_14156,N_14025);
or UO_875 (O_875,N_14657,N_14760);
xor UO_876 (O_876,N_14594,N_14250);
nor UO_877 (O_877,N_14466,N_14207);
and UO_878 (O_878,N_14686,N_14459);
or UO_879 (O_879,N_14226,N_14209);
xnor UO_880 (O_880,N_14027,N_14616);
nor UO_881 (O_881,N_14121,N_14281);
and UO_882 (O_882,N_14096,N_14401);
nor UO_883 (O_883,N_14618,N_14133);
nand UO_884 (O_884,N_14732,N_14428);
or UO_885 (O_885,N_14551,N_14896);
nand UO_886 (O_886,N_14503,N_14548);
xnor UO_887 (O_887,N_14337,N_14200);
nor UO_888 (O_888,N_14216,N_14145);
and UO_889 (O_889,N_14719,N_14132);
nor UO_890 (O_890,N_14315,N_14128);
and UO_891 (O_891,N_14063,N_14519);
nand UO_892 (O_892,N_14839,N_14962);
nand UO_893 (O_893,N_14811,N_14309);
xnor UO_894 (O_894,N_14738,N_14312);
or UO_895 (O_895,N_14893,N_14233);
and UO_896 (O_896,N_14626,N_14093);
nor UO_897 (O_897,N_14969,N_14255);
or UO_898 (O_898,N_14268,N_14504);
xnor UO_899 (O_899,N_14108,N_14283);
xnor UO_900 (O_900,N_14518,N_14140);
xnor UO_901 (O_901,N_14828,N_14152);
nand UO_902 (O_902,N_14466,N_14746);
and UO_903 (O_903,N_14674,N_14361);
xor UO_904 (O_904,N_14630,N_14275);
or UO_905 (O_905,N_14642,N_14399);
nor UO_906 (O_906,N_14081,N_14677);
or UO_907 (O_907,N_14235,N_14933);
and UO_908 (O_908,N_14874,N_14140);
and UO_909 (O_909,N_14223,N_14826);
or UO_910 (O_910,N_14616,N_14605);
xor UO_911 (O_911,N_14085,N_14511);
and UO_912 (O_912,N_14513,N_14324);
nand UO_913 (O_913,N_14471,N_14993);
nand UO_914 (O_914,N_14821,N_14439);
xnor UO_915 (O_915,N_14287,N_14090);
or UO_916 (O_916,N_14253,N_14831);
xor UO_917 (O_917,N_14695,N_14809);
nor UO_918 (O_918,N_14897,N_14354);
or UO_919 (O_919,N_14169,N_14654);
or UO_920 (O_920,N_14636,N_14303);
or UO_921 (O_921,N_14924,N_14504);
or UO_922 (O_922,N_14054,N_14133);
and UO_923 (O_923,N_14501,N_14574);
and UO_924 (O_924,N_14960,N_14502);
xor UO_925 (O_925,N_14639,N_14771);
and UO_926 (O_926,N_14192,N_14132);
nor UO_927 (O_927,N_14193,N_14943);
nand UO_928 (O_928,N_14841,N_14589);
xnor UO_929 (O_929,N_14357,N_14408);
nand UO_930 (O_930,N_14329,N_14119);
nor UO_931 (O_931,N_14270,N_14573);
nand UO_932 (O_932,N_14231,N_14188);
nor UO_933 (O_933,N_14786,N_14934);
xor UO_934 (O_934,N_14447,N_14411);
and UO_935 (O_935,N_14325,N_14670);
or UO_936 (O_936,N_14203,N_14283);
nor UO_937 (O_937,N_14165,N_14269);
nand UO_938 (O_938,N_14196,N_14852);
xnor UO_939 (O_939,N_14749,N_14832);
nand UO_940 (O_940,N_14858,N_14880);
nor UO_941 (O_941,N_14946,N_14184);
nor UO_942 (O_942,N_14044,N_14945);
xor UO_943 (O_943,N_14416,N_14650);
xnor UO_944 (O_944,N_14587,N_14993);
xor UO_945 (O_945,N_14539,N_14198);
xnor UO_946 (O_946,N_14805,N_14377);
xnor UO_947 (O_947,N_14741,N_14817);
nor UO_948 (O_948,N_14878,N_14760);
xor UO_949 (O_949,N_14733,N_14885);
and UO_950 (O_950,N_14634,N_14727);
nor UO_951 (O_951,N_14730,N_14032);
and UO_952 (O_952,N_14378,N_14152);
nand UO_953 (O_953,N_14555,N_14718);
nor UO_954 (O_954,N_14484,N_14140);
xnor UO_955 (O_955,N_14191,N_14992);
and UO_956 (O_956,N_14772,N_14679);
nand UO_957 (O_957,N_14378,N_14060);
or UO_958 (O_958,N_14260,N_14658);
xor UO_959 (O_959,N_14556,N_14059);
nor UO_960 (O_960,N_14183,N_14697);
nand UO_961 (O_961,N_14149,N_14654);
or UO_962 (O_962,N_14882,N_14852);
or UO_963 (O_963,N_14489,N_14305);
nor UO_964 (O_964,N_14642,N_14975);
xor UO_965 (O_965,N_14993,N_14754);
or UO_966 (O_966,N_14155,N_14552);
nand UO_967 (O_967,N_14183,N_14399);
nor UO_968 (O_968,N_14933,N_14490);
nand UO_969 (O_969,N_14816,N_14602);
or UO_970 (O_970,N_14412,N_14575);
or UO_971 (O_971,N_14586,N_14188);
nor UO_972 (O_972,N_14144,N_14997);
or UO_973 (O_973,N_14646,N_14820);
nand UO_974 (O_974,N_14910,N_14978);
and UO_975 (O_975,N_14452,N_14446);
nand UO_976 (O_976,N_14791,N_14579);
nor UO_977 (O_977,N_14074,N_14951);
nor UO_978 (O_978,N_14539,N_14360);
or UO_979 (O_979,N_14040,N_14706);
nor UO_980 (O_980,N_14535,N_14928);
and UO_981 (O_981,N_14884,N_14814);
nor UO_982 (O_982,N_14382,N_14136);
and UO_983 (O_983,N_14365,N_14574);
nor UO_984 (O_984,N_14080,N_14742);
nor UO_985 (O_985,N_14475,N_14657);
nand UO_986 (O_986,N_14153,N_14192);
or UO_987 (O_987,N_14853,N_14875);
xnor UO_988 (O_988,N_14724,N_14768);
xor UO_989 (O_989,N_14769,N_14716);
or UO_990 (O_990,N_14074,N_14765);
xor UO_991 (O_991,N_14229,N_14649);
nor UO_992 (O_992,N_14843,N_14256);
xnor UO_993 (O_993,N_14013,N_14531);
or UO_994 (O_994,N_14453,N_14466);
nor UO_995 (O_995,N_14923,N_14651);
and UO_996 (O_996,N_14489,N_14110);
and UO_997 (O_997,N_14751,N_14069);
and UO_998 (O_998,N_14910,N_14612);
nor UO_999 (O_999,N_14281,N_14609);
nand UO_1000 (O_1000,N_14547,N_14180);
or UO_1001 (O_1001,N_14490,N_14228);
or UO_1002 (O_1002,N_14928,N_14851);
or UO_1003 (O_1003,N_14289,N_14718);
nor UO_1004 (O_1004,N_14373,N_14245);
nor UO_1005 (O_1005,N_14897,N_14298);
nand UO_1006 (O_1006,N_14261,N_14820);
nand UO_1007 (O_1007,N_14795,N_14285);
xor UO_1008 (O_1008,N_14989,N_14250);
and UO_1009 (O_1009,N_14591,N_14815);
and UO_1010 (O_1010,N_14988,N_14465);
and UO_1011 (O_1011,N_14887,N_14737);
nand UO_1012 (O_1012,N_14931,N_14694);
nand UO_1013 (O_1013,N_14125,N_14095);
nand UO_1014 (O_1014,N_14787,N_14724);
nand UO_1015 (O_1015,N_14096,N_14510);
and UO_1016 (O_1016,N_14318,N_14265);
xnor UO_1017 (O_1017,N_14996,N_14112);
nand UO_1018 (O_1018,N_14868,N_14920);
or UO_1019 (O_1019,N_14830,N_14039);
nand UO_1020 (O_1020,N_14859,N_14477);
or UO_1021 (O_1021,N_14123,N_14207);
or UO_1022 (O_1022,N_14362,N_14075);
nand UO_1023 (O_1023,N_14593,N_14110);
or UO_1024 (O_1024,N_14637,N_14241);
or UO_1025 (O_1025,N_14275,N_14043);
xor UO_1026 (O_1026,N_14033,N_14182);
nor UO_1027 (O_1027,N_14697,N_14551);
or UO_1028 (O_1028,N_14378,N_14384);
nor UO_1029 (O_1029,N_14766,N_14953);
or UO_1030 (O_1030,N_14248,N_14132);
and UO_1031 (O_1031,N_14692,N_14102);
or UO_1032 (O_1032,N_14599,N_14839);
xor UO_1033 (O_1033,N_14763,N_14261);
or UO_1034 (O_1034,N_14415,N_14282);
nand UO_1035 (O_1035,N_14084,N_14473);
or UO_1036 (O_1036,N_14716,N_14043);
nor UO_1037 (O_1037,N_14823,N_14613);
nor UO_1038 (O_1038,N_14133,N_14763);
nand UO_1039 (O_1039,N_14429,N_14298);
nor UO_1040 (O_1040,N_14767,N_14703);
xnor UO_1041 (O_1041,N_14695,N_14093);
and UO_1042 (O_1042,N_14301,N_14070);
or UO_1043 (O_1043,N_14186,N_14034);
nand UO_1044 (O_1044,N_14573,N_14435);
nand UO_1045 (O_1045,N_14403,N_14531);
xnor UO_1046 (O_1046,N_14236,N_14458);
nand UO_1047 (O_1047,N_14542,N_14168);
and UO_1048 (O_1048,N_14241,N_14167);
and UO_1049 (O_1049,N_14689,N_14835);
xor UO_1050 (O_1050,N_14326,N_14786);
xnor UO_1051 (O_1051,N_14414,N_14564);
or UO_1052 (O_1052,N_14914,N_14317);
nand UO_1053 (O_1053,N_14661,N_14732);
nand UO_1054 (O_1054,N_14079,N_14790);
nor UO_1055 (O_1055,N_14660,N_14964);
and UO_1056 (O_1056,N_14818,N_14629);
nor UO_1057 (O_1057,N_14337,N_14959);
and UO_1058 (O_1058,N_14688,N_14869);
nor UO_1059 (O_1059,N_14724,N_14977);
nor UO_1060 (O_1060,N_14169,N_14235);
xnor UO_1061 (O_1061,N_14992,N_14864);
nand UO_1062 (O_1062,N_14119,N_14687);
xnor UO_1063 (O_1063,N_14289,N_14599);
xor UO_1064 (O_1064,N_14393,N_14167);
nor UO_1065 (O_1065,N_14947,N_14136);
nand UO_1066 (O_1066,N_14221,N_14011);
nor UO_1067 (O_1067,N_14813,N_14761);
nor UO_1068 (O_1068,N_14742,N_14302);
or UO_1069 (O_1069,N_14307,N_14499);
or UO_1070 (O_1070,N_14517,N_14727);
and UO_1071 (O_1071,N_14504,N_14226);
and UO_1072 (O_1072,N_14400,N_14114);
or UO_1073 (O_1073,N_14635,N_14022);
nor UO_1074 (O_1074,N_14156,N_14879);
nand UO_1075 (O_1075,N_14278,N_14898);
or UO_1076 (O_1076,N_14004,N_14716);
xnor UO_1077 (O_1077,N_14651,N_14000);
nor UO_1078 (O_1078,N_14570,N_14284);
nand UO_1079 (O_1079,N_14339,N_14850);
or UO_1080 (O_1080,N_14602,N_14383);
or UO_1081 (O_1081,N_14455,N_14433);
or UO_1082 (O_1082,N_14029,N_14333);
nor UO_1083 (O_1083,N_14977,N_14364);
nor UO_1084 (O_1084,N_14210,N_14064);
and UO_1085 (O_1085,N_14063,N_14093);
or UO_1086 (O_1086,N_14975,N_14686);
and UO_1087 (O_1087,N_14234,N_14795);
nand UO_1088 (O_1088,N_14788,N_14384);
nand UO_1089 (O_1089,N_14156,N_14478);
and UO_1090 (O_1090,N_14084,N_14591);
or UO_1091 (O_1091,N_14406,N_14810);
nand UO_1092 (O_1092,N_14502,N_14499);
nor UO_1093 (O_1093,N_14037,N_14624);
or UO_1094 (O_1094,N_14714,N_14625);
or UO_1095 (O_1095,N_14148,N_14591);
nor UO_1096 (O_1096,N_14616,N_14279);
or UO_1097 (O_1097,N_14625,N_14300);
xnor UO_1098 (O_1098,N_14692,N_14669);
and UO_1099 (O_1099,N_14029,N_14082);
xnor UO_1100 (O_1100,N_14395,N_14402);
and UO_1101 (O_1101,N_14359,N_14711);
nor UO_1102 (O_1102,N_14059,N_14770);
xnor UO_1103 (O_1103,N_14915,N_14173);
and UO_1104 (O_1104,N_14256,N_14263);
or UO_1105 (O_1105,N_14366,N_14204);
and UO_1106 (O_1106,N_14864,N_14970);
or UO_1107 (O_1107,N_14467,N_14084);
or UO_1108 (O_1108,N_14094,N_14099);
nor UO_1109 (O_1109,N_14947,N_14235);
and UO_1110 (O_1110,N_14465,N_14810);
nand UO_1111 (O_1111,N_14077,N_14634);
and UO_1112 (O_1112,N_14966,N_14203);
nand UO_1113 (O_1113,N_14068,N_14823);
xnor UO_1114 (O_1114,N_14778,N_14853);
and UO_1115 (O_1115,N_14336,N_14879);
xnor UO_1116 (O_1116,N_14325,N_14289);
nor UO_1117 (O_1117,N_14111,N_14398);
or UO_1118 (O_1118,N_14573,N_14031);
and UO_1119 (O_1119,N_14676,N_14903);
or UO_1120 (O_1120,N_14060,N_14246);
xnor UO_1121 (O_1121,N_14843,N_14847);
nor UO_1122 (O_1122,N_14169,N_14125);
nand UO_1123 (O_1123,N_14593,N_14194);
xnor UO_1124 (O_1124,N_14246,N_14956);
nor UO_1125 (O_1125,N_14512,N_14489);
xor UO_1126 (O_1126,N_14927,N_14445);
nor UO_1127 (O_1127,N_14783,N_14730);
or UO_1128 (O_1128,N_14130,N_14619);
nor UO_1129 (O_1129,N_14472,N_14191);
and UO_1130 (O_1130,N_14677,N_14238);
xor UO_1131 (O_1131,N_14556,N_14612);
nor UO_1132 (O_1132,N_14255,N_14190);
nor UO_1133 (O_1133,N_14202,N_14475);
nor UO_1134 (O_1134,N_14680,N_14907);
nor UO_1135 (O_1135,N_14968,N_14751);
and UO_1136 (O_1136,N_14417,N_14508);
or UO_1137 (O_1137,N_14895,N_14603);
xor UO_1138 (O_1138,N_14365,N_14183);
nor UO_1139 (O_1139,N_14689,N_14353);
and UO_1140 (O_1140,N_14946,N_14083);
xor UO_1141 (O_1141,N_14960,N_14758);
nor UO_1142 (O_1142,N_14029,N_14683);
and UO_1143 (O_1143,N_14428,N_14940);
or UO_1144 (O_1144,N_14651,N_14310);
xor UO_1145 (O_1145,N_14351,N_14413);
or UO_1146 (O_1146,N_14524,N_14324);
or UO_1147 (O_1147,N_14482,N_14591);
nor UO_1148 (O_1148,N_14339,N_14419);
or UO_1149 (O_1149,N_14573,N_14920);
nand UO_1150 (O_1150,N_14822,N_14833);
nor UO_1151 (O_1151,N_14616,N_14417);
or UO_1152 (O_1152,N_14130,N_14496);
and UO_1153 (O_1153,N_14406,N_14660);
nand UO_1154 (O_1154,N_14173,N_14571);
nand UO_1155 (O_1155,N_14571,N_14001);
and UO_1156 (O_1156,N_14978,N_14875);
or UO_1157 (O_1157,N_14161,N_14498);
xnor UO_1158 (O_1158,N_14410,N_14910);
nand UO_1159 (O_1159,N_14141,N_14314);
nor UO_1160 (O_1160,N_14654,N_14401);
or UO_1161 (O_1161,N_14440,N_14237);
xor UO_1162 (O_1162,N_14184,N_14093);
xor UO_1163 (O_1163,N_14870,N_14347);
and UO_1164 (O_1164,N_14217,N_14565);
and UO_1165 (O_1165,N_14314,N_14870);
nand UO_1166 (O_1166,N_14237,N_14616);
and UO_1167 (O_1167,N_14591,N_14254);
and UO_1168 (O_1168,N_14902,N_14722);
or UO_1169 (O_1169,N_14342,N_14836);
nor UO_1170 (O_1170,N_14881,N_14005);
xor UO_1171 (O_1171,N_14963,N_14307);
or UO_1172 (O_1172,N_14181,N_14606);
and UO_1173 (O_1173,N_14881,N_14454);
nand UO_1174 (O_1174,N_14802,N_14189);
xor UO_1175 (O_1175,N_14791,N_14619);
xnor UO_1176 (O_1176,N_14410,N_14847);
nor UO_1177 (O_1177,N_14693,N_14724);
xor UO_1178 (O_1178,N_14324,N_14778);
or UO_1179 (O_1179,N_14527,N_14874);
nor UO_1180 (O_1180,N_14189,N_14938);
or UO_1181 (O_1181,N_14113,N_14691);
nor UO_1182 (O_1182,N_14236,N_14053);
xnor UO_1183 (O_1183,N_14722,N_14380);
nor UO_1184 (O_1184,N_14488,N_14249);
or UO_1185 (O_1185,N_14768,N_14016);
and UO_1186 (O_1186,N_14128,N_14883);
nor UO_1187 (O_1187,N_14244,N_14709);
nand UO_1188 (O_1188,N_14937,N_14025);
or UO_1189 (O_1189,N_14680,N_14230);
or UO_1190 (O_1190,N_14386,N_14425);
or UO_1191 (O_1191,N_14726,N_14092);
nand UO_1192 (O_1192,N_14216,N_14991);
and UO_1193 (O_1193,N_14366,N_14035);
xor UO_1194 (O_1194,N_14146,N_14861);
or UO_1195 (O_1195,N_14028,N_14678);
or UO_1196 (O_1196,N_14409,N_14030);
or UO_1197 (O_1197,N_14609,N_14934);
nor UO_1198 (O_1198,N_14464,N_14566);
xnor UO_1199 (O_1199,N_14387,N_14257);
nor UO_1200 (O_1200,N_14378,N_14856);
nand UO_1201 (O_1201,N_14997,N_14614);
or UO_1202 (O_1202,N_14133,N_14930);
or UO_1203 (O_1203,N_14593,N_14638);
nand UO_1204 (O_1204,N_14041,N_14308);
and UO_1205 (O_1205,N_14563,N_14526);
and UO_1206 (O_1206,N_14338,N_14822);
nor UO_1207 (O_1207,N_14541,N_14945);
nand UO_1208 (O_1208,N_14864,N_14306);
nand UO_1209 (O_1209,N_14314,N_14712);
and UO_1210 (O_1210,N_14587,N_14815);
and UO_1211 (O_1211,N_14886,N_14115);
and UO_1212 (O_1212,N_14151,N_14512);
or UO_1213 (O_1213,N_14538,N_14678);
nand UO_1214 (O_1214,N_14215,N_14242);
nor UO_1215 (O_1215,N_14999,N_14406);
or UO_1216 (O_1216,N_14046,N_14321);
or UO_1217 (O_1217,N_14805,N_14686);
nand UO_1218 (O_1218,N_14114,N_14079);
xnor UO_1219 (O_1219,N_14897,N_14713);
xor UO_1220 (O_1220,N_14925,N_14696);
nor UO_1221 (O_1221,N_14901,N_14303);
xor UO_1222 (O_1222,N_14073,N_14949);
nand UO_1223 (O_1223,N_14997,N_14884);
nand UO_1224 (O_1224,N_14346,N_14178);
xor UO_1225 (O_1225,N_14609,N_14866);
nor UO_1226 (O_1226,N_14173,N_14523);
xor UO_1227 (O_1227,N_14441,N_14210);
nor UO_1228 (O_1228,N_14892,N_14422);
nor UO_1229 (O_1229,N_14460,N_14318);
nor UO_1230 (O_1230,N_14599,N_14985);
and UO_1231 (O_1231,N_14268,N_14746);
and UO_1232 (O_1232,N_14411,N_14673);
xor UO_1233 (O_1233,N_14595,N_14766);
and UO_1234 (O_1234,N_14212,N_14818);
nand UO_1235 (O_1235,N_14682,N_14128);
or UO_1236 (O_1236,N_14688,N_14506);
or UO_1237 (O_1237,N_14409,N_14336);
nand UO_1238 (O_1238,N_14805,N_14554);
xor UO_1239 (O_1239,N_14841,N_14114);
nand UO_1240 (O_1240,N_14983,N_14386);
nand UO_1241 (O_1241,N_14289,N_14384);
nor UO_1242 (O_1242,N_14676,N_14333);
or UO_1243 (O_1243,N_14256,N_14007);
and UO_1244 (O_1244,N_14853,N_14980);
and UO_1245 (O_1245,N_14136,N_14140);
xnor UO_1246 (O_1246,N_14220,N_14100);
and UO_1247 (O_1247,N_14859,N_14772);
nand UO_1248 (O_1248,N_14322,N_14657);
nor UO_1249 (O_1249,N_14718,N_14543);
xor UO_1250 (O_1250,N_14955,N_14058);
and UO_1251 (O_1251,N_14573,N_14700);
nand UO_1252 (O_1252,N_14651,N_14645);
xnor UO_1253 (O_1253,N_14658,N_14934);
nand UO_1254 (O_1254,N_14035,N_14589);
nor UO_1255 (O_1255,N_14015,N_14626);
nor UO_1256 (O_1256,N_14122,N_14314);
xor UO_1257 (O_1257,N_14062,N_14855);
nand UO_1258 (O_1258,N_14715,N_14997);
nand UO_1259 (O_1259,N_14308,N_14115);
and UO_1260 (O_1260,N_14899,N_14317);
and UO_1261 (O_1261,N_14337,N_14011);
and UO_1262 (O_1262,N_14137,N_14315);
or UO_1263 (O_1263,N_14430,N_14833);
or UO_1264 (O_1264,N_14122,N_14655);
or UO_1265 (O_1265,N_14552,N_14356);
xor UO_1266 (O_1266,N_14464,N_14980);
or UO_1267 (O_1267,N_14299,N_14162);
nand UO_1268 (O_1268,N_14316,N_14304);
xnor UO_1269 (O_1269,N_14983,N_14072);
nor UO_1270 (O_1270,N_14005,N_14529);
and UO_1271 (O_1271,N_14020,N_14536);
or UO_1272 (O_1272,N_14263,N_14825);
xnor UO_1273 (O_1273,N_14929,N_14600);
or UO_1274 (O_1274,N_14948,N_14985);
and UO_1275 (O_1275,N_14667,N_14003);
nor UO_1276 (O_1276,N_14697,N_14438);
nor UO_1277 (O_1277,N_14986,N_14474);
nand UO_1278 (O_1278,N_14110,N_14642);
nand UO_1279 (O_1279,N_14855,N_14220);
or UO_1280 (O_1280,N_14877,N_14890);
or UO_1281 (O_1281,N_14916,N_14740);
nand UO_1282 (O_1282,N_14655,N_14825);
xnor UO_1283 (O_1283,N_14606,N_14151);
xnor UO_1284 (O_1284,N_14375,N_14702);
or UO_1285 (O_1285,N_14468,N_14008);
and UO_1286 (O_1286,N_14059,N_14658);
xor UO_1287 (O_1287,N_14943,N_14617);
nor UO_1288 (O_1288,N_14335,N_14012);
and UO_1289 (O_1289,N_14531,N_14605);
or UO_1290 (O_1290,N_14238,N_14047);
and UO_1291 (O_1291,N_14404,N_14477);
xor UO_1292 (O_1292,N_14065,N_14344);
and UO_1293 (O_1293,N_14289,N_14370);
and UO_1294 (O_1294,N_14460,N_14281);
nor UO_1295 (O_1295,N_14959,N_14079);
nand UO_1296 (O_1296,N_14147,N_14727);
and UO_1297 (O_1297,N_14157,N_14517);
xnor UO_1298 (O_1298,N_14981,N_14326);
and UO_1299 (O_1299,N_14831,N_14737);
nor UO_1300 (O_1300,N_14289,N_14945);
nand UO_1301 (O_1301,N_14276,N_14817);
xor UO_1302 (O_1302,N_14419,N_14846);
or UO_1303 (O_1303,N_14179,N_14602);
xor UO_1304 (O_1304,N_14845,N_14163);
or UO_1305 (O_1305,N_14383,N_14283);
xnor UO_1306 (O_1306,N_14337,N_14794);
and UO_1307 (O_1307,N_14467,N_14372);
or UO_1308 (O_1308,N_14024,N_14604);
nor UO_1309 (O_1309,N_14044,N_14676);
xnor UO_1310 (O_1310,N_14025,N_14050);
nand UO_1311 (O_1311,N_14289,N_14853);
nor UO_1312 (O_1312,N_14569,N_14022);
and UO_1313 (O_1313,N_14420,N_14340);
or UO_1314 (O_1314,N_14410,N_14216);
and UO_1315 (O_1315,N_14172,N_14510);
and UO_1316 (O_1316,N_14290,N_14270);
and UO_1317 (O_1317,N_14384,N_14815);
xor UO_1318 (O_1318,N_14064,N_14293);
or UO_1319 (O_1319,N_14697,N_14888);
nor UO_1320 (O_1320,N_14352,N_14350);
nand UO_1321 (O_1321,N_14042,N_14669);
xnor UO_1322 (O_1322,N_14237,N_14634);
xnor UO_1323 (O_1323,N_14150,N_14056);
nand UO_1324 (O_1324,N_14056,N_14616);
and UO_1325 (O_1325,N_14930,N_14258);
and UO_1326 (O_1326,N_14243,N_14783);
or UO_1327 (O_1327,N_14823,N_14166);
xor UO_1328 (O_1328,N_14687,N_14657);
xnor UO_1329 (O_1329,N_14655,N_14927);
nor UO_1330 (O_1330,N_14113,N_14794);
xor UO_1331 (O_1331,N_14608,N_14909);
nand UO_1332 (O_1332,N_14557,N_14249);
and UO_1333 (O_1333,N_14813,N_14004);
xor UO_1334 (O_1334,N_14554,N_14009);
xor UO_1335 (O_1335,N_14167,N_14625);
or UO_1336 (O_1336,N_14261,N_14290);
xor UO_1337 (O_1337,N_14725,N_14572);
nand UO_1338 (O_1338,N_14231,N_14759);
and UO_1339 (O_1339,N_14062,N_14029);
xnor UO_1340 (O_1340,N_14439,N_14867);
xnor UO_1341 (O_1341,N_14370,N_14780);
nor UO_1342 (O_1342,N_14249,N_14498);
or UO_1343 (O_1343,N_14141,N_14892);
nand UO_1344 (O_1344,N_14089,N_14240);
or UO_1345 (O_1345,N_14510,N_14290);
and UO_1346 (O_1346,N_14001,N_14385);
and UO_1347 (O_1347,N_14478,N_14751);
nand UO_1348 (O_1348,N_14704,N_14055);
nand UO_1349 (O_1349,N_14763,N_14881);
xor UO_1350 (O_1350,N_14023,N_14059);
and UO_1351 (O_1351,N_14028,N_14710);
nand UO_1352 (O_1352,N_14837,N_14215);
or UO_1353 (O_1353,N_14083,N_14964);
nor UO_1354 (O_1354,N_14710,N_14790);
nand UO_1355 (O_1355,N_14835,N_14801);
xor UO_1356 (O_1356,N_14457,N_14717);
or UO_1357 (O_1357,N_14886,N_14784);
nand UO_1358 (O_1358,N_14246,N_14391);
or UO_1359 (O_1359,N_14799,N_14470);
nand UO_1360 (O_1360,N_14210,N_14092);
nand UO_1361 (O_1361,N_14679,N_14888);
and UO_1362 (O_1362,N_14986,N_14217);
nor UO_1363 (O_1363,N_14748,N_14728);
nand UO_1364 (O_1364,N_14801,N_14445);
or UO_1365 (O_1365,N_14193,N_14188);
or UO_1366 (O_1366,N_14082,N_14507);
nand UO_1367 (O_1367,N_14947,N_14056);
nor UO_1368 (O_1368,N_14227,N_14331);
nor UO_1369 (O_1369,N_14750,N_14943);
xor UO_1370 (O_1370,N_14844,N_14588);
or UO_1371 (O_1371,N_14672,N_14975);
or UO_1372 (O_1372,N_14863,N_14721);
nor UO_1373 (O_1373,N_14499,N_14318);
and UO_1374 (O_1374,N_14763,N_14159);
xor UO_1375 (O_1375,N_14353,N_14274);
nand UO_1376 (O_1376,N_14752,N_14116);
or UO_1377 (O_1377,N_14860,N_14638);
xnor UO_1378 (O_1378,N_14012,N_14734);
nor UO_1379 (O_1379,N_14965,N_14208);
nand UO_1380 (O_1380,N_14942,N_14432);
nand UO_1381 (O_1381,N_14991,N_14633);
and UO_1382 (O_1382,N_14863,N_14355);
and UO_1383 (O_1383,N_14711,N_14066);
or UO_1384 (O_1384,N_14483,N_14979);
nor UO_1385 (O_1385,N_14897,N_14795);
or UO_1386 (O_1386,N_14906,N_14956);
or UO_1387 (O_1387,N_14366,N_14854);
nand UO_1388 (O_1388,N_14571,N_14630);
and UO_1389 (O_1389,N_14407,N_14699);
nor UO_1390 (O_1390,N_14538,N_14312);
nor UO_1391 (O_1391,N_14360,N_14713);
nand UO_1392 (O_1392,N_14794,N_14086);
xor UO_1393 (O_1393,N_14813,N_14931);
nand UO_1394 (O_1394,N_14988,N_14598);
or UO_1395 (O_1395,N_14362,N_14101);
and UO_1396 (O_1396,N_14117,N_14219);
and UO_1397 (O_1397,N_14010,N_14389);
or UO_1398 (O_1398,N_14866,N_14427);
nand UO_1399 (O_1399,N_14163,N_14569);
nor UO_1400 (O_1400,N_14860,N_14296);
nand UO_1401 (O_1401,N_14390,N_14941);
xor UO_1402 (O_1402,N_14238,N_14708);
nor UO_1403 (O_1403,N_14289,N_14303);
xor UO_1404 (O_1404,N_14134,N_14777);
xor UO_1405 (O_1405,N_14486,N_14382);
xor UO_1406 (O_1406,N_14432,N_14768);
xnor UO_1407 (O_1407,N_14371,N_14735);
nor UO_1408 (O_1408,N_14097,N_14151);
or UO_1409 (O_1409,N_14962,N_14885);
or UO_1410 (O_1410,N_14389,N_14657);
nor UO_1411 (O_1411,N_14086,N_14758);
nand UO_1412 (O_1412,N_14777,N_14708);
nor UO_1413 (O_1413,N_14883,N_14314);
and UO_1414 (O_1414,N_14000,N_14855);
and UO_1415 (O_1415,N_14170,N_14744);
xnor UO_1416 (O_1416,N_14578,N_14831);
and UO_1417 (O_1417,N_14719,N_14064);
or UO_1418 (O_1418,N_14793,N_14671);
or UO_1419 (O_1419,N_14740,N_14836);
xor UO_1420 (O_1420,N_14800,N_14727);
or UO_1421 (O_1421,N_14718,N_14985);
nand UO_1422 (O_1422,N_14394,N_14235);
nand UO_1423 (O_1423,N_14125,N_14554);
and UO_1424 (O_1424,N_14800,N_14679);
nand UO_1425 (O_1425,N_14492,N_14262);
xnor UO_1426 (O_1426,N_14313,N_14896);
nand UO_1427 (O_1427,N_14181,N_14582);
or UO_1428 (O_1428,N_14886,N_14862);
nor UO_1429 (O_1429,N_14725,N_14660);
xor UO_1430 (O_1430,N_14879,N_14207);
or UO_1431 (O_1431,N_14780,N_14335);
or UO_1432 (O_1432,N_14826,N_14322);
and UO_1433 (O_1433,N_14782,N_14414);
or UO_1434 (O_1434,N_14890,N_14608);
xnor UO_1435 (O_1435,N_14601,N_14433);
or UO_1436 (O_1436,N_14335,N_14971);
nor UO_1437 (O_1437,N_14791,N_14166);
nor UO_1438 (O_1438,N_14423,N_14197);
nor UO_1439 (O_1439,N_14828,N_14134);
nand UO_1440 (O_1440,N_14901,N_14828);
xor UO_1441 (O_1441,N_14758,N_14765);
or UO_1442 (O_1442,N_14029,N_14954);
nor UO_1443 (O_1443,N_14536,N_14549);
nand UO_1444 (O_1444,N_14635,N_14411);
or UO_1445 (O_1445,N_14295,N_14101);
or UO_1446 (O_1446,N_14283,N_14494);
xor UO_1447 (O_1447,N_14244,N_14336);
nor UO_1448 (O_1448,N_14625,N_14901);
or UO_1449 (O_1449,N_14760,N_14286);
and UO_1450 (O_1450,N_14005,N_14755);
and UO_1451 (O_1451,N_14757,N_14249);
or UO_1452 (O_1452,N_14890,N_14493);
xor UO_1453 (O_1453,N_14906,N_14318);
or UO_1454 (O_1454,N_14506,N_14601);
and UO_1455 (O_1455,N_14721,N_14568);
and UO_1456 (O_1456,N_14013,N_14300);
xnor UO_1457 (O_1457,N_14091,N_14019);
xor UO_1458 (O_1458,N_14566,N_14218);
and UO_1459 (O_1459,N_14627,N_14457);
nor UO_1460 (O_1460,N_14887,N_14853);
and UO_1461 (O_1461,N_14332,N_14203);
nand UO_1462 (O_1462,N_14363,N_14719);
xnor UO_1463 (O_1463,N_14372,N_14802);
or UO_1464 (O_1464,N_14304,N_14314);
nand UO_1465 (O_1465,N_14616,N_14301);
or UO_1466 (O_1466,N_14498,N_14232);
xnor UO_1467 (O_1467,N_14675,N_14484);
xnor UO_1468 (O_1468,N_14274,N_14586);
and UO_1469 (O_1469,N_14051,N_14087);
or UO_1470 (O_1470,N_14641,N_14261);
and UO_1471 (O_1471,N_14074,N_14558);
nor UO_1472 (O_1472,N_14821,N_14515);
xor UO_1473 (O_1473,N_14464,N_14852);
nor UO_1474 (O_1474,N_14955,N_14038);
and UO_1475 (O_1475,N_14554,N_14613);
and UO_1476 (O_1476,N_14864,N_14683);
and UO_1477 (O_1477,N_14341,N_14661);
nand UO_1478 (O_1478,N_14610,N_14094);
xnor UO_1479 (O_1479,N_14486,N_14650);
xor UO_1480 (O_1480,N_14113,N_14221);
or UO_1481 (O_1481,N_14226,N_14705);
and UO_1482 (O_1482,N_14659,N_14125);
nor UO_1483 (O_1483,N_14516,N_14688);
nor UO_1484 (O_1484,N_14764,N_14724);
or UO_1485 (O_1485,N_14316,N_14659);
xnor UO_1486 (O_1486,N_14948,N_14895);
or UO_1487 (O_1487,N_14588,N_14458);
xor UO_1488 (O_1488,N_14282,N_14260);
nor UO_1489 (O_1489,N_14655,N_14308);
or UO_1490 (O_1490,N_14626,N_14296);
nor UO_1491 (O_1491,N_14124,N_14628);
xnor UO_1492 (O_1492,N_14922,N_14622);
xor UO_1493 (O_1493,N_14860,N_14375);
xor UO_1494 (O_1494,N_14158,N_14456);
nand UO_1495 (O_1495,N_14953,N_14722);
or UO_1496 (O_1496,N_14108,N_14004);
or UO_1497 (O_1497,N_14063,N_14315);
or UO_1498 (O_1498,N_14535,N_14934);
nand UO_1499 (O_1499,N_14070,N_14775);
nor UO_1500 (O_1500,N_14765,N_14920);
nand UO_1501 (O_1501,N_14893,N_14449);
xnor UO_1502 (O_1502,N_14374,N_14360);
nand UO_1503 (O_1503,N_14547,N_14809);
nand UO_1504 (O_1504,N_14383,N_14703);
xnor UO_1505 (O_1505,N_14632,N_14918);
or UO_1506 (O_1506,N_14965,N_14268);
or UO_1507 (O_1507,N_14009,N_14788);
xor UO_1508 (O_1508,N_14456,N_14446);
nand UO_1509 (O_1509,N_14881,N_14807);
nand UO_1510 (O_1510,N_14151,N_14084);
and UO_1511 (O_1511,N_14239,N_14358);
xnor UO_1512 (O_1512,N_14685,N_14238);
or UO_1513 (O_1513,N_14391,N_14552);
xnor UO_1514 (O_1514,N_14735,N_14004);
and UO_1515 (O_1515,N_14189,N_14817);
nor UO_1516 (O_1516,N_14653,N_14926);
nor UO_1517 (O_1517,N_14795,N_14829);
nand UO_1518 (O_1518,N_14195,N_14888);
nor UO_1519 (O_1519,N_14205,N_14504);
or UO_1520 (O_1520,N_14276,N_14980);
or UO_1521 (O_1521,N_14711,N_14757);
nand UO_1522 (O_1522,N_14572,N_14524);
nor UO_1523 (O_1523,N_14357,N_14235);
xor UO_1524 (O_1524,N_14037,N_14323);
nor UO_1525 (O_1525,N_14280,N_14207);
and UO_1526 (O_1526,N_14860,N_14531);
xor UO_1527 (O_1527,N_14117,N_14127);
and UO_1528 (O_1528,N_14352,N_14996);
nand UO_1529 (O_1529,N_14259,N_14703);
nor UO_1530 (O_1530,N_14143,N_14215);
xor UO_1531 (O_1531,N_14000,N_14013);
and UO_1532 (O_1532,N_14391,N_14036);
or UO_1533 (O_1533,N_14762,N_14003);
and UO_1534 (O_1534,N_14449,N_14909);
xor UO_1535 (O_1535,N_14344,N_14855);
xor UO_1536 (O_1536,N_14533,N_14688);
nand UO_1537 (O_1537,N_14044,N_14934);
nor UO_1538 (O_1538,N_14026,N_14049);
nor UO_1539 (O_1539,N_14908,N_14354);
or UO_1540 (O_1540,N_14544,N_14444);
nor UO_1541 (O_1541,N_14694,N_14644);
or UO_1542 (O_1542,N_14531,N_14501);
and UO_1543 (O_1543,N_14550,N_14812);
nor UO_1544 (O_1544,N_14928,N_14882);
or UO_1545 (O_1545,N_14110,N_14912);
xnor UO_1546 (O_1546,N_14566,N_14576);
nor UO_1547 (O_1547,N_14709,N_14142);
nand UO_1548 (O_1548,N_14167,N_14754);
nand UO_1549 (O_1549,N_14165,N_14086);
nand UO_1550 (O_1550,N_14012,N_14453);
xnor UO_1551 (O_1551,N_14370,N_14962);
and UO_1552 (O_1552,N_14246,N_14629);
xnor UO_1553 (O_1553,N_14059,N_14909);
or UO_1554 (O_1554,N_14666,N_14867);
and UO_1555 (O_1555,N_14555,N_14539);
nor UO_1556 (O_1556,N_14602,N_14974);
and UO_1557 (O_1557,N_14905,N_14820);
xnor UO_1558 (O_1558,N_14960,N_14333);
and UO_1559 (O_1559,N_14281,N_14720);
or UO_1560 (O_1560,N_14529,N_14361);
and UO_1561 (O_1561,N_14175,N_14123);
or UO_1562 (O_1562,N_14795,N_14482);
nor UO_1563 (O_1563,N_14929,N_14626);
xor UO_1564 (O_1564,N_14068,N_14873);
or UO_1565 (O_1565,N_14880,N_14172);
xor UO_1566 (O_1566,N_14579,N_14795);
and UO_1567 (O_1567,N_14333,N_14767);
or UO_1568 (O_1568,N_14686,N_14285);
xnor UO_1569 (O_1569,N_14118,N_14880);
xor UO_1570 (O_1570,N_14235,N_14890);
nor UO_1571 (O_1571,N_14784,N_14241);
nor UO_1572 (O_1572,N_14254,N_14854);
xnor UO_1573 (O_1573,N_14494,N_14427);
xor UO_1574 (O_1574,N_14208,N_14398);
nand UO_1575 (O_1575,N_14634,N_14575);
nand UO_1576 (O_1576,N_14616,N_14150);
or UO_1577 (O_1577,N_14117,N_14803);
nand UO_1578 (O_1578,N_14726,N_14158);
and UO_1579 (O_1579,N_14745,N_14574);
xnor UO_1580 (O_1580,N_14063,N_14731);
and UO_1581 (O_1581,N_14246,N_14679);
xor UO_1582 (O_1582,N_14778,N_14869);
nand UO_1583 (O_1583,N_14624,N_14450);
xnor UO_1584 (O_1584,N_14614,N_14825);
or UO_1585 (O_1585,N_14693,N_14864);
xnor UO_1586 (O_1586,N_14398,N_14716);
xnor UO_1587 (O_1587,N_14993,N_14369);
nor UO_1588 (O_1588,N_14854,N_14278);
and UO_1589 (O_1589,N_14164,N_14178);
nor UO_1590 (O_1590,N_14555,N_14092);
and UO_1591 (O_1591,N_14932,N_14074);
nand UO_1592 (O_1592,N_14372,N_14100);
nor UO_1593 (O_1593,N_14860,N_14544);
nor UO_1594 (O_1594,N_14316,N_14148);
or UO_1595 (O_1595,N_14681,N_14452);
nand UO_1596 (O_1596,N_14013,N_14655);
or UO_1597 (O_1597,N_14482,N_14103);
xor UO_1598 (O_1598,N_14227,N_14365);
nor UO_1599 (O_1599,N_14304,N_14923);
xnor UO_1600 (O_1600,N_14436,N_14640);
nand UO_1601 (O_1601,N_14513,N_14641);
or UO_1602 (O_1602,N_14838,N_14182);
nor UO_1603 (O_1603,N_14290,N_14560);
nand UO_1604 (O_1604,N_14718,N_14428);
nor UO_1605 (O_1605,N_14170,N_14950);
and UO_1606 (O_1606,N_14078,N_14513);
xor UO_1607 (O_1607,N_14759,N_14564);
xor UO_1608 (O_1608,N_14202,N_14737);
or UO_1609 (O_1609,N_14276,N_14925);
xnor UO_1610 (O_1610,N_14970,N_14320);
nand UO_1611 (O_1611,N_14463,N_14526);
nor UO_1612 (O_1612,N_14998,N_14988);
nand UO_1613 (O_1613,N_14425,N_14085);
nand UO_1614 (O_1614,N_14590,N_14139);
or UO_1615 (O_1615,N_14579,N_14130);
and UO_1616 (O_1616,N_14947,N_14789);
nor UO_1617 (O_1617,N_14683,N_14465);
nand UO_1618 (O_1618,N_14010,N_14447);
and UO_1619 (O_1619,N_14228,N_14297);
nor UO_1620 (O_1620,N_14327,N_14371);
or UO_1621 (O_1621,N_14414,N_14324);
or UO_1622 (O_1622,N_14415,N_14853);
xor UO_1623 (O_1623,N_14175,N_14359);
and UO_1624 (O_1624,N_14502,N_14057);
or UO_1625 (O_1625,N_14988,N_14311);
or UO_1626 (O_1626,N_14929,N_14991);
or UO_1627 (O_1627,N_14193,N_14853);
xor UO_1628 (O_1628,N_14171,N_14507);
xor UO_1629 (O_1629,N_14948,N_14572);
and UO_1630 (O_1630,N_14906,N_14765);
or UO_1631 (O_1631,N_14963,N_14647);
nand UO_1632 (O_1632,N_14788,N_14423);
nand UO_1633 (O_1633,N_14824,N_14754);
xor UO_1634 (O_1634,N_14732,N_14876);
or UO_1635 (O_1635,N_14441,N_14965);
nand UO_1636 (O_1636,N_14356,N_14453);
xnor UO_1637 (O_1637,N_14462,N_14114);
nor UO_1638 (O_1638,N_14397,N_14027);
xnor UO_1639 (O_1639,N_14451,N_14890);
nand UO_1640 (O_1640,N_14367,N_14210);
and UO_1641 (O_1641,N_14734,N_14244);
nor UO_1642 (O_1642,N_14061,N_14954);
nand UO_1643 (O_1643,N_14095,N_14870);
and UO_1644 (O_1644,N_14766,N_14137);
nor UO_1645 (O_1645,N_14685,N_14527);
and UO_1646 (O_1646,N_14434,N_14176);
nor UO_1647 (O_1647,N_14655,N_14445);
nor UO_1648 (O_1648,N_14440,N_14486);
nand UO_1649 (O_1649,N_14231,N_14184);
nor UO_1650 (O_1650,N_14446,N_14828);
xnor UO_1651 (O_1651,N_14364,N_14631);
nand UO_1652 (O_1652,N_14821,N_14597);
and UO_1653 (O_1653,N_14248,N_14675);
nor UO_1654 (O_1654,N_14504,N_14372);
nor UO_1655 (O_1655,N_14840,N_14758);
xor UO_1656 (O_1656,N_14753,N_14710);
or UO_1657 (O_1657,N_14327,N_14722);
or UO_1658 (O_1658,N_14217,N_14601);
or UO_1659 (O_1659,N_14563,N_14119);
nor UO_1660 (O_1660,N_14327,N_14869);
nand UO_1661 (O_1661,N_14220,N_14364);
nand UO_1662 (O_1662,N_14625,N_14862);
nand UO_1663 (O_1663,N_14566,N_14323);
nand UO_1664 (O_1664,N_14750,N_14744);
xnor UO_1665 (O_1665,N_14227,N_14896);
nand UO_1666 (O_1666,N_14036,N_14871);
nand UO_1667 (O_1667,N_14670,N_14139);
nor UO_1668 (O_1668,N_14070,N_14599);
xor UO_1669 (O_1669,N_14023,N_14173);
xor UO_1670 (O_1670,N_14406,N_14611);
or UO_1671 (O_1671,N_14398,N_14460);
nor UO_1672 (O_1672,N_14851,N_14975);
nand UO_1673 (O_1673,N_14021,N_14829);
xor UO_1674 (O_1674,N_14286,N_14296);
nor UO_1675 (O_1675,N_14101,N_14973);
and UO_1676 (O_1676,N_14130,N_14976);
nor UO_1677 (O_1677,N_14420,N_14522);
nand UO_1678 (O_1678,N_14005,N_14651);
xor UO_1679 (O_1679,N_14277,N_14983);
or UO_1680 (O_1680,N_14185,N_14070);
xor UO_1681 (O_1681,N_14156,N_14455);
and UO_1682 (O_1682,N_14952,N_14700);
xor UO_1683 (O_1683,N_14057,N_14266);
or UO_1684 (O_1684,N_14658,N_14001);
nand UO_1685 (O_1685,N_14429,N_14006);
nand UO_1686 (O_1686,N_14146,N_14976);
nand UO_1687 (O_1687,N_14881,N_14898);
xnor UO_1688 (O_1688,N_14387,N_14720);
and UO_1689 (O_1689,N_14259,N_14485);
or UO_1690 (O_1690,N_14059,N_14262);
nand UO_1691 (O_1691,N_14642,N_14011);
or UO_1692 (O_1692,N_14322,N_14559);
xor UO_1693 (O_1693,N_14709,N_14770);
xor UO_1694 (O_1694,N_14970,N_14117);
or UO_1695 (O_1695,N_14675,N_14258);
and UO_1696 (O_1696,N_14759,N_14063);
and UO_1697 (O_1697,N_14273,N_14203);
nand UO_1698 (O_1698,N_14476,N_14833);
xor UO_1699 (O_1699,N_14258,N_14827);
and UO_1700 (O_1700,N_14137,N_14325);
xnor UO_1701 (O_1701,N_14047,N_14221);
xnor UO_1702 (O_1702,N_14097,N_14547);
nand UO_1703 (O_1703,N_14248,N_14642);
xnor UO_1704 (O_1704,N_14618,N_14206);
xor UO_1705 (O_1705,N_14830,N_14312);
or UO_1706 (O_1706,N_14851,N_14546);
or UO_1707 (O_1707,N_14656,N_14832);
nor UO_1708 (O_1708,N_14810,N_14279);
and UO_1709 (O_1709,N_14851,N_14280);
xor UO_1710 (O_1710,N_14829,N_14810);
and UO_1711 (O_1711,N_14138,N_14488);
or UO_1712 (O_1712,N_14829,N_14731);
xnor UO_1713 (O_1713,N_14781,N_14601);
nor UO_1714 (O_1714,N_14427,N_14219);
nor UO_1715 (O_1715,N_14018,N_14702);
nand UO_1716 (O_1716,N_14627,N_14218);
and UO_1717 (O_1717,N_14965,N_14047);
and UO_1718 (O_1718,N_14757,N_14565);
and UO_1719 (O_1719,N_14773,N_14061);
xnor UO_1720 (O_1720,N_14219,N_14913);
nor UO_1721 (O_1721,N_14672,N_14899);
and UO_1722 (O_1722,N_14297,N_14254);
nand UO_1723 (O_1723,N_14341,N_14243);
xnor UO_1724 (O_1724,N_14285,N_14629);
nor UO_1725 (O_1725,N_14060,N_14873);
or UO_1726 (O_1726,N_14619,N_14885);
and UO_1727 (O_1727,N_14946,N_14626);
or UO_1728 (O_1728,N_14778,N_14724);
nand UO_1729 (O_1729,N_14142,N_14075);
nand UO_1730 (O_1730,N_14639,N_14098);
xnor UO_1731 (O_1731,N_14115,N_14289);
nor UO_1732 (O_1732,N_14250,N_14699);
nand UO_1733 (O_1733,N_14123,N_14774);
xor UO_1734 (O_1734,N_14527,N_14808);
or UO_1735 (O_1735,N_14803,N_14960);
and UO_1736 (O_1736,N_14504,N_14080);
nor UO_1737 (O_1737,N_14319,N_14101);
or UO_1738 (O_1738,N_14972,N_14165);
nand UO_1739 (O_1739,N_14923,N_14840);
or UO_1740 (O_1740,N_14773,N_14025);
xnor UO_1741 (O_1741,N_14762,N_14482);
xnor UO_1742 (O_1742,N_14066,N_14898);
nor UO_1743 (O_1743,N_14981,N_14952);
and UO_1744 (O_1744,N_14776,N_14546);
or UO_1745 (O_1745,N_14773,N_14858);
xnor UO_1746 (O_1746,N_14085,N_14898);
nor UO_1747 (O_1747,N_14120,N_14341);
or UO_1748 (O_1748,N_14196,N_14426);
nor UO_1749 (O_1749,N_14082,N_14982);
xor UO_1750 (O_1750,N_14045,N_14367);
nand UO_1751 (O_1751,N_14840,N_14233);
nor UO_1752 (O_1752,N_14085,N_14809);
xnor UO_1753 (O_1753,N_14609,N_14924);
nand UO_1754 (O_1754,N_14878,N_14087);
nand UO_1755 (O_1755,N_14625,N_14308);
or UO_1756 (O_1756,N_14589,N_14185);
nor UO_1757 (O_1757,N_14037,N_14373);
and UO_1758 (O_1758,N_14699,N_14386);
nand UO_1759 (O_1759,N_14917,N_14279);
xor UO_1760 (O_1760,N_14358,N_14058);
xor UO_1761 (O_1761,N_14686,N_14036);
xor UO_1762 (O_1762,N_14547,N_14935);
nor UO_1763 (O_1763,N_14504,N_14017);
xnor UO_1764 (O_1764,N_14259,N_14179);
nor UO_1765 (O_1765,N_14840,N_14130);
nor UO_1766 (O_1766,N_14434,N_14108);
nor UO_1767 (O_1767,N_14567,N_14337);
and UO_1768 (O_1768,N_14851,N_14838);
nor UO_1769 (O_1769,N_14589,N_14934);
nor UO_1770 (O_1770,N_14697,N_14957);
or UO_1771 (O_1771,N_14302,N_14632);
xor UO_1772 (O_1772,N_14980,N_14027);
xor UO_1773 (O_1773,N_14127,N_14818);
and UO_1774 (O_1774,N_14332,N_14375);
and UO_1775 (O_1775,N_14679,N_14319);
and UO_1776 (O_1776,N_14396,N_14041);
and UO_1777 (O_1777,N_14843,N_14420);
nand UO_1778 (O_1778,N_14009,N_14901);
and UO_1779 (O_1779,N_14530,N_14706);
or UO_1780 (O_1780,N_14026,N_14771);
nor UO_1781 (O_1781,N_14808,N_14101);
nand UO_1782 (O_1782,N_14770,N_14719);
nor UO_1783 (O_1783,N_14351,N_14971);
or UO_1784 (O_1784,N_14029,N_14413);
nor UO_1785 (O_1785,N_14169,N_14062);
nor UO_1786 (O_1786,N_14922,N_14439);
xnor UO_1787 (O_1787,N_14734,N_14040);
or UO_1788 (O_1788,N_14156,N_14068);
or UO_1789 (O_1789,N_14856,N_14875);
xnor UO_1790 (O_1790,N_14662,N_14675);
xnor UO_1791 (O_1791,N_14575,N_14196);
and UO_1792 (O_1792,N_14438,N_14830);
or UO_1793 (O_1793,N_14081,N_14586);
or UO_1794 (O_1794,N_14880,N_14081);
and UO_1795 (O_1795,N_14196,N_14415);
xnor UO_1796 (O_1796,N_14443,N_14406);
xnor UO_1797 (O_1797,N_14263,N_14607);
or UO_1798 (O_1798,N_14701,N_14709);
nand UO_1799 (O_1799,N_14829,N_14484);
and UO_1800 (O_1800,N_14488,N_14990);
xnor UO_1801 (O_1801,N_14857,N_14104);
nand UO_1802 (O_1802,N_14725,N_14542);
or UO_1803 (O_1803,N_14053,N_14123);
xor UO_1804 (O_1804,N_14092,N_14362);
xor UO_1805 (O_1805,N_14322,N_14150);
and UO_1806 (O_1806,N_14158,N_14735);
nand UO_1807 (O_1807,N_14078,N_14224);
nand UO_1808 (O_1808,N_14197,N_14754);
nor UO_1809 (O_1809,N_14538,N_14700);
xor UO_1810 (O_1810,N_14205,N_14483);
or UO_1811 (O_1811,N_14022,N_14037);
nor UO_1812 (O_1812,N_14310,N_14605);
and UO_1813 (O_1813,N_14339,N_14808);
or UO_1814 (O_1814,N_14801,N_14844);
nor UO_1815 (O_1815,N_14811,N_14814);
xnor UO_1816 (O_1816,N_14535,N_14557);
xnor UO_1817 (O_1817,N_14471,N_14875);
or UO_1818 (O_1818,N_14536,N_14709);
nor UO_1819 (O_1819,N_14870,N_14490);
or UO_1820 (O_1820,N_14162,N_14902);
nor UO_1821 (O_1821,N_14947,N_14503);
xnor UO_1822 (O_1822,N_14970,N_14704);
xor UO_1823 (O_1823,N_14679,N_14555);
nor UO_1824 (O_1824,N_14443,N_14919);
and UO_1825 (O_1825,N_14459,N_14928);
nand UO_1826 (O_1826,N_14484,N_14404);
and UO_1827 (O_1827,N_14786,N_14901);
nor UO_1828 (O_1828,N_14412,N_14979);
xor UO_1829 (O_1829,N_14196,N_14111);
and UO_1830 (O_1830,N_14785,N_14846);
or UO_1831 (O_1831,N_14691,N_14920);
nand UO_1832 (O_1832,N_14317,N_14595);
nor UO_1833 (O_1833,N_14315,N_14079);
xor UO_1834 (O_1834,N_14614,N_14731);
xor UO_1835 (O_1835,N_14769,N_14330);
xor UO_1836 (O_1836,N_14203,N_14571);
xnor UO_1837 (O_1837,N_14426,N_14537);
xnor UO_1838 (O_1838,N_14322,N_14988);
and UO_1839 (O_1839,N_14837,N_14051);
nor UO_1840 (O_1840,N_14343,N_14441);
nand UO_1841 (O_1841,N_14735,N_14642);
and UO_1842 (O_1842,N_14467,N_14576);
and UO_1843 (O_1843,N_14067,N_14572);
nor UO_1844 (O_1844,N_14574,N_14832);
and UO_1845 (O_1845,N_14321,N_14097);
and UO_1846 (O_1846,N_14597,N_14477);
or UO_1847 (O_1847,N_14038,N_14332);
and UO_1848 (O_1848,N_14178,N_14628);
or UO_1849 (O_1849,N_14585,N_14085);
nand UO_1850 (O_1850,N_14052,N_14513);
or UO_1851 (O_1851,N_14445,N_14929);
and UO_1852 (O_1852,N_14838,N_14285);
nand UO_1853 (O_1853,N_14770,N_14375);
or UO_1854 (O_1854,N_14739,N_14113);
and UO_1855 (O_1855,N_14304,N_14176);
nor UO_1856 (O_1856,N_14103,N_14707);
and UO_1857 (O_1857,N_14059,N_14416);
nor UO_1858 (O_1858,N_14193,N_14631);
nor UO_1859 (O_1859,N_14828,N_14816);
nor UO_1860 (O_1860,N_14579,N_14321);
nand UO_1861 (O_1861,N_14441,N_14236);
and UO_1862 (O_1862,N_14379,N_14721);
and UO_1863 (O_1863,N_14385,N_14750);
nor UO_1864 (O_1864,N_14225,N_14804);
xnor UO_1865 (O_1865,N_14946,N_14328);
and UO_1866 (O_1866,N_14967,N_14775);
nand UO_1867 (O_1867,N_14449,N_14690);
nand UO_1868 (O_1868,N_14607,N_14215);
nor UO_1869 (O_1869,N_14508,N_14513);
nor UO_1870 (O_1870,N_14290,N_14919);
xnor UO_1871 (O_1871,N_14988,N_14605);
and UO_1872 (O_1872,N_14182,N_14096);
nand UO_1873 (O_1873,N_14037,N_14027);
nor UO_1874 (O_1874,N_14302,N_14349);
nor UO_1875 (O_1875,N_14828,N_14710);
or UO_1876 (O_1876,N_14009,N_14306);
and UO_1877 (O_1877,N_14290,N_14314);
or UO_1878 (O_1878,N_14007,N_14017);
or UO_1879 (O_1879,N_14154,N_14103);
and UO_1880 (O_1880,N_14292,N_14852);
or UO_1881 (O_1881,N_14839,N_14051);
or UO_1882 (O_1882,N_14484,N_14039);
nor UO_1883 (O_1883,N_14457,N_14516);
nand UO_1884 (O_1884,N_14210,N_14507);
xor UO_1885 (O_1885,N_14623,N_14511);
and UO_1886 (O_1886,N_14000,N_14436);
xnor UO_1887 (O_1887,N_14403,N_14048);
nand UO_1888 (O_1888,N_14101,N_14443);
or UO_1889 (O_1889,N_14650,N_14231);
xor UO_1890 (O_1890,N_14827,N_14473);
nor UO_1891 (O_1891,N_14479,N_14136);
and UO_1892 (O_1892,N_14021,N_14120);
xor UO_1893 (O_1893,N_14641,N_14222);
and UO_1894 (O_1894,N_14393,N_14577);
xor UO_1895 (O_1895,N_14091,N_14963);
and UO_1896 (O_1896,N_14286,N_14368);
nor UO_1897 (O_1897,N_14265,N_14355);
nand UO_1898 (O_1898,N_14811,N_14177);
xnor UO_1899 (O_1899,N_14513,N_14428);
or UO_1900 (O_1900,N_14289,N_14097);
nor UO_1901 (O_1901,N_14081,N_14236);
nand UO_1902 (O_1902,N_14563,N_14903);
or UO_1903 (O_1903,N_14803,N_14192);
or UO_1904 (O_1904,N_14826,N_14704);
and UO_1905 (O_1905,N_14276,N_14708);
or UO_1906 (O_1906,N_14432,N_14129);
nand UO_1907 (O_1907,N_14547,N_14756);
nand UO_1908 (O_1908,N_14105,N_14702);
nor UO_1909 (O_1909,N_14530,N_14796);
nor UO_1910 (O_1910,N_14217,N_14895);
and UO_1911 (O_1911,N_14810,N_14508);
xor UO_1912 (O_1912,N_14311,N_14059);
or UO_1913 (O_1913,N_14814,N_14168);
xnor UO_1914 (O_1914,N_14042,N_14239);
xnor UO_1915 (O_1915,N_14899,N_14485);
nand UO_1916 (O_1916,N_14925,N_14108);
and UO_1917 (O_1917,N_14994,N_14968);
nor UO_1918 (O_1918,N_14807,N_14350);
and UO_1919 (O_1919,N_14067,N_14262);
nor UO_1920 (O_1920,N_14810,N_14696);
or UO_1921 (O_1921,N_14704,N_14266);
xnor UO_1922 (O_1922,N_14095,N_14763);
nor UO_1923 (O_1923,N_14156,N_14872);
xor UO_1924 (O_1924,N_14073,N_14543);
nor UO_1925 (O_1925,N_14169,N_14747);
xnor UO_1926 (O_1926,N_14631,N_14303);
xnor UO_1927 (O_1927,N_14549,N_14878);
and UO_1928 (O_1928,N_14905,N_14817);
xnor UO_1929 (O_1929,N_14274,N_14014);
nand UO_1930 (O_1930,N_14915,N_14851);
or UO_1931 (O_1931,N_14250,N_14948);
nand UO_1932 (O_1932,N_14987,N_14306);
xnor UO_1933 (O_1933,N_14297,N_14893);
and UO_1934 (O_1934,N_14205,N_14890);
and UO_1935 (O_1935,N_14800,N_14873);
or UO_1936 (O_1936,N_14570,N_14708);
and UO_1937 (O_1937,N_14248,N_14874);
nand UO_1938 (O_1938,N_14968,N_14550);
nor UO_1939 (O_1939,N_14136,N_14574);
and UO_1940 (O_1940,N_14708,N_14127);
and UO_1941 (O_1941,N_14261,N_14191);
xnor UO_1942 (O_1942,N_14272,N_14177);
nor UO_1943 (O_1943,N_14458,N_14028);
nor UO_1944 (O_1944,N_14195,N_14524);
or UO_1945 (O_1945,N_14218,N_14110);
xnor UO_1946 (O_1946,N_14603,N_14683);
or UO_1947 (O_1947,N_14418,N_14354);
and UO_1948 (O_1948,N_14937,N_14446);
nand UO_1949 (O_1949,N_14646,N_14080);
nand UO_1950 (O_1950,N_14046,N_14846);
nand UO_1951 (O_1951,N_14823,N_14132);
nand UO_1952 (O_1952,N_14254,N_14787);
nor UO_1953 (O_1953,N_14713,N_14794);
or UO_1954 (O_1954,N_14701,N_14775);
xnor UO_1955 (O_1955,N_14819,N_14924);
and UO_1956 (O_1956,N_14164,N_14793);
or UO_1957 (O_1957,N_14903,N_14014);
and UO_1958 (O_1958,N_14780,N_14518);
and UO_1959 (O_1959,N_14942,N_14033);
nand UO_1960 (O_1960,N_14252,N_14093);
xnor UO_1961 (O_1961,N_14637,N_14784);
nor UO_1962 (O_1962,N_14041,N_14879);
nand UO_1963 (O_1963,N_14148,N_14202);
nand UO_1964 (O_1964,N_14698,N_14904);
xor UO_1965 (O_1965,N_14047,N_14656);
and UO_1966 (O_1966,N_14333,N_14487);
nand UO_1967 (O_1967,N_14993,N_14199);
nand UO_1968 (O_1968,N_14944,N_14961);
and UO_1969 (O_1969,N_14016,N_14892);
xnor UO_1970 (O_1970,N_14971,N_14887);
nor UO_1971 (O_1971,N_14510,N_14431);
nor UO_1972 (O_1972,N_14729,N_14797);
nand UO_1973 (O_1973,N_14470,N_14179);
xor UO_1974 (O_1974,N_14078,N_14047);
and UO_1975 (O_1975,N_14729,N_14284);
nor UO_1976 (O_1976,N_14601,N_14365);
or UO_1977 (O_1977,N_14016,N_14566);
and UO_1978 (O_1978,N_14803,N_14641);
and UO_1979 (O_1979,N_14662,N_14873);
and UO_1980 (O_1980,N_14179,N_14795);
nor UO_1981 (O_1981,N_14455,N_14709);
xnor UO_1982 (O_1982,N_14898,N_14680);
and UO_1983 (O_1983,N_14634,N_14178);
xnor UO_1984 (O_1984,N_14856,N_14058);
nand UO_1985 (O_1985,N_14824,N_14382);
xnor UO_1986 (O_1986,N_14367,N_14930);
nand UO_1987 (O_1987,N_14015,N_14376);
and UO_1988 (O_1988,N_14885,N_14821);
nand UO_1989 (O_1989,N_14185,N_14804);
and UO_1990 (O_1990,N_14185,N_14869);
nand UO_1991 (O_1991,N_14508,N_14264);
and UO_1992 (O_1992,N_14982,N_14604);
nand UO_1993 (O_1993,N_14943,N_14442);
or UO_1994 (O_1994,N_14290,N_14150);
or UO_1995 (O_1995,N_14766,N_14269);
or UO_1996 (O_1996,N_14566,N_14012);
xnor UO_1997 (O_1997,N_14058,N_14635);
xor UO_1998 (O_1998,N_14908,N_14319);
xor UO_1999 (O_1999,N_14384,N_14240);
endmodule