module basic_1500_15000_2000_20_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
or U0 (N_0,In_627,In_1239);
xor U1 (N_1,In_314,In_769);
nand U2 (N_2,In_849,In_1093);
nand U3 (N_3,In_1253,In_923);
nand U4 (N_4,In_817,In_1418);
and U5 (N_5,In_1163,In_1073);
nand U6 (N_6,In_1077,In_1096);
nand U7 (N_7,In_1429,In_10);
xor U8 (N_8,In_774,In_130);
nand U9 (N_9,In_1472,In_789);
or U10 (N_10,In_641,In_688);
and U11 (N_11,In_625,In_982);
xnor U12 (N_12,In_327,In_341);
nand U13 (N_13,In_374,In_1101);
nor U14 (N_14,In_349,In_494);
and U15 (N_15,In_1082,In_167);
nor U16 (N_16,In_368,In_850);
xor U17 (N_17,In_1285,In_1311);
xor U18 (N_18,In_123,In_1030);
nor U19 (N_19,In_164,In_809);
nand U20 (N_20,In_237,In_1259);
and U21 (N_21,In_903,In_1432);
xnor U22 (N_22,In_560,In_978);
nand U23 (N_23,In_82,In_686);
xor U24 (N_24,In_1074,In_615);
nand U25 (N_25,In_800,In_1105);
xnor U26 (N_26,In_1111,In_523);
nand U27 (N_27,In_929,In_1463);
or U28 (N_28,In_997,In_1498);
nor U29 (N_29,In_537,In_1245);
or U30 (N_30,In_525,In_369);
nand U31 (N_31,In_410,In_1002);
or U32 (N_32,In_1161,In_70);
and U33 (N_33,In_1068,In_587);
or U34 (N_34,In_1388,In_415);
xor U35 (N_35,In_1294,In_1181);
nor U36 (N_36,In_440,In_475);
and U37 (N_37,In_348,In_746);
nor U38 (N_38,In_1042,In_1116);
nand U39 (N_39,In_512,In_947);
nor U40 (N_40,In_313,In_701);
and U41 (N_41,In_553,In_78);
nand U42 (N_42,In_1070,In_631);
or U43 (N_43,In_976,In_943);
nor U44 (N_44,In_1410,In_222);
nand U45 (N_45,In_1075,In_502);
xnor U46 (N_46,In_1129,In_71);
or U47 (N_47,In_1492,In_216);
and U48 (N_48,In_75,In_205);
or U49 (N_49,In_1089,In_1480);
and U50 (N_50,In_672,In_1489);
nand U51 (N_51,In_268,In_687);
nand U52 (N_52,In_810,In_964);
or U53 (N_53,In_791,In_1321);
and U54 (N_54,In_870,In_1197);
or U55 (N_55,In_1295,In_258);
or U56 (N_56,In_198,In_15);
and U57 (N_57,In_148,In_1015);
xor U58 (N_58,In_1466,In_320);
nor U59 (N_59,In_1112,In_516);
xor U60 (N_60,In_1423,In_1355);
xor U61 (N_61,In_1187,In_33);
xor U62 (N_62,In_482,In_526);
and U63 (N_63,In_232,In_499);
nand U64 (N_64,In_51,In_85);
and U65 (N_65,In_690,In_1099);
nor U66 (N_66,In_111,In_531);
nand U67 (N_67,In_1144,In_1141);
xnor U68 (N_68,In_115,In_491);
and U69 (N_69,In_127,In_1287);
and U70 (N_70,In_1292,In_804);
nor U71 (N_71,In_411,In_1020);
nor U72 (N_72,In_533,In_1189);
nor U73 (N_73,In_1350,In_110);
and U74 (N_74,In_729,In_354);
or U75 (N_75,In_1199,In_67);
nor U76 (N_76,In_728,In_1431);
nor U77 (N_77,In_893,In_1453);
nand U78 (N_78,In_206,In_1476);
nor U79 (N_79,In_501,In_240);
nor U80 (N_80,In_284,In_1336);
and U81 (N_81,In_614,In_611);
xor U82 (N_82,In_14,In_759);
xor U83 (N_83,In_955,In_973);
xor U84 (N_84,In_933,In_53);
xnor U85 (N_85,In_1190,In_1404);
or U86 (N_86,In_89,In_795);
or U87 (N_87,In_1014,In_596);
xor U88 (N_88,In_433,In_267);
nor U89 (N_89,In_694,In_1215);
and U90 (N_90,In_1449,In_382);
and U91 (N_91,In_1125,In_898);
xor U92 (N_92,In_1227,In_487);
nor U93 (N_93,In_852,In_1216);
and U94 (N_94,In_1102,In_364);
nand U95 (N_95,In_1145,In_1038);
nor U96 (N_96,In_1054,In_813);
xor U97 (N_97,In_266,In_1369);
or U98 (N_98,In_254,In_191);
xor U99 (N_99,In_609,In_202);
nand U100 (N_100,In_243,In_639);
and U101 (N_101,In_146,In_233);
nand U102 (N_102,In_763,In_1446);
nor U103 (N_103,In_176,In_1098);
or U104 (N_104,In_1450,In_397);
or U105 (N_105,In_918,In_801);
and U106 (N_106,In_981,In_151);
and U107 (N_107,In_782,In_542);
or U108 (N_108,In_1044,In_959);
or U109 (N_109,In_536,In_885);
xor U110 (N_110,In_541,In_58);
xnor U111 (N_111,In_432,In_527);
or U112 (N_112,In_477,In_478);
nand U113 (N_113,In_1314,In_373);
nand U114 (N_114,In_17,In_1346);
and U115 (N_115,In_335,In_102);
nand U116 (N_116,In_437,In_1400);
nand U117 (N_117,In_384,In_293);
and U118 (N_118,In_31,In_901);
or U119 (N_119,In_1313,In_294);
or U120 (N_120,In_913,In_90);
nor U121 (N_121,In_1322,In_704);
xnor U122 (N_122,In_1209,In_161);
nand U123 (N_123,In_696,In_949);
and U124 (N_124,In_1375,In_731);
and U125 (N_125,In_806,In_1288);
nand U126 (N_126,In_361,In_948);
nor U127 (N_127,In_922,In_498);
and U128 (N_128,In_50,In_1152);
xnor U129 (N_129,In_1135,In_1303);
nand U130 (N_130,In_117,In_304);
xor U131 (N_131,In_758,In_908);
and U132 (N_132,In_214,In_896);
xor U133 (N_133,In_1348,In_43);
or U134 (N_134,In_668,In_507);
nand U135 (N_135,In_1195,In_1034);
nor U136 (N_136,In_1132,In_1156);
xor U137 (N_137,In_911,In_986);
xnor U138 (N_138,In_174,In_86);
or U139 (N_139,In_504,In_428);
or U140 (N_140,In_100,In_57);
nand U141 (N_141,In_680,In_707);
nand U142 (N_142,In_888,In_967);
or U143 (N_143,In_339,In_917);
and U144 (N_144,In_640,In_952);
or U145 (N_145,In_841,In_204);
nor U146 (N_146,In_832,In_851);
nor U147 (N_147,In_509,In_878);
nor U148 (N_148,In_965,In_711);
or U149 (N_149,In_855,In_595);
and U150 (N_150,In_626,In_1424);
and U151 (N_151,In_1003,In_1155);
xnor U152 (N_152,In_653,In_1010);
nand U153 (N_153,In_916,In_462);
or U154 (N_154,In_407,In_788);
nand U155 (N_155,In_288,In_565);
nor U156 (N_156,In_289,In_1270);
or U157 (N_157,In_49,In_378);
xor U158 (N_158,In_1403,In_340);
or U159 (N_159,In_657,In_1159);
xor U160 (N_160,In_377,In_492);
nand U161 (N_161,In_875,In_332);
or U162 (N_162,In_1205,In_449);
or U163 (N_163,In_356,In_1071);
or U164 (N_164,In_1267,In_1301);
or U165 (N_165,In_996,In_26);
or U166 (N_166,In_1177,In_173);
and U167 (N_167,In_760,In_1256);
xor U168 (N_168,In_309,In_1234);
and U169 (N_169,In_963,In_941);
nand U170 (N_170,In_235,In_582);
and U171 (N_171,In_1006,In_1000);
nor U172 (N_172,In_617,In_1334);
or U173 (N_173,In_671,In_262);
xor U174 (N_174,In_27,In_107);
or U175 (N_175,In_141,In_969);
nor U176 (N_176,In_353,In_1291);
nand U177 (N_177,In_1276,In_66);
nand U178 (N_178,In_826,In_1327);
nand U179 (N_179,In_909,In_474);
nand U180 (N_180,In_37,In_1248);
or U181 (N_181,In_444,In_693);
or U182 (N_182,In_281,In_46);
nor U183 (N_183,In_140,In_834);
and U184 (N_184,In_403,In_305);
or U185 (N_185,In_1384,In_131);
or U186 (N_186,In_508,In_1078);
nor U187 (N_187,In_464,In_497);
nand U188 (N_188,In_94,In_1352);
and U189 (N_189,In_301,In_616);
nor U190 (N_190,In_914,In_1490);
nor U191 (N_191,In_1494,In_417);
nand U192 (N_192,In_456,In_1377);
nand U193 (N_193,In_1307,In_710);
xor U194 (N_194,In_1207,In_1457);
or U195 (N_195,In_1019,In_1376);
and U196 (N_196,In_580,In_956);
nor U197 (N_197,In_1139,In_1039);
nand U198 (N_198,In_158,In_1442);
nor U199 (N_199,In_521,In_39);
or U200 (N_200,In_1341,In_1421);
and U201 (N_201,In_1368,In_358);
nor U202 (N_202,In_264,In_257);
nand U203 (N_203,In_1485,In_29);
nor U204 (N_204,In_730,In_1232);
and U205 (N_205,In_613,In_472);
nand U206 (N_206,In_128,In_942);
xnor U207 (N_207,In_1488,In_346);
xor U208 (N_208,In_1005,In_726);
xor U209 (N_209,In_674,In_1395);
or U210 (N_210,In_194,In_1343);
nand U211 (N_211,In_578,In_1175);
and U212 (N_212,In_180,In_196);
nand U213 (N_213,In_16,In_1242);
nand U214 (N_214,In_1436,In_669);
nor U215 (N_215,In_253,In_594);
and U216 (N_216,In_786,In_621);
and U217 (N_217,In_54,In_8);
and U218 (N_218,In_1394,In_485);
nand U219 (N_219,In_1275,In_1304);
nor U220 (N_220,In_610,In_261);
or U221 (N_221,In_351,In_524);
nor U222 (N_222,In_650,In_290);
nor U223 (N_223,In_576,In_87);
and U224 (N_224,In_818,In_1086);
xor U225 (N_225,In_227,In_457);
or U226 (N_226,In_388,In_925);
nor U227 (N_227,In_1241,In_1133);
and U228 (N_228,In_1185,In_877);
and U229 (N_229,In_1076,In_139);
nand U230 (N_230,In_239,In_22);
and U231 (N_231,In_318,In_4);
and U232 (N_232,In_1188,In_514);
nor U233 (N_233,In_292,In_1059);
nor U234 (N_234,In_1122,In_1496);
xnor U235 (N_235,In_793,In_1481);
nand U236 (N_236,In_276,In_298);
nand U237 (N_237,In_404,In_1251);
nand U238 (N_238,In_28,In_566);
and U239 (N_239,In_633,In_995);
and U240 (N_240,In_463,In_1290);
xnor U241 (N_241,In_13,In_1069);
and U242 (N_242,In_300,In_242);
and U243 (N_243,In_11,In_904);
nand U244 (N_244,In_459,In_977);
nor U245 (N_245,In_334,In_836);
xnor U246 (N_246,In_329,In_951);
nor U247 (N_247,In_315,In_1254);
or U248 (N_248,In_1374,In_859);
or U249 (N_249,In_530,In_1398);
and U250 (N_250,In_418,In_1339);
nor U251 (N_251,In_0,In_980);
and U252 (N_252,In_495,In_455);
nor U253 (N_253,In_1470,In_1);
or U254 (N_254,In_819,In_628);
nand U255 (N_255,In_988,In_224);
and U256 (N_256,In_775,In_231);
nand U257 (N_257,In_30,In_1130);
nor U258 (N_258,In_953,In_355);
xnor U259 (N_259,In_717,In_1153);
nand U260 (N_260,In_9,In_520);
nand U261 (N_261,In_143,In_1140);
and U262 (N_262,In_1060,In_1171);
nand U263 (N_263,In_1306,In_1312);
or U264 (N_264,In_894,In_38);
and U265 (N_265,In_1486,In_557);
xnor U266 (N_266,In_1338,In_116);
nand U267 (N_267,In_1057,In_1027);
nor U268 (N_268,In_1382,In_1411);
nand U269 (N_269,In_714,In_220);
or U270 (N_270,In_1021,In_23);
nor U271 (N_271,In_1084,In_1274);
or U272 (N_272,In_1357,In_466);
and U273 (N_273,In_394,In_1447);
and U274 (N_274,In_550,In_1366);
xnor U275 (N_275,In_1364,In_559);
xnor U276 (N_276,In_752,In_1316);
and U277 (N_277,In_1178,In_109);
and U278 (N_278,In_658,In_1249);
nor U279 (N_279,In_145,In_427);
or U280 (N_280,In_776,In_480);
nor U281 (N_281,In_745,In_1217);
or U282 (N_282,In_751,In_259);
or U283 (N_283,In_957,In_1220);
or U284 (N_284,In_1337,In_519);
nand U285 (N_285,In_436,In_376);
and U286 (N_286,In_1271,In_1407);
xnor U287 (N_287,In_1479,In_544);
and U288 (N_288,In_405,In_1219);
nor U289 (N_289,In_844,In_842);
and U290 (N_290,In_121,In_175);
xor U291 (N_291,In_1041,In_853);
or U292 (N_292,In_372,In_134);
or U293 (N_293,In_63,In_1087);
xnor U294 (N_294,In_390,In_1058);
nor U295 (N_295,In_907,In_814);
and U296 (N_296,In_581,In_1113);
and U297 (N_297,In_1218,In_119);
or U298 (N_298,In_1162,In_858);
or U299 (N_299,In_60,In_347);
nor U300 (N_300,In_764,In_920);
or U301 (N_301,In_638,In_1282);
nor U302 (N_302,In_169,In_476);
nand U303 (N_303,In_1465,In_825);
nand U304 (N_304,In_1151,In_719);
and U305 (N_305,In_45,In_1438);
xnor U306 (N_306,In_919,In_811);
or U307 (N_307,In_1443,In_1298);
xor U308 (N_308,In_1356,In_1333);
and U309 (N_309,In_1131,In_664);
or U310 (N_310,In_165,In_1370);
xor U311 (N_311,In_207,In_568);
or U312 (N_312,In_186,In_551);
xor U313 (N_313,In_310,In_1016);
or U314 (N_314,In_1229,In_518);
or U315 (N_315,In_381,In_1154);
xor U316 (N_316,In_794,In_1428);
or U317 (N_317,In_398,In_1260);
nand U318 (N_318,In_1280,In_839);
and U319 (N_319,In_932,In_25);
xor U320 (N_320,In_352,In_150);
nor U321 (N_321,In_1007,In_984);
or U322 (N_322,In_879,In_1426);
and U323 (N_323,In_589,In_1097);
nor U324 (N_324,In_448,In_1286);
and U325 (N_325,In_77,In_881);
nor U326 (N_326,In_83,In_172);
and U327 (N_327,In_153,In_1165);
and U328 (N_328,In_425,In_871);
xnor U329 (N_329,In_748,In_64);
nor U330 (N_330,In_1167,In_891);
or U331 (N_331,In_387,In_935);
xor U332 (N_332,In_159,In_273);
and U333 (N_333,In_992,In_1080);
and U334 (N_334,In_1458,In_1250);
xnor U335 (N_335,In_35,In_692);
or U336 (N_336,In_1401,In_451);
nor U337 (N_337,In_213,In_1179);
xor U338 (N_338,In_1422,In_1115);
and U339 (N_339,In_212,In_777);
nor U340 (N_340,In_649,In_168);
nor U341 (N_341,In_241,In_856);
and U342 (N_342,In_635,In_47);
or U343 (N_343,In_1103,In_838);
nor U344 (N_344,In_6,In_1226);
or U345 (N_345,In_1067,In_36);
and U346 (N_346,In_249,In_781);
xnor U347 (N_347,In_1186,In_156);
or U348 (N_348,In_1385,In_431);
nor U349 (N_349,In_92,In_979);
nand U350 (N_350,In_602,In_1104);
xor U351 (N_351,In_337,In_1092);
and U352 (N_352,In_829,In_1347);
xor U353 (N_353,In_990,In_256);
nand U354 (N_354,In_1491,In_97);
nand U355 (N_355,In_319,In_489);
nor U356 (N_356,In_1011,In_438);
xnor U357 (N_357,In_152,In_221);
or U358 (N_358,In_265,In_24);
xor U359 (N_359,In_586,In_210);
nand U360 (N_360,In_506,In_286);
xnor U361 (N_361,In_647,In_1149);
nor U362 (N_362,In_1473,In_197);
nor U363 (N_363,In_467,In_744);
nand U364 (N_364,In_1127,In_229);
or U365 (N_365,In_816,In_1389);
nor U366 (N_366,In_1191,In_481);
xnor U367 (N_367,In_424,In_1469);
nor U368 (N_368,In_81,In_723);
nor U369 (N_369,In_890,In_74);
or U370 (N_370,In_753,In_1224);
and U371 (N_371,In_1325,In_252);
or U372 (N_372,In_488,In_588);
or U373 (N_373,In_685,In_307);
or U374 (N_374,In_1056,In_399);
xnor U375 (N_375,In_1413,In_648);
nor U376 (N_376,In_246,In_99);
nand U377 (N_377,In_848,In_303);
and U378 (N_378,In_446,In_938);
nand U379 (N_379,In_503,In_208);
nor U380 (N_380,In_426,In_1383);
or U381 (N_381,In_600,In_1213);
or U382 (N_382,In_1420,In_865);
nor U383 (N_383,In_326,In_473);
or U384 (N_384,In_385,In_1117);
xnor U385 (N_385,In_715,In_190);
or U386 (N_386,In_1497,In_1150);
and U387 (N_387,In_1246,In_940);
nor U388 (N_388,In_802,In_987);
xor U389 (N_389,In_867,In_366);
xor U390 (N_390,In_1048,In_1182);
or U391 (N_391,In_742,In_178);
nand U392 (N_392,In_1397,In_691);
xor U393 (N_393,In_539,In_285);
nand U394 (N_394,In_1063,In_934);
nor U395 (N_395,In_154,In_652);
or U396 (N_396,In_1045,In_924);
nor U397 (N_397,In_972,In_593);
nand U398 (N_398,In_1425,In_1354);
and U399 (N_399,In_113,In_1387);
nor U400 (N_400,In_654,In_423);
nor U401 (N_401,In_1430,In_106);
or U402 (N_402,In_1004,In_958);
xor U403 (N_403,In_72,In_1261);
nand U404 (N_404,In_1289,In_831);
xor U405 (N_405,In_1483,In_1362);
and U406 (N_406,In_768,In_1172);
xor U407 (N_407,In_1192,In_443);
and U408 (N_408,In_1123,In_1022);
nor U409 (N_409,In_549,In_400);
and U410 (N_410,In_590,In_359);
nor U411 (N_411,In_961,In_1464);
nor U412 (N_412,In_93,In_1475);
nand U413 (N_413,In_177,In_1367);
xnor U414 (N_414,In_1085,In_391);
and U415 (N_415,In_608,In_211);
xor U416 (N_416,In_1157,In_389);
nand U417 (N_417,In_637,In_1353);
and U418 (N_418,In_357,In_1128);
nand U419 (N_419,In_529,In_1296);
xnor U420 (N_420,In_234,In_325);
xor U421 (N_421,In_413,In_135);
and U422 (N_422,In_486,In_705);
nor U423 (N_423,In_269,In_1444);
or U424 (N_424,In_1221,In_732);
nand U425 (N_425,In_822,In_328);
and U426 (N_426,In_659,In_1033);
nor U427 (N_427,In_1342,In_338);
nand U428 (N_428,In_287,In_1416);
or U429 (N_429,In_755,In_906);
xor U430 (N_430,In_414,In_708);
nor U431 (N_431,In_1462,In_721);
nor U432 (N_432,In_716,In_584);
xnor U433 (N_433,In_1110,In_163);
nand U434 (N_434,In_749,In_1134);
nor U435 (N_435,In_1029,In_160);
xnor U436 (N_436,In_564,In_567);
and U437 (N_437,In_324,In_279);
xor U438 (N_438,In_1440,In_624);
xnor U439 (N_439,In_1499,In_496);
xor U440 (N_440,In_461,In_189);
nand U441 (N_441,In_968,In_629);
nor U442 (N_442,In_741,In_569);
or U443 (N_443,In_767,In_452);
or U444 (N_444,In_1380,In_720);
and U445 (N_445,In_681,In_1456);
or U446 (N_446,In_792,In_251);
xnor U447 (N_447,In_1448,In_1210);
nor U448 (N_448,In_62,In_1028);
or U449 (N_449,In_662,In_1433);
xor U450 (N_450,In_1332,In_114);
nand U451 (N_451,In_306,In_447);
nor U452 (N_452,In_1378,In_170);
nor U453 (N_453,In_157,In_1240);
or U454 (N_454,In_55,In_944);
xnor U455 (N_455,In_606,In_736);
nand U456 (N_456,In_1351,In_1090);
and U457 (N_457,In_1441,In_1247);
or U458 (N_458,In_1281,In_700);
and U459 (N_459,In_579,In_620);
and U460 (N_460,In_695,In_500);
xor U461 (N_461,In_401,In_236);
xor U462 (N_462,In_1393,In_1166);
and U463 (N_463,In_702,In_1273);
nand U464 (N_464,In_845,In_1230);
nand U465 (N_465,In_311,In_1434);
nor U466 (N_466,In_750,In_651);
or U467 (N_467,In_740,In_607);
or U468 (N_468,In_1032,In_228);
nand U469 (N_469,In_270,In_666);
or U470 (N_470,In_1238,In_954);
xor U471 (N_471,In_1231,In_623);
nand U472 (N_472,In_395,In_96);
nor U473 (N_473,In_1451,In_69);
nor U474 (N_474,In_192,In_1050);
nor U475 (N_475,In_59,In_1083);
nor U476 (N_476,In_1244,In_644);
xnor U477 (N_477,In_188,In_1202);
nand U478 (N_478,In_1065,In_622);
and U479 (N_479,In_209,In_1459);
nand U480 (N_480,In_677,In_846);
and U481 (N_481,In_678,In_1373);
nand U482 (N_482,In_1108,In_1168);
and U483 (N_483,In_910,In_103);
nor U484 (N_484,In_840,In_1262);
xnor U485 (N_485,In_317,In_316);
and U486 (N_486,In_1066,In_773);
xnor U487 (N_487,In_928,In_833);
nand U488 (N_488,In_1064,In_291);
nor U489 (N_489,In_703,In_808);
or U490 (N_490,In_634,In_603);
xor U491 (N_491,In_1452,In_1236);
or U492 (N_492,In_713,In_528);
nand U493 (N_493,In_470,In_375);
and U494 (N_494,In_921,In_815);
or U495 (N_495,In_1164,In_902);
xnor U496 (N_496,In_718,In_484);
nand U497 (N_497,In_1062,In_430);
and U498 (N_498,In_1300,In_857);
nand U499 (N_499,In_183,In_412);
or U500 (N_500,In_1297,In_80);
xnor U501 (N_501,In_1265,In_343);
or U502 (N_502,In_860,In_812);
nand U503 (N_503,In_1468,In_863);
nor U504 (N_504,In_1158,In_493);
xor U505 (N_505,In_998,In_563);
nand U506 (N_506,In_126,In_1467);
nand U507 (N_507,In_321,In_670);
nand U508 (N_508,In_667,In_1121);
xor U509 (N_509,In_517,In_962);
and U510 (N_510,In_761,In_556);
xor U511 (N_511,In_380,In_835);
xor U512 (N_512,In_1235,In_747);
and U513 (N_513,In_999,In_612);
and U514 (N_514,In_660,In_547);
nand U515 (N_515,In_1257,In_724);
nand U516 (N_516,In_483,In_1212);
xor U517 (N_517,In_1208,In_420);
or U518 (N_518,In_1174,In_960);
nand U519 (N_519,In_76,In_575);
nand U520 (N_520,In_1317,In_1169);
or U521 (N_521,In_278,In_1435);
and U522 (N_522,In_739,In_1204);
xor U523 (N_523,In_1495,In_383);
and U524 (N_524,In_1318,In_1049);
nand U525 (N_525,In_7,In_296);
or U526 (N_526,In_555,In_248);
xnor U527 (N_527,In_1417,In_737);
or U528 (N_528,In_989,In_283);
and U529 (N_529,In_510,In_1439);
and U530 (N_530,In_479,In_827);
nor U531 (N_531,In_854,In_709);
xnor U532 (N_532,In_323,In_84);
xnor U533 (N_533,In_1255,In_1143);
xor U534 (N_534,In_1017,In_201);
or U535 (N_535,In_1361,In_441);
or U536 (N_536,In_895,In_915);
or U537 (N_537,In_280,In_44);
or U538 (N_538,In_469,In_866);
and U539 (N_539,In_1088,In_125);
nor U540 (N_540,In_1414,In_68);
xor U541 (N_541,In_1478,In_785);
nor U542 (N_542,In_861,In_112);
nand U543 (N_543,In_1461,In_545);
nor U544 (N_544,In_1419,In_1148);
and U545 (N_545,In_683,In_129);
xor U546 (N_546,In_1040,In_1477);
and U547 (N_547,In_421,In_886);
xnor U548 (N_548,In_1319,In_1126);
nand U549 (N_549,In_926,In_630);
and U550 (N_550,In_226,In_422);
nand U551 (N_551,In_1035,In_181);
nand U552 (N_552,In_350,In_1379);
nor U553 (N_553,In_618,In_274);
and U554 (N_554,In_874,In_1046);
or U555 (N_555,In_20,In_561);
or U556 (N_556,In_673,In_892);
nor U557 (N_557,In_558,In_105);
or U558 (N_558,In_1008,In_676);
xnor U559 (N_559,In_179,In_873);
nor U560 (N_560,In_598,In_120);
nand U561 (N_561,In_1018,In_1079);
or U562 (N_562,In_1454,In_402);
or U563 (N_563,In_98,In_1091);
xnor U564 (N_564,In_1269,In_1284);
nand U565 (N_565,In_950,In_73);
or U566 (N_566,In_1176,In_52);
and U567 (N_567,In_1358,In_1043);
xor U568 (N_568,In_684,In_1302);
and U569 (N_569,In_2,In_522);
or U570 (N_570,In_458,In_661);
or U571 (N_571,In_1460,In_454);
xnor U572 (N_572,In_245,In_1237);
and U573 (N_573,In_1493,In_884);
nor U574 (N_574,In_665,In_1359);
or U575 (N_575,In_738,In_939);
nor U576 (N_576,In_1228,In_679);
xnor U577 (N_577,In_936,In_142);
and U578 (N_578,In_770,In_1335);
xor U579 (N_579,In_1363,In_880);
xnor U580 (N_580,In_757,In_439);
or U581 (N_581,In_505,In_682);
xor U582 (N_582,In_1243,In_689);
nor U583 (N_583,In_1399,In_552);
xor U584 (N_584,In_434,In_540);
nand U585 (N_585,In_1258,In_1194);
nand U586 (N_586,In_727,In_19);
nand U587 (N_587,In_577,In_1206);
nor U588 (N_588,In_572,In_435);
or U589 (N_589,In_193,In_805);
and U590 (N_590,In_765,In_619);
or U591 (N_591,In_133,In_1391);
nand U592 (N_592,In_1119,In_797);
nor U593 (N_593,In_1036,In_780);
nor U594 (N_594,In_396,In_101);
nand U595 (N_595,In_1201,In_1412);
and U596 (N_596,In_1408,In_1309);
or U597 (N_597,In_42,In_445);
nor U598 (N_598,In_820,In_1106);
nor U599 (N_599,In_429,In_1160);
nand U600 (N_600,In_419,In_535);
nor U601 (N_601,In_460,In_41);
xnor U602 (N_602,In_1026,In_271);
nor U603 (N_603,In_725,In_147);
or U604 (N_604,In_1047,In_118);
and U605 (N_605,In_3,In_543);
nor U606 (N_606,In_735,In_548);
and U607 (N_607,In_1455,In_991);
nor U608 (N_608,In_342,In_371);
nor U609 (N_609,In_897,In_697);
or U610 (N_610,In_1013,In_122);
xnor U611 (N_611,In_330,In_1427);
and U612 (N_612,In_1372,In_1081);
nor U613 (N_613,In_406,In_370);
or U614 (N_614,In_937,In_1471);
and U615 (N_615,In_1445,In_975);
xor U616 (N_616,In_302,In_1308);
xnor U617 (N_617,In_591,In_1137);
nor U618 (N_618,In_1180,In_1329);
or U619 (N_619,In_1252,In_699);
nand U620 (N_620,In_48,In_1114);
and U621 (N_621,In_1196,In_187);
xor U622 (N_622,In_756,In_1120);
or U623 (N_623,In_642,In_255);
nand U624 (N_624,In_538,In_970);
or U625 (N_625,In_821,In_1198);
or U626 (N_626,In_344,In_1396);
nand U627 (N_627,In_1183,In_787);
or U628 (N_628,In_1406,In_1415);
xor U629 (N_629,In_1340,In_468);
xnor U630 (N_630,In_1283,In_513);
and U631 (N_631,In_91,In_312);
nand U632 (N_632,In_345,In_1344);
xnor U633 (N_633,In_966,In_362);
nor U634 (N_634,In_471,In_1107);
nor U635 (N_635,In_1381,In_766);
nor U636 (N_636,In_1025,In_1263);
and U637 (N_637,In_1233,In_1225);
or U638 (N_638,In_546,In_574);
nand U639 (N_639,In_333,In_706);
nand U640 (N_640,In_946,In_636);
xnor U641 (N_641,In_1001,In_199);
nand U642 (N_642,In_1484,In_1012);
nand U643 (N_643,In_225,In_263);
xnor U644 (N_644,In_367,In_930);
or U645 (N_645,In_1147,In_260);
xor U646 (N_646,In_1331,In_883);
xnor U647 (N_647,In_772,In_1474);
xor U648 (N_648,In_1055,In_570);
xnor U649 (N_649,In_1223,In_1326);
and U650 (N_650,In_643,In_945);
nand U651 (N_651,In_453,In_1037);
and U652 (N_652,In_983,In_1094);
and U653 (N_653,In_1371,In_889);
nor U654 (N_654,In_386,In_778);
nand U655 (N_655,In_882,In_656);
nand U656 (N_656,In_104,In_132);
nand U657 (N_657,In_88,In_1328);
nand U658 (N_658,In_1072,In_1193);
nand U659 (N_659,In_1136,In_994);
or U660 (N_660,In_790,In_230);
xnor U661 (N_661,In_61,In_1138);
or U662 (N_662,In_900,In_899);
nor U663 (N_663,In_828,In_605);
nand U664 (N_664,In_218,In_416);
nor U665 (N_665,In_250,In_1009);
xor U666 (N_666,In_12,In_675);
xnor U667 (N_667,In_1365,In_864);
and U668 (N_668,In_21,In_162);
or U669 (N_669,In_217,In_1214);
xnor U670 (N_670,In_379,In_365);
and U671 (N_671,In_1487,In_779);
nand U672 (N_672,In_511,In_138);
or U673 (N_673,In_1109,In_1031);
xor U674 (N_674,In_872,In_95);
or U675 (N_675,In_655,In_830);
or U676 (N_676,In_1173,In_184);
nand U677 (N_677,In_823,In_645);
xor U678 (N_678,In_712,In_247);
and U679 (N_679,In_331,In_1277);
nor U680 (N_680,In_297,In_796);
xnor U681 (N_681,In_409,In_79);
and U682 (N_682,In_1293,In_108);
nor U683 (N_683,In_223,In_1272);
xor U684 (N_684,In_974,In_585);
nor U685 (N_685,In_985,In_5);
nor U686 (N_686,In_868,In_807);
or U687 (N_687,In_1390,In_597);
or U688 (N_688,In_393,In_1052);
nand U689 (N_689,In_203,In_905);
or U690 (N_690,In_771,In_124);
or U691 (N_691,In_155,In_1200);
xnor U692 (N_692,In_698,In_604);
xor U693 (N_693,In_784,In_465);
nand U694 (N_694,In_244,In_646);
nor U695 (N_695,In_562,In_734);
and U696 (N_696,In_632,In_144);
xor U697 (N_697,In_322,In_1402);
or U698 (N_698,In_408,In_869);
or U699 (N_699,In_532,In_1024);
nand U700 (N_700,In_1124,In_363);
or U701 (N_701,In_573,In_34);
or U702 (N_702,In_137,In_1305);
nor U703 (N_703,In_490,In_277);
nor U704 (N_704,In_1051,In_182);
xnor U705 (N_705,In_1222,In_299);
nor U706 (N_706,In_336,In_733);
and U707 (N_707,In_238,In_722);
or U708 (N_708,In_56,In_185);
and U709 (N_709,In_515,In_837);
nand U710 (N_710,In_360,In_912);
and U711 (N_711,In_65,In_1324);
nand U712 (N_712,In_783,In_663);
and U713 (N_713,In_40,In_1268);
nand U714 (N_714,In_803,In_927);
xnor U715 (N_715,In_847,In_1299);
and U716 (N_716,In_1211,In_1118);
xor U717 (N_717,In_1095,In_32);
xor U718 (N_718,In_1266,In_136);
nor U719 (N_719,In_1320,In_1100);
xnor U720 (N_720,In_1405,In_1184);
and U721 (N_721,In_1323,In_762);
nand U722 (N_722,In_1061,In_282);
nor U723 (N_723,In_1349,In_1203);
and U724 (N_724,In_798,In_272);
or U725 (N_725,In_1142,In_534);
or U726 (N_726,In_1310,In_1360);
or U727 (N_727,In_392,In_601);
and U728 (N_728,In_1330,In_200);
and U729 (N_729,In_1279,In_171);
nor U730 (N_730,In_1264,In_824);
nand U731 (N_731,In_195,In_931);
or U732 (N_732,In_876,In_1392);
xnor U733 (N_733,In_554,In_18);
nor U734 (N_734,In_295,In_1278);
and U735 (N_735,In_592,In_1482);
nor U736 (N_736,In_1053,In_862);
xor U737 (N_737,In_843,In_1315);
nor U738 (N_738,In_219,In_571);
nand U739 (N_739,In_1023,In_166);
or U740 (N_740,In_993,In_442);
nor U741 (N_741,In_450,In_743);
or U742 (N_742,In_1437,In_215);
nor U743 (N_743,In_599,In_149);
and U744 (N_744,In_754,In_887);
nor U745 (N_745,In_275,In_1170);
xnor U746 (N_746,In_1386,In_583);
or U747 (N_747,In_308,In_1146);
nand U748 (N_748,In_799,In_1409);
and U749 (N_749,In_971,In_1345);
xnor U750 (N_750,N_349,N_505);
nor U751 (N_751,N_248,N_458);
nand U752 (N_752,N_176,N_744);
and U753 (N_753,N_296,N_160);
and U754 (N_754,N_312,N_132);
and U755 (N_755,N_613,N_181);
nor U756 (N_756,N_179,N_426);
xnor U757 (N_757,N_182,N_95);
nand U758 (N_758,N_609,N_249);
and U759 (N_759,N_114,N_136);
and U760 (N_760,N_237,N_428);
xor U761 (N_761,N_251,N_683);
nor U762 (N_762,N_516,N_412);
nand U763 (N_763,N_39,N_134);
or U764 (N_764,N_702,N_605);
or U765 (N_765,N_603,N_684);
and U766 (N_766,N_719,N_653);
nand U767 (N_767,N_654,N_642);
nand U768 (N_768,N_727,N_746);
nand U769 (N_769,N_690,N_451);
and U770 (N_770,N_229,N_682);
xor U771 (N_771,N_445,N_588);
nor U772 (N_772,N_265,N_630);
or U773 (N_773,N_26,N_244);
and U774 (N_774,N_224,N_383);
xor U775 (N_775,N_479,N_706);
nand U776 (N_776,N_292,N_128);
nor U777 (N_777,N_663,N_1);
nand U778 (N_778,N_384,N_679);
xnor U779 (N_779,N_204,N_146);
or U780 (N_780,N_531,N_396);
xor U781 (N_781,N_44,N_511);
xor U782 (N_782,N_632,N_199);
and U783 (N_783,N_133,N_164);
nand U784 (N_784,N_722,N_156);
nor U785 (N_785,N_194,N_404);
and U786 (N_786,N_638,N_636);
nor U787 (N_787,N_582,N_370);
and U788 (N_788,N_266,N_567);
nand U789 (N_789,N_232,N_399);
nor U790 (N_790,N_593,N_703);
or U791 (N_791,N_489,N_96);
nor U792 (N_792,N_523,N_284);
and U793 (N_793,N_621,N_358);
and U794 (N_794,N_619,N_587);
nand U795 (N_795,N_540,N_267);
xnor U796 (N_796,N_355,N_65);
nand U797 (N_797,N_699,N_502);
nor U798 (N_798,N_450,N_219);
nand U799 (N_799,N_749,N_692);
nor U800 (N_800,N_446,N_416);
and U801 (N_801,N_611,N_477);
or U802 (N_802,N_569,N_554);
nor U803 (N_803,N_592,N_409);
or U804 (N_804,N_51,N_710);
or U805 (N_805,N_165,N_467);
nand U806 (N_806,N_282,N_623);
nor U807 (N_807,N_71,N_549);
and U808 (N_808,N_131,N_494);
nand U809 (N_809,N_375,N_685);
xor U810 (N_810,N_264,N_483);
or U811 (N_811,N_741,N_138);
or U812 (N_812,N_401,N_414);
xnor U813 (N_813,N_308,N_303);
nand U814 (N_814,N_646,N_658);
xnor U815 (N_815,N_58,N_697);
xor U816 (N_816,N_336,N_7);
xnor U817 (N_817,N_513,N_640);
nor U818 (N_818,N_328,N_177);
or U819 (N_819,N_413,N_575);
nor U820 (N_820,N_148,N_661);
and U821 (N_821,N_88,N_22);
or U822 (N_822,N_363,N_717);
and U823 (N_823,N_166,N_147);
nor U824 (N_824,N_572,N_274);
nor U825 (N_825,N_2,N_493);
or U826 (N_826,N_535,N_169);
nor U827 (N_827,N_31,N_82);
nor U828 (N_828,N_422,N_288);
xnor U829 (N_829,N_651,N_610);
or U830 (N_830,N_634,N_258);
xnor U831 (N_831,N_120,N_631);
nor U832 (N_832,N_113,N_628);
xnor U833 (N_833,N_454,N_434);
nor U834 (N_834,N_544,N_55);
nand U835 (N_835,N_231,N_537);
nor U836 (N_836,N_298,N_254);
xor U837 (N_837,N_740,N_712);
xor U838 (N_838,N_589,N_217);
or U839 (N_839,N_691,N_644);
nand U840 (N_840,N_443,N_47);
nand U841 (N_841,N_559,N_275);
or U842 (N_842,N_607,N_686);
nand U843 (N_843,N_129,N_257);
or U844 (N_844,N_221,N_552);
xor U845 (N_845,N_294,N_645);
nand U846 (N_846,N_180,N_50);
or U847 (N_847,N_627,N_85);
nor U848 (N_848,N_102,N_208);
and U849 (N_849,N_243,N_361);
nor U850 (N_850,N_448,N_724);
nand U851 (N_851,N_737,N_36);
nand U852 (N_852,N_253,N_571);
or U853 (N_853,N_67,N_590);
and U854 (N_854,N_614,N_121);
or U855 (N_855,N_444,N_207);
nand U856 (N_856,N_551,N_186);
nand U857 (N_857,N_301,N_408);
nor U858 (N_858,N_564,N_704);
xnor U859 (N_859,N_256,N_278);
nand U860 (N_860,N_557,N_144);
or U861 (N_861,N_393,N_581);
or U862 (N_862,N_18,N_337);
xnor U863 (N_863,N_488,N_678);
nor U864 (N_864,N_512,N_608);
nor U865 (N_865,N_236,N_106);
and U866 (N_866,N_343,N_713);
nor U867 (N_867,N_385,N_565);
and U868 (N_868,N_212,N_570);
nand U869 (N_869,N_98,N_373);
or U870 (N_870,N_93,N_16);
and U871 (N_871,N_595,N_500);
xor U872 (N_872,N_46,N_354);
xor U873 (N_873,N_339,N_118);
or U874 (N_874,N_123,N_624);
xnor U875 (N_875,N_429,N_211);
nor U876 (N_876,N_470,N_9);
nor U877 (N_877,N_518,N_318);
and U878 (N_878,N_541,N_174);
and U879 (N_879,N_742,N_60);
and U880 (N_880,N_504,N_299);
xor U881 (N_881,N_352,N_226);
and U882 (N_882,N_140,N_234);
or U883 (N_883,N_24,N_492);
and U884 (N_884,N_242,N_161);
and U885 (N_885,N_364,N_250);
or U886 (N_886,N_472,N_302);
nand U887 (N_887,N_407,N_524);
nor U888 (N_888,N_320,N_379);
or U889 (N_889,N_525,N_403);
nand U890 (N_890,N_732,N_149);
nor U891 (N_891,N_402,N_708);
nand U892 (N_892,N_261,N_545);
or U893 (N_893,N_167,N_405);
and U894 (N_894,N_550,N_29);
nor U895 (N_895,N_272,N_304);
nand U896 (N_896,N_716,N_233);
or U897 (N_897,N_660,N_395);
xor U898 (N_898,N_69,N_720);
xnor U899 (N_899,N_455,N_476);
and U900 (N_900,N_707,N_310);
nand U901 (N_901,N_57,N_291);
nor U902 (N_902,N_345,N_473);
nor U903 (N_903,N_322,N_526);
nand U904 (N_904,N_745,N_17);
nor U905 (N_905,N_536,N_641);
or U906 (N_906,N_616,N_568);
and U907 (N_907,N_112,N_410);
and U908 (N_908,N_687,N_676);
nor U909 (N_909,N_425,N_665);
or U910 (N_910,N_681,N_73);
nor U911 (N_911,N_246,N_220);
and U912 (N_912,N_748,N_64);
nand U913 (N_913,N_319,N_270);
or U914 (N_914,N_184,N_225);
and U915 (N_915,N_10,N_306);
or U916 (N_916,N_81,N_464);
and U917 (N_917,N_323,N_91);
xor U918 (N_918,N_466,N_63);
and U919 (N_919,N_269,N_360);
xor U920 (N_920,N_675,N_390);
xor U921 (N_921,N_255,N_441);
nand U922 (N_922,N_736,N_152);
and U923 (N_923,N_538,N_259);
or U924 (N_924,N_239,N_327);
xor U925 (N_925,N_452,N_387);
nand U926 (N_926,N_490,N_100);
xor U927 (N_927,N_347,N_45);
and U928 (N_928,N_629,N_437);
and U929 (N_929,N_12,N_580);
nor U930 (N_930,N_594,N_200);
nand U931 (N_931,N_48,N_637);
or U932 (N_932,N_117,N_689);
xnor U933 (N_933,N_419,N_394);
nand U934 (N_934,N_725,N_238);
xor U935 (N_935,N_171,N_508);
nor U936 (N_936,N_438,N_190);
and U937 (N_937,N_203,N_87);
nor U938 (N_938,N_89,N_290);
nand U939 (N_939,N_101,N_596);
or U940 (N_940,N_527,N_78);
nand U941 (N_941,N_321,N_378);
or U942 (N_942,N_49,N_726);
nor U943 (N_943,N_427,N_421);
or U944 (N_944,N_655,N_365);
or U945 (N_945,N_649,N_617);
or U946 (N_946,N_4,N_701);
xor U947 (N_947,N_8,N_639);
and U948 (N_948,N_420,N_210);
or U949 (N_949,N_216,N_521);
xor U950 (N_950,N_397,N_495);
nand U951 (N_951,N_700,N_19);
xnor U952 (N_952,N_316,N_430);
or U953 (N_953,N_435,N_743);
xnor U954 (N_954,N_126,N_34);
or U955 (N_955,N_245,N_597);
nand U956 (N_956,N_626,N_280);
xnor U957 (N_957,N_356,N_546);
xor U958 (N_958,N_215,N_436);
or U959 (N_959,N_271,N_13);
nor U960 (N_960,N_417,N_670);
or U961 (N_961,N_656,N_547);
and U962 (N_962,N_664,N_75);
nand U963 (N_963,N_262,N_474);
nand U964 (N_964,N_730,N_372);
nand U965 (N_965,N_585,N_400);
nor U966 (N_966,N_449,N_173);
nor U967 (N_967,N_709,N_197);
nor U968 (N_968,N_315,N_469);
or U969 (N_969,N_62,N_103);
or U970 (N_970,N_108,N_20);
and U971 (N_971,N_38,N_612);
nand U972 (N_972,N_90,N_591);
or U973 (N_973,N_80,N_485);
nor U974 (N_974,N_558,N_346);
xnor U975 (N_975,N_507,N_159);
xnor U976 (N_976,N_309,N_622);
or U977 (N_977,N_137,N_53);
or U978 (N_978,N_520,N_338);
nor U979 (N_979,N_440,N_61);
nor U980 (N_980,N_382,N_293);
and U981 (N_981,N_295,N_528);
xor U982 (N_982,N_723,N_388);
or U983 (N_983,N_105,N_311);
nand U984 (N_984,N_335,N_668);
or U985 (N_985,N_718,N_84);
or U986 (N_986,N_353,N_579);
and U987 (N_987,N_228,N_139);
nor U988 (N_988,N_602,N_647);
or U989 (N_989,N_487,N_235);
and U990 (N_990,N_300,N_289);
xor U991 (N_991,N_68,N_556);
and U992 (N_992,N_94,N_42);
xnor U993 (N_993,N_344,N_202);
xnor U994 (N_994,N_715,N_209);
and U995 (N_995,N_376,N_178);
xnor U996 (N_996,N_462,N_35);
or U997 (N_997,N_650,N_460);
nand U998 (N_998,N_688,N_497);
nand U999 (N_999,N_643,N_56);
nor U1000 (N_1000,N_468,N_366);
or U1001 (N_1001,N_424,N_482);
xnor U1002 (N_1002,N_155,N_277);
or U1003 (N_1003,N_86,N_27);
or U1004 (N_1004,N_110,N_307);
or U1005 (N_1005,N_705,N_76);
and U1006 (N_1006,N_693,N_30);
and U1007 (N_1007,N_496,N_130);
and U1008 (N_1008,N_11,N_738);
nand U1009 (N_1009,N_386,N_195);
nor U1010 (N_1010,N_677,N_350);
nor U1011 (N_1011,N_368,N_423);
or U1012 (N_1012,N_331,N_442);
nand U1013 (N_1013,N_729,N_486);
xor U1014 (N_1014,N_620,N_187);
nor U1015 (N_1015,N_0,N_324);
nor U1016 (N_1016,N_14,N_218);
nand U1017 (N_1017,N_330,N_519);
xnor U1018 (N_1018,N_714,N_260);
nand U1019 (N_1019,N_533,N_534);
xnor U1020 (N_1020,N_247,N_97);
and U1021 (N_1021,N_21,N_584);
nand U1022 (N_1022,N_652,N_711);
and U1023 (N_1023,N_40,N_465);
xnor U1024 (N_1024,N_530,N_672);
nand U1025 (N_1025,N_15,N_453);
or U1026 (N_1026,N_532,N_633);
nand U1027 (N_1027,N_578,N_317);
nor U1028 (N_1028,N_214,N_109);
nand U1029 (N_1029,N_432,N_514);
or U1030 (N_1030,N_392,N_457);
xor U1031 (N_1031,N_124,N_111);
nor U1032 (N_1032,N_456,N_325);
xnor U1033 (N_1033,N_555,N_509);
nor U1034 (N_1034,N_380,N_116);
and U1035 (N_1035,N_285,N_539);
nor U1036 (N_1036,N_314,N_188);
nand U1037 (N_1037,N_566,N_189);
nor U1038 (N_1038,N_377,N_625);
nand U1039 (N_1039,N_433,N_41);
nor U1040 (N_1040,N_305,N_499);
xnor U1041 (N_1041,N_193,N_739);
xor U1042 (N_1042,N_598,N_562);
xnor U1043 (N_1043,N_600,N_279);
nand U1044 (N_1044,N_143,N_230);
nor U1045 (N_1045,N_313,N_475);
or U1046 (N_1046,N_406,N_669);
nor U1047 (N_1047,N_747,N_168);
xor U1048 (N_1048,N_104,N_563);
or U1049 (N_1049,N_601,N_28);
nor U1050 (N_1050,N_157,N_503);
nand U1051 (N_1051,N_150,N_648);
xor U1052 (N_1052,N_119,N_135);
and U1053 (N_1053,N_52,N_506);
and U1054 (N_1054,N_560,N_72);
nand U1055 (N_1055,N_240,N_471);
nand U1056 (N_1056,N_734,N_162);
and U1057 (N_1057,N_151,N_99);
nor U1058 (N_1058,N_79,N_59);
xor U1059 (N_1059,N_329,N_501);
nand U1060 (N_1060,N_498,N_359);
or U1061 (N_1061,N_192,N_342);
or U1062 (N_1062,N_674,N_273);
and U1063 (N_1063,N_6,N_107);
and U1064 (N_1064,N_543,N_696);
and U1065 (N_1065,N_695,N_389);
or U1066 (N_1066,N_206,N_721);
xor U1067 (N_1067,N_32,N_635);
nor U1068 (N_1068,N_196,N_263);
nor U1069 (N_1069,N_83,N_586);
nor U1070 (N_1070,N_334,N_573);
or U1071 (N_1071,N_680,N_43);
or U1072 (N_1072,N_276,N_333);
xor U1073 (N_1073,N_367,N_348);
xnor U1074 (N_1074,N_576,N_733);
nand U1075 (N_1075,N_529,N_3);
or U1076 (N_1076,N_418,N_115);
nand U1077 (N_1077,N_583,N_37);
nand U1078 (N_1078,N_522,N_542);
nand U1079 (N_1079,N_141,N_213);
and U1080 (N_1080,N_351,N_671);
nor U1081 (N_1081,N_698,N_172);
and U1082 (N_1082,N_369,N_731);
nor U1083 (N_1083,N_728,N_223);
nor U1084 (N_1084,N_125,N_183);
and U1085 (N_1085,N_23,N_25);
nor U1086 (N_1086,N_659,N_283);
nand U1087 (N_1087,N_484,N_510);
and U1088 (N_1088,N_371,N_574);
and U1089 (N_1089,N_175,N_381);
or U1090 (N_1090,N_415,N_252);
or U1091 (N_1091,N_673,N_326);
and U1092 (N_1092,N_158,N_447);
nand U1093 (N_1093,N_411,N_374);
nor U1094 (N_1094,N_548,N_205);
or U1095 (N_1095,N_201,N_145);
xor U1096 (N_1096,N_340,N_163);
xor U1097 (N_1097,N_153,N_478);
and U1098 (N_1098,N_599,N_77);
xnor U1099 (N_1099,N_281,N_391);
xor U1100 (N_1100,N_517,N_515);
nor U1101 (N_1101,N_694,N_431);
nand U1102 (N_1102,N_480,N_122);
nor U1103 (N_1103,N_463,N_222);
nand U1104 (N_1104,N_604,N_662);
nor U1105 (N_1105,N_92,N_170);
and U1106 (N_1106,N_398,N_54);
nand U1107 (N_1107,N_142,N_74);
xor U1108 (N_1108,N_666,N_577);
or U1109 (N_1109,N_481,N_198);
nor U1110 (N_1110,N_615,N_362);
nor U1111 (N_1111,N_561,N_268);
nor U1112 (N_1112,N_461,N_667);
nand U1113 (N_1113,N_227,N_297);
xor U1114 (N_1114,N_191,N_127);
or U1115 (N_1115,N_185,N_357);
or U1116 (N_1116,N_657,N_154);
nor U1117 (N_1117,N_491,N_439);
and U1118 (N_1118,N_287,N_66);
nand U1119 (N_1119,N_286,N_341);
or U1120 (N_1120,N_459,N_70);
nor U1121 (N_1121,N_735,N_618);
nand U1122 (N_1122,N_5,N_606);
or U1123 (N_1123,N_33,N_553);
or U1124 (N_1124,N_241,N_332);
xnor U1125 (N_1125,N_567,N_450);
nand U1126 (N_1126,N_318,N_462);
and U1127 (N_1127,N_362,N_688);
nand U1128 (N_1128,N_117,N_741);
or U1129 (N_1129,N_188,N_106);
or U1130 (N_1130,N_609,N_469);
and U1131 (N_1131,N_170,N_441);
nor U1132 (N_1132,N_150,N_256);
or U1133 (N_1133,N_350,N_35);
or U1134 (N_1134,N_287,N_54);
or U1135 (N_1135,N_317,N_504);
and U1136 (N_1136,N_633,N_456);
or U1137 (N_1137,N_527,N_354);
xnor U1138 (N_1138,N_520,N_304);
and U1139 (N_1139,N_24,N_578);
nor U1140 (N_1140,N_421,N_193);
or U1141 (N_1141,N_660,N_733);
nor U1142 (N_1142,N_640,N_358);
and U1143 (N_1143,N_616,N_476);
xor U1144 (N_1144,N_70,N_228);
and U1145 (N_1145,N_216,N_738);
xor U1146 (N_1146,N_503,N_613);
xor U1147 (N_1147,N_433,N_391);
xor U1148 (N_1148,N_385,N_199);
xnor U1149 (N_1149,N_411,N_239);
and U1150 (N_1150,N_60,N_319);
nor U1151 (N_1151,N_177,N_150);
nor U1152 (N_1152,N_649,N_586);
and U1153 (N_1153,N_247,N_180);
nand U1154 (N_1154,N_677,N_66);
or U1155 (N_1155,N_636,N_418);
or U1156 (N_1156,N_188,N_744);
nor U1157 (N_1157,N_37,N_267);
or U1158 (N_1158,N_234,N_288);
or U1159 (N_1159,N_496,N_299);
xor U1160 (N_1160,N_386,N_150);
xor U1161 (N_1161,N_583,N_719);
and U1162 (N_1162,N_630,N_45);
xnor U1163 (N_1163,N_84,N_342);
nand U1164 (N_1164,N_560,N_46);
xnor U1165 (N_1165,N_39,N_33);
nand U1166 (N_1166,N_267,N_352);
nor U1167 (N_1167,N_162,N_252);
nand U1168 (N_1168,N_484,N_377);
xor U1169 (N_1169,N_493,N_206);
or U1170 (N_1170,N_71,N_124);
or U1171 (N_1171,N_431,N_214);
nor U1172 (N_1172,N_133,N_645);
nor U1173 (N_1173,N_407,N_165);
xnor U1174 (N_1174,N_731,N_470);
and U1175 (N_1175,N_546,N_298);
nand U1176 (N_1176,N_504,N_231);
nand U1177 (N_1177,N_241,N_621);
or U1178 (N_1178,N_697,N_376);
and U1179 (N_1179,N_241,N_482);
xor U1180 (N_1180,N_488,N_605);
and U1181 (N_1181,N_90,N_253);
nor U1182 (N_1182,N_495,N_719);
or U1183 (N_1183,N_590,N_439);
xor U1184 (N_1184,N_292,N_84);
nor U1185 (N_1185,N_588,N_261);
or U1186 (N_1186,N_346,N_414);
nor U1187 (N_1187,N_563,N_157);
nand U1188 (N_1188,N_173,N_435);
or U1189 (N_1189,N_644,N_544);
xor U1190 (N_1190,N_293,N_356);
and U1191 (N_1191,N_100,N_530);
and U1192 (N_1192,N_529,N_164);
nor U1193 (N_1193,N_487,N_73);
nor U1194 (N_1194,N_255,N_695);
xor U1195 (N_1195,N_30,N_92);
nor U1196 (N_1196,N_375,N_336);
nor U1197 (N_1197,N_47,N_98);
and U1198 (N_1198,N_491,N_237);
nand U1199 (N_1199,N_94,N_334);
and U1200 (N_1200,N_559,N_240);
nand U1201 (N_1201,N_40,N_351);
nor U1202 (N_1202,N_239,N_216);
nor U1203 (N_1203,N_627,N_557);
xnor U1204 (N_1204,N_437,N_61);
and U1205 (N_1205,N_176,N_728);
xnor U1206 (N_1206,N_425,N_743);
nor U1207 (N_1207,N_155,N_642);
nand U1208 (N_1208,N_525,N_660);
nor U1209 (N_1209,N_449,N_122);
nor U1210 (N_1210,N_20,N_726);
nor U1211 (N_1211,N_10,N_289);
or U1212 (N_1212,N_150,N_195);
nor U1213 (N_1213,N_520,N_502);
xor U1214 (N_1214,N_662,N_278);
or U1215 (N_1215,N_644,N_632);
nand U1216 (N_1216,N_95,N_502);
and U1217 (N_1217,N_412,N_511);
nor U1218 (N_1218,N_726,N_512);
and U1219 (N_1219,N_160,N_608);
and U1220 (N_1220,N_32,N_37);
or U1221 (N_1221,N_274,N_129);
nand U1222 (N_1222,N_483,N_608);
and U1223 (N_1223,N_140,N_36);
nand U1224 (N_1224,N_244,N_91);
xnor U1225 (N_1225,N_238,N_533);
nand U1226 (N_1226,N_430,N_460);
xor U1227 (N_1227,N_399,N_569);
xnor U1228 (N_1228,N_638,N_218);
nand U1229 (N_1229,N_746,N_127);
and U1230 (N_1230,N_359,N_356);
nor U1231 (N_1231,N_192,N_170);
or U1232 (N_1232,N_103,N_625);
nor U1233 (N_1233,N_613,N_347);
or U1234 (N_1234,N_502,N_86);
or U1235 (N_1235,N_278,N_655);
nand U1236 (N_1236,N_590,N_456);
and U1237 (N_1237,N_704,N_45);
nor U1238 (N_1238,N_572,N_23);
nor U1239 (N_1239,N_58,N_65);
nand U1240 (N_1240,N_553,N_425);
or U1241 (N_1241,N_723,N_681);
nor U1242 (N_1242,N_171,N_716);
xnor U1243 (N_1243,N_19,N_163);
and U1244 (N_1244,N_69,N_640);
nand U1245 (N_1245,N_652,N_531);
nor U1246 (N_1246,N_378,N_309);
and U1247 (N_1247,N_312,N_310);
xnor U1248 (N_1248,N_571,N_427);
nor U1249 (N_1249,N_427,N_8);
nor U1250 (N_1250,N_24,N_47);
and U1251 (N_1251,N_349,N_234);
nor U1252 (N_1252,N_356,N_533);
xnor U1253 (N_1253,N_694,N_362);
and U1254 (N_1254,N_313,N_172);
nor U1255 (N_1255,N_309,N_160);
nor U1256 (N_1256,N_634,N_293);
or U1257 (N_1257,N_440,N_317);
and U1258 (N_1258,N_433,N_120);
and U1259 (N_1259,N_369,N_248);
nand U1260 (N_1260,N_172,N_515);
nor U1261 (N_1261,N_576,N_256);
nor U1262 (N_1262,N_78,N_346);
nor U1263 (N_1263,N_396,N_588);
or U1264 (N_1264,N_65,N_376);
nand U1265 (N_1265,N_282,N_67);
or U1266 (N_1266,N_204,N_227);
or U1267 (N_1267,N_520,N_265);
and U1268 (N_1268,N_688,N_748);
or U1269 (N_1269,N_205,N_130);
or U1270 (N_1270,N_166,N_283);
and U1271 (N_1271,N_315,N_484);
and U1272 (N_1272,N_44,N_451);
nor U1273 (N_1273,N_135,N_89);
nor U1274 (N_1274,N_668,N_539);
or U1275 (N_1275,N_585,N_411);
or U1276 (N_1276,N_525,N_117);
or U1277 (N_1277,N_258,N_332);
xor U1278 (N_1278,N_380,N_626);
and U1279 (N_1279,N_45,N_190);
or U1280 (N_1280,N_154,N_584);
or U1281 (N_1281,N_135,N_272);
and U1282 (N_1282,N_76,N_463);
nor U1283 (N_1283,N_140,N_492);
nand U1284 (N_1284,N_363,N_691);
xnor U1285 (N_1285,N_592,N_383);
nor U1286 (N_1286,N_695,N_680);
nor U1287 (N_1287,N_470,N_743);
xnor U1288 (N_1288,N_101,N_536);
xor U1289 (N_1289,N_430,N_532);
and U1290 (N_1290,N_505,N_216);
and U1291 (N_1291,N_491,N_652);
nor U1292 (N_1292,N_518,N_133);
and U1293 (N_1293,N_264,N_74);
xnor U1294 (N_1294,N_35,N_145);
nor U1295 (N_1295,N_524,N_691);
nand U1296 (N_1296,N_124,N_364);
nor U1297 (N_1297,N_579,N_642);
nand U1298 (N_1298,N_176,N_501);
xnor U1299 (N_1299,N_86,N_620);
nor U1300 (N_1300,N_474,N_62);
or U1301 (N_1301,N_543,N_358);
and U1302 (N_1302,N_498,N_642);
and U1303 (N_1303,N_309,N_731);
nand U1304 (N_1304,N_470,N_459);
or U1305 (N_1305,N_205,N_598);
nand U1306 (N_1306,N_216,N_23);
nor U1307 (N_1307,N_115,N_667);
and U1308 (N_1308,N_151,N_690);
or U1309 (N_1309,N_234,N_548);
nor U1310 (N_1310,N_185,N_657);
and U1311 (N_1311,N_206,N_249);
xnor U1312 (N_1312,N_749,N_268);
nand U1313 (N_1313,N_350,N_409);
and U1314 (N_1314,N_147,N_640);
xor U1315 (N_1315,N_617,N_226);
nand U1316 (N_1316,N_278,N_550);
or U1317 (N_1317,N_105,N_366);
nor U1318 (N_1318,N_158,N_477);
or U1319 (N_1319,N_400,N_453);
nor U1320 (N_1320,N_114,N_227);
nand U1321 (N_1321,N_480,N_186);
and U1322 (N_1322,N_102,N_658);
nor U1323 (N_1323,N_451,N_610);
or U1324 (N_1324,N_178,N_365);
and U1325 (N_1325,N_664,N_487);
and U1326 (N_1326,N_411,N_525);
nand U1327 (N_1327,N_607,N_138);
nor U1328 (N_1328,N_687,N_525);
xnor U1329 (N_1329,N_528,N_109);
and U1330 (N_1330,N_119,N_237);
or U1331 (N_1331,N_672,N_274);
xnor U1332 (N_1332,N_115,N_311);
nor U1333 (N_1333,N_196,N_579);
nor U1334 (N_1334,N_609,N_2);
and U1335 (N_1335,N_377,N_145);
and U1336 (N_1336,N_252,N_503);
and U1337 (N_1337,N_632,N_76);
nand U1338 (N_1338,N_644,N_158);
xor U1339 (N_1339,N_83,N_216);
or U1340 (N_1340,N_415,N_169);
xnor U1341 (N_1341,N_382,N_555);
or U1342 (N_1342,N_397,N_12);
nor U1343 (N_1343,N_624,N_724);
and U1344 (N_1344,N_17,N_119);
nand U1345 (N_1345,N_242,N_303);
xnor U1346 (N_1346,N_444,N_10);
and U1347 (N_1347,N_405,N_694);
or U1348 (N_1348,N_403,N_266);
xor U1349 (N_1349,N_463,N_335);
nand U1350 (N_1350,N_276,N_445);
and U1351 (N_1351,N_421,N_711);
nand U1352 (N_1352,N_422,N_387);
xnor U1353 (N_1353,N_511,N_278);
or U1354 (N_1354,N_71,N_428);
nand U1355 (N_1355,N_592,N_349);
and U1356 (N_1356,N_610,N_691);
xor U1357 (N_1357,N_332,N_226);
or U1358 (N_1358,N_24,N_142);
nand U1359 (N_1359,N_407,N_564);
xor U1360 (N_1360,N_329,N_365);
nor U1361 (N_1361,N_111,N_362);
or U1362 (N_1362,N_89,N_170);
xor U1363 (N_1363,N_108,N_88);
nor U1364 (N_1364,N_385,N_239);
nand U1365 (N_1365,N_256,N_325);
nor U1366 (N_1366,N_327,N_294);
nand U1367 (N_1367,N_467,N_511);
or U1368 (N_1368,N_32,N_60);
nor U1369 (N_1369,N_697,N_318);
and U1370 (N_1370,N_315,N_530);
nor U1371 (N_1371,N_670,N_512);
xor U1372 (N_1372,N_357,N_548);
nor U1373 (N_1373,N_535,N_349);
xor U1374 (N_1374,N_633,N_747);
and U1375 (N_1375,N_657,N_173);
nand U1376 (N_1376,N_735,N_484);
or U1377 (N_1377,N_64,N_683);
nor U1378 (N_1378,N_288,N_64);
nor U1379 (N_1379,N_107,N_367);
nor U1380 (N_1380,N_404,N_389);
nand U1381 (N_1381,N_629,N_405);
or U1382 (N_1382,N_228,N_311);
nand U1383 (N_1383,N_486,N_453);
xnor U1384 (N_1384,N_181,N_91);
and U1385 (N_1385,N_131,N_675);
or U1386 (N_1386,N_463,N_433);
xnor U1387 (N_1387,N_97,N_424);
or U1388 (N_1388,N_484,N_197);
or U1389 (N_1389,N_523,N_701);
nand U1390 (N_1390,N_15,N_663);
nor U1391 (N_1391,N_4,N_89);
nand U1392 (N_1392,N_491,N_586);
nand U1393 (N_1393,N_371,N_711);
nand U1394 (N_1394,N_719,N_702);
xor U1395 (N_1395,N_525,N_274);
xnor U1396 (N_1396,N_731,N_415);
xor U1397 (N_1397,N_91,N_49);
xnor U1398 (N_1398,N_170,N_372);
nor U1399 (N_1399,N_93,N_546);
and U1400 (N_1400,N_738,N_364);
and U1401 (N_1401,N_549,N_512);
xor U1402 (N_1402,N_444,N_57);
and U1403 (N_1403,N_680,N_673);
nand U1404 (N_1404,N_220,N_270);
or U1405 (N_1405,N_213,N_597);
nor U1406 (N_1406,N_475,N_739);
and U1407 (N_1407,N_120,N_351);
nor U1408 (N_1408,N_193,N_420);
xor U1409 (N_1409,N_363,N_321);
nand U1410 (N_1410,N_432,N_613);
and U1411 (N_1411,N_93,N_678);
or U1412 (N_1412,N_557,N_340);
nand U1413 (N_1413,N_15,N_449);
xor U1414 (N_1414,N_151,N_570);
xor U1415 (N_1415,N_642,N_540);
or U1416 (N_1416,N_30,N_149);
or U1417 (N_1417,N_416,N_259);
and U1418 (N_1418,N_271,N_212);
nand U1419 (N_1419,N_405,N_141);
nand U1420 (N_1420,N_240,N_440);
nand U1421 (N_1421,N_523,N_322);
nor U1422 (N_1422,N_484,N_311);
and U1423 (N_1423,N_235,N_700);
or U1424 (N_1424,N_306,N_198);
xor U1425 (N_1425,N_254,N_85);
and U1426 (N_1426,N_488,N_634);
nand U1427 (N_1427,N_410,N_252);
nand U1428 (N_1428,N_501,N_550);
nor U1429 (N_1429,N_709,N_590);
nand U1430 (N_1430,N_354,N_538);
xnor U1431 (N_1431,N_418,N_187);
or U1432 (N_1432,N_728,N_692);
xor U1433 (N_1433,N_342,N_19);
or U1434 (N_1434,N_668,N_715);
or U1435 (N_1435,N_409,N_38);
nor U1436 (N_1436,N_290,N_706);
and U1437 (N_1437,N_239,N_526);
nand U1438 (N_1438,N_405,N_93);
or U1439 (N_1439,N_567,N_273);
or U1440 (N_1440,N_736,N_711);
nand U1441 (N_1441,N_83,N_747);
nor U1442 (N_1442,N_347,N_600);
and U1443 (N_1443,N_62,N_308);
and U1444 (N_1444,N_223,N_152);
nand U1445 (N_1445,N_324,N_218);
nand U1446 (N_1446,N_709,N_699);
and U1447 (N_1447,N_678,N_112);
nor U1448 (N_1448,N_701,N_362);
xor U1449 (N_1449,N_80,N_561);
nand U1450 (N_1450,N_373,N_81);
nand U1451 (N_1451,N_303,N_668);
nand U1452 (N_1452,N_670,N_495);
xnor U1453 (N_1453,N_359,N_271);
xnor U1454 (N_1454,N_50,N_173);
nand U1455 (N_1455,N_503,N_711);
nand U1456 (N_1456,N_740,N_608);
nand U1457 (N_1457,N_459,N_588);
or U1458 (N_1458,N_447,N_511);
and U1459 (N_1459,N_11,N_585);
nor U1460 (N_1460,N_202,N_375);
xnor U1461 (N_1461,N_722,N_21);
xor U1462 (N_1462,N_720,N_325);
or U1463 (N_1463,N_358,N_126);
xnor U1464 (N_1464,N_727,N_123);
nor U1465 (N_1465,N_365,N_455);
and U1466 (N_1466,N_170,N_108);
nand U1467 (N_1467,N_702,N_0);
nand U1468 (N_1468,N_547,N_220);
nand U1469 (N_1469,N_718,N_524);
or U1470 (N_1470,N_99,N_285);
or U1471 (N_1471,N_68,N_535);
and U1472 (N_1472,N_690,N_547);
nand U1473 (N_1473,N_612,N_615);
or U1474 (N_1474,N_175,N_179);
xor U1475 (N_1475,N_316,N_709);
or U1476 (N_1476,N_18,N_594);
nand U1477 (N_1477,N_525,N_297);
and U1478 (N_1478,N_85,N_570);
nor U1479 (N_1479,N_698,N_188);
nand U1480 (N_1480,N_456,N_434);
xor U1481 (N_1481,N_243,N_183);
or U1482 (N_1482,N_452,N_323);
and U1483 (N_1483,N_366,N_633);
xnor U1484 (N_1484,N_273,N_697);
and U1485 (N_1485,N_407,N_629);
nand U1486 (N_1486,N_732,N_291);
xnor U1487 (N_1487,N_642,N_69);
or U1488 (N_1488,N_655,N_516);
xnor U1489 (N_1489,N_80,N_567);
and U1490 (N_1490,N_328,N_654);
or U1491 (N_1491,N_460,N_162);
xnor U1492 (N_1492,N_513,N_566);
nor U1493 (N_1493,N_640,N_25);
and U1494 (N_1494,N_196,N_435);
nor U1495 (N_1495,N_122,N_571);
xnor U1496 (N_1496,N_401,N_127);
nor U1497 (N_1497,N_481,N_328);
or U1498 (N_1498,N_107,N_84);
or U1499 (N_1499,N_237,N_0);
nor U1500 (N_1500,N_990,N_762);
and U1501 (N_1501,N_954,N_1051);
and U1502 (N_1502,N_1323,N_831);
nor U1503 (N_1503,N_1476,N_1057);
nand U1504 (N_1504,N_1473,N_1143);
or U1505 (N_1505,N_1201,N_1089);
and U1506 (N_1506,N_1156,N_1078);
xnor U1507 (N_1507,N_1029,N_1064);
xor U1508 (N_1508,N_1460,N_1387);
xor U1509 (N_1509,N_952,N_1413);
xnor U1510 (N_1510,N_1260,N_1146);
nand U1511 (N_1511,N_1025,N_785);
nand U1512 (N_1512,N_1477,N_889);
nand U1513 (N_1513,N_1242,N_801);
or U1514 (N_1514,N_783,N_1395);
nor U1515 (N_1515,N_977,N_764);
and U1516 (N_1516,N_828,N_886);
or U1517 (N_1517,N_1498,N_1044);
xnor U1518 (N_1518,N_1152,N_1119);
and U1519 (N_1519,N_837,N_1141);
nor U1520 (N_1520,N_765,N_971);
and U1521 (N_1521,N_923,N_1104);
nand U1522 (N_1522,N_1014,N_798);
xnor U1523 (N_1523,N_998,N_888);
nor U1524 (N_1524,N_880,N_1344);
xnor U1525 (N_1525,N_1045,N_1332);
nor U1526 (N_1526,N_1264,N_962);
or U1527 (N_1527,N_942,N_1422);
nor U1528 (N_1528,N_1324,N_984);
xor U1529 (N_1529,N_1243,N_985);
xor U1530 (N_1530,N_915,N_1094);
nand U1531 (N_1531,N_1191,N_1306);
or U1532 (N_1532,N_814,N_1273);
and U1533 (N_1533,N_1289,N_1252);
or U1534 (N_1534,N_1442,N_768);
and U1535 (N_1535,N_1147,N_938);
or U1536 (N_1536,N_1174,N_1012);
and U1537 (N_1537,N_1457,N_1354);
or U1538 (N_1538,N_779,N_1463);
nand U1539 (N_1539,N_909,N_997);
or U1540 (N_1540,N_1282,N_1231);
nand U1541 (N_1541,N_1056,N_918);
nor U1542 (N_1542,N_1085,N_1298);
or U1543 (N_1543,N_1401,N_1224);
xnor U1544 (N_1544,N_1479,N_944);
nand U1545 (N_1545,N_1164,N_1493);
nor U1546 (N_1546,N_1385,N_1000);
xnor U1547 (N_1547,N_1368,N_1420);
nand U1548 (N_1548,N_898,N_838);
and U1549 (N_1549,N_1386,N_817);
nor U1550 (N_1550,N_910,N_1378);
nand U1551 (N_1551,N_849,N_1337);
nand U1552 (N_1552,N_1482,N_1183);
or U1553 (N_1553,N_1226,N_1281);
xnor U1554 (N_1554,N_1375,N_948);
nand U1555 (N_1555,N_919,N_1421);
xor U1556 (N_1556,N_966,N_782);
nor U1557 (N_1557,N_1053,N_772);
nand U1558 (N_1558,N_1061,N_1123);
nor U1559 (N_1559,N_921,N_1038);
or U1560 (N_1560,N_1023,N_867);
or U1561 (N_1561,N_896,N_1266);
xor U1562 (N_1562,N_1039,N_1329);
xnor U1563 (N_1563,N_1139,N_1162);
xnor U1564 (N_1564,N_1200,N_1022);
or U1565 (N_1565,N_1275,N_787);
nand U1566 (N_1566,N_1178,N_1322);
nor U1567 (N_1567,N_1219,N_1336);
xnor U1568 (N_1568,N_1013,N_1373);
xnor U1569 (N_1569,N_857,N_820);
and U1570 (N_1570,N_1213,N_790);
or U1571 (N_1571,N_963,N_974);
nand U1572 (N_1572,N_1155,N_906);
nand U1573 (N_1573,N_975,N_1445);
nand U1574 (N_1574,N_1090,N_1112);
xnor U1575 (N_1575,N_1163,N_970);
xnor U1576 (N_1576,N_1254,N_1189);
xor U1577 (N_1577,N_1425,N_1220);
and U1578 (N_1578,N_1389,N_881);
and U1579 (N_1579,N_839,N_1233);
xnor U1580 (N_1580,N_1302,N_1443);
or U1581 (N_1581,N_1048,N_850);
or U1582 (N_1582,N_1449,N_1431);
nor U1583 (N_1583,N_1184,N_1295);
and U1584 (N_1584,N_1232,N_1228);
or U1585 (N_1585,N_1384,N_1127);
xnor U1586 (N_1586,N_1440,N_1113);
nand U1587 (N_1587,N_874,N_1392);
xnor U1588 (N_1588,N_928,N_1317);
xnor U1589 (N_1589,N_1204,N_810);
or U1590 (N_1590,N_1497,N_1483);
nor U1591 (N_1591,N_1081,N_1432);
xnor U1592 (N_1592,N_1492,N_846);
or U1593 (N_1593,N_1453,N_1403);
nand U1594 (N_1594,N_879,N_1303);
and U1595 (N_1595,N_1372,N_1157);
xnor U1596 (N_1596,N_1076,N_1080);
and U1597 (N_1597,N_1304,N_1125);
xnor U1598 (N_1598,N_951,N_1364);
and U1599 (N_1599,N_781,N_949);
and U1600 (N_1600,N_1207,N_802);
nor U1601 (N_1601,N_1217,N_1287);
xnor U1602 (N_1602,N_1446,N_822);
xnor U1603 (N_1603,N_860,N_1404);
or U1604 (N_1604,N_1103,N_1390);
and U1605 (N_1605,N_1283,N_856);
nor U1606 (N_1606,N_1426,N_755);
xor U1607 (N_1607,N_1280,N_1454);
xnor U1608 (N_1608,N_1314,N_758);
nand U1609 (N_1609,N_1239,N_1316);
nand U1610 (N_1610,N_973,N_893);
nor U1611 (N_1611,N_1101,N_1247);
nor U1612 (N_1612,N_1333,N_979);
nor U1613 (N_1613,N_1459,N_826);
and U1614 (N_1614,N_1236,N_1185);
nand U1615 (N_1615,N_1255,N_1009);
nor U1616 (N_1616,N_812,N_1108);
nand U1617 (N_1617,N_1414,N_1248);
nand U1618 (N_1618,N_961,N_1307);
nand U1619 (N_1619,N_996,N_903);
and U1620 (N_1620,N_1394,N_958);
or U1621 (N_1621,N_892,N_1257);
nand U1622 (N_1622,N_760,N_1343);
xnor U1623 (N_1623,N_1409,N_1251);
xor U1624 (N_1624,N_847,N_1376);
and U1625 (N_1625,N_870,N_1202);
xor U1626 (N_1626,N_1002,N_1391);
or U1627 (N_1627,N_1423,N_1424);
xor U1628 (N_1628,N_929,N_967);
and U1629 (N_1629,N_993,N_1340);
nor U1630 (N_1630,N_836,N_1030);
or U1631 (N_1631,N_815,N_1438);
or U1632 (N_1632,N_1270,N_1106);
nor U1633 (N_1633,N_1010,N_1196);
nand U1634 (N_1634,N_1465,N_1097);
or U1635 (N_1635,N_1172,N_1145);
xor U1636 (N_1636,N_941,N_968);
and U1637 (N_1637,N_1227,N_1008);
xor U1638 (N_1638,N_1182,N_752);
and U1639 (N_1639,N_1456,N_1176);
nand U1640 (N_1640,N_953,N_1109);
nor U1641 (N_1641,N_763,N_862);
xnor U1642 (N_1642,N_885,N_1096);
and U1643 (N_1643,N_1494,N_1334);
nand U1644 (N_1644,N_854,N_1429);
or U1645 (N_1645,N_1199,N_1487);
nor U1646 (N_1646,N_805,N_1111);
or U1647 (N_1647,N_1007,N_1190);
nand U1648 (N_1648,N_1297,N_827);
nand U1649 (N_1649,N_1188,N_1475);
nand U1650 (N_1650,N_1259,N_1070);
nor U1651 (N_1651,N_1117,N_859);
nor U1652 (N_1652,N_994,N_1160);
and U1653 (N_1653,N_873,N_1165);
nand U1654 (N_1654,N_940,N_1077);
xnor U1655 (N_1655,N_1293,N_1100);
or U1656 (N_1656,N_1458,N_1299);
or U1657 (N_1657,N_842,N_806);
xnor U1658 (N_1658,N_1073,N_1168);
or U1659 (N_1659,N_1462,N_1399);
or U1660 (N_1660,N_1320,N_1218);
nor U1661 (N_1661,N_1159,N_1262);
xnor U1662 (N_1662,N_767,N_1197);
or U1663 (N_1663,N_947,N_1427);
nand U1664 (N_1664,N_1355,N_1467);
nor U1665 (N_1665,N_982,N_1279);
xnor U1666 (N_1666,N_1338,N_1120);
and U1667 (N_1667,N_1102,N_1330);
nand U1668 (N_1668,N_1067,N_803);
nor U1669 (N_1669,N_1206,N_1003);
and U1670 (N_1670,N_845,N_991);
nand U1671 (N_1671,N_916,N_1328);
or U1672 (N_1672,N_1065,N_1210);
nand U1673 (N_1673,N_816,N_1407);
xnor U1674 (N_1674,N_1169,N_1198);
and U1675 (N_1675,N_1122,N_808);
and U1676 (N_1676,N_1049,N_1031);
nor U1677 (N_1677,N_972,N_786);
nor U1678 (N_1678,N_858,N_1194);
and U1679 (N_1679,N_784,N_775);
nand U1680 (N_1680,N_1411,N_1063);
and U1681 (N_1681,N_1419,N_1181);
and U1682 (N_1682,N_1211,N_1474);
nand U1683 (N_1683,N_1225,N_1140);
xnor U1684 (N_1684,N_1246,N_1229);
nand U1685 (N_1685,N_1367,N_1265);
nand U1686 (N_1686,N_1398,N_1291);
and U1687 (N_1687,N_1046,N_965);
and U1688 (N_1688,N_936,N_1471);
nand U1689 (N_1689,N_920,N_1059);
xnor U1690 (N_1690,N_829,N_756);
and U1691 (N_1691,N_912,N_876);
and U1692 (N_1692,N_848,N_861);
nand U1693 (N_1693,N_937,N_1092);
xnor U1694 (N_1694,N_1245,N_1312);
or U1695 (N_1695,N_1105,N_1091);
nor U1696 (N_1696,N_1310,N_1305);
and U1697 (N_1697,N_960,N_1033);
nand U1698 (N_1698,N_1074,N_871);
or U1699 (N_1699,N_1346,N_935);
nand U1700 (N_1700,N_863,N_789);
nand U1701 (N_1701,N_1035,N_1491);
nand U1702 (N_1702,N_1488,N_1380);
nand U1703 (N_1703,N_1034,N_943);
nor U1704 (N_1704,N_1341,N_1167);
xor U1705 (N_1705,N_1240,N_1216);
and U1706 (N_1706,N_811,N_1018);
nand U1707 (N_1707,N_1235,N_791);
nor U1708 (N_1708,N_1315,N_1087);
or U1709 (N_1709,N_771,N_1495);
xor U1710 (N_1710,N_1365,N_804);
nand U1711 (N_1711,N_1084,N_1026);
nor U1712 (N_1712,N_1138,N_753);
xnor U1713 (N_1713,N_934,N_1161);
nand U1714 (N_1714,N_1472,N_1441);
nor U1715 (N_1715,N_1203,N_1261);
nand U1716 (N_1716,N_1144,N_1041);
and U1717 (N_1717,N_794,N_999);
nor U1718 (N_1718,N_884,N_891);
nand U1719 (N_1719,N_1052,N_1377);
or U1720 (N_1720,N_1093,N_1208);
or U1721 (N_1721,N_1321,N_1437);
xnor U1722 (N_1722,N_883,N_1110);
and U1723 (N_1723,N_1086,N_1170);
or U1724 (N_1724,N_1179,N_877);
xnor U1725 (N_1725,N_957,N_924);
nand U1726 (N_1726,N_946,N_1433);
and U1727 (N_1727,N_1095,N_1195);
and U1728 (N_1728,N_1402,N_926);
nand U1729 (N_1729,N_1418,N_1017);
nand U1730 (N_1730,N_1166,N_1066);
or U1731 (N_1731,N_1047,N_1277);
nor U1732 (N_1732,N_841,N_989);
xnor U1733 (N_1733,N_1024,N_1050);
xnor U1734 (N_1734,N_986,N_778);
or U1735 (N_1735,N_757,N_1192);
xnor U1736 (N_1736,N_799,N_1158);
nor U1737 (N_1737,N_955,N_927);
nor U1738 (N_1738,N_1062,N_1249);
xnor U1739 (N_1739,N_1128,N_1335);
nand U1740 (N_1740,N_1301,N_1331);
and U1741 (N_1741,N_1371,N_907);
nand U1742 (N_1742,N_1083,N_1326);
or U1743 (N_1743,N_1186,N_1481);
or U1744 (N_1744,N_875,N_1461);
and U1745 (N_1745,N_1374,N_853);
nor U1746 (N_1746,N_1071,N_1075);
and U1747 (N_1747,N_1244,N_1388);
xor U1748 (N_1748,N_932,N_1011);
and U1749 (N_1749,N_980,N_1148);
xor U1750 (N_1750,N_956,N_1253);
nand U1751 (N_1751,N_895,N_844);
nor U1752 (N_1752,N_978,N_1132);
nand U1753 (N_1753,N_1400,N_1116);
nor U1754 (N_1754,N_1366,N_914);
or U1755 (N_1755,N_1339,N_823);
and U1756 (N_1756,N_1484,N_922);
xnor U1757 (N_1757,N_1134,N_761);
nand U1758 (N_1758,N_1327,N_1153);
xor U1759 (N_1759,N_1383,N_866);
and U1760 (N_1760,N_1359,N_1450);
nand U1761 (N_1761,N_800,N_1319);
or U1762 (N_1762,N_899,N_1114);
or U1763 (N_1763,N_807,N_1350);
nor U1764 (N_1764,N_988,N_1032);
xnor U1765 (N_1765,N_1250,N_1434);
nor U1766 (N_1766,N_1363,N_769);
and U1767 (N_1767,N_911,N_1269);
or U1768 (N_1768,N_1223,N_1300);
and U1769 (N_1769,N_1318,N_1175);
and U1770 (N_1770,N_777,N_793);
and U1771 (N_1771,N_865,N_1271);
or U1772 (N_1772,N_843,N_825);
nand U1773 (N_1773,N_1027,N_933);
or U1774 (N_1774,N_950,N_1180);
and U1775 (N_1775,N_809,N_797);
or U1776 (N_1776,N_1069,N_887);
xnor U1777 (N_1777,N_913,N_1309);
nand U1778 (N_1778,N_1313,N_905);
nand U1779 (N_1779,N_1130,N_1215);
xor U1780 (N_1780,N_1238,N_1360);
and U1781 (N_1781,N_1149,N_1177);
and U1782 (N_1782,N_1358,N_1209);
or U1783 (N_1783,N_1499,N_1263);
nand U1784 (N_1784,N_1005,N_976);
nor U1785 (N_1785,N_1016,N_1370);
or U1786 (N_1786,N_931,N_824);
nor U1787 (N_1787,N_1396,N_1278);
nor U1788 (N_1788,N_1288,N_1221);
xor U1789 (N_1789,N_869,N_1382);
nor U1790 (N_1790,N_1468,N_1131);
nor U1791 (N_1791,N_1020,N_1121);
nand U1792 (N_1792,N_1415,N_1342);
or U1793 (N_1793,N_1072,N_773);
nand U1794 (N_1794,N_819,N_1410);
nand U1795 (N_1795,N_1036,N_1444);
or U1796 (N_1796,N_900,N_1436);
or U1797 (N_1797,N_864,N_1469);
xor U1798 (N_1798,N_1369,N_901);
nand U1799 (N_1799,N_1021,N_818);
nor U1800 (N_1800,N_1448,N_1397);
xnor U1801 (N_1801,N_1040,N_868);
or U1802 (N_1802,N_983,N_1489);
xor U1803 (N_1803,N_1060,N_1362);
nand U1804 (N_1804,N_1126,N_1272);
nor U1805 (N_1805,N_788,N_1361);
xnor U1806 (N_1806,N_969,N_1470);
and U1807 (N_1807,N_1054,N_832);
nor U1808 (N_1808,N_1296,N_1439);
nand U1809 (N_1809,N_1478,N_796);
nor U1810 (N_1810,N_1079,N_834);
xor U1811 (N_1811,N_1351,N_1004);
or U1812 (N_1812,N_894,N_1258);
nand U1813 (N_1813,N_1349,N_1311);
xor U1814 (N_1814,N_1345,N_1435);
xnor U1815 (N_1815,N_1135,N_1006);
nand U1816 (N_1816,N_917,N_1136);
nand U1817 (N_1817,N_1416,N_1151);
nand U1818 (N_1818,N_1124,N_1118);
nand U1819 (N_1819,N_1058,N_964);
and U1820 (N_1820,N_1408,N_1274);
nor U1821 (N_1821,N_1082,N_766);
xnor U1822 (N_1822,N_1212,N_1356);
nor U1823 (N_1823,N_1357,N_751);
nor U1824 (N_1824,N_821,N_840);
nor U1825 (N_1825,N_1379,N_1430);
xor U1826 (N_1826,N_1285,N_1171);
nor U1827 (N_1827,N_1055,N_1001);
xor U1828 (N_1828,N_1286,N_776);
nand U1829 (N_1829,N_1268,N_1193);
and U1830 (N_1830,N_1486,N_1150);
or U1831 (N_1831,N_1037,N_855);
or U1832 (N_1832,N_813,N_1405);
xor U1833 (N_1833,N_890,N_1256);
nor U1834 (N_1834,N_1417,N_1042);
nor U1835 (N_1835,N_882,N_750);
or U1836 (N_1836,N_1237,N_1412);
nand U1837 (N_1837,N_1205,N_959);
nor U1838 (N_1838,N_1241,N_878);
nor U1839 (N_1839,N_897,N_1137);
nand U1840 (N_1840,N_1019,N_904);
or U1841 (N_1841,N_1451,N_1276);
and U1842 (N_1842,N_1043,N_851);
or U1843 (N_1843,N_1267,N_1222);
nand U1844 (N_1844,N_1325,N_1455);
and U1845 (N_1845,N_992,N_1348);
xnor U1846 (N_1846,N_1347,N_1290);
xor U1847 (N_1847,N_1353,N_1187);
or U1848 (N_1848,N_835,N_1015);
nor U1849 (N_1849,N_1308,N_908);
nor U1850 (N_1850,N_770,N_833);
or U1851 (N_1851,N_1098,N_1294);
and U1852 (N_1852,N_792,N_1466);
xor U1853 (N_1853,N_759,N_1406);
and U1854 (N_1854,N_981,N_1393);
xnor U1855 (N_1855,N_1485,N_902);
nor U1856 (N_1856,N_1214,N_930);
nand U1857 (N_1857,N_795,N_1234);
nand U1858 (N_1858,N_1173,N_1068);
xor U1859 (N_1859,N_780,N_1480);
nor U1860 (N_1860,N_1292,N_1154);
xnor U1861 (N_1861,N_754,N_774);
nor U1862 (N_1862,N_1352,N_925);
nand U1863 (N_1863,N_1284,N_1381);
xnor U1864 (N_1864,N_945,N_1129);
or U1865 (N_1865,N_1447,N_1452);
nor U1866 (N_1866,N_1230,N_987);
or U1867 (N_1867,N_1028,N_1464);
xnor U1868 (N_1868,N_1496,N_1133);
nor U1869 (N_1869,N_995,N_1428);
nand U1870 (N_1870,N_1115,N_830);
and U1871 (N_1871,N_1107,N_872);
or U1872 (N_1872,N_1099,N_1088);
nor U1873 (N_1873,N_852,N_1490);
and U1874 (N_1874,N_939,N_1142);
nor U1875 (N_1875,N_1206,N_1231);
or U1876 (N_1876,N_1283,N_1085);
xnor U1877 (N_1877,N_1036,N_1407);
or U1878 (N_1878,N_946,N_1153);
or U1879 (N_1879,N_977,N_1238);
xnor U1880 (N_1880,N_793,N_1202);
nor U1881 (N_1881,N_1057,N_903);
and U1882 (N_1882,N_899,N_895);
xnor U1883 (N_1883,N_1177,N_1210);
nor U1884 (N_1884,N_790,N_963);
or U1885 (N_1885,N_1499,N_1385);
or U1886 (N_1886,N_1103,N_978);
and U1887 (N_1887,N_1422,N_1441);
xnor U1888 (N_1888,N_899,N_1392);
nand U1889 (N_1889,N_902,N_819);
and U1890 (N_1890,N_1038,N_822);
or U1891 (N_1891,N_831,N_1495);
nand U1892 (N_1892,N_1304,N_1225);
nand U1893 (N_1893,N_1247,N_1307);
or U1894 (N_1894,N_1330,N_847);
xor U1895 (N_1895,N_855,N_1461);
and U1896 (N_1896,N_974,N_905);
nand U1897 (N_1897,N_1475,N_1027);
and U1898 (N_1898,N_979,N_828);
or U1899 (N_1899,N_1178,N_901);
or U1900 (N_1900,N_1059,N_1464);
nor U1901 (N_1901,N_1476,N_1362);
or U1902 (N_1902,N_1116,N_796);
or U1903 (N_1903,N_919,N_955);
xnor U1904 (N_1904,N_1189,N_1075);
nor U1905 (N_1905,N_1365,N_1479);
or U1906 (N_1906,N_842,N_1186);
or U1907 (N_1907,N_1230,N_1479);
and U1908 (N_1908,N_1211,N_1172);
nand U1909 (N_1909,N_1259,N_1453);
and U1910 (N_1910,N_1236,N_980);
or U1911 (N_1911,N_813,N_1205);
xnor U1912 (N_1912,N_837,N_1133);
xor U1913 (N_1913,N_776,N_952);
nand U1914 (N_1914,N_1396,N_1257);
nand U1915 (N_1915,N_821,N_1198);
or U1916 (N_1916,N_853,N_1090);
nor U1917 (N_1917,N_1447,N_1317);
nor U1918 (N_1918,N_918,N_1238);
nand U1919 (N_1919,N_790,N_1198);
nor U1920 (N_1920,N_955,N_767);
nand U1921 (N_1921,N_1183,N_1185);
xor U1922 (N_1922,N_825,N_1007);
nand U1923 (N_1923,N_897,N_964);
nor U1924 (N_1924,N_975,N_1110);
and U1925 (N_1925,N_1420,N_1389);
and U1926 (N_1926,N_1123,N_1338);
xnor U1927 (N_1927,N_768,N_1203);
nand U1928 (N_1928,N_806,N_1085);
or U1929 (N_1929,N_1357,N_972);
nand U1930 (N_1930,N_1232,N_965);
or U1931 (N_1931,N_1026,N_1301);
and U1932 (N_1932,N_1126,N_1046);
and U1933 (N_1933,N_1107,N_1400);
or U1934 (N_1934,N_833,N_1360);
or U1935 (N_1935,N_796,N_935);
or U1936 (N_1936,N_1178,N_1079);
nor U1937 (N_1937,N_1455,N_1429);
nand U1938 (N_1938,N_991,N_1387);
nand U1939 (N_1939,N_1448,N_934);
or U1940 (N_1940,N_1210,N_1151);
nand U1941 (N_1941,N_1201,N_839);
or U1942 (N_1942,N_1355,N_897);
or U1943 (N_1943,N_845,N_1194);
or U1944 (N_1944,N_1257,N_1123);
nand U1945 (N_1945,N_1106,N_1145);
nor U1946 (N_1946,N_1128,N_1339);
nor U1947 (N_1947,N_909,N_1257);
or U1948 (N_1948,N_1264,N_1058);
xnor U1949 (N_1949,N_1158,N_1084);
or U1950 (N_1950,N_934,N_1105);
nand U1951 (N_1951,N_1470,N_1119);
nand U1952 (N_1952,N_1065,N_1103);
nand U1953 (N_1953,N_1190,N_1282);
or U1954 (N_1954,N_835,N_1232);
or U1955 (N_1955,N_1092,N_1236);
xor U1956 (N_1956,N_1238,N_1008);
nor U1957 (N_1957,N_1305,N_1421);
and U1958 (N_1958,N_1213,N_853);
nor U1959 (N_1959,N_909,N_1411);
nand U1960 (N_1960,N_1152,N_1386);
xor U1961 (N_1961,N_1423,N_1032);
nor U1962 (N_1962,N_1024,N_1476);
nor U1963 (N_1963,N_1233,N_1103);
and U1964 (N_1964,N_1278,N_1495);
or U1965 (N_1965,N_1043,N_1146);
and U1966 (N_1966,N_970,N_1004);
xor U1967 (N_1967,N_809,N_1085);
and U1968 (N_1968,N_1322,N_1144);
or U1969 (N_1969,N_890,N_1434);
nand U1970 (N_1970,N_887,N_816);
nand U1971 (N_1971,N_1196,N_950);
and U1972 (N_1972,N_1277,N_1174);
nand U1973 (N_1973,N_991,N_1391);
or U1974 (N_1974,N_1147,N_1458);
or U1975 (N_1975,N_1339,N_869);
nand U1976 (N_1976,N_1058,N_926);
nand U1977 (N_1977,N_955,N_1229);
xnor U1978 (N_1978,N_1299,N_1464);
or U1979 (N_1979,N_1389,N_918);
nand U1980 (N_1980,N_970,N_1077);
nor U1981 (N_1981,N_1413,N_912);
or U1982 (N_1982,N_1439,N_1376);
nor U1983 (N_1983,N_1375,N_970);
or U1984 (N_1984,N_1153,N_824);
and U1985 (N_1985,N_1328,N_1218);
and U1986 (N_1986,N_1404,N_1037);
nand U1987 (N_1987,N_1052,N_837);
nor U1988 (N_1988,N_1367,N_1462);
and U1989 (N_1989,N_874,N_930);
and U1990 (N_1990,N_1273,N_1062);
and U1991 (N_1991,N_1456,N_1028);
nor U1992 (N_1992,N_1127,N_995);
or U1993 (N_1993,N_1218,N_796);
nand U1994 (N_1994,N_1084,N_1495);
and U1995 (N_1995,N_1486,N_954);
nand U1996 (N_1996,N_1210,N_1300);
nand U1997 (N_1997,N_972,N_1295);
nor U1998 (N_1998,N_1490,N_990);
or U1999 (N_1999,N_1252,N_1384);
and U2000 (N_2000,N_1394,N_1260);
nor U2001 (N_2001,N_830,N_787);
or U2002 (N_2002,N_1256,N_829);
nand U2003 (N_2003,N_1059,N_1336);
and U2004 (N_2004,N_1020,N_1414);
or U2005 (N_2005,N_1198,N_909);
or U2006 (N_2006,N_1375,N_832);
nand U2007 (N_2007,N_1252,N_868);
nand U2008 (N_2008,N_1006,N_899);
nand U2009 (N_2009,N_1107,N_931);
nor U2010 (N_2010,N_1231,N_820);
nor U2011 (N_2011,N_912,N_1175);
and U2012 (N_2012,N_757,N_1473);
nor U2013 (N_2013,N_1000,N_1052);
xor U2014 (N_2014,N_1109,N_972);
and U2015 (N_2015,N_1373,N_1406);
and U2016 (N_2016,N_1224,N_1294);
or U2017 (N_2017,N_1246,N_964);
xor U2018 (N_2018,N_1207,N_1290);
or U2019 (N_2019,N_1253,N_1029);
xor U2020 (N_2020,N_1321,N_1165);
and U2021 (N_2021,N_1399,N_947);
and U2022 (N_2022,N_1367,N_1006);
or U2023 (N_2023,N_1120,N_1242);
nor U2024 (N_2024,N_1005,N_1223);
nand U2025 (N_2025,N_1400,N_1240);
and U2026 (N_2026,N_1377,N_1222);
nand U2027 (N_2027,N_1016,N_1457);
nor U2028 (N_2028,N_821,N_1056);
xnor U2029 (N_2029,N_1052,N_1178);
and U2030 (N_2030,N_1215,N_1069);
nand U2031 (N_2031,N_1254,N_1490);
nand U2032 (N_2032,N_1131,N_1272);
or U2033 (N_2033,N_949,N_1396);
and U2034 (N_2034,N_894,N_1243);
and U2035 (N_2035,N_841,N_1291);
and U2036 (N_2036,N_1258,N_1301);
and U2037 (N_2037,N_939,N_895);
nor U2038 (N_2038,N_1478,N_1378);
nand U2039 (N_2039,N_982,N_869);
nand U2040 (N_2040,N_1054,N_1393);
xnor U2041 (N_2041,N_882,N_1301);
nand U2042 (N_2042,N_846,N_763);
xor U2043 (N_2043,N_833,N_1416);
nor U2044 (N_2044,N_1043,N_1260);
or U2045 (N_2045,N_1328,N_1480);
xor U2046 (N_2046,N_1070,N_1255);
xnor U2047 (N_2047,N_1082,N_1295);
nand U2048 (N_2048,N_1335,N_1409);
nor U2049 (N_2049,N_1435,N_1004);
and U2050 (N_2050,N_1297,N_1381);
xnor U2051 (N_2051,N_873,N_1005);
xor U2052 (N_2052,N_996,N_924);
xor U2053 (N_2053,N_1465,N_1130);
or U2054 (N_2054,N_1153,N_1384);
nand U2055 (N_2055,N_1068,N_1143);
xnor U2056 (N_2056,N_1192,N_1282);
xor U2057 (N_2057,N_1016,N_1319);
nor U2058 (N_2058,N_1024,N_1382);
nand U2059 (N_2059,N_964,N_1492);
nor U2060 (N_2060,N_1374,N_1338);
nand U2061 (N_2061,N_1107,N_961);
or U2062 (N_2062,N_1399,N_783);
or U2063 (N_2063,N_1488,N_1430);
nor U2064 (N_2064,N_1232,N_1215);
nand U2065 (N_2065,N_1312,N_805);
xor U2066 (N_2066,N_1082,N_1072);
nor U2067 (N_2067,N_909,N_1079);
xor U2068 (N_2068,N_1211,N_953);
nor U2069 (N_2069,N_1177,N_1386);
nand U2070 (N_2070,N_1472,N_1031);
and U2071 (N_2071,N_1429,N_1435);
and U2072 (N_2072,N_955,N_1470);
and U2073 (N_2073,N_1037,N_1395);
xnor U2074 (N_2074,N_1130,N_766);
or U2075 (N_2075,N_1236,N_1016);
nand U2076 (N_2076,N_1402,N_1223);
nand U2077 (N_2077,N_1252,N_757);
or U2078 (N_2078,N_1040,N_950);
or U2079 (N_2079,N_895,N_978);
nand U2080 (N_2080,N_1323,N_816);
xor U2081 (N_2081,N_1139,N_1241);
xnor U2082 (N_2082,N_1305,N_1036);
xor U2083 (N_2083,N_1102,N_844);
xor U2084 (N_2084,N_984,N_835);
nand U2085 (N_2085,N_905,N_1345);
nand U2086 (N_2086,N_1099,N_1127);
and U2087 (N_2087,N_1336,N_886);
xnor U2088 (N_2088,N_1383,N_816);
nand U2089 (N_2089,N_1366,N_1439);
and U2090 (N_2090,N_855,N_1256);
or U2091 (N_2091,N_1324,N_1162);
nor U2092 (N_2092,N_1182,N_767);
nand U2093 (N_2093,N_1421,N_1139);
xor U2094 (N_2094,N_959,N_1067);
nand U2095 (N_2095,N_1429,N_852);
nor U2096 (N_2096,N_1377,N_849);
nor U2097 (N_2097,N_870,N_1042);
or U2098 (N_2098,N_1040,N_817);
xnor U2099 (N_2099,N_1390,N_934);
nor U2100 (N_2100,N_873,N_1013);
or U2101 (N_2101,N_1097,N_1269);
nor U2102 (N_2102,N_1192,N_1279);
xor U2103 (N_2103,N_1436,N_1337);
and U2104 (N_2104,N_1104,N_1442);
xor U2105 (N_2105,N_1103,N_994);
xnor U2106 (N_2106,N_1377,N_878);
or U2107 (N_2107,N_1361,N_1267);
xnor U2108 (N_2108,N_1158,N_1277);
nand U2109 (N_2109,N_828,N_764);
nor U2110 (N_2110,N_863,N_930);
nand U2111 (N_2111,N_818,N_896);
nor U2112 (N_2112,N_817,N_996);
nand U2113 (N_2113,N_1257,N_896);
and U2114 (N_2114,N_1334,N_924);
xor U2115 (N_2115,N_824,N_1244);
nand U2116 (N_2116,N_1025,N_816);
xnor U2117 (N_2117,N_1143,N_773);
xor U2118 (N_2118,N_1314,N_1173);
or U2119 (N_2119,N_793,N_1215);
nand U2120 (N_2120,N_1023,N_1107);
and U2121 (N_2121,N_961,N_1096);
and U2122 (N_2122,N_1234,N_1252);
and U2123 (N_2123,N_925,N_803);
or U2124 (N_2124,N_1321,N_925);
nor U2125 (N_2125,N_1440,N_981);
or U2126 (N_2126,N_1487,N_1404);
or U2127 (N_2127,N_1034,N_930);
nor U2128 (N_2128,N_1393,N_1026);
nor U2129 (N_2129,N_958,N_864);
and U2130 (N_2130,N_1104,N_898);
nand U2131 (N_2131,N_934,N_1180);
or U2132 (N_2132,N_978,N_1110);
and U2133 (N_2133,N_1041,N_1107);
and U2134 (N_2134,N_1209,N_1286);
xor U2135 (N_2135,N_1164,N_1183);
or U2136 (N_2136,N_827,N_1096);
xnor U2137 (N_2137,N_1199,N_973);
or U2138 (N_2138,N_845,N_1008);
nand U2139 (N_2139,N_907,N_1035);
nor U2140 (N_2140,N_1103,N_980);
and U2141 (N_2141,N_842,N_1047);
and U2142 (N_2142,N_1181,N_1472);
nor U2143 (N_2143,N_1109,N_1494);
and U2144 (N_2144,N_1403,N_1160);
nand U2145 (N_2145,N_1023,N_1252);
nor U2146 (N_2146,N_1398,N_1479);
nor U2147 (N_2147,N_1217,N_796);
or U2148 (N_2148,N_1438,N_897);
nor U2149 (N_2149,N_897,N_1359);
nor U2150 (N_2150,N_1169,N_1057);
nand U2151 (N_2151,N_885,N_1370);
or U2152 (N_2152,N_1344,N_776);
nand U2153 (N_2153,N_1105,N_1371);
or U2154 (N_2154,N_1032,N_1311);
and U2155 (N_2155,N_1335,N_789);
or U2156 (N_2156,N_1051,N_892);
nand U2157 (N_2157,N_890,N_1079);
nand U2158 (N_2158,N_1220,N_1296);
nor U2159 (N_2159,N_1399,N_875);
xor U2160 (N_2160,N_1025,N_1069);
nor U2161 (N_2161,N_896,N_1268);
nor U2162 (N_2162,N_844,N_1158);
or U2163 (N_2163,N_1113,N_1054);
xnor U2164 (N_2164,N_1112,N_1382);
nand U2165 (N_2165,N_1270,N_867);
nor U2166 (N_2166,N_1094,N_1011);
or U2167 (N_2167,N_1063,N_1401);
nor U2168 (N_2168,N_1411,N_869);
and U2169 (N_2169,N_973,N_1083);
nor U2170 (N_2170,N_1457,N_1305);
nor U2171 (N_2171,N_1476,N_862);
nor U2172 (N_2172,N_1318,N_866);
xor U2173 (N_2173,N_1364,N_803);
and U2174 (N_2174,N_1149,N_1459);
xor U2175 (N_2175,N_980,N_794);
and U2176 (N_2176,N_1494,N_1108);
and U2177 (N_2177,N_1406,N_1162);
nand U2178 (N_2178,N_1315,N_1023);
and U2179 (N_2179,N_790,N_1108);
nand U2180 (N_2180,N_952,N_1369);
nor U2181 (N_2181,N_1185,N_1497);
or U2182 (N_2182,N_1316,N_1043);
and U2183 (N_2183,N_993,N_1307);
or U2184 (N_2184,N_1119,N_1384);
nor U2185 (N_2185,N_1478,N_1203);
nand U2186 (N_2186,N_804,N_1013);
or U2187 (N_2187,N_1157,N_1032);
xor U2188 (N_2188,N_1462,N_1406);
nor U2189 (N_2189,N_994,N_1497);
and U2190 (N_2190,N_1105,N_1418);
xnor U2191 (N_2191,N_1294,N_1013);
nand U2192 (N_2192,N_1256,N_1106);
or U2193 (N_2193,N_1221,N_1363);
nand U2194 (N_2194,N_1104,N_1363);
and U2195 (N_2195,N_1441,N_808);
nand U2196 (N_2196,N_1165,N_1107);
xnor U2197 (N_2197,N_1371,N_836);
nand U2198 (N_2198,N_1258,N_1250);
and U2199 (N_2199,N_753,N_1310);
nand U2200 (N_2200,N_1445,N_1323);
xnor U2201 (N_2201,N_1220,N_1013);
or U2202 (N_2202,N_1270,N_1239);
nor U2203 (N_2203,N_1491,N_859);
xor U2204 (N_2204,N_1231,N_1219);
nand U2205 (N_2205,N_1153,N_1075);
or U2206 (N_2206,N_992,N_1285);
and U2207 (N_2207,N_1415,N_961);
nor U2208 (N_2208,N_956,N_1161);
nand U2209 (N_2209,N_783,N_1177);
or U2210 (N_2210,N_811,N_755);
and U2211 (N_2211,N_870,N_1389);
nor U2212 (N_2212,N_1134,N_960);
and U2213 (N_2213,N_1378,N_904);
or U2214 (N_2214,N_1461,N_1364);
and U2215 (N_2215,N_1122,N_1163);
and U2216 (N_2216,N_968,N_1482);
nor U2217 (N_2217,N_1154,N_1187);
nor U2218 (N_2218,N_1185,N_1189);
xor U2219 (N_2219,N_1318,N_1156);
and U2220 (N_2220,N_1211,N_1278);
or U2221 (N_2221,N_963,N_1169);
and U2222 (N_2222,N_804,N_1283);
xnor U2223 (N_2223,N_1310,N_1008);
xnor U2224 (N_2224,N_1195,N_862);
nand U2225 (N_2225,N_1407,N_1481);
xor U2226 (N_2226,N_1035,N_1218);
nand U2227 (N_2227,N_830,N_1394);
or U2228 (N_2228,N_971,N_1263);
nor U2229 (N_2229,N_1404,N_1260);
or U2230 (N_2230,N_1457,N_847);
nand U2231 (N_2231,N_855,N_1465);
xor U2232 (N_2232,N_1199,N_888);
nand U2233 (N_2233,N_1211,N_817);
nor U2234 (N_2234,N_832,N_955);
nand U2235 (N_2235,N_804,N_853);
and U2236 (N_2236,N_978,N_1114);
or U2237 (N_2237,N_1376,N_1400);
nor U2238 (N_2238,N_769,N_886);
or U2239 (N_2239,N_1093,N_784);
nor U2240 (N_2240,N_1055,N_1192);
and U2241 (N_2241,N_1064,N_847);
and U2242 (N_2242,N_1494,N_1317);
nor U2243 (N_2243,N_1242,N_919);
or U2244 (N_2244,N_1085,N_1264);
or U2245 (N_2245,N_1025,N_1057);
nor U2246 (N_2246,N_856,N_1139);
or U2247 (N_2247,N_881,N_1080);
nand U2248 (N_2248,N_1173,N_1164);
nand U2249 (N_2249,N_1333,N_903);
nor U2250 (N_2250,N_1676,N_2102);
nor U2251 (N_2251,N_1706,N_2185);
nand U2252 (N_2252,N_1965,N_2061);
nand U2253 (N_2253,N_1626,N_2156);
nand U2254 (N_2254,N_1636,N_2077);
nand U2255 (N_2255,N_1821,N_1526);
nand U2256 (N_2256,N_1950,N_2037);
xnor U2257 (N_2257,N_2134,N_2201);
and U2258 (N_2258,N_1937,N_1785);
xnor U2259 (N_2259,N_2206,N_1985);
nor U2260 (N_2260,N_1682,N_2232);
and U2261 (N_2261,N_2241,N_2090);
and U2262 (N_2262,N_1705,N_1554);
nor U2263 (N_2263,N_1579,N_1936);
or U2264 (N_2264,N_1601,N_1565);
or U2265 (N_2265,N_1522,N_1661);
and U2266 (N_2266,N_1786,N_2174);
and U2267 (N_2267,N_1769,N_2175);
nor U2268 (N_2268,N_1688,N_1831);
and U2269 (N_2269,N_1544,N_1764);
nand U2270 (N_2270,N_1960,N_1852);
nor U2271 (N_2271,N_1845,N_2111);
nand U2272 (N_2272,N_2179,N_2167);
xor U2273 (N_2273,N_1832,N_2135);
or U2274 (N_2274,N_1798,N_1864);
or U2275 (N_2275,N_2023,N_2049);
nor U2276 (N_2276,N_2073,N_2162);
nor U2277 (N_2277,N_2169,N_1557);
and U2278 (N_2278,N_1805,N_2123);
or U2279 (N_2279,N_1815,N_1904);
nand U2280 (N_2280,N_2119,N_1635);
or U2281 (N_2281,N_1595,N_1602);
nor U2282 (N_2282,N_2198,N_1730);
nor U2283 (N_2283,N_1508,N_2035);
nand U2284 (N_2284,N_1703,N_1589);
and U2285 (N_2285,N_1935,N_1925);
nand U2286 (N_2286,N_1511,N_1613);
xor U2287 (N_2287,N_1963,N_1837);
and U2288 (N_2288,N_2126,N_2074);
nand U2289 (N_2289,N_2099,N_1799);
nor U2290 (N_2290,N_1712,N_1701);
or U2291 (N_2291,N_1932,N_1759);
nor U2292 (N_2292,N_1674,N_2033);
and U2293 (N_2293,N_1671,N_1809);
nand U2294 (N_2294,N_1829,N_1572);
and U2295 (N_2295,N_1934,N_2030);
nor U2296 (N_2296,N_1578,N_1717);
or U2297 (N_2297,N_1833,N_2181);
or U2298 (N_2298,N_1765,N_1728);
nand U2299 (N_2299,N_1693,N_1859);
nand U2300 (N_2300,N_1581,N_1916);
or U2301 (N_2301,N_1822,N_1690);
nand U2302 (N_2302,N_1814,N_2170);
xnor U2303 (N_2303,N_2207,N_1617);
xnor U2304 (N_2304,N_1996,N_1760);
nor U2305 (N_2305,N_1774,N_2021);
and U2306 (N_2306,N_2212,N_1723);
nand U2307 (N_2307,N_2108,N_2112);
nor U2308 (N_2308,N_2139,N_2041);
or U2309 (N_2309,N_2053,N_1640);
xor U2310 (N_2310,N_2187,N_2022);
or U2311 (N_2311,N_1952,N_2028);
or U2312 (N_2312,N_1742,N_1747);
nand U2313 (N_2313,N_1881,N_1862);
and U2314 (N_2314,N_1750,N_1551);
nor U2315 (N_2315,N_1560,N_1724);
nand U2316 (N_2316,N_1989,N_2000);
nor U2317 (N_2317,N_1860,N_2248);
nand U2318 (N_2318,N_2199,N_1642);
xnor U2319 (N_2319,N_2116,N_1625);
xor U2320 (N_2320,N_1888,N_2226);
or U2321 (N_2321,N_2117,N_1972);
and U2322 (N_2322,N_1933,N_1539);
or U2323 (N_2323,N_2032,N_2208);
or U2324 (N_2324,N_1830,N_1971);
nor U2325 (N_2325,N_1944,N_1899);
nand U2326 (N_2326,N_1917,N_1926);
nand U2327 (N_2327,N_1949,N_2018);
nand U2328 (N_2328,N_1974,N_2089);
nand U2329 (N_2329,N_1641,N_1791);
nand U2330 (N_2330,N_1561,N_1817);
nor U2331 (N_2331,N_1722,N_1719);
xnor U2332 (N_2332,N_2164,N_1923);
xor U2333 (N_2333,N_2147,N_1748);
and U2334 (N_2334,N_1930,N_1726);
nand U2335 (N_2335,N_1873,N_1536);
or U2336 (N_2336,N_1563,N_2088);
nor U2337 (N_2337,N_1895,N_1892);
and U2338 (N_2338,N_2106,N_1962);
xor U2339 (N_2339,N_1983,N_1976);
nand U2340 (N_2340,N_1751,N_1597);
nor U2341 (N_2341,N_1796,N_1507);
xor U2342 (N_2342,N_1546,N_2230);
and U2343 (N_2343,N_1919,N_1615);
and U2344 (N_2344,N_1583,N_1900);
xor U2345 (N_2345,N_1826,N_1623);
nand U2346 (N_2346,N_2034,N_1503);
nor U2347 (N_2347,N_1608,N_2245);
and U2348 (N_2348,N_2157,N_1753);
and U2349 (N_2349,N_1953,N_1677);
nor U2350 (N_2350,N_2211,N_1782);
and U2351 (N_2351,N_2184,N_1891);
and U2352 (N_2352,N_1869,N_2075);
and U2353 (N_2353,N_1848,N_1756);
xor U2354 (N_2354,N_1954,N_1741);
nor U2355 (N_2355,N_1847,N_2015);
or U2356 (N_2356,N_2140,N_1681);
and U2357 (N_2357,N_1787,N_2127);
nor U2358 (N_2358,N_1858,N_2224);
nand U2359 (N_2359,N_1992,N_2081);
xor U2360 (N_2360,N_1649,N_2069);
and U2361 (N_2361,N_1594,N_1889);
nand U2362 (N_2362,N_1841,N_2062);
xnor U2363 (N_2363,N_2060,N_1530);
and U2364 (N_2364,N_1757,N_1844);
nand U2365 (N_2365,N_2122,N_2039);
nor U2366 (N_2366,N_1646,N_1927);
nand U2367 (N_2367,N_1660,N_1509);
nand U2368 (N_2368,N_1611,N_1694);
nand U2369 (N_2369,N_1633,N_1648);
nand U2370 (N_2370,N_1905,N_1721);
and U2371 (N_2371,N_2192,N_2209);
nor U2372 (N_2372,N_2172,N_1713);
nor U2373 (N_2373,N_1975,N_1700);
xnor U2374 (N_2374,N_1910,N_1886);
xnor U2375 (N_2375,N_2159,N_1567);
nand U2376 (N_2376,N_2031,N_2176);
xnor U2377 (N_2377,N_1877,N_1518);
or U2378 (N_2378,N_1811,N_1697);
nor U2379 (N_2379,N_2228,N_2138);
or U2380 (N_2380,N_1644,N_1991);
nor U2381 (N_2381,N_1547,N_1995);
or U2382 (N_2382,N_2197,N_1999);
nor U2383 (N_2383,N_1593,N_2001);
nor U2384 (N_2384,N_1612,N_1616);
and U2385 (N_2385,N_1691,N_1915);
and U2386 (N_2386,N_1564,N_2130);
xor U2387 (N_2387,N_1740,N_1708);
and U2388 (N_2388,N_2050,N_2136);
nor U2389 (N_2389,N_2163,N_1857);
or U2390 (N_2390,N_2141,N_1559);
nor U2391 (N_2391,N_2210,N_1780);
and U2392 (N_2392,N_1773,N_1537);
nand U2393 (N_2393,N_1851,N_2182);
nand U2394 (N_2394,N_1793,N_2244);
nand U2395 (N_2395,N_1973,N_1590);
xor U2396 (N_2396,N_1808,N_1517);
xnor U2397 (N_2397,N_1984,N_2149);
and U2398 (N_2398,N_2205,N_1928);
or U2399 (N_2399,N_2144,N_1619);
or U2400 (N_2400,N_1874,N_1970);
nand U2401 (N_2401,N_1894,N_1823);
and U2402 (N_2402,N_1737,N_2124);
xnor U2403 (N_2403,N_1727,N_1512);
or U2404 (N_2404,N_1761,N_1631);
and U2405 (N_2405,N_1609,N_2100);
nand U2406 (N_2406,N_1824,N_2151);
or U2407 (N_2407,N_2150,N_2243);
xnor U2408 (N_2408,N_1659,N_1948);
nor U2409 (N_2409,N_2171,N_2012);
nor U2410 (N_2410,N_2056,N_2084);
nand U2411 (N_2411,N_1673,N_1587);
and U2412 (N_2412,N_1513,N_1678);
xor U2413 (N_2413,N_2190,N_1825);
or U2414 (N_2414,N_1943,N_1592);
nand U2415 (N_2415,N_2045,N_1977);
and U2416 (N_2416,N_2038,N_2096);
and U2417 (N_2417,N_1630,N_1654);
and U2418 (N_2418,N_1647,N_1779);
or U2419 (N_2419,N_1846,N_1994);
nand U2420 (N_2420,N_1514,N_1997);
nand U2421 (N_2421,N_2177,N_1913);
or U2422 (N_2422,N_1951,N_1867);
nor U2423 (N_2423,N_1739,N_1875);
and U2424 (N_2424,N_1502,N_2242);
and U2425 (N_2425,N_1734,N_2145);
nor U2426 (N_2426,N_1736,N_1887);
and U2427 (N_2427,N_1806,N_1820);
nor U2428 (N_2428,N_1692,N_1655);
nor U2429 (N_2429,N_1819,N_1763);
nand U2430 (N_2430,N_1569,N_2218);
nand U2431 (N_2431,N_1622,N_1607);
or U2432 (N_2432,N_1929,N_2026);
nor U2433 (N_2433,N_1783,N_1665);
xnor U2434 (N_2434,N_1709,N_1529);
nor U2435 (N_2435,N_2173,N_2098);
and U2436 (N_2436,N_1521,N_2189);
nor U2437 (N_2437,N_1532,N_1663);
xnor U2438 (N_2438,N_1911,N_1909);
nand U2439 (N_2439,N_2095,N_2233);
and U2440 (N_2440,N_1922,N_2063);
nand U2441 (N_2441,N_2191,N_1777);
or U2442 (N_2442,N_1548,N_2065);
xnor U2443 (N_2443,N_1967,N_1651);
and U2444 (N_2444,N_2094,N_1586);
or U2445 (N_2445,N_1884,N_1657);
xnor U2446 (N_2446,N_1714,N_1772);
nor U2447 (N_2447,N_1800,N_1501);
nand U2448 (N_2448,N_1941,N_1969);
or U2449 (N_2449,N_1901,N_1988);
and U2450 (N_2450,N_2086,N_2082);
nand U2451 (N_2451,N_1638,N_2161);
nor U2452 (N_2452,N_1978,N_1902);
and U2453 (N_2453,N_1543,N_1792);
or U2454 (N_2454,N_1525,N_1653);
or U2455 (N_2455,N_1842,N_1666);
nor U2456 (N_2456,N_2017,N_1542);
xor U2457 (N_2457,N_2165,N_1684);
and U2458 (N_2458,N_2068,N_1720);
xnor U2459 (N_2459,N_2046,N_2129);
nor U2460 (N_2460,N_2066,N_1675);
xnor U2461 (N_2461,N_1998,N_1850);
nand U2462 (N_2462,N_2080,N_2109);
xor U2463 (N_2463,N_1632,N_1614);
and U2464 (N_2464,N_1855,N_1966);
nand U2465 (N_2465,N_2216,N_1744);
or U2466 (N_2466,N_1629,N_1510);
or U2467 (N_2467,N_1685,N_2042);
nand U2468 (N_2468,N_2036,N_1520);
or U2469 (N_2469,N_1914,N_2143);
xnor U2470 (N_2470,N_2019,N_1921);
nand U2471 (N_2471,N_2006,N_1766);
xnor U2472 (N_2472,N_1770,N_1549);
xnor U2473 (N_2473,N_1788,N_1898);
xor U2474 (N_2474,N_1794,N_2220);
xor U2475 (N_2475,N_1880,N_1606);
and U2476 (N_2476,N_2168,N_1958);
and U2477 (N_2477,N_1816,N_1893);
or U2478 (N_2478,N_2240,N_1667);
nand U2479 (N_2479,N_1957,N_2087);
nor U2480 (N_2480,N_2235,N_1696);
and U2481 (N_2481,N_1545,N_2107);
xnor U2482 (N_2482,N_2043,N_1584);
or U2483 (N_2483,N_2152,N_2047);
or U2484 (N_2484,N_2183,N_1679);
or U2485 (N_2485,N_2104,N_1687);
nor U2486 (N_2486,N_1812,N_1868);
xor U2487 (N_2487,N_1878,N_1729);
or U2488 (N_2488,N_1781,N_2079);
xnor U2489 (N_2489,N_1552,N_2202);
nand U2490 (N_2490,N_2203,N_2180);
and U2491 (N_2491,N_1870,N_1840);
nor U2492 (N_2492,N_2057,N_1643);
or U2493 (N_2493,N_1504,N_1573);
nand U2494 (N_2494,N_1818,N_1577);
xnor U2495 (N_2495,N_2221,N_1804);
xor U2496 (N_2496,N_2002,N_1968);
nand U2497 (N_2497,N_2227,N_1531);
or U2498 (N_2498,N_1890,N_1882);
and U2499 (N_2499,N_2091,N_1856);
nor U2500 (N_2500,N_1789,N_1803);
and U2501 (N_2501,N_1698,N_1658);
and U2502 (N_2502,N_2154,N_2114);
nor U2503 (N_2503,N_1735,N_1797);
nor U2504 (N_2504,N_1524,N_1876);
nor U2505 (N_2505,N_2118,N_2029);
or U2506 (N_2506,N_1527,N_2166);
and U2507 (N_2507,N_2016,N_2246);
and U2508 (N_2508,N_1942,N_1515);
and U2509 (N_2509,N_1940,N_2103);
xnor U2510 (N_2510,N_1528,N_1600);
nor U2511 (N_2511,N_1863,N_1538);
and U2512 (N_2512,N_1645,N_2215);
nor U2513 (N_2513,N_1924,N_1585);
and U2514 (N_2514,N_1964,N_1668);
and U2515 (N_2515,N_2219,N_1827);
nand U2516 (N_2516,N_1879,N_2196);
nor U2517 (N_2517,N_2067,N_2051);
and U2518 (N_2518,N_1908,N_2148);
nor U2519 (N_2519,N_1866,N_2040);
xor U2520 (N_2520,N_1986,N_2110);
or U2521 (N_2521,N_1711,N_1566);
or U2522 (N_2522,N_1505,N_1907);
or U2523 (N_2523,N_1699,N_1795);
and U2524 (N_2524,N_1540,N_1835);
nand U2525 (N_2525,N_2249,N_1990);
and U2526 (N_2526,N_2133,N_1749);
nand U2527 (N_2527,N_2153,N_1725);
xnor U2528 (N_2528,N_1634,N_2005);
xor U2529 (N_2529,N_1885,N_1716);
or U2530 (N_2530,N_1621,N_1982);
nor U2531 (N_2531,N_2009,N_1981);
xor U2532 (N_2532,N_2229,N_1775);
nand U2533 (N_2533,N_1523,N_1776);
or U2534 (N_2534,N_2200,N_2217);
xnor U2535 (N_2535,N_1519,N_1556);
and U2536 (N_2536,N_1650,N_1656);
nand U2537 (N_2537,N_2125,N_1738);
nor U2538 (N_2538,N_2078,N_2115);
and U2539 (N_2539,N_1807,N_1550);
nand U2540 (N_2540,N_2083,N_1516);
or U2541 (N_2541,N_1979,N_2113);
nand U2542 (N_2542,N_1718,N_2158);
nor U2543 (N_2543,N_2223,N_1596);
nor U2544 (N_2544,N_2054,N_1627);
nand U2545 (N_2545,N_1534,N_1624);
nand U2546 (N_2546,N_2014,N_2142);
nand U2547 (N_2547,N_1500,N_2193);
and U2548 (N_2548,N_2072,N_2239);
xor U2549 (N_2549,N_1872,N_1506);
nand U2550 (N_2550,N_1733,N_1576);
and U2551 (N_2551,N_1746,N_2178);
nand U2552 (N_2552,N_1903,N_1664);
nand U2553 (N_2553,N_1752,N_1838);
or U2554 (N_2554,N_1810,N_1669);
nor U2555 (N_2555,N_1828,N_1767);
or U2556 (N_2556,N_1670,N_2236);
nor U2557 (N_2557,N_1768,N_2237);
or U2558 (N_2558,N_1853,N_1865);
or U2559 (N_2559,N_1758,N_2238);
and U2560 (N_2560,N_1993,N_1672);
nor U2561 (N_2561,N_1591,N_1707);
nand U2562 (N_2562,N_1562,N_2222);
xnor U2563 (N_2563,N_2186,N_1553);
and U2564 (N_2564,N_2093,N_1689);
and U2565 (N_2565,N_1604,N_2120);
xnor U2566 (N_2566,N_1871,N_2146);
nor U2567 (N_2567,N_2092,N_2204);
xor U2568 (N_2568,N_1784,N_1956);
or U2569 (N_2569,N_2234,N_1732);
or U2570 (N_2570,N_1987,N_1686);
nand U2571 (N_2571,N_2231,N_2105);
xor U2572 (N_2572,N_1906,N_1662);
and U2573 (N_2573,N_1535,N_2052);
nand U2574 (N_2574,N_1704,N_1743);
xor U2575 (N_2575,N_1598,N_1778);
or U2576 (N_2576,N_1813,N_2071);
or U2577 (N_2577,N_1618,N_1558);
nand U2578 (N_2578,N_2247,N_1588);
nor U2579 (N_2579,N_2055,N_2013);
nor U2580 (N_2580,N_1574,N_2064);
nand U2581 (N_2581,N_2194,N_2008);
nor U2582 (N_2582,N_1637,N_2132);
xnor U2583 (N_2583,N_2044,N_1945);
xor U2584 (N_2584,N_2059,N_2010);
or U2585 (N_2585,N_2048,N_1883);
nor U2586 (N_2586,N_1939,N_1610);
nand U2587 (N_2587,N_1580,N_2131);
and U2588 (N_2588,N_1555,N_1599);
nand U2589 (N_2589,N_2213,N_2137);
nor U2590 (N_2590,N_2003,N_1710);
nor U2591 (N_2591,N_1959,N_2020);
and U2592 (N_2592,N_1920,N_1571);
or U2593 (N_2593,N_2004,N_1861);
nand U2594 (N_2594,N_1754,N_1802);
xor U2595 (N_2595,N_1980,N_2070);
nand U2596 (N_2596,N_1762,N_1533);
and U2597 (N_2597,N_1582,N_1575);
or U2598 (N_2598,N_1790,N_1843);
and U2599 (N_2599,N_1715,N_2128);
xnor U2600 (N_2600,N_2024,N_1695);
xnor U2601 (N_2601,N_2101,N_2188);
and U2602 (N_2602,N_1755,N_1639);
xnor U2603 (N_2603,N_1702,N_1849);
or U2604 (N_2604,N_2085,N_1896);
xnor U2605 (N_2605,N_1839,N_1683);
nor U2606 (N_2606,N_2214,N_1745);
or U2607 (N_2607,N_1955,N_1961);
and U2608 (N_2608,N_1771,N_1568);
and U2609 (N_2609,N_1620,N_1801);
nand U2610 (N_2610,N_1570,N_1834);
or U2611 (N_2611,N_2025,N_2097);
nor U2612 (N_2612,N_1912,N_2027);
or U2613 (N_2613,N_2058,N_1938);
nor U2614 (N_2614,N_1946,N_1603);
nor U2615 (N_2615,N_1605,N_1628);
or U2616 (N_2616,N_1680,N_1652);
nor U2617 (N_2617,N_2011,N_2007);
or U2618 (N_2618,N_1918,N_1947);
xor U2619 (N_2619,N_2160,N_1731);
nor U2620 (N_2620,N_1836,N_2155);
nand U2621 (N_2621,N_2121,N_2195);
xor U2622 (N_2622,N_1541,N_2076);
nor U2623 (N_2623,N_1931,N_1854);
or U2624 (N_2624,N_1897,N_2225);
nand U2625 (N_2625,N_2241,N_2203);
nor U2626 (N_2626,N_1640,N_1693);
nor U2627 (N_2627,N_2119,N_1637);
nand U2628 (N_2628,N_1564,N_2178);
or U2629 (N_2629,N_1703,N_1954);
nand U2630 (N_2630,N_1911,N_1781);
or U2631 (N_2631,N_1792,N_2094);
nor U2632 (N_2632,N_1525,N_1754);
nor U2633 (N_2633,N_1927,N_1941);
xnor U2634 (N_2634,N_1853,N_1693);
xnor U2635 (N_2635,N_1742,N_1637);
and U2636 (N_2636,N_1821,N_2171);
nand U2637 (N_2637,N_1849,N_1850);
xnor U2638 (N_2638,N_1701,N_1690);
xnor U2639 (N_2639,N_1977,N_1562);
xor U2640 (N_2640,N_1509,N_1926);
nand U2641 (N_2641,N_1690,N_1829);
nand U2642 (N_2642,N_1621,N_1762);
nand U2643 (N_2643,N_2174,N_1874);
xor U2644 (N_2644,N_2215,N_1557);
and U2645 (N_2645,N_1606,N_1770);
nand U2646 (N_2646,N_2078,N_1651);
nand U2647 (N_2647,N_2001,N_2148);
and U2648 (N_2648,N_1990,N_1712);
nor U2649 (N_2649,N_2231,N_1524);
xor U2650 (N_2650,N_1592,N_1528);
or U2651 (N_2651,N_2054,N_2019);
and U2652 (N_2652,N_2063,N_2190);
and U2653 (N_2653,N_1995,N_1934);
xor U2654 (N_2654,N_1529,N_2155);
or U2655 (N_2655,N_1538,N_2061);
xnor U2656 (N_2656,N_2233,N_2134);
nor U2657 (N_2657,N_1634,N_1619);
nor U2658 (N_2658,N_2082,N_2045);
nand U2659 (N_2659,N_2232,N_1698);
or U2660 (N_2660,N_2220,N_1763);
xnor U2661 (N_2661,N_1506,N_2210);
xnor U2662 (N_2662,N_1972,N_2219);
and U2663 (N_2663,N_1985,N_1652);
nand U2664 (N_2664,N_2017,N_2200);
xnor U2665 (N_2665,N_1817,N_1846);
and U2666 (N_2666,N_1658,N_1558);
nor U2667 (N_2667,N_1776,N_1983);
nor U2668 (N_2668,N_2160,N_1606);
or U2669 (N_2669,N_1779,N_1633);
nor U2670 (N_2670,N_1846,N_1573);
or U2671 (N_2671,N_1921,N_1929);
and U2672 (N_2672,N_1679,N_1617);
xor U2673 (N_2673,N_1705,N_1817);
nand U2674 (N_2674,N_1924,N_1797);
or U2675 (N_2675,N_1918,N_1718);
and U2676 (N_2676,N_2084,N_1608);
nor U2677 (N_2677,N_2117,N_2223);
nand U2678 (N_2678,N_1723,N_2220);
and U2679 (N_2679,N_1862,N_2159);
and U2680 (N_2680,N_2004,N_1954);
xor U2681 (N_2681,N_1995,N_1892);
or U2682 (N_2682,N_1729,N_1614);
nand U2683 (N_2683,N_1514,N_2151);
nor U2684 (N_2684,N_1761,N_1935);
nor U2685 (N_2685,N_1857,N_1768);
or U2686 (N_2686,N_1997,N_1532);
and U2687 (N_2687,N_1857,N_1815);
or U2688 (N_2688,N_2004,N_1566);
or U2689 (N_2689,N_1754,N_1548);
and U2690 (N_2690,N_2043,N_2073);
xnor U2691 (N_2691,N_2030,N_2057);
and U2692 (N_2692,N_1823,N_1587);
nand U2693 (N_2693,N_1885,N_1538);
nor U2694 (N_2694,N_2094,N_2132);
nor U2695 (N_2695,N_2153,N_1689);
nor U2696 (N_2696,N_1515,N_1694);
nand U2697 (N_2697,N_2151,N_1965);
xnor U2698 (N_2698,N_1857,N_2025);
nand U2699 (N_2699,N_1874,N_2085);
xnor U2700 (N_2700,N_1947,N_2221);
nand U2701 (N_2701,N_2153,N_1743);
xor U2702 (N_2702,N_1954,N_1895);
nor U2703 (N_2703,N_1953,N_1936);
xor U2704 (N_2704,N_1734,N_2077);
nor U2705 (N_2705,N_2001,N_2248);
and U2706 (N_2706,N_1973,N_1912);
nor U2707 (N_2707,N_1684,N_1682);
nand U2708 (N_2708,N_1613,N_2196);
or U2709 (N_2709,N_1642,N_1950);
and U2710 (N_2710,N_1680,N_1722);
and U2711 (N_2711,N_1980,N_1986);
xor U2712 (N_2712,N_1912,N_1638);
and U2713 (N_2713,N_1573,N_1505);
nand U2714 (N_2714,N_1851,N_1852);
nand U2715 (N_2715,N_1836,N_2191);
or U2716 (N_2716,N_2232,N_1701);
xnor U2717 (N_2717,N_1900,N_1603);
and U2718 (N_2718,N_1858,N_1857);
nand U2719 (N_2719,N_1810,N_1998);
or U2720 (N_2720,N_2245,N_1922);
or U2721 (N_2721,N_1631,N_1504);
nand U2722 (N_2722,N_1868,N_2152);
nor U2723 (N_2723,N_1705,N_1843);
and U2724 (N_2724,N_1522,N_1971);
nor U2725 (N_2725,N_1568,N_2059);
nor U2726 (N_2726,N_2103,N_1863);
xnor U2727 (N_2727,N_1979,N_1683);
nor U2728 (N_2728,N_2053,N_1814);
and U2729 (N_2729,N_2077,N_1765);
xor U2730 (N_2730,N_1963,N_2182);
nand U2731 (N_2731,N_1684,N_2072);
nor U2732 (N_2732,N_1832,N_1933);
nor U2733 (N_2733,N_1528,N_1926);
nor U2734 (N_2734,N_1503,N_2090);
and U2735 (N_2735,N_1899,N_1553);
and U2736 (N_2736,N_1554,N_1764);
nor U2737 (N_2737,N_1609,N_1881);
nand U2738 (N_2738,N_2075,N_1538);
or U2739 (N_2739,N_1687,N_2148);
or U2740 (N_2740,N_2108,N_1946);
xnor U2741 (N_2741,N_1891,N_2186);
and U2742 (N_2742,N_1556,N_1666);
xnor U2743 (N_2743,N_1970,N_1816);
and U2744 (N_2744,N_1671,N_1524);
nor U2745 (N_2745,N_1833,N_2188);
and U2746 (N_2746,N_1783,N_1813);
and U2747 (N_2747,N_1660,N_2165);
xor U2748 (N_2748,N_1713,N_1568);
and U2749 (N_2749,N_1738,N_2176);
and U2750 (N_2750,N_1923,N_1942);
nor U2751 (N_2751,N_1884,N_1768);
xor U2752 (N_2752,N_1823,N_1550);
and U2753 (N_2753,N_1689,N_1713);
and U2754 (N_2754,N_1679,N_1716);
nand U2755 (N_2755,N_2143,N_1933);
nor U2756 (N_2756,N_2023,N_1909);
nor U2757 (N_2757,N_2077,N_1815);
xnor U2758 (N_2758,N_1525,N_1938);
nand U2759 (N_2759,N_1879,N_1606);
nor U2760 (N_2760,N_1966,N_1501);
xnor U2761 (N_2761,N_1624,N_1978);
nor U2762 (N_2762,N_1813,N_1831);
or U2763 (N_2763,N_1864,N_1515);
nand U2764 (N_2764,N_1502,N_2118);
nand U2765 (N_2765,N_1750,N_1540);
nor U2766 (N_2766,N_2188,N_1987);
or U2767 (N_2767,N_1814,N_1982);
or U2768 (N_2768,N_2204,N_1509);
or U2769 (N_2769,N_1529,N_2240);
or U2770 (N_2770,N_1819,N_1701);
xor U2771 (N_2771,N_1531,N_2005);
or U2772 (N_2772,N_2106,N_1846);
or U2773 (N_2773,N_2134,N_1541);
nor U2774 (N_2774,N_1780,N_1591);
nor U2775 (N_2775,N_2171,N_1605);
or U2776 (N_2776,N_1950,N_1530);
or U2777 (N_2777,N_1983,N_2178);
nor U2778 (N_2778,N_1985,N_2091);
nand U2779 (N_2779,N_2220,N_2104);
or U2780 (N_2780,N_1964,N_1693);
xor U2781 (N_2781,N_1979,N_2197);
and U2782 (N_2782,N_2025,N_2020);
nand U2783 (N_2783,N_1570,N_1882);
and U2784 (N_2784,N_2095,N_1596);
and U2785 (N_2785,N_2057,N_2163);
xnor U2786 (N_2786,N_2239,N_1981);
nor U2787 (N_2787,N_2174,N_1960);
nand U2788 (N_2788,N_1516,N_1997);
or U2789 (N_2789,N_2163,N_2160);
nor U2790 (N_2790,N_1915,N_1608);
or U2791 (N_2791,N_1649,N_2124);
xor U2792 (N_2792,N_1604,N_2074);
xor U2793 (N_2793,N_1616,N_1915);
nor U2794 (N_2794,N_1822,N_1875);
nand U2795 (N_2795,N_1874,N_1964);
and U2796 (N_2796,N_2047,N_1711);
or U2797 (N_2797,N_1584,N_1738);
nand U2798 (N_2798,N_2068,N_2014);
and U2799 (N_2799,N_1715,N_2226);
nor U2800 (N_2800,N_1883,N_1761);
and U2801 (N_2801,N_2019,N_1892);
xor U2802 (N_2802,N_2037,N_1602);
and U2803 (N_2803,N_1845,N_2179);
or U2804 (N_2804,N_2010,N_1512);
xor U2805 (N_2805,N_1796,N_2046);
nor U2806 (N_2806,N_1654,N_1647);
nor U2807 (N_2807,N_1625,N_1885);
nand U2808 (N_2808,N_1945,N_1724);
and U2809 (N_2809,N_2198,N_1579);
or U2810 (N_2810,N_2196,N_1988);
nand U2811 (N_2811,N_1802,N_1667);
nor U2812 (N_2812,N_1964,N_1659);
xnor U2813 (N_2813,N_2155,N_1736);
nor U2814 (N_2814,N_1684,N_1604);
nand U2815 (N_2815,N_1672,N_2249);
nand U2816 (N_2816,N_1997,N_1789);
xor U2817 (N_2817,N_1637,N_1737);
or U2818 (N_2818,N_2054,N_1910);
xor U2819 (N_2819,N_1531,N_1627);
nor U2820 (N_2820,N_1856,N_1625);
or U2821 (N_2821,N_1727,N_1563);
and U2822 (N_2822,N_1577,N_1989);
nor U2823 (N_2823,N_2189,N_1788);
xor U2824 (N_2824,N_2209,N_1692);
or U2825 (N_2825,N_2231,N_1961);
nand U2826 (N_2826,N_2154,N_1888);
nand U2827 (N_2827,N_2249,N_1629);
nand U2828 (N_2828,N_1928,N_1685);
nor U2829 (N_2829,N_2150,N_1563);
xnor U2830 (N_2830,N_2011,N_2069);
xnor U2831 (N_2831,N_1712,N_1997);
and U2832 (N_2832,N_2103,N_1816);
nand U2833 (N_2833,N_1884,N_1778);
or U2834 (N_2834,N_1686,N_2106);
and U2835 (N_2835,N_1979,N_2037);
or U2836 (N_2836,N_1962,N_1907);
and U2837 (N_2837,N_1510,N_1631);
xor U2838 (N_2838,N_2240,N_1938);
nor U2839 (N_2839,N_1805,N_1611);
and U2840 (N_2840,N_1522,N_1857);
xor U2841 (N_2841,N_2118,N_2144);
or U2842 (N_2842,N_1587,N_1635);
nand U2843 (N_2843,N_2009,N_1576);
nor U2844 (N_2844,N_1543,N_1836);
or U2845 (N_2845,N_1529,N_1743);
nand U2846 (N_2846,N_1750,N_1729);
nand U2847 (N_2847,N_2046,N_2228);
nor U2848 (N_2848,N_2219,N_2135);
nand U2849 (N_2849,N_2093,N_1792);
and U2850 (N_2850,N_2229,N_2160);
xor U2851 (N_2851,N_1609,N_1569);
nand U2852 (N_2852,N_2192,N_2097);
or U2853 (N_2853,N_1921,N_2095);
or U2854 (N_2854,N_1754,N_1909);
and U2855 (N_2855,N_1658,N_2199);
and U2856 (N_2856,N_1937,N_2125);
and U2857 (N_2857,N_1943,N_1902);
nand U2858 (N_2858,N_2233,N_1863);
nor U2859 (N_2859,N_1521,N_1673);
and U2860 (N_2860,N_1949,N_2076);
xor U2861 (N_2861,N_2079,N_2068);
xor U2862 (N_2862,N_1703,N_1545);
or U2863 (N_2863,N_1805,N_2129);
nand U2864 (N_2864,N_1952,N_2016);
xor U2865 (N_2865,N_1748,N_1862);
xnor U2866 (N_2866,N_2107,N_1666);
and U2867 (N_2867,N_1715,N_1946);
nor U2868 (N_2868,N_2124,N_1665);
xor U2869 (N_2869,N_1530,N_1574);
nand U2870 (N_2870,N_1809,N_2092);
nand U2871 (N_2871,N_1898,N_1894);
nor U2872 (N_2872,N_1689,N_1780);
nor U2873 (N_2873,N_2117,N_1623);
or U2874 (N_2874,N_1737,N_1957);
nor U2875 (N_2875,N_2008,N_1559);
xnor U2876 (N_2876,N_1877,N_1723);
nand U2877 (N_2877,N_2103,N_1680);
nand U2878 (N_2878,N_1785,N_2048);
and U2879 (N_2879,N_1565,N_2161);
or U2880 (N_2880,N_2182,N_1921);
or U2881 (N_2881,N_2202,N_1519);
nor U2882 (N_2882,N_1608,N_1641);
and U2883 (N_2883,N_1553,N_2054);
nor U2884 (N_2884,N_1639,N_1972);
xor U2885 (N_2885,N_1741,N_1821);
nand U2886 (N_2886,N_2038,N_1722);
or U2887 (N_2887,N_1941,N_2207);
xnor U2888 (N_2888,N_1533,N_1684);
xor U2889 (N_2889,N_2156,N_1747);
or U2890 (N_2890,N_1988,N_1729);
nand U2891 (N_2891,N_2169,N_1821);
nor U2892 (N_2892,N_1500,N_1913);
or U2893 (N_2893,N_1927,N_2134);
and U2894 (N_2894,N_1583,N_2018);
nand U2895 (N_2895,N_2200,N_1566);
nor U2896 (N_2896,N_1865,N_1548);
or U2897 (N_2897,N_1709,N_2171);
nand U2898 (N_2898,N_1501,N_1670);
xor U2899 (N_2899,N_1852,N_1875);
xnor U2900 (N_2900,N_1565,N_1586);
nor U2901 (N_2901,N_2177,N_1791);
xor U2902 (N_2902,N_1760,N_1930);
nand U2903 (N_2903,N_1523,N_1811);
nand U2904 (N_2904,N_1908,N_2220);
nor U2905 (N_2905,N_2107,N_2001);
and U2906 (N_2906,N_1889,N_2046);
xnor U2907 (N_2907,N_1609,N_1885);
and U2908 (N_2908,N_1680,N_2206);
or U2909 (N_2909,N_1739,N_1975);
nand U2910 (N_2910,N_1997,N_1649);
nand U2911 (N_2911,N_1773,N_1774);
nand U2912 (N_2912,N_2137,N_1851);
xor U2913 (N_2913,N_1549,N_1931);
nor U2914 (N_2914,N_1680,N_2082);
nand U2915 (N_2915,N_1879,N_1706);
nand U2916 (N_2916,N_1927,N_1921);
xnor U2917 (N_2917,N_2170,N_2204);
xnor U2918 (N_2918,N_1535,N_1766);
or U2919 (N_2919,N_2044,N_2095);
xnor U2920 (N_2920,N_2232,N_1651);
or U2921 (N_2921,N_1760,N_2094);
or U2922 (N_2922,N_1732,N_1579);
nand U2923 (N_2923,N_1684,N_1542);
or U2924 (N_2924,N_1784,N_1965);
nand U2925 (N_2925,N_1966,N_2185);
nor U2926 (N_2926,N_2064,N_1694);
xnor U2927 (N_2927,N_2126,N_1967);
nand U2928 (N_2928,N_1667,N_2123);
nor U2929 (N_2929,N_2058,N_2100);
nor U2930 (N_2930,N_1690,N_2182);
nor U2931 (N_2931,N_2174,N_2112);
xor U2932 (N_2932,N_2053,N_1869);
nor U2933 (N_2933,N_1536,N_1741);
nor U2934 (N_2934,N_1537,N_2227);
nor U2935 (N_2935,N_1598,N_1517);
and U2936 (N_2936,N_1696,N_1645);
nor U2937 (N_2937,N_1666,N_1988);
nor U2938 (N_2938,N_1703,N_2246);
or U2939 (N_2939,N_2022,N_2244);
xor U2940 (N_2940,N_2004,N_1592);
nand U2941 (N_2941,N_1969,N_2065);
nor U2942 (N_2942,N_1781,N_1529);
or U2943 (N_2943,N_1506,N_2202);
nor U2944 (N_2944,N_1524,N_1613);
nand U2945 (N_2945,N_1614,N_2029);
or U2946 (N_2946,N_1834,N_2074);
or U2947 (N_2947,N_2117,N_2146);
and U2948 (N_2948,N_1796,N_2034);
and U2949 (N_2949,N_1694,N_1649);
xor U2950 (N_2950,N_1672,N_2244);
nor U2951 (N_2951,N_2219,N_2044);
or U2952 (N_2952,N_1637,N_1507);
nand U2953 (N_2953,N_1785,N_1768);
nor U2954 (N_2954,N_2205,N_1640);
and U2955 (N_2955,N_1740,N_1883);
xor U2956 (N_2956,N_1563,N_2012);
and U2957 (N_2957,N_1965,N_2145);
or U2958 (N_2958,N_1541,N_1991);
and U2959 (N_2959,N_1540,N_1687);
or U2960 (N_2960,N_1987,N_1578);
nand U2961 (N_2961,N_1865,N_1627);
xor U2962 (N_2962,N_2025,N_1775);
xor U2963 (N_2963,N_1932,N_2106);
nor U2964 (N_2964,N_1668,N_1526);
xor U2965 (N_2965,N_1552,N_2027);
and U2966 (N_2966,N_1798,N_1857);
nand U2967 (N_2967,N_1605,N_1953);
or U2968 (N_2968,N_1945,N_1510);
nor U2969 (N_2969,N_1960,N_2132);
nand U2970 (N_2970,N_1960,N_1797);
nand U2971 (N_2971,N_1932,N_1990);
xnor U2972 (N_2972,N_1753,N_1596);
nor U2973 (N_2973,N_1705,N_2029);
and U2974 (N_2974,N_2119,N_1775);
xor U2975 (N_2975,N_1700,N_2087);
nor U2976 (N_2976,N_1608,N_2075);
or U2977 (N_2977,N_1586,N_2244);
xor U2978 (N_2978,N_2199,N_1859);
and U2979 (N_2979,N_1719,N_1605);
nand U2980 (N_2980,N_1721,N_1722);
and U2981 (N_2981,N_1680,N_2139);
nor U2982 (N_2982,N_2179,N_2053);
nand U2983 (N_2983,N_2064,N_2131);
nand U2984 (N_2984,N_2048,N_1789);
xor U2985 (N_2985,N_1761,N_2239);
xor U2986 (N_2986,N_1679,N_1952);
or U2987 (N_2987,N_1845,N_1581);
nand U2988 (N_2988,N_1668,N_2122);
nor U2989 (N_2989,N_2154,N_1640);
and U2990 (N_2990,N_1736,N_1567);
or U2991 (N_2991,N_2031,N_1952);
nand U2992 (N_2992,N_1845,N_1621);
and U2993 (N_2993,N_2012,N_1602);
and U2994 (N_2994,N_1693,N_2152);
nand U2995 (N_2995,N_1904,N_2099);
nand U2996 (N_2996,N_1504,N_1989);
or U2997 (N_2997,N_2108,N_2202);
nor U2998 (N_2998,N_1645,N_1871);
nand U2999 (N_2999,N_1667,N_1697);
and U3000 (N_3000,N_2705,N_2315);
and U3001 (N_3001,N_2522,N_2472);
and U3002 (N_3002,N_2475,N_2911);
nand U3003 (N_3003,N_2785,N_2685);
xnor U3004 (N_3004,N_2893,N_2488);
or U3005 (N_3005,N_2840,N_2741);
or U3006 (N_3006,N_2393,N_2380);
or U3007 (N_3007,N_2977,N_2353);
or U3008 (N_3008,N_2336,N_2632);
and U3009 (N_3009,N_2426,N_2326);
xnor U3010 (N_3010,N_2777,N_2363);
and U3011 (N_3011,N_2787,N_2819);
or U3012 (N_3012,N_2409,N_2804);
nand U3013 (N_3013,N_2917,N_2290);
and U3014 (N_3014,N_2652,N_2394);
nor U3015 (N_3015,N_2993,N_2406);
xnor U3016 (N_3016,N_2817,N_2265);
or U3017 (N_3017,N_2355,N_2661);
xor U3018 (N_3018,N_2980,N_2562);
nand U3019 (N_3019,N_2937,N_2979);
and U3020 (N_3020,N_2465,N_2847);
or U3021 (N_3021,N_2384,N_2591);
and U3022 (N_3022,N_2533,N_2324);
nor U3023 (N_3023,N_2960,N_2619);
nor U3024 (N_3024,N_2594,N_2398);
nor U3025 (N_3025,N_2359,N_2816);
nor U3026 (N_3026,N_2833,N_2307);
nand U3027 (N_3027,N_2639,N_2318);
and U3028 (N_3028,N_2736,N_2293);
nor U3029 (N_3029,N_2779,N_2518);
xor U3030 (N_3030,N_2259,N_2669);
xor U3031 (N_3031,N_2373,N_2360);
and U3032 (N_3032,N_2545,N_2338);
nand U3033 (N_3033,N_2640,N_2861);
and U3034 (N_3034,N_2710,N_2614);
or U3035 (N_3035,N_2988,N_2728);
nand U3036 (N_3036,N_2814,N_2854);
nor U3037 (N_3037,N_2958,N_2752);
or U3038 (N_3038,N_2309,N_2289);
nor U3039 (N_3039,N_2953,N_2775);
nand U3040 (N_3040,N_2482,N_2744);
xor U3041 (N_3041,N_2948,N_2763);
xor U3042 (N_3042,N_2370,N_2949);
and U3043 (N_3043,N_2676,N_2994);
or U3044 (N_3044,N_2301,N_2633);
xnor U3045 (N_3045,N_2410,N_2497);
and U3046 (N_3046,N_2456,N_2564);
or U3047 (N_3047,N_2974,N_2563);
or U3048 (N_3048,N_2962,N_2824);
xnor U3049 (N_3049,N_2292,N_2449);
or U3050 (N_3050,N_2369,N_2534);
nand U3051 (N_3051,N_2478,N_2294);
or U3052 (N_3052,N_2670,N_2807);
nor U3053 (N_3053,N_2725,N_2759);
nand U3054 (N_3054,N_2445,N_2252);
and U3055 (N_3055,N_2646,N_2727);
xnor U3056 (N_3056,N_2895,N_2320);
nand U3057 (N_3057,N_2930,N_2490);
nand U3058 (N_3058,N_2766,N_2899);
and U3059 (N_3059,N_2712,N_2368);
xor U3060 (N_3060,N_2657,N_2417);
and U3061 (N_3061,N_2638,N_2890);
nor U3062 (N_3062,N_2595,N_2566);
and U3063 (N_3063,N_2365,N_2486);
or U3064 (N_3064,N_2623,N_2590);
nand U3065 (N_3065,N_2837,N_2715);
xnor U3066 (N_3066,N_2720,N_2733);
nand U3067 (N_3067,N_2458,N_2898);
nor U3068 (N_3068,N_2706,N_2946);
or U3069 (N_3069,N_2574,N_2656);
nand U3070 (N_3070,N_2622,N_2361);
xor U3071 (N_3071,N_2603,N_2922);
and U3072 (N_3072,N_2257,N_2467);
xnor U3073 (N_3073,N_2471,N_2615);
or U3074 (N_3074,N_2919,N_2910);
or U3075 (N_3075,N_2878,N_2912);
nand U3076 (N_3076,N_2538,N_2317);
nand U3077 (N_3077,N_2354,N_2892);
and U3078 (N_3078,N_2383,N_2653);
or U3079 (N_3079,N_2857,N_2978);
nand U3080 (N_3080,N_2842,N_2871);
or U3081 (N_3081,N_2726,N_2843);
xnor U3082 (N_3082,N_2966,N_2598);
xor U3083 (N_3083,N_2851,N_2902);
xor U3084 (N_3084,N_2561,N_2551);
or U3085 (N_3085,N_2802,N_2793);
xor U3086 (N_3086,N_2404,N_2516);
or U3087 (N_3087,N_2553,N_2631);
or U3088 (N_3088,N_2663,N_2778);
xor U3089 (N_3089,N_2424,N_2348);
xor U3090 (N_3090,N_2274,N_2378);
or U3091 (N_3091,N_2796,N_2375);
nor U3092 (N_3092,N_2511,N_2938);
and U3093 (N_3093,N_2700,N_2959);
xor U3094 (N_3094,N_2691,N_2675);
xnor U3095 (N_3095,N_2955,N_2961);
or U3096 (N_3096,N_2460,N_2846);
xor U3097 (N_3097,N_2559,N_2396);
nor U3098 (N_3098,N_2729,N_2903);
nand U3099 (N_3099,N_2602,N_2681);
and U3100 (N_3100,N_2283,N_2501);
nand U3101 (N_3101,N_2413,N_2957);
nor U3102 (N_3102,N_2434,N_2286);
and U3103 (N_3103,N_2331,N_2649);
nand U3104 (N_3104,N_2621,N_2399);
or U3105 (N_3105,N_2956,N_2818);
nand U3106 (N_3106,N_2872,N_2385);
xnor U3107 (N_3107,N_2708,N_2836);
or U3108 (N_3108,N_2476,N_2305);
or U3109 (N_3109,N_2341,N_2431);
xor U3110 (N_3110,N_2500,N_2342);
nor U3111 (N_3111,N_2769,N_2971);
nor U3112 (N_3112,N_2512,N_2882);
nand U3113 (N_3113,N_2717,N_2267);
and U3114 (N_3114,N_2481,N_2693);
and U3115 (N_3115,N_2666,N_2701);
and U3116 (N_3116,N_2635,N_2643);
nand U3117 (N_3117,N_2250,N_2584);
nor U3118 (N_3118,N_2346,N_2873);
xnor U3119 (N_3119,N_2269,N_2936);
xnor U3120 (N_3120,N_2514,N_2865);
nand U3121 (N_3121,N_2826,N_2419);
nand U3122 (N_3122,N_2548,N_2916);
nand U3123 (N_3123,N_2673,N_2783);
xnor U3124 (N_3124,N_2822,N_2254);
or U3125 (N_3125,N_2680,N_2592);
and U3126 (N_3126,N_2671,N_2862);
or U3127 (N_3127,N_2739,N_2894);
nand U3128 (N_3128,N_2414,N_2784);
nand U3129 (N_3129,N_2588,N_2925);
xor U3130 (N_3130,N_2255,N_2835);
nor U3131 (N_3131,N_2886,N_2698);
nor U3132 (N_3132,N_2637,N_2844);
xnor U3133 (N_3133,N_2299,N_2904);
and U3134 (N_3134,N_2811,N_2300);
xor U3135 (N_3135,N_2291,N_2374);
nand U3136 (N_3136,N_2275,N_2625);
nor U3137 (N_3137,N_2358,N_2996);
or U3138 (N_3138,N_2866,N_2770);
or U3139 (N_3139,N_2884,N_2780);
nor U3140 (N_3140,N_2907,N_2468);
xor U3141 (N_3141,N_2552,N_2998);
nor U3142 (N_3142,N_2343,N_2596);
and U3143 (N_3143,N_2483,N_2253);
nor U3144 (N_3144,N_2987,N_2513);
and U3145 (N_3145,N_2485,N_2823);
nand U3146 (N_3146,N_2412,N_2304);
nor U3147 (N_3147,N_2499,N_2968);
xnor U3148 (N_3148,N_2746,N_2812);
and U3149 (N_3149,N_2450,N_2423);
nor U3150 (N_3150,N_2609,N_2781);
and U3151 (N_3151,N_2427,N_2721);
or U3152 (N_3152,N_2992,N_2573);
and U3153 (N_3153,N_2947,N_2575);
and U3154 (N_3154,N_2913,N_2580);
xnor U3155 (N_3155,N_2755,N_2528);
xor U3156 (N_3156,N_2549,N_2703);
or U3157 (N_3157,N_2896,N_2487);
xnor U3158 (N_3158,N_2737,N_2768);
and U3159 (N_3159,N_2848,N_2757);
nand U3160 (N_3160,N_2760,N_2340);
nor U3161 (N_3161,N_2924,N_2489);
or U3162 (N_3162,N_2498,N_2422);
nand U3163 (N_3163,N_2734,N_2738);
xnor U3164 (N_3164,N_2352,N_2859);
nor U3165 (N_3165,N_2880,N_2745);
or U3166 (N_3166,N_2601,N_2525);
xnor U3167 (N_3167,N_2665,N_2690);
nor U3168 (N_3168,N_2443,N_2801);
xnor U3169 (N_3169,N_2923,N_2942);
or U3170 (N_3170,N_2897,N_2765);
nor U3171 (N_3171,N_2334,N_2918);
and U3172 (N_3172,N_2504,N_2654);
nor U3173 (N_3173,N_2664,N_2366);
xnor U3174 (N_3174,N_2411,N_2782);
nor U3175 (N_3175,N_2333,N_2628);
and U3176 (N_3176,N_2322,N_2277);
xnor U3177 (N_3177,N_2891,N_2287);
nor U3178 (N_3178,N_2810,N_2762);
or U3179 (N_3179,N_2403,N_2550);
and U3180 (N_3180,N_2767,N_2951);
and U3181 (N_3181,N_2952,N_2527);
nand U3182 (N_3182,N_2382,N_2448);
nand U3183 (N_3183,N_2695,N_2776);
nand U3184 (N_3184,N_2345,N_2532);
or U3185 (N_3185,N_2576,N_2735);
xnor U3186 (N_3186,N_2906,N_2935);
and U3187 (N_3187,N_2266,N_2418);
nand U3188 (N_3188,N_2672,N_2586);
nand U3189 (N_3189,N_2794,N_2932);
nand U3190 (N_3190,N_2707,N_2308);
nand U3191 (N_3191,N_2260,N_2644);
xnor U3192 (N_3192,N_2578,N_2477);
nor U3193 (N_3193,N_2507,N_2928);
or U3194 (N_3194,N_2986,N_2272);
or U3195 (N_3195,N_2647,N_2604);
nand U3196 (N_3196,N_2709,N_2539);
nand U3197 (N_3197,N_2645,N_2391);
xor U3198 (N_3198,N_2492,N_2428);
nor U3199 (N_3199,N_2885,N_2742);
xor U3200 (N_3200,N_2838,N_2941);
xor U3201 (N_3201,N_2756,N_2339);
nor U3202 (N_3202,N_2610,N_2839);
and U3203 (N_3203,N_2479,N_2876);
or U3204 (N_3204,N_2630,N_2641);
and U3205 (N_3205,N_2397,N_2557);
xnor U3206 (N_3206,N_2798,N_2616);
nand U3207 (N_3207,N_2909,N_2626);
nor U3208 (N_3208,N_2774,N_2939);
nor U3209 (N_3209,N_2929,N_2920);
xor U3210 (N_3210,N_2702,N_2599);
and U3211 (N_3211,N_2432,N_2276);
and U3212 (N_3212,N_2420,N_2852);
nand U3213 (N_3213,N_2668,N_2316);
and U3214 (N_3214,N_2459,N_2312);
or U3215 (N_3215,N_2439,N_2883);
or U3216 (N_3216,N_2350,N_2327);
nand U3217 (N_3217,N_2430,N_2901);
and U3218 (N_3218,N_2864,N_2560);
and U3219 (N_3219,N_2806,N_2808);
xnor U3220 (N_3220,N_2933,N_2973);
and U3221 (N_3221,N_2981,N_2392);
nor U3222 (N_3222,N_2674,N_2302);
and U3223 (N_3223,N_2461,N_2732);
xnor U3224 (N_3224,N_2803,N_2651);
xnor U3225 (N_3225,N_2473,N_2773);
or U3226 (N_3226,N_2634,N_2268);
and U3227 (N_3227,N_2743,N_2642);
xnor U3228 (N_3228,N_2323,N_2386);
xor U3229 (N_3229,N_2607,N_2570);
and U3230 (N_3230,N_2372,N_2261);
nor U3231 (N_3231,N_2758,N_2914);
and U3232 (N_3232,N_2335,N_2306);
nand U3233 (N_3233,N_2624,N_2694);
and U3234 (N_3234,N_2845,N_2531);
nand U3235 (N_3235,N_2815,N_2799);
nand U3236 (N_3236,N_2442,N_2658);
nor U3237 (N_3237,N_2696,N_2298);
xor U3238 (N_3238,N_2362,N_2530);
or U3239 (N_3239,N_2258,N_2526);
and U3240 (N_3240,N_2975,N_2853);
nand U3241 (N_3241,N_2889,N_2517);
or U3242 (N_3242,N_2496,N_2860);
nor U3243 (N_3243,N_2682,N_2569);
and U3244 (N_3244,N_2416,N_2699);
xor U3245 (N_3245,N_2377,N_2484);
xnor U3246 (N_3246,N_2888,N_2332);
nand U3247 (N_3247,N_2688,N_2795);
and U3248 (N_3248,N_2608,N_2466);
nand U3249 (N_3249,N_2985,N_2357);
or U3250 (N_3250,N_2470,N_2281);
nand U3251 (N_3251,N_2821,N_2521);
or U3252 (N_3252,N_2697,N_2510);
nor U3253 (N_3253,N_2515,N_2921);
xnor U3254 (N_3254,N_2263,N_2571);
and U3255 (N_3255,N_2667,N_2542);
and U3256 (N_3256,N_2991,N_2719);
nand U3257 (N_3257,N_2764,N_2344);
or U3258 (N_3258,N_2296,N_2612);
nor U3259 (N_3259,N_2330,N_2415);
nand U3260 (N_3260,N_2310,N_2792);
nor U3261 (N_3261,N_2444,N_2454);
nand U3262 (N_3262,N_2943,N_2648);
xnor U3263 (N_3263,N_2529,N_2905);
nand U3264 (N_3264,N_2827,N_2390);
and U3265 (N_3265,N_2984,N_2543);
nand U3266 (N_3266,N_2367,N_2683);
nand U3267 (N_3267,N_2704,N_2989);
nand U3268 (N_3268,N_2407,N_2435);
nor U3269 (N_3269,N_2867,N_2692);
nand U3270 (N_3270,N_2270,N_2753);
nand U3271 (N_3271,N_2789,N_2772);
xnor U3272 (N_3272,N_2313,N_2829);
xor U3273 (N_3273,N_2600,N_2718);
nor U3274 (N_3274,N_2446,N_2325);
nor U3275 (N_3275,N_2376,N_2967);
nor U3276 (N_3276,N_2650,N_2945);
nand U3277 (N_3277,N_2659,N_2877);
and U3278 (N_3278,N_2495,N_2438);
and U3279 (N_3279,N_2995,N_2617);
nand U3280 (N_3280,N_2965,N_2319);
nand U3281 (N_3281,N_2405,N_2425);
xor U3282 (N_3282,N_2856,N_2285);
or U3283 (N_3283,N_2329,N_2900);
xnor U3284 (N_3284,N_2474,N_2480);
nand U3285 (N_3285,N_2926,N_2536);
or U3286 (N_3286,N_2297,N_2972);
nor U3287 (N_3287,N_2711,N_2879);
or U3288 (N_3288,N_2679,N_2934);
and U3289 (N_3289,N_2321,N_2577);
xnor U3290 (N_3290,N_2251,N_2606);
xnor U3291 (N_3291,N_2832,N_2740);
nor U3292 (N_3292,N_2494,N_2520);
xor U3293 (N_3293,N_2786,N_2349);
and U3294 (N_3294,N_2805,N_2813);
nand U3295 (N_3295,N_2874,N_2589);
xor U3296 (N_3296,N_2453,N_2950);
or U3297 (N_3297,N_2731,N_2568);
nand U3298 (N_3298,N_2554,N_2686);
and U3299 (N_3299,N_2503,N_2303);
nand U3300 (N_3300,N_2469,N_2389);
nor U3301 (N_3301,N_2820,N_2678);
and U3302 (N_3302,N_2452,N_2611);
nor U3303 (N_3303,N_2915,N_2508);
or U3304 (N_3304,N_2523,N_2540);
xor U3305 (N_3305,N_2940,N_2620);
xnor U3306 (N_3306,N_2547,N_2713);
or U3307 (N_3307,N_2433,N_2558);
or U3308 (N_3308,N_2579,N_2583);
nand U3309 (N_3309,N_2556,N_2964);
nand U3310 (N_3310,N_2328,N_2855);
or U3311 (N_3311,N_2587,N_2401);
or U3312 (N_3312,N_2271,N_2724);
or U3313 (N_3313,N_2311,N_2748);
or U3314 (N_3314,N_2535,N_2502);
and U3315 (N_3315,N_2605,N_2581);
or U3316 (N_3316,N_2351,N_2969);
xor U3317 (N_3317,N_2800,N_2868);
xnor U3318 (N_3318,N_2388,N_2881);
nor U3319 (N_3319,N_2797,N_2749);
xnor U3320 (N_3320,N_2440,N_2402);
or U3321 (N_3321,N_2447,N_2264);
or U3322 (N_3322,N_2421,N_2970);
and U3323 (N_3323,N_2684,N_2716);
and U3324 (N_3324,N_2730,N_2273);
or U3325 (N_3325,N_2875,N_2280);
xor U3326 (N_3326,N_2597,N_2825);
and U3327 (N_3327,N_2629,N_2582);
or U3328 (N_3328,N_2436,N_2841);
nor U3329 (N_3329,N_2408,N_2537);
or U3330 (N_3330,N_2555,N_2284);
nor U3331 (N_3331,N_2660,N_2983);
xnor U3332 (N_3332,N_2999,N_2546);
and U3333 (N_3333,N_2544,N_2462);
or U3334 (N_3334,N_2636,N_2931);
xor U3335 (N_3335,N_2463,N_2689);
and U3336 (N_3336,N_2850,N_2505);
xor U3337 (N_3337,N_2747,N_2831);
xnor U3338 (N_3338,N_2618,N_2395);
xnor U3339 (N_3339,N_2809,N_2771);
and U3340 (N_3340,N_2451,N_2655);
xor U3341 (N_3341,N_2279,N_2927);
and U3342 (N_3342,N_2567,N_2262);
xnor U3343 (N_3343,N_2976,N_2387);
nor U3344 (N_3344,N_2751,N_2788);
nor U3345 (N_3345,N_2677,N_2722);
nor U3346 (N_3346,N_2381,N_2356);
or U3347 (N_3347,N_2565,N_2585);
nor U3348 (N_3348,N_2437,N_2288);
or U3349 (N_3349,N_2464,N_2541);
nand U3350 (N_3350,N_2400,N_2509);
nor U3351 (N_3351,N_2687,N_2627);
or U3352 (N_3352,N_2441,N_2750);
nand U3353 (N_3353,N_2790,N_2997);
or U3354 (N_3354,N_2869,N_2990);
or U3355 (N_3355,N_2572,N_2379);
nand U3356 (N_3356,N_2830,N_2963);
or U3357 (N_3357,N_2337,N_2371);
or U3358 (N_3358,N_2944,N_2256);
nand U3359 (N_3359,N_2714,N_2314);
xnor U3360 (N_3360,N_2613,N_2429);
xor U3361 (N_3361,N_2982,N_2455);
nand U3362 (N_3362,N_2849,N_2791);
nor U3363 (N_3363,N_2858,N_2278);
or U3364 (N_3364,N_2723,N_2908);
and U3365 (N_3365,N_2887,N_2491);
and U3366 (N_3366,N_2457,N_2519);
or U3367 (N_3367,N_2828,N_2754);
xor U3368 (N_3368,N_2593,N_2524);
or U3369 (N_3369,N_2364,N_2493);
and U3370 (N_3370,N_2761,N_2506);
nand U3371 (N_3371,N_2662,N_2295);
and U3372 (N_3372,N_2834,N_2282);
and U3373 (N_3373,N_2347,N_2954);
and U3374 (N_3374,N_2870,N_2863);
and U3375 (N_3375,N_2809,N_2749);
nor U3376 (N_3376,N_2790,N_2968);
nand U3377 (N_3377,N_2686,N_2591);
nor U3378 (N_3378,N_2937,N_2270);
xnor U3379 (N_3379,N_2896,N_2510);
nand U3380 (N_3380,N_2776,N_2838);
or U3381 (N_3381,N_2430,N_2973);
nor U3382 (N_3382,N_2577,N_2274);
xor U3383 (N_3383,N_2375,N_2346);
and U3384 (N_3384,N_2257,N_2510);
nand U3385 (N_3385,N_2683,N_2545);
and U3386 (N_3386,N_2837,N_2782);
xor U3387 (N_3387,N_2326,N_2893);
xor U3388 (N_3388,N_2499,N_2731);
nand U3389 (N_3389,N_2515,N_2703);
xor U3390 (N_3390,N_2639,N_2688);
or U3391 (N_3391,N_2927,N_2790);
nand U3392 (N_3392,N_2967,N_2466);
nand U3393 (N_3393,N_2480,N_2613);
or U3394 (N_3394,N_2504,N_2386);
and U3395 (N_3395,N_2331,N_2965);
nor U3396 (N_3396,N_2399,N_2874);
or U3397 (N_3397,N_2720,N_2357);
nand U3398 (N_3398,N_2521,N_2592);
nand U3399 (N_3399,N_2468,N_2702);
xnor U3400 (N_3400,N_2931,N_2412);
and U3401 (N_3401,N_2523,N_2726);
nor U3402 (N_3402,N_2785,N_2929);
and U3403 (N_3403,N_2309,N_2533);
xnor U3404 (N_3404,N_2815,N_2350);
and U3405 (N_3405,N_2486,N_2261);
or U3406 (N_3406,N_2453,N_2514);
xor U3407 (N_3407,N_2979,N_2539);
xnor U3408 (N_3408,N_2822,N_2872);
nor U3409 (N_3409,N_2689,N_2699);
xnor U3410 (N_3410,N_2540,N_2695);
or U3411 (N_3411,N_2850,N_2350);
xor U3412 (N_3412,N_2823,N_2491);
xor U3413 (N_3413,N_2496,N_2857);
or U3414 (N_3414,N_2617,N_2408);
nand U3415 (N_3415,N_2405,N_2995);
nor U3416 (N_3416,N_2671,N_2788);
and U3417 (N_3417,N_2866,N_2825);
nand U3418 (N_3418,N_2646,N_2655);
or U3419 (N_3419,N_2366,N_2457);
nand U3420 (N_3420,N_2946,N_2414);
nor U3421 (N_3421,N_2401,N_2361);
xor U3422 (N_3422,N_2783,N_2663);
nor U3423 (N_3423,N_2807,N_2485);
and U3424 (N_3424,N_2767,N_2359);
nor U3425 (N_3425,N_2402,N_2922);
and U3426 (N_3426,N_2828,N_2353);
xor U3427 (N_3427,N_2899,N_2574);
xor U3428 (N_3428,N_2478,N_2813);
xnor U3429 (N_3429,N_2484,N_2691);
and U3430 (N_3430,N_2593,N_2588);
nand U3431 (N_3431,N_2448,N_2376);
xor U3432 (N_3432,N_2775,N_2811);
and U3433 (N_3433,N_2997,N_2705);
nand U3434 (N_3434,N_2295,N_2290);
or U3435 (N_3435,N_2785,N_2531);
nor U3436 (N_3436,N_2801,N_2481);
nand U3437 (N_3437,N_2786,N_2735);
or U3438 (N_3438,N_2366,N_2684);
nor U3439 (N_3439,N_2902,N_2605);
or U3440 (N_3440,N_2620,N_2502);
or U3441 (N_3441,N_2585,N_2402);
or U3442 (N_3442,N_2941,N_2794);
nand U3443 (N_3443,N_2483,N_2641);
xor U3444 (N_3444,N_2719,N_2594);
xor U3445 (N_3445,N_2750,N_2965);
or U3446 (N_3446,N_2384,N_2798);
nand U3447 (N_3447,N_2905,N_2388);
xor U3448 (N_3448,N_2722,N_2624);
or U3449 (N_3449,N_2491,N_2540);
nor U3450 (N_3450,N_2510,N_2752);
xnor U3451 (N_3451,N_2334,N_2691);
or U3452 (N_3452,N_2663,N_2321);
or U3453 (N_3453,N_2370,N_2411);
or U3454 (N_3454,N_2749,N_2774);
nand U3455 (N_3455,N_2548,N_2909);
nand U3456 (N_3456,N_2336,N_2474);
nor U3457 (N_3457,N_2840,N_2450);
nand U3458 (N_3458,N_2413,N_2533);
or U3459 (N_3459,N_2254,N_2798);
xor U3460 (N_3460,N_2851,N_2278);
nor U3461 (N_3461,N_2986,N_2506);
nor U3462 (N_3462,N_2913,N_2816);
nor U3463 (N_3463,N_2357,N_2828);
and U3464 (N_3464,N_2309,N_2922);
nand U3465 (N_3465,N_2271,N_2660);
nand U3466 (N_3466,N_2715,N_2794);
and U3467 (N_3467,N_2813,N_2267);
and U3468 (N_3468,N_2728,N_2566);
or U3469 (N_3469,N_2485,N_2918);
and U3470 (N_3470,N_2285,N_2304);
nor U3471 (N_3471,N_2747,N_2629);
and U3472 (N_3472,N_2827,N_2894);
xnor U3473 (N_3473,N_2353,N_2777);
nor U3474 (N_3474,N_2525,N_2949);
and U3475 (N_3475,N_2464,N_2939);
nand U3476 (N_3476,N_2784,N_2446);
nand U3477 (N_3477,N_2924,N_2689);
nor U3478 (N_3478,N_2799,N_2566);
nor U3479 (N_3479,N_2759,N_2582);
nand U3480 (N_3480,N_2739,N_2751);
nor U3481 (N_3481,N_2649,N_2781);
xor U3482 (N_3482,N_2879,N_2516);
and U3483 (N_3483,N_2781,N_2760);
nand U3484 (N_3484,N_2328,N_2605);
nand U3485 (N_3485,N_2977,N_2452);
nand U3486 (N_3486,N_2786,N_2251);
xor U3487 (N_3487,N_2846,N_2743);
and U3488 (N_3488,N_2405,N_2270);
nand U3489 (N_3489,N_2997,N_2291);
nor U3490 (N_3490,N_2356,N_2713);
and U3491 (N_3491,N_2359,N_2817);
and U3492 (N_3492,N_2432,N_2588);
nor U3493 (N_3493,N_2890,N_2869);
xor U3494 (N_3494,N_2858,N_2495);
and U3495 (N_3495,N_2853,N_2703);
and U3496 (N_3496,N_2902,N_2479);
nand U3497 (N_3497,N_2514,N_2882);
nand U3498 (N_3498,N_2283,N_2376);
and U3499 (N_3499,N_2361,N_2581);
or U3500 (N_3500,N_2951,N_2251);
nand U3501 (N_3501,N_2404,N_2890);
nor U3502 (N_3502,N_2855,N_2798);
nand U3503 (N_3503,N_2718,N_2952);
or U3504 (N_3504,N_2281,N_2516);
nand U3505 (N_3505,N_2903,N_2957);
xnor U3506 (N_3506,N_2472,N_2415);
nand U3507 (N_3507,N_2319,N_2483);
nor U3508 (N_3508,N_2652,N_2464);
nand U3509 (N_3509,N_2418,N_2450);
nand U3510 (N_3510,N_2733,N_2825);
or U3511 (N_3511,N_2712,N_2538);
nor U3512 (N_3512,N_2552,N_2550);
xor U3513 (N_3513,N_2533,N_2596);
xnor U3514 (N_3514,N_2983,N_2526);
nor U3515 (N_3515,N_2661,N_2289);
nor U3516 (N_3516,N_2736,N_2788);
and U3517 (N_3517,N_2726,N_2472);
nand U3518 (N_3518,N_2806,N_2520);
nor U3519 (N_3519,N_2270,N_2438);
nor U3520 (N_3520,N_2574,N_2415);
nand U3521 (N_3521,N_2505,N_2650);
xnor U3522 (N_3522,N_2759,N_2346);
or U3523 (N_3523,N_2842,N_2721);
and U3524 (N_3524,N_2889,N_2724);
or U3525 (N_3525,N_2806,N_2496);
xor U3526 (N_3526,N_2254,N_2702);
nor U3527 (N_3527,N_2264,N_2836);
nor U3528 (N_3528,N_2542,N_2461);
or U3529 (N_3529,N_2696,N_2989);
xnor U3530 (N_3530,N_2251,N_2550);
or U3531 (N_3531,N_2665,N_2918);
nor U3532 (N_3532,N_2736,N_2739);
nand U3533 (N_3533,N_2620,N_2322);
and U3534 (N_3534,N_2632,N_2837);
nand U3535 (N_3535,N_2918,N_2619);
or U3536 (N_3536,N_2557,N_2755);
xor U3537 (N_3537,N_2491,N_2602);
xnor U3538 (N_3538,N_2787,N_2899);
nand U3539 (N_3539,N_2859,N_2505);
or U3540 (N_3540,N_2644,N_2438);
and U3541 (N_3541,N_2907,N_2531);
xor U3542 (N_3542,N_2976,N_2569);
nand U3543 (N_3543,N_2465,N_2307);
nand U3544 (N_3544,N_2926,N_2604);
or U3545 (N_3545,N_2793,N_2638);
nand U3546 (N_3546,N_2845,N_2369);
or U3547 (N_3547,N_2956,N_2302);
or U3548 (N_3548,N_2523,N_2664);
xnor U3549 (N_3549,N_2666,N_2756);
or U3550 (N_3550,N_2906,N_2910);
or U3551 (N_3551,N_2962,N_2500);
and U3552 (N_3552,N_2546,N_2604);
xor U3553 (N_3553,N_2656,N_2333);
nand U3554 (N_3554,N_2668,N_2920);
or U3555 (N_3555,N_2751,N_2926);
and U3556 (N_3556,N_2932,N_2966);
xnor U3557 (N_3557,N_2332,N_2259);
xor U3558 (N_3558,N_2307,N_2391);
xor U3559 (N_3559,N_2811,N_2318);
and U3560 (N_3560,N_2828,N_2410);
nor U3561 (N_3561,N_2813,N_2452);
xor U3562 (N_3562,N_2450,N_2477);
nor U3563 (N_3563,N_2349,N_2429);
nor U3564 (N_3564,N_2990,N_2693);
nor U3565 (N_3565,N_2731,N_2943);
nand U3566 (N_3566,N_2781,N_2964);
or U3567 (N_3567,N_2752,N_2887);
or U3568 (N_3568,N_2279,N_2869);
nand U3569 (N_3569,N_2430,N_2460);
nand U3570 (N_3570,N_2391,N_2354);
nor U3571 (N_3571,N_2469,N_2626);
nor U3572 (N_3572,N_2822,N_2361);
xor U3573 (N_3573,N_2948,N_2340);
and U3574 (N_3574,N_2434,N_2820);
nand U3575 (N_3575,N_2342,N_2530);
xnor U3576 (N_3576,N_2570,N_2461);
xnor U3577 (N_3577,N_2364,N_2687);
nor U3578 (N_3578,N_2411,N_2709);
nand U3579 (N_3579,N_2656,N_2686);
nor U3580 (N_3580,N_2254,N_2560);
and U3581 (N_3581,N_2428,N_2563);
and U3582 (N_3582,N_2678,N_2870);
nor U3583 (N_3583,N_2670,N_2544);
and U3584 (N_3584,N_2918,N_2773);
xnor U3585 (N_3585,N_2307,N_2999);
or U3586 (N_3586,N_2752,N_2898);
nor U3587 (N_3587,N_2804,N_2727);
and U3588 (N_3588,N_2830,N_2511);
nor U3589 (N_3589,N_2258,N_2743);
xnor U3590 (N_3590,N_2680,N_2740);
xnor U3591 (N_3591,N_2771,N_2576);
or U3592 (N_3592,N_2693,N_2955);
and U3593 (N_3593,N_2576,N_2506);
and U3594 (N_3594,N_2893,N_2636);
xnor U3595 (N_3595,N_2959,N_2517);
nor U3596 (N_3596,N_2299,N_2851);
xnor U3597 (N_3597,N_2276,N_2887);
and U3598 (N_3598,N_2660,N_2402);
or U3599 (N_3599,N_2735,N_2504);
nor U3600 (N_3600,N_2719,N_2302);
or U3601 (N_3601,N_2903,N_2704);
or U3602 (N_3602,N_2404,N_2305);
or U3603 (N_3603,N_2313,N_2748);
and U3604 (N_3604,N_2785,N_2362);
nand U3605 (N_3605,N_2868,N_2384);
or U3606 (N_3606,N_2831,N_2844);
nand U3607 (N_3607,N_2810,N_2500);
and U3608 (N_3608,N_2496,N_2596);
nand U3609 (N_3609,N_2383,N_2369);
or U3610 (N_3610,N_2309,N_2261);
nor U3611 (N_3611,N_2456,N_2749);
or U3612 (N_3612,N_2675,N_2523);
xnor U3613 (N_3613,N_2904,N_2870);
xnor U3614 (N_3614,N_2287,N_2932);
or U3615 (N_3615,N_2560,N_2983);
nand U3616 (N_3616,N_2673,N_2973);
nand U3617 (N_3617,N_2945,N_2353);
xor U3618 (N_3618,N_2550,N_2620);
xor U3619 (N_3619,N_2741,N_2727);
or U3620 (N_3620,N_2493,N_2576);
and U3621 (N_3621,N_2799,N_2931);
nor U3622 (N_3622,N_2583,N_2997);
xnor U3623 (N_3623,N_2984,N_2811);
xor U3624 (N_3624,N_2505,N_2289);
nand U3625 (N_3625,N_2443,N_2963);
and U3626 (N_3626,N_2566,N_2949);
and U3627 (N_3627,N_2828,N_2270);
nand U3628 (N_3628,N_2276,N_2849);
nand U3629 (N_3629,N_2444,N_2412);
nand U3630 (N_3630,N_2520,N_2926);
nor U3631 (N_3631,N_2705,N_2803);
nand U3632 (N_3632,N_2815,N_2914);
or U3633 (N_3633,N_2640,N_2985);
or U3634 (N_3634,N_2491,N_2364);
and U3635 (N_3635,N_2683,N_2681);
nor U3636 (N_3636,N_2576,N_2774);
or U3637 (N_3637,N_2252,N_2968);
or U3638 (N_3638,N_2358,N_2295);
nand U3639 (N_3639,N_2971,N_2849);
or U3640 (N_3640,N_2323,N_2250);
xor U3641 (N_3641,N_2694,N_2760);
nand U3642 (N_3642,N_2975,N_2389);
or U3643 (N_3643,N_2298,N_2527);
nor U3644 (N_3644,N_2636,N_2407);
and U3645 (N_3645,N_2373,N_2484);
and U3646 (N_3646,N_2501,N_2476);
and U3647 (N_3647,N_2951,N_2311);
and U3648 (N_3648,N_2864,N_2895);
and U3649 (N_3649,N_2902,N_2670);
or U3650 (N_3650,N_2894,N_2716);
or U3651 (N_3651,N_2625,N_2773);
nand U3652 (N_3652,N_2886,N_2674);
nor U3653 (N_3653,N_2798,N_2787);
xnor U3654 (N_3654,N_2457,N_2635);
or U3655 (N_3655,N_2827,N_2943);
nand U3656 (N_3656,N_2464,N_2405);
and U3657 (N_3657,N_2610,N_2960);
or U3658 (N_3658,N_2823,N_2930);
or U3659 (N_3659,N_2961,N_2276);
nand U3660 (N_3660,N_2512,N_2560);
and U3661 (N_3661,N_2474,N_2925);
or U3662 (N_3662,N_2503,N_2605);
and U3663 (N_3663,N_2377,N_2614);
nor U3664 (N_3664,N_2954,N_2416);
xnor U3665 (N_3665,N_2620,N_2574);
xor U3666 (N_3666,N_2480,N_2593);
nand U3667 (N_3667,N_2619,N_2356);
or U3668 (N_3668,N_2446,N_2833);
nand U3669 (N_3669,N_2863,N_2457);
nor U3670 (N_3670,N_2738,N_2581);
nor U3671 (N_3671,N_2252,N_2636);
xor U3672 (N_3672,N_2644,N_2302);
and U3673 (N_3673,N_2899,N_2336);
xnor U3674 (N_3674,N_2287,N_2741);
nand U3675 (N_3675,N_2398,N_2886);
xnor U3676 (N_3676,N_2671,N_2444);
xor U3677 (N_3677,N_2696,N_2495);
or U3678 (N_3678,N_2924,N_2835);
xnor U3679 (N_3679,N_2905,N_2547);
nand U3680 (N_3680,N_2699,N_2340);
nor U3681 (N_3681,N_2622,N_2678);
nand U3682 (N_3682,N_2515,N_2619);
nor U3683 (N_3683,N_2641,N_2618);
or U3684 (N_3684,N_2345,N_2593);
xor U3685 (N_3685,N_2281,N_2491);
nand U3686 (N_3686,N_2412,N_2765);
and U3687 (N_3687,N_2814,N_2963);
nor U3688 (N_3688,N_2917,N_2476);
nand U3689 (N_3689,N_2380,N_2357);
nand U3690 (N_3690,N_2361,N_2609);
or U3691 (N_3691,N_2465,N_2682);
nand U3692 (N_3692,N_2390,N_2597);
nand U3693 (N_3693,N_2720,N_2941);
and U3694 (N_3694,N_2306,N_2721);
or U3695 (N_3695,N_2277,N_2458);
nor U3696 (N_3696,N_2369,N_2969);
nor U3697 (N_3697,N_2726,N_2641);
nor U3698 (N_3698,N_2665,N_2984);
nand U3699 (N_3699,N_2530,N_2803);
xor U3700 (N_3700,N_2259,N_2869);
xor U3701 (N_3701,N_2368,N_2254);
nor U3702 (N_3702,N_2338,N_2316);
nand U3703 (N_3703,N_2536,N_2975);
or U3704 (N_3704,N_2927,N_2485);
nand U3705 (N_3705,N_2760,N_2682);
and U3706 (N_3706,N_2395,N_2261);
or U3707 (N_3707,N_2427,N_2600);
and U3708 (N_3708,N_2907,N_2673);
xnor U3709 (N_3709,N_2326,N_2739);
xor U3710 (N_3710,N_2357,N_2281);
and U3711 (N_3711,N_2784,N_2989);
nor U3712 (N_3712,N_2316,N_2255);
nand U3713 (N_3713,N_2449,N_2703);
and U3714 (N_3714,N_2899,N_2875);
nor U3715 (N_3715,N_2866,N_2597);
or U3716 (N_3716,N_2402,N_2912);
nor U3717 (N_3717,N_2581,N_2616);
or U3718 (N_3718,N_2508,N_2846);
xnor U3719 (N_3719,N_2514,N_2260);
or U3720 (N_3720,N_2756,N_2665);
or U3721 (N_3721,N_2491,N_2686);
or U3722 (N_3722,N_2328,N_2718);
nand U3723 (N_3723,N_2800,N_2752);
nor U3724 (N_3724,N_2732,N_2252);
nand U3725 (N_3725,N_2714,N_2459);
nor U3726 (N_3726,N_2291,N_2982);
xnor U3727 (N_3727,N_2811,N_2975);
xnor U3728 (N_3728,N_2453,N_2849);
and U3729 (N_3729,N_2851,N_2991);
nor U3730 (N_3730,N_2709,N_2540);
or U3731 (N_3731,N_2787,N_2435);
xnor U3732 (N_3732,N_2921,N_2266);
or U3733 (N_3733,N_2478,N_2334);
nor U3734 (N_3734,N_2545,N_2839);
or U3735 (N_3735,N_2878,N_2288);
nand U3736 (N_3736,N_2796,N_2347);
nand U3737 (N_3737,N_2632,N_2528);
nand U3738 (N_3738,N_2556,N_2368);
or U3739 (N_3739,N_2383,N_2753);
and U3740 (N_3740,N_2805,N_2303);
nor U3741 (N_3741,N_2474,N_2738);
or U3742 (N_3742,N_2272,N_2844);
xor U3743 (N_3743,N_2585,N_2322);
xor U3744 (N_3744,N_2476,N_2739);
and U3745 (N_3745,N_2848,N_2883);
or U3746 (N_3746,N_2961,N_2299);
nand U3747 (N_3747,N_2815,N_2366);
nand U3748 (N_3748,N_2411,N_2784);
xor U3749 (N_3749,N_2491,N_2935);
xor U3750 (N_3750,N_3662,N_3690);
and U3751 (N_3751,N_3578,N_3691);
nand U3752 (N_3752,N_3145,N_3537);
nand U3753 (N_3753,N_3558,N_3552);
nand U3754 (N_3754,N_3125,N_3361);
xnor U3755 (N_3755,N_3298,N_3381);
nand U3756 (N_3756,N_3417,N_3002);
and U3757 (N_3757,N_3720,N_3686);
nor U3758 (N_3758,N_3473,N_3083);
nand U3759 (N_3759,N_3626,N_3131);
nand U3760 (N_3760,N_3031,N_3744);
or U3761 (N_3761,N_3462,N_3390);
nor U3762 (N_3762,N_3664,N_3170);
nor U3763 (N_3763,N_3359,N_3114);
nor U3764 (N_3764,N_3588,N_3663);
or U3765 (N_3765,N_3240,N_3696);
nand U3766 (N_3766,N_3555,N_3583);
and U3767 (N_3767,N_3203,N_3076);
nor U3768 (N_3768,N_3709,N_3121);
and U3769 (N_3769,N_3159,N_3449);
or U3770 (N_3770,N_3331,N_3225);
or U3771 (N_3771,N_3502,N_3085);
or U3772 (N_3772,N_3737,N_3337);
and U3773 (N_3773,N_3429,N_3318);
nand U3774 (N_3774,N_3486,N_3130);
nand U3775 (N_3775,N_3579,N_3422);
xor U3776 (N_3776,N_3173,N_3183);
nand U3777 (N_3777,N_3453,N_3392);
or U3778 (N_3778,N_3053,N_3548);
nand U3779 (N_3779,N_3158,N_3250);
nor U3780 (N_3780,N_3036,N_3514);
xor U3781 (N_3781,N_3496,N_3009);
nor U3782 (N_3782,N_3202,N_3418);
and U3783 (N_3783,N_3119,N_3413);
nand U3784 (N_3784,N_3280,N_3096);
nand U3785 (N_3785,N_3373,N_3113);
and U3786 (N_3786,N_3127,N_3648);
nor U3787 (N_3787,N_3666,N_3345);
nand U3788 (N_3788,N_3168,N_3303);
or U3789 (N_3789,N_3748,N_3108);
and U3790 (N_3790,N_3556,N_3272);
or U3791 (N_3791,N_3704,N_3642);
nand U3792 (N_3792,N_3269,N_3654);
and U3793 (N_3793,N_3430,N_3024);
or U3794 (N_3794,N_3010,N_3148);
or U3795 (N_3795,N_3674,N_3103);
nor U3796 (N_3796,N_3469,N_3584);
xor U3797 (N_3797,N_3242,N_3622);
nand U3798 (N_3798,N_3695,N_3334);
nand U3799 (N_3799,N_3362,N_3068);
and U3800 (N_3800,N_3005,N_3377);
nor U3801 (N_3801,N_3197,N_3719);
nor U3802 (N_3802,N_3491,N_3100);
and U3803 (N_3803,N_3526,N_3154);
xnor U3804 (N_3804,N_3124,N_3482);
and U3805 (N_3805,N_3070,N_3027);
nor U3806 (N_3806,N_3647,N_3093);
nand U3807 (N_3807,N_3309,N_3138);
nand U3808 (N_3808,N_3435,N_3632);
and U3809 (N_3809,N_3320,N_3263);
xor U3810 (N_3810,N_3274,N_3178);
nor U3811 (N_3811,N_3290,N_3251);
nor U3812 (N_3812,N_3425,N_3445);
nand U3813 (N_3813,N_3045,N_3573);
nand U3814 (N_3814,N_3106,N_3650);
and U3815 (N_3815,N_3021,N_3658);
or U3816 (N_3816,N_3146,N_3735);
nor U3817 (N_3817,N_3593,N_3149);
nor U3818 (N_3818,N_3655,N_3079);
nor U3819 (N_3819,N_3568,N_3705);
xor U3820 (N_3820,N_3506,N_3421);
or U3821 (N_3821,N_3128,N_3505);
nand U3822 (N_3822,N_3637,N_3357);
nor U3823 (N_3823,N_3438,N_3501);
xor U3824 (N_3824,N_3388,N_3660);
and U3825 (N_3825,N_3694,N_3210);
and U3826 (N_3826,N_3039,N_3348);
or U3827 (N_3827,N_3446,N_3065);
nor U3828 (N_3828,N_3369,N_3329);
nand U3829 (N_3829,N_3325,N_3028);
or U3830 (N_3830,N_3315,N_3434);
and U3831 (N_3831,N_3199,N_3194);
xnor U3832 (N_3832,N_3101,N_3734);
nand U3833 (N_3833,N_3452,N_3166);
xor U3834 (N_3834,N_3220,N_3440);
or U3835 (N_3835,N_3094,N_3576);
nor U3836 (N_3836,N_3006,N_3436);
or U3837 (N_3837,N_3742,N_3195);
and U3838 (N_3838,N_3129,N_3466);
nor U3839 (N_3839,N_3625,N_3162);
and U3840 (N_3840,N_3447,N_3489);
nor U3841 (N_3841,N_3431,N_3545);
nand U3842 (N_3842,N_3344,N_3723);
or U3843 (N_3843,N_3456,N_3524);
or U3844 (N_3844,N_3564,N_3204);
and U3845 (N_3845,N_3547,N_3254);
and U3846 (N_3846,N_3693,N_3740);
or U3847 (N_3847,N_3287,N_3187);
xor U3848 (N_3848,N_3356,N_3400);
or U3849 (N_3849,N_3680,N_3386);
nor U3850 (N_3850,N_3364,N_3111);
or U3851 (N_3851,N_3741,N_3475);
xnor U3852 (N_3852,N_3252,N_3405);
xnor U3853 (N_3853,N_3518,N_3451);
nor U3854 (N_3854,N_3340,N_3708);
xnor U3855 (N_3855,N_3532,N_3196);
and U3856 (N_3856,N_3363,N_3351);
nand U3857 (N_3857,N_3281,N_3439);
and U3858 (N_3858,N_3126,N_3153);
and U3859 (N_3859,N_3278,N_3062);
xnor U3860 (N_3860,N_3721,N_3073);
or U3861 (N_3861,N_3627,N_3460);
nand U3862 (N_3862,N_3645,N_3619);
or U3863 (N_3863,N_3296,N_3536);
or U3864 (N_3864,N_3326,N_3087);
nor U3865 (N_3865,N_3464,N_3368);
and U3866 (N_3866,N_3732,N_3530);
nor U3867 (N_3867,N_3490,N_3268);
and U3868 (N_3868,N_3198,N_3729);
xor U3869 (N_3869,N_3415,N_3172);
and U3870 (N_3870,N_3353,N_3366);
nor U3871 (N_3871,N_3051,N_3504);
or U3872 (N_3872,N_3563,N_3285);
nand U3873 (N_3873,N_3058,N_3262);
and U3874 (N_3874,N_3015,N_3639);
xor U3875 (N_3875,N_3367,N_3712);
nor U3876 (N_3876,N_3286,N_3338);
and U3877 (N_3877,N_3008,N_3375);
or U3878 (N_3878,N_3059,N_3546);
nand U3879 (N_3879,N_3191,N_3401);
xnor U3880 (N_3880,N_3190,N_3160);
nor U3881 (N_3881,N_3284,N_3733);
and U3882 (N_3882,N_3201,N_3052);
and U3883 (N_3883,N_3683,N_3677);
nor U3884 (N_3884,N_3707,N_3410);
xor U3885 (N_3885,N_3212,N_3143);
or U3886 (N_3886,N_3617,N_3069);
xnor U3887 (N_3887,N_3403,N_3725);
and U3888 (N_3888,N_3688,N_3292);
nand U3889 (N_3889,N_3385,N_3266);
nor U3890 (N_3890,N_3597,N_3294);
or U3891 (N_3891,N_3509,N_3487);
xnor U3892 (N_3892,N_3606,N_3457);
or U3893 (N_3893,N_3595,N_3035);
xnor U3894 (N_3894,N_3300,N_3681);
nor U3895 (N_3895,N_3323,N_3739);
xor U3896 (N_3896,N_3186,N_3176);
nor U3897 (N_3897,N_3163,N_3507);
nand U3898 (N_3898,N_3221,N_3477);
xnor U3899 (N_3899,N_3480,N_3743);
and U3900 (N_3900,N_3156,N_3336);
nand U3901 (N_3901,N_3465,N_3665);
xnor U3902 (N_3902,N_3118,N_3525);
xnor U3903 (N_3903,N_3738,N_3454);
xor U3904 (N_3904,N_3311,N_3523);
or U3905 (N_3905,N_3517,N_3396);
nand U3906 (N_3906,N_3646,N_3533);
and U3907 (N_3907,N_3171,N_3048);
nand U3908 (N_3908,N_3382,N_3544);
nor U3909 (N_3909,N_3483,N_3044);
nor U3910 (N_3910,N_3378,N_3218);
nor U3911 (N_3911,N_3003,N_3569);
and U3912 (N_3912,N_3025,N_3519);
nand U3913 (N_3913,N_3253,N_3164);
and U3914 (N_3914,N_3335,N_3139);
and U3915 (N_3915,N_3342,N_3306);
and U3916 (N_3916,N_3152,N_3678);
and U3917 (N_3917,N_3217,N_3227);
nor U3918 (N_3918,N_3192,N_3511);
nor U3919 (N_3919,N_3673,N_3112);
nand U3920 (N_3920,N_3409,N_3016);
and U3921 (N_3921,N_3671,N_3142);
and U3922 (N_3922,N_3255,N_3550);
nand U3923 (N_3923,N_3245,N_3615);
or U3924 (N_3924,N_3706,N_3270);
xor U3925 (N_3925,N_3592,N_3535);
and U3926 (N_3926,N_3672,N_3497);
and U3927 (N_3927,N_3324,N_3060);
or U3928 (N_3928,N_3468,N_3554);
nor U3929 (N_3929,N_3596,N_3582);
and U3930 (N_3930,N_3717,N_3161);
nor U3931 (N_3931,N_3084,N_3577);
xnor U3932 (N_3932,N_3656,N_3551);
xor U3933 (N_3933,N_3267,N_3107);
and U3934 (N_3934,N_3703,N_3437);
or U3935 (N_3935,N_3557,N_3034);
nor U3936 (N_3936,N_3692,N_3715);
or U3937 (N_3937,N_3398,N_3589);
nand U3938 (N_3938,N_3040,N_3264);
nor U3939 (N_3939,N_3310,N_3301);
nor U3940 (N_3940,N_3246,N_3249);
nor U3941 (N_3941,N_3317,N_3455);
and U3942 (N_3942,N_3104,N_3167);
nand U3943 (N_3943,N_3638,N_3071);
nand U3944 (N_3944,N_3416,N_3177);
nor U3945 (N_3945,N_3207,N_3007);
and U3946 (N_3946,N_3488,N_3222);
xnor U3947 (N_3947,N_3586,N_3304);
nor U3948 (N_3948,N_3718,N_3132);
xor U3949 (N_3949,N_3443,N_3393);
or U3950 (N_3950,N_3411,N_3319);
nor U3951 (N_3951,N_3327,N_3470);
and U3952 (N_3952,N_3243,N_3219);
nand U3953 (N_3953,N_3407,N_3463);
xor U3954 (N_3954,N_3391,N_3432);
nand U3955 (N_3955,N_3591,N_3105);
and U3956 (N_3956,N_3669,N_3374);
or U3957 (N_3957,N_3259,N_3580);
or U3958 (N_3958,N_3376,N_3587);
nand U3959 (N_3959,N_3116,N_3046);
nand U3960 (N_3960,N_3231,N_3200);
and U3961 (N_3961,N_3621,N_3360);
xnor U3962 (N_3962,N_3384,N_3056);
xnor U3963 (N_3963,N_3305,N_3698);
and U3964 (N_3964,N_3140,N_3448);
or U3965 (N_3965,N_3063,N_3276);
and U3966 (N_3966,N_3258,N_3150);
or U3967 (N_3967,N_3019,N_3566);
nor U3968 (N_3968,N_3630,N_3636);
xor U3969 (N_3969,N_3022,N_3684);
nor U3970 (N_3970,N_3239,N_3283);
nand U3971 (N_3971,N_3610,N_3608);
and U3972 (N_3972,N_3018,N_3102);
nand U3973 (N_3973,N_3237,N_3075);
nand U3974 (N_3974,N_3224,N_3313);
or U3975 (N_3975,N_3498,N_3540);
and U3976 (N_3976,N_3289,N_3408);
xnor U3977 (N_3977,N_3001,N_3601);
and U3978 (N_3978,N_3749,N_3110);
and U3979 (N_3979,N_3653,N_3609);
xnor U3980 (N_3980,N_3134,N_3371);
or U3981 (N_3981,N_3082,N_3080);
or U3982 (N_3982,N_3341,N_3122);
nand U3983 (N_3983,N_3061,N_3144);
nand U3984 (N_3984,N_3716,N_3676);
or U3985 (N_3985,N_3029,N_3412);
or U3986 (N_3986,N_3299,N_3330);
nor U3987 (N_3987,N_3241,N_3643);
nor U3988 (N_3988,N_3529,N_3157);
nor U3989 (N_3989,N_3141,N_3321);
and U3990 (N_3990,N_3179,N_3618);
or U3991 (N_3991,N_3273,N_3699);
or U3992 (N_3992,N_3492,N_3604);
nand U3993 (N_3993,N_3380,N_3521);
or U3994 (N_3994,N_3049,N_3092);
and U3995 (N_3995,N_3649,N_3599);
nand U3996 (N_3996,N_3616,N_3339);
xnor U3997 (N_3997,N_3495,N_3520);
nand U3998 (N_3998,N_3020,N_3476);
xnor U3999 (N_3999,N_3651,N_3510);
nor U4000 (N_4000,N_3097,N_3135);
and U4001 (N_4001,N_3215,N_3038);
nand U4002 (N_4002,N_3667,N_3090);
xor U4003 (N_4003,N_3074,N_3508);
or U4004 (N_4004,N_3117,N_3624);
xor U4005 (N_4005,N_3328,N_3343);
nor U4006 (N_4006,N_3346,N_3333);
or U4007 (N_4007,N_3561,N_3355);
nand U4008 (N_4008,N_3426,N_3553);
xor U4009 (N_4009,N_3037,N_3472);
nand U4010 (N_4010,N_3644,N_3700);
nand U4011 (N_4011,N_3030,N_3017);
nor U4012 (N_4012,N_3394,N_3590);
and U4013 (N_4013,N_3011,N_3572);
or U4014 (N_4014,N_3032,N_3728);
nand U4015 (N_4015,N_3257,N_3297);
nor U4016 (N_4016,N_3613,N_3098);
or U4017 (N_4017,N_3628,N_3047);
nor U4018 (N_4018,N_3151,N_3226);
xor U4019 (N_4019,N_3261,N_3668);
and U4020 (N_4020,N_3652,N_3614);
nor U4021 (N_4021,N_3275,N_3516);
nor U4022 (N_4022,N_3659,N_3133);
or U4023 (N_4023,N_3347,N_3594);
and U4024 (N_4024,N_3088,N_3531);
nand U4025 (N_4025,N_3541,N_3685);
nor U4026 (N_4026,N_3670,N_3538);
xnor U4027 (N_4027,N_3387,N_3216);
or U4028 (N_4028,N_3598,N_3174);
xor U4029 (N_4029,N_3354,N_3657);
or U4030 (N_4030,N_3066,N_3302);
or U4031 (N_4031,N_3585,N_3050);
or U4032 (N_4032,N_3295,N_3099);
xor U4033 (N_4033,N_3562,N_3383);
nand U4034 (N_4034,N_3205,N_3014);
or U4035 (N_4035,N_3389,N_3077);
nor U4036 (N_4036,N_3235,N_3746);
nand U4037 (N_4037,N_3442,N_3702);
nor U4038 (N_4038,N_3402,N_3713);
nand U4039 (N_4039,N_3461,N_3370);
and U4040 (N_4040,N_3000,N_3542);
nor U4041 (N_4041,N_3322,N_3679);
nor U4042 (N_4042,N_3120,N_3155);
xor U4043 (N_4043,N_3682,N_3033);
xnor U4044 (N_4044,N_3730,N_3701);
nand U4045 (N_4045,N_3500,N_3271);
nor U4046 (N_4046,N_3549,N_3689);
xnor U4047 (N_4047,N_3697,N_3232);
nor U4048 (N_4048,N_3528,N_3265);
or U4049 (N_4049,N_3372,N_3213);
nor U4050 (N_4050,N_3406,N_3623);
xor U4051 (N_4051,N_3042,N_3395);
or U4052 (N_4052,N_3567,N_3640);
nand U4053 (N_4053,N_3414,N_3620);
or U4054 (N_4054,N_3710,N_3137);
nor U4055 (N_4055,N_3208,N_3420);
or U4056 (N_4056,N_3123,N_3012);
and U4057 (N_4057,N_3067,N_3474);
nand U4058 (N_4058,N_3184,N_3248);
nand U4059 (N_4059,N_3358,N_3189);
and U4060 (N_4060,N_3404,N_3481);
xor U4061 (N_4061,N_3316,N_3726);
nor U4062 (N_4062,N_3223,N_3458);
nor U4063 (N_4063,N_3234,N_3629);
or U4064 (N_4064,N_3419,N_3054);
and U4065 (N_4065,N_3236,N_3169);
xnor U4066 (N_4066,N_3399,N_3570);
xnor U4067 (N_4067,N_3424,N_3043);
or U4068 (N_4068,N_3057,N_3352);
and U4069 (N_4069,N_3308,N_3428);
xor U4070 (N_4070,N_3513,N_3312);
xnor U4071 (N_4071,N_3332,N_3745);
and U4072 (N_4072,N_3727,N_3379);
nand U4073 (N_4073,N_3293,N_3165);
nand U4074 (N_4074,N_3247,N_3288);
nand U4075 (N_4075,N_3041,N_3013);
xnor U4076 (N_4076,N_3349,N_3484);
and U4077 (N_4077,N_3602,N_3499);
xnor U4078 (N_4078,N_3055,N_3314);
or U4079 (N_4079,N_3147,N_3479);
nor U4080 (N_4080,N_3095,N_3136);
nand U4081 (N_4081,N_3365,N_3115);
nand U4082 (N_4082,N_3444,N_3605);
nand U4083 (N_4083,N_3214,N_3023);
xnor U4084 (N_4084,N_3291,N_3209);
or U4085 (N_4085,N_3467,N_3233);
and U4086 (N_4086,N_3731,N_3450);
or U4087 (N_4087,N_3091,N_3560);
nand U4088 (N_4088,N_3635,N_3634);
or U4089 (N_4089,N_3277,N_3724);
nand U4090 (N_4090,N_3575,N_3722);
and U4091 (N_4091,N_3175,N_3185);
and U4092 (N_4092,N_3109,N_3687);
and U4093 (N_4093,N_3279,N_3675);
nor U4094 (N_4094,N_3559,N_3512);
xnor U4095 (N_4095,N_3534,N_3072);
nand U4096 (N_4096,N_3747,N_3397);
xnor U4097 (N_4097,N_3527,N_3641);
nand U4098 (N_4098,N_3503,N_3571);
xor U4099 (N_4099,N_3607,N_3565);
or U4100 (N_4100,N_3064,N_3736);
nand U4101 (N_4101,N_3350,N_3193);
xnor U4102 (N_4102,N_3229,N_3433);
xor U4103 (N_4103,N_3260,N_3244);
nand U4104 (N_4104,N_3004,N_3307);
nor U4105 (N_4105,N_3600,N_3282);
xor U4106 (N_4106,N_3515,N_3493);
xor U4107 (N_4107,N_3543,N_3574);
nand U4108 (N_4108,N_3441,N_3423);
or U4109 (N_4109,N_3539,N_3611);
nor U4110 (N_4110,N_3256,N_3459);
nor U4111 (N_4111,N_3471,N_3714);
nand U4112 (N_4112,N_3182,N_3228);
nand U4113 (N_4113,N_3181,N_3494);
nand U4114 (N_4114,N_3026,N_3485);
nor U4115 (N_4115,N_3081,N_3603);
and U4116 (N_4116,N_3180,N_3633);
nand U4117 (N_4117,N_3631,N_3206);
and U4118 (N_4118,N_3661,N_3086);
nand U4119 (N_4119,N_3522,N_3089);
nand U4120 (N_4120,N_3711,N_3478);
nor U4121 (N_4121,N_3211,N_3230);
nand U4122 (N_4122,N_3078,N_3188);
nor U4123 (N_4123,N_3612,N_3427);
nand U4124 (N_4124,N_3581,N_3238);
nand U4125 (N_4125,N_3181,N_3042);
nor U4126 (N_4126,N_3593,N_3053);
or U4127 (N_4127,N_3074,N_3448);
xnor U4128 (N_4128,N_3120,N_3439);
nand U4129 (N_4129,N_3126,N_3491);
and U4130 (N_4130,N_3736,N_3337);
nand U4131 (N_4131,N_3711,N_3601);
and U4132 (N_4132,N_3110,N_3085);
or U4133 (N_4133,N_3664,N_3168);
nor U4134 (N_4134,N_3105,N_3564);
xor U4135 (N_4135,N_3212,N_3442);
or U4136 (N_4136,N_3046,N_3190);
nor U4137 (N_4137,N_3111,N_3443);
nand U4138 (N_4138,N_3654,N_3409);
xor U4139 (N_4139,N_3675,N_3097);
or U4140 (N_4140,N_3540,N_3198);
and U4141 (N_4141,N_3736,N_3054);
or U4142 (N_4142,N_3356,N_3699);
or U4143 (N_4143,N_3704,N_3076);
nand U4144 (N_4144,N_3310,N_3630);
and U4145 (N_4145,N_3109,N_3294);
or U4146 (N_4146,N_3739,N_3097);
xor U4147 (N_4147,N_3591,N_3130);
xnor U4148 (N_4148,N_3220,N_3407);
and U4149 (N_4149,N_3699,N_3611);
or U4150 (N_4150,N_3504,N_3622);
and U4151 (N_4151,N_3630,N_3500);
nand U4152 (N_4152,N_3081,N_3408);
or U4153 (N_4153,N_3098,N_3201);
nor U4154 (N_4154,N_3563,N_3602);
nand U4155 (N_4155,N_3272,N_3693);
xnor U4156 (N_4156,N_3063,N_3191);
or U4157 (N_4157,N_3304,N_3294);
xnor U4158 (N_4158,N_3438,N_3516);
xnor U4159 (N_4159,N_3509,N_3093);
nor U4160 (N_4160,N_3038,N_3302);
xor U4161 (N_4161,N_3678,N_3325);
xnor U4162 (N_4162,N_3420,N_3183);
nor U4163 (N_4163,N_3570,N_3376);
nor U4164 (N_4164,N_3045,N_3489);
nand U4165 (N_4165,N_3336,N_3618);
or U4166 (N_4166,N_3410,N_3506);
or U4167 (N_4167,N_3538,N_3444);
nand U4168 (N_4168,N_3264,N_3429);
or U4169 (N_4169,N_3524,N_3299);
and U4170 (N_4170,N_3591,N_3048);
nand U4171 (N_4171,N_3464,N_3592);
xnor U4172 (N_4172,N_3730,N_3454);
xnor U4173 (N_4173,N_3220,N_3138);
xnor U4174 (N_4174,N_3194,N_3320);
nand U4175 (N_4175,N_3500,N_3269);
xnor U4176 (N_4176,N_3727,N_3031);
and U4177 (N_4177,N_3076,N_3129);
and U4178 (N_4178,N_3141,N_3249);
xnor U4179 (N_4179,N_3528,N_3405);
nor U4180 (N_4180,N_3295,N_3533);
xnor U4181 (N_4181,N_3218,N_3671);
xnor U4182 (N_4182,N_3735,N_3315);
nand U4183 (N_4183,N_3735,N_3232);
and U4184 (N_4184,N_3256,N_3351);
nand U4185 (N_4185,N_3563,N_3420);
and U4186 (N_4186,N_3409,N_3175);
and U4187 (N_4187,N_3077,N_3484);
or U4188 (N_4188,N_3339,N_3670);
and U4189 (N_4189,N_3024,N_3154);
and U4190 (N_4190,N_3460,N_3515);
xor U4191 (N_4191,N_3215,N_3730);
nand U4192 (N_4192,N_3236,N_3057);
nor U4193 (N_4193,N_3324,N_3485);
nand U4194 (N_4194,N_3714,N_3432);
xnor U4195 (N_4195,N_3191,N_3093);
or U4196 (N_4196,N_3170,N_3745);
and U4197 (N_4197,N_3156,N_3196);
or U4198 (N_4198,N_3552,N_3159);
and U4199 (N_4199,N_3632,N_3495);
nand U4200 (N_4200,N_3494,N_3735);
or U4201 (N_4201,N_3321,N_3458);
xnor U4202 (N_4202,N_3180,N_3108);
and U4203 (N_4203,N_3675,N_3074);
or U4204 (N_4204,N_3268,N_3591);
and U4205 (N_4205,N_3595,N_3110);
or U4206 (N_4206,N_3532,N_3602);
and U4207 (N_4207,N_3535,N_3562);
nand U4208 (N_4208,N_3489,N_3415);
and U4209 (N_4209,N_3306,N_3637);
and U4210 (N_4210,N_3684,N_3361);
xor U4211 (N_4211,N_3506,N_3701);
or U4212 (N_4212,N_3430,N_3544);
or U4213 (N_4213,N_3278,N_3031);
nor U4214 (N_4214,N_3710,N_3359);
or U4215 (N_4215,N_3675,N_3217);
nand U4216 (N_4216,N_3572,N_3229);
xor U4217 (N_4217,N_3038,N_3441);
nand U4218 (N_4218,N_3427,N_3123);
and U4219 (N_4219,N_3236,N_3729);
nor U4220 (N_4220,N_3499,N_3551);
and U4221 (N_4221,N_3552,N_3704);
nor U4222 (N_4222,N_3191,N_3263);
xnor U4223 (N_4223,N_3273,N_3339);
xor U4224 (N_4224,N_3346,N_3001);
xor U4225 (N_4225,N_3544,N_3375);
nand U4226 (N_4226,N_3439,N_3270);
and U4227 (N_4227,N_3724,N_3092);
xor U4228 (N_4228,N_3273,N_3716);
and U4229 (N_4229,N_3540,N_3136);
nor U4230 (N_4230,N_3662,N_3483);
xor U4231 (N_4231,N_3630,N_3323);
xnor U4232 (N_4232,N_3312,N_3656);
xnor U4233 (N_4233,N_3714,N_3620);
xor U4234 (N_4234,N_3216,N_3401);
nor U4235 (N_4235,N_3264,N_3500);
xor U4236 (N_4236,N_3028,N_3350);
xnor U4237 (N_4237,N_3386,N_3149);
xor U4238 (N_4238,N_3171,N_3075);
nand U4239 (N_4239,N_3589,N_3743);
and U4240 (N_4240,N_3631,N_3606);
nor U4241 (N_4241,N_3054,N_3567);
nor U4242 (N_4242,N_3209,N_3556);
xor U4243 (N_4243,N_3030,N_3011);
nand U4244 (N_4244,N_3563,N_3132);
nand U4245 (N_4245,N_3385,N_3517);
nand U4246 (N_4246,N_3518,N_3101);
nand U4247 (N_4247,N_3739,N_3188);
nand U4248 (N_4248,N_3078,N_3211);
xnor U4249 (N_4249,N_3411,N_3420);
nor U4250 (N_4250,N_3199,N_3587);
or U4251 (N_4251,N_3235,N_3674);
nand U4252 (N_4252,N_3393,N_3591);
and U4253 (N_4253,N_3566,N_3039);
nand U4254 (N_4254,N_3705,N_3572);
and U4255 (N_4255,N_3128,N_3065);
nand U4256 (N_4256,N_3180,N_3432);
nand U4257 (N_4257,N_3539,N_3716);
nand U4258 (N_4258,N_3515,N_3748);
xnor U4259 (N_4259,N_3732,N_3308);
nand U4260 (N_4260,N_3169,N_3251);
nor U4261 (N_4261,N_3308,N_3368);
nor U4262 (N_4262,N_3276,N_3082);
nand U4263 (N_4263,N_3370,N_3540);
nand U4264 (N_4264,N_3295,N_3371);
or U4265 (N_4265,N_3136,N_3386);
or U4266 (N_4266,N_3289,N_3643);
nand U4267 (N_4267,N_3738,N_3078);
nor U4268 (N_4268,N_3742,N_3467);
nor U4269 (N_4269,N_3220,N_3014);
xor U4270 (N_4270,N_3167,N_3644);
nand U4271 (N_4271,N_3631,N_3282);
nand U4272 (N_4272,N_3583,N_3572);
or U4273 (N_4273,N_3322,N_3018);
nor U4274 (N_4274,N_3001,N_3283);
nand U4275 (N_4275,N_3674,N_3553);
xor U4276 (N_4276,N_3518,N_3314);
xor U4277 (N_4277,N_3161,N_3504);
xor U4278 (N_4278,N_3012,N_3269);
nand U4279 (N_4279,N_3570,N_3026);
and U4280 (N_4280,N_3267,N_3699);
nor U4281 (N_4281,N_3292,N_3536);
and U4282 (N_4282,N_3729,N_3131);
nand U4283 (N_4283,N_3002,N_3335);
and U4284 (N_4284,N_3675,N_3019);
xnor U4285 (N_4285,N_3321,N_3048);
or U4286 (N_4286,N_3229,N_3317);
nor U4287 (N_4287,N_3571,N_3637);
nand U4288 (N_4288,N_3205,N_3405);
or U4289 (N_4289,N_3438,N_3413);
and U4290 (N_4290,N_3347,N_3306);
nand U4291 (N_4291,N_3157,N_3472);
nand U4292 (N_4292,N_3309,N_3041);
and U4293 (N_4293,N_3553,N_3218);
nor U4294 (N_4294,N_3264,N_3062);
and U4295 (N_4295,N_3004,N_3414);
or U4296 (N_4296,N_3536,N_3225);
nand U4297 (N_4297,N_3674,N_3558);
nand U4298 (N_4298,N_3702,N_3545);
nor U4299 (N_4299,N_3169,N_3321);
nor U4300 (N_4300,N_3158,N_3486);
xnor U4301 (N_4301,N_3432,N_3211);
or U4302 (N_4302,N_3156,N_3449);
nor U4303 (N_4303,N_3634,N_3316);
nand U4304 (N_4304,N_3201,N_3401);
and U4305 (N_4305,N_3269,N_3746);
nand U4306 (N_4306,N_3401,N_3659);
nor U4307 (N_4307,N_3492,N_3728);
or U4308 (N_4308,N_3191,N_3111);
nor U4309 (N_4309,N_3604,N_3175);
or U4310 (N_4310,N_3204,N_3342);
xnor U4311 (N_4311,N_3062,N_3747);
nand U4312 (N_4312,N_3560,N_3040);
xnor U4313 (N_4313,N_3107,N_3052);
nand U4314 (N_4314,N_3120,N_3187);
and U4315 (N_4315,N_3657,N_3424);
nor U4316 (N_4316,N_3457,N_3421);
or U4317 (N_4317,N_3503,N_3403);
or U4318 (N_4318,N_3544,N_3012);
xnor U4319 (N_4319,N_3376,N_3647);
and U4320 (N_4320,N_3321,N_3311);
nand U4321 (N_4321,N_3699,N_3270);
nand U4322 (N_4322,N_3658,N_3569);
xnor U4323 (N_4323,N_3513,N_3350);
and U4324 (N_4324,N_3745,N_3659);
or U4325 (N_4325,N_3440,N_3377);
or U4326 (N_4326,N_3580,N_3330);
and U4327 (N_4327,N_3581,N_3685);
xor U4328 (N_4328,N_3091,N_3510);
or U4329 (N_4329,N_3563,N_3043);
or U4330 (N_4330,N_3450,N_3324);
nand U4331 (N_4331,N_3092,N_3719);
and U4332 (N_4332,N_3663,N_3277);
nor U4333 (N_4333,N_3611,N_3558);
xnor U4334 (N_4334,N_3643,N_3521);
nand U4335 (N_4335,N_3330,N_3389);
nor U4336 (N_4336,N_3058,N_3260);
or U4337 (N_4337,N_3372,N_3190);
nor U4338 (N_4338,N_3562,N_3071);
nand U4339 (N_4339,N_3507,N_3272);
nand U4340 (N_4340,N_3523,N_3066);
nor U4341 (N_4341,N_3664,N_3563);
nand U4342 (N_4342,N_3688,N_3277);
nand U4343 (N_4343,N_3293,N_3002);
nand U4344 (N_4344,N_3288,N_3573);
or U4345 (N_4345,N_3691,N_3018);
nor U4346 (N_4346,N_3736,N_3235);
or U4347 (N_4347,N_3167,N_3049);
nor U4348 (N_4348,N_3319,N_3653);
xnor U4349 (N_4349,N_3260,N_3487);
xor U4350 (N_4350,N_3519,N_3343);
and U4351 (N_4351,N_3727,N_3504);
or U4352 (N_4352,N_3587,N_3063);
and U4353 (N_4353,N_3412,N_3381);
or U4354 (N_4354,N_3594,N_3522);
and U4355 (N_4355,N_3291,N_3610);
and U4356 (N_4356,N_3406,N_3440);
and U4357 (N_4357,N_3561,N_3316);
xor U4358 (N_4358,N_3211,N_3075);
nand U4359 (N_4359,N_3650,N_3285);
xor U4360 (N_4360,N_3384,N_3044);
xor U4361 (N_4361,N_3546,N_3224);
xnor U4362 (N_4362,N_3640,N_3649);
nor U4363 (N_4363,N_3612,N_3738);
nor U4364 (N_4364,N_3479,N_3197);
or U4365 (N_4365,N_3118,N_3002);
nor U4366 (N_4366,N_3335,N_3186);
nor U4367 (N_4367,N_3654,N_3344);
nor U4368 (N_4368,N_3403,N_3623);
xnor U4369 (N_4369,N_3208,N_3328);
xor U4370 (N_4370,N_3525,N_3713);
xor U4371 (N_4371,N_3072,N_3531);
nand U4372 (N_4372,N_3267,N_3662);
nand U4373 (N_4373,N_3437,N_3720);
nor U4374 (N_4374,N_3230,N_3423);
and U4375 (N_4375,N_3084,N_3504);
nor U4376 (N_4376,N_3324,N_3666);
nand U4377 (N_4377,N_3193,N_3471);
or U4378 (N_4378,N_3355,N_3153);
xor U4379 (N_4379,N_3078,N_3256);
and U4380 (N_4380,N_3416,N_3202);
xnor U4381 (N_4381,N_3235,N_3387);
and U4382 (N_4382,N_3399,N_3723);
and U4383 (N_4383,N_3097,N_3497);
xnor U4384 (N_4384,N_3637,N_3711);
and U4385 (N_4385,N_3031,N_3011);
nor U4386 (N_4386,N_3219,N_3559);
and U4387 (N_4387,N_3634,N_3036);
or U4388 (N_4388,N_3450,N_3574);
nand U4389 (N_4389,N_3706,N_3282);
or U4390 (N_4390,N_3299,N_3156);
nand U4391 (N_4391,N_3041,N_3712);
or U4392 (N_4392,N_3747,N_3542);
and U4393 (N_4393,N_3345,N_3046);
and U4394 (N_4394,N_3367,N_3528);
nor U4395 (N_4395,N_3064,N_3192);
xnor U4396 (N_4396,N_3623,N_3706);
or U4397 (N_4397,N_3031,N_3125);
or U4398 (N_4398,N_3687,N_3147);
xor U4399 (N_4399,N_3358,N_3701);
xor U4400 (N_4400,N_3127,N_3084);
or U4401 (N_4401,N_3370,N_3157);
or U4402 (N_4402,N_3617,N_3171);
nand U4403 (N_4403,N_3292,N_3378);
nor U4404 (N_4404,N_3276,N_3674);
xnor U4405 (N_4405,N_3566,N_3264);
and U4406 (N_4406,N_3695,N_3266);
xor U4407 (N_4407,N_3150,N_3226);
or U4408 (N_4408,N_3518,N_3433);
nor U4409 (N_4409,N_3742,N_3648);
nor U4410 (N_4410,N_3083,N_3087);
or U4411 (N_4411,N_3398,N_3579);
xnor U4412 (N_4412,N_3735,N_3518);
or U4413 (N_4413,N_3286,N_3014);
xnor U4414 (N_4414,N_3353,N_3411);
nand U4415 (N_4415,N_3135,N_3447);
nand U4416 (N_4416,N_3348,N_3489);
or U4417 (N_4417,N_3352,N_3691);
nand U4418 (N_4418,N_3208,N_3462);
and U4419 (N_4419,N_3221,N_3103);
nand U4420 (N_4420,N_3189,N_3036);
and U4421 (N_4421,N_3260,N_3546);
nand U4422 (N_4422,N_3533,N_3220);
nor U4423 (N_4423,N_3379,N_3586);
or U4424 (N_4424,N_3029,N_3219);
nand U4425 (N_4425,N_3229,N_3365);
xnor U4426 (N_4426,N_3583,N_3620);
nor U4427 (N_4427,N_3526,N_3344);
nand U4428 (N_4428,N_3710,N_3525);
and U4429 (N_4429,N_3052,N_3194);
xor U4430 (N_4430,N_3054,N_3479);
xnor U4431 (N_4431,N_3332,N_3235);
xnor U4432 (N_4432,N_3603,N_3452);
nand U4433 (N_4433,N_3522,N_3263);
nor U4434 (N_4434,N_3583,N_3632);
nand U4435 (N_4435,N_3258,N_3520);
and U4436 (N_4436,N_3161,N_3108);
nand U4437 (N_4437,N_3143,N_3009);
and U4438 (N_4438,N_3047,N_3343);
nand U4439 (N_4439,N_3068,N_3330);
or U4440 (N_4440,N_3078,N_3178);
and U4441 (N_4441,N_3497,N_3526);
nand U4442 (N_4442,N_3214,N_3039);
xnor U4443 (N_4443,N_3268,N_3714);
xnor U4444 (N_4444,N_3391,N_3533);
nand U4445 (N_4445,N_3522,N_3247);
or U4446 (N_4446,N_3335,N_3136);
xnor U4447 (N_4447,N_3569,N_3273);
and U4448 (N_4448,N_3654,N_3611);
nor U4449 (N_4449,N_3458,N_3577);
nand U4450 (N_4450,N_3374,N_3296);
xor U4451 (N_4451,N_3713,N_3702);
or U4452 (N_4452,N_3008,N_3160);
nor U4453 (N_4453,N_3632,N_3129);
and U4454 (N_4454,N_3097,N_3449);
xor U4455 (N_4455,N_3265,N_3214);
nand U4456 (N_4456,N_3186,N_3130);
nor U4457 (N_4457,N_3672,N_3552);
or U4458 (N_4458,N_3111,N_3530);
and U4459 (N_4459,N_3593,N_3403);
and U4460 (N_4460,N_3660,N_3276);
or U4461 (N_4461,N_3511,N_3461);
or U4462 (N_4462,N_3221,N_3597);
nand U4463 (N_4463,N_3519,N_3065);
nand U4464 (N_4464,N_3204,N_3572);
and U4465 (N_4465,N_3076,N_3064);
nand U4466 (N_4466,N_3565,N_3064);
nor U4467 (N_4467,N_3129,N_3335);
xnor U4468 (N_4468,N_3739,N_3001);
or U4469 (N_4469,N_3665,N_3170);
nor U4470 (N_4470,N_3193,N_3570);
nor U4471 (N_4471,N_3609,N_3746);
xor U4472 (N_4472,N_3003,N_3731);
nand U4473 (N_4473,N_3067,N_3096);
or U4474 (N_4474,N_3205,N_3277);
nor U4475 (N_4475,N_3330,N_3691);
xor U4476 (N_4476,N_3281,N_3017);
nor U4477 (N_4477,N_3216,N_3262);
xor U4478 (N_4478,N_3309,N_3516);
or U4479 (N_4479,N_3225,N_3097);
or U4480 (N_4480,N_3347,N_3178);
xnor U4481 (N_4481,N_3578,N_3617);
nand U4482 (N_4482,N_3689,N_3114);
xnor U4483 (N_4483,N_3533,N_3317);
or U4484 (N_4484,N_3539,N_3418);
or U4485 (N_4485,N_3287,N_3679);
and U4486 (N_4486,N_3129,N_3036);
nand U4487 (N_4487,N_3557,N_3575);
or U4488 (N_4488,N_3561,N_3144);
and U4489 (N_4489,N_3743,N_3103);
and U4490 (N_4490,N_3434,N_3330);
or U4491 (N_4491,N_3145,N_3156);
and U4492 (N_4492,N_3344,N_3237);
nor U4493 (N_4493,N_3200,N_3435);
or U4494 (N_4494,N_3362,N_3005);
nor U4495 (N_4495,N_3223,N_3529);
nand U4496 (N_4496,N_3518,N_3726);
xnor U4497 (N_4497,N_3520,N_3170);
nand U4498 (N_4498,N_3040,N_3170);
or U4499 (N_4499,N_3132,N_3129);
nand U4500 (N_4500,N_3842,N_3789);
nand U4501 (N_4501,N_3763,N_4435);
nand U4502 (N_4502,N_3801,N_4432);
xor U4503 (N_4503,N_4447,N_3890);
nor U4504 (N_4504,N_3930,N_4354);
and U4505 (N_4505,N_4442,N_4171);
and U4506 (N_4506,N_4455,N_3822);
nand U4507 (N_4507,N_4034,N_3971);
nand U4508 (N_4508,N_3935,N_4230);
nor U4509 (N_4509,N_4199,N_4293);
and U4510 (N_4510,N_3885,N_4357);
or U4511 (N_4511,N_3876,N_3802);
and U4512 (N_4512,N_3828,N_4499);
and U4513 (N_4513,N_4489,N_4225);
or U4514 (N_4514,N_4267,N_4345);
xnor U4515 (N_4515,N_4468,N_4166);
nor U4516 (N_4516,N_4061,N_4071);
and U4517 (N_4517,N_3823,N_4042);
and U4518 (N_4518,N_3754,N_4215);
xor U4519 (N_4519,N_4223,N_3899);
or U4520 (N_4520,N_4309,N_4219);
nor U4521 (N_4521,N_3979,N_4367);
nor U4522 (N_4522,N_4068,N_4207);
xnor U4523 (N_4523,N_4399,N_4317);
xnor U4524 (N_4524,N_3922,N_4114);
and U4525 (N_4525,N_3883,N_3829);
or U4526 (N_4526,N_4433,N_3755);
and U4527 (N_4527,N_3938,N_3837);
xnor U4528 (N_4528,N_3900,N_3927);
and U4529 (N_4529,N_4465,N_4056);
nand U4530 (N_4530,N_4291,N_4406);
and U4531 (N_4531,N_4319,N_4244);
nor U4532 (N_4532,N_4161,N_4281);
and U4533 (N_4533,N_4402,N_4364);
nor U4534 (N_4534,N_3811,N_4213);
nand U4535 (N_4535,N_3821,N_4057);
and U4536 (N_4536,N_4492,N_3894);
xor U4537 (N_4537,N_4023,N_3879);
or U4538 (N_4538,N_3806,N_4016);
or U4539 (N_4539,N_4386,N_4158);
and U4540 (N_4540,N_4132,N_3937);
or U4541 (N_4541,N_3870,N_3907);
nand U4542 (N_4542,N_3924,N_3785);
nor U4543 (N_4543,N_4180,N_4106);
nor U4544 (N_4544,N_4024,N_3882);
nor U4545 (N_4545,N_4005,N_4390);
and U4546 (N_4546,N_3774,N_3861);
or U4547 (N_4547,N_3949,N_3803);
xnor U4548 (N_4548,N_4141,N_3758);
xor U4549 (N_4549,N_4487,N_3839);
nand U4550 (N_4550,N_4082,N_4113);
xor U4551 (N_4551,N_4064,N_3926);
nor U4552 (N_4552,N_4418,N_3916);
or U4553 (N_4553,N_4466,N_4160);
or U4554 (N_4554,N_4077,N_4246);
nor U4555 (N_4555,N_4374,N_3799);
nor U4556 (N_4556,N_4012,N_4181);
and U4557 (N_4557,N_3810,N_4471);
and U4558 (N_4558,N_4325,N_3874);
or U4559 (N_4559,N_3901,N_3860);
and U4560 (N_4560,N_4192,N_4209);
and U4561 (N_4561,N_4131,N_4172);
nand U4562 (N_4562,N_4051,N_3939);
and U4563 (N_4563,N_4282,N_4065);
xor U4564 (N_4564,N_4073,N_4279);
and U4565 (N_4565,N_4413,N_3943);
xnor U4566 (N_4566,N_4194,N_4186);
nand U4567 (N_4567,N_4198,N_3980);
xor U4568 (N_4568,N_4408,N_3794);
nor U4569 (N_4569,N_4273,N_4047);
and U4570 (N_4570,N_4119,N_4312);
and U4571 (N_4571,N_3972,N_4336);
and U4572 (N_4572,N_4294,N_4340);
nor U4573 (N_4573,N_3849,N_3996);
nor U4574 (N_4574,N_3830,N_4283);
and U4575 (N_4575,N_3845,N_4214);
or U4576 (N_4576,N_3859,N_4001);
nand U4577 (N_4577,N_4239,N_4038);
xnor U4578 (N_4578,N_4464,N_4189);
nand U4579 (N_4579,N_3807,N_4087);
and U4580 (N_4580,N_4368,N_4254);
nand U4581 (N_4581,N_3766,N_3910);
and U4582 (N_4582,N_4145,N_4216);
nor U4583 (N_4583,N_3771,N_4156);
xor U4584 (N_4584,N_4292,N_4008);
and U4585 (N_4585,N_4417,N_4481);
or U4586 (N_4586,N_4370,N_4338);
xnor U4587 (N_4587,N_4226,N_4062);
and U4588 (N_4588,N_3765,N_4070);
xor U4589 (N_4589,N_4391,N_4066);
and U4590 (N_4590,N_4006,N_4335);
and U4591 (N_4591,N_3950,N_3786);
or U4592 (N_4592,N_4098,N_3757);
or U4593 (N_4593,N_4228,N_3877);
nor U4594 (N_4594,N_3891,N_3800);
nand U4595 (N_4595,N_3791,N_4382);
nor U4596 (N_4596,N_4099,N_3976);
nand U4597 (N_4597,N_4152,N_4449);
nor U4598 (N_4598,N_3867,N_4453);
nand U4599 (N_4599,N_4304,N_4316);
and U4600 (N_4600,N_3779,N_3918);
xor U4601 (N_4601,N_4188,N_4249);
xor U4602 (N_4602,N_3793,N_4088);
nand U4603 (N_4603,N_3915,N_4346);
nor U4604 (N_4604,N_4422,N_4200);
nor U4605 (N_4605,N_4018,N_3853);
and U4606 (N_4606,N_4262,N_4372);
and U4607 (N_4607,N_4288,N_4380);
xnor U4608 (N_4608,N_3906,N_4121);
and U4609 (N_4609,N_4379,N_3816);
xnor U4610 (N_4610,N_3797,N_4067);
xnor U4611 (N_4611,N_4169,N_4494);
or U4612 (N_4612,N_4393,N_4478);
nand U4613 (N_4613,N_4229,N_4474);
nor U4614 (N_4614,N_3824,N_3989);
or U4615 (N_4615,N_4400,N_4222);
xor U4616 (N_4616,N_3967,N_4434);
and U4617 (N_4617,N_3970,N_4117);
or U4618 (N_4618,N_4348,N_3940);
and U4619 (N_4619,N_4302,N_4371);
nand U4620 (N_4620,N_4458,N_3869);
xor U4621 (N_4621,N_4125,N_3776);
nor U4622 (N_4622,N_4028,N_4448);
nor U4623 (N_4623,N_3985,N_4331);
nand U4624 (N_4624,N_3969,N_4389);
and U4625 (N_4625,N_4324,N_4352);
nand U4626 (N_4626,N_4050,N_4369);
nor U4627 (N_4627,N_4052,N_3848);
nand U4628 (N_4628,N_4086,N_4472);
or U4629 (N_4629,N_4060,N_4095);
xor U4630 (N_4630,N_3820,N_3852);
or U4631 (N_4631,N_3884,N_4303);
nand U4632 (N_4632,N_3769,N_4365);
or U4633 (N_4633,N_4040,N_4197);
xnor U4634 (N_4634,N_3977,N_4295);
xnor U4635 (N_4635,N_4355,N_3889);
or U4636 (N_4636,N_4101,N_3978);
nand U4637 (N_4637,N_3831,N_4440);
xor U4638 (N_4638,N_3951,N_3847);
xor U4639 (N_4639,N_4049,N_3973);
or U4640 (N_4640,N_4296,N_4360);
nor U4641 (N_4641,N_3932,N_4490);
and U4642 (N_4642,N_4456,N_3858);
nor U4643 (N_4643,N_4495,N_3984);
nand U4644 (N_4644,N_3875,N_4092);
and U4645 (N_4645,N_3986,N_4475);
and U4646 (N_4646,N_4412,N_3964);
and U4647 (N_4647,N_3813,N_4392);
nor U4648 (N_4648,N_4109,N_3960);
xor U4649 (N_4649,N_4168,N_3775);
nor U4650 (N_4650,N_4469,N_3954);
nand U4651 (N_4651,N_3783,N_3887);
xnor U4652 (N_4652,N_4224,N_4339);
nor U4653 (N_4653,N_4151,N_3934);
nor U4654 (N_4654,N_3817,N_4083);
nor U4655 (N_4655,N_4103,N_4165);
or U4656 (N_4656,N_3835,N_4253);
or U4657 (N_4657,N_3760,N_4031);
or U4658 (N_4658,N_4314,N_3772);
nor U4659 (N_4659,N_4286,N_3990);
nand U4660 (N_4660,N_4220,N_4270);
or U4661 (N_4661,N_3991,N_3944);
and U4662 (N_4662,N_3780,N_4381);
or U4663 (N_4663,N_3767,N_3905);
or U4664 (N_4664,N_3981,N_4497);
or U4665 (N_4665,N_4305,N_4410);
and U4666 (N_4666,N_4307,N_4055);
nand U4667 (N_4667,N_4461,N_4334);
nand U4668 (N_4668,N_3796,N_4470);
nor U4669 (N_4669,N_3925,N_4484);
xor U4670 (N_4670,N_3914,N_4009);
or U4671 (N_4671,N_4120,N_4091);
nand U4672 (N_4672,N_4377,N_4366);
nor U4673 (N_4673,N_4397,N_4261);
or U4674 (N_4674,N_3790,N_4078);
and U4675 (N_4675,N_3966,N_4232);
nor U4676 (N_4676,N_4446,N_4300);
and U4677 (N_4677,N_3881,N_3893);
and U4678 (N_4678,N_4190,N_3819);
or U4679 (N_4679,N_3841,N_4297);
nand U4680 (N_4680,N_3957,N_3764);
and U4681 (N_4681,N_4096,N_4248);
nor U4682 (N_4682,N_3908,N_4264);
or U4683 (N_4683,N_4327,N_4234);
or U4684 (N_4684,N_4419,N_4411);
and U4685 (N_4685,N_4157,N_4245);
nand U4686 (N_4686,N_3892,N_4477);
or U4687 (N_4687,N_4035,N_4473);
xnor U4688 (N_4688,N_4129,N_3836);
xnor U4689 (N_4689,N_3777,N_4444);
nand U4690 (N_4690,N_3994,N_3999);
and U4691 (N_4691,N_4424,N_3762);
or U4692 (N_4692,N_3788,N_4175);
or U4693 (N_4693,N_4404,N_4159);
or U4694 (N_4694,N_4277,N_4238);
or U4695 (N_4695,N_4425,N_4211);
nor U4696 (N_4696,N_4231,N_3752);
nor U4697 (N_4697,N_3770,N_4429);
nand U4698 (N_4698,N_3851,N_3809);
xor U4699 (N_4699,N_3896,N_4236);
nor U4700 (N_4700,N_4030,N_4395);
nand U4701 (N_4701,N_4208,N_4081);
nand U4702 (N_4702,N_4045,N_4138);
nor U4703 (N_4703,N_3888,N_4021);
xor U4704 (N_4704,N_4069,N_4170);
and U4705 (N_4705,N_3983,N_4266);
nand U4706 (N_4706,N_4112,N_4178);
xnor U4707 (N_4707,N_4420,N_4250);
nand U4708 (N_4708,N_4493,N_4085);
nor U4709 (N_4709,N_4322,N_4124);
or U4710 (N_4710,N_4255,N_3808);
nand U4711 (N_4711,N_3826,N_4054);
xnor U4712 (N_4712,N_4026,N_4491);
nor U4713 (N_4713,N_3902,N_3846);
and U4714 (N_4714,N_4451,N_4003);
nand U4715 (N_4715,N_4311,N_4041);
or U4716 (N_4716,N_4358,N_3958);
nand U4717 (N_4717,N_3818,N_4384);
and U4718 (N_4718,N_3992,N_4315);
and U4719 (N_4719,N_3855,N_4337);
nand U4720 (N_4720,N_4046,N_3856);
and U4721 (N_4721,N_4019,N_4206);
or U4722 (N_4722,N_4462,N_4241);
nand U4723 (N_4723,N_4356,N_4321);
xnor U4724 (N_4724,N_4276,N_4486);
nor U4725 (N_4725,N_4401,N_4405);
and U4726 (N_4726,N_4097,N_3963);
or U4727 (N_4727,N_4247,N_4265);
nor U4728 (N_4728,N_4278,N_3854);
or U4729 (N_4729,N_3959,N_4218);
or U4730 (N_4730,N_3751,N_4439);
and U4731 (N_4731,N_4394,N_4079);
and U4732 (N_4732,N_3850,N_4457);
nand U4733 (N_4733,N_4235,N_4496);
and U4734 (N_4734,N_4426,N_3965);
nor U4735 (N_4735,N_3920,N_4326);
nand U4736 (N_4736,N_3942,N_4122);
or U4737 (N_4737,N_3865,N_4454);
xor U4738 (N_4738,N_4011,N_3988);
nor U4739 (N_4739,N_4094,N_3945);
nor U4740 (N_4740,N_4361,N_4343);
or U4741 (N_4741,N_4020,N_4107);
nor U4742 (N_4742,N_4258,N_3864);
nor U4743 (N_4743,N_4090,N_3866);
or U4744 (N_4744,N_3756,N_4134);
nor U4745 (N_4745,N_3987,N_4205);
and U4746 (N_4746,N_4146,N_4155);
and U4747 (N_4747,N_4147,N_4164);
and U4748 (N_4748,N_4080,N_3929);
nand U4749 (N_4749,N_3948,N_4299);
nand U4750 (N_4750,N_3773,N_4460);
xor U4751 (N_4751,N_3955,N_3998);
and U4752 (N_4752,N_4268,N_4269);
xor U4753 (N_4753,N_4183,N_3953);
xor U4754 (N_4754,N_4259,N_4174);
and U4755 (N_4755,N_3995,N_3840);
nand U4756 (N_4756,N_4015,N_3931);
or U4757 (N_4757,N_4115,N_4310);
nor U4758 (N_4758,N_3947,N_4013);
nor U4759 (N_4759,N_4204,N_3895);
nand U4760 (N_4760,N_4000,N_3838);
or U4761 (N_4761,N_3815,N_4428);
nand U4762 (N_4762,N_4272,N_4378);
nand U4763 (N_4763,N_4427,N_4333);
or U4764 (N_4764,N_4036,N_4436);
xor U4765 (N_4765,N_4287,N_4251);
nand U4766 (N_4766,N_4184,N_3868);
nand U4767 (N_4767,N_4313,N_3933);
and U4768 (N_4768,N_4133,N_4328);
nor U4769 (N_4769,N_3857,N_4482);
or U4770 (N_4770,N_4140,N_3778);
and U4771 (N_4771,N_4443,N_4463);
xor U4772 (N_4772,N_3912,N_4480);
nand U4773 (N_4773,N_4483,N_4135);
nand U4774 (N_4774,N_4257,N_3946);
or U4775 (N_4775,N_4139,N_3759);
nor U4776 (N_4776,N_4306,N_4072);
nand U4777 (N_4777,N_4350,N_4240);
and U4778 (N_4778,N_4150,N_4010);
and U4779 (N_4779,N_4421,N_4318);
or U4780 (N_4780,N_4237,N_3753);
nor U4781 (N_4781,N_4341,N_3814);
xnor U4782 (N_4782,N_4438,N_4459);
xor U4783 (N_4783,N_3871,N_3941);
and U4784 (N_4784,N_4128,N_3974);
and U4785 (N_4785,N_4162,N_3844);
or U4786 (N_4786,N_4032,N_4467);
nor U4787 (N_4787,N_4388,N_4075);
nor U4788 (N_4788,N_3781,N_4376);
and U4789 (N_4789,N_4329,N_3787);
and U4790 (N_4790,N_3962,N_4344);
nand U4791 (N_4791,N_4039,N_4445);
nor U4792 (N_4792,N_4363,N_4153);
nand U4793 (N_4793,N_4332,N_4185);
nor U4794 (N_4794,N_4017,N_4403);
nor U4795 (N_4795,N_4126,N_4430);
and U4796 (N_4796,N_3898,N_4022);
xnor U4797 (N_4797,N_4025,N_4383);
and U4798 (N_4798,N_4243,N_3761);
xnor U4799 (N_4799,N_4398,N_3833);
and U4800 (N_4800,N_3812,N_4203);
or U4801 (N_4801,N_4108,N_4063);
nand U4802 (N_4802,N_4242,N_4349);
xnor U4803 (N_4803,N_3917,N_4351);
nor U4804 (N_4804,N_4176,N_3921);
or U4805 (N_4805,N_3768,N_4143);
nand U4806 (N_4806,N_3804,N_4284);
nor U4807 (N_4807,N_4100,N_3784);
nor U4808 (N_4808,N_3961,N_4387);
xor U4809 (N_4809,N_3880,N_4201);
nor U4810 (N_4810,N_3805,N_4173);
or U4811 (N_4811,N_3936,N_3975);
or U4812 (N_4812,N_4271,N_4202);
xor U4813 (N_4813,N_3792,N_4195);
xnor U4814 (N_4814,N_4217,N_4212);
or U4815 (N_4815,N_4347,N_4044);
xnor U4816 (N_4816,N_4330,N_4342);
nand U4817 (N_4817,N_4285,N_3993);
nor U4818 (N_4818,N_4452,N_3897);
nand U4819 (N_4819,N_4148,N_4260);
or U4820 (N_4820,N_4256,N_4123);
or U4821 (N_4821,N_4004,N_3911);
xnor U4822 (N_4822,N_4149,N_4275);
or U4823 (N_4823,N_4142,N_3919);
nand U4824 (N_4824,N_4373,N_4385);
nand U4825 (N_4825,N_4084,N_4053);
and U4826 (N_4826,N_4359,N_3872);
nor U4827 (N_4827,N_4210,N_4320);
or U4828 (N_4828,N_4076,N_4301);
and U4829 (N_4829,N_4136,N_3795);
nor U4830 (N_4830,N_3982,N_3909);
or U4831 (N_4831,N_4450,N_3903);
nand U4832 (N_4832,N_4252,N_4441);
nand U4833 (N_4833,N_3825,N_4102);
nand U4834 (N_4834,N_3956,N_4437);
or U4835 (N_4835,N_4227,N_4048);
nand U4836 (N_4836,N_4167,N_3873);
nor U4837 (N_4837,N_4414,N_4130);
nor U4838 (N_4838,N_4093,N_3834);
nand U4839 (N_4839,N_3997,N_4488);
nor U4840 (N_4840,N_4104,N_4179);
or U4841 (N_4841,N_4274,N_4233);
or U4842 (N_4842,N_3798,N_3904);
nor U4843 (N_4843,N_3827,N_3843);
nand U4844 (N_4844,N_4498,N_3928);
and U4845 (N_4845,N_4059,N_3750);
xnor U4846 (N_4846,N_4196,N_3782);
xnor U4847 (N_4847,N_4002,N_4137);
or U4848 (N_4848,N_3923,N_4407);
xor U4849 (N_4849,N_4423,N_4431);
or U4850 (N_4850,N_4353,N_4308);
nor U4851 (N_4851,N_4375,N_3863);
nand U4852 (N_4852,N_4479,N_4476);
nor U4853 (N_4853,N_4280,N_4007);
nand U4854 (N_4854,N_4409,N_4177);
nor U4855 (N_4855,N_4221,N_4144);
and U4856 (N_4856,N_4187,N_4290);
nor U4857 (N_4857,N_3832,N_4074);
nand U4858 (N_4858,N_3862,N_4014);
nor U4859 (N_4859,N_4110,N_4263);
xnor U4860 (N_4860,N_4027,N_4116);
xnor U4861 (N_4861,N_4154,N_3968);
nor U4862 (N_4862,N_3878,N_4415);
xnor U4863 (N_4863,N_3952,N_4105);
nand U4864 (N_4864,N_4029,N_4396);
xor U4865 (N_4865,N_4037,N_4289);
nand U4866 (N_4866,N_4163,N_4111);
or U4867 (N_4867,N_4118,N_4362);
nor U4868 (N_4868,N_3913,N_4182);
and U4869 (N_4869,N_4089,N_4127);
and U4870 (N_4870,N_4191,N_4058);
or U4871 (N_4871,N_4298,N_3886);
nor U4872 (N_4872,N_4043,N_4416);
or U4873 (N_4873,N_4193,N_4323);
or U4874 (N_4874,N_4033,N_4485);
nand U4875 (N_4875,N_3883,N_4343);
nand U4876 (N_4876,N_3976,N_4377);
nand U4877 (N_4877,N_4336,N_3929);
nor U4878 (N_4878,N_3955,N_4051);
nor U4879 (N_4879,N_4489,N_3762);
nor U4880 (N_4880,N_3855,N_4134);
nor U4881 (N_4881,N_3832,N_4137);
nor U4882 (N_4882,N_4469,N_4496);
xnor U4883 (N_4883,N_3884,N_4208);
nand U4884 (N_4884,N_3970,N_4275);
and U4885 (N_4885,N_4338,N_4007);
or U4886 (N_4886,N_4020,N_4151);
xnor U4887 (N_4887,N_4113,N_4370);
nand U4888 (N_4888,N_3925,N_4062);
or U4889 (N_4889,N_4280,N_4248);
or U4890 (N_4890,N_4037,N_4315);
nor U4891 (N_4891,N_4052,N_3955);
or U4892 (N_4892,N_4463,N_4003);
nor U4893 (N_4893,N_3855,N_4129);
nor U4894 (N_4894,N_4356,N_4250);
or U4895 (N_4895,N_4407,N_4341);
or U4896 (N_4896,N_3882,N_4263);
and U4897 (N_4897,N_4291,N_4040);
nand U4898 (N_4898,N_4099,N_4218);
or U4899 (N_4899,N_4366,N_4468);
xnor U4900 (N_4900,N_3917,N_3889);
xor U4901 (N_4901,N_4280,N_3923);
and U4902 (N_4902,N_4156,N_4331);
nor U4903 (N_4903,N_4375,N_4362);
and U4904 (N_4904,N_4423,N_3955);
nand U4905 (N_4905,N_4115,N_4185);
nand U4906 (N_4906,N_4446,N_4057);
xnor U4907 (N_4907,N_4054,N_4143);
and U4908 (N_4908,N_3954,N_3850);
and U4909 (N_4909,N_4426,N_3792);
and U4910 (N_4910,N_4146,N_3776);
nor U4911 (N_4911,N_3963,N_3909);
or U4912 (N_4912,N_3816,N_4375);
and U4913 (N_4913,N_3962,N_4241);
nor U4914 (N_4914,N_4227,N_3753);
or U4915 (N_4915,N_4273,N_3951);
nor U4916 (N_4916,N_4074,N_4047);
or U4917 (N_4917,N_4223,N_4346);
nand U4918 (N_4918,N_4237,N_3879);
or U4919 (N_4919,N_4180,N_3952);
xor U4920 (N_4920,N_4392,N_3881);
and U4921 (N_4921,N_3865,N_3870);
nand U4922 (N_4922,N_4306,N_4376);
and U4923 (N_4923,N_4495,N_4181);
nand U4924 (N_4924,N_3830,N_4408);
xnor U4925 (N_4925,N_3899,N_4273);
and U4926 (N_4926,N_4467,N_4493);
and U4927 (N_4927,N_4131,N_3857);
nand U4928 (N_4928,N_4458,N_4258);
and U4929 (N_4929,N_3886,N_3982);
xnor U4930 (N_4930,N_4430,N_4295);
nand U4931 (N_4931,N_3775,N_4437);
or U4932 (N_4932,N_3831,N_4482);
nor U4933 (N_4933,N_3969,N_3974);
and U4934 (N_4934,N_4345,N_3912);
xnor U4935 (N_4935,N_4405,N_4385);
xnor U4936 (N_4936,N_4386,N_4279);
xor U4937 (N_4937,N_3887,N_3789);
nor U4938 (N_4938,N_3837,N_4426);
nand U4939 (N_4939,N_4475,N_4111);
or U4940 (N_4940,N_4140,N_3871);
xor U4941 (N_4941,N_3919,N_4023);
nor U4942 (N_4942,N_3943,N_4074);
nor U4943 (N_4943,N_4257,N_4391);
or U4944 (N_4944,N_3787,N_3935);
and U4945 (N_4945,N_4085,N_3935);
xor U4946 (N_4946,N_3792,N_4029);
or U4947 (N_4947,N_4390,N_4491);
xnor U4948 (N_4948,N_4215,N_4091);
and U4949 (N_4949,N_3836,N_4350);
or U4950 (N_4950,N_4333,N_3927);
xor U4951 (N_4951,N_3991,N_4151);
xnor U4952 (N_4952,N_4049,N_3955);
nand U4953 (N_4953,N_4360,N_3998);
nand U4954 (N_4954,N_3979,N_3811);
or U4955 (N_4955,N_4457,N_4374);
and U4956 (N_4956,N_4473,N_3953);
xor U4957 (N_4957,N_4334,N_3884);
nand U4958 (N_4958,N_3953,N_4069);
and U4959 (N_4959,N_4002,N_4254);
and U4960 (N_4960,N_4401,N_4195);
and U4961 (N_4961,N_3763,N_4410);
or U4962 (N_4962,N_4051,N_4057);
xor U4963 (N_4963,N_4464,N_4364);
xnor U4964 (N_4964,N_3780,N_3958);
xnor U4965 (N_4965,N_4304,N_3806);
xor U4966 (N_4966,N_4162,N_4350);
or U4967 (N_4967,N_4113,N_3919);
xnor U4968 (N_4968,N_3797,N_4099);
xor U4969 (N_4969,N_4120,N_4306);
nor U4970 (N_4970,N_4276,N_4465);
nand U4971 (N_4971,N_4436,N_3758);
and U4972 (N_4972,N_4192,N_3880);
xor U4973 (N_4973,N_4092,N_4315);
and U4974 (N_4974,N_4479,N_4003);
nand U4975 (N_4975,N_4057,N_4113);
xnor U4976 (N_4976,N_4228,N_4085);
or U4977 (N_4977,N_4210,N_4039);
nand U4978 (N_4978,N_4407,N_3938);
nand U4979 (N_4979,N_4494,N_3847);
xnor U4980 (N_4980,N_4306,N_3858);
nand U4981 (N_4981,N_4036,N_4016);
or U4982 (N_4982,N_4329,N_4174);
and U4983 (N_4983,N_4292,N_3821);
or U4984 (N_4984,N_3787,N_4276);
nor U4985 (N_4985,N_3919,N_4337);
nor U4986 (N_4986,N_3959,N_3869);
xor U4987 (N_4987,N_4468,N_4439);
and U4988 (N_4988,N_4291,N_4472);
or U4989 (N_4989,N_4108,N_4000);
nand U4990 (N_4990,N_4300,N_3919);
nand U4991 (N_4991,N_4383,N_4090);
nand U4992 (N_4992,N_4119,N_3881);
nor U4993 (N_4993,N_4183,N_4146);
nor U4994 (N_4994,N_4410,N_4279);
and U4995 (N_4995,N_4447,N_4040);
or U4996 (N_4996,N_4442,N_4239);
nand U4997 (N_4997,N_4056,N_4171);
or U4998 (N_4998,N_4045,N_3852);
and U4999 (N_4999,N_4314,N_4221);
xnor U5000 (N_5000,N_4384,N_4275);
xnor U5001 (N_5001,N_4428,N_4060);
nand U5002 (N_5002,N_3853,N_3837);
or U5003 (N_5003,N_3978,N_3775);
nand U5004 (N_5004,N_3767,N_4089);
and U5005 (N_5005,N_4369,N_4493);
nor U5006 (N_5006,N_3953,N_4207);
nor U5007 (N_5007,N_4221,N_4151);
nand U5008 (N_5008,N_3764,N_4270);
and U5009 (N_5009,N_4100,N_4229);
or U5010 (N_5010,N_4050,N_4412);
xnor U5011 (N_5011,N_3972,N_4116);
xnor U5012 (N_5012,N_4473,N_4318);
nor U5013 (N_5013,N_4425,N_3891);
or U5014 (N_5014,N_3782,N_4069);
nand U5015 (N_5015,N_3819,N_3858);
nor U5016 (N_5016,N_4133,N_3903);
nand U5017 (N_5017,N_4402,N_4422);
nor U5018 (N_5018,N_3767,N_4428);
or U5019 (N_5019,N_4380,N_3806);
nor U5020 (N_5020,N_4198,N_4493);
nand U5021 (N_5021,N_3831,N_4062);
or U5022 (N_5022,N_4253,N_4051);
xnor U5023 (N_5023,N_3902,N_3795);
xnor U5024 (N_5024,N_3969,N_4357);
nor U5025 (N_5025,N_4379,N_4224);
xnor U5026 (N_5026,N_4403,N_4261);
nor U5027 (N_5027,N_4402,N_4067);
nor U5028 (N_5028,N_4493,N_4163);
or U5029 (N_5029,N_4170,N_4380);
and U5030 (N_5030,N_4110,N_4154);
nor U5031 (N_5031,N_4370,N_3770);
or U5032 (N_5032,N_4430,N_4194);
nor U5033 (N_5033,N_4038,N_4387);
and U5034 (N_5034,N_3896,N_3860);
xnor U5035 (N_5035,N_4096,N_3864);
or U5036 (N_5036,N_4212,N_3822);
or U5037 (N_5037,N_3788,N_4033);
nand U5038 (N_5038,N_4005,N_4187);
nand U5039 (N_5039,N_4467,N_4211);
nor U5040 (N_5040,N_4403,N_4484);
nand U5041 (N_5041,N_3790,N_3951);
nor U5042 (N_5042,N_4394,N_4339);
or U5043 (N_5043,N_4071,N_3919);
nand U5044 (N_5044,N_3939,N_4232);
nor U5045 (N_5045,N_4041,N_3986);
or U5046 (N_5046,N_4302,N_4240);
or U5047 (N_5047,N_4361,N_4221);
xor U5048 (N_5048,N_4009,N_4293);
or U5049 (N_5049,N_4334,N_4477);
nor U5050 (N_5050,N_4035,N_4381);
nor U5051 (N_5051,N_4166,N_4108);
or U5052 (N_5052,N_3821,N_3976);
and U5053 (N_5053,N_4317,N_3912);
and U5054 (N_5054,N_4471,N_4067);
and U5055 (N_5055,N_4459,N_4063);
or U5056 (N_5056,N_3828,N_3764);
nor U5057 (N_5057,N_4476,N_4077);
and U5058 (N_5058,N_3933,N_4454);
nand U5059 (N_5059,N_4273,N_4348);
xnor U5060 (N_5060,N_4273,N_3903);
and U5061 (N_5061,N_3818,N_4493);
nor U5062 (N_5062,N_3898,N_4362);
nor U5063 (N_5063,N_4480,N_3987);
or U5064 (N_5064,N_3995,N_4292);
or U5065 (N_5065,N_4066,N_3869);
nand U5066 (N_5066,N_3984,N_3845);
and U5067 (N_5067,N_4335,N_3862);
xor U5068 (N_5068,N_4358,N_4368);
nor U5069 (N_5069,N_4025,N_4361);
or U5070 (N_5070,N_4135,N_4299);
nor U5071 (N_5071,N_4056,N_3971);
nor U5072 (N_5072,N_3798,N_4022);
and U5073 (N_5073,N_4366,N_3961);
xnor U5074 (N_5074,N_4253,N_3883);
xnor U5075 (N_5075,N_3868,N_4425);
and U5076 (N_5076,N_3908,N_3785);
or U5077 (N_5077,N_4106,N_4174);
nor U5078 (N_5078,N_4275,N_4017);
nor U5079 (N_5079,N_4247,N_4483);
nor U5080 (N_5080,N_4233,N_3984);
nor U5081 (N_5081,N_4472,N_4314);
or U5082 (N_5082,N_4006,N_4014);
or U5083 (N_5083,N_4233,N_4208);
or U5084 (N_5084,N_4457,N_3782);
nor U5085 (N_5085,N_3889,N_4001);
and U5086 (N_5086,N_3753,N_4335);
nor U5087 (N_5087,N_3824,N_4001);
nand U5088 (N_5088,N_4187,N_4221);
nor U5089 (N_5089,N_4204,N_3809);
or U5090 (N_5090,N_3885,N_3832);
nor U5091 (N_5091,N_3763,N_4186);
and U5092 (N_5092,N_4372,N_3847);
or U5093 (N_5093,N_4322,N_4381);
nor U5094 (N_5094,N_4202,N_4483);
and U5095 (N_5095,N_4076,N_4125);
nand U5096 (N_5096,N_4414,N_4220);
and U5097 (N_5097,N_4250,N_4296);
xnor U5098 (N_5098,N_3914,N_4291);
or U5099 (N_5099,N_4005,N_4234);
nand U5100 (N_5100,N_3966,N_4415);
and U5101 (N_5101,N_3973,N_4312);
nand U5102 (N_5102,N_3809,N_4015);
nor U5103 (N_5103,N_4377,N_3932);
xnor U5104 (N_5104,N_4048,N_4121);
or U5105 (N_5105,N_3917,N_4447);
nand U5106 (N_5106,N_4146,N_3751);
or U5107 (N_5107,N_3972,N_4497);
nor U5108 (N_5108,N_4061,N_4155);
and U5109 (N_5109,N_4454,N_4033);
and U5110 (N_5110,N_4388,N_3938);
nor U5111 (N_5111,N_3797,N_4238);
nand U5112 (N_5112,N_4017,N_4208);
or U5113 (N_5113,N_4057,N_3922);
xnor U5114 (N_5114,N_4133,N_4275);
or U5115 (N_5115,N_4418,N_4062);
nor U5116 (N_5116,N_3982,N_4451);
and U5117 (N_5117,N_4272,N_4140);
nand U5118 (N_5118,N_3792,N_3778);
xnor U5119 (N_5119,N_4141,N_4453);
or U5120 (N_5120,N_3810,N_4447);
nand U5121 (N_5121,N_4246,N_4443);
nor U5122 (N_5122,N_3750,N_4273);
nand U5123 (N_5123,N_4421,N_4466);
xor U5124 (N_5124,N_4070,N_4357);
or U5125 (N_5125,N_3959,N_4350);
nor U5126 (N_5126,N_3771,N_4313);
and U5127 (N_5127,N_3803,N_4489);
xnor U5128 (N_5128,N_3827,N_3965);
xnor U5129 (N_5129,N_3985,N_4249);
or U5130 (N_5130,N_4033,N_4183);
nor U5131 (N_5131,N_3853,N_4201);
nand U5132 (N_5132,N_4309,N_3960);
xor U5133 (N_5133,N_4344,N_3766);
xnor U5134 (N_5134,N_4349,N_4292);
nor U5135 (N_5135,N_4458,N_3946);
xnor U5136 (N_5136,N_4499,N_4362);
and U5137 (N_5137,N_4494,N_3895);
and U5138 (N_5138,N_4137,N_4227);
nand U5139 (N_5139,N_4338,N_3786);
nand U5140 (N_5140,N_4237,N_4413);
nor U5141 (N_5141,N_3783,N_4340);
xnor U5142 (N_5142,N_4128,N_3906);
xor U5143 (N_5143,N_4037,N_3807);
nand U5144 (N_5144,N_3953,N_3966);
nor U5145 (N_5145,N_3993,N_4117);
and U5146 (N_5146,N_4301,N_4249);
xor U5147 (N_5147,N_3963,N_4471);
or U5148 (N_5148,N_4139,N_4166);
or U5149 (N_5149,N_4405,N_4437);
nand U5150 (N_5150,N_3924,N_4452);
or U5151 (N_5151,N_4418,N_4381);
or U5152 (N_5152,N_4185,N_4053);
or U5153 (N_5153,N_4356,N_3861);
nand U5154 (N_5154,N_4045,N_4198);
xnor U5155 (N_5155,N_3837,N_4279);
xnor U5156 (N_5156,N_4271,N_4342);
and U5157 (N_5157,N_4348,N_3997);
and U5158 (N_5158,N_4262,N_4487);
or U5159 (N_5159,N_4480,N_3990);
nor U5160 (N_5160,N_4336,N_3997);
and U5161 (N_5161,N_3905,N_4073);
xor U5162 (N_5162,N_4049,N_4453);
nor U5163 (N_5163,N_4099,N_3915);
xor U5164 (N_5164,N_4059,N_3985);
xor U5165 (N_5165,N_4236,N_4243);
nand U5166 (N_5166,N_3873,N_3855);
and U5167 (N_5167,N_4217,N_4453);
nor U5168 (N_5168,N_4093,N_4241);
nor U5169 (N_5169,N_4009,N_4010);
and U5170 (N_5170,N_4139,N_4222);
xor U5171 (N_5171,N_4435,N_3869);
xnor U5172 (N_5172,N_4301,N_3820);
nor U5173 (N_5173,N_4236,N_4180);
nor U5174 (N_5174,N_4311,N_3914);
xnor U5175 (N_5175,N_4144,N_3901);
nand U5176 (N_5176,N_3894,N_4279);
xnor U5177 (N_5177,N_4222,N_4118);
nor U5178 (N_5178,N_3799,N_3927);
nor U5179 (N_5179,N_4134,N_4019);
and U5180 (N_5180,N_4114,N_4374);
xnor U5181 (N_5181,N_4462,N_3947);
xnor U5182 (N_5182,N_3963,N_3784);
and U5183 (N_5183,N_4282,N_4478);
and U5184 (N_5184,N_4409,N_3927);
or U5185 (N_5185,N_3871,N_3957);
and U5186 (N_5186,N_3751,N_4388);
and U5187 (N_5187,N_4199,N_4197);
xnor U5188 (N_5188,N_3992,N_4012);
nor U5189 (N_5189,N_4060,N_4133);
xnor U5190 (N_5190,N_4379,N_4071);
nor U5191 (N_5191,N_3862,N_4411);
xor U5192 (N_5192,N_4117,N_3967);
and U5193 (N_5193,N_4019,N_4030);
nor U5194 (N_5194,N_3969,N_3848);
nor U5195 (N_5195,N_4123,N_4186);
xnor U5196 (N_5196,N_4193,N_3752);
nor U5197 (N_5197,N_3838,N_3884);
or U5198 (N_5198,N_4314,N_3839);
or U5199 (N_5199,N_4375,N_4109);
and U5200 (N_5200,N_3976,N_3854);
or U5201 (N_5201,N_4494,N_3946);
nor U5202 (N_5202,N_3773,N_4356);
nor U5203 (N_5203,N_4398,N_4469);
and U5204 (N_5204,N_4286,N_4041);
and U5205 (N_5205,N_4139,N_4383);
or U5206 (N_5206,N_3932,N_4097);
or U5207 (N_5207,N_4038,N_3935);
nand U5208 (N_5208,N_3942,N_4421);
and U5209 (N_5209,N_4341,N_4361);
xnor U5210 (N_5210,N_3789,N_4215);
xnor U5211 (N_5211,N_4306,N_3788);
nor U5212 (N_5212,N_3811,N_3945);
xnor U5213 (N_5213,N_4093,N_3844);
xor U5214 (N_5214,N_4390,N_4268);
nor U5215 (N_5215,N_4357,N_3974);
nor U5216 (N_5216,N_3827,N_3879);
nand U5217 (N_5217,N_4325,N_3808);
or U5218 (N_5218,N_3831,N_3974);
xor U5219 (N_5219,N_4047,N_4380);
nand U5220 (N_5220,N_3996,N_4306);
xnor U5221 (N_5221,N_4459,N_4481);
or U5222 (N_5222,N_3970,N_4004);
or U5223 (N_5223,N_3873,N_4225);
xnor U5224 (N_5224,N_4341,N_4405);
nor U5225 (N_5225,N_4461,N_3902);
xnor U5226 (N_5226,N_4249,N_3780);
and U5227 (N_5227,N_4072,N_4444);
or U5228 (N_5228,N_4018,N_4426);
or U5229 (N_5229,N_4008,N_4113);
nand U5230 (N_5230,N_3901,N_4089);
and U5231 (N_5231,N_3754,N_4369);
nand U5232 (N_5232,N_4430,N_4289);
xor U5233 (N_5233,N_3963,N_4152);
xor U5234 (N_5234,N_4420,N_3852);
and U5235 (N_5235,N_4374,N_4442);
nor U5236 (N_5236,N_4029,N_4126);
and U5237 (N_5237,N_3977,N_4497);
nand U5238 (N_5238,N_4145,N_4398);
nor U5239 (N_5239,N_3935,N_3860);
nor U5240 (N_5240,N_4153,N_4455);
xor U5241 (N_5241,N_4343,N_3939);
nor U5242 (N_5242,N_4195,N_4355);
or U5243 (N_5243,N_4143,N_4397);
nor U5244 (N_5244,N_3969,N_4047);
and U5245 (N_5245,N_3843,N_3764);
or U5246 (N_5246,N_4429,N_3825);
nand U5247 (N_5247,N_3944,N_3864);
nand U5248 (N_5248,N_3787,N_4045);
or U5249 (N_5249,N_3759,N_4410);
nand U5250 (N_5250,N_4808,N_4967);
xor U5251 (N_5251,N_4766,N_4831);
or U5252 (N_5252,N_4698,N_4796);
and U5253 (N_5253,N_5152,N_4537);
nand U5254 (N_5254,N_4954,N_5038);
and U5255 (N_5255,N_5098,N_5079);
nor U5256 (N_5256,N_5247,N_4754);
and U5257 (N_5257,N_4930,N_5165);
and U5258 (N_5258,N_4784,N_4869);
nand U5259 (N_5259,N_4673,N_4641);
nor U5260 (N_5260,N_4840,N_5199);
or U5261 (N_5261,N_4929,N_4826);
xnor U5262 (N_5262,N_5227,N_4927);
nand U5263 (N_5263,N_4968,N_5032);
nor U5264 (N_5264,N_4616,N_5125);
nor U5265 (N_5265,N_5031,N_4684);
nor U5266 (N_5266,N_5148,N_4696);
and U5267 (N_5267,N_5043,N_4891);
or U5268 (N_5268,N_4623,N_4664);
nor U5269 (N_5269,N_4941,N_4769);
xnor U5270 (N_5270,N_4986,N_4981);
nor U5271 (N_5271,N_4897,N_4645);
nand U5272 (N_5272,N_5062,N_5016);
nor U5273 (N_5273,N_4668,N_5244);
nand U5274 (N_5274,N_5163,N_5178);
and U5275 (N_5275,N_5249,N_4520);
or U5276 (N_5276,N_4579,N_4775);
nand U5277 (N_5277,N_4876,N_4566);
nand U5278 (N_5278,N_4875,N_4828);
nand U5279 (N_5279,N_5193,N_4987);
xnor U5280 (N_5280,N_4720,N_4874);
nor U5281 (N_5281,N_4745,N_4918);
nor U5282 (N_5282,N_4921,N_4822);
xnor U5283 (N_5283,N_4913,N_4719);
and U5284 (N_5284,N_5036,N_5101);
and U5285 (N_5285,N_4732,N_5023);
nor U5286 (N_5286,N_4586,N_4746);
xnor U5287 (N_5287,N_4750,N_5024);
and U5288 (N_5288,N_4847,N_5009);
nor U5289 (N_5289,N_4608,N_4820);
xor U5290 (N_5290,N_4815,N_5129);
nand U5291 (N_5291,N_5056,N_4649);
nor U5292 (N_5292,N_5145,N_4757);
and U5293 (N_5293,N_4912,N_5202);
xor U5294 (N_5294,N_5105,N_5215);
or U5295 (N_5295,N_4853,N_4888);
nor U5296 (N_5296,N_4924,N_5162);
xor U5297 (N_5297,N_4504,N_5059);
and U5298 (N_5298,N_4596,N_4838);
xor U5299 (N_5299,N_5216,N_5067);
and U5300 (N_5300,N_4980,N_4588);
and U5301 (N_5301,N_5205,N_5138);
or U5302 (N_5302,N_5046,N_5226);
nand U5303 (N_5303,N_5231,N_5096);
nand U5304 (N_5304,N_4584,N_4506);
nor U5305 (N_5305,N_5188,N_4546);
nand U5306 (N_5306,N_5189,N_4819);
and U5307 (N_5307,N_5166,N_5242);
xor U5308 (N_5308,N_4837,N_4679);
nor U5309 (N_5309,N_4574,N_5186);
and U5310 (N_5310,N_5159,N_5222);
xnor U5311 (N_5311,N_4501,N_5109);
and U5312 (N_5312,N_5080,N_4605);
xnor U5313 (N_5313,N_5173,N_4843);
or U5314 (N_5314,N_4812,N_4878);
and U5315 (N_5315,N_5124,N_5131);
or U5316 (N_5316,N_4667,N_4798);
nor U5317 (N_5317,N_4965,N_4681);
xnor U5318 (N_5318,N_4758,N_4799);
and U5319 (N_5319,N_4909,N_4829);
nor U5320 (N_5320,N_5097,N_4702);
nor U5321 (N_5321,N_4549,N_4627);
and U5322 (N_5322,N_5091,N_5030);
or U5323 (N_5323,N_4740,N_5183);
nor U5324 (N_5324,N_4656,N_5094);
xnor U5325 (N_5325,N_4850,N_4530);
and U5326 (N_5326,N_4614,N_4657);
nor U5327 (N_5327,N_5132,N_5116);
nor U5328 (N_5328,N_4594,N_4517);
xnor U5329 (N_5329,N_4979,N_5118);
nand U5330 (N_5330,N_4682,N_5089);
nor U5331 (N_5331,N_4917,N_4813);
and U5332 (N_5332,N_4742,N_5156);
or U5333 (N_5333,N_5157,N_4950);
xnor U5334 (N_5334,N_4782,N_4779);
nor U5335 (N_5335,N_4573,N_4639);
and U5336 (N_5336,N_4949,N_4933);
or U5337 (N_5337,N_4814,N_5100);
and U5338 (N_5338,N_5060,N_5200);
xor U5339 (N_5339,N_4728,N_4747);
nor U5340 (N_5340,N_5164,N_4845);
or U5341 (N_5341,N_5083,N_5246);
nand U5342 (N_5342,N_5190,N_5248);
or U5343 (N_5343,N_4772,N_4806);
xor U5344 (N_5344,N_5010,N_4893);
or U5345 (N_5345,N_4926,N_4695);
nand U5346 (N_5346,N_4633,N_5191);
nand U5347 (N_5347,N_5208,N_5114);
nor U5348 (N_5348,N_4866,N_5077);
xor U5349 (N_5349,N_4856,N_4522);
and U5350 (N_5350,N_4699,N_4810);
and U5351 (N_5351,N_4995,N_4857);
and U5352 (N_5352,N_5180,N_5237);
nor U5353 (N_5353,N_5245,N_4593);
nand U5354 (N_5354,N_4726,N_4722);
or U5355 (N_5355,N_4783,N_5185);
nor U5356 (N_5356,N_4983,N_4741);
nand U5357 (N_5357,N_4932,N_4789);
or U5358 (N_5358,N_5001,N_5184);
xor U5359 (N_5359,N_5084,N_4692);
nor U5360 (N_5360,N_4873,N_4727);
nor U5361 (N_5361,N_5135,N_4816);
xnor U5362 (N_5362,N_5017,N_4602);
nand U5363 (N_5363,N_5011,N_5206);
nand U5364 (N_5364,N_5015,N_5230);
xor U5365 (N_5365,N_4640,N_4872);
or U5366 (N_5366,N_4577,N_4825);
or U5367 (N_5367,N_4793,N_4744);
nand U5368 (N_5368,N_4703,N_5221);
nand U5369 (N_5369,N_5238,N_4663);
xor U5370 (N_5370,N_4529,N_4867);
and U5371 (N_5371,N_4567,N_4560);
nor U5372 (N_5372,N_5141,N_5219);
nand U5373 (N_5373,N_4958,N_5140);
nand U5374 (N_5374,N_4998,N_4846);
xor U5375 (N_5375,N_4800,N_5137);
and U5376 (N_5376,N_4778,N_5029);
and U5377 (N_5377,N_5013,N_4707);
and U5378 (N_5378,N_4675,N_4767);
nand U5379 (N_5379,N_5068,N_5171);
or U5380 (N_5380,N_4768,N_4851);
or U5381 (N_5381,N_4548,N_4961);
nand U5382 (N_5382,N_5217,N_5053);
xor U5383 (N_5383,N_5092,N_4672);
or U5384 (N_5384,N_4642,N_5233);
nor U5385 (N_5385,N_4585,N_4882);
nand U5386 (N_5386,N_4774,N_4559);
or U5387 (N_5387,N_5212,N_4561);
and U5388 (N_5388,N_4615,N_4944);
and U5389 (N_5389,N_4660,N_5058);
nand U5390 (N_5390,N_5181,N_4931);
or U5391 (N_5391,N_5050,N_4580);
xor U5392 (N_5392,N_5057,N_4599);
or U5393 (N_5393,N_5147,N_4571);
xor U5394 (N_5394,N_4895,N_4724);
nor U5395 (N_5395,N_4677,N_5134);
nand U5396 (N_5396,N_5161,N_4592);
or U5397 (N_5397,N_4734,N_5085);
nor U5398 (N_5398,N_4512,N_4666);
or U5399 (N_5399,N_4794,N_4948);
xor U5400 (N_5400,N_5123,N_4883);
and U5401 (N_5401,N_4786,N_5047);
xnor U5402 (N_5402,N_5153,N_4606);
or U5403 (N_5403,N_4945,N_4712);
nor U5404 (N_5404,N_4835,N_4992);
nor U5405 (N_5405,N_4646,N_5121);
nor U5406 (N_5406,N_5176,N_4653);
and U5407 (N_5407,N_4691,N_4790);
xor U5408 (N_5408,N_4557,N_4618);
or U5409 (N_5409,N_4532,N_4834);
nor U5410 (N_5410,N_4595,N_5025);
nand U5411 (N_5411,N_4509,N_4620);
xor U5412 (N_5412,N_4694,N_4538);
or U5413 (N_5413,N_4648,N_5063);
nor U5414 (N_5414,N_4871,N_4735);
or U5415 (N_5415,N_4870,N_4773);
or U5416 (N_5416,N_5090,N_4612);
xnor U5417 (N_5417,N_4565,N_4526);
nand U5418 (N_5418,N_4683,N_5055);
and U5419 (N_5419,N_4885,N_5167);
nand U5420 (N_5420,N_4920,N_4570);
nor U5421 (N_5421,N_4865,N_4705);
or U5422 (N_5422,N_4868,N_4964);
nand U5423 (N_5423,N_5104,N_4762);
or U5424 (N_5424,N_4609,N_4737);
nor U5425 (N_5425,N_4731,N_4984);
xnor U5426 (N_5426,N_5078,N_5229);
nand U5427 (N_5427,N_4797,N_4626);
nor U5428 (N_5428,N_5240,N_4988);
and U5429 (N_5429,N_4904,N_4710);
or U5430 (N_5430,N_5041,N_4858);
nor U5431 (N_5431,N_5115,N_4780);
or U5432 (N_5432,N_5127,N_4994);
nand U5433 (N_5433,N_4923,N_5220);
xnor U5434 (N_5434,N_5172,N_4937);
nor U5435 (N_5435,N_5155,N_5087);
and U5436 (N_5436,N_4634,N_4953);
xnor U5437 (N_5437,N_4562,N_4892);
xor U5438 (N_5438,N_4558,N_4951);
or U5439 (N_5439,N_4830,N_4952);
nor U5440 (N_5440,N_5005,N_5150);
nor U5441 (N_5441,N_4903,N_4823);
or U5442 (N_5442,N_4801,N_4598);
xor U5443 (N_5443,N_4622,N_4651);
xor U5444 (N_5444,N_4617,N_4670);
nor U5445 (N_5445,N_5214,N_4963);
and U5446 (N_5446,N_5075,N_4877);
xor U5447 (N_5447,N_4922,N_5102);
nor U5448 (N_5448,N_4502,N_5033);
xor U5449 (N_5449,N_4575,N_4889);
xor U5450 (N_5450,N_4827,N_5120);
xor U5451 (N_5451,N_5223,N_4503);
or U5452 (N_5452,N_4943,N_4978);
and U5453 (N_5453,N_4859,N_4836);
and U5454 (N_5454,N_4852,N_5144);
nand U5455 (N_5455,N_5113,N_4701);
and U5456 (N_5456,N_4514,N_4804);
xor U5457 (N_5457,N_5204,N_5061);
xor U5458 (N_5458,N_4591,N_4776);
and U5459 (N_5459,N_5143,N_4803);
and U5460 (N_5460,N_4807,N_4706);
nor U5461 (N_5461,N_4583,N_5210);
xor U5462 (N_5462,N_4781,N_4635);
xor U5463 (N_5463,N_4555,N_4603);
and U5464 (N_5464,N_5130,N_4908);
or U5465 (N_5465,N_4531,N_5065);
and U5466 (N_5466,N_4898,N_4542);
xnor U5467 (N_5467,N_4914,N_5196);
nor U5468 (N_5468,N_5241,N_5003);
and U5469 (N_5469,N_4686,N_5207);
nor U5470 (N_5470,N_4665,N_5234);
nand U5471 (N_5471,N_4824,N_4714);
and U5472 (N_5472,N_5197,N_5002);
xor U5473 (N_5473,N_5026,N_4659);
or U5474 (N_5474,N_4887,N_4650);
and U5475 (N_5475,N_4896,N_4975);
nand U5476 (N_5476,N_4690,N_5004);
and U5477 (N_5477,N_5095,N_5194);
nor U5478 (N_5478,N_4993,N_4907);
or U5479 (N_5479,N_5211,N_5110);
nand U5480 (N_5480,N_4547,N_5225);
and U5481 (N_5481,N_5107,N_5174);
or U5482 (N_5482,N_4525,N_4556);
and U5483 (N_5483,N_5236,N_4613);
nand U5484 (N_5484,N_5008,N_4832);
xnor U5485 (N_5485,N_5177,N_4721);
nor U5486 (N_5486,N_5112,N_5020);
or U5487 (N_5487,N_4507,N_4770);
and U5488 (N_5488,N_5239,N_4821);
or U5489 (N_5489,N_4534,N_5027);
and U5490 (N_5490,N_4966,N_5182);
nor U5491 (N_5491,N_5082,N_5175);
and U5492 (N_5492,N_5187,N_4552);
or U5493 (N_5493,N_4974,N_4787);
nor U5494 (N_5494,N_4637,N_4713);
nand U5495 (N_5495,N_4607,N_5228);
or U5496 (N_5496,N_4693,N_4711);
nor U5497 (N_5497,N_5128,N_4510);
nor U5498 (N_5498,N_5086,N_4733);
nand U5499 (N_5499,N_5195,N_5044);
xnor U5500 (N_5500,N_4861,N_4678);
or U5501 (N_5501,N_4523,N_5021);
nand U5502 (N_5502,N_4630,N_4500);
and U5503 (N_5503,N_5007,N_4674);
and U5504 (N_5504,N_4854,N_4553);
nor U5505 (N_5505,N_4545,N_4970);
nor U5506 (N_5506,N_5119,N_4533);
nand U5507 (N_5507,N_4905,N_5073);
and U5508 (N_5508,N_5006,N_4982);
nor U5509 (N_5509,N_5133,N_4755);
xnor U5510 (N_5510,N_4643,N_4972);
and U5511 (N_5511,N_5232,N_4515);
nor U5512 (N_5512,N_4676,N_4777);
nand U5513 (N_5513,N_4879,N_5201);
or U5514 (N_5514,N_4600,N_4971);
xnor U5515 (N_5515,N_4716,N_4928);
nor U5516 (N_5516,N_4881,N_5154);
xnor U5517 (N_5517,N_4669,N_4795);
or U5518 (N_5518,N_4541,N_5203);
xor U5519 (N_5519,N_4611,N_5106);
nand U5520 (N_5520,N_4708,N_4991);
and U5521 (N_5521,N_4925,N_4715);
or U5522 (N_5522,N_5160,N_4862);
or U5523 (N_5523,N_4680,N_5052);
and U5524 (N_5524,N_5051,N_5224);
nor U5525 (N_5525,N_4962,N_4911);
nor U5526 (N_5526,N_4576,N_5076);
nor U5527 (N_5527,N_4704,N_4860);
or U5528 (N_5528,N_5168,N_4685);
or U5529 (N_5529,N_4989,N_5179);
xnor U5530 (N_5530,N_4916,N_5074);
or U5531 (N_5531,N_5243,N_5209);
xnor U5532 (N_5532,N_4899,N_5045);
nand U5533 (N_5533,N_5146,N_4849);
nand U5534 (N_5534,N_4519,N_4977);
and U5535 (N_5535,N_4996,N_4884);
and U5536 (N_5536,N_5028,N_4619);
xnor U5537 (N_5537,N_5108,N_4818);
xnor U5538 (N_5538,N_4687,N_4902);
xnor U5539 (N_5539,N_4997,N_4671);
xor U5540 (N_5540,N_5158,N_4844);
and U5541 (N_5541,N_4842,N_4934);
xor U5542 (N_5542,N_4511,N_5099);
or U5543 (N_5543,N_4751,N_4880);
xor U5544 (N_5544,N_4906,N_4957);
xor U5545 (N_5545,N_4791,N_4535);
or U5546 (N_5546,N_4938,N_4654);
xor U5547 (N_5547,N_4811,N_4725);
xnor U5548 (N_5548,N_4540,N_4900);
and U5549 (N_5549,N_5071,N_4568);
nand U5550 (N_5550,N_4756,N_4946);
xnor U5551 (N_5551,N_5022,N_4940);
and U5552 (N_5552,N_4582,N_4662);
and U5553 (N_5553,N_4753,N_4809);
nor U5554 (N_5554,N_4947,N_4551);
nor U5555 (N_5555,N_4508,N_4792);
nand U5556 (N_5556,N_4973,N_5126);
nand U5557 (N_5557,N_4544,N_4739);
or U5558 (N_5558,N_4730,N_4802);
and U5559 (N_5559,N_5054,N_4655);
nor U5560 (N_5560,N_4505,N_5169);
or U5561 (N_5561,N_4894,N_5037);
and U5562 (N_5562,N_5139,N_5093);
and U5563 (N_5563,N_5040,N_4817);
nand U5564 (N_5564,N_4759,N_4890);
nor U5565 (N_5565,N_4625,N_4765);
nor U5566 (N_5566,N_5018,N_4915);
xnor U5567 (N_5567,N_5122,N_4833);
xnor U5568 (N_5568,N_4688,N_4942);
nand U5569 (N_5569,N_4554,N_4936);
and U5570 (N_5570,N_5142,N_5081);
and U5571 (N_5571,N_4841,N_4658);
xor U5572 (N_5572,N_4587,N_5117);
and U5573 (N_5573,N_4610,N_4839);
or U5574 (N_5574,N_4738,N_4955);
and U5575 (N_5575,N_5012,N_4632);
xnor U5576 (N_5576,N_4785,N_4631);
nand U5577 (N_5577,N_4736,N_4527);
nor U5578 (N_5578,N_4960,N_5192);
nand U5579 (N_5579,N_4999,N_5136);
or U5580 (N_5580,N_4521,N_4864);
or U5581 (N_5581,N_5149,N_4764);
xor U5582 (N_5582,N_4524,N_5235);
or U5583 (N_5583,N_5072,N_4661);
or U5584 (N_5584,N_4752,N_4539);
and U5585 (N_5585,N_4939,N_5111);
nand U5586 (N_5586,N_4604,N_4550);
xnor U5587 (N_5587,N_5070,N_4597);
nand U5588 (N_5588,N_4910,N_5066);
or U5589 (N_5589,N_4760,N_4763);
nor U5590 (N_5590,N_4935,N_4644);
and U5591 (N_5591,N_5039,N_4647);
and U5592 (N_5592,N_4564,N_4578);
or U5593 (N_5593,N_4717,N_5035);
and U5594 (N_5594,N_5069,N_4636);
and U5595 (N_5595,N_5034,N_4629);
xnor U5596 (N_5596,N_4729,N_4518);
nand U5597 (N_5597,N_4590,N_4536);
nor U5598 (N_5598,N_4743,N_4528);
nor U5599 (N_5599,N_4959,N_4718);
nor U5600 (N_5600,N_4771,N_4863);
nand U5601 (N_5601,N_5088,N_4624);
and U5602 (N_5602,N_4969,N_4513);
and U5603 (N_5603,N_4543,N_4601);
or U5604 (N_5604,N_5042,N_4709);
and U5605 (N_5605,N_4985,N_4700);
and U5606 (N_5606,N_5049,N_4749);
and U5607 (N_5607,N_5000,N_4748);
or U5608 (N_5608,N_4855,N_4919);
nor U5609 (N_5609,N_4652,N_4976);
nor U5610 (N_5610,N_4788,N_4572);
or U5611 (N_5611,N_5170,N_4628);
xor U5612 (N_5612,N_4569,N_4697);
nand U5613 (N_5613,N_4761,N_4805);
xor U5614 (N_5614,N_5064,N_4516);
and U5615 (N_5615,N_5151,N_5048);
nor U5616 (N_5616,N_4589,N_4956);
or U5617 (N_5617,N_5213,N_4563);
or U5618 (N_5618,N_4638,N_4886);
nand U5619 (N_5619,N_4848,N_4689);
xnor U5620 (N_5620,N_4621,N_4901);
nor U5621 (N_5621,N_5014,N_5218);
xnor U5622 (N_5622,N_5103,N_5198);
nor U5623 (N_5623,N_4723,N_4990);
nor U5624 (N_5624,N_5019,N_4581);
and U5625 (N_5625,N_4992,N_4930);
or U5626 (N_5626,N_5064,N_4943);
nor U5627 (N_5627,N_4663,N_4956);
and U5628 (N_5628,N_5142,N_5096);
and U5629 (N_5629,N_5119,N_4939);
nor U5630 (N_5630,N_4701,N_4751);
nand U5631 (N_5631,N_5115,N_5086);
nor U5632 (N_5632,N_5020,N_4893);
nand U5633 (N_5633,N_5244,N_5161);
or U5634 (N_5634,N_4775,N_4686);
and U5635 (N_5635,N_4596,N_4855);
nor U5636 (N_5636,N_4671,N_4916);
and U5637 (N_5637,N_5031,N_4730);
nand U5638 (N_5638,N_5042,N_4859);
nand U5639 (N_5639,N_4596,N_5202);
nand U5640 (N_5640,N_4502,N_4827);
or U5641 (N_5641,N_5101,N_5168);
and U5642 (N_5642,N_4573,N_4501);
nand U5643 (N_5643,N_4986,N_4849);
nand U5644 (N_5644,N_4540,N_5170);
or U5645 (N_5645,N_4922,N_4939);
nand U5646 (N_5646,N_4515,N_5191);
or U5647 (N_5647,N_4794,N_5094);
nand U5648 (N_5648,N_5180,N_4725);
or U5649 (N_5649,N_5090,N_4859);
nor U5650 (N_5650,N_5039,N_5134);
nand U5651 (N_5651,N_4534,N_4613);
and U5652 (N_5652,N_5007,N_4652);
or U5653 (N_5653,N_4763,N_4643);
and U5654 (N_5654,N_4915,N_4600);
nor U5655 (N_5655,N_4821,N_4774);
or U5656 (N_5656,N_4733,N_4547);
or U5657 (N_5657,N_4734,N_4686);
nand U5658 (N_5658,N_4648,N_4662);
xor U5659 (N_5659,N_4794,N_4925);
xor U5660 (N_5660,N_4520,N_4922);
or U5661 (N_5661,N_4874,N_5188);
nand U5662 (N_5662,N_4643,N_5157);
nand U5663 (N_5663,N_4838,N_4935);
nand U5664 (N_5664,N_4809,N_4935);
and U5665 (N_5665,N_4846,N_4943);
and U5666 (N_5666,N_4516,N_4897);
and U5667 (N_5667,N_5211,N_5118);
xor U5668 (N_5668,N_4891,N_4900);
and U5669 (N_5669,N_5175,N_4840);
nand U5670 (N_5670,N_4992,N_5053);
xnor U5671 (N_5671,N_4550,N_4531);
nand U5672 (N_5672,N_4915,N_4988);
or U5673 (N_5673,N_4899,N_4798);
nand U5674 (N_5674,N_4760,N_5104);
nor U5675 (N_5675,N_4778,N_4595);
xor U5676 (N_5676,N_4946,N_5006);
and U5677 (N_5677,N_4501,N_5127);
and U5678 (N_5678,N_4868,N_5205);
or U5679 (N_5679,N_4980,N_4929);
nand U5680 (N_5680,N_5013,N_4892);
and U5681 (N_5681,N_4743,N_4588);
nor U5682 (N_5682,N_4554,N_4695);
xor U5683 (N_5683,N_5155,N_4597);
nand U5684 (N_5684,N_4979,N_4697);
and U5685 (N_5685,N_5006,N_4615);
or U5686 (N_5686,N_4884,N_5117);
nor U5687 (N_5687,N_4587,N_4733);
nor U5688 (N_5688,N_4567,N_4582);
and U5689 (N_5689,N_5070,N_4527);
or U5690 (N_5690,N_4940,N_4740);
and U5691 (N_5691,N_4965,N_5120);
and U5692 (N_5692,N_4750,N_4679);
xor U5693 (N_5693,N_5156,N_5225);
nor U5694 (N_5694,N_4664,N_4730);
and U5695 (N_5695,N_4938,N_4860);
nand U5696 (N_5696,N_4606,N_4916);
nor U5697 (N_5697,N_5172,N_4534);
nand U5698 (N_5698,N_4817,N_4828);
nor U5699 (N_5699,N_5141,N_4638);
or U5700 (N_5700,N_4688,N_4678);
nand U5701 (N_5701,N_4636,N_4828);
xor U5702 (N_5702,N_4586,N_4601);
and U5703 (N_5703,N_4907,N_5066);
and U5704 (N_5704,N_5196,N_5132);
nand U5705 (N_5705,N_4573,N_5188);
nand U5706 (N_5706,N_4707,N_4584);
xor U5707 (N_5707,N_4533,N_5006);
nor U5708 (N_5708,N_4972,N_4887);
nand U5709 (N_5709,N_4697,N_4576);
nand U5710 (N_5710,N_4599,N_4641);
or U5711 (N_5711,N_4902,N_4805);
and U5712 (N_5712,N_5238,N_5129);
and U5713 (N_5713,N_4625,N_5005);
or U5714 (N_5714,N_4978,N_4671);
xor U5715 (N_5715,N_4963,N_4840);
nand U5716 (N_5716,N_5248,N_4522);
or U5717 (N_5717,N_4920,N_5054);
nand U5718 (N_5718,N_5180,N_4728);
nand U5719 (N_5719,N_4510,N_4526);
and U5720 (N_5720,N_5231,N_4811);
or U5721 (N_5721,N_4744,N_4923);
nor U5722 (N_5722,N_4685,N_4949);
nor U5723 (N_5723,N_4519,N_5102);
and U5724 (N_5724,N_4555,N_4913);
xor U5725 (N_5725,N_4865,N_5162);
nand U5726 (N_5726,N_4568,N_4612);
xnor U5727 (N_5727,N_5243,N_4694);
and U5728 (N_5728,N_4720,N_4783);
nor U5729 (N_5729,N_4889,N_4755);
or U5730 (N_5730,N_5241,N_5002);
or U5731 (N_5731,N_4969,N_5175);
and U5732 (N_5732,N_5149,N_5023);
xor U5733 (N_5733,N_4942,N_4921);
or U5734 (N_5734,N_4756,N_5101);
xnor U5735 (N_5735,N_4854,N_5222);
or U5736 (N_5736,N_4717,N_4858);
or U5737 (N_5737,N_5099,N_5061);
xor U5738 (N_5738,N_5146,N_5110);
and U5739 (N_5739,N_4699,N_4716);
or U5740 (N_5740,N_5222,N_5242);
and U5741 (N_5741,N_4524,N_4931);
xor U5742 (N_5742,N_5128,N_4738);
nand U5743 (N_5743,N_4610,N_4502);
nor U5744 (N_5744,N_5234,N_4719);
nor U5745 (N_5745,N_4674,N_4604);
nor U5746 (N_5746,N_5244,N_5148);
and U5747 (N_5747,N_4672,N_5228);
and U5748 (N_5748,N_5053,N_4627);
xor U5749 (N_5749,N_4994,N_5038);
xnor U5750 (N_5750,N_5020,N_4878);
and U5751 (N_5751,N_4877,N_4694);
nor U5752 (N_5752,N_5210,N_4814);
nor U5753 (N_5753,N_4804,N_4916);
nand U5754 (N_5754,N_4573,N_4841);
nand U5755 (N_5755,N_4749,N_4761);
and U5756 (N_5756,N_4868,N_4543);
and U5757 (N_5757,N_4762,N_4521);
nor U5758 (N_5758,N_4997,N_5027);
xnor U5759 (N_5759,N_4873,N_5113);
nand U5760 (N_5760,N_5234,N_5042);
nand U5761 (N_5761,N_5025,N_4682);
and U5762 (N_5762,N_5069,N_4818);
and U5763 (N_5763,N_4879,N_4932);
and U5764 (N_5764,N_4834,N_4575);
xor U5765 (N_5765,N_4779,N_4681);
nand U5766 (N_5766,N_5119,N_4767);
nor U5767 (N_5767,N_5155,N_4601);
and U5768 (N_5768,N_4704,N_5049);
nand U5769 (N_5769,N_4540,N_5037);
nor U5770 (N_5770,N_5059,N_4749);
nand U5771 (N_5771,N_4682,N_5053);
and U5772 (N_5772,N_4949,N_4695);
and U5773 (N_5773,N_5058,N_5076);
or U5774 (N_5774,N_4959,N_5219);
and U5775 (N_5775,N_4658,N_5039);
and U5776 (N_5776,N_4750,N_4741);
nand U5777 (N_5777,N_4929,N_4747);
xor U5778 (N_5778,N_4564,N_5202);
nor U5779 (N_5779,N_4701,N_4848);
and U5780 (N_5780,N_4714,N_4972);
nor U5781 (N_5781,N_5197,N_4673);
nor U5782 (N_5782,N_4701,N_4867);
and U5783 (N_5783,N_4566,N_4738);
xnor U5784 (N_5784,N_4596,N_4610);
and U5785 (N_5785,N_4873,N_4749);
nand U5786 (N_5786,N_5213,N_4957);
nand U5787 (N_5787,N_4861,N_4502);
nor U5788 (N_5788,N_5215,N_4593);
nand U5789 (N_5789,N_5248,N_5016);
nor U5790 (N_5790,N_5003,N_5119);
xor U5791 (N_5791,N_5114,N_5107);
nor U5792 (N_5792,N_4934,N_4902);
nor U5793 (N_5793,N_5094,N_4815);
or U5794 (N_5794,N_4781,N_4929);
nand U5795 (N_5795,N_4981,N_4707);
and U5796 (N_5796,N_4775,N_4892);
or U5797 (N_5797,N_5206,N_4809);
and U5798 (N_5798,N_4707,N_4716);
and U5799 (N_5799,N_4900,N_5002);
xnor U5800 (N_5800,N_4570,N_4533);
xor U5801 (N_5801,N_5194,N_5234);
and U5802 (N_5802,N_4646,N_4630);
nor U5803 (N_5803,N_4880,N_4661);
or U5804 (N_5804,N_5005,N_4745);
and U5805 (N_5805,N_5042,N_4926);
and U5806 (N_5806,N_5144,N_4507);
and U5807 (N_5807,N_5204,N_4994);
nor U5808 (N_5808,N_4935,N_4744);
xor U5809 (N_5809,N_4511,N_4961);
or U5810 (N_5810,N_4576,N_4529);
xor U5811 (N_5811,N_4568,N_4859);
or U5812 (N_5812,N_5140,N_4599);
nand U5813 (N_5813,N_4705,N_4517);
xor U5814 (N_5814,N_5195,N_4894);
or U5815 (N_5815,N_4834,N_5221);
nor U5816 (N_5816,N_4736,N_5051);
xor U5817 (N_5817,N_4515,N_4593);
nor U5818 (N_5818,N_5055,N_4523);
nand U5819 (N_5819,N_4826,N_4921);
and U5820 (N_5820,N_4757,N_5187);
and U5821 (N_5821,N_4616,N_4712);
xnor U5822 (N_5822,N_4760,N_5019);
nor U5823 (N_5823,N_4730,N_5086);
nor U5824 (N_5824,N_4680,N_5131);
xnor U5825 (N_5825,N_4972,N_4722);
or U5826 (N_5826,N_5000,N_4830);
and U5827 (N_5827,N_5127,N_5052);
xnor U5828 (N_5828,N_4597,N_5231);
and U5829 (N_5829,N_4939,N_4880);
xor U5830 (N_5830,N_4652,N_4904);
nand U5831 (N_5831,N_4838,N_4870);
nand U5832 (N_5832,N_4895,N_5122);
xor U5833 (N_5833,N_5011,N_4730);
xnor U5834 (N_5834,N_4557,N_4521);
and U5835 (N_5835,N_5048,N_4919);
nand U5836 (N_5836,N_5242,N_4668);
nand U5837 (N_5837,N_5229,N_4997);
nor U5838 (N_5838,N_4980,N_4841);
and U5839 (N_5839,N_5053,N_5203);
or U5840 (N_5840,N_4951,N_4947);
and U5841 (N_5841,N_4621,N_4592);
or U5842 (N_5842,N_5247,N_4920);
nand U5843 (N_5843,N_4633,N_4678);
or U5844 (N_5844,N_5027,N_4787);
xor U5845 (N_5845,N_5094,N_4571);
and U5846 (N_5846,N_4554,N_4919);
nor U5847 (N_5847,N_5146,N_5072);
or U5848 (N_5848,N_5070,N_4958);
xnor U5849 (N_5849,N_5244,N_4895);
nand U5850 (N_5850,N_5203,N_5046);
or U5851 (N_5851,N_5055,N_4791);
or U5852 (N_5852,N_4868,N_4668);
nand U5853 (N_5853,N_4599,N_4967);
nand U5854 (N_5854,N_4555,N_5049);
xnor U5855 (N_5855,N_4847,N_5014);
nand U5856 (N_5856,N_4560,N_4848);
nand U5857 (N_5857,N_4672,N_4905);
nand U5858 (N_5858,N_4510,N_5220);
nor U5859 (N_5859,N_4622,N_4644);
nor U5860 (N_5860,N_5107,N_4578);
nand U5861 (N_5861,N_4590,N_5001);
nor U5862 (N_5862,N_4595,N_4751);
and U5863 (N_5863,N_4981,N_4957);
nand U5864 (N_5864,N_5019,N_5133);
nand U5865 (N_5865,N_4760,N_4717);
xnor U5866 (N_5866,N_4627,N_5054);
and U5867 (N_5867,N_4757,N_4750);
or U5868 (N_5868,N_5108,N_5031);
and U5869 (N_5869,N_5210,N_5034);
and U5870 (N_5870,N_4678,N_5088);
nand U5871 (N_5871,N_5082,N_4668);
xnor U5872 (N_5872,N_4605,N_5099);
and U5873 (N_5873,N_4984,N_4589);
nor U5874 (N_5874,N_5022,N_4589);
nand U5875 (N_5875,N_4855,N_4801);
nand U5876 (N_5876,N_4640,N_5022);
nand U5877 (N_5877,N_4568,N_4797);
xor U5878 (N_5878,N_5158,N_4553);
xnor U5879 (N_5879,N_5209,N_4546);
nand U5880 (N_5880,N_5118,N_4869);
nand U5881 (N_5881,N_4545,N_4731);
nand U5882 (N_5882,N_4723,N_4743);
or U5883 (N_5883,N_4560,N_4855);
nand U5884 (N_5884,N_4601,N_5154);
xor U5885 (N_5885,N_5010,N_5033);
nand U5886 (N_5886,N_4693,N_5024);
nor U5887 (N_5887,N_4948,N_4566);
xnor U5888 (N_5888,N_4853,N_4844);
nand U5889 (N_5889,N_4704,N_4772);
or U5890 (N_5890,N_4978,N_4881);
xor U5891 (N_5891,N_5085,N_5237);
or U5892 (N_5892,N_4569,N_4794);
xor U5893 (N_5893,N_4516,N_4711);
or U5894 (N_5894,N_4510,N_4885);
xnor U5895 (N_5895,N_4580,N_4913);
or U5896 (N_5896,N_5146,N_5091);
xor U5897 (N_5897,N_4610,N_4572);
xor U5898 (N_5898,N_5204,N_5119);
or U5899 (N_5899,N_5084,N_5014);
and U5900 (N_5900,N_4870,N_4741);
and U5901 (N_5901,N_4739,N_5227);
nor U5902 (N_5902,N_5190,N_5219);
nand U5903 (N_5903,N_4586,N_5044);
and U5904 (N_5904,N_5011,N_4678);
xnor U5905 (N_5905,N_5160,N_4916);
xnor U5906 (N_5906,N_4750,N_4985);
xor U5907 (N_5907,N_4629,N_5175);
nand U5908 (N_5908,N_5090,N_5107);
and U5909 (N_5909,N_5050,N_4981);
xor U5910 (N_5910,N_4920,N_4512);
or U5911 (N_5911,N_5111,N_5158);
and U5912 (N_5912,N_4701,N_4595);
nor U5913 (N_5913,N_4899,N_5109);
nor U5914 (N_5914,N_5151,N_4976);
nor U5915 (N_5915,N_5020,N_5018);
nor U5916 (N_5916,N_4543,N_4578);
xor U5917 (N_5917,N_4622,N_5130);
and U5918 (N_5918,N_5102,N_4866);
nand U5919 (N_5919,N_5145,N_4995);
nand U5920 (N_5920,N_5087,N_4758);
xnor U5921 (N_5921,N_4930,N_5091);
and U5922 (N_5922,N_4638,N_4712);
or U5923 (N_5923,N_4764,N_5136);
xnor U5924 (N_5924,N_4766,N_4582);
nand U5925 (N_5925,N_5026,N_5186);
xor U5926 (N_5926,N_4806,N_4804);
or U5927 (N_5927,N_4730,N_5067);
nor U5928 (N_5928,N_5227,N_4786);
nand U5929 (N_5929,N_4506,N_4881);
nand U5930 (N_5930,N_5134,N_5028);
xnor U5931 (N_5931,N_4675,N_5246);
or U5932 (N_5932,N_5200,N_5034);
nor U5933 (N_5933,N_4970,N_5240);
and U5934 (N_5934,N_4968,N_5039);
and U5935 (N_5935,N_4848,N_4598);
and U5936 (N_5936,N_5238,N_5230);
or U5937 (N_5937,N_5242,N_4723);
nand U5938 (N_5938,N_4739,N_4656);
nor U5939 (N_5939,N_4951,N_4507);
xor U5940 (N_5940,N_4759,N_4838);
nand U5941 (N_5941,N_4768,N_5023);
nor U5942 (N_5942,N_4512,N_4899);
xnor U5943 (N_5943,N_4510,N_4572);
nor U5944 (N_5944,N_4798,N_5066);
nand U5945 (N_5945,N_5039,N_5226);
nor U5946 (N_5946,N_4870,N_4942);
nand U5947 (N_5947,N_4952,N_4834);
nor U5948 (N_5948,N_4856,N_5161);
or U5949 (N_5949,N_4827,N_5221);
or U5950 (N_5950,N_4617,N_5168);
xnor U5951 (N_5951,N_4518,N_4597);
and U5952 (N_5952,N_4739,N_5042);
and U5953 (N_5953,N_4957,N_4595);
nor U5954 (N_5954,N_5019,N_4579);
nand U5955 (N_5955,N_4777,N_4557);
nand U5956 (N_5956,N_4926,N_4892);
nor U5957 (N_5957,N_4973,N_5249);
or U5958 (N_5958,N_4859,N_4784);
xor U5959 (N_5959,N_4587,N_5111);
and U5960 (N_5960,N_4906,N_5121);
or U5961 (N_5961,N_5015,N_4633);
and U5962 (N_5962,N_4850,N_5180);
xnor U5963 (N_5963,N_5131,N_4867);
nor U5964 (N_5964,N_4740,N_4759);
and U5965 (N_5965,N_4700,N_5001);
and U5966 (N_5966,N_5130,N_4779);
nand U5967 (N_5967,N_5199,N_4866);
nor U5968 (N_5968,N_4894,N_5134);
nor U5969 (N_5969,N_4742,N_4673);
or U5970 (N_5970,N_4984,N_5007);
xnor U5971 (N_5971,N_4516,N_4555);
nand U5972 (N_5972,N_5009,N_4829);
xor U5973 (N_5973,N_5217,N_4558);
or U5974 (N_5974,N_5050,N_4605);
xnor U5975 (N_5975,N_4656,N_5020);
nor U5976 (N_5976,N_4687,N_5098);
or U5977 (N_5977,N_5204,N_4702);
xnor U5978 (N_5978,N_4804,N_4658);
and U5979 (N_5979,N_5151,N_5037);
or U5980 (N_5980,N_5176,N_4801);
nor U5981 (N_5981,N_5066,N_4929);
and U5982 (N_5982,N_5038,N_4631);
or U5983 (N_5983,N_5157,N_4705);
or U5984 (N_5984,N_4636,N_5131);
or U5985 (N_5985,N_4877,N_4594);
and U5986 (N_5986,N_5119,N_4711);
and U5987 (N_5987,N_5133,N_4751);
xor U5988 (N_5988,N_4546,N_4555);
nor U5989 (N_5989,N_5116,N_5120);
or U5990 (N_5990,N_4756,N_5216);
nor U5991 (N_5991,N_4524,N_4811);
and U5992 (N_5992,N_4920,N_4906);
or U5993 (N_5993,N_4944,N_4715);
and U5994 (N_5994,N_4864,N_5027);
xor U5995 (N_5995,N_4965,N_4775);
and U5996 (N_5996,N_5096,N_4985);
nor U5997 (N_5997,N_4636,N_4746);
or U5998 (N_5998,N_5033,N_4764);
and U5999 (N_5999,N_5110,N_5074);
nand U6000 (N_6000,N_5865,N_5873);
or U6001 (N_6001,N_5361,N_5836);
and U6002 (N_6002,N_5421,N_5714);
or U6003 (N_6003,N_5318,N_5300);
xor U6004 (N_6004,N_5552,N_5635);
xnor U6005 (N_6005,N_5584,N_5499);
nand U6006 (N_6006,N_5979,N_5955);
nand U6007 (N_6007,N_5463,N_5471);
and U6008 (N_6008,N_5350,N_5931);
nand U6009 (N_6009,N_5780,N_5653);
and U6010 (N_6010,N_5416,N_5700);
xor U6011 (N_6011,N_5451,N_5682);
xnor U6012 (N_6012,N_5749,N_5371);
nand U6013 (N_6013,N_5947,N_5967);
nand U6014 (N_6014,N_5397,N_5852);
nor U6015 (N_6015,N_5440,N_5418);
or U6016 (N_6016,N_5442,N_5790);
or U6017 (N_6017,N_5476,N_5285);
and U6018 (N_6018,N_5562,N_5566);
nand U6019 (N_6019,N_5255,N_5385);
xor U6020 (N_6020,N_5405,N_5553);
nor U6021 (N_6021,N_5448,N_5837);
or U6022 (N_6022,N_5815,N_5327);
xor U6023 (N_6023,N_5487,N_5480);
and U6024 (N_6024,N_5830,N_5525);
xor U6025 (N_6025,N_5725,N_5345);
nand U6026 (N_6026,N_5719,N_5274);
or U6027 (N_6027,N_5497,N_5379);
and U6028 (N_6028,N_5690,N_5520);
and U6029 (N_6029,N_5764,N_5641);
nor U6030 (N_6030,N_5608,N_5329);
or U6031 (N_6031,N_5828,N_5298);
xnor U6032 (N_6032,N_5545,N_5752);
xor U6033 (N_6033,N_5351,N_5378);
nand U6034 (N_6034,N_5945,N_5962);
nand U6035 (N_6035,N_5370,N_5992);
xnor U6036 (N_6036,N_5718,N_5796);
or U6037 (N_6037,N_5860,N_5994);
and U6038 (N_6038,N_5661,N_5910);
nor U6039 (N_6039,N_5841,N_5973);
or U6040 (N_6040,N_5468,N_5565);
xor U6041 (N_6041,N_5941,N_5976);
and U6042 (N_6042,N_5920,N_5786);
or U6043 (N_6043,N_5623,N_5891);
xor U6044 (N_6044,N_5369,N_5443);
and U6045 (N_6045,N_5722,N_5301);
nor U6046 (N_6046,N_5358,N_5490);
xor U6047 (N_6047,N_5498,N_5573);
and U6048 (N_6048,N_5612,N_5995);
or U6049 (N_6049,N_5568,N_5377);
nand U6050 (N_6050,N_5754,N_5362);
xnor U6051 (N_6051,N_5744,N_5289);
and U6052 (N_6052,N_5696,N_5892);
nand U6053 (N_6053,N_5311,N_5341);
nand U6054 (N_6054,N_5742,N_5849);
or U6055 (N_6055,N_5436,N_5328);
xnor U6056 (N_6056,N_5807,N_5654);
xor U6057 (N_6057,N_5262,N_5750);
xnor U6058 (N_6058,N_5425,N_5676);
nor U6059 (N_6059,N_5509,N_5856);
and U6060 (N_6060,N_5558,N_5561);
xnor U6061 (N_6061,N_5901,N_5616);
or U6062 (N_6062,N_5532,N_5672);
xnor U6063 (N_6063,N_5619,N_5768);
xor U6064 (N_6064,N_5814,N_5803);
and U6065 (N_6065,N_5896,N_5555);
and U6066 (N_6066,N_5581,N_5646);
or U6067 (N_6067,N_5634,N_5333);
nand U6068 (N_6068,N_5611,N_5567);
nor U6069 (N_6069,N_5829,N_5863);
or U6070 (N_6070,N_5670,N_5326);
or U6071 (N_6071,N_5753,N_5374);
and U6072 (N_6072,N_5337,N_5512);
or U6073 (N_6073,N_5938,N_5867);
or U6074 (N_6074,N_5927,N_5677);
nand U6075 (N_6075,N_5316,N_5999);
nand U6076 (N_6076,N_5946,N_5913);
nand U6077 (N_6077,N_5866,N_5514);
nand U6078 (N_6078,N_5348,N_5441);
nand U6079 (N_6079,N_5346,N_5275);
xnor U6080 (N_6080,N_5404,N_5368);
or U6081 (N_6081,N_5877,N_5844);
nor U6082 (N_6082,N_5642,N_5669);
or U6083 (N_6083,N_5615,N_5782);
and U6084 (N_6084,N_5317,N_5906);
nand U6085 (N_6085,N_5446,N_5762);
nand U6086 (N_6086,N_5688,N_5985);
nand U6087 (N_6087,N_5821,N_5548);
nor U6088 (N_6088,N_5689,N_5705);
nor U6089 (N_6089,N_5384,N_5338);
and U6090 (N_6090,N_5554,N_5465);
xnor U6091 (N_6091,N_5438,N_5734);
and U6092 (N_6092,N_5632,N_5454);
xnor U6093 (N_6093,N_5622,N_5953);
xor U6094 (N_6094,N_5702,N_5657);
nor U6095 (N_6095,N_5998,N_5388);
and U6096 (N_6096,N_5776,N_5420);
or U6097 (N_6097,N_5427,N_5492);
or U6098 (N_6098,N_5745,N_5406);
xor U6099 (N_6099,N_5957,N_5709);
xnor U6100 (N_6100,N_5894,N_5578);
nor U6101 (N_6101,N_5987,N_5680);
xor U6102 (N_6102,N_5902,N_5854);
or U6103 (N_6103,N_5574,N_5504);
nor U6104 (N_6104,N_5767,N_5850);
and U6105 (N_6105,N_5305,N_5394);
nor U6106 (N_6106,N_5312,N_5472);
nand U6107 (N_6107,N_5740,N_5602);
and U6108 (N_6108,N_5570,N_5510);
nor U6109 (N_6109,N_5543,N_5726);
xor U6110 (N_6110,N_5820,N_5899);
nor U6111 (N_6111,N_5452,N_5989);
nand U6112 (N_6112,N_5536,N_5589);
or U6113 (N_6113,N_5538,N_5339);
nand U6114 (N_6114,N_5952,N_5868);
or U6115 (N_6115,N_5785,N_5970);
or U6116 (N_6116,N_5335,N_5625);
nand U6117 (N_6117,N_5610,N_5271);
or U6118 (N_6118,N_5883,N_5518);
xnor U6119 (N_6119,N_5469,N_5295);
and U6120 (N_6120,N_5626,N_5769);
xnor U6121 (N_6121,N_5478,N_5942);
and U6122 (N_6122,N_5278,N_5569);
and U6123 (N_6123,N_5503,N_5884);
nand U6124 (N_6124,N_5864,N_5889);
nand U6125 (N_6125,N_5323,N_5784);
nand U6126 (N_6126,N_5313,N_5809);
and U6127 (N_6127,N_5280,N_5445);
and U6128 (N_6128,N_5297,N_5517);
xnor U6129 (N_6129,N_5412,N_5834);
and U6130 (N_6130,N_5692,N_5964);
and U6131 (N_6131,N_5426,N_5544);
nand U6132 (N_6132,N_5818,N_5652);
nor U6133 (N_6133,N_5281,N_5359);
xor U6134 (N_6134,N_5251,N_5594);
nor U6135 (N_6135,N_5708,N_5590);
xor U6136 (N_6136,N_5853,N_5325);
or U6137 (N_6137,N_5585,N_5331);
nand U6138 (N_6138,N_5732,N_5467);
or U6139 (N_6139,N_5971,N_5644);
and U6140 (N_6140,N_5876,N_5703);
nor U6141 (N_6141,N_5943,N_5975);
nor U6142 (N_6142,N_5712,N_5332);
or U6143 (N_6143,N_5269,N_5484);
nand U6144 (N_6144,N_5917,N_5758);
and U6145 (N_6145,N_5686,N_5481);
xor U6146 (N_6146,N_5314,N_5748);
or U6147 (N_6147,N_5813,N_5668);
or U6148 (N_6148,N_5811,N_5435);
or U6149 (N_6149,N_5423,N_5905);
xnor U6150 (N_6150,N_5355,N_5344);
or U6151 (N_6151,N_5586,N_5401);
and U6152 (N_6152,N_5546,N_5530);
xnor U6153 (N_6153,N_5766,N_5847);
and U6154 (N_6154,N_5290,N_5729);
nand U6155 (N_6155,N_5598,N_5673);
nand U6156 (N_6156,N_5595,N_5306);
and U6157 (N_6157,N_5851,N_5540);
and U6158 (N_6158,N_5483,N_5717);
or U6159 (N_6159,N_5526,N_5550);
or U6160 (N_6160,N_5888,N_5839);
nand U6161 (N_6161,N_5779,N_5870);
xor U6162 (N_6162,N_5637,N_5432);
nor U6163 (N_6163,N_5960,N_5264);
nand U6164 (N_6164,N_5800,N_5407);
nor U6165 (N_6165,N_5986,N_5933);
nor U6166 (N_6166,N_5287,N_5390);
nand U6167 (N_6167,N_5715,N_5485);
or U6168 (N_6168,N_5254,N_5663);
xor U6169 (N_6169,N_5763,N_5838);
nor U6170 (N_6170,N_5733,N_5523);
or U6171 (N_6171,N_5701,N_5577);
nand U6172 (N_6172,N_5479,N_5721);
xor U6173 (N_6173,N_5267,N_5473);
and U6174 (N_6174,N_5810,N_5618);
or U6175 (N_6175,N_5787,N_5356);
xor U6176 (N_6176,N_5893,N_5462);
nand U6177 (N_6177,N_5997,N_5659);
nand U6178 (N_6178,N_5699,N_5923);
and U6179 (N_6179,N_5541,N_5738);
xnor U6180 (N_6180,N_5831,N_5372);
and U6181 (N_6181,N_5904,N_5458);
and U6182 (N_6182,N_5593,N_5872);
and U6183 (N_6183,N_5835,N_5600);
xnor U6184 (N_6184,N_5772,N_5687);
xor U6185 (N_6185,N_5477,N_5575);
xnor U6186 (N_6186,N_5808,N_5706);
and U6187 (N_6187,N_5367,N_5391);
or U6188 (N_6188,N_5396,N_5324);
and U6189 (N_6189,N_5919,N_5697);
xnor U6190 (N_6190,N_5778,N_5507);
xnor U6191 (N_6191,N_5266,N_5789);
xnor U6192 (N_6192,N_5277,N_5886);
and U6193 (N_6193,N_5797,N_5263);
or U6194 (N_6194,N_5542,N_5879);
nor U6195 (N_6195,N_5691,N_5950);
and U6196 (N_6196,N_5310,N_5293);
xnor U6197 (N_6197,N_5417,N_5909);
or U6198 (N_6198,N_5430,N_5607);
or U6199 (N_6199,N_5456,N_5392);
or U6200 (N_6200,N_5320,N_5505);
xnor U6201 (N_6201,N_5832,N_5671);
nand U6202 (N_6202,N_5373,N_5674);
xor U6203 (N_6203,N_5424,N_5783);
xnor U6204 (N_6204,N_5439,N_5887);
and U6205 (N_6205,N_5824,N_5980);
nand U6206 (N_6206,N_5648,N_5609);
and U6207 (N_6207,N_5897,N_5400);
or U6208 (N_6208,N_5282,N_5825);
and U6209 (N_6209,N_5963,N_5730);
and U6210 (N_6210,N_5294,N_5665);
and U6211 (N_6211,N_5951,N_5991);
and U6212 (N_6212,N_5982,N_5583);
and U6213 (N_6213,N_5929,N_5954);
xor U6214 (N_6214,N_5827,N_5823);
and U6215 (N_6215,N_5912,N_5636);
xnor U6216 (N_6216,N_5524,N_5628);
nand U6217 (N_6217,N_5798,N_5679);
nand U6218 (N_6218,N_5268,N_5592);
or U6219 (N_6219,N_5793,N_5795);
xor U6220 (N_6220,N_5655,N_5539);
and U6221 (N_6221,N_5775,N_5258);
nor U6222 (N_6222,N_5513,N_5502);
and U6223 (N_6223,N_5747,N_5756);
and U6224 (N_6224,N_5981,N_5840);
nand U6225 (N_6225,N_5630,N_5788);
and U6226 (N_6226,N_5252,N_5460);
xnor U6227 (N_6227,N_5930,N_5645);
and U6228 (N_6228,N_5296,N_5587);
and U6229 (N_6229,N_5474,N_5489);
xor U6230 (N_6230,N_5988,N_5871);
and U6231 (N_6231,N_5916,N_5723);
nor U6232 (N_6232,N_5261,N_5681);
nor U6233 (N_6233,N_5650,N_5869);
nor U6234 (N_6234,N_5398,N_5382);
and U6235 (N_6235,N_5966,N_5651);
nor U6236 (N_6236,N_5433,N_5649);
nor U6237 (N_6237,N_5256,N_5855);
nor U6238 (N_6238,N_5253,N_5531);
or U6239 (N_6239,N_5667,N_5534);
xnor U6240 (N_6240,N_5434,N_5903);
xnor U6241 (N_6241,N_5826,N_5560);
or U6242 (N_6242,N_5773,N_5386);
nand U6243 (N_6243,N_5805,N_5940);
and U6244 (N_6244,N_5944,N_5878);
and U6245 (N_6245,N_5647,N_5961);
nor U6246 (N_6246,N_5354,N_5969);
nand U6247 (N_6247,N_5959,N_5349);
xnor U6248 (N_6248,N_5340,N_5322);
or U6249 (N_6249,N_5363,N_5631);
xor U6250 (N_6250,N_5704,N_5292);
nand U6251 (N_6251,N_5932,N_5627);
xnor U6252 (N_6252,N_5447,N_5496);
nand U6253 (N_6253,N_5336,N_5875);
nand U6254 (N_6254,N_5259,N_5413);
xor U6255 (N_6255,N_5547,N_5403);
and U6256 (N_6256,N_5713,N_5410);
and U6257 (N_6257,N_5928,N_5308);
nor U6258 (N_6258,N_5968,N_5770);
and U6259 (N_6259,N_5664,N_5731);
or U6260 (N_6260,N_5812,N_5457);
or U6261 (N_6261,N_5716,N_5605);
nand U6262 (N_6262,N_5279,N_5614);
nor U6263 (N_6263,N_5486,N_5741);
xor U6264 (N_6264,N_5303,N_5735);
xor U6265 (N_6265,N_5728,N_5521);
and U6266 (N_6266,N_5761,N_5914);
and U6267 (N_6267,N_5792,N_5848);
and U6268 (N_6268,N_5684,N_5972);
or U6269 (N_6269,N_5934,N_5765);
or U6270 (N_6270,N_5360,N_5307);
nand U6271 (N_6271,N_5470,N_5760);
nand U6272 (N_6272,N_5529,N_5613);
or U6273 (N_6273,N_5816,N_5774);
nor U6274 (N_6274,N_5675,N_5694);
and U6275 (N_6275,N_5389,N_5908);
xor U6276 (N_6276,N_5660,N_5501);
nand U6277 (N_6277,N_5475,N_5978);
nor U6278 (N_6278,N_5414,N_5408);
and U6279 (N_6279,N_5482,N_5949);
or U6280 (N_6280,N_5707,N_5381);
nor U6281 (N_6281,N_5522,N_5315);
nand U6282 (N_6282,N_5958,N_5781);
and U6283 (N_6283,N_5596,N_5387);
and U6284 (N_6284,N_5495,N_5617);
nand U6285 (N_6285,N_5399,N_5500);
nand U6286 (N_6286,N_5260,N_5343);
nor U6287 (N_6287,N_5597,N_5422);
or U6288 (N_6288,N_5819,N_5376);
and U6289 (N_6289,N_5563,N_5739);
and U6290 (N_6290,N_5857,N_5624);
and U6291 (N_6291,N_5450,N_5250);
or U6292 (N_6292,N_5845,N_5366);
nand U6293 (N_6293,N_5683,N_5859);
nand U6294 (N_6294,N_5288,N_5582);
nor U6295 (N_6295,N_5265,N_5506);
and U6296 (N_6296,N_5273,N_5572);
nor U6297 (N_6297,N_5334,N_5640);
xnor U6298 (N_6298,N_5757,N_5977);
nor U6299 (N_6299,N_5915,N_5347);
nor U6300 (N_6300,N_5606,N_5299);
and U6301 (N_6301,N_5270,N_5291);
nor U6302 (N_6302,N_5309,N_5535);
nor U6303 (N_6303,N_5755,N_5519);
nand U6304 (N_6304,N_5409,N_5579);
and U6305 (N_6305,N_5419,N_5638);
nor U6306 (N_6306,N_5759,N_5357);
xnor U6307 (N_6307,N_5528,N_5353);
and U6308 (N_6308,N_5918,N_5556);
and U6309 (N_6309,N_5629,N_5633);
nand U6310 (N_6310,N_5678,N_5571);
xor U6311 (N_6311,N_5777,N_5656);
nand U6312 (N_6312,N_5736,N_5411);
or U6313 (N_6313,N_5461,N_5576);
nand U6314 (N_6314,N_5907,N_5580);
nor U6315 (N_6315,N_5428,N_5993);
xor U6316 (N_6316,N_5319,N_5990);
and U6317 (N_6317,N_5415,N_5806);
nand U6318 (N_6318,N_5257,N_5603);
or U6319 (N_6319,N_5874,N_5453);
xor U6320 (N_6320,N_5794,N_5533);
xnor U6321 (N_6321,N_5685,N_5383);
nor U6322 (N_6322,N_5455,N_5983);
and U6323 (N_6323,N_5284,N_5984);
or U6324 (N_6324,N_5639,N_5895);
and U6325 (N_6325,N_5861,N_5936);
xor U6326 (N_6326,N_5304,N_5516);
nand U6327 (N_6327,N_5488,N_5921);
nand U6328 (N_6328,N_5737,N_5621);
and U6329 (N_6329,N_5286,N_5843);
nand U6330 (N_6330,N_5515,N_5604);
or U6331 (N_6331,N_5746,N_5666);
nor U6332 (N_6332,N_5276,N_5466);
and U6333 (N_6333,N_5527,N_5551);
or U6334 (N_6334,N_5493,N_5925);
and U6335 (N_6335,N_5491,N_5935);
xor U6336 (N_6336,N_5429,N_5771);
xor U6337 (N_6337,N_5375,N_5444);
or U6338 (N_6338,N_5431,N_5922);
and U6339 (N_6339,N_5710,N_5464);
and U6340 (N_6340,N_5822,N_5833);
or U6341 (N_6341,N_5693,N_5342);
nor U6342 (N_6342,N_5862,N_5791);
nand U6343 (N_6343,N_5996,N_5395);
nand U6344 (N_6344,N_5885,N_5564);
and U6345 (N_6345,N_5620,N_5662);
nand U6346 (N_6346,N_5364,N_5437);
nor U6347 (N_6347,N_5882,N_5711);
nor U6348 (N_6348,N_5743,N_5846);
or U6349 (N_6349,N_5402,N_5924);
xor U6350 (N_6350,N_5937,N_5549);
nand U6351 (N_6351,N_5658,N_5393);
xor U6352 (N_6352,N_5817,N_5751);
and U6353 (N_6353,N_5974,N_5449);
or U6354 (N_6354,N_5494,N_5321);
or U6355 (N_6355,N_5559,N_5643);
xor U6356 (N_6356,N_5880,N_5591);
nor U6357 (N_6357,N_5956,N_5557);
nand U6358 (N_6358,N_5890,N_5283);
and U6359 (N_6359,N_5601,N_5799);
xnor U6360 (N_6360,N_5365,N_5727);
and U6361 (N_6361,N_5858,N_5802);
xor U6362 (N_6362,N_5881,N_5508);
xnor U6363 (N_6363,N_5352,N_5926);
or U6364 (N_6364,N_5965,N_5801);
and U6365 (N_6365,N_5898,N_5804);
nand U6366 (N_6366,N_5272,N_5330);
or U6367 (N_6367,N_5698,N_5939);
and U6368 (N_6368,N_5724,N_5537);
nor U6369 (N_6369,N_5911,N_5459);
nand U6370 (N_6370,N_5948,N_5900);
nor U6371 (N_6371,N_5302,N_5720);
and U6372 (N_6372,N_5842,N_5511);
or U6373 (N_6373,N_5380,N_5599);
and U6374 (N_6374,N_5695,N_5588);
and U6375 (N_6375,N_5859,N_5362);
nor U6376 (N_6376,N_5700,N_5574);
and U6377 (N_6377,N_5534,N_5268);
or U6378 (N_6378,N_5280,N_5639);
nand U6379 (N_6379,N_5298,N_5267);
and U6380 (N_6380,N_5477,N_5952);
and U6381 (N_6381,N_5467,N_5435);
nand U6382 (N_6382,N_5568,N_5261);
xnor U6383 (N_6383,N_5380,N_5725);
and U6384 (N_6384,N_5362,N_5473);
and U6385 (N_6385,N_5927,N_5990);
or U6386 (N_6386,N_5700,N_5787);
xnor U6387 (N_6387,N_5856,N_5579);
nor U6388 (N_6388,N_5851,N_5872);
nand U6389 (N_6389,N_5969,N_5463);
nand U6390 (N_6390,N_5926,N_5414);
xnor U6391 (N_6391,N_5372,N_5536);
and U6392 (N_6392,N_5717,N_5825);
nand U6393 (N_6393,N_5779,N_5548);
xor U6394 (N_6394,N_5505,N_5252);
nor U6395 (N_6395,N_5636,N_5876);
nor U6396 (N_6396,N_5977,N_5365);
nor U6397 (N_6397,N_5403,N_5419);
and U6398 (N_6398,N_5969,N_5555);
xnor U6399 (N_6399,N_5270,N_5660);
and U6400 (N_6400,N_5551,N_5651);
and U6401 (N_6401,N_5832,N_5419);
and U6402 (N_6402,N_5355,N_5696);
or U6403 (N_6403,N_5309,N_5693);
nor U6404 (N_6404,N_5702,N_5820);
nor U6405 (N_6405,N_5431,N_5766);
nand U6406 (N_6406,N_5811,N_5533);
xnor U6407 (N_6407,N_5662,N_5693);
xnor U6408 (N_6408,N_5888,N_5674);
xor U6409 (N_6409,N_5684,N_5777);
or U6410 (N_6410,N_5820,N_5938);
or U6411 (N_6411,N_5870,N_5842);
and U6412 (N_6412,N_5420,N_5909);
nand U6413 (N_6413,N_5565,N_5946);
and U6414 (N_6414,N_5980,N_5807);
xor U6415 (N_6415,N_5298,N_5443);
and U6416 (N_6416,N_5786,N_5692);
xnor U6417 (N_6417,N_5626,N_5764);
nor U6418 (N_6418,N_5713,N_5560);
nor U6419 (N_6419,N_5901,N_5845);
or U6420 (N_6420,N_5329,N_5500);
and U6421 (N_6421,N_5290,N_5774);
nand U6422 (N_6422,N_5667,N_5978);
nor U6423 (N_6423,N_5866,N_5841);
and U6424 (N_6424,N_5688,N_5810);
and U6425 (N_6425,N_5407,N_5556);
xor U6426 (N_6426,N_5490,N_5408);
xor U6427 (N_6427,N_5808,N_5301);
or U6428 (N_6428,N_5437,N_5252);
nand U6429 (N_6429,N_5890,N_5298);
and U6430 (N_6430,N_5377,N_5809);
and U6431 (N_6431,N_5509,N_5654);
and U6432 (N_6432,N_5721,N_5589);
or U6433 (N_6433,N_5996,N_5905);
xnor U6434 (N_6434,N_5576,N_5310);
nor U6435 (N_6435,N_5463,N_5547);
xor U6436 (N_6436,N_5705,N_5880);
and U6437 (N_6437,N_5912,N_5745);
and U6438 (N_6438,N_5805,N_5269);
and U6439 (N_6439,N_5460,N_5274);
and U6440 (N_6440,N_5613,N_5811);
or U6441 (N_6441,N_5287,N_5885);
or U6442 (N_6442,N_5620,N_5381);
xor U6443 (N_6443,N_5463,N_5449);
nand U6444 (N_6444,N_5782,N_5683);
and U6445 (N_6445,N_5320,N_5839);
nand U6446 (N_6446,N_5831,N_5554);
xnor U6447 (N_6447,N_5908,N_5381);
or U6448 (N_6448,N_5909,N_5858);
and U6449 (N_6449,N_5251,N_5743);
nor U6450 (N_6450,N_5935,N_5689);
nand U6451 (N_6451,N_5900,N_5506);
or U6452 (N_6452,N_5445,N_5423);
or U6453 (N_6453,N_5976,N_5753);
or U6454 (N_6454,N_5420,N_5958);
nor U6455 (N_6455,N_5788,N_5724);
nor U6456 (N_6456,N_5278,N_5965);
and U6457 (N_6457,N_5792,N_5346);
and U6458 (N_6458,N_5988,N_5640);
nor U6459 (N_6459,N_5279,N_5340);
and U6460 (N_6460,N_5914,N_5656);
nand U6461 (N_6461,N_5772,N_5779);
nand U6462 (N_6462,N_5832,N_5409);
and U6463 (N_6463,N_5436,N_5747);
xnor U6464 (N_6464,N_5945,N_5640);
and U6465 (N_6465,N_5325,N_5387);
nand U6466 (N_6466,N_5997,N_5980);
and U6467 (N_6467,N_5460,N_5562);
nand U6468 (N_6468,N_5640,N_5757);
or U6469 (N_6469,N_5967,N_5389);
nor U6470 (N_6470,N_5926,N_5872);
or U6471 (N_6471,N_5792,N_5332);
nand U6472 (N_6472,N_5423,N_5630);
nor U6473 (N_6473,N_5325,N_5665);
or U6474 (N_6474,N_5540,N_5606);
xnor U6475 (N_6475,N_5871,N_5476);
or U6476 (N_6476,N_5795,N_5732);
or U6477 (N_6477,N_5441,N_5912);
or U6478 (N_6478,N_5997,N_5368);
xor U6479 (N_6479,N_5946,N_5853);
nor U6480 (N_6480,N_5641,N_5651);
nand U6481 (N_6481,N_5499,N_5392);
xnor U6482 (N_6482,N_5395,N_5462);
and U6483 (N_6483,N_5706,N_5858);
or U6484 (N_6484,N_5905,N_5720);
nand U6485 (N_6485,N_5339,N_5720);
and U6486 (N_6486,N_5913,N_5787);
xnor U6487 (N_6487,N_5281,N_5536);
or U6488 (N_6488,N_5475,N_5796);
nor U6489 (N_6489,N_5738,N_5403);
xnor U6490 (N_6490,N_5336,N_5469);
or U6491 (N_6491,N_5764,N_5943);
or U6492 (N_6492,N_5923,N_5575);
or U6493 (N_6493,N_5858,N_5886);
and U6494 (N_6494,N_5988,N_5566);
nand U6495 (N_6495,N_5767,N_5300);
or U6496 (N_6496,N_5449,N_5518);
nand U6497 (N_6497,N_5323,N_5676);
nor U6498 (N_6498,N_5312,N_5809);
or U6499 (N_6499,N_5766,N_5812);
nand U6500 (N_6500,N_5701,N_5529);
xor U6501 (N_6501,N_5635,N_5993);
nor U6502 (N_6502,N_5949,N_5431);
nor U6503 (N_6503,N_5346,N_5900);
and U6504 (N_6504,N_5913,N_5944);
or U6505 (N_6505,N_5808,N_5884);
xnor U6506 (N_6506,N_5639,N_5607);
and U6507 (N_6507,N_5686,N_5565);
or U6508 (N_6508,N_5964,N_5536);
and U6509 (N_6509,N_5858,N_5682);
xnor U6510 (N_6510,N_5720,N_5813);
or U6511 (N_6511,N_5879,N_5420);
nor U6512 (N_6512,N_5500,N_5292);
nand U6513 (N_6513,N_5374,N_5808);
xnor U6514 (N_6514,N_5942,N_5871);
nor U6515 (N_6515,N_5571,N_5982);
nand U6516 (N_6516,N_5594,N_5802);
nor U6517 (N_6517,N_5254,N_5821);
xnor U6518 (N_6518,N_5750,N_5616);
nand U6519 (N_6519,N_5488,N_5324);
xnor U6520 (N_6520,N_5334,N_5857);
and U6521 (N_6521,N_5968,N_5749);
nand U6522 (N_6522,N_5713,N_5980);
nor U6523 (N_6523,N_5471,N_5712);
nand U6524 (N_6524,N_5642,N_5992);
and U6525 (N_6525,N_5693,N_5932);
and U6526 (N_6526,N_5994,N_5912);
or U6527 (N_6527,N_5997,N_5490);
nor U6528 (N_6528,N_5895,N_5867);
or U6529 (N_6529,N_5729,N_5564);
and U6530 (N_6530,N_5495,N_5634);
nor U6531 (N_6531,N_5416,N_5254);
xnor U6532 (N_6532,N_5632,N_5592);
and U6533 (N_6533,N_5359,N_5931);
nand U6534 (N_6534,N_5254,N_5992);
and U6535 (N_6535,N_5727,N_5766);
and U6536 (N_6536,N_5488,N_5779);
nand U6537 (N_6537,N_5318,N_5462);
and U6538 (N_6538,N_5576,N_5375);
or U6539 (N_6539,N_5868,N_5698);
or U6540 (N_6540,N_5370,N_5845);
nor U6541 (N_6541,N_5921,N_5735);
xor U6542 (N_6542,N_5530,N_5759);
or U6543 (N_6543,N_5768,N_5740);
and U6544 (N_6544,N_5656,N_5795);
nor U6545 (N_6545,N_5934,N_5993);
nand U6546 (N_6546,N_5825,N_5876);
xor U6547 (N_6547,N_5778,N_5853);
and U6548 (N_6548,N_5639,N_5603);
or U6549 (N_6549,N_5873,N_5600);
or U6550 (N_6550,N_5741,N_5727);
nand U6551 (N_6551,N_5270,N_5930);
and U6552 (N_6552,N_5514,N_5651);
and U6553 (N_6553,N_5404,N_5619);
or U6554 (N_6554,N_5696,N_5705);
nand U6555 (N_6555,N_5422,N_5428);
and U6556 (N_6556,N_5660,N_5376);
or U6557 (N_6557,N_5955,N_5874);
nand U6558 (N_6558,N_5258,N_5765);
and U6559 (N_6559,N_5967,N_5979);
and U6560 (N_6560,N_5264,N_5861);
or U6561 (N_6561,N_5632,N_5294);
nand U6562 (N_6562,N_5781,N_5990);
nor U6563 (N_6563,N_5446,N_5458);
nand U6564 (N_6564,N_5641,N_5738);
nor U6565 (N_6565,N_5364,N_5633);
or U6566 (N_6566,N_5654,N_5764);
or U6567 (N_6567,N_5986,N_5399);
nor U6568 (N_6568,N_5844,N_5913);
nor U6569 (N_6569,N_5849,N_5905);
xnor U6570 (N_6570,N_5447,N_5697);
nand U6571 (N_6571,N_5266,N_5455);
nand U6572 (N_6572,N_5597,N_5366);
or U6573 (N_6573,N_5657,N_5910);
nor U6574 (N_6574,N_5712,N_5938);
and U6575 (N_6575,N_5411,N_5663);
or U6576 (N_6576,N_5283,N_5756);
xor U6577 (N_6577,N_5298,N_5915);
xnor U6578 (N_6578,N_5309,N_5410);
nor U6579 (N_6579,N_5284,N_5391);
nand U6580 (N_6580,N_5892,N_5559);
and U6581 (N_6581,N_5258,N_5766);
xnor U6582 (N_6582,N_5683,N_5431);
xnor U6583 (N_6583,N_5847,N_5784);
and U6584 (N_6584,N_5250,N_5343);
or U6585 (N_6585,N_5769,N_5918);
nand U6586 (N_6586,N_5537,N_5786);
or U6587 (N_6587,N_5316,N_5596);
nand U6588 (N_6588,N_5357,N_5273);
xor U6589 (N_6589,N_5862,N_5339);
and U6590 (N_6590,N_5465,N_5837);
nand U6591 (N_6591,N_5476,N_5653);
nand U6592 (N_6592,N_5567,N_5602);
or U6593 (N_6593,N_5854,N_5476);
nor U6594 (N_6594,N_5767,N_5499);
nor U6595 (N_6595,N_5692,N_5391);
nor U6596 (N_6596,N_5749,N_5923);
nor U6597 (N_6597,N_5809,N_5350);
xnor U6598 (N_6598,N_5613,N_5816);
nand U6599 (N_6599,N_5864,N_5761);
and U6600 (N_6600,N_5413,N_5323);
and U6601 (N_6601,N_5373,N_5941);
nor U6602 (N_6602,N_5530,N_5588);
and U6603 (N_6603,N_5372,N_5405);
or U6604 (N_6604,N_5715,N_5580);
nor U6605 (N_6605,N_5618,N_5505);
nand U6606 (N_6606,N_5393,N_5328);
xnor U6607 (N_6607,N_5680,N_5670);
nand U6608 (N_6608,N_5516,N_5486);
nor U6609 (N_6609,N_5707,N_5582);
nand U6610 (N_6610,N_5573,N_5927);
or U6611 (N_6611,N_5365,N_5799);
and U6612 (N_6612,N_5817,N_5939);
nor U6613 (N_6613,N_5558,N_5409);
or U6614 (N_6614,N_5317,N_5616);
xor U6615 (N_6615,N_5350,N_5639);
nor U6616 (N_6616,N_5972,N_5544);
xnor U6617 (N_6617,N_5554,N_5266);
nor U6618 (N_6618,N_5830,N_5841);
and U6619 (N_6619,N_5535,N_5328);
or U6620 (N_6620,N_5555,N_5318);
and U6621 (N_6621,N_5699,N_5520);
nand U6622 (N_6622,N_5761,N_5600);
xnor U6623 (N_6623,N_5807,N_5831);
xnor U6624 (N_6624,N_5598,N_5360);
and U6625 (N_6625,N_5711,N_5741);
and U6626 (N_6626,N_5915,N_5870);
xor U6627 (N_6627,N_5265,N_5737);
and U6628 (N_6628,N_5391,N_5397);
and U6629 (N_6629,N_5370,N_5842);
xnor U6630 (N_6630,N_5261,N_5320);
or U6631 (N_6631,N_5478,N_5665);
or U6632 (N_6632,N_5283,N_5470);
nor U6633 (N_6633,N_5628,N_5539);
or U6634 (N_6634,N_5940,N_5838);
or U6635 (N_6635,N_5434,N_5942);
nor U6636 (N_6636,N_5565,N_5743);
nand U6637 (N_6637,N_5369,N_5476);
or U6638 (N_6638,N_5643,N_5942);
xnor U6639 (N_6639,N_5541,N_5359);
or U6640 (N_6640,N_5582,N_5639);
nor U6641 (N_6641,N_5761,N_5501);
nor U6642 (N_6642,N_5873,N_5898);
or U6643 (N_6643,N_5490,N_5415);
xor U6644 (N_6644,N_5989,N_5573);
and U6645 (N_6645,N_5859,N_5931);
or U6646 (N_6646,N_5899,N_5616);
nor U6647 (N_6647,N_5872,N_5465);
xor U6648 (N_6648,N_5719,N_5538);
and U6649 (N_6649,N_5436,N_5762);
xnor U6650 (N_6650,N_5395,N_5382);
nand U6651 (N_6651,N_5464,N_5669);
and U6652 (N_6652,N_5691,N_5615);
nand U6653 (N_6653,N_5512,N_5279);
and U6654 (N_6654,N_5345,N_5923);
or U6655 (N_6655,N_5531,N_5877);
nand U6656 (N_6656,N_5482,N_5721);
or U6657 (N_6657,N_5299,N_5956);
or U6658 (N_6658,N_5357,N_5785);
nor U6659 (N_6659,N_5601,N_5556);
nor U6660 (N_6660,N_5748,N_5635);
nor U6661 (N_6661,N_5828,N_5597);
nand U6662 (N_6662,N_5517,N_5509);
nand U6663 (N_6663,N_5707,N_5797);
nand U6664 (N_6664,N_5533,N_5613);
nand U6665 (N_6665,N_5324,N_5783);
xnor U6666 (N_6666,N_5843,N_5485);
and U6667 (N_6667,N_5334,N_5579);
or U6668 (N_6668,N_5678,N_5708);
xor U6669 (N_6669,N_5254,N_5264);
nand U6670 (N_6670,N_5751,N_5911);
nor U6671 (N_6671,N_5370,N_5814);
or U6672 (N_6672,N_5947,N_5647);
nand U6673 (N_6673,N_5629,N_5787);
xor U6674 (N_6674,N_5295,N_5766);
nor U6675 (N_6675,N_5955,N_5756);
xor U6676 (N_6676,N_5960,N_5353);
xor U6677 (N_6677,N_5627,N_5497);
or U6678 (N_6678,N_5629,N_5810);
nor U6679 (N_6679,N_5681,N_5412);
or U6680 (N_6680,N_5298,N_5297);
and U6681 (N_6681,N_5872,N_5391);
nand U6682 (N_6682,N_5800,N_5422);
nor U6683 (N_6683,N_5496,N_5407);
nand U6684 (N_6684,N_5685,N_5608);
nand U6685 (N_6685,N_5317,N_5554);
xnor U6686 (N_6686,N_5387,N_5919);
nor U6687 (N_6687,N_5893,N_5666);
nand U6688 (N_6688,N_5716,N_5262);
xnor U6689 (N_6689,N_5590,N_5648);
nand U6690 (N_6690,N_5844,N_5507);
nor U6691 (N_6691,N_5747,N_5901);
nand U6692 (N_6692,N_5958,N_5384);
nand U6693 (N_6693,N_5991,N_5645);
nand U6694 (N_6694,N_5434,N_5475);
nand U6695 (N_6695,N_5291,N_5417);
nor U6696 (N_6696,N_5904,N_5322);
nand U6697 (N_6697,N_5326,N_5809);
or U6698 (N_6698,N_5295,N_5472);
or U6699 (N_6699,N_5287,N_5863);
nand U6700 (N_6700,N_5675,N_5547);
nand U6701 (N_6701,N_5876,N_5269);
and U6702 (N_6702,N_5520,N_5963);
or U6703 (N_6703,N_5564,N_5293);
xnor U6704 (N_6704,N_5364,N_5883);
nor U6705 (N_6705,N_5824,N_5663);
xnor U6706 (N_6706,N_5521,N_5494);
xor U6707 (N_6707,N_5730,N_5777);
xnor U6708 (N_6708,N_5863,N_5665);
xnor U6709 (N_6709,N_5422,N_5806);
nand U6710 (N_6710,N_5668,N_5910);
nand U6711 (N_6711,N_5690,N_5379);
xor U6712 (N_6712,N_5524,N_5446);
or U6713 (N_6713,N_5646,N_5289);
nor U6714 (N_6714,N_5587,N_5377);
or U6715 (N_6715,N_5844,N_5881);
and U6716 (N_6716,N_5327,N_5442);
and U6717 (N_6717,N_5311,N_5851);
and U6718 (N_6718,N_5801,N_5869);
nand U6719 (N_6719,N_5359,N_5647);
nor U6720 (N_6720,N_5433,N_5793);
and U6721 (N_6721,N_5388,N_5997);
and U6722 (N_6722,N_5349,N_5716);
nand U6723 (N_6723,N_5511,N_5720);
nand U6724 (N_6724,N_5255,N_5905);
or U6725 (N_6725,N_5376,N_5804);
xnor U6726 (N_6726,N_5347,N_5495);
nand U6727 (N_6727,N_5619,N_5302);
nand U6728 (N_6728,N_5559,N_5417);
nor U6729 (N_6729,N_5940,N_5533);
nand U6730 (N_6730,N_5754,N_5402);
xnor U6731 (N_6731,N_5505,N_5644);
nor U6732 (N_6732,N_5829,N_5760);
xnor U6733 (N_6733,N_5610,N_5959);
nor U6734 (N_6734,N_5577,N_5551);
nand U6735 (N_6735,N_5960,N_5701);
nand U6736 (N_6736,N_5259,N_5639);
or U6737 (N_6737,N_5921,N_5587);
and U6738 (N_6738,N_5717,N_5777);
or U6739 (N_6739,N_5672,N_5735);
or U6740 (N_6740,N_5725,N_5764);
or U6741 (N_6741,N_5697,N_5789);
or U6742 (N_6742,N_5605,N_5472);
and U6743 (N_6743,N_5963,N_5896);
and U6744 (N_6744,N_5271,N_5477);
and U6745 (N_6745,N_5570,N_5626);
nor U6746 (N_6746,N_5607,N_5930);
nor U6747 (N_6747,N_5317,N_5573);
nor U6748 (N_6748,N_5706,N_5346);
or U6749 (N_6749,N_5674,N_5462);
or U6750 (N_6750,N_6525,N_6561);
and U6751 (N_6751,N_6482,N_6650);
nand U6752 (N_6752,N_6740,N_6474);
and U6753 (N_6753,N_6660,N_6504);
nor U6754 (N_6754,N_6193,N_6331);
and U6755 (N_6755,N_6116,N_6015);
xnor U6756 (N_6756,N_6320,N_6487);
xor U6757 (N_6757,N_6510,N_6004);
or U6758 (N_6758,N_6665,N_6053);
or U6759 (N_6759,N_6663,N_6018);
nand U6760 (N_6760,N_6566,N_6257);
or U6761 (N_6761,N_6301,N_6600);
nor U6762 (N_6762,N_6213,N_6233);
and U6763 (N_6763,N_6730,N_6059);
or U6764 (N_6764,N_6542,N_6154);
xor U6765 (N_6765,N_6286,N_6009);
and U6766 (N_6766,N_6473,N_6584);
nand U6767 (N_6767,N_6447,N_6611);
nor U6768 (N_6768,N_6393,N_6071);
or U6769 (N_6769,N_6676,N_6242);
or U6770 (N_6770,N_6515,N_6028);
or U6771 (N_6771,N_6248,N_6014);
and U6772 (N_6772,N_6545,N_6489);
xnor U6773 (N_6773,N_6404,N_6132);
xnor U6774 (N_6774,N_6118,N_6604);
and U6775 (N_6775,N_6190,N_6728);
nor U6776 (N_6776,N_6606,N_6067);
nor U6777 (N_6777,N_6125,N_6544);
xor U6778 (N_6778,N_6044,N_6319);
nand U6779 (N_6779,N_6051,N_6653);
nor U6780 (N_6780,N_6005,N_6572);
nor U6781 (N_6781,N_6078,N_6289);
and U6782 (N_6782,N_6210,N_6052);
nor U6783 (N_6783,N_6098,N_6690);
and U6784 (N_6784,N_6141,N_6207);
xor U6785 (N_6785,N_6326,N_6469);
nor U6786 (N_6786,N_6072,N_6436);
or U6787 (N_6787,N_6491,N_6434);
nand U6788 (N_6788,N_6266,N_6414);
or U6789 (N_6789,N_6505,N_6008);
xnor U6790 (N_6790,N_6430,N_6106);
or U6791 (N_6791,N_6494,N_6252);
nor U6792 (N_6792,N_6462,N_6003);
or U6793 (N_6793,N_6138,N_6022);
nor U6794 (N_6794,N_6256,N_6222);
and U6795 (N_6795,N_6657,N_6696);
nor U6796 (N_6796,N_6457,N_6527);
or U6797 (N_6797,N_6365,N_6490);
or U6798 (N_6798,N_6360,N_6297);
nor U6799 (N_6799,N_6073,N_6038);
and U6800 (N_6800,N_6380,N_6352);
nand U6801 (N_6801,N_6047,N_6145);
or U6802 (N_6802,N_6272,N_6361);
nor U6803 (N_6803,N_6199,N_6020);
or U6804 (N_6804,N_6721,N_6423);
nand U6805 (N_6805,N_6672,N_6529);
and U6806 (N_6806,N_6415,N_6149);
and U6807 (N_6807,N_6565,N_6006);
or U6808 (N_6808,N_6277,N_6726);
nand U6809 (N_6809,N_6244,N_6559);
xor U6810 (N_6810,N_6049,N_6587);
and U6811 (N_6811,N_6736,N_6001);
xnor U6812 (N_6812,N_6610,N_6732);
xnor U6813 (N_6813,N_6113,N_6707);
and U6814 (N_6814,N_6713,N_6570);
nor U6815 (N_6815,N_6479,N_6114);
nand U6816 (N_6816,N_6029,N_6431);
nand U6817 (N_6817,N_6183,N_6498);
or U6818 (N_6818,N_6523,N_6030);
or U6819 (N_6819,N_6115,N_6481);
nor U6820 (N_6820,N_6236,N_6450);
and U6821 (N_6821,N_6167,N_6605);
or U6822 (N_6822,N_6658,N_6539);
xnor U6823 (N_6823,N_6219,N_6249);
nand U6824 (N_6824,N_6276,N_6554);
nor U6825 (N_6825,N_6285,N_6217);
nor U6826 (N_6826,N_6677,N_6321);
or U6827 (N_6827,N_6744,N_6358);
xor U6828 (N_6828,N_6381,N_6101);
or U6829 (N_6829,N_6461,N_6378);
nand U6830 (N_6830,N_6578,N_6151);
or U6831 (N_6831,N_6061,N_6274);
xor U6832 (N_6832,N_6254,N_6485);
and U6833 (N_6833,N_6636,N_6367);
nand U6834 (N_6834,N_6045,N_6557);
nor U6835 (N_6835,N_6019,N_6189);
xor U6836 (N_6836,N_6674,N_6577);
xor U6837 (N_6837,N_6172,N_6225);
and U6838 (N_6838,N_6284,N_6466);
xnor U6839 (N_6839,N_6214,N_6122);
nand U6840 (N_6840,N_6643,N_6507);
and U6841 (N_6841,N_6741,N_6405);
nor U6842 (N_6842,N_6234,N_6514);
xnor U6843 (N_6843,N_6619,N_6340);
or U6844 (N_6844,N_6317,N_6614);
nand U6845 (N_6845,N_6435,N_6399);
and U6846 (N_6846,N_6155,N_6120);
and U6847 (N_6847,N_6678,N_6299);
nor U6848 (N_6848,N_6410,N_6085);
nand U6849 (N_6849,N_6448,N_6328);
xor U6850 (N_6850,N_6166,N_6127);
and U6851 (N_6851,N_6452,N_6633);
nor U6852 (N_6852,N_6060,N_6638);
nand U6853 (N_6853,N_6235,N_6548);
xnor U6854 (N_6854,N_6205,N_6264);
and U6855 (N_6855,N_6439,N_6148);
nand U6856 (N_6856,N_6620,N_6041);
xnor U6857 (N_6857,N_6402,N_6621);
or U6858 (N_6858,N_6226,N_6232);
nor U6859 (N_6859,N_6348,N_6691);
nor U6860 (N_6860,N_6395,N_6050);
and U6861 (N_6861,N_6521,N_6699);
nand U6862 (N_6862,N_6412,N_6500);
or U6863 (N_6863,N_6451,N_6188);
nand U6864 (N_6864,N_6247,N_6586);
nand U6865 (N_6865,N_6516,N_6366);
nor U6866 (N_6866,N_6747,N_6720);
nor U6867 (N_6867,N_6419,N_6023);
and U6868 (N_6868,N_6255,N_6099);
and U6869 (N_6869,N_6283,N_6282);
nor U6870 (N_6870,N_6315,N_6314);
nand U6871 (N_6871,N_6520,N_6224);
or U6872 (N_6872,N_6689,N_6243);
and U6873 (N_6873,N_6094,N_6291);
and U6874 (N_6874,N_6409,N_6622);
nand U6875 (N_6875,N_6524,N_6237);
nor U6876 (N_6876,N_6056,N_6540);
nor U6877 (N_6877,N_6074,N_6583);
nand U6878 (N_6878,N_6270,N_6456);
and U6879 (N_6879,N_6316,N_6216);
xor U6880 (N_6880,N_6543,N_6556);
nand U6881 (N_6881,N_6648,N_6576);
xor U6882 (N_6882,N_6356,N_6323);
and U6883 (N_6883,N_6105,N_6704);
xnor U6884 (N_6884,N_6359,N_6344);
xor U6885 (N_6885,N_6631,N_6449);
nor U6886 (N_6886,N_6262,N_6693);
nand U6887 (N_6887,N_6089,N_6341);
nand U6888 (N_6888,N_6590,N_6396);
nor U6889 (N_6889,N_6308,N_6136);
nand U6890 (N_6890,N_6655,N_6594);
nor U6891 (N_6891,N_6722,N_6688);
and U6892 (N_6892,N_6275,N_6734);
nand U6893 (N_6893,N_6519,N_6281);
and U6894 (N_6894,N_6513,N_6311);
nand U6895 (N_6895,N_6706,N_6407);
nor U6896 (N_6896,N_6123,N_6201);
or U6897 (N_6897,N_6338,N_6377);
or U6898 (N_6898,N_6483,N_6669);
nand U6899 (N_6899,N_6342,N_6035);
xor U6900 (N_6900,N_6156,N_6608);
nand U6901 (N_6901,N_6593,N_6013);
nor U6902 (N_6902,N_6077,N_6108);
xor U6903 (N_6903,N_6273,N_6095);
and U6904 (N_6904,N_6468,N_6575);
nand U6905 (N_6905,N_6547,N_6304);
and U6906 (N_6906,N_6066,N_6162);
or U6907 (N_6907,N_6416,N_6422);
nor U6908 (N_6908,N_6421,N_6209);
and U6909 (N_6909,N_6097,N_6629);
xor U6910 (N_6910,N_6687,N_6170);
or U6911 (N_6911,N_6177,N_6695);
or U6912 (N_6912,N_6432,N_6502);
and U6913 (N_6913,N_6686,N_6470);
nor U6914 (N_6914,N_6215,N_6533);
or U6915 (N_6915,N_6692,N_6596);
nand U6916 (N_6916,N_6330,N_6288);
and U6917 (N_6917,N_6160,N_6580);
xnor U6918 (N_6918,N_6347,N_6454);
nor U6919 (N_6919,N_6157,N_6568);
nand U6920 (N_6920,N_6171,N_6159);
xnor U6921 (N_6921,N_6501,N_6639);
xnor U6922 (N_6922,N_6389,N_6163);
nor U6923 (N_6923,N_6144,N_6664);
nor U6924 (N_6924,N_6599,N_6312);
and U6925 (N_6925,N_6346,N_6103);
xnor U6926 (N_6926,N_6685,N_6191);
or U6927 (N_6927,N_6345,N_6265);
nand U6928 (N_6928,N_6362,N_6601);
and U6929 (N_6929,N_6518,N_6385);
nor U6930 (N_6930,N_6198,N_6550);
nand U6931 (N_6931,N_6735,N_6581);
or U6932 (N_6932,N_6534,N_6585);
xor U6933 (N_6933,N_6325,N_6387);
xnor U6934 (N_6934,N_6551,N_6475);
nor U6935 (N_6935,N_6012,N_6438);
xnor U6936 (N_6936,N_6339,N_6032);
and U6937 (N_6937,N_6698,N_6719);
xor U6938 (N_6938,N_6075,N_6091);
nor U6939 (N_6939,N_6709,N_6558);
nor U6940 (N_6940,N_6294,N_6303);
nand U6941 (N_6941,N_6645,N_6058);
xnor U6942 (N_6942,N_6647,N_6086);
nand U6943 (N_6943,N_6040,N_6368);
and U6944 (N_6944,N_6716,N_6522);
xor U6945 (N_6945,N_6202,N_6654);
or U6946 (N_6946,N_6745,N_6128);
xor U6947 (N_6947,N_6253,N_6261);
xor U6948 (N_6948,N_6227,N_6223);
or U6949 (N_6949,N_6287,N_6703);
nor U6950 (N_6950,N_6337,N_6441);
and U6951 (N_6951,N_6024,N_6714);
nor U6952 (N_6952,N_6598,N_6603);
and U6953 (N_6953,N_6589,N_6712);
nand U6954 (N_6954,N_6370,N_6532);
or U6955 (N_6955,N_6147,N_6530);
nand U6956 (N_6956,N_6492,N_6062);
nand U6957 (N_6957,N_6228,N_6503);
and U6958 (N_6958,N_6386,N_6673);
nor U6959 (N_6959,N_6644,N_6129);
nor U6960 (N_6960,N_6406,N_6135);
and U6961 (N_6961,N_6725,N_6618);
or U6962 (N_6962,N_6567,N_6184);
or U6963 (N_6963,N_6239,N_6700);
or U6964 (N_6964,N_6718,N_6302);
xor U6965 (N_6965,N_6652,N_6221);
nor U6966 (N_6966,N_6424,N_6597);
nand U6967 (N_6967,N_6295,N_6659);
nand U6968 (N_6968,N_6528,N_6057);
xor U6969 (N_6969,N_6573,N_6218);
nand U6970 (N_6970,N_6087,N_6371);
and U6971 (N_6971,N_6083,N_6322);
or U6972 (N_6972,N_6306,N_6443);
xor U6973 (N_6973,N_6746,N_6142);
xor U6974 (N_6974,N_6268,N_6175);
nand U6975 (N_6975,N_6446,N_6307);
xnor U6976 (N_6976,N_6104,N_6506);
xor U6977 (N_6977,N_6025,N_6496);
or U6978 (N_6978,N_6168,N_6632);
xnor U6979 (N_6979,N_6333,N_6488);
nor U6980 (N_6980,N_6169,N_6560);
or U6981 (N_6981,N_6382,N_6353);
xor U6982 (N_6982,N_6158,N_6472);
or U6983 (N_6983,N_6705,N_6354);
and U6984 (N_6984,N_6697,N_6511);
or U6985 (N_6985,N_6708,N_6016);
nor U6986 (N_6986,N_6039,N_6426);
xor U6987 (N_6987,N_6240,N_6027);
nor U6988 (N_6988,N_6195,N_6563);
and U6989 (N_6989,N_6335,N_6082);
xor U6990 (N_6990,N_6197,N_6553);
and U6991 (N_6991,N_6437,N_6204);
nor U6992 (N_6992,N_6748,N_6260);
nand U6993 (N_6993,N_6363,N_6220);
or U6994 (N_6994,N_6296,N_6508);
and U6995 (N_6995,N_6666,N_6467);
nand U6996 (N_6996,N_6392,N_6065);
nand U6997 (N_6997,N_6546,N_6139);
nor U6998 (N_6998,N_6310,N_6180);
or U6999 (N_6999,N_6174,N_6549);
xnor U7000 (N_7000,N_6208,N_6379);
xor U7001 (N_7001,N_6192,N_6376);
xor U7002 (N_7002,N_6607,N_6531);
xor U7003 (N_7003,N_6495,N_6609);
xor U7004 (N_7004,N_6634,N_6591);
xor U7005 (N_7005,N_6181,N_6715);
and U7006 (N_7006,N_6290,N_6476);
nor U7007 (N_7007,N_6384,N_6011);
and U7008 (N_7008,N_6034,N_6112);
nand U7009 (N_7009,N_6702,N_6364);
xnor U7010 (N_7010,N_6710,N_6111);
nor U7011 (N_7011,N_6334,N_6043);
nor U7012 (N_7012,N_6143,N_6178);
nand U7013 (N_7013,N_6656,N_6110);
nand U7014 (N_7014,N_6063,N_6497);
or U7015 (N_7015,N_6612,N_6343);
or U7016 (N_7016,N_6512,N_6313);
xnor U7017 (N_7017,N_6574,N_6717);
or U7018 (N_7018,N_6305,N_6683);
xor U7019 (N_7019,N_6121,N_6186);
or U7020 (N_7020,N_6250,N_6048);
nor U7021 (N_7021,N_6246,N_6068);
xor U7022 (N_7022,N_6084,N_6212);
and U7023 (N_7023,N_6153,N_6682);
nor U7024 (N_7024,N_6517,N_6427);
nor U7025 (N_7025,N_6464,N_6667);
and U7026 (N_7026,N_6055,N_6679);
xor U7027 (N_7027,N_6211,N_6231);
nand U7028 (N_7028,N_6592,N_6418);
and U7029 (N_7029,N_6397,N_6133);
nand U7030 (N_7030,N_6007,N_6164);
nand U7031 (N_7031,N_6300,N_6571);
and U7032 (N_7032,N_6743,N_6403);
or U7033 (N_7033,N_6420,N_6642);
or U7034 (N_7034,N_6458,N_6681);
nor U7035 (N_7035,N_6615,N_6017);
and U7036 (N_7036,N_6433,N_6684);
or U7037 (N_7037,N_6258,N_6079);
xor U7038 (N_7038,N_6651,N_6069);
nor U7039 (N_7039,N_6241,N_6613);
nand U7040 (N_7040,N_6411,N_6635);
xor U7041 (N_7041,N_6092,N_6727);
nand U7042 (N_7042,N_6137,N_6499);
or U7043 (N_7043,N_6109,N_6373);
nand U7044 (N_7044,N_6076,N_6538);
nand U7045 (N_7045,N_6054,N_6391);
and U7046 (N_7046,N_6640,N_6729);
nand U7047 (N_7047,N_6298,N_6680);
or U7048 (N_7048,N_6737,N_6429);
or U7049 (N_7049,N_6093,N_6662);
nor U7050 (N_7050,N_6440,N_6460);
nor U7051 (N_7051,N_6327,N_6002);
and U7052 (N_7052,N_6318,N_6046);
or U7053 (N_7053,N_6119,N_6624);
or U7054 (N_7054,N_6292,N_6269);
or U7055 (N_7055,N_6324,N_6185);
nor U7056 (N_7056,N_6671,N_6064);
nand U7057 (N_7057,N_6126,N_6602);
and U7058 (N_7058,N_6271,N_6465);
nand U7059 (N_7059,N_6649,N_6463);
nand U7060 (N_7060,N_6336,N_6628);
nand U7061 (N_7061,N_6357,N_6588);
or U7062 (N_7062,N_6401,N_6388);
nor U7063 (N_7063,N_6021,N_6595);
or U7064 (N_7064,N_6417,N_6131);
nand U7065 (N_7065,N_6230,N_6196);
xnor U7066 (N_7066,N_6161,N_6739);
nand U7067 (N_7067,N_6152,N_6723);
or U7068 (N_7068,N_6187,N_6478);
nand U7069 (N_7069,N_6641,N_6107);
or U7070 (N_7070,N_6579,N_6173);
and U7071 (N_7071,N_6203,N_6675);
nor U7072 (N_7072,N_6455,N_6140);
nand U7073 (N_7073,N_6000,N_6617);
and U7074 (N_7074,N_6130,N_6010);
nand U7075 (N_7075,N_6711,N_6569);
xor U7076 (N_7076,N_6355,N_6425);
or U7077 (N_7077,N_6150,N_6096);
nand U7078 (N_7078,N_6165,N_6245);
or U7079 (N_7079,N_6146,N_6627);
and U7080 (N_7080,N_6102,N_6280);
nand U7081 (N_7081,N_6372,N_6229);
nor U7082 (N_7082,N_6626,N_6637);
xor U7083 (N_7083,N_6279,N_6582);
nor U7084 (N_7084,N_6668,N_6444);
nor U7085 (N_7085,N_6749,N_6070);
or U7086 (N_7086,N_6293,N_6731);
nand U7087 (N_7087,N_6400,N_6349);
or U7088 (N_7088,N_6278,N_6200);
or U7089 (N_7089,N_6117,N_6484);
xor U7090 (N_7090,N_6724,N_6661);
nor U7091 (N_7091,N_6477,N_6670);
and U7092 (N_7092,N_6394,N_6374);
or U7093 (N_7093,N_6537,N_6471);
and U7094 (N_7094,N_6329,N_6134);
or U7095 (N_7095,N_6738,N_6251);
xnor U7096 (N_7096,N_6375,N_6493);
nand U7097 (N_7097,N_6332,N_6616);
nand U7098 (N_7098,N_6206,N_6486);
and U7099 (N_7099,N_6428,N_6625);
or U7100 (N_7100,N_6259,N_6562);
and U7101 (N_7101,N_6445,N_6459);
xnor U7102 (N_7102,N_6701,N_6398);
xnor U7103 (N_7103,N_6453,N_6033);
nand U7104 (N_7104,N_6026,N_6081);
and U7105 (N_7105,N_6555,N_6390);
xor U7106 (N_7106,N_6646,N_6536);
or U7107 (N_7107,N_6623,N_6031);
nor U7108 (N_7108,N_6194,N_6541);
and U7109 (N_7109,N_6733,N_6413);
nand U7110 (N_7110,N_6535,N_6509);
nor U7111 (N_7111,N_6351,N_6369);
nor U7112 (N_7112,N_6350,N_6742);
nor U7113 (N_7113,N_6036,N_6088);
xnor U7114 (N_7114,N_6042,N_6309);
nand U7115 (N_7115,N_6408,N_6100);
nor U7116 (N_7116,N_6182,N_6124);
xnor U7117 (N_7117,N_6090,N_6564);
and U7118 (N_7118,N_6176,N_6238);
xnor U7119 (N_7119,N_6179,N_6383);
nor U7120 (N_7120,N_6263,N_6694);
nor U7121 (N_7121,N_6552,N_6267);
nand U7122 (N_7122,N_6630,N_6526);
or U7123 (N_7123,N_6442,N_6037);
or U7124 (N_7124,N_6080,N_6480);
nor U7125 (N_7125,N_6424,N_6124);
xor U7126 (N_7126,N_6275,N_6378);
nor U7127 (N_7127,N_6083,N_6335);
and U7128 (N_7128,N_6055,N_6694);
and U7129 (N_7129,N_6543,N_6740);
nor U7130 (N_7130,N_6298,N_6395);
nor U7131 (N_7131,N_6374,N_6313);
or U7132 (N_7132,N_6372,N_6013);
nand U7133 (N_7133,N_6337,N_6471);
nor U7134 (N_7134,N_6453,N_6040);
and U7135 (N_7135,N_6090,N_6020);
nand U7136 (N_7136,N_6391,N_6342);
or U7137 (N_7137,N_6382,N_6565);
and U7138 (N_7138,N_6681,N_6231);
and U7139 (N_7139,N_6090,N_6636);
or U7140 (N_7140,N_6716,N_6092);
nor U7141 (N_7141,N_6054,N_6159);
nand U7142 (N_7142,N_6734,N_6017);
xor U7143 (N_7143,N_6480,N_6027);
nand U7144 (N_7144,N_6651,N_6019);
or U7145 (N_7145,N_6576,N_6688);
nor U7146 (N_7146,N_6285,N_6075);
nor U7147 (N_7147,N_6009,N_6724);
xor U7148 (N_7148,N_6046,N_6473);
or U7149 (N_7149,N_6559,N_6066);
nand U7150 (N_7150,N_6087,N_6126);
and U7151 (N_7151,N_6739,N_6547);
nand U7152 (N_7152,N_6254,N_6296);
and U7153 (N_7153,N_6657,N_6184);
and U7154 (N_7154,N_6160,N_6333);
nand U7155 (N_7155,N_6304,N_6420);
nor U7156 (N_7156,N_6262,N_6646);
xnor U7157 (N_7157,N_6033,N_6230);
and U7158 (N_7158,N_6319,N_6391);
or U7159 (N_7159,N_6288,N_6249);
nand U7160 (N_7160,N_6139,N_6677);
nand U7161 (N_7161,N_6442,N_6364);
nor U7162 (N_7162,N_6708,N_6268);
nand U7163 (N_7163,N_6333,N_6606);
and U7164 (N_7164,N_6101,N_6595);
nand U7165 (N_7165,N_6117,N_6706);
or U7166 (N_7166,N_6374,N_6414);
or U7167 (N_7167,N_6221,N_6414);
nor U7168 (N_7168,N_6420,N_6075);
nand U7169 (N_7169,N_6561,N_6142);
nor U7170 (N_7170,N_6404,N_6048);
nor U7171 (N_7171,N_6207,N_6606);
nor U7172 (N_7172,N_6286,N_6031);
xnor U7173 (N_7173,N_6683,N_6186);
and U7174 (N_7174,N_6127,N_6044);
xnor U7175 (N_7175,N_6338,N_6243);
nand U7176 (N_7176,N_6272,N_6457);
and U7177 (N_7177,N_6313,N_6352);
nor U7178 (N_7178,N_6493,N_6519);
and U7179 (N_7179,N_6165,N_6569);
nand U7180 (N_7180,N_6618,N_6510);
nor U7181 (N_7181,N_6728,N_6484);
nand U7182 (N_7182,N_6015,N_6525);
xor U7183 (N_7183,N_6195,N_6716);
xnor U7184 (N_7184,N_6145,N_6148);
and U7185 (N_7185,N_6071,N_6175);
nor U7186 (N_7186,N_6651,N_6668);
nor U7187 (N_7187,N_6310,N_6095);
and U7188 (N_7188,N_6627,N_6488);
xor U7189 (N_7189,N_6414,N_6357);
nand U7190 (N_7190,N_6504,N_6495);
xnor U7191 (N_7191,N_6428,N_6652);
nand U7192 (N_7192,N_6176,N_6599);
and U7193 (N_7193,N_6622,N_6394);
nor U7194 (N_7194,N_6618,N_6738);
and U7195 (N_7195,N_6296,N_6094);
or U7196 (N_7196,N_6500,N_6545);
nand U7197 (N_7197,N_6360,N_6344);
nand U7198 (N_7198,N_6333,N_6001);
nor U7199 (N_7199,N_6726,N_6591);
nor U7200 (N_7200,N_6161,N_6172);
or U7201 (N_7201,N_6517,N_6607);
and U7202 (N_7202,N_6367,N_6180);
nor U7203 (N_7203,N_6164,N_6025);
xnor U7204 (N_7204,N_6092,N_6058);
xor U7205 (N_7205,N_6005,N_6132);
and U7206 (N_7206,N_6220,N_6227);
or U7207 (N_7207,N_6140,N_6489);
and U7208 (N_7208,N_6365,N_6622);
xor U7209 (N_7209,N_6513,N_6089);
xor U7210 (N_7210,N_6160,N_6621);
and U7211 (N_7211,N_6334,N_6532);
nor U7212 (N_7212,N_6607,N_6027);
and U7213 (N_7213,N_6495,N_6312);
nand U7214 (N_7214,N_6186,N_6700);
xor U7215 (N_7215,N_6438,N_6472);
and U7216 (N_7216,N_6391,N_6702);
and U7217 (N_7217,N_6597,N_6612);
xor U7218 (N_7218,N_6480,N_6040);
nor U7219 (N_7219,N_6032,N_6219);
or U7220 (N_7220,N_6233,N_6523);
nor U7221 (N_7221,N_6665,N_6231);
xor U7222 (N_7222,N_6599,N_6722);
or U7223 (N_7223,N_6010,N_6550);
nor U7224 (N_7224,N_6016,N_6579);
nor U7225 (N_7225,N_6282,N_6549);
and U7226 (N_7226,N_6242,N_6314);
nor U7227 (N_7227,N_6552,N_6588);
and U7228 (N_7228,N_6641,N_6561);
xor U7229 (N_7229,N_6571,N_6468);
and U7230 (N_7230,N_6298,N_6208);
nor U7231 (N_7231,N_6251,N_6065);
nand U7232 (N_7232,N_6516,N_6651);
nand U7233 (N_7233,N_6491,N_6147);
nand U7234 (N_7234,N_6266,N_6116);
nand U7235 (N_7235,N_6523,N_6574);
nand U7236 (N_7236,N_6273,N_6047);
nor U7237 (N_7237,N_6161,N_6271);
xor U7238 (N_7238,N_6333,N_6694);
xnor U7239 (N_7239,N_6403,N_6052);
and U7240 (N_7240,N_6246,N_6008);
xnor U7241 (N_7241,N_6594,N_6730);
xnor U7242 (N_7242,N_6496,N_6218);
xor U7243 (N_7243,N_6013,N_6004);
xor U7244 (N_7244,N_6056,N_6087);
nor U7245 (N_7245,N_6345,N_6073);
or U7246 (N_7246,N_6630,N_6521);
and U7247 (N_7247,N_6529,N_6032);
nor U7248 (N_7248,N_6631,N_6132);
nor U7249 (N_7249,N_6544,N_6330);
and U7250 (N_7250,N_6012,N_6081);
xor U7251 (N_7251,N_6592,N_6585);
nand U7252 (N_7252,N_6597,N_6672);
and U7253 (N_7253,N_6274,N_6145);
or U7254 (N_7254,N_6203,N_6663);
or U7255 (N_7255,N_6212,N_6028);
or U7256 (N_7256,N_6677,N_6338);
nand U7257 (N_7257,N_6609,N_6195);
xnor U7258 (N_7258,N_6599,N_6721);
nor U7259 (N_7259,N_6371,N_6104);
and U7260 (N_7260,N_6668,N_6692);
nand U7261 (N_7261,N_6096,N_6629);
nand U7262 (N_7262,N_6248,N_6672);
or U7263 (N_7263,N_6001,N_6324);
or U7264 (N_7264,N_6680,N_6230);
nor U7265 (N_7265,N_6188,N_6311);
or U7266 (N_7266,N_6205,N_6086);
or U7267 (N_7267,N_6704,N_6071);
nor U7268 (N_7268,N_6719,N_6645);
or U7269 (N_7269,N_6590,N_6310);
xnor U7270 (N_7270,N_6429,N_6303);
xor U7271 (N_7271,N_6180,N_6033);
or U7272 (N_7272,N_6102,N_6724);
xnor U7273 (N_7273,N_6101,N_6286);
nand U7274 (N_7274,N_6459,N_6266);
or U7275 (N_7275,N_6647,N_6677);
or U7276 (N_7276,N_6304,N_6288);
xor U7277 (N_7277,N_6613,N_6416);
or U7278 (N_7278,N_6661,N_6279);
nor U7279 (N_7279,N_6608,N_6652);
and U7280 (N_7280,N_6472,N_6023);
and U7281 (N_7281,N_6191,N_6063);
or U7282 (N_7282,N_6198,N_6257);
or U7283 (N_7283,N_6156,N_6108);
nor U7284 (N_7284,N_6259,N_6428);
xor U7285 (N_7285,N_6042,N_6306);
nor U7286 (N_7286,N_6523,N_6483);
xnor U7287 (N_7287,N_6010,N_6199);
nor U7288 (N_7288,N_6044,N_6643);
nor U7289 (N_7289,N_6656,N_6183);
nand U7290 (N_7290,N_6535,N_6593);
nor U7291 (N_7291,N_6740,N_6095);
nor U7292 (N_7292,N_6021,N_6691);
xor U7293 (N_7293,N_6082,N_6118);
and U7294 (N_7294,N_6325,N_6512);
nand U7295 (N_7295,N_6394,N_6107);
and U7296 (N_7296,N_6377,N_6548);
or U7297 (N_7297,N_6227,N_6167);
and U7298 (N_7298,N_6553,N_6659);
nand U7299 (N_7299,N_6628,N_6152);
xor U7300 (N_7300,N_6338,N_6333);
nand U7301 (N_7301,N_6721,N_6700);
nand U7302 (N_7302,N_6698,N_6588);
nand U7303 (N_7303,N_6367,N_6440);
nor U7304 (N_7304,N_6626,N_6257);
and U7305 (N_7305,N_6371,N_6031);
nor U7306 (N_7306,N_6605,N_6105);
and U7307 (N_7307,N_6134,N_6641);
nor U7308 (N_7308,N_6217,N_6604);
and U7309 (N_7309,N_6604,N_6051);
nand U7310 (N_7310,N_6126,N_6343);
or U7311 (N_7311,N_6522,N_6580);
or U7312 (N_7312,N_6064,N_6102);
xor U7313 (N_7313,N_6131,N_6655);
xnor U7314 (N_7314,N_6673,N_6111);
xor U7315 (N_7315,N_6184,N_6749);
or U7316 (N_7316,N_6000,N_6598);
xnor U7317 (N_7317,N_6574,N_6120);
xnor U7318 (N_7318,N_6590,N_6227);
nor U7319 (N_7319,N_6695,N_6482);
xor U7320 (N_7320,N_6258,N_6318);
or U7321 (N_7321,N_6530,N_6214);
xnor U7322 (N_7322,N_6628,N_6457);
nor U7323 (N_7323,N_6705,N_6221);
and U7324 (N_7324,N_6478,N_6139);
nand U7325 (N_7325,N_6154,N_6404);
or U7326 (N_7326,N_6086,N_6157);
and U7327 (N_7327,N_6109,N_6176);
and U7328 (N_7328,N_6590,N_6327);
or U7329 (N_7329,N_6030,N_6586);
nor U7330 (N_7330,N_6326,N_6375);
xnor U7331 (N_7331,N_6612,N_6374);
xor U7332 (N_7332,N_6111,N_6644);
nand U7333 (N_7333,N_6074,N_6601);
nand U7334 (N_7334,N_6177,N_6511);
xor U7335 (N_7335,N_6683,N_6127);
nand U7336 (N_7336,N_6008,N_6407);
and U7337 (N_7337,N_6192,N_6397);
and U7338 (N_7338,N_6437,N_6174);
or U7339 (N_7339,N_6215,N_6049);
and U7340 (N_7340,N_6734,N_6607);
nand U7341 (N_7341,N_6184,N_6159);
nand U7342 (N_7342,N_6170,N_6250);
nand U7343 (N_7343,N_6569,N_6134);
or U7344 (N_7344,N_6274,N_6634);
nor U7345 (N_7345,N_6395,N_6537);
or U7346 (N_7346,N_6011,N_6225);
xnor U7347 (N_7347,N_6413,N_6728);
nand U7348 (N_7348,N_6448,N_6366);
nand U7349 (N_7349,N_6407,N_6364);
and U7350 (N_7350,N_6220,N_6349);
nand U7351 (N_7351,N_6060,N_6692);
and U7352 (N_7352,N_6269,N_6472);
or U7353 (N_7353,N_6080,N_6406);
or U7354 (N_7354,N_6515,N_6078);
xor U7355 (N_7355,N_6422,N_6025);
nand U7356 (N_7356,N_6695,N_6162);
nand U7357 (N_7357,N_6289,N_6061);
xor U7358 (N_7358,N_6260,N_6710);
nor U7359 (N_7359,N_6355,N_6367);
and U7360 (N_7360,N_6116,N_6117);
nand U7361 (N_7361,N_6339,N_6575);
xnor U7362 (N_7362,N_6032,N_6662);
xor U7363 (N_7363,N_6719,N_6726);
or U7364 (N_7364,N_6596,N_6110);
or U7365 (N_7365,N_6497,N_6433);
xnor U7366 (N_7366,N_6576,N_6085);
nor U7367 (N_7367,N_6662,N_6427);
or U7368 (N_7368,N_6394,N_6354);
xnor U7369 (N_7369,N_6495,N_6498);
xor U7370 (N_7370,N_6419,N_6482);
xor U7371 (N_7371,N_6149,N_6425);
nand U7372 (N_7372,N_6054,N_6147);
xor U7373 (N_7373,N_6447,N_6462);
nand U7374 (N_7374,N_6256,N_6523);
xnor U7375 (N_7375,N_6467,N_6011);
nor U7376 (N_7376,N_6126,N_6140);
nand U7377 (N_7377,N_6446,N_6207);
or U7378 (N_7378,N_6693,N_6243);
and U7379 (N_7379,N_6354,N_6091);
nor U7380 (N_7380,N_6083,N_6675);
nor U7381 (N_7381,N_6662,N_6697);
nand U7382 (N_7382,N_6300,N_6630);
nand U7383 (N_7383,N_6307,N_6098);
nor U7384 (N_7384,N_6511,N_6192);
xor U7385 (N_7385,N_6633,N_6625);
nand U7386 (N_7386,N_6704,N_6575);
nand U7387 (N_7387,N_6256,N_6531);
nor U7388 (N_7388,N_6377,N_6125);
or U7389 (N_7389,N_6722,N_6359);
or U7390 (N_7390,N_6115,N_6739);
xnor U7391 (N_7391,N_6385,N_6353);
xnor U7392 (N_7392,N_6450,N_6073);
or U7393 (N_7393,N_6237,N_6339);
nand U7394 (N_7394,N_6407,N_6462);
nor U7395 (N_7395,N_6006,N_6599);
or U7396 (N_7396,N_6640,N_6310);
nand U7397 (N_7397,N_6062,N_6633);
nand U7398 (N_7398,N_6007,N_6650);
nor U7399 (N_7399,N_6541,N_6247);
xnor U7400 (N_7400,N_6634,N_6426);
and U7401 (N_7401,N_6428,N_6517);
nand U7402 (N_7402,N_6178,N_6647);
or U7403 (N_7403,N_6378,N_6313);
and U7404 (N_7404,N_6202,N_6696);
and U7405 (N_7405,N_6618,N_6113);
and U7406 (N_7406,N_6294,N_6360);
nand U7407 (N_7407,N_6590,N_6642);
nand U7408 (N_7408,N_6268,N_6237);
and U7409 (N_7409,N_6483,N_6133);
xnor U7410 (N_7410,N_6464,N_6190);
nand U7411 (N_7411,N_6025,N_6726);
nand U7412 (N_7412,N_6080,N_6216);
xnor U7413 (N_7413,N_6106,N_6675);
xor U7414 (N_7414,N_6674,N_6710);
nor U7415 (N_7415,N_6336,N_6089);
or U7416 (N_7416,N_6652,N_6726);
and U7417 (N_7417,N_6553,N_6205);
xor U7418 (N_7418,N_6345,N_6206);
nor U7419 (N_7419,N_6511,N_6557);
nor U7420 (N_7420,N_6551,N_6035);
or U7421 (N_7421,N_6295,N_6451);
nand U7422 (N_7422,N_6308,N_6249);
nand U7423 (N_7423,N_6178,N_6229);
nand U7424 (N_7424,N_6511,N_6577);
or U7425 (N_7425,N_6442,N_6022);
or U7426 (N_7426,N_6268,N_6549);
nand U7427 (N_7427,N_6586,N_6205);
nand U7428 (N_7428,N_6316,N_6308);
or U7429 (N_7429,N_6267,N_6211);
xor U7430 (N_7430,N_6315,N_6703);
nor U7431 (N_7431,N_6120,N_6456);
nand U7432 (N_7432,N_6722,N_6204);
xor U7433 (N_7433,N_6319,N_6110);
nand U7434 (N_7434,N_6460,N_6029);
xnor U7435 (N_7435,N_6131,N_6533);
nor U7436 (N_7436,N_6321,N_6745);
or U7437 (N_7437,N_6658,N_6010);
and U7438 (N_7438,N_6173,N_6119);
or U7439 (N_7439,N_6171,N_6121);
nand U7440 (N_7440,N_6072,N_6245);
or U7441 (N_7441,N_6376,N_6642);
or U7442 (N_7442,N_6051,N_6245);
xnor U7443 (N_7443,N_6166,N_6260);
or U7444 (N_7444,N_6088,N_6472);
xor U7445 (N_7445,N_6044,N_6491);
or U7446 (N_7446,N_6462,N_6196);
nor U7447 (N_7447,N_6197,N_6561);
nor U7448 (N_7448,N_6510,N_6156);
nand U7449 (N_7449,N_6085,N_6132);
or U7450 (N_7450,N_6745,N_6037);
and U7451 (N_7451,N_6580,N_6575);
nor U7452 (N_7452,N_6142,N_6270);
xor U7453 (N_7453,N_6606,N_6365);
xor U7454 (N_7454,N_6131,N_6554);
or U7455 (N_7455,N_6392,N_6016);
xor U7456 (N_7456,N_6272,N_6001);
nor U7457 (N_7457,N_6467,N_6138);
or U7458 (N_7458,N_6031,N_6091);
nand U7459 (N_7459,N_6590,N_6684);
and U7460 (N_7460,N_6162,N_6454);
nand U7461 (N_7461,N_6170,N_6646);
and U7462 (N_7462,N_6583,N_6375);
nor U7463 (N_7463,N_6568,N_6160);
or U7464 (N_7464,N_6478,N_6285);
nand U7465 (N_7465,N_6367,N_6395);
and U7466 (N_7466,N_6075,N_6022);
xnor U7467 (N_7467,N_6589,N_6488);
or U7468 (N_7468,N_6691,N_6731);
nand U7469 (N_7469,N_6336,N_6692);
nand U7470 (N_7470,N_6273,N_6206);
and U7471 (N_7471,N_6235,N_6439);
nand U7472 (N_7472,N_6396,N_6059);
nand U7473 (N_7473,N_6039,N_6565);
nand U7474 (N_7474,N_6487,N_6131);
nand U7475 (N_7475,N_6652,N_6404);
or U7476 (N_7476,N_6675,N_6560);
nor U7477 (N_7477,N_6708,N_6363);
or U7478 (N_7478,N_6481,N_6059);
xor U7479 (N_7479,N_6136,N_6732);
or U7480 (N_7480,N_6010,N_6738);
and U7481 (N_7481,N_6049,N_6405);
nor U7482 (N_7482,N_6710,N_6298);
nor U7483 (N_7483,N_6270,N_6552);
or U7484 (N_7484,N_6401,N_6231);
or U7485 (N_7485,N_6606,N_6036);
or U7486 (N_7486,N_6317,N_6222);
nand U7487 (N_7487,N_6597,N_6409);
and U7488 (N_7488,N_6043,N_6179);
and U7489 (N_7489,N_6448,N_6194);
nor U7490 (N_7490,N_6322,N_6443);
nor U7491 (N_7491,N_6609,N_6318);
and U7492 (N_7492,N_6727,N_6175);
xor U7493 (N_7493,N_6171,N_6129);
xor U7494 (N_7494,N_6585,N_6018);
xor U7495 (N_7495,N_6731,N_6445);
or U7496 (N_7496,N_6732,N_6320);
nor U7497 (N_7497,N_6516,N_6002);
nand U7498 (N_7498,N_6194,N_6271);
nand U7499 (N_7499,N_6489,N_6142);
and U7500 (N_7500,N_7267,N_6847);
and U7501 (N_7501,N_7170,N_7002);
xnor U7502 (N_7502,N_7275,N_6930);
nor U7503 (N_7503,N_6890,N_7221);
xor U7504 (N_7504,N_7231,N_7158);
and U7505 (N_7505,N_6964,N_7253);
xor U7506 (N_7506,N_6953,N_6863);
nor U7507 (N_7507,N_6905,N_7204);
xor U7508 (N_7508,N_6972,N_7118);
xnor U7509 (N_7509,N_6815,N_6958);
nand U7510 (N_7510,N_7181,N_7058);
xor U7511 (N_7511,N_7168,N_6789);
xnor U7512 (N_7512,N_7139,N_7392);
and U7513 (N_7513,N_6976,N_7124);
or U7514 (N_7514,N_6891,N_6951);
and U7515 (N_7515,N_6817,N_7054);
nor U7516 (N_7516,N_6793,N_7013);
or U7517 (N_7517,N_6756,N_7029);
xnor U7518 (N_7518,N_6894,N_7256);
nand U7519 (N_7519,N_7085,N_7064);
and U7520 (N_7520,N_7127,N_7420);
nor U7521 (N_7521,N_6886,N_7414);
and U7522 (N_7522,N_7070,N_6868);
nand U7523 (N_7523,N_7217,N_6771);
and U7524 (N_7524,N_7192,N_6990);
xnor U7525 (N_7525,N_7095,N_6820);
nand U7526 (N_7526,N_6906,N_6980);
nand U7527 (N_7527,N_7362,N_6968);
nand U7528 (N_7528,N_7093,N_7378);
nand U7529 (N_7529,N_7130,N_7388);
and U7530 (N_7530,N_7012,N_6878);
nand U7531 (N_7531,N_6917,N_6816);
nor U7532 (N_7532,N_7228,N_7298);
nand U7533 (N_7533,N_6804,N_6995);
xor U7534 (N_7534,N_7036,N_7383);
nor U7535 (N_7535,N_7189,N_6773);
nand U7536 (N_7536,N_7358,N_7155);
or U7537 (N_7537,N_6967,N_7385);
and U7538 (N_7538,N_6851,N_6883);
nor U7539 (N_7539,N_7487,N_7235);
nor U7540 (N_7540,N_7238,N_6751);
nand U7541 (N_7541,N_7172,N_6956);
nand U7542 (N_7542,N_7164,N_6795);
nand U7543 (N_7543,N_7131,N_7350);
or U7544 (N_7544,N_7055,N_6943);
and U7545 (N_7545,N_6801,N_7083);
or U7546 (N_7546,N_7038,N_7003);
nor U7547 (N_7547,N_6857,N_7399);
or U7548 (N_7548,N_7101,N_7295);
nor U7549 (N_7549,N_7347,N_6777);
or U7550 (N_7550,N_6937,N_7240);
nand U7551 (N_7551,N_6952,N_6965);
and U7552 (N_7552,N_7318,N_7185);
nor U7553 (N_7553,N_7402,N_7480);
nand U7554 (N_7554,N_7020,N_7272);
nor U7555 (N_7555,N_7497,N_6781);
xnor U7556 (N_7556,N_7308,N_7113);
nor U7557 (N_7557,N_7486,N_7006);
xnor U7558 (N_7558,N_7413,N_6785);
xor U7559 (N_7559,N_7493,N_7452);
nor U7560 (N_7560,N_7367,N_6974);
xnor U7561 (N_7561,N_7326,N_7196);
or U7562 (N_7562,N_7442,N_7255);
nand U7563 (N_7563,N_7111,N_7395);
xor U7564 (N_7564,N_7454,N_7492);
or U7565 (N_7565,N_7068,N_6915);
nand U7566 (N_7566,N_6827,N_6970);
xor U7567 (N_7567,N_7306,N_7075);
nor U7568 (N_7568,N_6760,N_7490);
nor U7569 (N_7569,N_7444,N_7191);
and U7570 (N_7570,N_6860,N_7389);
nor U7571 (N_7571,N_6977,N_6838);
and U7572 (N_7572,N_7425,N_7474);
nand U7573 (N_7573,N_7488,N_7223);
nor U7574 (N_7574,N_7258,N_6918);
xnor U7575 (N_7575,N_7465,N_6866);
nor U7576 (N_7576,N_7129,N_7201);
and U7577 (N_7577,N_7321,N_6767);
nand U7578 (N_7578,N_7063,N_7135);
and U7579 (N_7579,N_6800,N_7432);
and U7580 (N_7580,N_6910,N_6901);
nand U7581 (N_7581,N_7343,N_6837);
and U7582 (N_7582,N_7222,N_7208);
nand U7583 (N_7583,N_7317,N_6790);
or U7584 (N_7584,N_7008,N_7257);
and U7585 (N_7585,N_6911,N_7122);
or U7586 (N_7586,N_7102,N_7180);
xnor U7587 (N_7587,N_6913,N_6830);
or U7588 (N_7588,N_7121,N_6884);
and U7589 (N_7589,N_7028,N_7471);
nand U7590 (N_7590,N_6971,N_7183);
xor U7591 (N_7591,N_7014,N_6850);
nand U7592 (N_7592,N_7056,N_7400);
or U7593 (N_7593,N_6836,N_7407);
nand U7594 (N_7594,N_7498,N_7381);
nor U7595 (N_7595,N_6859,N_7069);
or U7596 (N_7596,N_7355,N_7110);
xor U7597 (N_7597,N_7445,N_7470);
and U7598 (N_7598,N_6834,N_6784);
nand U7599 (N_7599,N_7220,N_6969);
nand U7600 (N_7600,N_7187,N_7346);
nand U7601 (N_7601,N_6854,N_7330);
xnor U7602 (N_7602,N_7186,N_7026);
or U7603 (N_7603,N_7265,N_7151);
nor U7604 (N_7604,N_7422,N_6875);
nand U7605 (N_7605,N_6908,N_7161);
xnor U7606 (N_7606,N_7276,N_6978);
xnor U7607 (N_7607,N_7067,N_6879);
nand U7608 (N_7608,N_7100,N_7132);
and U7609 (N_7609,N_7000,N_7489);
and U7610 (N_7610,N_7245,N_6931);
xor U7611 (N_7611,N_7401,N_7001);
nor U7612 (N_7612,N_7084,N_7019);
xor U7613 (N_7613,N_6809,N_7107);
and U7614 (N_7614,N_7173,N_7380);
and U7615 (N_7615,N_7299,N_6807);
and U7616 (N_7616,N_6842,N_7052);
and U7617 (N_7617,N_6973,N_7225);
and U7618 (N_7618,N_6870,N_7357);
nand U7619 (N_7619,N_7092,N_6833);
nand U7620 (N_7620,N_7334,N_7184);
xnor U7621 (N_7621,N_6902,N_6997);
nor U7622 (N_7622,N_6812,N_7426);
or U7623 (N_7623,N_6852,N_6981);
nor U7624 (N_7624,N_7441,N_7017);
xor U7625 (N_7625,N_7289,N_7244);
nand U7626 (N_7626,N_6869,N_7438);
xor U7627 (N_7627,N_6961,N_7212);
xnor U7628 (N_7628,N_6960,N_7246);
nor U7629 (N_7629,N_6946,N_6841);
xnor U7630 (N_7630,N_6754,N_7491);
or U7631 (N_7631,N_7300,N_7117);
or U7632 (N_7632,N_7496,N_7249);
nor U7633 (N_7633,N_6957,N_7448);
nand U7634 (N_7634,N_6761,N_7024);
or U7635 (N_7635,N_6787,N_7106);
nand U7636 (N_7636,N_7045,N_7352);
or U7637 (N_7637,N_7202,N_7162);
or U7638 (N_7638,N_7288,N_7284);
nor U7639 (N_7639,N_6853,N_6986);
nor U7640 (N_7640,N_6826,N_6979);
nand U7641 (N_7641,N_7462,N_7226);
nor U7642 (N_7642,N_7066,N_7485);
and U7643 (N_7643,N_6811,N_7022);
xor U7644 (N_7644,N_7287,N_7443);
nor U7645 (N_7645,N_7293,N_7379);
or U7646 (N_7646,N_6797,N_7283);
nand U7647 (N_7647,N_7171,N_7440);
nand U7648 (N_7648,N_7160,N_7262);
nand U7649 (N_7649,N_7169,N_7072);
or U7650 (N_7650,N_7112,N_6764);
xor U7651 (N_7651,N_7365,N_6765);
nor U7652 (N_7652,N_7133,N_7364);
and U7653 (N_7653,N_7123,N_6782);
or U7654 (N_7654,N_6947,N_7263);
xor U7655 (N_7655,N_6792,N_7412);
xor U7656 (N_7656,N_7354,N_6780);
nor U7657 (N_7657,N_7207,N_6880);
and U7658 (N_7658,N_7254,N_6923);
or U7659 (N_7659,N_6821,N_6938);
nand U7660 (N_7660,N_7370,N_7475);
or U7661 (N_7661,N_7053,N_7077);
or U7662 (N_7662,N_6993,N_7175);
nor U7663 (N_7663,N_7398,N_6994);
or U7664 (N_7664,N_7371,N_7197);
or U7665 (N_7665,N_7079,N_7232);
or U7666 (N_7666,N_6759,N_7406);
and U7667 (N_7667,N_6813,N_6825);
or U7668 (N_7668,N_6895,N_7335);
and U7669 (N_7669,N_7074,N_6962);
nor U7670 (N_7670,N_7153,N_6858);
nor U7671 (N_7671,N_7086,N_6755);
xnor U7672 (N_7672,N_7329,N_6832);
and U7673 (N_7673,N_7259,N_7034);
nor U7674 (N_7674,N_6983,N_7239);
or U7675 (N_7675,N_6776,N_6829);
and U7676 (N_7676,N_6881,N_7473);
and U7677 (N_7677,N_6885,N_7156);
nand U7678 (N_7678,N_7349,N_6892);
or U7679 (N_7679,N_7229,N_6955);
nor U7680 (N_7680,N_7405,N_7359);
or U7681 (N_7681,N_6909,N_7037);
nor U7682 (N_7682,N_7463,N_7224);
nor U7683 (N_7683,N_6802,N_6871);
nor U7684 (N_7684,N_7270,N_7433);
nand U7685 (N_7685,N_7097,N_7030);
and U7686 (N_7686,N_6779,N_7313);
nor U7687 (N_7687,N_6840,N_7057);
and U7688 (N_7688,N_7233,N_7430);
nor U7689 (N_7689,N_7458,N_7088);
nor U7690 (N_7690,N_7120,N_7176);
and U7691 (N_7691,N_7320,N_7499);
or U7692 (N_7692,N_7250,N_7091);
xnor U7693 (N_7693,N_7286,N_7073);
xnor U7694 (N_7694,N_7303,N_7126);
and U7695 (N_7695,N_7145,N_7331);
and U7696 (N_7696,N_7082,N_7198);
and U7697 (N_7697,N_6919,N_6935);
or U7698 (N_7698,N_7447,N_7495);
nor U7699 (N_7699,N_7345,N_6845);
or U7700 (N_7700,N_6904,N_6864);
nand U7701 (N_7701,N_7375,N_7437);
nor U7702 (N_7702,N_7435,N_7482);
or U7703 (N_7703,N_7309,N_7230);
xnor U7704 (N_7704,N_6877,N_6903);
or U7705 (N_7705,N_7149,N_6808);
xnor U7706 (N_7706,N_6975,N_7373);
xor U7707 (N_7707,N_7290,N_7418);
nor U7708 (N_7708,N_7025,N_6774);
or U7709 (N_7709,N_7115,N_7451);
xor U7710 (N_7710,N_7103,N_6862);
nor U7711 (N_7711,N_7339,N_7461);
xor U7712 (N_7712,N_6805,N_7188);
and U7713 (N_7713,N_7104,N_7050);
or U7714 (N_7714,N_7337,N_7146);
xor U7715 (N_7715,N_7087,N_6924);
and U7716 (N_7716,N_7165,N_7136);
and U7717 (N_7717,N_7140,N_7427);
nor U7718 (N_7718,N_6944,N_6873);
nor U7719 (N_7719,N_7033,N_6982);
nor U7720 (N_7720,N_7209,N_6999);
or U7721 (N_7721,N_6874,N_7341);
or U7722 (N_7722,N_7384,N_7377);
xor U7723 (N_7723,N_7312,N_7456);
or U7724 (N_7724,N_7179,N_7386);
nand U7725 (N_7725,N_7138,N_7046);
nand U7726 (N_7726,N_6932,N_6888);
nor U7727 (N_7727,N_6916,N_7166);
and U7728 (N_7728,N_7281,N_7148);
xnor U7729 (N_7729,N_7015,N_6819);
nand U7730 (N_7730,N_6988,N_7369);
nor U7731 (N_7731,N_7061,N_6896);
and U7732 (N_7732,N_7338,N_6933);
and U7733 (N_7733,N_6949,N_7089);
nor U7734 (N_7734,N_7062,N_7144);
or U7735 (N_7735,N_7382,N_7478);
and U7736 (N_7736,N_7206,N_7361);
or U7737 (N_7737,N_7472,N_7269);
xnor U7738 (N_7738,N_7051,N_6987);
nor U7739 (N_7739,N_6769,N_7154);
xnor U7740 (N_7740,N_7016,N_7237);
nor U7741 (N_7741,N_6803,N_7310);
and U7742 (N_7742,N_7348,N_7041);
or U7743 (N_7743,N_6856,N_7018);
and U7744 (N_7744,N_7446,N_7080);
nor U7745 (N_7745,N_7150,N_7457);
or U7746 (N_7746,N_7439,N_7271);
or U7747 (N_7747,N_7178,N_7043);
nand U7748 (N_7748,N_6912,N_6996);
or U7749 (N_7749,N_6899,N_7215);
nor U7750 (N_7750,N_6758,N_6936);
xnor U7751 (N_7751,N_7157,N_7356);
nand U7752 (N_7752,N_7049,N_7174);
nor U7753 (N_7753,N_7409,N_6775);
xnor U7754 (N_7754,N_7134,N_7469);
and U7755 (N_7755,N_7211,N_7429);
or U7756 (N_7756,N_6985,N_7419);
xnor U7757 (N_7757,N_7460,N_7009);
or U7758 (N_7758,N_7047,N_7416);
or U7759 (N_7759,N_7279,N_6752);
or U7760 (N_7760,N_6763,N_7251);
nand U7761 (N_7761,N_7214,N_7039);
xor U7762 (N_7762,N_7342,N_7415);
or U7763 (N_7763,N_6810,N_6984);
nor U7764 (N_7764,N_7116,N_7479);
or U7765 (N_7765,N_7322,N_6945);
or U7766 (N_7766,N_7213,N_6794);
nor U7767 (N_7767,N_6925,N_7340);
or U7768 (N_7768,N_7241,N_6929);
or U7769 (N_7769,N_7297,N_7125);
nor U7770 (N_7770,N_6788,N_6835);
nor U7771 (N_7771,N_7152,N_7261);
nor U7772 (N_7772,N_7203,N_6806);
and U7773 (N_7773,N_7076,N_7005);
or U7774 (N_7774,N_7459,N_6770);
or U7775 (N_7775,N_6959,N_6848);
xnor U7776 (N_7776,N_7408,N_7105);
nand U7777 (N_7777,N_7484,N_6900);
and U7778 (N_7778,N_7453,N_7021);
nor U7779 (N_7779,N_7351,N_7483);
or U7780 (N_7780,N_7247,N_6855);
and U7781 (N_7781,N_6766,N_7301);
nand U7782 (N_7782,N_7314,N_7332);
and U7783 (N_7783,N_7094,N_6798);
or U7784 (N_7784,N_6893,N_6867);
nand U7785 (N_7785,N_7007,N_7285);
nand U7786 (N_7786,N_6940,N_7032);
nor U7787 (N_7787,N_7182,N_6887);
or U7788 (N_7788,N_6839,N_7434);
and U7789 (N_7789,N_7060,N_6939);
and U7790 (N_7790,N_6998,N_6861);
xnor U7791 (N_7791,N_7199,N_6814);
nor U7792 (N_7792,N_7119,N_6822);
nor U7793 (N_7793,N_6950,N_7109);
xor U7794 (N_7794,N_7455,N_7044);
and U7795 (N_7795,N_7031,N_7494);
nor U7796 (N_7796,N_6786,N_7177);
and U7797 (N_7797,N_7081,N_7090);
or U7798 (N_7798,N_6920,N_7316);
or U7799 (N_7799,N_7048,N_7449);
and U7800 (N_7800,N_7328,N_7163);
and U7801 (N_7801,N_6828,N_7099);
and U7802 (N_7802,N_7167,N_7294);
nand U7803 (N_7803,N_7098,N_7344);
or U7804 (N_7804,N_7023,N_7227);
and U7805 (N_7805,N_7323,N_7307);
and U7806 (N_7806,N_7292,N_7372);
and U7807 (N_7807,N_7141,N_6934);
xnor U7808 (N_7808,N_7219,N_7436);
and U7809 (N_7809,N_7390,N_7142);
nor U7810 (N_7810,N_7305,N_7143);
or U7811 (N_7811,N_6948,N_6992);
xor U7812 (N_7812,N_7315,N_7476);
nor U7813 (N_7813,N_7387,N_6753);
nor U7814 (N_7814,N_7210,N_6963);
and U7815 (N_7815,N_7353,N_6926);
or U7816 (N_7816,N_6942,N_6922);
or U7817 (N_7817,N_6799,N_6823);
nand U7818 (N_7818,N_7302,N_6928);
and U7819 (N_7819,N_7266,N_7071);
and U7820 (N_7820,N_6768,N_7423);
or U7821 (N_7821,N_6927,N_7391);
nor U7822 (N_7822,N_7236,N_6783);
nor U7823 (N_7823,N_7376,N_7327);
or U7824 (N_7824,N_7243,N_7374);
xnor U7825 (N_7825,N_6849,N_7394);
or U7826 (N_7826,N_7278,N_6876);
and U7827 (N_7827,N_7159,N_7333);
and U7828 (N_7828,N_7324,N_7195);
nand U7829 (N_7829,N_6921,N_7190);
xnor U7830 (N_7830,N_7114,N_7304);
or U7831 (N_7831,N_7410,N_7466);
xor U7832 (N_7832,N_7366,N_7268);
and U7833 (N_7833,N_7040,N_6991);
and U7834 (N_7834,N_7424,N_6750);
nand U7835 (N_7835,N_7252,N_7078);
nor U7836 (N_7836,N_7218,N_6762);
xor U7837 (N_7837,N_7200,N_7467);
or U7838 (N_7838,N_7193,N_6818);
nor U7839 (N_7839,N_6844,N_7397);
nand U7840 (N_7840,N_7481,N_7011);
nand U7841 (N_7841,N_7147,N_6941);
nor U7842 (N_7842,N_6889,N_7325);
nand U7843 (N_7843,N_7194,N_6831);
and U7844 (N_7844,N_7296,N_6914);
nand U7845 (N_7845,N_7428,N_7360);
nor U7846 (N_7846,N_7065,N_7421);
or U7847 (N_7847,N_7205,N_7363);
xor U7848 (N_7848,N_7280,N_7477);
and U7849 (N_7849,N_7411,N_7004);
nand U7850 (N_7850,N_7282,N_7260);
or U7851 (N_7851,N_7396,N_6872);
and U7852 (N_7852,N_7417,N_7319);
or U7853 (N_7853,N_7108,N_7277);
nor U7854 (N_7854,N_7042,N_6882);
nand U7855 (N_7855,N_7450,N_6843);
nand U7856 (N_7856,N_6796,N_7393);
and U7857 (N_7857,N_7035,N_7368);
and U7858 (N_7858,N_6989,N_6954);
and U7859 (N_7859,N_7336,N_7273);
and U7860 (N_7860,N_7216,N_7431);
and U7861 (N_7861,N_6966,N_6778);
nand U7862 (N_7862,N_7404,N_6865);
and U7863 (N_7863,N_6846,N_7137);
or U7864 (N_7864,N_6824,N_7464);
or U7865 (N_7865,N_7096,N_7027);
nor U7866 (N_7866,N_7274,N_7311);
and U7867 (N_7867,N_6898,N_6897);
or U7868 (N_7868,N_7403,N_6791);
or U7869 (N_7869,N_7248,N_7242);
nand U7870 (N_7870,N_7234,N_7291);
and U7871 (N_7871,N_6772,N_7059);
and U7872 (N_7872,N_7264,N_7128);
and U7873 (N_7873,N_7468,N_6907);
and U7874 (N_7874,N_7010,N_6757);
xnor U7875 (N_7875,N_7336,N_7313);
nand U7876 (N_7876,N_7196,N_6860);
or U7877 (N_7877,N_7037,N_7015);
and U7878 (N_7878,N_7291,N_6912);
and U7879 (N_7879,N_7396,N_7096);
nand U7880 (N_7880,N_6888,N_7206);
or U7881 (N_7881,N_7495,N_7099);
or U7882 (N_7882,N_6941,N_7419);
nor U7883 (N_7883,N_6965,N_6932);
xor U7884 (N_7884,N_7258,N_7195);
nor U7885 (N_7885,N_6983,N_7336);
or U7886 (N_7886,N_7443,N_7363);
xor U7887 (N_7887,N_7014,N_6816);
nand U7888 (N_7888,N_7396,N_6917);
or U7889 (N_7889,N_7384,N_6812);
xnor U7890 (N_7890,N_7136,N_7064);
nor U7891 (N_7891,N_7322,N_7069);
or U7892 (N_7892,N_7141,N_7358);
and U7893 (N_7893,N_7385,N_7348);
and U7894 (N_7894,N_7478,N_7385);
nor U7895 (N_7895,N_7113,N_7022);
xor U7896 (N_7896,N_6952,N_7483);
nand U7897 (N_7897,N_7255,N_6781);
xnor U7898 (N_7898,N_7099,N_7025);
xnor U7899 (N_7899,N_6755,N_6784);
xnor U7900 (N_7900,N_7014,N_7475);
nand U7901 (N_7901,N_7121,N_6800);
nand U7902 (N_7902,N_7414,N_7213);
xor U7903 (N_7903,N_6803,N_7026);
and U7904 (N_7904,N_7267,N_7030);
xnor U7905 (N_7905,N_7390,N_7018);
nor U7906 (N_7906,N_7211,N_7389);
nor U7907 (N_7907,N_7380,N_7120);
nand U7908 (N_7908,N_6845,N_6967);
nor U7909 (N_7909,N_6939,N_7498);
xnor U7910 (N_7910,N_7023,N_7196);
and U7911 (N_7911,N_7186,N_7496);
xnor U7912 (N_7912,N_6948,N_6857);
and U7913 (N_7913,N_7448,N_6924);
or U7914 (N_7914,N_7270,N_6896);
and U7915 (N_7915,N_6968,N_7160);
xnor U7916 (N_7916,N_7186,N_6935);
nand U7917 (N_7917,N_7033,N_7368);
or U7918 (N_7918,N_6764,N_7339);
and U7919 (N_7919,N_6912,N_6809);
or U7920 (N_7920,N_7076,N_7329);
nand U7921 (N_7921,N_6766,N_7497);
nor U7922 (N_7922,N_6963,N_7396);
or U7923 (N_7923,N_7125,N_7256);
and U7924 (N_7924,N_7255,N_7147);
nor U7925 (N_7925,N_7337,N_7031);
and U7926 (N_7926,N_7293,N_7029);
xnor U7927 (N_7927,N_7074,N_7110);
nand U7928 (N_7928,N_6828,N_7199);
or U7929 (N_7929,N_6873,N_7487);
nand U7930 (N_7930,N_6752,N_7381);
nor U7931 (N_7931,N_7034,N_7262);
nand U7932 (N_7932,N_7212,N_6901);
nor U7933 (N_7933,N_6888,N_6793);
nand U7934 (N_7934,N_6881,N_6813);
xor U7935 (N_7935,N_7097,N_7351);
nand U7936 (N_7936,N_7322,N_7113);
xnor U7937 (N_7937,N_6762,N_7131);
or U7938 (N_7938,N_7368,N_6770);
nor U7939 (N_7939,N_7093,N_7347);
xnor U7940 (N_7940,N_7190,N_6815);
or U7941 (N_7941,N_7294,N_7315);
and U7942 (N_7942,N_6824,N_7123);
xor U7943 (N_7943,N_7265,N_7146);
or U7944 (N_7944,N_7202,N_7242);
nand U7945 (N_7945,N_6920,N_7200);
or U7946 (N_7946,N_7006,N_7133);
nor U7947 (N_7947,N_7331,N_7015);
xnor U7948 (N_7948,N_6929,N_7096);
nand U7949 (N_7949,N_7284,N_6771);
and U7950 (N_7950,N_6953,N_7394);
xnor U7951 (N_7951,N_6963,N_7112);
or U7952 (N_7952,N_7192,N_6844);
xnor U7953 (N_7953,N_6963,N_6854);
nand U7954 (N_7954,N_7125,N_7014);
xnor U7955 (N_7955,N_6772,N_7041);
or U7956 (N_7956,N_6801,N_6862);
nand U7957 (N_7957,N_7317,N_6816);
and U7958 (N_7958,N_7459,N_7244);
xor U7959 (N_7959,N_7319,N_6907);
xor U7960 (N_7960,N_7082,N_7409);
or U7961 (N_7961,N_7485,N_7018);
nand U7962 (N_7962,N_6828,N_7433);
and U7963 (N_7963,N_7094,N_6769);
and U7964 (N_7964,N_6793,N_7329);
nand U7965 (N_7965,N_7366,N_7383);
nand U7966 (N_7966,N_7057,N_7338);
xnor U7967 (N_7967,N_7116,N_6920);
xnor U7968 (N_7968,N_7040,N_7422);
nor U7969 (N_7969,N_6853,N_7018);
xnor U7970 (N_7970,N_7117,N_6833);
nand U7971 (N_7971,N_7330,N_6905);
xor U7972 (N_7972,N_6753,N_6986);
nor U7973 (N_7973,N_6970,N_7024);
nor U7974 (N_7974,N_7068,N_7373);
nand U7975 (N_7975,N_6867,N_7438);
xnor U7976 (N_7976,N_6797,N_7057);
and U7977 (N_7977,N_7047,N_6992);
and U7978 (N_7978,N_7343,N_6856);
nor U7979 (N_7979,N_6911,N_7242);
nand U7980 (N_7980,N_7221,N_6767);
and U7981 (N_7981,N_7093,N_6806);
nand U7982 (N_7982,N_6956,N_6760);
and U7983 (N_7983,N_7149,N_7239);
nor U7984 (N_7984,N_7427,N_7375);
and U7985 (N_7985,N_6968,N_7471);
nor U7986 (N_7986,N_7175,N_7461);
nand U7987 (N_7987,N_6878,N_6995);
or U7988 (N_7988,N_7141,N_7250);
xor U7989 (N_7989,N_6892,N_7499);
nor U7990 (N_7990,N_6887,N_7410);
nor U7991 (N_7991,N_6903,N_7445);
nor U7992 (N_7992,N_6893,N_6821);
nor U7993 (N_7993,N_6774,N_6851);
xnor U7994 (N_7994,N_7262,N_7473);
or U7995 (N_7995,N_6885,N_6839);
xor U7996 (N_7996,N_6951,N_7204);
xnor U7997 (N_7997,N_7259,N_7102);
or U7998 (N_7998,N_6827,N_6932);
and U7999 (N_7999,N_7146,N_7250);
nand U8000 (N_8000,N_7404,N_7067);
nor U8001 (N_8001,N_7227,N_6922);
nor U8002 (N_8002,N_7029,N_6825);
nand U8003 (N_8003,N_7291,N_6893);
nand U8004 (N_8004,N_7497,N_6898);
or U8005 (N_8005,N_7391,N_7254);
nand U8006 (N_8006,N_7431,N_7204);
xor U8007 (N_8007,N_6951,N_6944);
nand U8008 (N_8008,N_6782,N_6774);
and U8009 (N_8009,N_7286,N_6984);
nor U8010 (N_8010,N_7441,N_6893);
nor U8011 (N_8011,N_6840,N_6751);
nand U8012 (N_8012,N_7155,N_7146);
xor U8013 (N_8013,N_7148,N_7046);
nand U8014 (N_8014,N_7441,N_7178);
or U8015 (N_8015,N_7248,N_6978);
nand U8016 (N_8016,N_7370,N_7489);
xnor U8017 (N_8017,N_7076,N_7169);
nor U8018 (N_8018,N_6898,N_7238);
nand U8019 (N_8019,N_7485,N_6767);
nor U8020 (N_8020,N_7081,N_7386);
or U8021 (N_8021,N_7328,N_7420);
and U8022 (N_8022,N_6791,N_7190);
nor U8023 (N_8023,N_7483,N_7190);
xnor U8024 (N_8024,N_6865,N_7159);
nand U8025 (N_8025,N_6992,N_7182);
or U8026 (N_8026,N_7278,N_7396);
xnor U8027 (N_8027,N_7167,N_6803);
or U8028 (N_8028,N_7193,N_7415);
nor U8029 (N_8029,N_6855,N_6908);
nor U8030 (N_8030,N_6870,N_6941);
and U8031 (N_8031,N_6976,N_6758);
nand U8032 (N_8032,N_7299,N_7298);
or U8033 (N_8033,N_7202,N_7203);
xnor U8034 (N_8034,N_7384,N_7144);
and U8035 (N_8035,N_7452,N_7346);
nor U8036 (N_8036,N_6773,N_7388);
and U8037 (N_8037,N_7305,N_7114);
nor U8038 (N_8038,N_7461,N_7118);
nor U8039 (N_8039,N_7213,N_7391);
or U8040 (N_8040,N_6931,N_7333);
and U8041 (N_8041,N_7210,N_7376);
and U8042 (N_8042,N_7209,N_6770);
and U8043 (N_8043,N_6876,N_7051);
nor U8044 (N_8044,N_7109,N_7017);
or U8045 (N_8045,N_7477,N_6901);
or U8046 (N_8046,N_6841,N_7100);
xnor U8047 (N_8047,N_7385,N_7263);
nor U8048 (N_8048,N_7195,N_7264);
nor U8049 (N_8049,N_7053,N_7262);
nor U8050 (N_8050,N_7161,N_7235);
nand U8051 (N_8051,N_6967,N_6835);
or U8052 (N_8052,N_7067,N_6979);
nor U8053 (N_8053,N_7067,N_6792);
nand U8054 (N_8054,N_7270,N_6836);
or U8055 (N_8055,N_7236,N_7142);
xnor U8056 (N_8056,N_6982,N_7278);
or U8057 (N_8057,N_6990,N_7361);
and U8058 (N_8058,N_6863,N_6949);
nor U8059 (N_8059,N_7125,N_6868);
nor U8060 (N_8060,N_7241,N_7202);
nand U8061 (N_8061,N_7470,N_7491);
xor U8062 (N_8062,N_7032,N_7441);
xnor U8063 (N_8063,N_7431,N_7268);
and U8064 (N_8064,N_6793,N_6883);
or U8065 (N_8065,N_7477,N_7225);
xnor U8066 (N_8066,N_7304,N_6827);
and U8067 (N_8067,N_6878,N_6855);
nor U8068 (N_8068,N_7019,N_7416);
nor U8069 (N_8069,N_7340,N_7217);
nand U8070 (N_8070,N_6777,N_7244);
nor U8071 (N_8071,N_7375,N_7324);
nand U8072 (N_8072,N_6932,N_6901);
xor U8073 (N_8073,N_7388,N_7391);
xnor U8074 (N_8074,N_7077,N_6803);
nor U8075 (N_8075,N_7184,N_7431);
nor U8076 (N_8076,N_6888,N_7188);
nor U8077 (N_8077,N_7201,N_6833);
and U8078 (N_8078,N_6996,N_7351);
and U8079 (N_8079,N_7290,N_6907);
or U8080 (N_8080,N_6795,N_6779);
xnor U8081 (N_8081,N_7081,N_7476);
nand U8082 (N_8082,N_7027,N_7397);
and U8083 (N_8083,N_7231,N_6847);
or U8084 (N_8084,N_7448,N_7265);
nor U8085 (N_8085,N_7059,N_7498);
nand U8086 (N_8086,N_7196,N_7247);
xor U8087 (N_8087,N_7467,N_7217);
and U8088 (N_8088,N_6784,N_7063);
or U8089 (N_8089,N_7300,N_6975);
nor U8090 (N_8090,N_7339,N_7382);
or U8091 (N_8091,N_6751,N_6821);
nand U8092 (N_8092,N_6818,N_7412);
nor U8093 (N_8093,N_7190,N_7160);
or U8094 (N_8094,N_7006,N_7069);
nor U8095 (N_8095,N_7128,N_6770);
xnor U8096 (N_8096,N_7049,N_6871);
or U8097 (N_8097,N_6909,N_7486);
nand U8098 (N_8098,N_7002,N_7280);
and U8099 (N_8099,N_7160,N_7373);
xor U8100 (N_8100,N_7466,N_6920);
and U8101 (N_8101,N_6986,N_6887);
and U8102 (N_8102,N_7334,N_7228);
and U8103 (N_8103,N_7412,N_7380);
nor U8104 (N_8104,N_6904,N_7191);
nor U8105 (N_8105,N_6859,N_6784);
or U8106 (N_8106,N_6905,N_7454);
and U8107 (N_8107,N_6900,N_6970);
xnor U8108 (N_8108,N_7093,N_7062);
and U8109 (N_8109,N_6944,N_7226);
and U8110 (N_8110,N_6995,N_6870);
xnor U8111 (N_8111,N_7164,N_7389);
or U8112 (N_8112,N_7202,N_6807);
xor U8113 (N_8113,N_7462,N_7277);
xnor U8114 (N_8114,N_6869,N_7305);
or U8115 (N_8115,N_7130,N_6910);
nor U8116 (N_8116,N_7498,N_7137);
xnor U8117 (N_8117,N_7342,N_7203);
or U8118 (N_8118,N_6811,N_7448);
or U8119 (N_8119,N_7420,N_7168);
and U8120 (N_8120,N_6952,N_6992);
nor U8121 (N_8121,N_6872,N_6848);
and U8122 (N_8122,N_7468,N_6997);
and U8123 (N_8123,N_7252,N_6944);
or U8124 (N_8124,N_6869,N_7153);
nor U8125 (N_8125,N_6812,N_7080);
nand U8126 (N_8126,N_7472,N_7140);
nor U8127 (N_8127,N_7315,N_7140);
nand U8128 (N_8128,N_7060,N_7424);
nand U8129 (N_8129,N_7117,N_6764);
nand U8130 (N_8130,N_6869,N_7297);
xnor U8131 (N_8131,N_7482,N_7260);
and U8132 (N_8132,N_7272,N_7205);
or U8133 (N_8133,N_7199,N_7197);
nor U8134 (N_8134,N_7393,N_7442);
nor U8135 (N_8135,N_7318,N_7203);
nand U8136 (N_8136,N_7428,N_6777);
xor U8137 (N_8137,N_7197,N_6793);
nor U8138 (N_8138,N_7399,N_7329);
nor U8139 (N_8139,N_7156,N_7307);
or U8140 (N_8140,N_7451,N_7311);
or U8141 (N_8141,N_6933,N_6878);
nor U8142 (N_8142,N_7398,N_6925);
nand U8143 (N_8143,N_6761,N_7337);
xnor U8144 (N_8144,N_7058,N_7432);
xnor U8145 (N_8145,N_6761,N_7328);
nor U8146 (N_8146,N_7133,N_7042);
or U8147 (N_8147,N_7046,N_7406);
nand U8148 (N_8148,N_7288,N_7124);
or U8149 (N_8149,N_7073,N_7110);
nor U8150 (N_8150,N_7408,N_7417);
nor U8151 (N_8151,N_7186,N_7309);
nor U8152 (N_8152,N_6887,N_7067);
nor U8153 (N_8153,N_6963,N_6829);
and U8154 (N_8154,N_6997,N_7349);
and U8155 (N_8155,N_6873,N_7171);
nor U8156 (N_8156,N_7229,N_7312);
nand U8157 (N_8157,N_7372,N_6876);
and U8158 (N_8158,N_6977,N_6879);
nor U8159 (N_8159,N_7326,N_7021);
nor U8160 (N_8160,N_7362,N_7184);
nand U8161 (N_8161,N_7481,N_7132);
xor U8162 (N_8162,N_6805,N_6843);
xor U8163 (N_8163,N_6943,N_7180);
nor U8164 (N_8164,N_7240,N_6964);
or U8165 (N_8165,N_7417,N_7172);
nor U8166 (N_8166,N_7286,N_7000);
nand U8167 (N_8167,N_7211,N_6953);
or U8168 (N_8168,N_7323,N_6876);
nor U8169 (N_8169,N_6890,N_6986);
and U8170 (N_8170,N_7235,N_7312);
nor U8171 (N_8171,N_7236,N_7011);
nand U8172 (N_8172,N_7174,N_7173);
nand U8173 (N_8173,N_7312,N_7031);
nand U8174 (N_8174,N_6785,N_6995);
xor U8175 (N_8175,N_7281,N_7339);
and U8176 (N_8176,N_6919,N_7452);
or U8177 (N_8177,N_7358,N_6769);
or U8178 (N_8178,N_7192,N_6833);
xnor U8179 (N_8179,N_7282,N_7210);
nor U8180 (N_8180,N_6914,N_6929);
nand U8181 (N_8181,N_7346,N_6916);
xnor U8182 (N_8182,N_7277,N_7404);
nor U8183 (N_8183,N_6896,N_6923);
or U8184 (N_8184,N_7238,N_6845);
nand U8185 (N_8185,N_6825,N_6757);
nor U8186 (N_8186,N_7494,N_7467);
and U8187 (N_8187,N_7432,N_6797);
and U8188 (N_8188,N_7418,N_7197);
xnor U8189 (N_8189,N_6925,N_7438);
nand U8190 (N_8190,N_6881,N_7312);
nor U8191 (N_8191,N_7011,N_7048);
or U8192 (N_8192,N_7346,N_6892);
xnor U8193 (N_8193,N_6899,N_7136);
and U8194 (N_8194,N_7331,N_7226);
nand U8195 (N_8195,N_7007,N_7348);
nand U8196 (N_8196,N_6883,N_6869);
nor U8197 (N_8197,N_7318,N_7387);
xnor U8198 (N_8198,N_7372,N_6972);
or U8199 (N_8199,N_6755,N_7232);
xor U8200 (N_8200,N_7170,N_7264);
nand U8201 (N_8201,N_7097,N_7416);
or U8202 (N_8202,N_7022,N_6806);
nand U8203 (N_8203,N_7041,N_7390);
nor U8204 (N_8204,N_7303,N_6957);
nand U8205 (N_8205,N_6810,N_7238);
xor U8206 (N_8206,N_7361,N_7121);
or U8207 (N_8207,N_7269,N_6934);
xor U8208 (N_8208,N_7148,N_7487);
and U8209 (N_8209,N_7295,N_6874);
nand U8210 (N_8210,N_6837,N_7380);
nor U8211 (N_8211,N_7396,N_7073);
and U8212 (N_8212,N_7277,N_6751);
or U8213 (N_8213,N_7475,N_6877);
nor U8214 (N_8214,N_6974,N_6949);
nor U8215 (N_8215,N_7380,N_6969);
nand U8216 (N_8216,N_7452,N_7286);
xnor U8217 (N_8217,N_7182,N_6888);
xnor U8218 (N_8218,N_7327,N_6800);
and U8219 (N_8219,N_7316,N_7391);
or U8220 (N_8220,N_7194,N_7460);
nand U8221 (N_8221,N_7224,N_6850);
and U8222 (N_8222,N_6839,N_6761);
xnor U8223 (N_8223,N_6940,N_7076);
or U8224 (N_8224,N_7423,N_6773);
nand U8225 (N_8225,N_7140,N_7062);
and U8226 (N_8226,N_7057,N_7418);
nand U8227 (N_8227,N_6782,N_7121);
xor U8228 (N_8228,N_7458,N_6858);
nand U8229 (N_8229,N_7308,N_7316);
nor U8230 (N_8230,N_7320,N_7178);
xor U8231 (N_8231,N_7256,N_7200);
xor U8232 (N_8232,N_7392,N_6942);
xnor U8233 (N_8233,N_6918,N_7226);
nand U8234 (N_8234,N_7253,N_7481);
and U8235 (N_8235,N_7358,N_7053);
xnor U8236 (N_8236,N_7178,N_7050);
or U8237 (N_8237,N_6959,N_7130);
nand U8238 (N_8238,N_7484,N_6961);
and U8239 (N_8239,N_6835,N_7043);
or U8240 (N_8240,N_7255,N_6989);
nand U8241 (N_8241,N_7440,N_7373);
nor U8242 (N_8242,N_7015,N_7252);
nand U8243 (N_8243,N_7361,N_6793);
xor U8244 (N_8244,N_6901,N_6918);
nand U8245 (N_8245,N_7313,N_7402);
nor U8246 (N_8246,N_7245,N_7315);
xnor U8247 (N_8247,N_7273,N_7223);
or U8248 (N_8248,N_6826,N_6949);
and U8249 (N_8249,N_7205,N_6854);
nor U8250 (N_8250,N_8149,N_7837);
and U8251 (N_8251,N_7519,N_8191);
xor U8252 (N_8252,N_7642,N_7629);
xnor U8253 (N_8253,N_7862,N_7786);
or U8254 (N_8254,N_7823,N_7876);
xor U8255 (N_8255,N_7684,N_7576);
xnor U8256 (N_8256,N_7963,N_7880);
nand U8257 (N_8257,N_7841,N_7778);
and U8258 (N_8258,N_8181,N_7831);
nand U8259 (N_8259,N_7705,N_8169);
nor U8260 (N_8260,N_8027,N_8141);
and U8261 (N_8261,N_8050,N_7545);
nand U8262 (N_8262,N_7985,N_7975);
nor U8263 (N_8263,N_8016,N_7733);
and U8264 (N_8264,N_7503,N_7991);
or U8265 (N_8265,N_7795,N_7799);
nand U8266 (N_8266,N_7518,N_7577);
and U8267 (N_8267,N_8119,N_7660);
or U8268 (N_8268,N_8020,N_8182);
nand U8269 (N_8269,N_7744,N_8045);
or U8270 (N_8270,N_8057,N_8185);
or U8271 (N_8271,N_7633,N_7704);
and U8272 (N_8272,N_8039,N_7555);
nand U8273 (N_8273,N_8052,N_7513);
or U8274 (N_8274,N_7996,N_7520);
or U8275 (N_8275,N_8116,N_7643);
and U8276 (N_8276,N_8161,N_8097);
nor U8277 (N_8277,N_8004,N_7878);
nor U8278 (N_8278,N_7726,N_7822);
or U8279 (N_8279,N_8222,N_7649);
nand U8280 (N_8280,N_8217,N_7716);
xnor U8281 (N_8281,N_7804,N_8196);
xor U8282 (N_8282,N_7916,N_8211);
nor U8283 (N_8283,N_7685,N_7839);
nor U8284 (N_8284,N_7801,N_8018);
xor U8285 (N_8285,N_7510,N_7937);
nand U8286 (N_8286,N_7912,N_7508);
nor U8287 (N_8287,N_8112,N_8208);
nand U8288 (N_8288,N_8021,N_7693);
or U8289 (N_8289,N_7534,N_7748);
and U8290 (N_8290,N_8105,N_7775);
or U8291 (N_8291,N_7770,N_8127);
and U8292 (N_8292,N_7547,N_8066);
xnor U8293 (N_8293,N_7857,N_7600);
or U8294 (N_8294,N_8079,N_8044);
nor U8295 (N_8295,N_8240,N_7608);
xnor U8296 (N_8296,N_8114,N_7853);
or U8297 (N_8297,N_8213,N_7917);
xor U8298 (N_8298,N_7583,N_8029);
xor U8299 (N_8299,N_7724,N_7535);
or U8300 (N_8300,N_8201,N_7615);
xnor U8301 (N_8301,N_7550,N_7815);
or U8302 (N_8302,N_8022,N_8062);
and U8303 (N_8303,N_7502,N_7667);
or U8304 (N_8304,N_7607,N_7955);
xnor U8305 (N_8305,N_7983,N_8015);
or U8306 (N_8306,N_8153,N_7552);
xor U8307 (N_8307,N_7883,N_7563);
nor U8308 (N_8308,N_7903,N_7720);
and U8309 (N_8309,N_7929,N_7570);
xor U8310 (N_8310,N_8071,N_8162);
and U8311 (N_8311,N_7790,N_7905);
and U8312 (N_8312,N_7665,N_7617);
or U8313 (N_8313,N_7678,N_7889);
nor U8314 (N_8314,N_7741,N_8233);
nor U8315 (N_8315,N_7793,N_7967);
and U8316 (N_8316,N_7509,N_8229);
or U8317 (N_8317,N_8049,N_7962);
and U8318 (N_8318,N_8134,N_8058);
nor U8319 (N_8319,N_7779,N_7925);
nand U8320 (N_8320,N_8001,N_7868);
or U8321 (N_8321,N_7578,N_7906);
or U8322 (N_8322,N_8085,N_7700);
nor U8323 (N_8323,N_8108,N_7637);
nand U8324 (N_8324,N_8171,N_7900);
nand U8325 (N_8325,N_8013,N_8140);
xor U8326 (N_8326,N_7528,N_7611);
nand U8327 (N_8327,N_7689,N_7899);
nor U8328 (N_8328,N_7663,N_8006);
nor U8329 (N_8329,N_7904,N_7543);
nor U8330 (N_8330,N_7956,N_8040);
and U8331 (N_8331,N_8073,N_7585);
nand U8332 (N_8332,N_7625,N_8231);
or U8333 (N_8333,N_8170,N_8129);
nor U8334 (N_8334,N_7834,N_7910);
and U8335 (N_8335,N_7859,N_7881);
nand U8336 (N_8336,N_7957,N_7673);
and U8337 (N_8337,N_7527,N_7877);
nor U8338 (N_8338,N_7734,N_8163);
and U8339 (N_8339,N_8106,N_8035);
nand U8340 (N_8340,N_7674,N_8008);
xor U8341 (N_8341,N_7610,N_7539);
nor U8342 (N_8342,N_7742,N_7768);
xnor U8343 (N_8343,N_7845,N_7976);
xor U8344 (N_8344,N_8028,N_7544);
xnor U8345 (N_8345,N_8246,N_7747);
nand U8346 (N_8346,N_7875,N_8056);
or U8347 (N_8347,N_7767,N_8175);
or U8348 (N_8348,N_8184,N_7556);
xor U8349 (N_8349,N_7788,N_7909);
xnor U8350 (N_8350,N_7927,N_7773);
nand U8351 (N_8351,N_7864,N_8000);
nand U8352 (N_8352,N_7749,N_7719);
nor U8353 (N_8353,N_7698,N_7706);
nand U8354 (N_8354,N_7567,N_8226);
xnor U8355 (N_8355,N_7970,N_8143);
and U8356 (N_8356,N_7536,N_7952);
nand U8357 (N_8357,N_7800,N_8032);
nor U8358 (N_8358,N_7626,N_7943);
nand U8359 (N_8359,N_7817,N_7592);
xor U8360 (N_8360,N_8077,N_7670);
and U8361 (N_8361,N_7558,N_7683);
and U8362 (N_8362,N_7731,N_7870);
or U8363 (N_8363,N_7701,N_8033);
nand U8364 (N_8364,N_7695,N_8247);
nor U8365 (N_8365,N_7762,N_7710);
or U8366 (N_8366,N_7727,N_8099);
and U8367 (N_8367,N_7814,N_7761);
nand U8368 (N_8368,N_7968,N_7812);
nor U8369 (N_8369,N_8068,N_7833);
nor U8370 (N_8370,N_8051,N_7691);
or U8371 (N_8371,N_7500,N_7818);
nor U8372 (N_8372,N_8160,N_8053);
xnor U8373 (N_8373,N_8124,N_7995);
and U8374 (N_8374,N_7715,N_7802);
xor U8375 (N_8375,N_8227,N_8224);
nor U8376 (N_8376,N_8003,N_7998);
xnor U8377 (N_8377,N_8121,N_8123);
xor U8378 (N_8378,N_7789,N_8195);
and U8379 (N_8379,N_7714,N_8002);
nor U8380 (N_8380,N_7803,N_7753);
xor U8381 (N_8381,N_7908,N_7791);
nand U8382 (N_8382,N_8054,N_7581);
xnor U8383 (N_8383,N_7948,N_7918);
or U8384 (N_8384,N_7627,N_7921);
nand U8385 (N_8385,N_8237,N_8120);
and U8386 (N_8386,N_7553,N_7892);
nand U8387 (N_8387,N_7882,N_7939);
nor U8388 (N_8388,N_8094,N_7897);
nor U8389 (N_8389,N_7588,N_7901);
xnor U8390 (N_8390,N_7688,N_8088);
or U8391 (N_8391,N_7835,N_7754);
or U8392 (N_8392,N_7636,N_8210);
xor U8393 (N_8393,N_8212,N_7532);
or U8394 (N_8394,N_8133,N_8074);
and U8395 (N_8395,N_7584,N_7538);
nor U8396 (N_8396,N_7923,N_7632);
nand U8397 (N_8397,N_8135,N_8194);
or U8398 (N_8398,N_8243,N_7507);
and U8399 (N_8399,N_7737,N_7711);
xor U8400 (N_8400,N_7751,N_8207);
xnor U8401 (N_8401,N_7650,N_7755);
nand U8402 (N_8402,N_7736,N_7809);
nor U8403 (N_8403,N_8087,N_7554);
xnor U8404 (N_8404,N_8216,N_7646);
and U8405 (N_8405,N_7568,N_8014);
xnor U8406 (N_8406,N_7512,N_7722);
nor U8407 (N_8407,N_7590,N_7657);
nand U8408 (N_8408,N_7707,N_7992);
nand U8409 (N_8409,N_7846,N_7517);
nor U8410 (N_8410,N_7565,N_8089);
xnor U8411 (N_8411,N_7514,N_7913);
and U8412 (N_8412,N_7863,N_7758);
and U8413 (N_8413,N_8091,N_7609);
xor U8414 (N_8414,N_7990,N_7529);
xnor U8415 (N_8415,N_7915,N_7690);
and U8416 (N_8416,N_7603,N_7622);
nor U8417 (N_8417,N_7630,N_7907);
and U8418 (N_8418,N_7564,N_7887);
and U8419 (N_8419,N_8158,N_7573);
and U8420 (N_8420,N_7652,N_8046);
or U8421 (N_8421,N_7838,N_7946);
or U8422 (N_8422,N_7858,N_8197);
xnor U8423 (N_8423,N_8131,N_8178);
nand U8424 (N_8424,N_7890,N_7951);
and U8425 (N_8425,N_7807,N_8125);
nand U8426 (N_8426,N_8138,N_7679);
xnor U8427 (N_8427,N_7774,N_7559);
xnor U8428 (N_8428,N_7624,N_7813);
nand U8429 (N_8429,N_8036,N_7826);
xnor U8430 (N_8430,N_7505,N_7666);
nand U8431 (N_8431,N_7548,N_8236);
or U8432 (N_8432,N_7856,N_7647);
xnor U8433 (N_8433,N_7816,N_7993);
or U8434 (N_8434,N_7732,N_7628);
or U8435 (N_8435,N_7787,N_8188);
and U8436 (N_8436,N_8193,N_7885);
xnor U8437 (N_8437,N_7501,N_8220);
nor U8438 (N_8438,N_7954,N_7780);
and U8439 (N_8439,N_7523,N_7965);
xor U8440 (N_8440,N_7551,N_7797);
nand U8441 (N_8441,N_7926,N_7709);
nand U8442 (N_8442,N_7728,N_7824);
xor U8443 (N_8443,N_7852,N_7825);
nand U8444 (N_8444,N_8168,N_7641);
xor U8445 (N_8445,N_8147,N_7855);
and U8446 (N_8446,N_7860,N_7723);
and U8447 (N_8447,N_7572,N_7756);
nor U8448 (N_8448,N_7596,N_7966);
or U8449 (N_8449,N_8031,N_7785);
xor U8450 (N_8450,N_8144,N_8078);
xnor U8451 (N_8451,N_7886,N_7934);
nand U8452 (N_8452,N_7949,N_7871);
nand U8453 (N_8453,N_8174,N_7595);
nor U8454 (N_8454,N_7696,N_7606);
nand U8455 (N_8455,N_7664,N_8048);
or U8456 (N_8456,N_7594,N_7618);
nand U8457 (N_8457,N_7542,N_8239);
and U8458 (N_8458,N_8249,N_7644);
nor U8459 (N_8459,N_8214,N_8146);
or U8460 (N_8460,N_7953,N_7869);
nand U8461 (N_8461,N_8081,N_8159);
or U8462 (N_8462,N_8202,N_8061);
nor U8463 (N_8463,N_7729,N_8083);
xnor U8464 (N_8464,N_7989,N_7879);
or U8465 (N_8465,N_7922,N_7671);
xnor U8466 (N_8466,N_8041,N_7999);
nor U8467 (N_8467,N_8245,N_8086);
and U8468 (N_8468,N_7524,N_7763);
xor U8469 (N_8469,N_8165,N_7602);
nand U8470 (N_8470,N_8037,N_7920);
and U8471 (N_8471,N_7546,N_7911);
or U8472 (N_8472,N_8228,N_8157);
xnor U8473 (N_8473,N_8187,N_7979);
and U8474 (N_8474,N_8019,N_7827);
or U8475 (N_8475,N_7792,N_7702);
xnor U8476 (N_8476,N_7589,N_7672);
or U8477 (N_8477,N_7634,N_7866);
xnor U8478 (N_8478,N_8065,N_7593);
or U8479 (N_8479,N_7506,N_7677);
or U8480 (N_8480,N_7764,N_7531);
nand U8481 (N_8481,N_7540,N_8180);
or U8482 (N_8482,N_7516,N_7977);
nor U8483 (N_8483,N_7687,N_8166);
nand U8484 (N_8484,N_8173,N_7692);
nor U8485 (N_8485,N_7840,N_7895);
and U8486 (N_8486,N_7619,N_7614);
and U8487 (N_8487,N_8010,N_7504);
nor U8488 (N_8488,N_7560,N_7743);
or U8489 (N_8489,N_7924,N_7574);
xnor U8490 (N_8490,N_8219,N_7562);
xnor U8491 (N_8491,N_8067,N_7638);
nor U8492 (N_8492,N_8012,N_7851);
xor U8493 (N_8493,N_8110,N_7654);
or U8494 (N_8494,N_7575,N_7694);
and U8495 (N_8495,N_8023,N_7675);
nand U8496 (N_8496,N_8192,N_8164);
xnor U8497 (N_8497,N_7530,N_8090);
nor U8498 (N_8498,N_8132,N_7865);
nand U8499 (N_8499,N_8200,N_8230);
and U8500 (N_8500,N_8177,N_8025);
or U8501 (N_8501,N_7896,N_7712);
xor U8502 (N_8502,N_7725,N_7776);
and U8503 (N_8503,N_7888,N_7783);
or U8504 (N_8504,N_7902,N_7784);
nand U8505 (N_8505,N_8076,N_8156);
nor U8506 (N_8506,N_7891,N_8232);
or U8507 (N_8507,N_7919,N_8244);
nand U8508 (N_8508,N_7668,N_7940);
or U8509 (N_8509,N_7735,N_7944);
and U8510 (N_8510,N_8095,N_7645);
nand U8511 (N_8511,N_8167,N_8223);
or U8512 (N_8512,N_7537,N_8055);
and U8513 (N_8513,N_8183,N_8204);
and U8514 (N_8514,N_7854,N_8069);
xor U8515 (N_8515,N_7580,N_7681);
nand U8516 (N_8516,N_8142,N_7935);
nand U8517 (N_8517,N_8093,N_8092);
and U8518 (N_8518,N_7661,N_7794);
xor U8519 (N_8519,N_7680,N_8203);
and U8520 (N_8520,N_7522,N_7601);
or U8521 (N_8521,N_8139,N_8155);
and U8522 (N_8522,N_7806,N_7525);
or U8523 (N_8523,N_7988,N_7697);
xnor U8524 (N_8524,N_7836,N_8070);
xor U8525 (N_8525,N_8107,N_7557);
or U8526 (N_8526,N_7750,N_7586);
xor U8527 (N_8527,N_8011,N_7829);
nand U8528 (N_8528,N_7867,N_8005);
nand U8529 (N_8529,N_8118,N_7936);
nand U8530 (N_8530,N_8064,N_8104);
nor U8531 (N_8531,N_8126,N_7969);
nand U8532 (N_8532,N_8047,N_7623);
and U8533 (N_8533,N_7947,N_7997);
xnor U8534 (N_8534,N_7811,N_8130);
nand U8535 (N_8535,N_8238,N_8242);
and U8536 (N_8536,N_8122,N_7682);
nand U8537 (N_8537,N_7740,N_8063);
nand U8538 (N_8538,N_8080,N_8024);
and U8539 (N_8539,N_7579,N_7676);
nand U8540 (N_8540,N_7861,N_7959);
or U8541 (N_8541,N_7850,N_7781);
and U8542 (N_8542,N_8206,N_7930);
or U8543 (N_8543,N_7766,N_7821);
nor U8544 (N_8544,N_8209,N_8096);
nor U8545 (N_8545,N_7810,N_7639);
nor U8546 (N_8546,N_7808,N_8218);
or U8547 (N_8547,N_8225,N_8234);
and U8548 (N_8548,N_8152,N_7961);
nor U8549 (N_8549,N_7739,N_7928);
nor U8550 (N_8550,N_7769,N_7777);
xor U8551 (N_8551,N_8154,N_7942);
nand U8552 (N_8552,N_7604,N_8101);
and U8553 (N_8553,N_7541,N_7658);
and U8554 (N_8554,N_7805,N_7587);
or U8555 (N_8555,N_7616,N_7842);
or U8556 (N_8556,N_7958,N_8038);
nor U8557 (N_8557,N_7964,N_7938);
nand U8558 (N_8558,N_8082,N_8215);
nor U8559 (N_8559,N_7721,N_7757);
or U8560 (N_8560,N_7987,N_7960);
and U8561 (N_8561,N_8241,N_7894);
and U8562 (N_8562,N_7566,N_7653);
nor U8563 (N_8563,N_7669,N_7655);
or U8564 (N_8564,N_7561,N_7598);
and U8565 (N_8565,N_8026,N_8009);
or U8566 (N_8566,N_7848,N_8199);
and U8567 (N_8567,N_8098,N_7945);
nor U8568 (N_8568,N_7708,N_7893);
or U8569 (N_8569,N_8186,N_7613);
nand U8570 (N_8570,N_7752,N_7772);
and U8571 (N_8571,N_7932,N_7873);
xnor U8572 (N_8572,N_7984,N_7974);
nand U8573 (N_8573,N_8172,N_7686);
nand U8574 (N_8574,N_7599,N_7651);
or U8575 (N_8575,N_7746,N_7759);
and U8576 (N_8576,N_7981,N_7832);
nor U8577 (N_8577,N_7612,N_7621);
xor U8578 (N_8578,N_7933,N_7914);
or U8579 (N_8579,N_8189,N_8136);
nor U8580 (N_8580,N_7745,N_7874);
nand U8581 (N_8581,N_7656,N_7526);
xor U8582 (N_8582,N_7549,N_8084);
nor U8583 (N_8583,N_8205,N_8111);
xnor U8584 (N_8584,N_7798,N_7978);
xnor U8585 (N_8585,N_7980,N_7640);
and U8586 (N_8586,N_8007,N_7703);
nor U8587 (N_8587,N_8075,N_8109);
nor U8588 (N_8588,N_7819,N_7931);
xnor U8589 (N_8589,N_7994,N_8179);
nand U8590 (N_8590,N_7771,N_8176);
or U8591 (N_8591,N_8043,N_8148);
xor U8592 (N_8592,N_7631,N_7620);
xnor U8593 (N_8593,N_7843,N_7648);
or U8594 (N_8594,N_7718,N_8103);
and U8595 (N_8595,N_8151,N_7971);
xnor U8596 (N_8596,N_7973,N_8235);
nor U8597 (N_8597,N_7591,N_7533);
or U8598 (N_8598,N_7847,N_7820);
nand U8599 (N_8599,N_8060,N_8150);
and U8600 (N_8600,N_7571,N_7849);
nand U8601 (N_8601,N_8145,N_7605);
and U8602 (N_8602,N_7730,N_7872);
nand U8603 (N_8603,N_7765,N_7635);
nor U8604 (N_8604,N_8059,N_7972);
nor U8605 (N_8605,N_8017,N_8072);
or U8606 (N_8606,N_7515,N_7796);
nand U8607 (N_8607,N_7950,N_8190);
nor U8608 (N_8608,N_8030,N_8117);
nor U8609 (N_8609,N_7782,N_7511);
or U8610 (N_8610,N_8102,N_7830);
xor U8611 (N_8611,N_7828,N_7569);
and U8612 (N_8612,N_7898,N_7662);
nand U8613 (N_8613,N_8042,N_7521);
nor U8614 (N_8614,N_7760,N_8115);
nand U8615 (N_8615,N_7844,N_7659);
xnor U8616 (N_8616,N_7699,N_8034);
nor U8617 (N_8617,N_7941,N_7738);
nand U8618 (N_8618,N_8113,N_8137);
xnor U8619 (N_8619,N_8128,N_7884);
nor U8620 (N_8620,N_7986,N_7982);
and U8621 (N_8621,N_7582,N_8221);
and U8622 (N_8622,N_7717,N_7597);
xor U8623 (N_8623,N_7713,N_8100);
nor U8624 (N_8624,N_8198,N_8248);
nand U8625 (N_8625,N_8056,N_8032);
and U8626 (N_8626,N_7626,N_7997);
or U8627 (N_8627,N_8064,N_8089);
nand U8628 (N_8628,N_8180,N_8056);
nor U8629 (N_8629,N_7769,N_7763);
nand U8630 (N_8630,N_7731,N_8007);
nor U8631 (N_8631,N_7823,N_7769);
xnor U8632 (N_8632,N_7584,N_8142);
nor U8633 (N_8633,N_7725,N_7641);
nand U8634 (N_8634,N_7873,N_7831);
nand U8635 (N_8635,N_8212,N_7621);
nand U8636 (N_8636,N_8010,N_7751);
nand U8637 (N_8637,N_7869,N_7708);
nand U8638 (N_8638,N_7983,N_8007);
nor U8639 (N_8639,N_8201,N_7993);
nand U8640 (N_8640,N_7778,N_7587);
or U8641 (N_8641,N_7581,N_7945);
nand U8642 (N_8642,N_7607,N_8110);
and U8643 (N_8643,N_8132,N_7932);
xnor U8644 (N_8644,N_7944,N_7662);
and U8645 (N_8645,N_7828,N_7652);
xnor U8646 (N_8646,N_7803,N_8160);
nor U8647 (N_8647,N_7888,N_7645);
and U8648 (N_8648,N_8007,N_8036);
nor U8649 (N_8649,N_7653,N_7728);
xor U8650 (N_8650,N_7745,N_7566);
xnor U8651 (N_8651,N_7989,N_8231);
nor U8652 (N_8652,N_8051,N_7892);
nand U8653 (N_8653,N_7898,N_8215);
xnor U8654 (N_8654,N_8005,N_7802);
nor U8655 (N_8655,N_7571,N_8169);
nand U8656 (N_8656,N_7656,N_7790);
and U8657 (N_8657,N_8245,N_8148);
xnor U8658 (N_8658,N_7659,N_7909);
or U8659 (N_8659,N_8155,N_7561);
xor U8660 (N_8660,N_7986,N_7914);
xnor U8661 (N_8661,N_7783,N_7720);
and U8662 (N_8662,N_7833,N_8173);
nor U8663 (N_8663,N_8209,N_7500);
or U8664 (N_8664,N_8161,N_7818);
nor U8665 (N_8665,N_8199,N_8133);
nor U8666 (N_8666,N_7980,N_7533);
or U8667 (N_8667,N_7862,N_7951);
and U8668 (N_8668,N_7773,N_7677);
xor U8669 (N_8669,N_7593,N_7781);
nand U8670 (N_8670,N_7838,N_8183);
and U8671 (N_8671,N_8142,N_8183);
or U8672 (N_8672,N_7769,N_8099);
nand U8673 (N_8673,N_7969,N_8000);
nor U8674 (N_8674,N_7766,N_7741);
and U8675 (N_8675,N_7639,N_8100);
and U8676 (N_8676,N_8149,N_8014);
and U8677 (N_8677,N_7766,N_8102);
nor U8678 (N_8678,N_7634,N_8231);
nor U8679 (N_8679,N_7516,N_8123);
or U8680 (N_8680,N_7555,N_7604);
or U8681 (N_8681,N_7929,N_7709);
nor U8682 (N_8682,N_8057,N_8072);
nor U8683 (N_8683,N_7673,N_7828);
nand U8684 (N_8684,N_7589,N_7950);
nor U8685 (N_8685,N_7552,N_8068);
nand U8686 (N_8686,N_8025,N_7850);
nor U8687 (N_8687,N_7926,N_7689);
nand U8688 (N_8688,N_7879,N_7719);
nor U8689 (N_8689,N_7560,N_7529);
or U8690 (N_8690,N_7703,N_7994);
or U8691 (N_8691,N_8136,N_8181);
nand U8692 (N_8692,N_7777,N_8187);
nand U8693 (N_8693,N_8135,N_7560);
or U8694 (N_8694,N_8236,N_7927);
nand U8695 (N_8695,N_7533,N_7504);
xnor U8696 (N_8696,N_7799,N_7615);
and U8697 (N_8697,N_8194,N_7635);
and U8698 (N_8698,N_8030,N_7673);
nand U8699 (N_8699,N_7662,N_7820);
xnor U8700 (N_8700,N_7685,N_8057);
nand U8701 (N_8701,N_7607,N_8005);
or U8702 (N_8702,N_7917,N_7602);
or U8703 (N_8703,N_7750,N_7761);
and U8704 (N_8704,N_7973,N_7524);
xor U8705 (N_8705,N_7608,N_8044);
or U8706 (N_8706,N_8021,N_7935);
nor U8707 (N_8707,N_8124,N_8132);
nor U8708 (N_8708,N_7977,N_8044);
or U8709 (N_8709,N_8207,N_8150);
and U8710 (N_8710,N_7608,N_8056);
or U8711 (N_8711,N_7804,N_7502);
xnor U8712 (N_8712,N_7669,N_8073);
and U8713 (N_8713,N_7604,N_7639);
nand U8714 (N_8714,N_7676,N_7838);
or U8715 (N_8715,N_8016,N_7534);
or U8716 (N_8716,N_7555,N_8137);
and U8717 (N_8717,N_8112,N_8030);
or U8718 (N_8718,N_7586,N_7666);
nor U8719 (N_8719,N_7991,N_7774);
or U8720 (N_8720,N_7630,N_7758);
xor U8721 (N_8721,N_7972,N_7697);
nand U8722 (N_8722,N_8119,N_7928);
and U8723 (N_8723,N_8164,N_7817);
or U8724 (N_8724,N_7862,N_7549);
and U8725 (N_8725,N_7686,N_7781);
and U8726 (N_8726,N_8197,N_7517);
or U8727 (N_8727,N_7688,N_8173);
nor U8728 (N_8728,N_7604,N_7715);
nor U8729 (N_8729,N_7753,N_8095);
nor U8730 (N_8730,N_8083,N_7925);
or U8731 (N_8731,N_7556,N_7716);
and U8732 (N_8732,N_8067,N_7965);
or U8733 (N_8733,N_7553,N_7696);
nand U8734 (N_8734,N_8113,N_7819);
and U8735 (N_8735,N_7605,N_7878);
and U8736 (N_8736,N_7679,N_7656);
xnor U8737 (N_8737,N_7695,N_7981);
or U8738 (N_8738,N_7992,N_7794);
or U8739 (N_8739,N_7920,N_8094);
nand U8740 (N_8740,N_8187,N_7590);
or U8741 (N_8741,N_7519,N_7830);
xor U8742 (N_8742,N_7912,N_7757);
or U8743 (N_8743,N_7810,N_8175);
or U8744 (N_8744,N_8001,N_7598);
nand U8745 (N_8745,N_7852,N_7978);
nor U8746 (N_8746,N_8049,N_7725);
xor U8747 (N_8747,N_7808,N_8225);
nor U8748 (N_8748,N_7677,N_8017);
or U8749 (N_8749,N_8016,N_7511);
xnor U8750 (N_8750,N_7946,N_7836);
nor U8751 (N_8751,N_7889,N_8042);
and U8752 (N_8752,N_7669,N_8044);
xor U8753 (N_8753,N_8145,N_8126);
xor U8754 (N_8754,N_7980,N_7793);
nor U8755 (N_8755,N_7917,N_7783);
nand U8756 (N_8756,N_8147,N_8101);
nand U8757 (N_8757,N_7634,N_7752);
xor U8758 (N_8758,N_8149,N_7728);
nor U8759 (N_8759,N_7790,N_7614);
or U8760 (N_8760,N_7504,N_8103);
xnor U8761 (N_8761,N_8195,N_7923);
nor U8762 (N_8762,N_7994,N_8139);
nor U8763 (N_8763,N_7529,N_7568);
nand U8764 (N_8764,N_7501,N_7736);
xor U8765 (N_8765,N_7976,N_7925);
xnor U8766 (N_8766,N_7951,N_7917);
xor U8767 (N_8767,N_7619,N_8142);
nor U8768 (N_8768,N_7765,N_7873);
or U8769 (N_8769,N_7705,N_7642);
nand U8770 (N_8770,N_8067,N_7754);
nand U8771 (N_8771,N_7612,N_7834);
nor U8772 (N_8772,N_7674,N_7729);
nor U8773 (N_8773,N_8100,N_7602);
nor U8774 (N_8774,N_8111,N_8206);
xnor U8775 (N_8775,N_8211,N_7578);
and U8776 (N_8776,N_8111,N_7781);
nor U8777 (N_8777,N_8070,N_7564);
or U8778 (N_8778,N_8105,N_7821);
or U8779 (N_8779,N_7924,N_8109);
nor U8780 (N_8780,N_7946,N_8069);
and U8781 (N_8781,N_7983,N_8082);
and U8782 (N_8782,N_8025,N_7956);
and U8783 (N_8783,N_7937,N_7593);
and U8784 (N_8784,N_7697,N_7927);
or U8785 (N_8785,N_7501,N_7984);
xor U8786 (N_8786,N_8191,N_8067);
and U8787 (N_8787,N_8198,N_7816);
nor U8788 (N_8788,N_8146,N_8126);
nand U8789 (N_8789,N_7923,N_7736);
or U8790 (N_8790,N_7685,N_7852);
nand U8791 (N_8791,N_8017,N_7860);
nor U8792 (N_8792,N_8219,N_7519);
and U8793 (N_8793,N_7572,N_7709);
nand U8794 (N_8794,N_7638,N_8026);
nand U8795 (N_8795,N_7594,N_7810);
xnor U8796 (N_8796,N_8051,N_7895);
nor U8797 (N_8797,N_7511,N_8088);
xor U8798 (N_8798,N_8011,N_8017);
nand U8799 (N_8799,N_7696,N_7715);
nand U8800 (N_8800,N_7569,N_7647);
xor U8801 (N_8801,N_7739,N_7822);
xnor U8802 (N_8802,N_7713,N_7887);
nand U8803 (N_8803,N_7904,N_7736);
nor U8804 (N_8804,N_7879,N_7728);
or U8805 (N_8805,N_8082,N_7721);
nand U8806 (N_8806,N_8076,N_7501);
nor U8807 (N_8807,N_7820,N_8064);
nand U8808 (N_8808,N_7540,N_7548);
and U8809 (N_8809,N_7803,N_8052);
or U8810 (N_8810,N_7522,N_7663);
xnor U8811 (N_8811,N_7931,N_7912);
and U8812 (N_8812,N_7658,N_7660);
xor U8813 (N_8813,N_8115,N_7866);
nand U8814 (N_8814,N_8224,N_7774);
nand U8815 (N_8815,N_8172,N_8073);
xor U8816 (N_8816,N_7695,N_8170);
and U8817 (N_8817,N_7568,N_7823);
nand U8818 (N_8818,N_7685,N_7521);
xnor U8819 (N_8819,N_7828,N_8034);
nand U8820 (N_8820,N_7986,N_7582);
nand U8821 (N_8821,N_7771,N_7866);
nand U8822 (N_8822,N_7649,N_8214);
or U8823 (N_8823,N_8117,N_7583);
and U8824 (N_8824,N_7885,N_7570);
nor U8825 (N_8825,N_7694,N_7885);
nor U8826 (N_8826,N_8196,N_7513);
nor U8827 (N_8827,N_8060,N_8248);
nor U8828 (N_8828,N_8091,N_8232);
and U8829 (N_8829,N_7631,N_7932);
and U8830 (N_8830,N_7996,N_7994);
or U8831 (N_8831,N_7951,N_7582);
xnor U8832 (N_8832,N_8240,N_8158);
and U8833 (N_8833,N_7706,N_7930);
or U8834 (N_8834,N_8097,N_8079);
or U8835 (N_8835,N_7552,N_7502);
nand U8836 (N_8836,N_7555,N_8158);
nand U8837 (N_8837,N_8239,N_7672);
nand U8838 (N_8838,N_7831,N_8012);
or U8839 (N_8839,N_7942,N_7867);
and U8840 (N_8840,N_8113,N_7820);
or U8841 (N_8841,N_7551,N_7588);
xor U8842 (N_8842,N_7543,N_8094);
nor U8843 (N_8843,N_7881,N_7590);
nand U8844 (N_8844,N_8209,N_7584);
or U8845 (N_8845,N_7868,N_7911);
nor U8846 (N_8846,N_8179,N_8245);
nand U8847 (N_8847,N_8228,N_7569);
xnor U8848 (N_8848,N_7705,N_7656);
or U8849 (N_8849,N_7889,N_7865);
nor U8850 (N_8850,N_7775,N_8016);
xor U8851 (N_8851,N_7520,N_8235);
or U8852 (N_8852,N_7521,N_7775);
xnor U8853 (N_8853,N_8120,N_7857);
or U8854 (N_8854,N_7757,N_7988);
nand U8855 (N_8855,N_7653,N_7886);
xnor U8856 (N_8856,N_8207,N_7654);
nor U8857 (N_8857,N_8151,N_7627);
xor U8858 (N_8858,N_7794,N_7510);
xor U8859 (N_8859,N_7678,N_8217);
nand U8860 (N_8860,N_7554,N_7854);
xor U8861 (N_8861,N_8179,N_8010);
nand U8862 (N_8862,N_7944,N_7994);
nand U8863 (N_8863,N_7881,N_7598);
and U8864 (N_8864,N_7735,N_8179);
nor U8865 (N_8865,N_8014,N_7634);
or U8866 (N_8866,N_8203,N_7641);
nand U8867 (N_8867,N_8170,N_8049);
nor U8868 (N_8868,N_8109,N_7911);
xnor U8869 (N_8869,N_8246,N_8192);
nor U8870 (N_8870,N_7824,N_8055);
nor U8871 (N_8871,N_7535,N_8049);
and U8872 (N_8872,N_7980,N_7987);
or U8873 (N_8873,N_7587,N_8245);
nor U8874 (N_8874,N_7906,N_8222);
xnor U8875 (N_8875,N_8172,N_7981);
nand U8876 (N_8876,N_7652,N_8125);
and U8877 (N_8877,N_7534,N_7966);
or U8878 (N_8878,N_8120,N_8127);
nor U8879 (N_8879,N_7904,N_7834);
nor U8880 (N_8880,N_8198,N_8184);
or U8881 (N_8881,N_8129,N_7508);
nor U8882 (N_8882,N_7548,N_7725);
xor U8883 (N_8883,N_7538,N_8007);
and U8884 (N_8884,N_7697,N_7932);
or U8885 (N_8885,N_7681,N_8214);
nand U8886 (N_8886,N_7817,N_7961);
nor U8887 (N_8887,N_7830,N_7899);
or U8888 (N_8888,N_7957,N_7982);
nor U8889 (N_8889,N_8025,N_8134);
xor U8890 (N_8890,N_7902,N_8182);
nand U8891 (N_8891,N_7682,N_7902);
nor U8892 (N_8892,N_8039,N_7853);
or U8893 (N_8893,N_7706,N_7542);
or U8894 (N_8894,N_8187,N_7645);
nand U8895 (N_8895,N_8246,N_8035);
xnor U8896 (N_8896,N_7794,N_7629);
or U8897 (N_8897,N_7946,N_8090);
or U8898 (N_8898,N_8143,N_7735);
or U8899 (N_8899,N_7739,N_8050);
and U8900 (N_8900,N_7764,N_7885);
or U8901 (N_8901,N_7772,N_7907);
nand U8902 (N_8902,N_8007,N_8141);
and U8903 (N_8903,N_8076,N_7803);
xnor U8904 (N_8904,N_8210,N_7838);
or U8905 (N_8905,N_7679,N_7504);
xor U8906 (N_8906,N_8023,N_8127);
nand U8907 (N_8907,N_7522,N_8186);
xor U8908 (N_8908,N_8092,N_8156);
xor U8909 (N_8909,N_7806,N_7946);
or U8910 (N_8910,N_8042,N_7929);
xnor U8911 (N_8911,N_7648,N_7683);
nand U8912 (N_8912,N_7859,N_7878);
and U8913 (N_8913,N_8190,N_7540);
or U8914 (N_8914,N_8205,N_7863);
nand U8915 (N_8915,N_7904,N_8056);
nand U8916 (N_8916,N_8002,N_7567);
nand U8917 (N_8917,N_8063,N_7793);
xnor U8918 (N_8918,N_7897,N_8080);
nor U8919 (N_8919,N_7884,N_8147);
nor U8920 (N_8920,N_7879,N_7557);
nand U8921 (N_8921,N_7637,N_7524);
and U8922 (N_8922,N_7574,N_7992);
nor U8923 (N_8923,N_7540,N_7946);
nor U8924 (N_8924,N_7726,N_7680);
nand U8925 (N_8925,N_7687,N_8046);
xnor U8926 (N_8926,N_8112,N_7918);
nor U8927 (N_8927,N_7709,N_8098);
xnor U8928 (N_8928,N_7851,N_7529);
nor U8929 (N_8929,N_7805,N_7964);
nor U8930 (N_8930,N_7585,N_8059);
nor U8931 (N_8931,N_7983,N_7829);
or U8932 (N_8932,N_8057,N_7966);
and U8933 (N_8933,N_7608,N_8238);
and U8934 (N_8934,N_7566,N_7638);
or U8935 (N_8935,N_7821,N_8235);
or U8936 (N_8936,N_8053,N_7953);
or U8937 (N_8937,N_7535,N_7698);
or U8938 (N_8938,N_8145,N_7697);
xor U8939 (N_8939,N_7916,N_8012);
nor U8940 (N_8940,N_8121,N_7778);
and U8941 (N_8941,N_8059,N_7679);
xnor U8942 (N_8942,N_8232,N_7963);
nand U8943 (N_8943,N_7682,N_7784);
xnor U8944 (N_8944,N_8071,N_8005);
nor U8945 (N_8945,N_7527,N_7723);
nor U8946 (N_8946,N_7568,N_8185);
or U8947 (N_8947,N_8234,N_7770);
or U8948 (N_8948,N_7802,N_7936);
and U8949 (N_8949,N_7936,N_7509);
nor U8950 (N_8950,N_7731,N_7626);
nand U8951 (N_8951,N_7756,N_7708);
nor U8952 (N_8952,N_7700,N_8034);
and U8953 (N_8953,N_7798,N_7634);
nor U8954 (N_8954,N_7864,N_8043);
or U8955 (N_8955,N_7837,N_7615);
xor U8956 (N_8956,N_7500,N_7526);
or U8957 (N_8957,N_7526,N_7738);
nor U8958 (N_8958,N_7648,N_8005);
and U8959 (N_8959,N_8112,N_8015);
nor U8960 (N_8960,N_7799,N_8113);
or U8961 (N_8961,N_8036,N_7927);
xnor U8962 (N_8962,N_7908,N_7671);
nor U8963 (N_8963,N_7547,N_7885);
or U8964 (N_8964,N_7979,N_7582);
nand U8965 (N_8965,N_7736,N_7946);
nor U8966 (N_8966,N_7817,N_8003);
or U8967 (N_8967,N_7946,N_7979);
or U8968 (N_8968,N_8198,N_8073);
nand U8969 (N_8969,N_8055,N_7593);
and U8970 (N_8970,N_7915,N_7692);
and U8971 (N_8971,N_8086,N_8043);
and U8972 (N_8972,N_8061,N_8211);
nor U8973 (N_8973,N_7621,N_7941);
or U8974 (N_8974,N_8045,N_7697);
and U8975 (N_8975,N_7544,N_7935);
xnor U8976 (N_8976,N_8143,N_8166);
xnor U8977 (N_8977,N_8181,N_7950);
nand U8978 (N_8978,N_8051,N_7734);
nand U8979 (N_8979,N_7872,N_7947);
and U8980 (N_8980,N_8234,N_7733);
or U8981 (N_8981,N_7849,N_7672);
and U8982 (N_8982,N_7535,N_7582);
and U8983 (N_8983,N_7944,N_7942);
or U8984 (N_8984,N_8166,N_7928);
nand U8985 (N_8985,N_7902,N_7749);
nand U8986 (N_8986,N_7966,N_8204);
xnor U8987 (N_8987,N_8184,N_8200);
nand U8988 (N_8988,N_7739,N_7762);
or U8989 (N_8989,N_7804,N_7839);
nor U8990 (N_8990,N_8203,N_7528);
nand U8991 (N_8991,N_7964,N_7980);
and U8992 (N_8992,N_7759,N_8026);
nand U8993 (N_8993,N_7621,N_8096);
nor U8994 (N_8994,N_8107,N_7701);
xor U8995 (N_8995,N_8056,N_7816);
xor U8996 (N_8996,N_7928,N_7701);
or U8997 (N_8997,N_8168,N_7685);
and U8998 (N_8998,N_7765,N_8122);
nand U8999 (N_8999,N_8020,N_7978);
xor U9000 (N_9000,N_8632,N_8811);
or U9001 (N_9001,N_8521,N_8756);
nor U9002 (N_9002,N_8305,N_8358);
or U9003 (N_9003,N_8751,N_8735);
xor U9004 (N_9004,N_8889,N_8458);
nor U9005 (N_9005,N_8444,N_8495);
or U9006 (N_9006,N_8609,N_8368);
nand U9007 (N_9007,N_8283,N_8800);
or U9008 (N_9008,N_8586,N_8380);
or U9009 (N_9009,N_8834,N_8562);
or U9010 (N_9010,N_8804,N_8369);
and U9011 (N_9011,N_8456,N_8560);
nor U9012 (N_9012,N_8610,N_8439);
or U9013 (N_9013,N_8443,N_8440);
or U9014 (N_9014,N_8436,N_8429);
and U9015 (N_9015,N_8888,N_8573);
nand U9016 (N_9016,N_8294,N_8809);
and U9017 (N_9017,N_8943,N_8907);
and U9018 (N_9018,N_8359,N_8490);
nor U9019 (N_9019,N_8334,N_8664);
nand U9020 (N_9020,N_8396,N_8445);
nand U9021 (N_9021,N_8417,N_8281);
xnor U9022 (N_9022,N_8864,N_8308);
nor U9023 (N_9023,N_8416,N_8386);
nand U9024 (N_9024,N_8457,N_8556);
xnor U9025 (N_9025,N_8506,N_8652);
xnor U9026 (N_9026,N_8718,N_8851);
and U9027 (N_9027,N_8534,N_8553);
and U9028 (N_9028,N_8975,N_8381);
or U9029 (N_9029,N_8746,N_8651);
nor U9030 (N_9030,N_8934,N_8961);
xor U9031 (N_9031,N_8401,N_8295);
xnor U9032 (N_9032,N_8977,N_8917);
xnor U9033 (N_9033,N_8788,N_8335);
nand U9034 (N_9034,N_8894,N_8402);
or U9035 (N_9035,N_8845,N_8284);
nor U9036 (N_9036,N_8450,N_8503);
or U9037 (N_9037,N_8611,N_8320);
and U9038 (N_9038,N_8944,N_8302);
nor U9039 (N_9039,N_8715,N_8557);
nor U9040 (N_9040,N_8890,N_8647);
nor U9041 (N_9041,N_8345,N_8683);
and U9042 (N_9042,N_8668,N_8307);
xnor U9043 (N_9043,N_8828,N_8921);
xnor U9044 (N_9044,N_8790,N_8929);
nand U9045 (N_9045,N_8676,N_8687);
nand U9046 (N_9046,N_8291,N_8625);
xor U9047 (N_9047,N_8517,N_8862);
nand U9048 (N_9048,N_8914,N_8780);
xor U9049 (N_9049,N_8645,N_8777);
nor U9050 (N_9050,N_8985,N_8261);
nand U9051 (N_9051,N_8768,N_8903);
and U9052 (N_9052,N_8707,N_8466);
nand U9053 (N_9053,N_8955,N_8564);
nand U9054 (N_9054,N_8455,N_8460);
and U9055 (N_9055,N_8518,N_8839);
nand U9056 (N_9056,N_8689,N_8430);
nor U9057 (N_9057,N_8354,N_8824);
nand U9058 (N_9058,N_8877,N_8315);
xnor U9059 (N_9059,N_8761,N_8940);
nor U9060 (N_9060,N_8298,N_8960);
or U9061 (N_9061,N_8974,N_8920);
nand U9062 (N_9062,N_8542,N_8885);
xor U9063 (N_9063,N_8643,N_8304);
nor U9064 (N_9064,N_8447,N_8323);
or U9065 (N_9065,N_8759,N_8696);
and U9066 (N_9066,N_8962,N_8479);
and U9067 (N_9067,N_8372,N_8478);
xor U9068 (N_9068,N_8724,N_8822);
or U9069 (N_9069,N_8523,N_8462);
or U9070 (N_9070,N_8282,N_8438);
xor U9071 (N_9071,N_8277,N_8814);
and U9072 (N_9072,N_8448,N_8374);
nand U9073 (N_9073,N_8679,N_8391);
nor U9074 (N_9074,N_8700,N_8898);
nand U9075 (N_9075,N_8642,N_8474);
xor U9076 (N_9076,N_8451,N_8719);
or U9077 (N_9077,N_8978,N_8703);
xnor U9078 (N_9078,N_8883,N_8485);
and U9079 (N_9079,N_8784,N_8729);
and U9080 (N_9080,N_8522,N_8615);
xnor U9081 (N_9081,N_8584,N_8398);
nor U9082 (N_9082,N_8858,N_8312);
nor U9083 (N_9083,N_8856,N_8730);
and U9084 (N_9084,N_8721,N_8336);
and U9085 (N_9085,N_8293,N_8774);
xnor U9086 (N_9086,N_8971,N_8531);
xor U9087 (N_9087,N_8324,N_8952);
and U9088 (N_9088,N_8484,N_8525);
nand U9089 (N_9089,N_8410,N_8569);
or U9090 (N_9090,N_8966,N_8378);
and U9091 (N_9091,N_8434,N_8734);
nor U9092 (N_9092,N_8453,N_8633);
and U9093 (N_9093,N_8594,N_8502);
nor U9094 (N_9094,N_8912,N_8639);
nand U9095 (N_9095,N_8526,N_8829);
xnor U9096 (N_9096,N_8667,N_8988);
nor U9097 (N_9097,N_8379,N_8571);
xor U9098 (N_9098,N_8566,N_8861);
nand U9099 (N_9099,N_8798,N_8841);
or U9100 (N_9100,N_8793,N_8688);
nand U9101 (N_9101,N_8904,N_8637);
or U9102 (N_9102,N_8537,N_8911);
or U9103 (N_9103,N_8626,N_8675);
nand U9104 (N_9104,N_8886,N_8329);
nand U9105 (N_9105,N_8390,N_8420);
nor U9106 (N_9106,N_8548,N_8674);
xnor U9107 (N_9107,N_8599,N_8601);
or U9108 (N_9108,N_8343,N_8844);
or U9109 (N_9109,N_8749,N_8596);
and U9110 (N_9110,N_8579,N_8412);
and U9111 (N_9111,N_8499,N_8832);
nand U9112 (N_9112,N_8972,N_8692);
and U9113 (N_9113,N_8252,N_8946);
xor U9114 (N_9114,N_8909,N_8311);
xnor U9115 (N_9115,N_8538,N_8422);
or U9116 (N_9116,N_8899,N_8426);
or U9117 (N_9117,N_8635,N_8303);
nor U9118 (N_9118,N_8591,N_8658);
nor U9119 (N_9119,N_8551,N_8792);
nand U9120 (N_9120,N_8547,N_8810);
nor U9121 (N_9121,N_8482,N_8732);
nor U9122 (N_9122,N_8554,N_8980);
xnor U9123 (N_9123,N_8684,N_8661);
xor U9124 (N_9124,N_8605,N_8701);
xnor U9125 (N_9125,N_8278,N_8769);
xor U9126 (N_9126,N_8949,N_8736);
or U9127 (N_9127,N_8857,N_8916);
xor U9128 (N_9128,N_8737,N_8322);
nor U9129 (N_9129,N_8817,N_8991);
and U9130 (N_9130,N_8572,N_8570);
nor U9131 (N_9131,N_8698,N_8640);
nand U9132 (N_9132,N_8338,N_8748);
and U9133 (N_9133,N_8446,N_8775);
xnor U9134 (N_9134,N_8519,N_8947);
and U9135 (N_9135,N_8382,N_8357);
nor U9136 (N_9136,N_8849,N_8567);
and U9137 (N_9137,N_8908,N_8987);
nand U9138 (N_9138,N_8470,N_8835);
and U9139 (N_9139,N_8452,N_8404);
nand U9140 (N_9140,N_8831,N_8901);
or U9141 (N_9141,N_8956,N_8524);
xor U9142 (N_9142,N_8848,N_8257);
or U9143 (N_9143,N_8937,N_8654);
and U9144 (N_9144,N_8863,N_8648);
xnor U9145 (N_9145,N_8767,N_8913);
nand U9146 (N_9146,N_8786,N_8589);
or U9147 (N_9147,N_8866,N_8253);
nand U9148 (N_9148,N_8339,N_8353);
and U9149 (N_9149,N_8942,N_8580);
and U9150 (N_9150,N_8672,N_8500);
nor U9151 (N_9151,N_8896,N_8869);
and U9152 (N_9152,N_8906,N_8389);
nor U9153 (N_9153,N_8649,N_8799);
or U9154 (N_9154,N_8879,N_8982);
xor U9155 (N_9155,N_8263,N_8623);
xnor U9156 (N_9156,N_8710,N_8983);
and U9157 (N_9157,N_8530,N_8431);
or U9158 (N_9158,N_8641,N_8424);
xnor U9159 (N_9159,N_8833,N_8741);
or U9160 (N_9160,N_8527,N_8405);
or U9161 (N_9161,N_8878,N_8581);
or U9162 (N_9162,N_8301,N_8875);
nand U9163 (N_9163,N_8744,N_8680);
or U9164 (N_9164,N_8990,N_8691);
xnor U9165 (N_9165,N_8273,N_8384);
and U9166 (N_9166,N_8319,N_8747);
nand U9167 (N_9167,N_8475,N_8727);
nor U9168 (N_9168,N_8627,N_8363);
nand U9169 (N_9169,N_8976,N_8763);
nand U9170 (N_9170,N_8713,N_8468);
nand U9171 (N_9171,N_8331,N_8510);
or U9172 (N_9172,N_8613,N_8771);
and U9173 (N_9173,N_8840,N_8669);
xnor U9174 (N_9174,N_8598,N_8264);
xor U9175 (N_9175,N_8481,N_8393);
xnor U9176 (N_9176,N_8532,N_8954);
xnor U9177 (N_9177,N_8826,N_8433);
nor U9178 (N_9178,N_8583,N_8435);
xor U9179 (N_9179,N_8418,N_8483);
or U9180 (N_9180,N_8789,N_8493);
nand U9181 (N_9181,N_8770,N_8967);
or U9182 (N_9182,N_8515,N_8344);
nor U9183 (N_9183,N_8795,N_8272);
or U9184 (N_9184,N_8997,N_8620);
nand U9185 (N_9185,N_8529,N_8590);
nand U9186 (N_9186,N_8881,N_8803);
and U9187 (N_9187,N_8406,N_8365);
xor U9188 (N_9188,N_8816,N_8708);
or U9189 (N_9189,N_8773,N_8340);
xor U9190 (N_9190,N_8563,N_8373);
nor U9191 (N_9191,N_8663,N_8449);
or U9192 (N_9192,N_8876,N_8853);
nand U9193 (N_9193,N_8606,N_8818);
and U9194 (N_9194,N_8964,N_8267);
or U9195 (N_9195,N_8738,N_8656);
nor U9196 (N_9196,N_8309,N_8604);
xor U9197 (N_9197,N_8544,N_8859);
and U9198 (N_9198,N_8505,N_8758);
nand U9199 (N_9199,N_8603,N_8720);
nor U9200 (N_9200,N_8965,N_8897);
and U9201 (N_9201,N_8860,N_8677);
xor U9202 (N_9202,N_8797,N_8552);
nand U9203 (N_9203,N_8880,N_8593);
and U9204 (N_9204,N_8968,N_8785);
or U9205 (N_9205,N_8513,N_8993);
nor U9206 (N_9206,N_8614,N_8694);
nor U9207 (N_9207,N_8480,N_8351);
nand U9208 (N_9208,N_8926,N_8815);
or U9209 (N_9209,N_8995,N_8948);
xnor U9210 (N_9210,N_8459,N_8884);
nor U9211 (N_9211,N_8731,N_8671);
xor U9212 (N_9212,N_8388,N_8313);
xor U9213 (N_9213,N_8910,N_8805);
nand U9214 (N_9214,N_8742,N_8998);
nand U9215 (N_9215,N_8427,N_8699);
nand U9216 (N_9216,N_8260,N_8408);
and U9217 (N_9217,N_8992,N_8873);
nor U9218 (N_9218,N_8726,N_8289);
nand U9219 (N_9219,N_8488,N_8394);
xnor U9220 (N_9220,N_8508,N_8565);
nor U9221 (N_9221,N_8621,N_8932);
or U9222 (N_9222,N_8546,N_8709);
nor U9223 (N_9223,N_8516,N_8489);
nor U9224 (N_9224,N_8825,N_8356);
and U9225 (N_9225,N_8745,N_8791);
xnor U9226 (N_9226,N_8270,N_8855);
nand U9227 (N_9227,N_8360,N_8364);
or U9228 (N_9228,N_8938,N_8778);
or U9229 (N_9229,N_8782,N_8653);
and U9230 (N_9230,N_8690,N_8256);
and U9231 (N_9231,N_8491,N_8600);
and U9232 (N_9232,N_8325,N_8755);
nand U9233 (N_9233,N_8963,N_8612);
xnor U9234 (N_9234,N_8595,N_8843);
nand U9235 (N_9235,N_8285,N_8712);
and U9236 (N_9236,N_8678,N_8919);
xor U9237 (N_9237,N_8432,N_8650);
or U9238 (N_9238,N_8695,N_8941);
nand U9239 (N_9239,N_8762,N_8865);
nor U9240 (N_9240,N_8414,N_8882);
and U9241 (N_9241,N_8383,N_8628);
or U9242 (N_9242,N_8801,N_8662);
nand U9243 (N_9243,N_8413,N_8437);
nor U9244 (N_9244,N_8366,N_8665);
and U9245 (N_9245,N_8409,N_8629);
and U9246 (N_9246,N_8574,N_8617);
and U9247 (N_9247,N_8918,N_8607);
nor U9248 (N_9248,N_8922,N_8870);
xnor U9249 (N_9249,N_8415,N_8387);
xnor U9250 (N_9250,N_8928,N_8330);
xnor U9251 (N_9251,N_8268,N_8300);
nand U9252 (N_9252,N_8702,N_8332);
nand U9253 (N_9253,N_8924,N_8631);
xor U9254 (N_9254,N_8638,N_8830);
xnor U9255 (N_9255,N_8504,N_8706);
and U9256 (N_9256,N_8492,N_8874);
and U9257 (N_9257,N_8765,N_8403);
nand U9258 (N_9258,N_8397,N_8867);
and U9259 (N_9259,N_8314,N_8464);
nor U9260 (N_9260,N_8266,N_8535);
xnor U9261 (N_9261,N_8723,N_8717);
xnor U9262 (N_9262,N_8469,N_8827);
or U9263 (N_9263,N_8578,N_8370);
nor U9264 (N_9264,N_8346,N_8276);
or U9265 (N_9265,N_8711,N_8931);
xor U9266 (N_9266,N_8984,N_8528);
or U9267 (N_9267,N_8533,N_8757);
and U9268 (N_9268,N_8377,N_8655);
or U9269 (N_9269,N_8618,N_8539);
or U9270 (N_9270,N_8644,N_8986);
or U9271 (N_9271,N_8872,N_8476);
nand U9272 (N_9272,N_8685,N_8520);
xor U9273 (N_9273,N_8622,N_8561);
and U9274 (N_9274,N_8395,N_8750);
or U9275 (N_9275,N_8821,N_8487);
and U9276 (N_9276,N_8996,N_8673);
nand U9277 (N_9277,N_8959,N_8576);
nor U9278 (N_9278,N_8902,N_8250);
or U9279 (N_9279,N_8787,N_8989);
or U9280 (N_9280,N_8740,N_8496);
or U9281 (N_9281,N_8477,N_8682);
or U9282 (N_9282,N_8973,N_8465);
or U9283 (N_9283,N_8288,N_8296);
and U9284 (N_9284,N_8779,N_8287);
xnor U9285 (N_9285,N_8497,N_8321);
nor U9286 (N_9286,N_8752,N_8543);
nor U9287 (N_9287,N_8616,N_8290);
nand U9288 (N_9288,N_8292,N_8802);
xor U9289 (N_9289,N_8254,N_8498);
nor U9290 (N_9290,N_8341,N_8274);
xnor U9291 (N_9291,N_8636,N_8507);
nor U9292 (N_9292,N_8392,N_8355);
and U9293 (N_9293,N_8608,N_8582);
or U9294 (N_9294,N_8969,N_8597);
or U9295 (N_9295,N_8783,N_8286);
xor U9296 (N_9296,N_8999,N_8419);
or U9297 (N_9297,N_8349,N_8316);
nand U9298 (N_9298,N_8352,N_8258);
or U9299 (N_9299,N_8697,N_8933);
or U9300 (N_9300,N_8299,N_8850);
or U9301 (N_9301,N_8714,N_8776);
and U9302 (N_9302,N_8337,N_8376);
xor U9303 (N_9303,N_8945,N_8951);
and U9304 (N_9304,N_8753,N_8536);
xnor U9305 (N_9305,N_8385,N_8900);
xor U9306 (N_9306,N_8754,N_8838);
nor U9307 (N_9307,N_8494,N_8820);
xnor U9308 (N_9308,N_8550,N_8486);
or U9309 (N_9309,N_8808,N_8472);
nand U9310 (N_9310,N_8425,N_8887);
nand U9311 (N_9311,N_8326,N_8255);
nor U9312 (N_9312,N_8297,N_8367);
nor U9313 (N_9313,N_8812,N_8407);
or U9314 (N_9314,N_8442,N_8950);
and U9315 (N_9315,N_8362,N_8588);
xor U9316 (N_9316,N_8743,N_8939);
xor U9317 (N_9317,N_8957,N_8893);
nor U9318 (N_9318,N_8265,N_8807);
xor U9319 (N_9319,N_8927,N_8577);
nor U9320 (N_9320,N_8806,N_8936);
xnor U9321 (N_9321,N_8471,N_8994);
or U9322 (N_9322,N_8657,N_8728);
xnor U9323 (N_9323,N_8852,N_8646);
or U9324 (N_9324,N_8764,N_8411);
nand U9325 (N_9325,N_8371,N_8318);
nand U9326 (N_9326,N_8423,N_8514);
xnor U9327 (N_9327,N_8558,N_8251);
nor U9328 (N_9328,N_8509,N_8512);
nor U9329 (N_9329,N_8630,N_8819);
nor U9330 (N_9330,N_8733,N_8361);
nand U9331 (N_9331,N_8935,N_8327);
and U9332 (N_9332,N_8794,N_8463);
or U9333 (N_9333,N_8634,N_8905);
nor U9334 (N_9334,N_8399,N_8317);
and U9335 (N_9335,N_8739,N_8953);
nor U9336 (N_9336,N_8400,N_8259);
nand U9337 (N_9337,N_8280,N_8979);
xor U9338 (N_9338,N_8306,N_8823);
and U9339 (N_9339,N_8541,N_8781);
xnor U9340 (N_9340,N_8981,N_8347);
and U9341 (N_9341,N_8722,N_8310);
xor U9342 (N_9342,N_8846,N_8915);
nand U9343 (N_9343,N_8847,N_8842);
and U9344 (N_9344,N_8568,N_8836);
nand U9345 (N_9345,N_8725,N_8421);
nor U9346 (N_9346,N_8660,N_8624);
nor U9347 (N_9347,N_8587,N_8760);
nor U9348 (N_9348,N_8559,N_8585);
and U9349 (N_9349,N_8441,N_8473);
nor U9350 (N_9350,N_8958,N_8461);
and U9351 (N_9351,N_8271,N_8333);
and U9352 (N_9352,N_8930,N_8545);
nor U9353 (N_9353,N_8262,N_8813);
nand U9354 (N_9354,N_8923,N_8467);
or U9355 (N_9355,N_8895,N_8275);
nand U9356 (N_9356,N_8837,N_8772);
nor U9357 (N_9357,N_8348,N_8269);
nand U9358 (N_9358,N_8892,N_8511);
xor U9359 (N_9359,N_8350,N_8619);
or U9360 (N_9360,N_8659,N_8375);
and U9361 (N_9361,N_8705,N_8681);
nor U9362 (N_9362,N_8970,N_8549);
nor U9363 (N_9363,N_8575,N_8501);
xnor U9364 (N_9364,N_8540,N_8454);
nor U9365 (N_9365,N_8328,N_8796);
nand U9366 (N_9366,N_8555,N_8592);
xnor U9367 (N_9367,N_8871,N_8686);
xnor U9368 (N_9368,N_8704,N_8666);
or U9369 (N_9369,N_8693,N_8279);
or U9370 (N_9370,N_8602,N_8854);
and U9371 (N_9371,N_8891,N_8428);
nand U9372 (N_9372,N_8716,N_8868);
nand U9373 (N_9373,N_8670,N_8766);
or U9374 (N_9374,N_8342,N_8925);
nor U9375 (N_9375,N_8880,N_8294);
or U9376 (N_9376,N_8722,N_8812);
xnor U9377 (N_9377,N_8845,N_8913);
or U9378 (N_9378,N_8895,N_8954);
nor U9379 (N_9379,N_8566,N_8500);
nor U9380 (N_9380,N_8678,N_8579);
xor U9381 (N_9381,N_8470,N_8299);
xor U9382 (N_9382,N_8907,N_8350);
and U9383 (N_9383,N_8981,N_8665);
nor U9384 (N_9384,N_8768,N_8532);
nor U9385 (N_9385,N_8281,N_8428);
or U9386 (N_9386,N_8881,N_8636);
nor U9387 (N_9387,N_8698,N_8728);
nand U9388 (N_9388,N_8644,N_8621);
nand U9389 (N_9389,N_8545,N_8838);
or U9390 (N_9390,N_8642,N_8899);
nor U9391 (N_9391,N_8687,N_8440);
nor U9392 (N_9392,N_8364,N_8467);
or U9393 (N_9393,N_8483,N_8704);
xor U9394 (N_9394,N_8344,N_8724);
nand U9395 (N_9395,N_8758,N_8616);
xnor U9396 (N_9396,N_8707,N_8728);
or U9397 (N_9397,N_8322,N_8272);
nor U9398 (N_9398,N_8681,N_8574);
xnor U9399 (N_9399,N_8656,N_8851);
nor U9400 (N_9400,N_8863,N_8401);
or U9401 (N_9401,N_8272,N_8703);
or U9402 (N_9402,N_8832,N_8866);
xnor U9403 (N_9403,N_8822,N_8543);
or U9404 (N_9404,N_8595,N_8760);
nor U9405 (N_9405,N_8532,N_8673);
nand U9406 (N_9406,N_8879,N_8872);
and U9407 (N_9407,N_8317,N_8876);
xor U9408 (N_9408,N_8535,N_8690);
nand U9409 (N_9409,N_8565,N_8322);
and U9410 (N_9410,N_8329,N_8714);
xnor U9411 (N_9411,N_8796,N_8486);
and U9412 (N_9412,N_8866,N_8294);
or U9413 (N_9413,N_8545,N_8826);
nor U9414 (N_9414,N_8529,N_8592);
xnor U9415 (N_9415,N_8889,N_8499);
xor U9416 (N_9416,N_8487,N_8793);
xor U9417 (N_9417,N_8674,N_8319);
nand U9418 (N_9418,N_8398,N_8771);
nand U9419 (N_9419,N_8688,N_8356);
and U9420 (N_9420,N_8583,N_8814);
nor U9421 (N_9421,N_8516,N_8476);
nor U9422 (N_9422,N_8824,N_8741);
or U9423 (N_9423,N_8689,N_8329);
and U9424 (N_9424,N_8580,N_8562);
nand U9425 (N_9425,N_8953,N_8429);
nor U9426 (N_9426,N_8678,N_8663);
nor U9427 (N_9427,N_8674,N_8934);
or U9428 (N_9428,N_8252,N_8701);
nand U9429 (N_9429,N_8829,N_8911);
or U9430 (N_9430,N_8866,N_8471);
xor U9431 (N_9431,N_8271,N_8693);
nor U9432 (N_9432,N_8261,N_8862);
nor U9433 (N_9433,N_8644,N_8788);
xor U9434 (N_9434,N_8854,N_8379);
nor U9435 (N_9435,N_8385,N_8268);
or U9436 (N_9436,N_8661,N_8845);
xnor U9437 (N_9437,N_8918,N_8799);
nand U9438 (N_9438,N_8348,N_8315);
xnor U9439 (N_9439,N_8998,N_8918);
nand U9440 (N_9440,N_8927,N_8425);
nor U9441 (N_9441,N_8515,N_8430);
nor U9442 (N_9442,N_8795,N_8877);
or U9443 (N_9443,N_8728,N_8759);
or U9444 (N_9444,N_8487,N_8569);
and U9445 (N_9445,N_8292,N_8865);
nor U9446 (N_9446,N_8994,N_8535);
and U9447 (N_9447,N_8291,N_8712);
xnor U9448 (N_9448,N_8658,N_8302);
and U9449 (N_9449,N_8760,N_8265);
xor U9450 (N_9450,N_8319,N_8548);
nand U9451 (N_9451,N_8997,N_8417);
xnor U9452 (N_9452,N_8567,N_8680);
xnor U9453 (N_9453,N_8483,N_8326);
or U9454 (N_9454,N_8500,N_8847);
nor U9455 (N_9455,N_8306,N_8759);
or U9456 (N_9456,N_8722,N_8645);
nand U9457 (N_9457,N_8763,N_8845);
and U9458 (N_9458,N_8718,N_8974);
xnor U9459 (N_9459,N_8692,N_8308);
or U9460 (N_9460,N_8573,N_8715);
nor U9461 (N_9461,N_8778,N_8639);
nor U9462 (N_9462,N_8329,N_8986);
xnor U9463 (N_9463,N_8834,N_8299);
nand U9464 (N_9464,N_8937,N_8966);
nand U9465 (N_9465,N_8823,N_8976);
xor U9466 (N_9466,N_8968,N_8721);
and U9467 (N_9467,N_8562,N_8469);
xor U9468 (N_9468,N_8899,N_8491);
or U9469 (N_9469,N_8436,N_8542);
nand U9470 (N_9470,N_8374,N_8464);
or U9471 (N_9471,N_8290,N_8760);
nor U9472 (N_9472,N_8709,N_8831);
and U9473 (N_9473,N_8340,N_8477);
or U9474 (N_9474,N_8577,N_8493);
xor U9475 (N_9475,N_8767,N_8709);
xor U9476 (N_9476,N_8943,N_8502);
nand U9477 (N_9477,N_8607,N_8565);
nor U9478 (N_9478,N_8928,N_8887);
nor U9479 (N_9479,N_8695,N_8309);
nor U9480 (N_9480,N_8564,N_8660);
nor U9481 (N_9481,N_8835,N_8383);
or U9482 (N_9482,N_8596,N_8815);
nor U9483 (N_9483,N_8976,N_8256);
nand U9484 (N_9484,N_8287,N_8373);
and U9485 (N_9485,N_8537,N_8276);
nor U9486 (N_9486,N_8989,N_8467);
xor U9487 (N_9487,N_8534,N_8515);
nor U9488 (N_9488,N_8634,N_8859);
and U9489 (N_9489,N_8444,N_8335);
or U9490 (N_9490,N_8831,N_8793);
xnor U9491 (N_9491,N_8423,N_8810);
nand U9492 (N_9492,N_8877,N_8573);
xor U9493 (N_9493,N_8498,N_8257);
and U9494 (N_9494,N_8760,N_8653);
and U9495 (N_9495,N_8464,N_8511);
nor U9496 (N_9496,N_8955,N_8898);
and U9497 (N_9497,N_8898,N_8584);
xnor U9498 (N_9498,N_8558,N_8550);
nor U9499 (N_9499,N_8884,N_8390);
nor U9500 (N_9500,N_8359,N_8312);
xnor U9501 (N_9501,N_8735,N_8302);
nor U9502 (N_9502,N_8351,N_8310);
and U9503 (N_9503,N_8989,N_8524);
and U9504 (N_9504,N_8371,N_8761);
or U9505 (N_9505,N_8567,N_8394);
nor U9506 (N_9506,N_8397,N_8759);
nand U9507 (N_9507,N_8566,N_8467);
or U9508 (N_9508,N_8903,N_8327);
nor U9509 (N_9509,N_8386,N_8992);
or U9510 (N_9510,N_8546,N_8586);
xnor U9511 (N_9511,N_8363,N_8431);
or U9512 (N_9512,N_8804,N_8327);
nand U9513 (N_9513,N_8443,N_8869);
and U9514 (N_9514,N_8509,N_8984);
and U9515 (N_9515,N_8650,N_8816);
or U9516 (N_9516,N_8636,N_8753);
and U9517 (N_9517,N_8763,N_8697);
nand U9518 (N_9518,N_8471,N_8911);
or U9519 (N_9519,N_8680,N_8463);
and U9520 (N_9520,N_8701,N_8552);
nor U9521 (N_9521,N_8864,N_8497);
or U9522 (N_9522,N_8341,N_8380);
nor U9523 (N_9523,N_8345,N_8724);
xnor U9524 (N_9524,N_8798,N_8286);
or U9525 (N_9525,N_8481,N_8764);
nor U9526 (N_9526,N_8955,N_8571);
xor U9527 (N_9527,N_8265,N_8874);
or U9528 (N_9528,N_8533,N_8510);
and U9529 (N_9529,N_8759,N_8385);
or U9530 (N_9530,N_8867,N_8365);
xor U9531 (N_9531,N_8307,N_8542);
or U9532 (N_9532,N_8600,N_8578);
and U9533 (N_9533,N_8363,N_8910);
nand U9534 (N_9534,N_8392,N_8827);
nand U9535 (N_9535,N_8455,N_8881);
and U9536 (N_9536,N_8757,N_8272);
or U9537 (N_9537,N_8753,N_8577);
xnor U9538 (N_9538,N_8875,N_8408);
or U9539 (N_9539,N_8628,N_8901);
nand U9540 (N_9540,N_8629,N_8318);
and U9541 (N_9541,N_8390,N_8769);
nand U9542 (N_9542,N_8702,N_8980);
or U9543 (N_9543,N_8926,N_8950);
nor U9544 (N_9544,N_8361,N_8661);
xor U9545 (N_9545,N_8798,N_8980);
xnor U9546 (N_9546,N_8659,N_8888);
nor U9547 (N_9547,N_8656,N_8476);
xnor U9548 (N_9548,N_8259,N_8351);
nor U9549 (N_9549,N_8425,N_8575);
or U9550 (N_9550,N_8990,N_8386);
nand U9551 (N_9551,N_8666,N_8760);
and U9552 (N_9552,N_8986,N_8322);
nand U9553 (N_9553,N_8784,N_8302);
nand U9554 (N_9554,N_8882,N_8575);
xor U9555 (N_9555,N_8630,N_8796);
nor U9556 (N_9556,N_8349,N_8809);
and U9557 (N_9557,N_8357,N_8455);
or U9558 (N_9558,N_8299,N_8677);
xnor U9559 (N_9559,N_8787,N_8920);
nand U9560 (N_9560,N_8412,N_8334);
or U9561 (N_9561,N_8707,N_8809);
or U9562 (N_9562,N_8644,N_8431);
nor U9563 (N_9563,N_8930,N_8725);
xnor U9564 (N_9564,N_8320,N_8890);
xnor U9565 (N_9565,N_8312,N_8347);
or U9566 (N_9566,N_8887,N_8791);
nor U9567 (N_9567,N_8900,N_8675);
or U9568 (N_9568,N_8331,N_8436);
nor U9569 (N_9569,N_8265,N_8753);
nor U9570 (N_9570,N_8484,N_8956);
nor U9571 (N_9571,N_8886,N_8539);
xor U9572 (N_9572,N_8711,N_8591);
xor U9573 (N_9573,N_8256,N_8899);
and U9574 (N_9574,N_8842,N_8349);
nor U9575 (N_9575,N_8692,N_8258);
nor U9576 (N_9576,N_8625,N_8392);
nand U9577 (N_9577,N_8676,N_8667);
nor U9578 (N_9578,N_8614,N_8396);
nor U9579 (N_9579,N_8741,N_8349);
xnor U9580 (N_9580,N_8499,N_8463);
nand U9581 (N_9581,N_8851,N_8953);
nor U9582 (N_9582,N_8512,N_8754);
nor U9583 (N_9583,N_8854,N_8958);
and U9584 (N_9584,N_8462,N_8262);
or U9585 (N_9585,N_8762,N_8501);
nand U9586 (N_9586,N_8319,N_8568);
nor U9587 (N_9587,N_8802,N_8918);
and U9588 (N_9588,N_8877,N_8913);
xor U9589 (N_9589,N_8505,N_8989);
nand U9590 (N_9590,N_8536,N_8539);
or U9591 (N_9591,N_8520,N_8944);
nor U9592 (N_9592,N_8430,N_8334);
and U9593 (N_9593,N_8262,N_8406);
or U9594 (N_9594,N_8619,N_8841);
nor U9595 (N_9595,N_8275,N_8368);
and U9596 (N_9596,N_8864,N_8615);
and U9597 (N_9597,N_8989,N_8259);
or U9598 (N_9598,N_8349,N_8479);
nand U9599 (N_9599,N_8895,N_8392);
xnor U9600 (N_9600,N_8516,N_8450);
and U9601 (N_9601,N_8910,N_8295);
and U9602 (N_9602,N_8266,N_8378);
nor U9603 (N_9603,N_8932,N_8360);
or U9604 (N_9604,N_8551,N_8734);
nand U9605 (N_9605,N_8494,N_8734);
xor U9606 (N_9606,N_8743,N_8855);
nor U9607 (N_9607,N_8964,N_8504);
and U9608 (N_9608,N_8307,N_8514);
or U9609 (N_9609,N_8510,N_8529);
nand U9610 (N_9610,N_8710,N_8587);
nand U9611 (N_9611,N_8652,N_8522);
xnor U9612 (N_9612,N_8710,N_8679);
nand U9613 (N_9613,N_8260,N_8703);
or U9614 (N_9614,N_8452,N_8390);
or U9615 (N_9615,N_8574,N_8625);
or U9616 (N_9616,N_8812,N_8321);
nor U9617 (N_9617,N_8925,N_8816);
nor U9618 (N_9618,N_8873,N_8954);
xnor U9619 (N_9619,N_8796,N_8460);
nor U9620 (N_9620,N_8955,N_8828);
nor U9621 (N_9621,N_8927,N_8728);
and U9622 (N_9622,N_8408,N_8688);
and U9623 (N_9623,N_8272,N_8584);
xnor U9624 (N_9624,N_8330,N_8477);
nor U9625 (N_9625,N_8569,N_8806);
nor U9626 (N_9626,N_8805,N_8519);
xor U9627 (N_9627,N_8563,N_8850);
nand U9628 (N_9628,N_8694,N_8259);
xor U9629 (N_9629,N_8569,N_8948);
or U9630 (N_9630,N_8295,N_8646);
nand U9631 (N_9631,N_8990,N_8288);
and U9632 (N_9632,N_8883,N_8764);
or U9633 (N_9633,N_8644,N_8982);
nand U9634 (N_9634,N_8795,N_8766);
nand U9635 (N_9635,N_8380,N_8927);
and U9636 (N_9636,N_8508,N_8313);
or U9637 (N_9637,N_8753,N_8946);
and U9638 (N_9638,N_8922,N_8634);
or U9639 (N_9639,N_8597,N_8432);
and U9640 (N_9640,N_8935,N_8797);
nand U9641 (N_9641,N_8603,N_8946);
nand U9642 (N_9642,N_8258,N_8646);
xnor U9643 (N_9643,N_8617,N_8695);
xnor U9644 (N_9644,N_8673,N_8388);
and U9645 (N_9645,N_8500,N_8867);
nor U9646 (N_9646,N_8895,N_8992);
nor U9647 (N_9647,N_8741,N_8761);
and U9648 (N_9648,N_8785,N_8468);
and U9649 (N_9649,N_8895,N_8744);
nor U9650 (N_9650,N_8622,N_8790);
and U9651 (N_9651,N_8721,N_8307);
and U9652 (N_9652,N_8318,N_8608);
and U9653 (N_9653,N_8950,N_8307);
nor U9654 (N_9654,N_8408,N_8988);
and U9655 (N_9655,N_8850,N_8790);
nor U9656 (N_9656,N_8314,N_8474);
and U9657 (N_9657,N_8701,N_8699);
nor U9658 (N_9658,N_8360,N_8917);
nor U9659 (N_9659,N_8956,N_8833);
xor U9660 (N_9660,N_8271,N_8574);
or U9661 (N_9661,N_8309,N_8331);
nor U9662 (N_9662,N_8439,N_8882);
nand U9663 (N_9663,N_8888,N_8639);
or U9664 (N_9664,N_8523,N_8959);
nand U9665 (N_9665,N_8780,N_8575);
xor U9666 (N_9666,N_8806,N_8755);
and U9667 (N_9667,N_8572,N_8325);
or U9668 (N_9668,N_8918,N_8741);
and U9669 (N_9669,N_8534,N_8568);
xnor U9670 (N_9670,N_8341,N_8634);
nor U9671 (N_9671,N_8889,N_8997);
and U9672 (N_9672,N_8678,N_8881);
nor U9673 (N_9673,N_8731,N_8775);
nand U9674 (N_9674,N_8948,N_8606);
or U9675 (N_9675,N_8489,N_8396);
xnor U9676 (N_9676,N_8481,N_8968);
nand U9677 (N_9677,N_8748,N_8741);
xor U9678 (N_9678,N_8763,N_8715);
and U9679 (N_9679,N_8641,N_8253);
nand U9680 (N_9680,N_8985,N_8676);
and U9681 (N_9681,N_8335,N_8690);
or U9682 (N_9682,N_8268,N_8311);
or U9683 (N_9683,N_8764,N_8634);
or U9684 (N_9684,N_8995,N_8496);
nor U9685 (N_9685,N_8544,N_8674);
xnor U9686 (N_9686,N_8280,N_8807);
or U9687 (N_9687,N_8354,N_8450);
xor U9688 (N_9688,N_8263,N_8464);
and U9689 (N_9689,N_8913,N_8663);
nor U9690 (N_9690,N_8569,N_8858);
xor U9691 (N_9691,N_8258,N_8314);
nor U9692 (N_9692,N_8575,N_8732);
nor U9693 (N_9693,N_8297,N_8958);
xnor U9694 (N_9694,N_8272,N_8740);
nor U9695 (N_9695,N_8777,N_8607);
xnor U9696 (N_9696,N_8919,N_8293);
xor U9697 (N_9697,N_8355,N_8845);
nand U9698 (N_9698,N_8730,N_8565);
or U9699 (N_9699,N_8320,N_8894);
nand U9700 (N_9700,N_8645,N_8664);
nor U9701 (N_9701,N_8663,N_8514);
xnor U9702 (N_9702,N_8372,N_8819);
nor U9703 (N_9703,N_8333,N_8687);
nand U9704 (N_9704,N_8452,N_8606);
nor U9705 (N_9705,N_8793,N_8540);
nor U9706 (N_9706,N_8482,N_8818);
xor U9707 (N_9707,N_8586,N_8439);
and U9708 (N_9708,N_8543,N_8747);
xor U9709 (N_9709,N_8263,N_8752);
or U9710 (N_9710,N_8449,N_8500);
nand U9711 (N_9711,N_8361,N_8443);
or U9712 (N_9712,N_8595,N_8410);
or U9713 (N_9713,N_8307,N_8300);
nand U9714 (N_9714,N_8310,N_8551);
nand U9715 (N_9715,N_8836,N_8471);
nand U9716 (N_9716,N_8287,N_8448);
nand U9717 (N_9717,N_8520,N_8642);
nor U9718 (N_9718,N_8998,N_8806);
or U9719 (N_9719,N_8407,N_8845);
nand U9720 (N_9720,N_8746,N_8890);
and U9721 (N_9721,N_8717,N_8463);
nand U9722 (N_9722,N_8653,N_8548);
nand U9723 (N_9723,N_8544,N_8384);
nor U9724 (N_9724,N_8840,N_8601);
and U9725 (N_9725,N_8269,N_8991);
nor U9726 (N_9726,N_8581,N_8656);
and U9727 (N_9727,N_8619,N_8672);
or U9728 (N_9728,N_8893,N_8720);
xor U9729 (N_9729,N_8988,N_8786);
or U9730 (N_9730,N_8629,N_8875);
xnor U9731 (N_9731,N_8919,N_8253);
or U9732 (N_9732,N_8672,N_8965);
nor U9733 (N_9733,N_8412,N_8971);
xnor U9734 (N_9734,N_8727,N_8748);
or U9735 (N_9735,N_8861,N_8798);
nor U9736 (N_9736,N_8347,N_8554);
or U9737 (N_9737,N_8299,N_8831);
nand U9738 (N_9738,N_8489,N_8450);
and U9739 (N_9739,N_8839,N_8955);
nor U9740 (N_9740,N_8507,N_8841);
nor U9741 (N_9741,N_8788,N_8554);
and U9742 (N_9742,N_8579,N_8670);
or U9743 (N_9743,N_8942,N_8310);
or U9744 (N_9744,N_8539,N_8610);
or U9745 (N_9745,N_8283,N_8705);
nand U9746 (N_9746,N_8890,N_8876);
or U9747 (N_9747,N_8698,N_8327);
xor U9748 (N_9748,N_8871,N_8342);
nor U9749 (N_9749,N_8420,N_8564);
nor U9750 (N_9750,N_9363,N_9519);
nand U9751 (N_9751,N_9581,N_9611);
xnor U9752 (N_9752,N_9465,N_9466);
nand U9753 (N_9753,N_9485,N_9595);
xor U9754 (N_9754,N_9240,N_9554);
and U9755 (N_9755,N_9027,N_9518);
and U9756 (N_9756,N_9710,N_9580);
nand U9757 (N_9757,N_9103,N_9443);
and U9758 (N_9758,N_9314,N_9319);
and U9759 (N_9759,N_9736,N_9480);
nand U9760 (N_9760,N_9698,N_9468);
xnor U9761 (N_9761,N_9345,N_9128);
and U9762 (N_9762,N_9083,N_9113);
xnor U9763 (N_9763,N_9610,N_9202);
nand U9764 (N_9764,N_9009,N_9396);
nor U9765 (N_9765,N_9278,N_9725);
xnor U9766 (N_9766,N_9476,N_9196);
nand U9767 (N_9767,N_9135,N_9184);
nand U9768 (N_9768,N_9272,N_9087);
and U9769 (N_9769,N_9367,N_9530);
nand U9770 (N_9770,N_9534,N_9604);
and U9771 (N_9771,N_9420,N_9579);
nand U9772 (N_9772,N_9681,N_9139);
nand U9773 (N_9773,N_9385,N_9620);
or U9774 (N_9774,N_9423,N_9689);
nand U9775 (N_9775,N_9719,N_9539);
and U9776 (N_9776,N_9024,N_9360);
and U9777 (N_9777,N_9479,N_9524);
xor U9778 (N_9778,N_9043,N_9356);
xnor U9779 (N_9779,N_9086,N_9721);
nor U9780 (N_9780,N_9093,N_9603);
nand U9781 (N_9781,N_9124,N_9696);
and U9782 (N_9782,N_9526,N_9259);
nor U9783 (N_9783,N_9134,N_9436);
or U9784 (N_9784,N_9183,N_9156);
xor U9785 (N_9785,N_9566,N_9335);
xor U9786 (N_9786,N_9407,N_9462);
xor U9787 (N_9787,N_9256,N_9712);
nor U9788 (N_9788,N_9732,N_9310);
nand U9789 (N_9789,N_9711,N_9447);
or U9790 (N_9790,N_9397,N_9121);
or U9791 (N_9791,N_9295,N_9585);
or U9792 (N_9792,N_9498,N_9383);
and U9793 (N_9793,N_9442,N_9469);
nand U9794 (N_9794,N_9193,N_9174);
and U9795 (N_9795,N_9654,N_9302);
nand U9796 (N_9796,N_9692,N_9075);
nand U9797 (N_9797,N_9321,N_9582);
nor U9798 (N_9798,N_9092,N_9602);
and U9799 (N_9799,N_9616,N_9392);
nor U9800 (N_9800,N_9630,N_9413);
nor U9801 (N_9801,N_9746,N_9735);
xnor U9802 (N_9802,N_9490,N_9003);
xnor U9803 (N_9803,N_9250,N_9600);
nand U9804 (N_9804,N_9399,N_9085);
nand U9805 (N_9805,N_9238,N_9133);
xor U9806 (N_9806,N_9486,N_9509);
and U9807 (N_9807,N_9271,N_9306);
nand U9808 (N_9808,N_9512,N_9069);
and U9809 (N_9809,N_9346,N_9727);
or U9810 (N_9810,N_9629,N_9340);
nor U9811 (N_9811,N_9362,N_9058);
or U9812 (N_9812,N_9672,N_9145);
nor U9813 (N_9813,N_9459,N_9403);
and U9814 (N_9814,N_9387,N_9264);
or U9815 (N_9815,N_9018,N_9343);
or U9816 (N_9816,N_9263,N_9576);
nor U9817 (N_9817,N_9749,N_9472);
nor U9818 (N_9818,N_9538,N_9679);
nor U9819 (N_9819,N_9042,N_9636);
nand U9820 (N_9820,N_9214,N_9702);
nor U9821 (N_9821,N_9211,N_9478);
and U9822 (N_9822,N_9705,N_9663);
xnor U9823 (N_9823,N_9587,N_9546);
xnor U9824 (N_9824,N_9647,N_9007);
nand U9825 (N_9825,N_9531,N_9557);
nor U9826 (N_9826,N_9082,N_9073);
nor U9827 (N_9827,N_9528,N_9109);
xor U9828 (N_9828,N_9406,N_9516);
and U9829 (N_9829,N_9562,N_9243);
nand U9830 (N_9830,N_9617,N_9701);
and U9831 (N_9831,N_9285,N_9274);
nor U9832 (N_9832,N_9350,N_9066);
nor U9833 (N_9833,N_9612,N_9523);
nand U9834 (N_9834,N_9270,N_9461);
nor U9835 (N_9835,N_9181,N_9635);
or U9836 (N_9836,N_9170,N_9687);
or U9837 (N_9837,N_9716,N_9354);
or U9838 (N_9838,N_9670,N_9598);
or U9839 (N_9839,N_9703,N_9568);
nor U9840 (N_9840,N_9563,N_9377);
xnor U9841 (N_9841,N_9195,N_9107);
xor U9842 (N_9842,N_9079,N_9279);
xnor U9843 (N_9843,N_9567,N_9502);
nand U9844 (N_9844,N_9064,N_9448);
and U9845 (N_9845,N_9694,N_9400);
and U9846 (N_9846,N_9334,N_9475);
xor U9847 (N_9847,N_9232,N_9014);
nand U9848 (N_9848,N_9412,N_9305);
nand U9849 (N_9849,N_9313,N_9661);
nand U9850 (N_9850,N_9723,N_9381);
nor U9851 (N_9851,N_9105,N_9717);
nor U9852 (N_9852,N_9000,N_9131);
nor U9853 (N_9853,N_9021,N_9633);
nand U9854 (N_9854,N_9312,N_9266);
and U9855 (N_9855,N_9456,N_9347);
xnor U9856 (N_9856,N_9148,N_9330);
nand U9857 (N_9857,N_9159,N_9393);
or U9858 (N_9858,N_9618,N_9382);
and U9859 (N_9859,N_9741,N_9571);
nor U9860 (N_9860,N_9303,N_9218);
nand U9861 (N_9861,N_9053,N_9682);
nor U9862 (N_9862,N_9676,N_9652);
xnor U9863 (N_9863,N_9558,N_9414);
or U9864 (N_9864,N_9144,N_9594);
nand U9865 (N_9865,N_9253,N_9226);
or U9866 (N_9866,N_9147,N_9258);
and U9867 (N_9867,N_9451,N_9157);
and U9868 (N_9868,N_9119,N_9275);
nand U9869 (N_9869,N_9130,N_9641);
xor U9870 (N_9870,N_9491,N_9228);
nor U9871 (N_9871,N_9433,N_9287);
or U9872 (N_9872,N_9707,N_9158);
xnor U9873 (N_9873,N_9143,N_9318);
xor U9874 (N_9874,N_9316,N_9054);
nor U9875 (N_9875,N_9031,N_9065);
nor U9876 (N_9876,N_9495,N_9208);
or U9877 (N_9877,N_9199,N_9596);
or U9878 (N_9878,N_9541,N_9213);
or U9879 (N_9879,N_9146,N_9039);
or U9880 (N_9880,N_9660,N_9536);
and U9881 (N_9881,N_9508,N_9637);
nor U9882 (N_9882,N_9080,N_9578);
nor U9883 (N_9883,N_9188,N_9435);
xor U9884 (N_9884,N_9230,N_9187);
nor U9885 (N_9885,N_9454,N_9570);
and U9886 (N_9886,N_9200,N_9575);
or U9887 (N_9887,N_9606,N_9527);
or U9888 (N_9888,N_9477,N_9235);
xnor U9889 (N_9889,N_9336,N_9678);
nand U9890 (N_9890,N_9619,N_9391);
xor U9891 (N_9891,N_9368,N_9185);
xnor U9892 (N_9892,N_9004,N_9572);
nor U9893 (N_9893,N_9650,N_9286);
or U9894 (N_9894,N_9722,N_9482);
and U9895 (N_9895,N_9507,N_9683);
nor U9896 (N_9896,N_9012,N_9640);
nand U9897 (N_9897,N_9704,N_9653);
nor U9898 (N_9898,N_9201,N_9470);
xnor U9899 (N_9899,N_9709,N_9255);
or U9900 (N_9900,N_9223,N_9005);
nand U9901 (N_9901,N_9730,N_9118);
nor U9902 (N_9902,N_9658,N_9239);
nor U9903 (N_9903,N_9553,N_9404);
nor U9904 (N_9904,N_9010,N_9590);
xnor U9905 (N_9905,N_9720,N_9252);
nand U9906 (N_9906,N_9608,N_9511);
or U9907 (N_9907,N_9150,N_9104);
nor U9908 (N_9908,N_9639,N_9422);
nor U9909 (N_9909,N_9520,N_9375);
and U9910 (N_9910,N_9671,N_9047);
or U9911 (N_9911,N_9379,N_9745);
nand U9912 (N_9912,N_9055,N_9292);
and U9913 (N_9913,N_9028,N_9168);
or U9914 (N_9914,N_9550,N_9555);
nand U9915 (N_9915,N_9593,N_9645);
nand U9916 (N_9916,N_9097,N_9674);
and U9917 (N_9917,N_9127,N_9493);
and U9918 (N_9918,N_9029,N_9708);
xor U9919 (N_9919,N_9463,N_9685);
or U9920 (N_9920,N_9298,N_9409);
and U9921 (N_9921,N_9634,N_9718);
xnor U9922 (N_9922,N_9378,N_9045);
xor U9923 (N_9923,N_9438,N_9050);
nand U9924 (N_9924,N_9607,N_9457);
and U9925 (N_9925,N_9601,N_9370);
nand U9926 (N_9926,N_9338,N_9544);
nand U9927 (N_9927,N_9540,N_9504);
nor U9928 (N_9928,N_9020,N_9351);
nor U9929 (N_9929,N_9289,N_9398);
xnor U9930 (N_9930,N_9076,N_9455);
nor U9931 (N_9931,N_9388,N_9624);
nand U9932 (N_9932,N_9341,N_9237);
xor U9933 (N_9933,N_9680,N_9323);
nand U9934 (N_9934,N_9352,N_9657);
and U9935 (N_9935,N_9430,N_9098);
xor U9936 (N_9936,N_9584,N_9025);
nor U9937 (N_9937,N_9162,N_9686);
and U9938 (N_9938,N_9744,N_9215);
or U9939 (N_9939,N_9062,N_9190);
nand U9940 (N_9940,N_9372,N_9206);
or U9941 (N_9941,N_9155,N_9048);
nor U9942 (N_9942,N_9405,N_9609);
nor U9943 (N_9943,N_9434,N_9699);
nand U9944 (N_9944,N_9091,N_9643);
nand U9945 (N_9945,N_9328,N_9163);
nor U9946 (N_9946,N_9026,N_9357);
and U9947 (N_9947,N_9123,N_9090);
xnor U9948 (N_9948,N_9153,N_9551);
and U9949 (N_9949,N_9138,N_9233);
or U9950 (N_9950,N_9673,N_9542);
nor U9951 (N_9951,N_9344,N_9171);
or U9952 (N_9952,N_9577,N_9293);
nand U9953 (N_9953,N_9445,N_9217);
or U9954 (N_9954,N_9549,N_9548);
or U9955 (N_9955,N_9440,N_9458);
and U9956 (N_9956,N_9309,N_9389);
and U9957 (N_9957,N_9733,N_9429);
and U9958 (N_9958,N_9561,N_9122);
and U9959 (N_9959,N_9742,N_9591);
xnor U9960 (N_9960,N_9496,N_9160);
xor U9961 (N_9961,N_9499,N_9339);
nor U9962 (N_9962,N_9327,N_9269);
or U9963 (N_9963,N_9189,N_9035);
nand U9964 (N_9964,N_9614,N_9724);
nor U9965 (N_9965,N_9739,N_9556);
and U9966 (N_9966,N_9695,N_9222);
xor U9967 (N_9967,N_9384,N_9165);
nand U9968 (N_9968,N_9142,N_9471);
nand U9969 (N_9969,N_9311,N_9078);
or U9970 (N_9970,N_9514,N_9016);
nor U9971 (N_9971,N_9329,N_9627);
nor U9972 (N_9972,N_9547,N_9446);
and U9973 (N_9973,N_9715,N_9033);
nor U9974 (N_9974,N_9729,N_9615);
and U9975 (N_9975,N_9056,N_9517);
xor U9976 (N_9976,N_9194,N_9212);
or U9977 (N_9977,N_9693,N_9084);
nand U9978 (N_9978,N_9651,N_9236);
nand U9979 (N_9979,N_9251,N_9573);
nand U9980 (N_9980,N_9281,N_9140);
nand U9981 (N_9981,N_9649,N_9642);
nor U9982 (N_9982,N_9613,N_9592);
xor U9983 (N_9983,N_9747,N_9564);
nand U9984 (N_9984,N_9301,N_9697);
nand U9985 (N_9985,N_9129,N_9424);
nor U9986 (N_9986,N_9565,N_9099);
nor U9987 (N_9987,N_9268,N_9167);
xor U9988 (N_9988,N_9364,N_9172);
and U9989 (N_9989,N_9525,N_9068);
xor U9990 (N_9990,N_9041,N_9220);
and U9991 (N_9991,N_9116,N_9169);
and U9992 (N_9992,N_9205,N_9102);
and U9993 (N_9993,N_9246,N_9307);
and U9994 (N_9994,N_9662,N_9738);
or U9995 (N_9995,N_9605,N_9529);
nor U9996 (N_9996,N_9111,N_9728);
or U9997 (N_9997,N_9522,N_9437);
xnor U9998 (N_9998,N_9543,N_9365);
nand U9999 (N_9999,N_9115,N_9489);
nand U10000 (N_10000,N_9366,N_9164);
xor U10001 (N_10001,N_9484,N_9441);
or U10002 (N_10002,N_9234,N_9125);
and U10003 (N_10003,N_9320,N_9052);
xnor U10004 (N_10004,N_9487,N_9369);
nor U10005 (N_10005,N_9373,N_9209);
or U10006 (N_10006,N_9094,N_9261);
nand U10007 (N_10007,N_9110,N_9358);
xnor U10008 (N_10008,N_9100,N_9532);
nand U10009 (N_10009,N_9374,N_9284);
or U10010 (N_10010,N_9006,N_9081);
nor U10011 (N_10011,N_9060,N_9467);
nor U10012 (N_10012,N_9583,N_9049);
or U10013 (N_10013,N_9667,N_9276);
xnor U10014 (N_10014,N_9656,N_9108);
or U10015 (N_10015,N_9186,N_9178);
nor U10016 (N_10016,N_9669,N_9586);
xor U10017 (N_10017,N_9402,N_9452);
nand U10018 (N_10018,N_9513,N_9664);
xnor U10019 (N_10019,N_9559,N_9154);
nor U10020 (N_10020,N_9265,N_9371);
xnor U10021 (N_10021,N_9588,N_9114);
xnor U10022 (N_10022,N_9691,N_9473);
xnor U10023 (N_10023,N_9072,N_9503);
or U10024 (N_10024,N_9734,N_9057);
and U10025 (N_10025,N_9324,N_9015);
nand U10026 (N_10026,N_9501,N_9337);
or U10027 (N_10027,N_9040,N_9177);
nand U10028 (N_10028,N_9428,N_9229);
nand U10029 (N_10029,N_9515,N_9247);
or U10030 (N_10030,N_9277,N_9282);
or U10031 (N_10031,N_9677,N_9242);
nor U10032 (N_10032,N_9359,N_9019);
and U10033 (N_10033,N_9297,N_9219);
and U10034 (N_10034,N_9096,N_9149);
xor U10035 (N_10035,N_9179,N_9063);
or U10036 (N_10036,N_9221,N_9421);
and U10037 (N_10037,N_9067,N_9349);
or U10038 (N_10038,N_9101,N_9173);
nor U10039 (N_10039,N_9161,N_9488);
and U10040 (N_10040,N_9071,N_9684);
xor U10041 (N_10041,N_9304,N_9740);
nor U10042 (N_10042,N_9380,N_9748);
xor U10043 (N_10043,N_9151,N_9017);
nand U10044 (N_10044,N_9418,N_9638);
nand U10045 (N_10045,N_9227,N_9089);
xnor U10046 (N_10046,N_9700,N_9244);
or U10047 (N_10047,N_9688,N_9132);
xnor U10048 (N_10048,N_9574,N_9262);
or U10049 (N_10049,N_9023,N_9464);
nand U10050 (N_10050,N_9631,N_9505);
xor U10051 (N_10051,N_9315,N_9248);
and U10052 (N_10052,N_9494,N_9648);
or U10053 (N_10053,N_9552,N_9037);
xnor U10054 (N_10054,N_9492,N_9714);
nor U10055 (N_10055,N_9342,N_9355);
nand U10056 (N_10056,N_9506,N_9419);
xnor U10057 (N_10057,N_9521,N_9535);
or U10058 (N_10058,N_9326,N_9175);
and U10059 (N_10059,N_9308,N_9432);
and U10060 (N_10060,N_9411,N_9322);
nand U10061 (N_10061,N_9126,N_9537);
nor U10062 (N_10062,N_9625,N_9245);
nor U10063 (N_10063,N_9361,N_9449);
nand U10064 (N_10064,N_9299,N_9296);
xnor U10065 (N_10065,N_9348,N_9013);
and U10066 (N_10066,N_9626,N_9417);
or U10067 (N_10067,N_9002,N_9241);
and U10068 (N_10068,N_9332,N_9415);
and U10069 (N_10069,N_9008,N_9112);
and U10070 (N_10070,N_9300,N_9260);
xnor U10071 (N_10071,N_9408,N_9273);
nand U10072 (N_10072,N_9207,N_9401);
or U10073 (N_10073,N_9597,N_9095);
or U10074 (N_10074,N_9141,N_9666);
nor U10075 (N_10075,N_9290,N_9545);
and U10076 (N_10076,N_9569,N_9166);
xnor U10077 (N_10077,N_9197,N_9192);
xor U10078 (N_10078,N_9001,N_9743);
nor U10079 (N_10079,N_9210,N_9483);
xor U10080 (N_10080,N_9410,N_9533);
nor U10081 (N_10081,N_9152,N_9628);
xor U10082 (N_10082,N_9032,N_9390);
nor U10083 (N_10083,N_9038,N_9182);
nor U10084 (N_10084,N_9450,N_9560);
nand U10085 (N_10085,N_9386,N_9120);
and U10086 (N_10086,N_9731,N_9426);
xor U10087 (N_10087,N_9137,N_9453);
and U10088 (N_10088,N_9046,N_9225);
nor U10089 (N_10089,N_9726,N_9198);
and U10090 (N_10090,N_9257,N_9030);
nor U10091 (N_10091,N_9059,N_9621);
nor U10092 (N_10092,N_9283,N_9632);
xor U10093 (N_10093,N_9136,N_9589);
nor U10094 (N_10094,N_9706,N_9331);
or U10095 (N_10095,N_9646,N_9737);
nand U10096 (N_10096,N_9481,N_9061);
and U10097 (N_10097,N_9254,N_9077);
and U10098 (N_10098,N_9074,N_9317);
nand U10099 (N_10099,N_9249,N_9622);
or U10100 (N_10100,N_9713,N_9106);
nor U10101 (N_10101,N_9665,N_9510);
nand U10102 (N_10102,N_9325,N_9117);
and U10103 (N_10103,N_9655,N_9690);
xor U10104 (N_10104,N_9599,N_9191);
or U10105 (N_10105,N_9497,N_9288);
or U10106 (N_10106,N_9431,N_9180);
or U10107 (N_10107,N_9034,N_9036);
nand U10108 (N_10108,N_9623,N_9460);
and U10109 (N_10109,N_9394,N_9204);
nor U10110 (N_10110,N_9291,N_9659);
nor U10111 (N_10111,N_9395,N_9203);
or U10112 (N_10112,N_9231,N_9267);
nand U10113 (N_10113,N_9333,N_9376);
xor U10114 (N_10114,N_9425,N_9500);
xnor U10115 (N_10115,N_9070,N_9051);
nand U10116 (N_10116,N_9176,N_9011);
xnor U10117 (N_10117,N_9280,N_9668);
nand U10118 (N_10118,N_9444,N_9353);
and U10119 (N_10119,N_9427,N_9088);
and U10120 (N_10120,N_9416,N_9224);
and U10121 (N_10121,N_9675,N_9644);
xor U10122 (N_10122,N_9022,N_9474);
nor U10123 (N_10123,N_9216,N_9294);
and U10124 (N_10124,N_9439,N_9044);
and U10125 (N_10125,N_9471,N_9311);
nor U10126 (N_10126,N_9588,N_9671);
and U10127 (N_10127,N_9258,N_9354);
or U10128 (N_10128,N_9660,N_9520);
xnor U10129 (N_10129,N_9691,N_9059);
or U10130 (N_10130,N_9268,N_9077);
nand U10131 (N_10131,N_9250,N_9299);
or U10132 (N_10132,N_9662,N_9498);
xnor U10133 (N_10133,N_9153,N_9255);
xnor U10134 (N_10134,N_9094,N_9738);
nand U10135 (N_10135,N_9222,N_9101);
nor U10136 (N_10136,N_9390,N_9585);
xor U10137 (N_10137,N_9173,N_9412);
nor U10138 (N_10138,N_9257,N_9700);
nor U10139 (N_10139,N_9500,N_9084);
and U10140 (N_10140,N_9242,N_9715);
or U10141 (N_10141,N_9581,N_9135);
nor U10142 (N_10142,N_9671,N_9216);
xnor U10143 (N_10143,N_9527,N_9276);
or U10144 (N_10144,N_9639,N_9632);
nor U10145 (N_10145,N_9182,N_9690);
xnor U10146 (N_10146,N_9735,N_9110);
and U10147 (N_10147,N_9275,N_9579);
or U10148 (N_10148,N_9331,N_9113);
and U10149 (N_10149,N_9130,N_9347);
xnor U10150 (N_10150,N_9456,N_9606);
nor U10151 (N_10151,N_9355,N_9127);
xnor U10152 (N_10152,N_9645,N_9008);
nand U10153 (N_10153,N_9623,N_9608);
nand U10154 (N_10154,N_9375,N_9054);
nand U10155 (N_10155,N_9321,N_9567);
and U10156 (N_10156,N_9263,N_9431);
xor U10157 (N_10157,N_9190,N_9610);
xor U10158 (N_10158,N_9350,N_9526);
and U10159 (N_10159,N_9670,N_9658);
or U10160 (N_10160,N_9197,N_9499);
and U10161 (N_10161,N_9347,N_9689);
and U10162 (N_10162,N_9294,N_9295);
or U10163 (N_10163,N_9578,N_9692);
nand U10164 (N_10164,N_9254,N_9643);
and U10165 (N_10165,N_9365,N_9442);
nand U10166 (N_10166,N_9557,N_9172);
or U10167 (N_10167,N_9651,N_9704);
and U10168 (N_10168,N_9029,N_9443);
nand U10169 (N_10169,N_9569,N_9303);
or U10170 (N_10170,N_9621,N_9331);
or U10171 (N_10171,N_9661,N_9144);
and U10172 (N_10172,N_9291,N_9449);
or U10173 (N_10173,N_9232,N_9533);
xnor U10174 (N_10174,N_9310,N_9301);
and U10175 (N_10175,N_9458,N_9599);
xnor U10176 (N_10176,N_9063,N_9548);
nor U10177 (N_10177,N_9069,N_9041);
nor U10178 (N_10178,N_9384,N_9532);
xor U10179 (N_10179,N_9470,N_9539);
or U10180 (N_10180,N_9619,N_9296);
nand U10181 (N_10181,N_9732,N_9551);
or U10182 (N_10182,N_9367,N_9374);
xor U10183 (N_10183,N_9010,N_9157);
or U10184 (N_10184,N_9436,N_9313);
or U10185 (N_10185,N_9576,N_9427);
and U10186 (N_10186,N_9223,N_9268);
nand U10187 (N_10187,N_9466,N_9301);
and U10188 (N_10188,N_9694,N_9593);
and U10189 (N_10189,N_9510,N_9598);
xor U10190 (N_10190,N_9425,N_9092);
and U10191 (N_10191,N_9027,N_9062);
nor U10192 (N_10192,N_9461,N_9527);
and U10193 (N_10193,N_9062,N_9693);
xnor U10194 (N_10194,N_9079,N_9443);
xor U10195 (N_10195,N_9172,N_9163);
nand U10196 (N_10196,N_9003,N_9629);
nor U10197 (N_10197,N_9567,N_9488);
xnor U10198 (N_10198,N_9576,N_9397);
xor U10199 (N_10199,N_9628,N_9521);
and U10200 (N_10200,N_9489,N_9635);
nand U10201 (N_10201,N_9628,N_9126);
and U10202 (N_10202,N_9154,N_9535);
xor U10203 (N_10203,N_9484,N_9358);
nor U10204 (N_10204,N_9368,N_9352);
and U10205 (N_10205,N_9408,N_9553);
nor U10206 (N_10206,N_9454,N_9235);
and U10207 (N_10207,N_9743,N_9088);
or U10208 (N_10208,N_9237,N_9379);
nand U10209 (N_10209,N_9041,N_9447);
and U10210 (N_10210,N_9224,N_9143);
nor U10211 (N_10211,N_9295,N_9342);
and U10212 (N_10212,N_9547,N_9103);
or U10213 (N_10213,N_9549,N_9592);
nand U10214 (N_10214,N_9069,N_9121);
nor U10215 (N_10215,N_9075,N_9214);
xor U10216 (N_10216,N_9130,N_9036);
and U10217 (N_10217,N_9462,N_9438);
or U10218 (N_10218,N_9398,N_9230);
and U10219 (N_10219,N_9586,N_9430);
or U10220 (N_10220,N_9536,N_9097);
xnor U10221 (N_10221,N_9349,N_9077);
or U10222 (N_10222,N_9580,N_9444);
and U10223 (N_10223,N_9658,N_9447);
or U10224 (N_10224,N_9696,N_9289);
or U10225 (N_10225,N_9391,N_9035);
or U10226 (N_10226,N_9006,N_9550);
xnor U10227 (N_10227,N_9523,N_9527);
xor U10228 (N_10228,N_9108,N_9485);
and U10229 (N_10229,N_9632,N_9159);
nor U10230 (N_10230,N_9535,N_9405);
nand U10231 (N_10231,N_9278,N_9722);
and U10232 (N_10232,N_9150,N_9043);
or U10233 (N_10233,N_9180,N_9736);
nor U10234 (N_10234,N_9256,N_9526);
and U10235 (N_10235,N_9122,N_9513);
nor U10236 (N_10236,N_9488,N_9153);
nand U10237 (N_10237,N_9117,N_9573);
nor U10238 (N_10238,N_9661,N_9486);
nand U10239 (N_10239,N_9657,N_9300);
and U10240 (N_10240,N_9174,N_9031);
xor U10241 (N_10241,N_9050,N_9509);
nor U10242 (N_10242,N_9558,N_9554);
or U10243 (N_10243,N_9035,N_9701);
xor U10244 (N_10244,N_9437,N_9549);
or U10245 (N_10245,N_9202,N_9432);
and U10246 (N_10246,N_9149,N_9545);
nand U10247 (N_10247,N_9362,N_9421);
or U10248 (N_10248,N_9582,N_9094);
xnor U10249 (N_10249,N_9452,N_9215);
nand U10250 (N_10250,N_9215,N_9187);
and U10251 (N_10251,N_9337,N_9676);
nor U10252 (N_10252,N_9716,N_9164);
and U10253 (N_10253,N_9127,N_9655);
xor U10254 (N_10254,N_9668,N_9061);
nor U10255 (N_10255,N_9171,N_9124);
and U10256 (N_10256,N_9056,N_9009);
xor U10257 (N_10257,N_9102,N_9397);
or U10258 (N_10258,N_9662,N_9001);
and U10259 (N_10259,N_9271,N_9073);
xnor U10260 (N_10260,N_9722,N_9144);
nand U10261 (N_10261,N_9520,N_9675);
xnor U10262 (N_10262,N_9676,N_9227);
or U10263 (N_10263,N_9459,N_9684);
xnor U10264 (N_10264,N_9553,N_9438);
nor U10265 (N_10265,N_9583,N_9356);
and U10266 (N_10266,N_9400,N_9540);
or U10267 (N_10267,N_9236,N_9647);
and U10268 (N_10268,N_9633,N_9206);
xnor U10269 (N_10269,N_9298,N_9731);
nor U10270 (N_10270,N_9229,N_9252);
or U10271 (N_10271,N_9277,N_9725);
nand U10272 (N_10272,N_9515,N_9017);
xnor U10273 (N_10273,N_9152,N_9338);
nand U10274 (N_10274,N_9301,N_9411);
and U10275 (N_10275,N_9689,N_9377);
or U10276 (N_10276,N_9731,N_9007);
xor U10277 (N_10277,N_9025,N_9446);
and U10278 (N_10278,N_9335,N_9564);
xnor U10279 (N_10279,N_9538,N_9243);
and U10280 (N_10280,N_9087,N_9172);
or U10281 (N_10281,N_9269,N_9049);
and U10282 (N_10282,N_9562,N_9557);
nor U10283 (N_10283,N_9731,N_9154);
and U10284 (N_10284,N_9587,N_9566);
xnor U10285 (N_10285,N_9074,N_9114);
nand U10286 (N_10286,N_9052,N_9626);
xor U10287 (N_10287,N_9220,N_9296);
and U10288 (N_10288,N_9118,N_9617);
and U10289 (N_10289,N_9704,N_9207);
and U10290 (N_10290,N_9067,N_9663);
and U10291 (N_10291,N_9721,N_9294);
or U10292 (N_10292,N_9263,N_9098);
xor U10293 (N_10293,N_9576,N_9587);
and U10294 (N_10294,N_9213,N_9201);
and U10295 (N_10295,N_9585,N_9112);
nand U10296 (N_10296,N_9281,N_9110);
nand U10297 (N_10297,N_9151,N_9249);
nand U10298 (N_10298,N_9300,N_9321);
nor U10299 (N_10299,N_9149,N_9052);
xnor U10300 (N_10300,N_9597,N_9208);
nor U10301 (N_10301,N_9275,N_9298);
or U10302 (N_10302,N_9621,N_9493);
or U10303 (N_10303,N_9370,N_9244);
nor U10304 (N_10304,N_9502,N_9494);
xor U10305 (N_10305,N_9423,N_9078);
xnor U10306 (N_10306,N_9735,N_9216);
nand U10307 (N_10307,N_9592,N_9355);
or U10308 (N_10308,N_9044,N_9509);
nor U10309 (N_10309,N_9308,N_9075);
xnor U10310 (N_10310,N_9258,N_9173);
xnor U10311 (N_10311,N_9559,N_9003);
or U10312 (N_10312,N_9102,N_9489);
nand U10313 (N_10313,N_9238,N_9154);
nor U10314 (N_10314,N_9205,N_9054);
and U10315 (N_10315,N_9119,N_9192);
nand U10316 (N_10316,N_9386,N_9156);
nor U10317 (N_10317,N_9528,N_9370);
or U10318 (N_10318,N_9160,N_9290);
and U10319 (N_10319,N_9339,N_9163);
nand U10320 (N_10320,N_9510,N_9694);
nand U10321 (N_10321,N_9147,N_9162);
nor U10322 (N_10322,N_9080,N_9533);
or U10323 (N_10323,N_9244,N_9028);
nand U10324 (N_10324,N_9005,N_9709);
or U10325 (N_10325,N_9001,N_9337);
nor U10326 (N_10326,N_9320,N_9747);
or U10327 (N_10327,N_9402,N_9094);
and U10328 (N_10328,N_9169,N_9257);
xor U10329 (N_10329,N_9456,N_9517);
nor U10330 (N_10330,N_9685,N_9583);
xor U10331 (N_10331,N_9006,N_9242);
nand U10332 (N_10332,N_9415,N_9043);
nor U10333 (N_10333,N_9465,N_9521);
nand U10334 (N_10334,N_9263,N_9372);
nand U10335 (N_10335,N_9594,N_9147);
nand U10336 (N_10336,N_9311,N_9415);
and U10337 (N_10337,N_9326,N_9295);
nand U10338 (N_10338,N_9625,N_9275);
nand U10339 (N_10339,N_9720,N_9087);
or U10340 (N_10340,N_9736,N_9012);
and U10341 (N_10341,N_9669,N_9648);
and U10342 (N_10342,N_9344,N_9510);
nand U10343 (N_10343,N_9746,N_9749);
nand U10344 (N_10344,N_9272,N_9377);
and U10345 (N_10345,N_9392,N_9665);
nor U10346 (N_10346,N_9308,N_9186);
and U10347 (N_10347,N_9495,N_9326);
xnor U10348 (N_10348,N_9391,N_9026);
or U10349 (N_10349,N_9172,N_9263);
nand U10350 (N_10350,N_9391,N_9511);
nand U10351 (N_10351,N_9041,N_9726);
nor U10352 (N_10352,N_9487,N_9530);
or U10353 (N_10353,N_9192,N_9591);
and U10354 (N_10354,N_9054,N_9645);
or U10355 (N_10355,N_9293,N_9575);
xnor U10356 (N_10356,N_9656,N_9280);
and U10357 (N_10357,N_9243,N_9227);
and U10358 (N_10358,N_9602,N_9701);
or U10359 (N_10359,N_9156,N_9530);
and U10360 (N_10360,N_9157,N_9747);
nand U10361 (N_10361,N_9316,N_9405);
nand U10362 (N_10362,N_9098,N_9176);
or U10363 (N_10363,N_9748,N_9407);
xor U10364 (N_10364,N_9133,N_9742);
nor U10365 (N_10365,N_9361,N_9372);
nor U10366 (N_10366,N_9717,N_9274);
or U10367 (N_10367,N_9428,N_9478);
and U10368 (N_10368,N_9028,N_9293);
or U10369 (N_10369,N_9067,N_9462);
nand U10370 (N_10370,N_9475,N_9220);
or U10371 (N_10371,N_9079,N_9385);
and U10372 (N_10372,N_9037,N_9120);
or U10373 (N_10373,N_9711,N_9259);
nor U10374 (N_10374,N_9045,N_9368);
xor U10375 (N_10375,N_9404,N_9062);
nand U10376 (N_10376,N_9268,N_9511);
xor U10377 (N_10377,N_9029,N_9529);
or U10378 (N_10378,N_9510,N_9699);
and U10379 (N_10379,N_9394,N_9571);
or U10380 (N_10380,N_9492,N_9263);
and U10381 (N_10381,N_9456,N_9408);
xnor U10382 (N_10382,N_9651,N_9161);
and U10383 (N_10383,N_9239,N_9018);
and U10384 (N_10384,N_9559,N_9106);
xor U10385 (N_10385,N_9534,N_9711);
nand U10386 (N_10386,N_9323,N_9232);
nand U10387 (N_10387,N_9241,N_9309);
xor U10388 (N_10388,N_9190,N_9131);
nor U10389 (N_10389,N_9240,N_9645);
nand U10390 (N_10390,N_9745,N_9711);
and U10391 (N_10391,N_9384,N_9426);
and U10392 (N_10392,N_9039,N_9620);
xnor U10393 (N_10393,N_9069,N_9219);
nor U10394 (N_10394,N_9204,N_9131);
nor U10395 (N_10395,N_9358,N_9620);
nand U10396 (N_10396,N_9182,N_9053);
nand U10397 (N_10397,N_9723,N_9140);
and U10398 (N_10398,N_9167,N_9540);
and U10399 (N_10399,N_9411,N_9538);
and U10400 (N_10400,N_9038,N_9435);
xor U10401 (N_10401,N_9334,N_9528);
or U10402 (N_10402,N_9050,N_9302);
and U10403 (N_10403,N_9715,N_9445);
nand U10404 (N_10404,N_9418,N_9539);
or U10405 (N_10405,N_9115,N_9116);
and U10406 (N_10406,N_9256,N_9098);
nand U10407 (N_10407,N_9483,N_9243);
xnor U10408 (N_10408,N_9300,N_9651);
or U10409 (N_10409,N_9334,N_9462);
nor U10410 (N_10410,N_9494,N_9026);
xnor U10411 (N_10411,N_9181,N_9288);
and U10412 (N_10412,N_9443,N_9329);
nand U10413 (N_10413,N_9570,N_9639);
and U10414 (N_10414,N_9072,N_9312);
nand U10415 (N_10415,N_9176,N_9081);
and U10416 (N_10416,N_9082,N_9333);
nand U10417 (N_10417,N_9595,N_9395);
nor U10418 (N_10418,N_9447,N_9172);
or U10419 (N_10419,N_9081,N_9234);
or U10420 (N_10420,N_9219,N_9152);
or U10421 (N_10421,N_9257,N_9090);
xor U10422 (N_10422,N_9025,N_9175);
nand U10423 (N_10423,N_9271,N_9448);
or U10424 (N_10424,N_9728,N_9482);
and U10425 (N_10425,N_9701,N_9225);
xor U10426 (N_10426,N_9182,N_9100);
nand U10427 (N_10427,N_9373,N_9270);
nand U10428 (N_10428,N_9155,N_9392);
or U10429 (N_10429,N_9565,N_9647);
nor U10430 (N_10430,N_9731,N_9655);
nand U10431 (N_10431,N_9529,N_9421);
nand U10432 (N_10432,N_9036,N_9075);
xnor U10433 (N_10433,N_9028,N_9001);
nor U10434 (N_10434,N_9390,N_9186);
nand U10435 (N_10435,N_9187,N_9232);
or U10436 (N_10436,N_9255,N_9319);
or U10437 (N_10437,N_9682,N_9531);
nand U10438 (N_10438,N_9735,N_9423);
xnor U10439 (N_10439,N_9502,N_9307);
and U10440 (N_10440,N_9682,N_9187);
nand U10441 (N_10441,N_9287,N_9358);
nand U10442 (N_10442,N_9316,N_9363);
or U10443 (N_10443,N_9391,N_9305);
and U10444 (N_10444,N_9132,N_9183);
xor U10445 (N_10445,N_9628,N_9654);
xnor U10446 (N_10446,N_9697,N_9345);
xor U10447 (N_10447,N_9126,N_9067);
or U10448 (N_10448,N_9726,N_9437);
and U10449 (N_10449,N_9267,N_9289);
or U10450 (N_10450,N_9560,N_9409);
nor U10451 (N_10451,N_9170,N_9628);
or U10452 (N_10452,N_9059,N_9421);
xor U10453 (N_10453,N_9094,N_9164);
and U10454 (N_10454,N_9671,N_9432);
and U10455 (N_10455,N_9051,N_9499);
or U10456 (N_10456,N_9320,N_9229);
xnor U10457 (N_10457,N_9489,N_9186);
nor U10458 (N_10458,N_9162,N_9071);
or U10459 (N_10459,N_9110,N_9011);
nor U10460 (N_10460,N_9385,N_9382);
nor U10461 (N_10461,N_9440,N_9230);
or U10462 (N_10462,N_9511,N_9559);
nand U10463 (N_10463,N_9049,N_9703);
and U10464 (N_10464,N_9184,N_9567);
and U10465 (N_10465,N_9088,N_9573);
nor U10466 (N_10466,N_9211,N_9624);
or U10467 (N_10467,N_9160,N_9621);
nor U10468 (N_10468,N_9250,N_9416);
nor U10469 (N_10469,N_9594,N_9730);
and U10470 (N_10470,N_9121,N_9677);
and U10471 (N_10471,N_9445,N_9430);
nand U10472 (N_10472,N_9142,N_9438);
or U10473 (N_10473,N_9397,N_9685);
and U10474 (N_10474,N_9267,N_9398);
xor U10475 (N_10475,N_9128,N_9188);
xor U10476 (N_10476,N_9681,N_9301);
nand U10477 (N_10477,N_9042,N_9695);
nor U10478 (N_10478,N_9590,N_9411);
or U10479 (N_10479,N_9296,N_9172);
nand U10480 (N_10480,N_9129,N_9417);
xnor U10481 (N_10481,N_9221,N_9449);
nor U10482 (N_10482,N_9543,N_9584);
nand U10483 (N_10483,N_9102,N_9628);
nor U10484 (N_10484,N_9724,N_9316);
and U10485 (N_10485,N_9668,N_9366);
or U10486 (N_10486,N_9136,N_9235);
xor U10487 (N_10487,N_9318,N_9230);
nand U10488 (N_10488,N_9307,N_9154);
nor U10489 (N_10489,N_9436,N_9650);
and U10490 (N_10490,N_9137,N_9643);
and U10491 (N_10491,N_9201,N_9554);
nor U10492 (N_10492,N_9183,N_9563);
xnor U10493 (N_10493,N_9647,N_9331);
xnor U10494 (N_10494,N_9463,N_9363);
nand U10495 (N_10495,N_9498,N_9497);
and U10496 (N_10496,N_9627,N_9078);
nor U10497 (N_10497,N_9018,N_9026);
and U10498 (N_10498,N_9458,N_9333);
nor U10499 (N_10499,N_9021,N_9108);
xnor U10500 (N_10500,N_10117,N_9995);
nand U10501 (N_10501,N_9880,N_10337);
or U10502 (N_10502,N_10198,N_9760);
nand U10503 (N_10503,N_10147,N_9978);
nand U10504 (N_10504,N_9953,N_10199);
and U10505 (N_10505,N_10395,N_9772);
nand U10506 (N_10506,N_9860,N_9915);
and U10507 (N_10507,N_9952,N_10392);
xor U10508 (N_10508,N_10153,N_10068);
nand U10509 (N_10509,N_10164,N_10412);
nor U10510 (N_10510,N_9771,N_10225);
nor U10511 (N_10511,N_10282,N_10010);
nand U10512 (N_10512,N_10071,N_10353);
xnor U10513 (N_10513,N_10079,N_9791);
nor U10514 (N_10514,N_10294,N_9938);
nand U10515 (N_10515,N_10108,N_9956);
or U10516 (N_10516,N_10475,N_10341);
nand U10517 (N_10517,N_9873,N_10038);
nand U10518 (N_10518,N_9810,N_10291);
xor U10519 (N_10519,N_10106,N_9750);
xnor U10520 (N_10520,N_10460,N_10192);
nand U10521 (N_10521,N_9993,N_10231);
xnor U10522 (N_10522,N_9814,N_10466);
and U10523 (N_10523,N_9851,N_10271);
nor U10524 (N_10524,N_10154,N_9936);
xor U10525 (N_10525,N_10037,N_10381);
or U10526 (N_10526,N_10358,N_9874);
and U10527 (N_10527,N_9821,N_10495);
xor U10528 (N_10528,N_9804,N_10461);
nand U10529 (N_10529,N_10126,N_10321);
nand U10530 (N_10530,N_10133,N_10411);
or U10531 (N_10531,N_10263,N_9923);
or U10532 (N_10532,N_9913,N_9968);
nor U10533 (N_10533,N_10202,N_10129);
and U10534 (N_10534,N_9783,N_10131);
and U10535 (N_10535,N_10423,N_10367);
nand U10536 (N_10536,N_10484,N_9929);
nand U10537 (N_10537,N_9802,N_10284);
nand U10538 (N_10538,N_10360,N_10141);
xnor U10539 (N_10539,N_9872,N_10030);
or U10540 (N_10540,N_10171,N_9881);
xnor U10541 (N_10541,N_9912,N_10176);
nor U10542 (N_10542,N_9795,N_10174);
and U10543 (N_10543,N_10144,N_10086);
and U10544 (N_10544,N_9835,N_10157);
nor U10545 (N_10545,N_10436,N_10128);
nor U10546 (N_10546,N_9815,N_9755);
nand U10547 (N_10547,N_9752,N_9761);
or U10548 (N_10548,N_10022,N_9972);
nor U10549 (N_10549,N_9803,N_10327);
or U10550 (N_10550,N_10017,N_9800);
nand U10551 (N_10551,N_9957,N_9834);
xor U10552 (N_10552,N_9899,N_10338);
nor U10553 (N_10553,N_10494,N_10309);
nand U10554 (N_10554,N_10318,N_10464);
nor U10555 (N_10555,N_10437,N_9766);
and U10556 (N_10556,N_10322,N_9777);
xnor U10557 (N_10557,N_9924,N_10127);
or U10558 (N_10558,N_10215,N_9914);
and U10559 (N_10559,N_9843,N_9981);
or U10560 (N_10560,N_10113,N_10182);
nor U10561 (N_10561,N_9959,N_10000);
nand U10562 (N_10562,N_10351,N_10339);
and U10563 (N_10563,N_9866,N_10214);
and U10564 (N_10564,N_10384,N_9960);
or U10565 (N_10565,N_9871,N_9986);
nor U10566 (N_10566,N_9909,N_10414);
or U10567 (N_10567,N_9838,N_10472);
or U10568 (N_10568,N_10259,N_9989);
or U10569 (N_10569,N_10146,N_10346);
and U10570 (N_10570,N_10389,N_9976);
or U10571 (N_10571,N_10145,N_9827);
xnor U10572 (N_10572,N_9982,N_10306);
nor U10573 (N_10573,N_9824,N_10021);
nand U10574 (N_10574,N_10344,N_9879);
or U10575 (N_10575,N_10057,N_9862);
nor U10576 (N_10576,N_9831,N_10115);
nand U10577 (N_10577,N_10228,N_10122);
and U10578 (N_10578,N_10029,N_9868);
nand U10579 (N_10579,N_10486,N_10100);
nand U10580 (N_10580,N_9850,N_10201);
and U10581 (N_10581,N_10204,N_10219);
nand U10582 (N_10582,N_10102,N_10480);
or U10583 (N_10583,N_9939,N_10270);
nand U10584 (N_10584,N_10006,N_9798);
xnor U10585 (N_10585,N_10211,N_10380);
xor U10586 (N_10586,N_9935,N_10386);
or U10587 (N_10587,N_10413,N_10250);
xor U10588 (N_10588,N_10462,N_9820);
nand U10589 (N_10589,N_10454,N_10451);
and U10590 (N_10590,N_10487,N_10240);
nand U10591 (N_10591,N_9920,N_10498);
xor U10592 (N_10592,N_9948,N_10123);
or U10593 (N_10593,N_10187,N_9849);
and U10594 (N_10594,N_10433,N_10292);
and U10595 (N_10595,N_10234,N_10378);
nand U10596 (N_10596,N_10355,N_10398);
nand U10597 (N_10597,N_10168,N_9819);
nor U10598 (N_10598,N_9756,N_9758);
or U10599 (N_10599,N_9916,N_10424);
xnor U10600 (N_10600,N_10160,N_10104);
xor U10601 (N_10601,N_10172,N_10312);
and U10602 (N_10602,N_10042,N_10492);
nor U10603 (N_10603,N_10333,N_9779);
and U10604 (N_10604,N_10082,N_10136);
nor U10605 (N_10605,N_9751,N_10459);
nor U10606 (N_10606,N_10098,N_9809);
nand U10607 (N_10607,N_10148,N_9934);
or U10608 (N_10608,N_10298,N_9770);
nor U10609 (N_10609,N_10249,N_10336);
or U10610 (N_10610,N_10237,N_9921);
and U10611 (N_10611,N_10391,N_9994);
nor U10612 (N_10612,N_10425,N_10111);
nand U10613 (N_10613,N_10383,N_10328);
nor U10614 (N_10614,N_9947,N_10223);
nand U10615 (N_10615,N_9896,N_9966);
or U10616 (N_10616,N_10090,N_10279);
nor U10617 (N_10617,N_10257,N_10331);
or U10618 (N_10618,N_10130,N_10458);
xor U10619 (N_10619,N_9759,N_9906);
xor U10620 (N_10620,N_9992,N_9951);
xor U10621 (N_10621,N_10352,N_10499);
and U10622 (N_10622,N_9863,N_9840);
xnor U10623 (N_10623,N_9917,N_10340);
nand U10624 (N_10624,N_10200,N_10216);
and U10625 (N_10625,N_10166,N_9890);
xnor U10626 (N_10626,N_9904,N_10359);
or U10627 (N_10627,N_10177,N_10286);
and U10628 (N_10628,N_10097,N_10422);
nor U10629 (N_10629,N_10114,N_10163);
or U10630 (N_10630,N_10008,N_10138);
nor U10631 (N_10631,N_10046,N_10132);
and U10632 (N_10632,N_10450,N_9886);
or U10633 (N_10633,N_10348,N_10137);
nand U10634 (N_10634,N_10024,N_10072);
nand U10635 (N_10635,N_9757,N_10239);
xnor U10636 (N_10636,N_10262,N_10476);
or U10637 (N_10637,N_10094,N_10264);
xnor U10638 (N_10638,N_10385,N_10307);
or U10639 (N_10639,N_10406,N_10419);
nor U10640 (N_10640,N_10374,N_10434);
nor U10641 (N_10641,N_10335,N_9898);
nand U10642 (N_10642,N_10330,N_10009);
nand U10643 (N_10643,N_10305,N_10236);
or U10644 (N_10644,N_10238,N_10426);
or U10645 (N_10645,N_9839,N_9996);
or U10646 (N_10646,N_10197,N_10015);
nand U10647 (N_10647,N_10295,N_9856);
nand U10648 (N_10648,N_9829,N_9937);
or U10649 (N_10649,N_10405,N_10287);
and U10650 (N_10650,N_10077,N_10449);
or U10651 (N_10651,N_10326,N_9782);
nor U10652 (N_10652,N_10345,N_10053);
nor U10653 (N_10653,N_10039,N_10260);
nand U10654 (N_10654,N_10035,N_10261);
or U10655 (N_10655,N_9786,N_9908);
nor U10656 (N_10656,N_9781,N_10368);
xor U10657 (N_10657,N_10169,N_9979);
nand U10658 (N_10658,N_10455,N_10364);
and U10659 (N_10659,N_9826,N_9894);
nor U10660 (N_10660,N_10315,N_10101);
or U10661 (N_10661,N_9846,N_9907);
nor U10662 (N_10662,N_10440,N_9983);
xor U10663 (N_10663,N_9943,N_10099);
or U10664 (N_10664,N_10296,N_9971);
or U10665 (N_10665,N_10427,N_10350);
nor U10666 (N_10666,N_10470,N_10156);
nand U10667 (N_10667,N_10161,N_10377);
xor U10668 (N_10668,N_10005,N_9778);
or U10669 (N_10669,N_10408,N_10226);
nand U10670 (N_10670,N_10273,N_10203);
and U10671 (N_10671,N_10087,N_10052);
or U10672 (N_10672,N_10444,N_10329);
or U10673 (N_10673,N_10045,N_9776);
nand U10674 (N_10674,N_10034,N_9876);
nand U10675 (N_10675,N_10469,N_10151);
xor U10676 (N_10676,N_10073,N_10059);
nor U10677 (N_10677,N_10076,N_10061);
xor U10678 (N_10678,N_10402,N_10293);
nand U10679 (N_10679,N_10242,N_10445);
xnor U10680 (N_10680,N_10290,N_10212);
and U10681 (N_10681,N_10183,N_10421);
xnor U10682 (N_10682,N_10400,N_10063);
xnor U10683 (N_10683,N_10004,N_10317);
or U10684 (N_10684,N_9892,N_10230);
nor U10685 (N_10685,N_9855,N_9869);
or U10686 (N_10686,N_9964,N_10442);
nor U10687 (N_10687,N_10075,N_10220);
and U10688 (N_10688,N_10447,N_9852);
nor U10689 (N_10689,N_10471,N_10334);
nand U10690 (N_10690,N_9864,N_9784);
or U10691 (N_10691,N_10103,N_9969);
and U10692 (N_10692,N_10342,N_10371);
nand U10693 (N_10693,N_9762,N_10258);
nor U10694 (N_10694,N_10050,N_10185);
nor U10695 (N_10695,N_10430,N_9888);
nor U10696 (N_10696,N_9987,N_10382);
nand U10697 (N_10697,N_9818,N_10049);
xnor U10698 (N_10698,N_9808,N_9997);
nand U10699 (N_10699,N_10483,N_10105);
xor U10700 (N_10700,N_10431,N_9836);
nor U10701 (N_10701,N_10221,N_10366);
nor U10702 (N_10702,N_10404,N_10417);
nand U10703 (N_10703,N_10224,N_10055);
and U10704 (N_10704,N_9807,N_10323);
or U10705 (N_10705,N_10121,N_10418);
and U10706 (N_10706,N_9897,N_10474);
and U10707 (N_10707,N_10116,N_10388);
or U10708 (N_10708,N_9999,N_10477);
or U10709 (N_10709,N_9822,N_10482);
nand U10710 (N_10710,N_10403,N_9805);
and U10711 (N_10711,N_10248,N_9845);
and U10712 (N_10712,N_10362,N_10142);
or U10713 (N_10713,N_10452,N_10416);
and U10714 (N_10714,N_9985,N_10302);
xor U10715 (N_10715,N_9844,N_10194);
or U10716 (N_10716,N_10020,N_9980);
or U10717 (N_10717,N_10301,N_9789);
nor U10718 (N_10718,N_9865,N_10319);
xor U10719 (N_10719,N_9990,N_10170);
nor U10720 (N_10720,N_10397,N_10372);
nor U10721 (N_10721,N_10051,N_10297);
xor U10722 (N_10722,N_10218,N_10195);
nor U10723 (N_10723,N_10396,N_9790);
nand U10724 (N_10724,N_10095,N_9891);
and U10725 (N_10725,N_10446,N_10375);
and U10726 (N_10726,N_9945,N_9903);
nand U10727 (N_10727,N_10489,N_10308);
or U10728 (N_10728,N_10190,N_10083);
or U10729 (N_10729,N_10158,N_9785);
nor U10730 (N_10730,N_10457,N_9882);
or U10731 (N_10731,N_10180,N_10031);
or U10732 (N_10732,N_9988,N_10274);
nor U10733 (N_10733,N_9801,N_10265);
nor U10734 (N_10734,N_10361,N_10186);
xnor U10735 (N_10735,N_9788,N_10088);
or U10736 (N_10736,N_9753,N_10175);
nand U10737 (N_10737,N_9926,N_10268);
nor U10738 (N_10738,N_10018,N_10435);
xor U10739 (N_10739,N_9774,N_9870);
nand U10740 (N_10740,N_9875,N_10438);
or U10741 (N_10741,N_10165,N_10140);
nor U10742 (N_10742,N_10189,N_10109);
and U10743 (N_10743,N_9911,N_9857);
nand U10744 (N_10744,N_10316,N_10266);
xor U10745 (N_10745,N_10139,N_10056);
xnor U10746 (N_10746,N_10354,N_10379);
xnor U10747 (N_10747,N_9933,N_10032);
xor U10748 (N_10748,N_10409,N_10014);
nor U10749 (N_10749,N_10357,N_10428);
or U10750 (N_10750,N_10179,N_9963);
nor U10751 (N_10751,N_10304,N_10481);
nor U10752 (N_10752,N_9885,N_9763);
xor U10753 (N_10753,N_10300,N_10205);
nor U10754 (N_10754,N_10178,N_10181);
xor U10755 (N_10755,N_9787,N_10096);
nand U10756 (N_10756,N_10119,N_10019);
nor U10757 (N_10757,N_10283,N_9949);
xor U10758 (N_10758,N_10047,N_10001);
xor U10759 (N_10759,N_10276,N_10048);
xnor U10760 (N_10760,N_10227,N_10478);
or U10761 (N_10761,N_10497,N_9830);
and U10762 (N_10762,N_9806,N_9837);
or U10763 (N_10763,N_10058,N_10496);
and U10764 (N_10764,N_9883,N_10089);
nand U10765 (N_10765,N_10280,N_10155);
xor U10766 (N_10766,N_10493,N_10347);
and U10767 (N_10767,N_10325,N_9984);
or U10768 (N_10768,N_10324,N_10107);
and U10769 (N_10769,N_10043,N_9941);
nor U10770 (N_10770,N_10093,N_10085);
and U10771 (N_10771,N_10252,N_10432);
nor U10772 (N_10772,N_10376,N_10363);
and U10773 (N_10773,N_9925,N_9975);
nor U10774 (N_10774,N_10209,N_9901);
or U10775 (N_10775,N_10288,N_10251);
or U10776 (N_10776,N_10003,N_10028);
nor U10777 (N_10777,N_9833,N_9887);
nand U10778 (N_10778,N_9965,N_10054);
and U10779 (N_10779,N_9967,N_9946);
or U10780 (N_10780,N_10448,N_10060);
xor U10781 (N_10781,N_9977,N_10278);
nor U10782 (N_10782,N_9841,N_9793);
xor U10783 (N_10783,N_10429,N_9816);
xor U10784 (N_10784,N_10023,N_9754);
and U10785 (N_10785,N_9961,N_9828);
and U10786 (N_10786,N_9853,N_10255);
and U10787 (N_10787,N_9765,N_9811);
nor U10788 (N_10788,N_10150,N_9813);
xnor U10789 (N_10789,N_9942,N_9930);
xor U10790 (N_10790,N_9944,N_9842);
nand U10791 (N_10791,N_10012,N_10233);
nor U10792 (N_10792,N_10162,N_10208);
or U10793 (N_10793,N_10026,N_10479);
and U10794 (N_10794,N_10245,N_10369);
nor U10795 (N_10795,N_10036,N_10394);
nor U10796 (N_10796,N_10210,N_10453);
or U10797 (N_10797,N_10149,N_10465);
nor U10798 (N_10798,N_9825,N_9927);
xnor U10799 (N_10799,N_9858,N_10415);
nand U10800 (N_10800,N_9867,N_10407);
nand U10801 (N_10801,N_10332,N_10491);
xor U10802 (N_10802,N_10488,N_10256);
and U10803 (N_10803,N_10112,N_9958);
or U10804 (N_10804,N_9991,N_10393);
nand U10805 (N_10805,N_10473,N_9922);
or U10806 (N_10806,N_9764,N_10490);
nand U10807 (N_10807,N_10011,N_10485);
nor U10808 (N_10808,N_10246,N_9773);
nand U10809 (N_10809,N_10311,N_10235);
and U10810 (N_10810,N_10184,N_9796);
and U10811 (N_10811,N_10196,N_10084);
nand U10812 (N_10812,N_9767,N_10081);
nor U10813 (N_10813,N_10091,N_10222);
xor U10814 (N_10814,N_10349,N_10420);
xor U10815 (N_10815,N_10247,N_10269);
or U10816 (N_10816,N_10213,N_10410);
xor U10817 (N_10817,N_10159,N_10467);
nand U10818 (N_10818,N_10066,N_10027);
nand U10819 (N_10819,N_10092,N_10070);
xor U10820 (N_10820,N_10399,N_10025);
nor U10821 (N_10821,N_9905,N_10310);
nand U10822 (N_10822,N_10356,N_9998);
nand U10823 (N_10823,N_9950,N_9902);
nor U10824 (N_10824,N_10007,N_9794);
and U10825 (N_10825,N_10401,N_9884);
or U10826 (N_10826,N_9895,N_10033);
and U10827 (N_10827,N_10232,N_9799);
and U10828 (N_10828,N_10002,N_10253);
nor U10829 (N_10829,N_10013,N_10229);
nor U10830 (N_10830,N_9780,N_9832);
or U10831 (N_10831,N_9878,N_10370);
nor U10832 (N_10832,N_10143,N_10152);
nor U10833 (N_10833,N_10277,N_10134);
or U10834 (N_10834,N_10343,N_10016);
nor U10835 (N_10835,N_9940,N_10267);
and U10836 (N_10836,N_10365,N_10303);
and U10837 (N_10837,N_10167,N_10439);
nor U10838 (N_10838,N_10217,N_10468);
or U10839 (N_10839,N_9928,N_10118);
or U10840 (N_10840,N_9955,N_9859);
and U10841 (N_10841,N_9877,N_9970);
nor U10842 (N_10842,N_10275,N_10040);
nand U10843 (N_10843,N_10390,N_9974);
or U10844 (N_10844,N_10206,N_9900);
nor U10845 (N_10845,N_10173,N_10244);
or U10846 (N_10846,N_10067,N_10373);
and U10847 (N_10847,N_10243,N_10080);
or U10848 (N_10848,N_9797,N_10044);
or U10849 (N_10849,N_10314,N_10188);
or U10850 (N_10850,N_9823,N_10441);
and U10851 (N_10851,N_10387,N_9910);
or U10852 (N_10852,N_9812,N_10078);
and U10853 (N_10853,N_10041,N_10289);
xor U10854 (N_10854,N_10285,N_9954);
or U10855 (N_10855,N_10241,N_9962);
and U10856 (N_10856,N_9932,N_10124);
or U10857 (N_10857,N_10125,N_9775);
nor U10858 (N_10858,N_10320,N_9817);
or U10859 (N_10859,N_9931,N_10065);
nand U10860 (N_10860,N_10463,N_9889);
nor U10861 (N_10861,N_9973,N_10062);
and U10862 (N_10862,N_10281,N_9847);
xor U10863 (N_10863,N_10110,N_10193);
xor U10864 (N_10864,N_10120,N_9854);
nand U10865 (N_10865,N_10456,N_9768);
and U10866 (N_10866,N_10064,N_10254);
nand U10867 (N_10867,N_10135,N_10191);
xnor U10868 (N_10868,N_9848,N_10069);
nand U10869 (N_10869,N_9893,N_10299);
nor U10870 (N_10870,N_10272,N_9769);
and U10871 (N_10871,N_9792,N_9918);
xor U10872 (N_10872,N_10207,N_10313);
nand U10873 (N_10873,N_9861,N_9919);
nor U10874 (N_10874,N_10074,N_10443);
xnor U10875 (N_10875,N_9889,N_10253);
and U10876 (N_10876,N_10307,N_9962);
and U10877 (N_10877,N_10142,N_10491);
and U10878 (N_10878,N_9838,N_9952);
and U10879 (N_10879,N_9954,N_10017);
nand U10880 (N_10880,N_10303,N_9797);
xnor U10881 (N_10881,N_10475,N_10323);
nor U10882 (N_10882,N_10473,N_10468);
nand U10883 (N_10883,N_10336,N_10264);
or U10884 (N_10884,N_10376,N_10250);
nor U10885 (N_10885,N_9753,N_9886);
nand U10886 (N_10886,N_10074,N_10255);
nand U10887 (N_10887,N_10174,N_10020);
and U10888 (N_10888,N_10415,N_9778);
or U10889 (N_10889,N_9937,N_10209);
xnor U10890 (N_10890,N_9995,N_10329);
and U10891 (N_10891,N_9928,N_10400);
or U10892 (N_10892,N_10124,N_10240);
and U10893 (N_10893,N_9852,N_10179);
xnor U10894 (N_10894,N_10153,N_9786);
or U10895 (N_10895,N_10483,N_9938);
and U10896 (N_10896,N_10191,N_10192);
xnor U10897 (N_10897,N_10064,N_10442);
nor U10898 (N_10898,N_10445,N_10383);
xnor U10899 (N_10899,N_9924,N_10092);
nand U10900 (N_10900,N_10172,N_9815);
xnor U10901 (N_10901,N_10297,N_10195);
and U10902 (N_10902,N_10047,N_10245);
or U10903 (N_10903,N_9836,N_10363);
nand U10904 (N_10904,N_9771,N_10288);
and U10905 (N_10905,N_10483,N_9751);
xor U10906 (N_10906,N_10300,N_9960);
and U10907 (N_10907,N_10385,N_9829);
xor U10908 (N_10908,N_10282,N_10293);
xnor U10909 (N_10909,N_9874,N_10197);
or U10910 (N_10910,N_9938,N_10393);
and U10911 (N_10911,N_10374,N_10008);
nor U10912 (N_10912,N_10434,N_10085);
nor U10913 (N_10913,N_9819,N_10064);
and U10914 (N_10914,N_10162,N_10158);
and U10915 (N_10915,N_10372,N_10203);
or U10916 (N_10916,N_10406,N_10342);
and U10917 (N_10917,N_10041,N_10234);
nor U10918 (N_10918,N_10487,N_9878);
nand U10919 (N_10919,N_9933,N_10106);
xnor U10920 (N_10920,N_9841,N_9883);
xnor U10921 (N_10921,N_10247,N_9939);
nand U10922 (N_10922,N_10128,N_9905);
nor U10923 (N_10923,N_10009,N_9936);
nand U10924 (N_10924,N_10497,N_9955);
nand U10925 (N_10925,N_9902,N_10490);
nand U10926 (N_10926,N_10076,N_10242);
nor U10927 (N_10927,N_9846,N_9884);
and U10928 (N_10928,N_9888,N_10453);
nor U10929 (N_10929,N_10024,N_10354);
or U10930 (N_10930,N_9963,N_9868);
xnor U10931 (N_10931,N_10493,N_10490);
nor U10932 (N_10932,N_10365,N_9884);
or U10933 (N_10933,N_10213,N_10067);
nand U10934 (N_10934,N_10030,N_9906);
and U10935 (N_10935,N_9766,N_10184);
or U10936 (N_10936,N_10249,N_10219);
nor U10937 (N_10937,N_10429,N_10255);
nor U10938 (N_10938,N_10362,N_10100);
xor U10939 (N_10939,N_10417,N_10180);
and U10940 (N_10940,N_9885,N_10283);
nor U10941 (N_10941,N_10449,N_10441);
or U10942 (N_10942,N_10020,N_9958);
nor U10943 (N_10943,N_10254,N_10147);
or U10944 (N_10944,N_10395,N_9912);
nor U10945 (N_10945,N_9903,N_10070);
xor U10946 (N_10946,N_10496,N_9966);
xnor U10947 (N_10947,N_10499,N_10390);
and U10948 (N_10948,N_10005,N_10078);
and U10949 (N_10949,N_10101,N_10463);
or U10950 (N_10950,N_10341,N_10480);
or U10951 (N_10951,N_10406,N_10001);
xor U10952 (N_10952,N_9994,N_10155);
nor U10953 (N_10953,N_9829,N_10239);
or U10954 (N_10954,N_10333,N_10102);
or U10955 (N_10955,N_10159,N_9798);
xnor U10956 (N_10956,N_10485,N_9893);
nor U10957 (N_10957,N_10168,N_10205);
xor U10958 (N_10958,N_10308,N_10036);
nor U10959 (N_10959,N_10349,N_10025);
nor U10960 (N_10960,N_10217,N_9986);
xnor U10961 (N_10961,N_10146,N_10278);
or U10962 (N_10962,N_10095,N_10264);
xor U10963 (N_10963,N_10004,N_9945);
nand U10964 (N_10964,N_9949,N_10450);
xnor U10965 (N_10965,N_10014,N_10398);
nand U10966 (N_10966,N_10206,N_10285);
and U10967 (N_10967,N_10138,N_10100);
nand U10968 (N_10968,N_9866,N_9790);
nand U10969 (N_10969,N_9919,N_10249);
nor U10970 (N_10970,N_10014,N_10141);
xnor U10971 (N_10971,N_10161,N_10007);
nand U10972 (N_10972,N_10404,N_10282);
and U10973 (N_10973,N_9752,N_9930);
or U10974 (N_10974,N_10069,N_9808);
or U10975 (N_10975,N_9968,N_10139);
and U10976 (N_10976,N_10049,N_10363);
nand U10977 (N_10977,N_9793,N_10384);
nand U10978 (N_10978,N_10022,N_9979);
and U10979 (N_10979,N_10083,N_10413);
nor U10980 (N_10980,N_10308,N_10062);
xnor U10981 (N_10981,N_9969,N_10266);
and U10982 (N_10982,N_10076,N_10405);
and U10983 (N_10983,N_9846,N_10470);
nor U10984 (N_10984,N_9833,N_9789);
and U10985 (N_10985,N_10263,N_10227);
nor U10986 (N_10986,N_10081,N_9909);
xor U10987 (N_10987,N_10037,N_9875);
nand U10988 (N_10988,N_10158,N_10026);
or U10989 (N_10989,N_10362,N_10484);
xor U10990 (N_10990,N_10321,N_10471);
and U10991 (N_10991,N_9932,N_10002);
and U10992 (N_10992,N_10230,N_10010);
or U10993 (N_10993,N_10129,N_10425);
nor U10994 (N_10994,N_9971,N_10450);
or U10995 (N_10995,N_10169,N_10477);
nand U10996 (N_10996,N_9825,N_10099);
and U10997 (N_10997,N_10228,N_10291);
nand U10998 (N_10998,N_10215,N_10441);
and U10999 (N_10999,N_10407,N_10153);
and U11000 (N_11000,N_9961,N_10113);
nand U11001 (N_11001,N_9809,N_10499);
nor U11002 (N_11002,N_10349,N_9800);
or U11003 (N_11003,N_10163,N_10432);
nand U11004 (N_11004,N_10321,N_10342);
xor U11005 (N_11005,N_10346,N_10019);
and U11006 (N_11006,N_10395,N_9862);
nor U11007 (N_11007,N_10166,N_9807);
and U11008 (N_11008,N_9849,N_10160);
or U11009 (N_11009,N_9996,N_10444);
xnor U11010 (N_11010,N_10051,N_9952);
and U11011 (N_11011,N_10362,N_10297);
nand U11012 (N_11012,N_10188,N_9839);
nor U11013 (N_11013,N_10454,N_9954);
or U11014 (N_11014,N_9988,N_10429);
xnor U11015 (N_11015,N_10265,N_10230);
and U11016 (N_11016,N_9805,N_10195);
nor U11017 (N_11017,N_9835,N_10408);
nand U11018 (N_11018,N_10331,N_9796);
nand U11019 (N_11019,N_10072,N_10248);
nand U11020 (N_11020,N_10026,N_10183);
xnor U11021 (N_11021,N_9925,N_10148);
nand U11022 (N_11022,N_10146,N_10337);
or U11023 (N_11023,N_10070,N_10085);
nand U11024 (N_11024,N_10145,N_9935);
and U11025 (N_11025,N_9795,N_10361);
nand U11026 (N_11026,N_10011,N_9844);
nand U11027 (N_11027,N_10036,N_9974);
and U11028 (N_11028,N_10026,N_9750);
nor U11029 (N_11029,N_10444,N_10109);
or U11030 (N_11030,N_10252,N_9909);
nor U11031 (N_11031,N_10438,N_10297);
nand U11032 (N_11032,N_10372,N_10300);
or U11033 (N_11033,N_10488,N_9929);
nand U11034 (N_11034,N_10338,N_10082);
or U11035 (N_11035,N_10341,N_10111);
nand U11036 (N_11036,N_10475,N_10073);
nand U11037 (N_11037,N_10095,N_10482);
and U11038 (N_11038,N_10073,N_9868);
or U11039 (N_11039,N_9803,N_10445);
xor U11040 (N_11040,N_9882,N_9879);
and U11041 (N_11041,N_10383,N_9756);
and U11042 (N_11042,N_9887,N_9840);
nor U11043 (N_11043,N_9962,N_9993);
nor U11044 (N_11044,N_10092,N_10408);
nand U11045 (N_11045,N_9939,N_9948);
nand U11046 (N_11046,N_10410,N_10431);
and U11047 (N_11047,N_9954,N_10299);
and U11048 (N_11048,N_9777,N_10416);
xnor U11049 (N_11049,N_10391,N_10277);
nand U11050 (N_11050,N_10220,N_10215);
xor U11051 (N_11051,N_10228,N_10287);
nand U11052 (N_11052,N_10162,N_10475);
and U11053 (N_11053,N_10386,N_10341);
or U11054 (N_11054,N_10281,N_10260);
nor U11055 (N_11055,N_10120,N_10176);
nand U11056 (N_11056,N_9974,N_9959);
and U11057 (N_11057,N_9999,N_10007);
or U11058 (N_11058,N_10219,N_10089);
nor U11059 (N_11059,N_9861,N_9763);
or U11060 (N_11060,N_9909,N_9961);
xor U11061 (N_11061,N_10118,N_9957);
nor U11062 (N_11062,N_10030,N_10118);
or U11063 (N_11063,N_10039,N_9978);
nand U11064 (N_11064,N_10264,N_9938);
nand U11065 (N_11065,N_10335,N_10061);
nor U11066 (N_11066,N_10180,N_10474);
and U11067 (N_11067,N_10035,N_10170);
nand U11068 (N_11068,N_9983,N_9893);
nand U11069 (N_11069,N_9931,N_9761);
nand U11070 (N_11070,N_9832,N_9973);
xor U11071 (N_11071,N_9825,N_10113);
and U11072 (N_11072,N_10160,N_9843);
nand U11073 (N_11073,N_10243,N_10094);
and U11074 (N_11074,N_10367,N_10263);
nor U11075 (N_11075,N_10447,N_9778);
nor U11076 (N_11076,N_10177,N_10030);
nor U11077 (N_11077,N_9867,N_9895);
or U11078 (N_11078,N_10348,N_10370);
xnor U11079 (N_11079,N_10202,N_9943);
or U11080 (N_11080,N_10214,N_10266);
and U11081 (N_11081,N_9965,N_9776);
nand U11082 (N_11082,N_10409,N_10015);
nor U11083 (N_11083,N_9785,N_10109);
xor U11084 (N_11084,N_10186,N_10003);
nand U11085 (N_11085,N_10138,N_9829);
nand U11086 (N_11086,N_9798,N_10146);
xor U11087 (N_11087,N_10338,N_9774);
xor U11088 (N_11088,N_9847,N_9856);
and U11089 (N_11089,N_10282,N_10465);
and U11090 (N_11090,N_9797,N_10091);
xnor U11091 (N_11091,N_10395,N_10036);
xnor U11092 (N_11092,N_9828,N_10194);
and U11093 (N_11093,N_9776,N_9940);
nand U11094 (N_11094,N_9779,N_10097);
nor U11095 (N_11095,N_10150,N_10335);
and U11096 (N_11096,N_10023,N_9931);
nor U11097 (N_11097,N_9941,N_10077);
nor U11098 (N_11098,N_9951,N_9812);
nor U11099 (N_11099,N_10013,N_10382);
nor U11100 (N_11100,N_10059,N_10286);
nand U11101 (N_11101,N_9836,N_10149);
nor U11102 (N_11102,N_10110,N_10078);
nor U11103 (N_11103,N_10411,N_10463);
and U11104 (N_11104,N_9921,N_10007);
xor U11105 (N_11105,N_9897,N_10398);
and U11106 (N_11106,N_10275,N_10087);
and U11107 (N_11107,N_10404,N_10434);
or U11108 (N_11108,N_9903,N_10065);
nand U11109 (N_11109,N_10133,N_10318);
and U11110 (N_11110,N_9892,N_10333);
nor U11111 (N_11111,N_10277,N_10303);
nand U11112 (N_11112,N_9881,N_9826);
or U11113 (N_11113,N_10188,N_9946);
nor U11114 (N_11114,N_10107,N_10100);
nor U11115 (N_11115,N_9876,N_9864);
or U11116 (N_11116,N_10464,N_10478);
nand U11117 (N_11117,N_10004,N_9849);
nor U11118 (N_11118,N_9785,N_10312);
xor U11119 (N_11119,N_10242,N_10133);
nand U11120 (N_11120,N_10071,N_10006);
and U11121 (N_11121,N_10094,N_10481);
and U11122 (N_11122,N_10142,N_10236);
nand U11123 (N_11123,N_10343,N_9844);
nor U11124 (N_11124,N_10257,N_10199);
xnor U11125 (N_11125,N_10472,N_10238);
nand U11126 (N_11126,N_9895,N_10477);
nor U11127 (N_11127,N_9989,N_9789);
or U11128 (N_11128,N_9768,N_10380);
xnor U11129 (N_11129,N_10093,N_9813);
xnor U11130 (N_11130,N_9857,N_10033);
and U11131 (N_11131,N_10209,N_10472);
and U11132 (N_11132,N_9808,N_9917);
or U11133 (N_11133,N_9894,N_10043);
nor U11134 (N_11134,N_9877,N_10225);
and U11135 (N_11135,N_9882,N_9954);
or U11136 (N_11136,N_10417,N_10401);
nor U11137 (N_11137,N_9854,N_10440);
and U11138 (N_11138,N_10207,N_9951);
and U11139 (N_11139,N_9965,N_10288);
and U11140 (N_11140,N_9763,N_10471);
xnor U11141 (N_11141,N_9951,N_10080);
nand U11142 (N_11142,N_10055,N_10022);
and U11143 (N_11143,N_10048,N_10280);
nor U11144 (N_11144,N_9815,N_9850);
nand U11145 (N_11145,N_9778,N_10101);
or U11146 (N_11146,N_10015,N_10007);
or U11147 (N_11147,N_10432,N_9962);
nor U11148 (N_11148,N_10479,N_10085);
nor U11149 (N_11149,N_9860,N_10292);
and U11150 (N_11150,N_9971,N_9769);
nor U11151 (N_11151,N_10376,N_9917);
xor U11152 (N_11152,N_10071,N_9799);
nor U11153 (N_11153,N_10106,N_10225);
or U11154 (N_11154,N_10169,N_10226);
nand U11155 (N_11155,N_9906,N_9754);
and U11156 (N_11156,N_10113,N_10255);
nor U11157 (N_11157,N_9796,N_10378);
xnor U11158 (N_11158,N_10210,N_10062);
xor U11159 (N_11159,N_10444,N_10308);
or U11160 (N_11160,N_9958,N_10485);
nand U11161 (N_11161,N_10344,N_10008);
and U11162 (N_11162,N_10084,N_10488);
xnor U11163 (N_11163,N_9886,N_10063);
or U11164 (N_11164,N_10289,N_9799);
nand U11165 (N_11165,N_10108,N_10181);
or U11166 (N_11166,N_9751,N_10144);
or U11167 (N_11167,N_10480,N_9901);
or U11168 (N_11168,N_10412,N_10102);
nand U11169 (N_11169,N_10015,N_10133);
nand U11170 (N_11170,N_10415,N_9842);
or U11171 (N_11171,N_10074,N_10115);
nand U11172 (N_11172,N_10033,N_10269);
and U11173 (N_11173,N_10358,N_10324);
xor U11174 (N_11174,N_9872,N_9882);
xnor U11175 (N_11175,N_10197,N_10042);
nand U11176 (N_11176,N_10085,N_10030);
nor U11177 (N_11177,N_10246,N_10477);
nand U11178 (N_11178,N_10385,N_9771);
nand U11179 (N_11179,N_9932,N_10256);
and U11180 (N_11180,N_9969,N_9953);
xor U11181 (N_11181,N_9851,N_10027);
nor U11182 (N_11182,N_10261,N_10402);
and U11183 (N_11183,N_10194,N_9826);
or U11184 (N_11184,N_9961,N_10201);
xor U11185 (N_11185,N_10160,N_10116);
and U11186 (N_11186,N_9863,N_9759);
or U11187 (N_11187,N_10370,N_10170);
and U11188 (N_11188,N_9764,N_10080);
or U11189 (N_11189,N_10337,N_10336);
xnor U11190 (N_11190,N_10437,N_10151);
nand U11191 (N_11191,N_10266,N_10475);
nor U11192 (N_11192,N_9782,N_9843);
nand U11193 (N_11193,N_10258,N_10035);
nor U11194 (N_11194,N_9884,N_10446);
and U11195 (N_11195,N_10218,N_10333);
or U11196 (N_11196,N_9802,N_9760);
or U11197 (N_11197,N_10385,N_10199);
nor U11198 (N_11198,N_10391,N_9753);
and U11199 (N_11199,N_10181,N_10372);
nor U11200 (N_11200,N_9940,N_10349);
or U11201 (N_11201,N_10392,N_10213);
or U11202 (N_11202,N_10426,N_10188);
or U11203 (N_11203,N_10093,N_9939);
nor U11204 (N_11204,N_9915,N_9898);
or U11205 (N_11205,N_10230,N_9960);
nor U11206 (N_11206,N_10000,N_10239);
nor U11207 (N_11207,N_10170,N_10104);
or U11208 (N_11208,N_10449,N_10257);
and U11209 (N_11209,N_10412,N_9761);
nand U11210 (N_11210,N_9896,N_10284);
xor U11211 (N_11211,N_10484,N_10183);
nand U11212 (N_11212,N_9939,N_9754);
xnor U11213 (N_11213,N_10121,N_10011);
nor U11214 (N_11214,N_10457,N_10126);
nand U11215 (N_11215,N_10005,N_9834);
nand U11216 (N_11216,N_10181,N_10358);
nor U11217 (N_11217,N_10081,N_9895);
and U11218 (N_11218,N_10286,N_10110);
nand U11219 (N_11219,N_10027,N_10185);
and U11220 (N_11220,N_10468,N_10070);
and U11221 (N_11221,N_9892,N_10332);
nand U11222 (N_11222,N_9990,N_10029);
xor U11223 (N_11223,N_10108,N_9992);
or U11224 (N_11224,N_10370,N_10428);
nand U11225 (N_11225,N_10095,N_10365);
nor U11226 (N_11226,N_10106,N_9906);
or U11227 (N_11227,N_10247,N_9949);
xor U11228 (N_11228,N_10035,N_10234);
and U11229 (N_11229,N_10211,N_10326);
nand U11230 (N_11230,N_10225,N_9970);
nor U11231 (N_11231,N_9870,N_10384);
nand U11232 (N_11232,N_10061,N_10085);
nor U11233 (N_11233,N_10309,N_10111);
or U11234 (N_11234,N_10054,N_10140);
and U11235 (N_11235,N_10217,N_10330);
or U11236 (N_11236,N_9999,N_10361);
nor U11237 (N_11237,N_10024,N_10086);
and U11238 (N_11238,N_10006,N_9885);
nand U11239 (N_11239,N_10134,N_10202);
nor U11240 (N_11240,N_10496,N_10195);
and U11241 (N_11241,N_10483,N_9789);
nand U11242 (N_11242,N_10312,N_10004);
and U11243 (N_11243,N_10259,N_9750);
or U11244 (N_11244,N_10132,N_10175);
nand U11245 (N_11245,N_10006,N_9860);
and U11246 (N_11246,N_9931,N_10315);
nor U11247 (N_11247,N_9857,N_10250);
xor U11248 (N_11248,N_10390,N_10056);
nand U11249 (N_11249,N_10418,N_10303);
nor U11250 (N_11250,N_10677,N_10765);
xnor U11251 (N_11251,N_10894,N_10833);
nand U11252 (N_11252,N_10545,N_10718);
nor U11253 (N_11253,N_11090,N_10671);
and U11254 (N_11254,N_10883,N_10820);
nor U11255 (N_11255,N_10739,N_10508);
or U11256 (N_11256,N_11100,N_11223);
nor U11257 (N_11257,N_10547,N_11075);
and U11258 (N_11258,N_11246,N_10890);
nor U11259 (N_11259,N_10683,N_10904);
or U11260 (N_11260,N_11077,N_11050);
xor U11261 (N_11261,N_10663,N_10939);
nand U11262 (N_11262,N_10875,N_10798);
nand U11263 (N_11263,N_10744,N_10692);
or U11264 (N_11264,N_11024,N_11093);
and U11265 (N_11265,N_10937,N_10988);
nor U11266 (N_11266,N_11056,N_10566);
xor U11267 (N_11267,N_10582,N_11009);
and U11268 (N_11268,N_10655,N_10747);
nand U11269 (N_11269,N_10788,N_11025);
xor U11270 (N_11270,N_11207,N_10579);
and U11271 (N_11271,N_10843,N_11117);
nor U11272 (N_11272,N_10598,N_11082);
and U11273 (N_11273,N_10910,N_10604);
xor U11274 (N_11274,N_10537,N_11163);
nor U11275 (N_11275,N_10501,N_11191);
nor U11276 (N_11276,N_10999,N_11181);
nor U11277 (N_11277,N_10821,N_11079);
xor U11278 (N_11278,N_10926,N_10803);
nor U11279 (N_11279,N_10854,N_11130);
and U11280 (N_11280,N_11213,N_10542);
nor U11281 (N_11281,N_11195,N_10993);
nand U11282 (N_11282,N_10913,N_10757);
and U11283 (N_11283,N_10578,N_10963);
nor U11284 (N_11284,N_10981,N_10942);
xnor U11285 (N_11285,N_10546,N_11189);
xnor U11286 (N_11286,N_11027,N_10672);
xor U11287 (N_11287,N_10940,N_10530);
or U11288 (N_11288,N_11046,N_10882);
or U11289 (N_11289,N_11132,N_11118);
xnor U11290 (N_11290,N_11186,N_11228);
and U11291 (N_11291,N_10505,N_11164);
nor U11292 (N_11292,N_11111,N_11206);
or U11293 (N_11293,N_11174,N_10896);
and U11294 (N_11294,N_10580,N_11198);
xnor U11295 (N_11295,N_10748,N_10838);
and U11296 (N_11296,N_10657,N_11249);
or U11297 (N_11297,N_10811,N_11108);
xnor U11298 (N_11298,N_10727,N_11070);
or U11299 (N_11299,N_11154,N_10835);
and U11300 (N_11300,N_11088,N_11052);
and U11301 (N_11301,N_10893,N_11190);
or U11302 (N_11302,N_10573,N_10664);
xnor U11303 (N_11303,N_10624,N_10852);
or U11304 (N_11304,N_10526,N_10769);
nand U11305 (N_11305,N_11156,N_11146);
and U11306 (N_11306,N_11153,N_10707);
nand U11307 (N_11307,N_10889,N_10538);
or U11308 (N_11308,N_10534,N_10916);
nor U11309 (N_11309,N_10515,N_10620);
nand U11310 (N_11310,N_10575,N_10878);
nand U11311 (N_11311,N_11109,N_11140);
xnor U11312 (N_11312,N_10698,N_10553);
nor U11313 (N_11313,N_10613,N_10502);
and U11314 (N_11314,N_10584,N_11067);
xor U11315 (N_11315,N_11044,N_10715);
nand U11316 (N_11316,N_10702,N_10522);
and U11317 (N_11317,N_11201,N_10750);
nand U11318 (N_11318,N_10592,N_10531);
xor U11319 (N_11319,N_10679,N_11063);
and U11320 (N_11320,N_10756,N_10927);
xor U11321 (N_11321,N_11105,N_11176);
and U11322 (N_11322,N_10549,N_11107);
nand U11323 (N_11323,N_10709,N_11203);
nand U11324 (N_11324,N_11101,N_11241);
nor U11325 (N_11325,N_10642,N_10654);
nor U11326 (N_11326,N_10895,N_11102);
nand U11327 (N_11327,N_10749,N_11012);
or U11328 (N_11328,N_11248,N_10902);
or U11329 (N_11329,N_11196,N_11006);
nand U11330 (N_11330,N_10851,N_11216);
and U11331 (N_11331,N_10638,N_11084);
and U11332 (N_11332,N_10569,N_11187);
or U11333 (N_11333,N_10631,N_10858);
nand U11334 (N_11334,N_10636,N_10509);
xnor U11335 (N_11335,N_11225,N_10724);
nand U11336 (N_11336,N_10831,N_11169);
nor U11337 (N_11337,N_11208,N_11222);
nor U11338 (N_11338,N_11162,N_10876);
nor U11339 (N_11339,N_10871,N_10797);
xnor U11340 (N_11340,N_11110,N_10911);
or U11341 (N_11341,N_11112,N_11144);
nor U11342 (N_11342,N_10690,N_11188);
nand U11343 (N_11343,N_10703,N_10759);
and U11344 (N_11344,N_10958,N_10775);
and U11345 (N_11345,N_11094,N_11014);
nand U11346 (N_11346,N_10887,N_10816);
or U11347 (N_11347,N_11098,N_10639);
or U11348 (N_11348,N_10565,N_10799);
and U11349 (N_11349,N_11182,N_10610);
nor U11350 (N_11350,N_10694,N_11149);
and U11351 (N_11351,N_11022,N_10825);
xor U11352 (N_11352,N_10609,N_11097);
xor U11353 (N_11353,N_11114,N_10667);
nand U11354 (N_11354,N_10752,N_10730);
nor U11355 (N_11355,N_10983,N_10539);
xor U11356 (N_11356,N_10777,N_10784);
nor U11357 (N_11357,N_10527,N_10929);
xnor U11358 (N_11358,N_10706,N_10771);
nand U11359 (N_11359,N_10746,N_10701);
or U11360 (N_11360,N_10848,N_10712);
xor U11361 (N_11361,N_11010,N_10994);
or U11362 (N_11362,N_10614,N_10836);
nor U11363 (N_11363,N_10812,N_11037);
xor U11364 (N_11364,N_11124,N_10961);
and U11365 (N_11365,N_10901,N_10984);
or U11366 (N_11366,N_11159,N_11120);
nor U11367 (N_11367,N_10517,N_11166);
or U11368 (N_11368,N_11167,N_10572);
or U11369 (N_11369,N_10837,N_10951);
and U11370 (N_11370,N_10947,N_10523);
and U11371 (N_11371,N_10800,N_11237);
and U11372 (N_11372,N_11038,N_10669);
and U11373 (N_11373,N_10529,N_10753);
and U11374 (N_11374,N_11217,N_11123);
and U11375 (N_11375,N_11180,N_10990);
or U11376 (N_11376,N_10814,N_10968);
nor U11377 (N_11377,N_10595,N_10924);
nand U11378 (N_11378,N_10934,N_10783);
or U11379 (N_11379,N_10818,N_11071);
nand U11380 (N_11380,N_10944,N_10810);
and U11381 (N_11381,N_10932,N_10596);
xor U11382 (N_11382,N_11205,N_10869);
nor U11383 (N_11383,N_10528,N_10972);
nor U11384 (N_11384,N_10844,N_10828);
nand U11385 (N_11385,N_10689,N_10697);
or U11386 (N_11386,N_10608,N_10964);
xnor U11387 (N_11387,N_10891,N_10533);
or U11388 (N_11388,N_10905,N_11137);
nor U11389 (N_11389,N_11016,N_10661);
xnor U11390 (N_11390,N_10541,N_10659);
or U11391 (N_11391,N_11019,N_10686);
nand U11392 (N_11392,N_10870,N_10807);
and U11393 (N_11393,N_10770,N_10822);
nand U11394 (N_11394,N_11091,N_10949);
nor U11395 (N_11395,N_11240,N_10633);
nand U11396 (N_11396,N_11041,N_11175);
nor U11397 (N_11397,N_10935,N_10699);
or U11398 (N_11398,N_10884,N_10601);
nor U11399 (N_11399,N_10605,N_10995);
xnor U11400 (N_11400,N_10866,N_10625);
or U11401 (N_11401,N_10977,N_10918);
xor U11402 (N_11402,N_11230,N_10830);
and U11403 (N_11403,N_11099,N_11200);
nand U11404 (N_11404,N_10808,N_10863);
nand U11405 (N_11405,N_10510,N_10741);
xnor U11406 (N_11406,N_10774,N_10500);
nand U11407 (N_11407,N_10789,N_10540);
xnor U11408 (N_11408,N_10559,N_11125);
xor U11409 (N_11409,N_11076,N_10776);
and U11410 (N_11410,N_11209,N_10550);
and U11411 (N_11411,N_10568,N_10503);
nand U11412 (N_11412,N_11008,N_10950);
nor U11413 (N_11413,N_10643,N_10680);
or U11414 (N_11414,N_10773,N_10980);
and U11415 (N_11415,N_10743,N_10646);
nand U11416 (N_11416,N_10742,N_10617);
xor U11417 (N_11417,N_10966,N_10576);
and U11418 (N_11418,N_11194,N_11129);
nor U11419 (N_11419,N_11030,N_11005);
and U11420 (N_11420,N_10589,N_11211);
or U11421 (N_11421,N_10726,N_10665);
nand U11422 (N_11422,N_11160,N_10829);
xor U11423 (N_11423,N_10511,N_11247);
and U11424 (N_11424,N_10591,N_11141);
or U11425 (N_11425,N_11229,N_11001);
or U11426 (N_11426,N_10960,N_10570);
or U11427 (N_11427,N_10754,N_10745);
nand U11428 (N_11428,N_11131,N_11126);
nand U11429 (N_11429,N_10612,N_10768);
nor U11430 (N_11430,N_10917,N_11212);
xor U11431 (N_11431,N_11015,N_10532);
nand U11432 (N_11432,N_10524,N_10758);
xnor U11433 (N_11433,N_10615,N_11007);
nand U11434 (N_11434,N_10513,N_11066);
and U11435 (N_11435,N_10735,N_10815);
xnor U11436 (N_11436,N_10946,N_10606);
nor U11437 (N_11437,N_10861,N_10857);
xnor U11438 (N_11438,N_10920,N_10886);
nand U11439 (N_11439,N_11078,N_10785);
xnor U11440 (N_11440,N_10717,N_10982);
nand U11441 (N_11441,N_10725,N_10953);
xor U11442 (N_11442,N_10720,N_10859);
nand U11443 (N_11443,N_11151,N_10907);
xnor U11444 (N_11444,N_11103,N_10865);
and U11445 (N_11445,N_10733,N_11226);
xor U11446 (N_11446,N_11028,N_10996);
or U11447 (N_11447,N_10974,N_11032);
nor U11448 (N_11448,N_11029,N_10778);
nor U11449 (N_11449,N_10520,N_10536);
xor U11450 (N_11450,N_11138,N_11049);
xnor U11451 (N_11451,N_10856,N_10897);
xnor U11452 (N_11452,N_10948,N_11199);
nand U11453 (N_11453,N_10928,N_10597);
and U11454 (N_11454,N_10594,N_11026);
or U11455 (N_11455,N_10574,N_10599);
and U11456 (N_11456,N_11134,N_11000);
xnor U11457 (N_11457,N_10973,N_10713);
nand U11458 (N_11458,N_11085,N_10872);
xor U11459 (N_11459,N_11143,N_11224);
nor U11460 (N_11460,N_10687,N_10802);
nor U11461 (N_11461,N_10847,N_11034);
nand U11462 (N_11462,N_10855,N_11036);
xnor U11463 (N_11463,N_10903,N_10954);
or U11464 (N_11464,N_11245,N_10734);
nand U11465 (N_11465,N_10877,N_10933);
and U11466 (N_11466,N_10737,N_10845);
nand U11467 (N_11467,N_10938,N_10806);
nor U11468 (N_11468,N_10967,N_10627);
and U11469 (N_11469,N_11221,N_10728);
nand U11470 (N_11470,N_10696,N_10585);
xnor U11471 (N_11471,N_10767,N_10751);
xnor U11472 (N_11472,N_11157,N_11239);
nand U11473 (N_11473,N_10558,N_10987);
nor U11474 (N_11474,N_10824,N_10618);
nand U11475 (N_11475,N_10853,N_10989);
nand U11476 (N_11476,N_11086,N_10931);
nor U11477 (N_11477,N_10652,N_11047);
or U11478 (N_11478,N_10885,N_11092);
nand U11479 (N_11479,N_10656,N_11227);
xnor U11480 (N_11480,N_10556,N_10881);
and U11481 (N_11481,N_10834,N_10782);
nand U11482 (N_11482,N_10640,N_10586);
nand U11483 (N_11483,N_11218,N_11035);
and U11484 (N_11484,N_10554,N_11128);
or U11485 (N_11485,N_10850,N_10674);
and U11486 (N_11486,N_10673,N_11039);
nand U11487 (N_11487,N_10704,N_10662);
nor U11488 (N_11488,N_11233,N_11045);
nor U11489 (N_11489,N_11113,N_11148);
or U11490 (N_11490,N_10603,N_10602);
xnor U11491 (N_11491,N_10676,N_10764);
xnor U11492 (N_11492,N_10930,N_11106);
nor U11493 (N_11493,N_10826,N_11115);
nand U11494 (N_11494,N_10864,N_11238);
nand U11495 (N_11495,N_11145,N_10675);
and U11496 (N_11496,N_11104,N_10979);
or U11497 (N_11497,N_10685,N_10827);
nor U11498 (N_11498,N_11150,N_10868);
or U11499 (N_11499,N_11214,N_11122);
and U11500 (N_11500,N_10772,N_10779);
xnor U11501 (N_11501,N_11018,N_10763);
xor U11502 (N_11502,N_10719,N_10849);
and U11503 (N_11503,N_10985,N_10970);
xor U11504 (N_11504,N_11121,N_10738);
or U11505 (N_11505,N_10888,N_10957);
nand U11506 (N_11506,N_10711,N_10562);
and U11507 (N_11507,N_11061,N_10922);
nand U11508 (N_11508,N_10941,N_11060);
nand U11509 (N_11509,N_10666,N_11170);
nand U11510 (N_11510,N_10516,N_11043);
nand U11511 (N_11511,N_10621,N_10684);
nand U11512 (N_11512,N_10991,N_11058);
nor U11513 (N_11513,N_10760,N_10908);
xnor U11514 (N_11514,N_11119,N_11048);
xnor U11515 (N_11515,N_11051,N_10841);
nand U11516 (N_11516,N_10860,N_10943);
xnor U11517 (N_11517,N_10965,N_10846);
or U11518 (N_11518,N_10632,N_10906);
or U11519 (N_11519,N_10832,N_10682);
nor U11520 (N_11520,N_11072,N_10915);
nor U11521 (N_11521,N_11059,N_11152);
or U11522 (N_11522,N_11197,N_10731);
nand U11523 (N_11523,N_11087,N_10716);
or U11524 (N_11524,N_10912,N_11033);
and U11525 (N_11525,N_10790,N_10645);
and U11526 (N_11526,N_11192,N_10879);
nor U11527 (N_11527,N_10792,N_11202);
nand U11528 (N_11528,N_11081,N_10914);
and U11529 (N_11529,N_10563,N_10809);
nor U11530 (N_11530,N_10504,N_10766);
or U11531 (N_11531,N_10678,N_10705);
nor U11532 (N_11532,N_10560,N_11136);
nor U11533 (N_11533,N_10793,N_10819);
or U11534 (N_11534,N_10971,N_10571);
or U11535 (N_11535,N_10660,N_10623);
nor U11536 (N_11536,N_11158,N_10583);
and U11537 (N_11537,N_11083,N_10732);
xor U11538 (N_11538,N_10619,N_10781);
nor U11539 (N_11539,N_10796,N_10628);
or U11540 (N_11540,N_10588,N_10975);
and U11541 (N_11541,N_10992,N_10691);
nor U11542 (N_11542,N_10969,N_10688);
xnor U11543 (N_11543,N_11168,N_10544);
nor U11544 (N_11544,N_11133,N_11040);
nor U11545 (N_11545,N_11185,N_11065);
nand U11546 (N_11546,N_10813,N_10653);
xor U11547 (N_11547,N_11183,N_10693);
nand U11548 (N_11548,N_10525,N_10721);
nor U11549 (N_11549,N_10512,N_11127);
xnor U11550 (N_11550,N_10804,N_11234);
or U11551 (N_11551,N_11073,N_10923);
nor U11552 (N_11552,N_10607,N_10521);
nor U11553 (N_11553,N_11242,N_11179);
nand U11554 (N_11554,N_10551,N_11054);
or U11555 (N_11555,N_11235,N_10561);
xnor U11556 (N_11556,N_10670,N_11243);
xor U11557 (N_11557,N_10761,N_10644);
or U11558 (N_11558,N_10543,N_11165);
xor U11559 (N_11559,N_10630,N_11219);
and U11560 (N_11560,N_10710,N_11171);
and U11561 (N_11561,N_10658,N_10714);
and U11562 (N_11562,N_10755,N_10956);
xor U11563 (N_11563,N_10874,N_10548);
xor U11564 (N_11564,N_11204,N_10557);
or U11565 (N_11565,N_11057,N_10976);
and U11566 (N_11566,N_10805,N_10593);
xor U11567 (N_11567,N_11095,N_10506);
xor U11568 (N_11568,N_10823,N_10955);
xnor U11569 (N_11569,N_10740,N_10962);
and U11570 (N_11570,N_10647,N_10986);
and U11571 (N_11571,N_10587,N_11017);
nor U11572 (N_11572,N_11021,N_11116);
nor U11573 (N_11573,N_11055,N_10634);
nor U11574 (N_11574,N_10681,N_10668);
xor U11575 (N_11575,N_11232,N_11231);
nand U11576 (N_11576,N_11155,N_10919);
and U11577 (N_11577,N_10708,N_10898);
nand U11578 (N_11578,N_10650,N_10862);
nand U11579 (N_11579,N_10626,N_11096);
xor U11580 (N_11580,N_11042,N_10581);
nor U11581 (N_11581,N_10590,N_10892);
nand U11582 (N_11582,N_11074,N_10649);
xor U11583 (N_11583,N_10867,N_11023);
nand U11584 (N_11584,N_11020,N_11053);
nor U11585 (N_11585,N_10959,N_11013);
or U11586 (N_11586,N_10722,N_11080);
nand U11587 (N_11587,N_11089,N_10507);
and U11588 (N_11588,N_10921,N_11215);
or U11589 (N_11589,N_10997,N_11002);
xor U11590 (N_11590,N_10555,N_11147);
xor U11591 (N_11591,N_10651,N_11064);
xnor U11592 (N_11592,N_10552,N_11173);
nand U11593 (N_11593,N_11069,N_10945);
or U11594 (N_11594,N_10909,N_11220);
and U11595 (N_11595,N_10611,N_11177);
nand U11596 (N_11596,N_10900,N_10729);
nand U11597 (N_11597,N_10801,N_10648);
xnor U11598 (N_11598,N_10925,N_10567);
xnor U11599 (N_11599,N_10577,N_10564);
nor U11600 (N_11600,N_10873,N_11031);
xor U11601 (N_11601,N_10641,N_11068);
nand U11602 (N_11602,N_11161,N_10952);
xor U11603 (N_11603,N_10794,N_10514);
nand U11604 (N_11604,N_10635,N_10978);
or U11605 (N_11605,N_10840,N_10880);
and U11606 (N_11606,N_10842,N_10787);
or U11607 (N_11607,N_11011,N_11184);
xnor U11608 (N_11608,N_11062,N_11139);
and U11609 (N_11609,N_11142,N_10936);
and U11610 (N_11610,N_10795,N_11178);
or U11611 (N_11611,N_10723,N_10622);
or U11612 (N_11612,N_10791,N_10998);
nand U11613 (N_11613,N_10700,N_10535);
or U11614 (N_11614,N_10762,N_10839);
nand U11615 (N_11615,N_11172,N_10600);
xnor U11616 (N_11616,N_11004,N_11236);
xnor U11617 (N_11617,N_11193,N_11135);
xnor U11618 (N_11618,N_10780,N_10736);
nand U11619 (N_11619,N_11210,N_10899);
nand U11620 (N_11620,N_10629,N_10616);
nand U11621 (N_11621,N_10519,N_11244);
or U11622 (N_11622,N_10817,N_10695);
and U11623 (N_11623,N_10637,N_10518);
or U11624 (N_11624,N_10786,N_11003);
xor U11625 (N_11625,N_10653,N_10922);
or U11626 (N_11626,N_10577,N_11212);
or U11627 (N_11627,N_10721,N_10977);
xor U11628 (N_11628,N_10922,N_10569);
nor U11629 (N_11629,N_10822,N_11060);
xnor U11630 (N_11630,N_10614,N_11164);
nand U11631 (N_11631,N_11009,N_11080);
nand U11632 (N_11632,N_11174,N_10518);
and U11633 (N_11633,N_11092,N_10565);
nor U11634 (N_11634,N_10623,N_10530);
or U11635 (N_11635,N_10926,N_10724);
nand U11636 (N_11636,N_10716,N_11166);
xor U11637 (N_11637,N_11116,N_11128);
nand U11638 (N_11638,N_10952,N_11229);
nor U11639 (N_11639,N_11047,N_11187);
nor U11640 (N_11640,N_10975,N_10692);
nand U11641 (N_11641,N_11044,N_11208);
xnor U11642 (N_11642,N_10783,N_11240);
nand U11643 (N_11643,N_10714,N_10866);
nor U11644 (N_11644,N_11006,N_10552);
nor U11645 (N_11645,N_11226,N_10754);
xor U11646 (N_11646,N_10767,N_10608);
nand U11647 (N_11647,N_10549,N_10728);
or U11648 (N_11648,N_10890,N_10765);
nor U11649 (N_11649,N_10681,N_10738);
nor U11650 (N_11650,N_10680,N_10565);
xnor U11651 (N_11651,N_11025,N_10769);
xor U11652 (N_11652,N_10695,N_10735);
nor U11653 (N_11653,N_10758,N_10814);
xnor U11654 (N_11654,N_10837,N_10772);
xor U11655 (N_11655,N_11169,N_10575);
nand U11656 (N_11656,N_10534,N_11237);
and U11657 (N_11657,N_10568,N_11158);
or U11658 (N_11658,N_10890,N_11100);
nor U11659 (N_11659,N_11000,N_10632);
and U11660 (N_11660,N_11180,N_11224);
nand U11661 (N_11661,N_11047,N_10615);
or U11662 (N_11662,N_11220,N_10975);
and U11663 (N_11663,N_10985,N_10565);
and U11664 (N_11664,N_10918,N_10609);
nor U11665 (N_11665,N_10990,N_11237);
or U11666 (N_11666,N_10662,N_10736);
or U11667 (N_11667,N_10809,N_11050);
xor U11668 (N_11668,N_10910,N_10992);
nand U11669 (N_11669,N_10514,N_10657);
or U11670 (N_11670,N_11085,N_10803);
nand U11671 (N_11671,N_10620,N_10837);
nor U11672 (N_11672,N_10921,N_11005);
nor U11673 (N_11673,N_11144,N_10517);
and U11674 (N_11674,N_10945,N_11162);
and U11675 (N_11675,N_10538,N_10800);
nor U11676 (N_11676,N_11125,N_10667);
nor U11677 (N_11677,N_11029,N_10754);
xnor U11678 (N_11678,N_10828,N_11236);
or U11679 (N_11679,N_10977,N_10806);
and U11680 (N_11680,N_10774,N_10904);
nand U11681 (N_11681,N_10575,N_10811);
or U11682 (N_11682,N_10836,N_11207);
and U11683 (N_11683,N_10599,N_10823);
or U11684 (N_11684,N_10745,N_10807);
nand U11685 (N_11685,N_11198,N_11064);
nand U11686 (N_11686,N_10515,N_10765);
nor U11687 (N_11687,N_10578,N_10857);
or U11688 (N_11688,N_10882,N_10610);
xnor U11689 (N_11689,N_10873,N_11093);
and U11690 (N_11690,N_11020,N_11035);
nand U11691 (N_11691,N_10511,N_10940);
nand U11692 (N_11692,N_10723,N_10961);
or U11693 (N_11693,N_10960,N_10966);
and U11694 (N_11694,N_10617,N_11190);
nand U11695 (N_11695,N_10604,N_10766);
nor U11696 (N_11696,N_10769,N_10707);
or U11697 (N_11697,N_10973,N_10756);
nand U11698 (N_11698,N_10989,N_10517);
nand U11699 (N_11699,N_10799,N_11232);
xnor U11700 (N_11700,N_10864,N_11063);
xnor U11701 (N_11701,N_11212,N_11105);
or U11702 (N_11702,N_10988,N_10858);
nor U11703 (N_11703,N_10608,N_10500);
nor U11704 (N_11704,N_10576,N_10891);
or U11705 (N_11705,N_10682,N_10911);
nor U11706 (N_11706,N_11098,N_11082);
xor U11707 (N_11707,N_10548,N_10884);
xnor U11708 (N_11708,N_10774,N_10706);
or U11709 (N_11709,N_11127,N_11202);
or U11710 (N_11710,N_10974,N_11106);
xor U11711 (N_11711,N_11166,N_10650);
or U11712 (N_11712,N_10775,N_10795);
xor U11713 (N_11713,N_10622,N_10963);
and U11714 (N_11714,N_10831,N_10940);
nand U11715 (N_11715,N_11143,N_10917);
nor U11716 (N_11716,N_11197,N_10987);
and U11717 (N_11717,N_10991,N_10928);
xnor U11718 (N_11718,N_10569,N_11190);
or U11719 (N_11719,N_10584,N_10678);
nor U11720 (N_11720,N_10578,N_10924);
nand U11721 (N_11721,N_10872,N_10978);
nor U11722 (N_11722,N_11168,N_10518);
nand U11723 (N_11723,N_10939,N_10737);
nand U11724 (N_11724,N_10982,N_10933);
and U11725 (N_11725,N_11116,N_11120);
nor U11726 (N_11726,N_10503,N_11064);
nor U11727 (N_11727,N_10752,N_10764);
nand U11728 (N_11728,N_11058,N_10616);
or U11729 (N_11729,N_11130,N_10550);
nor U11730 (N_11730,N_11027,N_10917);
or U11731 (N_11731,N_10702,N_11055);
xnor U11732 (N_11732,N_10726,N_10675);
nand U11733 (N_11733,N_10639,N_11236);
nor U11734 (N_11734,N_11181,N_10945);
or U11735 (N_11735,N_10870,N_10905);
and U11736 (N_11736,N_10578,N_10954);
nor U11737 (N_11737,N_11043,N_10971);
and U11738 (N_11738,N_10591,N_10751);
xnor U11739 (N_11739,N_10528,N_11113);
xnor U11740 (N_11740,N_10546,N_10624);
and U11741 (N_11741,N_10711,N_10634);
and U11742 (N_11742,N_11153,N_10592);
xnor U11743 (N_11743,N_10688,N_10950);
xnor U11744 (N_11744,N_11032,N_10894);
and U11745 (N_11745,N_10958,N_11124);
or U11746 (N_11746,N_10825,N_10801);
xnor U11747 (N_11747,N_11123,N_10903);
xnor U11748 (N_11748,N_10817,N_10867);
nor U11749 (N_11749,N_10656,N_11222);
or U11750 (N_11750,N_10698,N_10866);
and U11751 (N_11751,N_11083,N_10545);
and U11752 (N_11752,N_10795,N_10907);
or U11753 (N_11753,N_11131,N_10638);
xor U11754 (N_11754,N_10765,N_11079);
or U11755 (N_11755,N_11071,N_11134);
and U11756 (N_11756,N_11194,N_10944);
nor U11757 (N_11757,N_10978,N_10685);
or U11758 (N_11758,N_10842,N_10726);
nor U11759 (N_11759,N_11120,N_10520);
nand U11760 (N_11760,N_10571,N_11223);
xnor U11761 (N_11761,N_10858,N_11163);
nand U11762 (N_11762,N_11049,N_10528);
and U11763 (N_11763,N_10792,N_10503);
nand U11764 (N_11764,N_11115,N_11193);
or U11765 (N_11765,N_10796,N_10688);
nand U11766 (N_11766,N_10912,N_10880);
nor U11767 (N_11767,N_10943,N_11098);
xnor U11768 (N_11768,N_10672,N_10666);
and U11769 (N_11769,N_10850,N_10763);
xnor U11770 (N_11770,N_10852,N_10949);
and U11771 (N_11771,N_11064,N_10914);
xor U11772 (N_11772,N_10722,N_10773);
xnor U11773 (N_11773,N_11181,N_11220);
or U11774 (N_11774,N_11025,N_10721);
or U11775 (N_11775,N_10850,N_10857);
nand U11776 (N_11776,N_10660,N_10944);
and U11777 (N_11777,N_11033,N_10714);
and U11778 (N_11778,N_10575,N_10599);
xnor U11779 (N_11779,N_11031,N_10920);
or U11780 (N_11780,N_10997,N_10846);
and U11781 (N_11781,N_10673,N_10753);
and U11782 (N_11782,N_11212,N_11119);
or U11783 (N_11783,N_11044,N_10950);
nand U11784 (N_11784,N_11180,N_10687);
or U11785 (N_11785,N_11117,N_10971);
and U11786 (N_11786,N_10950,N_10574);
nor U11787 (N_11787,N_11178,N_11050);
nand U11788 (N_11788,N_11206,N_11165);
and U11789 (N_11789,N_10760,N_10599);
xnor U11790 (N_11790,N_10562,N_11160);
nand U11791 (N_11791,N_11034,N_10997);
nor U11792 (N_11792,N_10546,N_11057);
and U11793 (N_11793,N_10506,N_10500);
and U11794 (N_11794,N_11196,N_10592);
nor U11795 (N_11795,N_10902,N_11012);
nand U11796 (N_11796,N_11135,N_10569);
nand U11797 (N_11797,N_10820,N_10730);
xor U11798 (N_11798,N_10599,N_11086);
and U11799 (N_11799,N_10529,N_11159);
and U11800 (N_11800,N_10863,N_10942);
and U11801 (N_11801,N_10976,N_10512);
and U11802 (N_11802,N_11098,N_10503);
nand U11803 (N_11803,N_11046,N_10922);
nor U11804 (N_11804,N_10968,N_11146);
xnor U11805 (N_11805,N_11163,N_11124);
or U11806 (N_11806,N_11238,N_10651);
xor U11807 (N_11807,N_11039,N_10669);
and U11808 (N_11808,N_11016,N_11223);
nor U11809 (N_11809,N_10983,N_10595);
nand U11810 (N_11810,N_10590,N_10517);
and U11811 (N_11811,N_11241,N_10950);
nand U11812 (N_11812,N_10757,N_10624);
and U11813 (N_11813,N_10591,N_10978);
nand U11814 (N_11814,N_10846,N_11042);
and U11815 (N_11815,N_10817,N_11069);
nand U11816 (N_11816,N_10739,N_10846);
nand U11817 (N_11817,N_11166,N_10676);
xor U11818 (N_11818,N_10869,N_10785);
or U11819 (N_11819,N_10759,N_11094);
xnor U11820 (N_11820,N_10540,N_10859);
nand U11821 (N_11821,N_10736,N_10593);
nand U11822 (N_11822,N_11039,N_11229);
xor U11823 (N_11823,N_10936,N_11076);
and U11824 (N_11824,N_11112,N_10689);
nor U11825 (N_11825,N_10577,N_10882);
xnor U11826 (N_11826,N_10639,N_10972);
or U11827 (N_11827,N_10823,N_10679);
xor U11828 (N_11828,N_11134,N_11155);
nand U11829 (N_11829,N_10830,N_11102);
nand U11830 (N_11830,N_10869,N_10769);
and U11831 (N_11831,N_10774,N_10681);
and U11832 (N_11832,N_11213,N_10561);
nor U11833 (N_11833,N_11136,N_11107);
nor U11834 (N_11834,N_10674,N_11060);
xor U11835 (N_11835,N_10769,N_11042);
and U11836 (N_11836,N_10829,N_10907);
and U11837 (N_11837,N_11196,N_11223);
or U11838 (N_11838,N_10743,N_11171);
nand U11839 (N_11839,N_10961,N_11138);
and U11840 (N_11840,N_11240,N_11158);
and U11841 (N_11841,N_11209,N_11114);
xor U11842 (N_11842,N_10554,N_10973);
xnor U11843 (N_11843,N_10557,N_11013);
or U11844 (N_11844,N_10807,N_10552);
or U11845 (N_11845,N_11025,N_10512);
nand U11846 (N_11846,N_11152,N_10721);
nor U11847 (N_11847,N_10602,N_11188);
and U11848 (N_11848,N_11076,N_10989);
xor U11849 (N_11849,N_10550,N_10814);
nand U11850 (N_11850,N_10979,N_10862);
nand U11851 (N_11851,N_10962,N_11181);
nor U11852 (N_11852,N_10958,N_11167);
or U11853 (N_11853,N_11048,N_10535);
xor U11854 (N_11854,N_11163,N_10962);
nor U11855 (N_11855,N_11044,N_11206);
or U11856 (N_11856,N_10649,N_10994);
nand U11857 (N_11857,N_10584,N_10798);
nand U11858 (N_11858,N_10948,N_11071);
and U11859 (N_11859,N_10984,N_11121);
nor U11860 (N_11860,N_10792,N_10946);
or U11861 (N_11861,N_10783,N_10864);
nand U11862 (N_11862,N_10817,N_10865);
or U11863 (N_11863,N_10665,N_10787);
nand U11864 (N_11864,N_10790,N_10745);
nor U11865 (N_11865,N_11243,N_11165);
and U11866 (N_11866,N_11124,N_10746);
and U11867 (N_11867,N_11183,N_11042);
and U11868 (N_11868,N_10605,N_10715);
nor U11869 (N_11869,N_10748,N_11186);
or U11870 (N_11870,N_10659,N_11014);
or U11871 (N_11871,N_10619,N_10737);
xor U11872 (N_11872,N_10517,N_10832);
and U11873 (N_11873,N_11113,N_10689);
and U11874 (N_11874,N_10832,N_11194);
nand U11875 (N_11875,N_11009,N_10594);
or U11876 (N_11876,N_10801,N_11104);
nor U11877 (N_11877,N_10660,N_10522);
and U11878 (N_11878,N_10570,N_10916);
xnor U11879 (N_11879,N_10610,N_10581);
and U11880 (N_11880,N_10796,N_10947);
and U11881 (N_11881,N_11246,N_11046);
xnor U11882 (N_11882,N_11171,N_11191);
nand U11883 (N_11883,N_10561,N_10922);
or U11884 (N_11884,N_10901,N_10559);
xor U11885 (N_11885,N_11181,N_10688);
and U11886 (N_11886,N_10748,N_11229);
nand U11887 (N_11887,N_10885,N_11072);
and U11888 (N_11888,N_10505,N_10977);
nand U11889 (N_11889,N_10932,N_11159);
xor U11890 (N_11890,N_10782,N_11218);
nand U11891 (N_11891,N_10810,N_10795);
xnor U11892 (N_11892,N_10905,N_11173);
or U11893 (N_11893,N_10556,N_11051);
or U11894 (N_11894,N_11026,N_11087);
nor U11895 (N_11895,N_11233,N_10536);
xor U11896 (N_11896,N_10851,N_10926);
and U11897 (N_11897,N_10785,N_10714);
or U11898 (N_11898,N_11218,N_11051);
nor U11899 (N_11899,N_10540,N_10824);
and U11900 (N_11900,N_10898,N_10938);
or U11901 (N_11901,N_10701,N_11154);
and U11902 (N_11902,N_10829,N_11029);
nand U11903 (N_11903,N_10950,N_10946);
nor U11904 (N_11904,N_10661,N_11059);
nor U11905 (N_11905,N_10643,N_11092);
and U11906 (N_11906,N_11073,N_10664);
or U11907 (N_11907,N_11184,N_11231);
or U11908 (N_11908,N_10784,N_10797);
nor U11909 (N_11909,N_10655,N_10901);
nor U11910 (N_11910,N_11116,N_10545);
xnor U11911 (N_11911,N_10723,N_11234);
or U11912 (N_11912,N_10587,N_11104);
or U11913 (N_11913,N_10760,N_11226);
xnor U11914 (N_11914,N_10756,N_11082);
nand U11915 (N_11915,N_10834,N_10933);
and U11916 (N_11916,N_10570,N_11123);
nand U11917 (N_11917,N_10899,N_11230);
or U11918 (N_11918,N_10819,N_11243);
xor U11919 (N_11919,N_10648,N_11173);
or U11920 (N_11920,N_11036,N_10920);
xnor U11921 (N_11921,N_10700,N_11153);
or U11922 (N_11922,N_10780,N_11087);
xnor U11923 (N_11923,N_11082,N_11127);
nor U11924 (N_11924,N_10762,N_10519);
and U11925 (N_11925,N_11206,N_11153);
nor U11926 (N_11926,N_10989,N_10947);
nor U11927 (N_11927,N_10550,N_10676);
nor U11928 (N_11928,N_11172,N_10553);
or U11929 (N_11929,N_11013,N_11113);
nor U11930 (N_11930,N_11008,N_11229);
or U11931 (N_11931,N_11009,N_10668);
xnor U11932 (N_11932,N_10514,N_11238);
xnor U11933 (N_11933,N_10582,N_10887);
nand U11934 (N_11934,N_10783,N_11244);
nor U11935 (N_11935,N_11249,N_10574);
xnor U11936 (N_11936,N_11141,N_11055);
xnor U11937 (N_11937,N_10536,N_10715);
and U11938 (N_11938,N_10999,N_11207);
nand U11939 (N_11939,N_10936,N_10625);
nor U11940 (N_11940,N_10731,N_10824);
or U11941 (N_11941,N_11024,N_10508);
nor U11942 (N_11942,N_10882,N_10523);
xor U11943 (N_11943,N_11092,N_10570);
xor U11944 (N_11944,N_10820,N_11154);
nand U11945 (N_11945,N_11099,N_10998);
nor U11946 (N_11946,N_10879,N_11073);
and U11947 (N_11947,N_10991,N_10957);
nand U11948 (N_11948,N_10532,N_10720);
nor U11949 (N_11949,N_10548,N_10859);
nand U11950 (N_11950,N_10560,N_11181);
xnor U11951 (N_11951,N_10868,N_10873);
xnor U11952 (N_11952,N_10841,N_10931);
or U11953 (N_11953,N_10874,N_11216);
and U11954 (N_11954,N_10642,N_10689);
nand U11955 (N_11955,N_10544,N_11146);
nand U11956 (N_11956,N_10703,N_11193);
and U11957 (N_11957,N_10622,N_10680);
and U11958 (N_11958,N_11135,N_11239);
and U11959 (N_11959,N_10508,N_10590);
nand U11960 (N_11960,N_11205,N_10747);
nand U11961 (N_11961,N_10922,N_10671);
nand U11962 (N_11962,N_11114,N_10570);
xor U11963 (N_11963,N_10555,N_10719);
nor U11964 (N_11964,N_11183,N_10748);
nand U11965 (N_11965,N_10775,N_11040);
and U11966 (N_11966,N_10776,N_10953);
or U11967 (N_11967,N_10510,N_11161);
xnor U11968 (N_11968,N_10642,N_10887);
or U11969 (N_11969,N_10740,N_10984);
or U11970 (N_11970,N_11090,N_10500);
nor U11971 (N_11971,N_10637,N_11130);
xor U11972 (N_11972,N_10843,N_11144);
nor U11973 (N_11973,N_11207,N_10673);
xnor U11974 (N_11974,N_11055,N_11077);
xor U11975 (N_11975,N_10622,N_10989);
xnor U11976 (N_11976,N_10955,N_10885);
or U11977 (N_11977,N_10694,N_10944);
nor U11978 (N_11978,N_11219,N_10527);
and U11979 (N_11979,N_11049,N_11157);
and U11980 (N_11980,N_10504,N_10948);
nor U11981 (N_11981,N_10915,N_10945);
nand U11982 (N_11982,N_10985,N_10528);
and U11983 (N_11983,N_10994,N_10942);
nand U11984 (N_11984,N_10605,N_10502);
xor U11985 (N_11985,N_11236,N_10773);
or U11986 (N_11986,N_10851,N_11028);
nor U11987 (N_11987,N_11181,N_11182);
nor U11988 (N_11988,N_11241,N_11029);
nand U11989 (N_11989,N_10832,N_10611);
xor U11990 (N_11990,N_11019,N_11145);
nand U11991 (N_11991,N_10707,N_10717);
and U11992 (N_11992,N_10545,N_11201);
nand U11993 (N_11993,N_11015,N_10953);
nand U11994 (N_11994,N_10724,N_10864);
nand U11995 (N_11995,N_11158,N_11097);
nand U11996 (N_11996,N_10815,N_11043);
xor U11997 (N_11997,N_10853,N_11134);
xor U11998 (N_11998,N_11197,N_10927);
xor U11999 (N_11999,N_10756,N_11103);
nand U12000 (N_12000,N_11582,N_11886);
nor U12001 (N_12001,N_11774,N_11725);
nand U12002 (N_12002,N_11601,N_11669);
and U12003 (N_12003,N_11777,N_11987);
nor U12004 (N_12004,N_11898,N_11876);
nor U12005 (N_12005,N_11361,N_11716);
nand U12006 (N_12006,N_11834,N_11383);
or U12007 (N_12007,N_11400,N_11972);
xor U12008 (N_12008,N_11457,N_11874);
nand U12009 (N_12009,N_11757,N_11707);
or U12010 (N_12010,N_11465,N_11281);
xnor U12011 (N_12011,N_11598,N_11830);
and U12012 (N_12012,N_11971,N_11862);
or U12013 (N_12013,N_11866,N_11753);
nor U12014 (N_12014,N_11856,N_11515);
nand U12015 (N_12015,N_11736,N_11307);
nor U12016 (N_12016,N_11375,N_11890);
xnor U12017 (N_12017,N_11634,N_11430);
nand U12018 (N_12018,N_11351,N_11333);
nor U12019 (N_12019,N_11626,N_11259);
nand U12020 (N_12020,N_11426,N_11906);
nor U12021 (N_12021,N_11620,N_11592);
or U12022 (N_12022,N_11917,N_11904);
nand U12023 (N_12023,N_11937,N_11966);
or U12024 (N_12024,N_11415,N_11536);
and U12025 (N_12025,N_11294,N_11401);
nand U12026 (N_12026,N_11545,N_11570);
nand U12027 (N_12027,N_11732,N_11493);
xor U12028 (N_12028,N_11702,N_11782);
nand U12029 (N_12029,N_11901,N_11595);
nand U12030 (N_12030,N_11900,N_11655);
nand U12031 (N_12031,N_11588,N_11377);
nand U12032 (N_12032,N_11758,N_11916);
or U12033 (N_12033,N_11995,N_11389);
nor U12034 (N_12034,N_11612,N_11529);
or U12035 (N_12035,N_11583,N_11441);
nand U12036 (N_12036,N_11387,N_11839);
and U12037 (N_12037,N_11539,N_11662);
nand U12038 (N_12038,N_11823,N_11791);
nor U12039 (N_12039,N_11799,N_11310);
or U12040 (N_12040,N_11433,N_11396);
and U12041 (N_12041,N_11747,N_11462);
and U12042 (N_12042,N_11501,N_11522);
or U12043 (N_12043,N_11704,N_11836);
and U12044 (N_12044,N_11269,N_11502);
or U12045 (N_12045,N_11721,N_11981);
and U12046 (N_12046,N_11825,N_11684);
xor U12047 (N_12047,N_11558,N_11474);
nor U12048 (N_12048,N_11727,N_11434);
nand U12049 (N_12049,N_11820,N_11413);
nand U12050 (N_12050,N_11359,N_11802);
and U12051 (N_12051,N_11309,N_11629);
nand U12052 (N_12052,N_11475,N_11258);
nor U12053 (N_12053,N_11844,N_11533);
nor U12054 (N_12054,N_11745,N_11718);
or U12055 (N_12055,N_11445,N_11977);
nor U12056 (N_12056,N_11879,N_11869);
and U12057 (N_12057,N_11665,N_11391);
or U12058 (N_12058,N_11499,N_11819);
xor U12059 (N_12059,N_11689,N_11305);
or U12060 (N_12060,N_11978,N_11509);
and U12061 (N_12061,N_11677,N_11323);
or U12062 (N_12062,N_11255,N_11503);
nand U12063 (N_12063,N_11720,N_11970);
nand U12064 (N_12064,N_11518,N_11764);
nor U12065 (N_12065,N_11930,N_11451);
or U12066 (N_12066,N_11691,N_11628);
or U12067 (N_12067,N_11708,N_11311);
nand U12068 (N_12068,N_11602,N_11342);
or U12069 (N_12069,N_11479,N_11286);
and U12070 (N_12070,N_11822,N_11840);
nor U12071 (N_12071,N_11454,N_11641);
nor U12072 (N_12072,N_11306,N_11251);
nor U12073 (N_12073,N_11636,N_11722);
and U12074 (N_12074,N_11557,N_11423);
nand U12075 (N_12075,N_11642,N_11374);
or U12076 (N_12076,N_11428,N_11644);
or U12077 (N_12077,N_11394,N_11650);
nand U12078 (N_12078,N_11399,N_11292);
nand U12079 (N_12079,N_11811,N_11594);
nor U12080 (N_12080,N_11769,N_11974);
xnor U12081 (N_12081,N_11914,N_11440);
or U12082 (N_12082,N_11637,N_11431);
nand U12083 (N_12083,N_11951,N_11439);
xnor U12084 (N_12084,N_11315,N_11339);
nand U12085 (N_12085,N_11562,N_11550);
xor U12086 (N_12086,N_11591,N_11920);
nor U12087 (N_12087,N_11861,N_11523);
or U12088 (N_12088,N_11918,N_11770);
and U12089 (N_12089,N_11297,N_11700);
or U12090 (N_12090,N_11646,N_11670);
and U12091 (N_12091,N_11982,N_11663);
and U12092 (N_12092,N_11997,N_11902);
or U12093 (N_12093,N_11751,N_11723);
xnor U12094 (N_12094,N_11907,N_11794);
or U12095 (N_12095,N_11809,N_11291);
and U12096 (N_12096,N_11976,N_11318);
nand U12097 (N_12097,N_11340,N_11468);
or U12098 (N_12098,N_11638,N_11345);
and U12099 (N_12099,N_11553,N_11657);
nand U12100 (N_12100,N_11572,N_11910);
nand U12101 (N_12101,N_11453,N_11568);
or U12102 (N_12102,N_11991,N_11923);
nand U12103 (N_12103,N_11563,N_11382);
xor U12104 (N_12104,N_11576,N_11648);
or U12105 (N_12105,N_11633,N_11565);
xor U12106 (N_12106,N_11875,N_11487);
and U12107 (N_12107,N_11537,N_11776);
xor U12108 (N_12108,N_11762,N_11852);
nor U12109 (N_12109,N_11754,N_11541);
nand U12110 (N_12110,N_11504,N_11372);
nor U12111 (N_12111,N_11936,N_11506);
nand U12112 (N_12112,N_11596,N_11765);
nor U12113 (N_12113,N_11253,N_11488);
or U12114 (N_12114,N_11327,N_11711);
xor U12115 (N_12115,N_11336,N_11485);
or U12116 (N_12116,N_11321,N_11514);
or U12117 (N_12117,N_11337,N_11276);
and U12118 (N_12118,N_11527,N_11380);
nor U12119 (N_12119,N_11800,N_11385);
and U12120 (N_12120,N_11694,N_11410);
xor U12121 (N_12121,N_11969,N_11760);
and U12122 (N_12122,N_11405,N_11960);
nor U12123 (N_12123,N_11889,N_11835);
nor U12124 (N_12124,N_11486,N_11731);
nor U12125 (N_12125,N_11567,N_11350);
nor U12126 (N_12126,N_11585,N_11639);
and U12127 (N_12127,N_11324,N_11797);
or U12128 (N_12128,N_11482,N_11564);
nand U12129 (N_12129,N_11547,N_11561);
nand U12130 (N_12130,N_11710,N_11845);
and U12131 (N_12131,N_11632,N_11697);
or U12132 (N_12132,N_11470,N_11891);
and U12133 (N_12133,N_11801,N_11744);
nand U12134 (N_12134,N_11322,N_11416);
and U12135 (N_12135,N_11554,N_11609);
nor U12136 (N_12136,N_11832,N_11579);
nand U12137 (N_12137,N_11614,N_11645);
nor U12138 (N_12138,N_11773,N_11566);
and U12139 (N_12139,N_11535,N_11544);
and U12140 (N_12140,N_11922,N_11422);
xor U12141 (N_12141,N_11654,N_11386);
xor U12142 (N_12142,N_11356,N_11792);
nand U12143 (N_12143,N_11290,N_11552);
or U12144 (N_12144,N_11652,N_11334);
and U12145 (N_12145,N_11548,N_11967);
or U12146 (N_12146,N_11301,N_11640);
or U12147 (N_12147,N_11685,N_11517);
nor U12148 (N_12148,N_11784,N_11709);
or U12149 (N_12149,N_11328,N_11540);
and U12150 (N_12150,N_11384,N_11667);
or U12151 (N_12151,N_11953,N_11962);
or U12152 (N_12152,N_11432,N_11429);
or U12153 (N_12153,N_11607,N_11894);
nor U12154 (N_12154,N_11559,N_11414);
nor U12155 (N_12155,N_11575,N_11473);
or U12156 (N_12156,N_11489,N_11870);
nand U12157 (N_12157,N_11302,N_11740);
and U12158 (N_12158,N_11942,N_11926);
nor U12159 (N_12159,N_11279,N_11829);
nand U12160 (N_12160,N_11603,N_11796);
xor U12161 (N_12161,N_11534,N_11887);
xor U12162 (N_12162,N_11980,N_11524);
nand U12163 (N_12163,N_11419,N_11938);
or U12164 (N_12164,N_11477,N_11590);
xor U12165 (N_12165,N_11409,N_11463);
or U12166 (N_12166,N_11376,N_11673);
and U12167 (N_12167,N_11947,N_11927);
or U12168 (N_12168,N_11828,N_11363);
nand U12169 (N_12169,N_11768,N_11883);
or U12170 (N_12170,N_11338,N_11466);
or U12171 (N_12171,N_11779,N_11317);
nand U12172 (N_12172,N_11521,N_11360);
nand U12173 (N_12173,N_11686,N_11846);
nor U12174 (N_12174,N_11847,N_11756);
xnor U12175 (N_12175,N_11480,N_11672);
xnor U12176 (N_12176,N_11516,N_11683);
or U12177 (N_12177,N_11742,N_11491);
xnor U12178 (N_12178,N_11934,N_11647);
xnor U12179 (N_12179,N_11873,N_11510);
xor U12180 (N_12180,N_11586,N_11366);
xnor U12181 (N_12181,N_11319,N_11496);
or U12182 (N_12182,N_11444,N_11717);
and U12183 (N_12183,N_11530,N_11734);
and U12184 (N_12184,N_11406,N_11701);
nor U12185 (N_12185,N_11417,N_11274);
xor U12186 (N_12186,N_11806,N_11420);
and U12187 (N_12187,N_11965,N_11766);
nor U12188 (N_12188,N_11332,N_11945);
nand U12189 (N_12189,N_11881,N_11355);
xnor U12190 (N_12190,N_11508,N_11824);
and U12191 (N_12191,N_11767,N_11743);
nand U12192 (N_12192,N_11330,N_11346);
nor U12193 (N_12193,N_11984,N_11619);
or U12194 (N_12194,N_11999,N_11868);
xor U12195 (N_12195,N_11312,N_11625);
or U12196 (N_12196,N_11343,N_11706);
nand U12197 (N_12197,N_11958,N_11313);
or U12198 (N_12198,N_11741,N_11909);
and U12199 (N_12199,N_11955,N_11812);
nand U12200 (N_12200,N_11378,N_11994);
and U12201 (N_12201,N_11495,N_11271);
nor U12202 (N_12202,N_11880,N_11421);
nor U12203 (N_12203,N_11364,N_11471);
nor U12204 (N_12204,N_11948,N_11816);
or U12205 (N_12205,N_11660,N_11989);
nand U12206 (N_12206,N_11831,N_11808);
xor U12207 (N_12207,N_11858,N_11273);
or U12208 (N_12208,N_11810,N_11737);
or U12209 (N_12209,N_11885,N_11608);
nor U12210 (N_12210,N_11975,N_11528);
nor U12211 (N_12211,N_11293,N_11573);
nor U12212 (N_12212,N_11878,N_11726);
xnor U12213 (N_12213,N_11775,N_11735);
xor U12214 (N_12214,N_11983,N_11497);
or U12215 (N_12215,N_11705,N_11261);
and U12216 (N_12216,N_11699,N_11492);
nor U12217 (N_12217,N_11940,N_11959);
or U12218 (N_12218,N_11865,N_11954);
xor U12219 (N_12219,N_11365,N_11928);
nor U12220 (N_12220,N_11733,N_11746);
and U12221 (N_12221,N_11973,N_11803);
nand U12222 (N_12222,N_11818,N_11838);
xor U12223 (N_12223,N_11266,N_11854);
nand U12224 (N_12224,N_11988,N_11814);
and U12225 (N_12225,N_11783,N_11450);
and U12226 (N_12226,N_11759,N_11915);
or U12227 (N_12227,N_11956,N_11262);
xnor U12228 (N_12228,N_11448,N_11863);
xnor U12229 (N_12229,N_11649,N_11690);
nor U12230 (N_12230,N_11623,N_11352);
nor U12231 (N_12231,N_11848,N_11621);
nor U12232 (N_12232,N_11577,N_11919);
xnor U12233 (N_12233,N_11484,N_11872);
or U12234 (N_12234,N_11892,N_11659);
xnor U12235 (N_12235,N_11551,N_11884);
nand U12236 (N_12236,N_11675,N_11857);
or U12237 (N_12237,N_11739,N_11996);
nor U12238 (N_12238,N_11442,N_11631);
and U12239 (N_12239,N_11584,N_11455);
xor U12240 (N_12240,N_11461,N_11467);
xnor U12241 (N_12241,N_11331,N_11289);
xor U12242 (N_12242,N_11635,N_11896);
or U12243 (N_12243,N_11452,N_11481);
nand U12244 (N_12244,N_11821,N_11908);
and U12245 (N_12245,N_11578,N_11505);
nor U12246 (N_12246,N_11285,N_11913);
or U12247 (N_12247,N_11263,N_11664);
nand U12248 (N_12248,N_11320,N_11786);
or U12249 (N_12249,N_11371,N_11925);
nand U12250 (N_12250,N_11304,N_11569);
or U12251 (N_12251,N_11341,N_11864);
nand U12252 (N_12252,N_11580,N_11693);
and U12253 (N_12253,N_11787,N_11682);
nand U12254 (N_12254,N_11763,N_11932);
or U12255 (N_12255,N_11254,N_11893);
nor U12256 (N_12256,N_11348,N_11671);
nand U12257 (N_12257,N_11494,N_11656);
nand U12258 (N_12258,N_11935,N_11265);
nand U12259 (N_12259,N_11469,N_11730);
and U12260 (N_12260,N_11618,N_11851);
nor U12261 (N_12261,N_11714,N_11986);
and U12262 (N_12262,N_11519,N_11833);
nand U12263 (N_12263,N_11687,N_11729);
or U12264 (N_12264,N_11257,N_11950);
nand U12265 (N_12265,N_11713,N_11354);
nor U12266 (N_12266,N_11793,N_11347);
and U12267 (N_12267,N_11903,N_11456);
nand U12268 (N_12268,N_11606,N_11611);
and U12269 (N_12269,N_11277,N_11616);
nor U12270 (N_12270,N_11437,N_11931);
or U12271 (N_12271,N_11888,N_11532);
or U12272 (N_12272,N_11867,N_11300);
and U12273 (N_12273,N_11895,N_11270);
and U12274 (N_12274,N_11546,N_11357);
or U12275 (N_12275,N_11264,N_11458);
nand U12276 (N_12276,N_11761,N_11666);
xnor U12277 (N_12277,N_11388,N_11842);
and U12278 (N_12278,N_11600,N_11587);
and U12279 (N_12279,N_11849,N_11531);
nor U12280 (N_12280,N_11256,N_11778);
nand U12281 (N_12281,N_11651,N_11911);
xor U12282 (N_12282,N_11680,N_11853);
xor U12283 (N_12283,N_11703,N_11556);
nor U12284 (N_12284,N_11772,N_11622);
xor U12285 (N_12285,N_11815,N_11795);
nand U12286 (N_12286,N_11859,N_11369);
nor U12287 (N_12287,N_11512,N_11957);
nor U12288 (N_12288,N_11335,N_11946);
nor U12289 (N_12289,N_11476,N_11610);
or U12290 (N_12290,N_11921,N_11789);
or U12291 (N_12291,N_11715,N_11882);
nor U12292 (N_12292,N_11373,N_11571);
and U12293 (N_12293,N_11941,N_11728);
xnor U12294 (N_12294,N_11443,N_11449);
and U12295 (N_12295,N_11738,N_11963);
or U12296 (N_12296,N_11678,N_11615);
nor U12297 (N_12297,N_11418,N_11933);
xor U12298 (N_12298,N_11446,N_11924);
xor U12299 (N_12299,N_11397,N_11555);
nor U12300 (N_12300,N_11712,N_11617);
or U12301 (N_12301,N_11288,N_11929);
nand U12302 (N_12302,N_11368,N_11695);
xnor U12303 (N_12303,N_11513,N_11483);
or U12304 (N_12304,N_11992,N_11298);
nor U12305 (N_12305,N_11964,N_11748);
and U12306 (N_12306,N_11472,N_11282);
or U12307 (N_12307,N_11459,N_11605);
nor U12308 (N_12308,N_11398,N_11589);
or U12309 (N_12309,N_11643,N_11688);
or U12310 (N_12310,N_11771,N_11407);
and U12311 (N_12311,N_11877,N_11303);
and U12312 (N_12312,N_11574,N_11905);
xnor U12313 (N_12313,N_11299,N_11827);
or U12314 (N_12314,N_11507,N_11788);
and U12315 (N_12315,N_11817,N_11275);
nand U12316 (N_12316,N_11408,N_11990);
and U12317 (N_12317,N_11511,N_11344);
xnor U12318 (N_12318,N_11549,N_11676);
nand U12319 (N_12319,N_11899,N_11679);
or U12320 (N_12320,N_11411,N_11939);
and U12321 (N_12321,N_11944,N_11460);
xor U12322 (N_12322,N_11278,N_11805);
nand U12323 (N_12323,N_11952,N_11314);
nor U12324 (N_12324,N_11425,N_11798);
xnor U12325 (N_12325,N_11719,N_11500);
xor U12326 (N_12326,N_11252,N_11807);
xnor U12327 (N_12327,N_11404,N_11979);
xnor U12328 (N_12328,N_11284,N_11390);
or U12329 (N_12329,N_11447,N_11698);
nand U12330 (N_12330,N_11843,N_11630);
nand U12331 (N_12331,N_11993,N_11785);
or U12332 (N_12332,N_11260,N_11581);
nor U12333 (N_12333,N_11604,N_11624);
nor U12334 (N_12334,N_11755,N_11326);
or U12335 (N_12335,N_11402,N_11438);
nand U12336 (N_12336,N_11837,N_11464);
xor U12337 (N_12337,N_11855,N_11370);
or U12338 (N_12338,N_11985,N_11395);
nor U12339 (N_12339,N_11781,N_11696);
and U12340 (N_12340,N_11349,N_11543);
or U12341 (N_12341,N_11436,N_11597);
nor U12342 (N_12342,N_11542,N_11272);
and U12343 (N_12343,N_11295,N_11525);
nand U12344 (N_12344,N_11424,N_11381);
or U12345 (N_12345,N_11538,N_11296);
or U12346 (N_12346,N_11860,N_11283);
xnor U12347 (N_12347,N_11750,N_11627);
xnor U12348 (N_12348,N_11478,N_11287);
or U12349 (N_12349,N_11393,N_11427);
nand U12350 (N_12350,N_11412,N_11613);
and U12351 (N_12351,N_11780,N_11841);
nor U12352 (N_12352,N_11520,N_11308);
or U12353 (N_12353,N_11379,N_11813);
xnor U12354 (N_12354,N_11943,N_11403);
nand U12355 (N_12355,N_11681,N_11653);
nor U12356 (N_12356,N_11593,N_11498);
and U12357 (N_12357,N_11871,N_11362);
xnor U12358 (N_12358,N_11804,N_11724);
and U12359 (N_12359,N_11850,N_11749);
and U12360 (N_12360,N_11490,N_11961);
nor U12361 (N_12361,N_11367,N_11897);
and U12362 (N_12362,N_11692,N_11353);
or U12363 (N_12363,N_11790,N_11392);
and U12364 (N_12364,N_11949,N_11752);
xnor U12365 (N_12365,N_11280,N_11998);
and U12366 (N_12366,N_11668,N_11599);
nand U12367 (N_12367,N_11826,N_11661);
nand U12368 (N_12368,N_11358,N_11325);
nand U12369 (N_12369,N_11250,N_11658);
and U12370 (N_12370,N_11912,N_11268);
and U12371 (N_12371,N_11267,N_11329);
nand U12372 (N_12372,N_11674,N_11526);
nand U12373 (N_12373,N_11968,N_11435);
or U12374 (N_12374,N_11316,N_11560);
nand U12375 (N_12375,N_11661,N_11295);
nor U12376 (N_12376,N_11995,N_11299);
nand U12377 (N_12377,N_11675,N_11384);
nor U12378 (N_12378,N_11546,N_11369);
xor U12379 (N_12379,N_11901,N_11767);
xnor U12380 (N_12380,N_11269,N_11652);
xor U12381 (N_12381,N_11254,N_11568);
nand U12382 (N_12382,N_11825,N_11832);
and U12383 (N_12383,N_11874,N_11490);
nand U12384 (N_12384,N_11429,N_11507);
or U12385 (N_12385,N_11611,N_11254);
nand U12386 (N_12386,N_11848,N_11262);
xnor U12387 (N_12387,N_11406,N_11747);
xor U12388 (N_12388,N_11914,N_11668);
nor U12389 (N_12389,N_11472,N_11454);
and U12390 (N_12390,N_11624,N_11597);
nand U12391 (N_12391,N_11288,N_11362);
and U12392 (N_12392,N_11989,N_11565);
nor U12393 (N_12393,N_11598,N_11954);
xor U12394 (N_12394,N_11775,N_11350);
and U12395 (N_12395,N_11423,N_11667);
and U12396 (N_12396,N_11270,N_11844);
or U12397 (N_12397,N_11262,N_11706);
nand U12398 (N_12398,N_11538,N_11977);
nor U12399 (N_12399,N_11718,N_11653);
xnor U12400 (N_12400,N_11503,N_11839);
xnor U12401 (N_12401,N_11861,N_11924);
xor U12402 (N_12402,N_11583,N_11397);
xor U12403 (N_12403,N_11730,N_11697);
nor U12404 (N_12404,N_11574,N_11513);
nor U12405 (N_12405,N_11324,N_11281);
nor U12406 (N_12406,N_11492,N_11666);
xor U12407 (N_12407,N_11644,N_11762);
nand U12408 (N_12408,N_11494,N_11431);
xor U12409 (N_12409,N_11483,N_11477);
xnor U12410 (N_12410,N_11949,N_11883);
xor U12411 (N_12411,N_11726,N_11783);
or U12412 (N_12412,N_11980,N_11926);
or U12413 (N_12413,N_11584,N_11569);
xor U12414 (N_12414,N_11546,N_11567);
xnor U12415 (N_12415,N_11621,N_11584);
nand U12416 (N_12416,N_11359,N_11908);
nor U12417 (N_12417,N_11296,N_11587);
nand U12418 (N_12418,N_11271,N_11533);
nand U12419 (N_12419,N_11751,N_11896);
nand U12420 (N_12420,N_11696,N_11577);
or U12421 (N_12421,N_11492,N_11522);
or U12422 (N_12422,N_11332,N_11853);
xnor U12423 (N_12423,N_11336,N_11894);
nand U12424 (N_12424,N_11287,N_11332);
nand U12425 (N_12425,N_11380,N_11384);
nor U12426 (N_12426,N_11361,N_11410);
xor U12427 (N_12427,N_11750,N_11703);
and U12428 (N_12428,N_11908,N_11296);
xnor U12429 (N_12429,N_11977,N_11717);
or U12430 (N_12430,N_11293,N_11479);
nand U12431 (N_12431,N_11375,N_11468);
nand U12432 (N_12432,N_11977,N_11922);
nor U12433 (N_12433,N_11371,N_11948);
or U12434 (N_12434,N_11503,N_11637);
xnor U12435 (N_12435,N_11947,N_11364);
and U12436 (N_12436,N_11730,N_11967);
or U12437 (N_12437,N_11417,N_11359);
nand U12438 (N_12438,N_11377,N_11517);
nor U12439 (N_12439,N_11798,N_11688);
or U12440 (N_12440,N_11801,N_11542);
xnor U12441 (N_12441,N_11926,N_11276);
and U12442 (N_12442,N_11910,N_11644);
and U12443 (N_12443,N_11515,N_11282);
xnor U12444 (N_12444,N_11381,N_11306);
nor U12445 (N_12445,N_11402,N_11918);
or U12446 (N_12446,N_11374,N_11397);
nor U12447 (N_12447,N_11358,N_11970);
and U12448 (N_12448,N_11415,N_11605);
and U12449 (N_12449,N_11645,N_11275);
nor U12450 (N_12450,N_11426,N_11589);
and U12451 (N_12451,N_11466,N_11477);
nor U12452 (N_12452,N_11912,N_11983);
or U12453 (N_12453,N_11449,N_11900);
nor U12454 (N_12454,N_11864,N_11255);
or U12455 (N_12455,N_11297,N_11387);
nor U12456 (N_12456,N_11533,N_11466);
nand U12457 (N_12457,N_11915,N_11756);
or U12458 (N_12458,N_11517,N_11933);
nand U12459 (N_12459,N_11308,N_11396);
nor U12460 (N_12460,N_11704,N_11711);
xnor U12461 (N_12461,N_11950,N_11827);
xnor U12462 (N_12462,N_11478,N_11907);
or U12463 (N_12463,N_11354,N_11861);
nand U12464 (N_12464,N_11334,N_11529);
xnor U12465 (N_12465,N_11396,N_11940);
nand U12466 (N_12466,N_11998,N_11497);
and U12467 (N_12467,N_11718,N_11812);
or U12468 (N_12468,N_11591,N_11341);
xnor U12469 (N_12469,N_11866,N_11457);
nand U12470 (N_12470,N_11433,N_11281);
nor U12471 (N_12471,N_11788,N_11567);
nor U12472 (N_12472,N_11696,N_11627);
nand U12473 (N_12473,N_11348,N_11913);
xnor U12474 (N_12474,N_11254,N_11370);
nor U12475 (N_12475,N_11722,N_11668);
nor U12476 (N_12476,N_11965,N_11851);
or U12477 (N_12477,N_11997,N_11252);
or U12478 (N_12478,N_11919,N_11293);
or U12479 (N_12479,N_11796,N_11269);
xor U12480 (N_12480,N_11364,N_11923);
xnor U12481 (N_12481,N_11540,N_11632);
nand U12482 (N_12482,N_11515,N_11977);
or U12483 (N_12483,N_11438,N_11299);
and U12484 (N_12484,N_11582,N_11533);
and U12485 (N_12485,N_11834,N_11577);
nor U12486 (N_12486,N_11420,N_11558);
nor U12487 (N_12487,N_11884,N_11627);
nand U12488 (N_12488,N_11409,N_11965);
xnor U12489 (N_12489,N_11456,N_11875);
xor U12490 (N_12490,N_11321,N_11680);
xor U12491 (N_12491,N_11750,N_11426);
xor U12492 (N_12492,N_11660,N_11662);
and U12493 (N_12493,N_11339,N_11304);
xnor U12494 (N_12494,N_11648,N_11874);
or U12495 (N_12495,N_11315,N_11965);
nor U12496 (N_12496,N_11543,N_11555);
xor U12497 (N_12497,N_11562,N_11316);
or U12498 (N_12498,N_11862,N_11960);
and U12499 (N_12499,N_11505,N_11924);
xnor U12500 (N_12500,N_11937,N_11960);
nand U12501 (N_12501,N_11840,N_11953);
nand U12502 (N_12502,N_11587,N_11837);
nor U12503 (N_12503,N_11369,N_11691);
nand U12504 (N_12504,N_11507,N_11344);
nor U12505 (N_12505,N_11353,N_11638);
xor U12506 (N_12506,N_11761,N_11681);
nand U12507 (N_12507,N_11581,N_11751);
nor U12508 (N_12508,N_11594,N_11685);
or U12509 (N_12509,N_11575,N_11679);
and U12510 (N_12510,N_11572,N_11834);
nor U12511 (N_12511,N_11854,N_11746);
or U12512 (N_12512,N_11924,N_11788);
nor U12513 (N_12513,N_11460,N_11620);
nor U12514 (N_12514,N_11682,N_11814);
or U12515 (N_12515,N_11874,N_11531);
xor U12516 (N_12516,N_11488,N_11481);
nand U12517 (N_12517,N_11280,N_11913);
and U12518 (N_12518,N_11466,N_11649);
nor U12519 (N_12519,N_11475,N_11366);
xor U12520 (N_12520,N_11649,N_11418);
nor U12521 (N_12521,N_11261,N_11522);
or U12522 (N_12522,N_11374,N_11265);
nand U12523 (N_12523,N_11654,N_11301);
or U12524 (N_12524,N_11299,N_11583);
or U12525 (N_12525,N_11469,N_11436);
nor U12526 (N_12526,N_11547,N_11326);
or U12527 (N_12527,N_11647,N_11321);
and U12528 (N_12528,N_11654,N_11744);
and U12529 (N_12529,N_11561,N_11898);
or U12530 (N_12530,N_11555,N_11845);
or U12531 (N_12531,N_11304,N_11390);
xnor U12532 (N_12532,N_11892,N_11793);
nor U12533 (N_12533,N_11805,N_11785);
xnor U12534 (N_12534,N_11623,N_11815);
or U12535 (N_12535,N_11311,N_11977);
and U12536 (N_12536,N_11571,N_11593);
xnor U12537 (N_12537,N_11430,N_11739);
nand U12538 (N_12538,N_11805,N_11464);
xor U12539 (N_12539,N_11337,N_11535);
and U12540 (N_12540,N_11530,N_11434);
or U12541 (N_12541,N_11465,N_11440);
and U12542 (N_12542,N_11824,N_11463);
or U12543 (N_12543,N_11258,N_11982);
nor U12544 (N_12544,N_11489,N_11690);
xor U12545 (N_12545,N_11538,N_11982);
and U12546 (N_12546,N_11552,N_11353);
nand U12547 (N_12547,N_11938,N_11950);
nand U12548 (N_12548,N_11847,N_11981);
nand U12549 (N_12549,N_11864,N_11742);
nand U12550 (N_12550,N_11545,N_11352);
nand U12551 (N_12551,N_11343,N_11963);
or U12552 (N_12552,N_11645,N_11732);
xor U12553 (N_12553,N_11959,N_11533);
or U12554 (N_12554,N_11277,N_11851);
and U12555 (N_12555,N_11741,N_11901);
nand U12556 (N_12556,N_11673,N_11607);
or U12557 (N_12557,N_11432,N_11305);
nor U12558 (N_12558,N_11798,N_11487);
or U12559 (N_12559,N_11704,N_11816);
and U12560 (N_12560,N_11416,N_11294);
or U12561 (N_12561,N_11948,N_11649);
nand U12562 (N_12562,N_11313,N_11261);
nor U12563 (N_12563,N_11793,N_11934);
and U12564 (N_12564,N_11781,N_11463);
nor U12565 (N_12565,N_11781,N_11869);
xnor U12566 (N_12566,N_11575,N_11664);
xnor U12567 (N_12567,N_11757,N_11266);
xnor U12568 (N_12568,N_11854,N_11434);
nand U12569 (N_12569,N_11476,N_11979);
and U12570 (N_12570,N_11390,N_11550);
nor U12571 (N_12571,N_11928,N_11512);
and U12572 (N_12572,N_11884,N_11819);
xor U12573 (N_12573,N_11990,N_11939);
nor U12574 (N_12574,N_11932,N_11857);
or U12575 (N_12575,N_11825,N_11638);
xor U12576 (N_12576,N_11619,N_11542);
xnor U12577 (N_12577,N_11411,N_11831);
nor U12578 (N_12578,N_11852,N_11662);
and U12579 (N_12579,N_11352,N_11256);
nor U12580 (N_12580,N_11529,N_11616);
xnor U12581 (N_12581,N_11472,N_11683);
and U12582 (N_12582,N_11849,N_11965);
xor U12583 (N_12583,N_11408,N_11728);
and U12584 (N_12584,N_11789,N_11931);
and U12585 (N_12585,N_11278,N_11877);
or U12586 (N_12586,N_11393,N_11331);
nand U12587 (N_12587,N_11553,N_11462);
and U12588 (N_12588,N_11371,N_11595);
xor U12589 (N_12589,N_11501,N_11732);
or U12590 (N_12590,N_11622,N_11336);
and U12591 (N_12591,N_11612,N_11689);
and U12592 (N_12592,N_11428,N_11818);
or U12593 (N_12593,N_11905,N_11928);
xnor U12594 (N_12594,N_11782,N_11993);
nand U12595 (N_12595,N_11284,N_11799);
and U12596 (N_12596,N_11909,N_11878);
xor U12597 (N_12597,N_11379,N_11938);
nor U12598 (N_12598,N_11554,N_11314);
and U12599 (N_12599,N_11294,N_11651);
nor U12600 (N_12600,N_11745,N_11458);
nor U12601 (N_12601,N_11400,N_11688);
xnor U12602 (N_12602,N_11269,N_11723);
xnor U12603 (N_12603,N_11815,N_11882);
xor U12604 (N_12604,N_11529,N_11976);
nor U12605 (N_12605,N_11715,N_11428);
xnor U12606 (N_12606,N_11666,N_11326);
xor U12607 (N_12607,N_11319,N_11779);
or U12608 (N_12608,N_11358,N_11415);
xor U12609 (N_12609,N_11293,N_11794);
or U12610 (N_12610,N_11596,N_11557);
or U12611 (N_12611,N_11267,N_11884);
or U12612 (N_12612,N_11323,N_11670);
and U12613 (N_12613,N_11343,N_11262);
or U12614 (N_12614,N_11378,N_11324);
xor U12615 (N_12615,N_11454,N_11677);
or U12616 (N_12616,N_11735,N_11668);
and U12617 (N_12617,N_11327,N_11979);
xor U12618 (N_12618,N_11848,N_11876);
and U12619 (N_12619,N_11675,N_11611);
and U12620 (N_12620,N_11945,N_11396);
or U12621 (N_12621,N_11312,N_11463);
xor U12622 (N_12622,N_11309,N_11992);
xor U12623 (N_12623,N_11871,N_11997);
or U12624 (N_12624,N_11493,N_11901);
xor U12625 (N_12625,N_11604,N_11332);
nor U12626 (N_12626,N_11880,N_11576);
and U12627 (N_12627,N_11880,N_11358);
or U12628 (N_12628,N_11415,N_11507);
or U12629 (N_12629,N_11819,N_11851);
nand U12630 (N_12630,N_11421,N_11424);
nand U12631 (N_12631,N_11335,N_11953);
or U12632 (N_12632,N_11724,N_11592);
xnor U12633 (N_12633,N_11520,N_11978);
or U12634 (N_12634,N_11258,N_11578);
and U12635 (N_12635,N_11783,N_11872);
xnor U12636 (N_12636,N_11709,N_11819);
or U12637 (N_12637,N_11824,N_11874);
or U12638 (N_12638,N_11924,N_11668);
nor U12639 (N_12639,N_11817,N_11356);
nor U12640 (N_12640,N_11440,N_11749);
or U12641 (N_12641,N_11624,N_11893);
and U12642 (N_12642,N_11255,N_11438);
nand U12643 (N_12643,N_11940,N_11675);
nor U12644 (N_12644,N_11657,N_11457);
nand U12645 (N_12645,N_11754,N_11471);
or U12646 (N_12646,N_11663,N_11342);
nor U12647 (N_12647,N_11800,N_11771);
nand U12648 (N_12648,N_11423,N_11981);
nor U12649 (N_12649,N_11878,N_11276);
nor U12650 (N_12650,N_11696,N_11617);
nand U12651 (N_12651,N_11788,N_11961);
or U12652 (N_12652,N_11600,N_11698);
nand U12653 (N_12653,N_11740,N_11478);
nor U12654 (N_12654,N_11440,N_11970);
xor U12655 (N_12655,N_11446,N_11774);
or U12656 (N_12656,N_11815,N_11983);
and U12657 (N_12657,N_11704,N_11883);
and U12658 (N_12658,N_11690,N_11822);
xnor U12659 (N_12659,N_11862,N_11832);
and U12660 (N_12660,N_11643,N_11652);
and U12661 (N_12661,N_11883,N_11760);
nor U12662 (N_12662,N_11913,N_11621);
nand U12663 (N_12663,N_11688,N_11744);
and U12664 (N_12664,N_11630,N_11440);
and U12665 (N_12665,N_11532,N_11536);
nor U12666 (N_12666,N_11669,N_11804);
and U12667 (N_12667,N_11306,N_11522);
nor U12668 (N_12668,N_11290,N_11657);
or U12669 (N_12669,N_11871,N_11952);
xnor U12670 (N_12670,N_11583,N_11700);
or U12671 (N_12671,N_11649,N_11345);
or U12672 (N_12672,N_11452,N_11547);
nor U12673 (N_12673,N_11742,N_11338);
xor U12674 (N_12674,N_11899,N_11359);
nor U12675 (N_12675,N_11555,N_11961);
and U12676 (N_12676,N_11575,N_11936);
nand U12677 (N_12677,N_11930,N_11958);
nor U12678 (N_12678,N_11373,N_11404);
xor U12679 (N_12679,N_11442,N_11928);
or U12680 (N_12680,N_11469,N_11841);
nor U12681 (N_12681,N_11605,N_11528);
nor U12682 (N_12682,N_11882,N_11820);
or U12683 (N_12683,N_11998,N_11877);
or U12684 (N_12684,N_11557,N_11979);
nor U12685 (N_12685,N_11537,N_11957);
or U12686 (N_12686,N_11982,N_11285);
or U12687 (N_12687,N_11422,N_11407);
nand U12688 (N_12688,N_11764,N_11892);
xor U12689 (N_12689,N_11383,N_11430);
and U12690 (N_12690,N_11967,N_11986);
nand U12691 (N_12691,N_11477,N_11981);
and U12692 (N_12692,N_11413,N_11617);
nor U12693 (N_12693,N_11703,N_11998);
xnor U12694 (N_12694,N_11594,N_11552);
or U12695 (N_12695,N_11663,N_11409);
nor U12696 (N_12696,N_11643,N_11440);
xnor U12697 (N_12697,N_11334,N_11966);
nand U12698 (N_12698,N_11401,N_11509);
xor U12699 (N_12699,N_11546,N_11356);
or U12700 (N_12700,N_11546,N_11670);
nor U12701 (N_12701,N_11378,N_11696);
or U12702 (N_12702,N_11868,N_11830);
xor U12703 (N_12703,N_11517,N_11922);
xor U12704 (N_12704,N_11997,N_11836);
xor U12705 (N_12705,N_11551,N_11636);
or U12706 (N_12706,N_11397,N_11553);
xor U12707 (N_12707,N_11372,N_11963);
nor U12708 (N_12708,N_11783,N_11420);
xnor U12709 (N_12709,N_11515,N_11605);
nor U12710 (N_12710,N_11949,N_11488);
and U12711 (N_12711,N_11637,N_11747);
and U12712 (N_12712,N_11662,N_11536);
nor U12713 (N_12713,N_11633,N_11439);
or U12714 (N_12714,N_11715,N_11599);
nand U12715 (N_12715,N_11931,N_11410);
nor U12716 (N_12716,N_11389,N_11443);
nor U12717 (N_12717,N_11773,N_11646);
nand U12718 (N_12718,N_11430,N_11641);
nand U12719 (N_12719,N_11673,N_11313);
and U12720 (N_12720,N_11348,N_11598);
nor U12721 (N_12721,N_11813,N_11608);
or U12722 (N_12722,N_11617,N_11918);
and U12723 (N_12723,N_11315,N_11555);
xnor U12724 (N_12724,N_11549,N_11548);
nand U12725 (N_12725,N_11748,N_11548);
nand U12726 (N_12726,N_11758,N_11357);
or U12727 (N_12727,N_11442,N_11703);
and U12728 (N_12728,N_11379,N_11731);
xnor U12729 (N_12729,N_11428,N_11667);
and U12730 (N_12730,N_11859,N_11550);
xnor U12731 (N_12731,N_11407,N_11379);
nor U12732 (N_12732,N_11455,N_11260);
nand U12733 (N_12733,N_11492,N_11441);
xnor U12734 (N_12734,N_11763,N_11783);
nor U12735 (N_12735,N_11616,N_11810);
xor U12736 (N_12736,N_11639,N_11917);
nor U12737 (N_12737,N_11594,N_11711);
nand U12738 (N_12738,N_11888,N_11302);
nor U12739 (N_12739,N_11381,N_11301);
or U12740 (N_12740,N_11796,N_11439);
nand U12741 (N_12741,N_11996,N_11892);
nand U12742 (N_12742,N_11781,N_11842);
nand U12743 (N_12743,N_11674,N_11664);
or U12744 (N_12744,N_11254,N_11873);
or U12745 (N_12745,N_11512,N_11876);
nand U12746 (N_12746,N_11565,N_11308);
and U12747 (N_12747,N_11339,N_11723);
nor U12748 (N_12748,N_11287,N_11701);
nand U12749 (N_12749,N_11561,N_11788);
nand U12750 (N_12750,N_12544,N_12603);
and U12751 (N_12751,N_12707,N_12389);
nand U12752 (N_12752,N_12106,N_12209);
or U12753 (N_12753,N_12672,N_12711);
nand U12754 (N_12754,N_12427,N_12325);
xnor U12755 (N_12755,N_12018,N_12240);
nor U12756 (N_12756,N_12673,N_12190);
and U12757 (N_12757,N_12744,N_12742);
nor U12758 (N_12758,N_12695,N_12599);
or U12759 (N_12759,N_12729,N_12355);
or U12760 (N_12760,N_12388,N_12456);
and U12761 (N_12761,N_12260,N_12386);
or U12762 (N_12762,N_12627,N_12368);
nor U12763 (N_12763,N_12741,N_12461);
or U12764 (N_12764,N_12358,N_12737);
nand U12765 (N_12765,N_12273,N_12490);
or U12766 (N_12766,N_12479,N_12526);
nor U12767 (N_12767,N_12558,N_12146);
xnor U12768 (N_12768,N_12020,N_12238);
xnor U12769 (N_12769,N_12195,N_12489);
nor U12770 (N_12770,N_12025,N_12044);
nand U12771 (N_12771,N_12323,N_12166);
nor U12772 (N_12772,N_12374,N_12118);
or U12773 (N_12773,N_12563,N_12459);
nand U12774 (N_12774,N_12621,N_12609);
or U12775 (N_12775,N_12727,N_12108);
nor U12776 (N_12776,N_12067,N_12442);
nand U12777 (N_12777,N_12587,N_12124);
nor U12778 (N_12778,N_12275,N_12411);
xor U12779 (N_12779,N_12600,N_12602);
xor U12780 (N_12780,N_12253,N_12441);
xnor U12781 (N_12781,N_12132,N_12364);
xnor U12782 (N_12782,N_12152,N_12467);
nor U12783 (N_12783,N_12568,N_12090);
or U12784 (N_12784,N_12213,N_12099);
nand U12785 (N_12785,N_12278,N_12197);
nand U12786 (N_12786,N_12270,N_12585);
or U12787 (N_12787,N_12538,N_12431);
xor U12788 (N_12788,N_12588,N_12282);
nor U12789 (N_12789,N_12159,N_12165);
or U12790 (N_12790,N_12307,N_12516);
xor U12791 (N_12791,N_12077,N_12685);
nor U12792 (N_12792,N_12066,N_12128);
and U12793 (N_12793,N_12652,N_12351);
or U12794 (N_12794,N_12206,N_12419);
and U12795 (N_12795,N_12092,N_12281);
nor U12796 (N_12796,N_12674,N_12300);
or U12797 (N_12797,N_12519,N_12584);
and U12798 (N_12798,N_12148,N_12367);
xnor U12799 (N_12799,N_12341,N_12085);
nor U12800 (N_12800,N_12503,N_12357);
nand U12801 (N_12801,N_12229,N_12175);
and U12802 (N_12802,N_12015,N_12384);
nor U12803 (N_12803,N_12397,N_12696);
xnor U12804 (N_12804,N_12342,N_12043);
nor U12805 (N_12805,N_12614,N_12518);
nand U12806 (N_12806,N_12523,N_12022);
xor U12807 (N_12807,N_12413,N_12064);
xnor U12808 (N_12808,N_12283,N_12626);
xor U12809 (N_12809,N_12036,N_12613);
or U12810 (N_12810,N_12595,N_12403);
xnor U12811 (N_12811,N_12482,N_12097);
or U12812 (N_12812,N_12458,N_12453);
nand U12813 (N_12813,N_12428,N_12701);
xnor U12814 (N_12814,N_12059,N_12514);
and U12815 (N_12815,N_12535,N_12537);
and U12816 (N_12816,N_12130,N_12002);
or U12817 (N_12817,N_12634,N_12034);
nor U12818 (N_12818,N_12623,N_12136);
nor U12819 (N_12819,N_12713,N_12566);
nand U12820 (N_12820,N_12414,N_12593);
or U12821 (N_12821,N_12265,N_12610);
nor U12822 (N_12822,N_12380,N_12030);
xnor U12823 (N_12823,N_12472,N_12122);
nor U12824 (N_12824,N_12725,N_12207);
nand U12825 (N_12825,N_12115,N_12455);
or U12826 (N_12826,N_12072,N_12271);
nand U12827 (N_12827,N_12668,N_12167);
and U12828 (N_12828,N_12259,N_12013);
nor U12829 (N_12829,N_12655,N_12338);
xnor U12830 (N_12830,N_12263,N_12163);
xor U12831 (N_12831,N_12572,N_12606);
or U12832 (N_12832,N_12199,N_12501);
nor U12833 (N_12833,N_12290,N_12079);
nor U12834 (N_12834,N_12356,N_12372);
and U12835 (N_12835,N_12645,N_12474);
and U12836 (N_12836,N_12087,N_12715);
and U12837 (N_12837,N_12109,N_12258);
and U12838 (N_12838,N_12399,N_12532);
xor U12839 (N_12839,N_12377,N_12716);
or U12840 (N_12840,N_12484,N_12636);
nor U12841 (N_12841,N_12415,N_12451);
or U12842 (N_12842,N_12352,N_12155);
nand U12843 (N_12843,N_12512,N_12447);
and U12844 (N_12844,N_12313,N_12202);
or U12845 (N_12845,N_12251,N_12590);
or U12846 (N_12846,N_12317,N_12511);
or U12847 (N_12847,N_12465,N_12050);
xnor U12848 (N_12848,N_12406,N_12549);
xor U12849 (N_12849,N_12158,N_12294);
and U12850 (N_12850,N_12344,N_12638);
xor U12851 (N_12851,N_12140,N_12346);
nand U12852 (N_12852,N_12131,N_12348);
nor U12853 (N_12853,N_12493,N_12049);
or U12854 (N_12854,N_12733,N_12252);
nand U12855 (N_12855,N_12042,N_12055);
nand U12856 (N_12856,N_12378,N_12021);
or U12857 (N_12857,N_12201,N_12745);
and U12858 (N_12858,N_12222,N_12463);
nor U12859 (N_12859,N_12683,N_12712);
nand U12860 (N_12860,N_12576,N_12095);
nand U12861 (N_12861,N_12394,N_12666);
and U12862 (N_12862,N_12284,N_12006);
and U12863 (N_12863,N_12464,N_12228);
and U12864 (N_12864,N_12226,N_12470);
or U12865 (N_12865,N_12533,N_12671);
or U12866 (N_12866,N_12393,N_12094);
or U12867 (N_12867,N_12429,N_12530);
nor U12868 (N_12868,N_12731,N_12524);
or U12869 (N_12869,N_12142,N_12506);
nand U12870 (N_12870,N_12723,N_12249);
nand U12871 (N_12871,N_12436,N_12345);
and U12872 (N_12872,N_12417,N_12738);
and U12873 (N_12873,N_12037,N_12257);
nand U12874 (N_12874,N_12350,N_12457);
or U12875 (N_12875,N_12440,N_12542);
and U12876 (N_12876,N_12041,N_12187);
nand U12877 (N_12877,N_12363,N_12365);
nor U12878 (N_12878,N_12204,N_12054);
xnor U12879 (N_12879,N_12646,N_12515);
nor U12880 (N_12880,N_12310,N_12242);
and U12881 (N_12881,N_12147,N_12183);
xnor U12882 (N_12882,N_12089,N_12302);
nand U12883 (N_12883,N_12071,N_12268);
or U12884 (N_12884,N_12560,N_12579);
nand U12885 (N_12885,N_12379,N_12214);
nor U12886 (N_12886,N_12293,N_12318);
nor U12887 (N_12887,N_12174,N_12589);
nor U12888 (N_12888,N_12382,N_12404);
xnor U12889 (N_12889,N_12091,N_12137);
or U12890 (N_12890,N_12297,N_12004);
and U12891 (N_12891,N_12211,N_12637);
xnor U12892 (N_12892,N_12126,N_12477);
and U12893 (N_12893,N_12121,N_12123);
or U12894 (N_12894,N_12694,N_12084);
xor U12895 (N_12895,N_12557,N_12076);
nor U12896 (N_12896,N_12179,N_12188);
nor U12897 (N_12897,N_12139,N_12320);
nor U12898 (N_12898,N_12279,N_12185);
or U12899 (N_12899,N_12517,N_12657);
nor U12900 (N_12900,N_12027,N_12040);
or U12901 (N_12901,N_12045,N_12150);
and U12902 (N_12902,N_12475,N_12728);
or U12903 (N_12903,N_12048,N_12616);
and U12904 (N_12904,N_12105,N_12628);
and U12905 (N_12905,N_12507,N_12629);
nand U12906 (N_12906,N_12522,N_12019);
xnor U12907 (N_12907,N_12462,N_12193);
or U12908 (N_12908,N_12541,N_12141);
nor U12909 (N_12909,N_12697,N_12651);
nand U12910 (N_12910,N_12432,N_12687);
and U12911 (N_12911,N_12486,N_12650);
nand U12912 (N_12912,N_12420,N_12395);
or U12913 (N_12913,N_12662,N_12385);
xor U12914 (N_12914,N_12660,N_12497);
xnor U12915 (N_12915,N_12722,N_12081);
nor U12916 (N_12916,N_12096,N_12144);
and U12917 (N_12917,N_12306,N_12513);
xnor U12918 (N_12918,N_12192,N_12704);
or U12919 (N_12919,N_12292,N_12008);
nand U12920 (N_12920,N_12012,N_12033);
and U12921 (N_12921,N_12031,N_12659);
or U12922 (N_12922,N_12700,N_12418);
or U12923 (N_12923,N_12369,N_12658);
or U12924 (N_12924,N_12303,N_12254);
or U12925 (N_12925,N_12653,N_12597);
or U12926 (N_12926,N_12443,N_12119);
nor U12927 (N_12927,N_12581,N_12721);
nor U12928 (N_12928,N_12264,N_12127);
or U12929 (N_12929,N_12011,N_12161);
nand U12930 (N_12930,N_12028,N_12110);
nand U12931 (N_12931,N_12112,N_12277);
and U12932 (N_12932,N_12422,N_12145);
or U12933 (N_12933,N_12434,N_12505);
nand U12934 (N_12934,N_12000,N_12334);
or U12935 (N_12935,N_12649,N_12408);
nor U12936 (N_12936,N_12337,N_12304);
nor U12937 (N_12937,N_12104,N_12604);
or U12938 (N_12938,N_12746,N_12133);
and U12939 (N_12939,N_12619,N_12003);
or U12940 (N_12940,N_12551,N_12135);
nor U12941 (N_12941,N_12327,N_12691);
xor U12942 (N_12942,N_12156,N_12200);
or U12943 (N_12943,N_12117,N_12340);
nand U12944 (N_12944,N_12499,N_12680);
nor U12945 (N_12945,N_12101,N_12615);
and U12946 (N_12946,N_12171,N_12564);
or U12947 (N_12947,N_12640,N_12439);
or U12948 (N_12948,N_12682,N_12098);
or U12949 (N_12949,N_12578,N_12164);
xor U12950 (N_12950,N_12366,N_12433);
and U12951 (N_12951,N_12539,N_12631);
nand U12952 (N_12952,N_12485,N_12308);
nor U12953 (N_12953,N_12329,N_12509);
xnor U12954 (N_12954,N_12218,N_12483);
and U12955 (N_12955,N_12577,N_12138);
xor U12956 (N_12956,N_12359,N_12491);
and U12957 (N_12957,N_12675,N_12469);
nor U12958 (N_12958,N_12232,N_12567);
xnor U12959 (N_12959,N_12245,N_12113);
xnor U12960 (N_12960,N_12702,N_12035);
or U12961 (N_12961,N_12014,N_12051);
nor U12962 (N_12962,N_12452,N_12740);
nand U12963 (N_12963,N_12029,N_12219);
and U12964 (N_12964,N_12169,N_12554);
nand U12965 (N_12965,N_12339,N_12500);
xnor U12966 (N_12966,N_12208,N_12714);
and U12967 (N_12967,N_12748,N_12416);
nand U12968 (N_12968,N_12052,N_12561);
nor U12969 (N_12969,N_12719,N_12319);
and U12970 (N_12970,N_12726,N_12371);
nor U12971 (N_12971,N_12543,N_12047);
or U12972 (N_12972,N_12559,N_12210);
and U12973 (N_12973,N_12227,N_12749);
or U12974 (N_12974,N_12056,N_12068);
nor U12975 (N_12975,N_12181,N_12468);
nand U12976 (N_12976,N_12445,N_12592);
nand U12977 (N_12977,N_12335,N_12625);
xor U12978 (N_12978,N_12534,N_12699);
or U12979 (N_12979,N_12550,N_12070);
xnor U12980 (N_12980,N_12178,N_12693);
xnor U12981 (N_12981,N_12060,N_12032);
or U12982 (N_12982,N_12120,N_12446);
nand U12983 (N_12983,N_12409,N_12556);
xor U12984 (N_12984,N_12648,N_12663);
xnor U12985 (N_12985,N_12360,N_12487);
and U12986 (N_12986,N_12669,N_12476);
and U12987 (N_12987,N_12521,N_12423);
and U12988 (N_12988,N_12644,N_12225);
and U12989 (N_12989,N_12312,N_12250);
xor U12990 (N_12990,N_12678,N_12046);
nand U12991 (N_12991,N_12189,N_12009);
xnor U12992 (N_12992,N_12633,N_12296);
and U12993 (N_12993,N_12545,N_12703);
and U12994 (N_12994,N_12495,N_12286);
nor U12995 (N_12995,N_12361,N_12168);
nand U12996 (N_12996,N_12488,N_12665);
or U12997 (N_12997,N_12692,N_12480);
or U12998 (N_12998,N_12449,N_12058);
or U12999 (N_12999,N_12582,N_12654);
xnor U13000 (N_13000,N_12311,N_12336);
or U13001 (N_13001,N_12315,N_12546);
and U13002 (N_13002,N_12435,N_12362);
and U13003 (N_13003,N_12698,N_12053);
xor U13004 (N_13004,N_12093,N_12285);
nor U13005 (N_13005,N_12580,N_12233);
xnor U13006 (N_13006,N_12223,N_12343);
xnor U13007 (N_13007,N_12583,N_12314);
xor U13008 (N_13008,N_12412,N_12017);
and U13009 (N_13009,N_12402,N_12262);
nor U13010 (N_13010,N_12024,N_12180);
nand U13011 (N_13011,N_12689,N_12272);
and U13012 (N_13012,N_12005,N_12743);
and U13013 (N_13013,N_12016,N_12157);
nand U13014 (N_13014,N_12073,N_12732);
nor U13015 (N_13015,N_12437,N_12617);
nand U13016 (N_13016,N_12287,N_12276);
xor U13017 (N_13017,N_12129,N_12591);
nand U13018 (N_13018,N_12291,N_12639);
and U13019 (N_13019,N_12390,N_12607);
nand U13020 (N_13020,N_12620,N_12596);
and U13021 (N_13021,N_12221,N_12570);
xnor U13022 (N_13022,N_12494,N_12224);
xnor U13023 (N_13023,N_12326,N_12706);
and U13024 (N_13024,N_12205,N_12736);
nor U13025 (N_13025,N_12574,N_12065);
or U13026 (N_13026,N_12594,N_12237);
nor U13027 (N_13027,N_12642,N_12547);
and U13028 (N_13028,N_12234,N_12734);
or U13029 (N_13029,N_12527,N_12410);
or U13030 (N_13030,N_12216,N_12632);
xnor U13031 (N_13031,N_12392,N_12316);
and U13032 (N_13032,N_12198,N_12280);
nand U13033 (N_13033,N_12375,N_12170);
or U13034 (N_13034,N_12667,N_12063);
xnor U13035 (N_13035,N_12421,N_12010);
and U13036 (N_13036,N_12575,N_12353);
xnor U13037 (N_13037,N_12154,N_12391);
nand U13038 (N_13038,N_12062,N_12215);
xor U13039 (N_13039,N_12618,N_12239);
and U13040 (N_13040,N_12525,N_12075);
nand U13041 (N_13041,N_12681,N_12705);
nand U13042 (N_13042,N_12424,N_12730);
and U13043 (N_13043,N_12354,N_12540);
nor U13044 (N_13044,N_12641,N_12177);
nand U13045 (N_13045,N_12153,N_12330);
and U13046 (N_13046,N_12332,N_12677);
nand U13047 (N_13047,N_12688,N_12196);
nor U13048 (N_13048,N_12194,N_12502);
or U13049 (N_13049,N_12686,N_12114);
xnor U13050 (N_13050,N_12478,N_12266);
nand U13051 (N_13051,N_12038,N_12598);
nor U13052 (N_13052,N_12498,N_12396);
or U13053 (N_13053,N_12690,N_12548);
xnor U13054 (N_13054,N_12407,N_12039);
xnor U13055 (N_13055,N_12160,N_12536);
or U13056 (N_13056,N_12529,N_12611);
xnor U13057 (N_13057,N_12612,N_12710);
nand U13058 (N_13058,N_12309,N_12444);
xnor U13059 (N_13059,N_12496,N_12643);
nor U13060 (N_13060,N_12608,N_12247);
and U13061 (N_13061,N_12088,N_12471);
or U13062 (N_13062,N_12684,N_12508);
or U13063 (N_13063,N_12565,N_12082);
nor U13064 (N_13064,N_12670,N_12492);
nand U13065 (N_13065,N_12173,N_12107);
and U13066 (N_13066,N_12069,N_12001);
nand U13067 (N_13067,N_12601,N_12256);
or U13068 (N_13068,N_12747,N_12605);
nor U13069 (N_13069,N_12301,N_12400);
and U13070 (N_13070,N_12724,N_12274);
nand U13071 (N_13071,N_12269,N_12676);
nand U13072 (N_13072,N_12405,N_12562);
nor U13073 (N_13073,N_12246,N_12255);
nand U13074 (N_13074,N_12381,N_12241);
nand U13075 (N_13075,N_12708,N_12217);
and U13076 (N_13076,N_12116,N_12295);
or U13077 (N_13077,N_12387,N_12347);
and U13078 (N_13078,N_12647,N_12026);
or U13079 (N_13079,N_12134,N_12236);
nand U13080 (N_13080,N_12331,N_12555);
and U13081 (N_13081,N_12438,N_12324);
xor U13082 (N_13082,N_12305,N_12635);
nand U13083 (N_13083,N_12454,N_12383);
xor U13084 (N_13084,N_12718,N_12373);
xor U13085 (N_13085,N_12078,N_12086);
nor U13086 (N_13086,N_12267,N_12074);
nand U13087 (N_13087,N_12007,N_12466);
and U13088 (N_13088,N_12661,N_12573);
nand U13089 (N_13089,N_12630,N_12664);
xor U13090 (N_13090,N_12481,N_12230);
xor U13091 (N_13091,N_12244,N_12151);
xnor U13092 (N_13092,N_12111,N_12261);
or U13093 (N_13093,N_12231,N_12656);
and U13094 (N_13094,N_12298,N_12125);
xor U13095 (N_13095,N_12735,N_12100);
or U13096 (N_13096,N_12328,N_12520);
nand U13097 (N_13097,N_12401,N_12288);
nand U13098 (N_13098,N_12709,N_12510);
xnor U13099 (N_13099,N_12426,N_12176);
or U13100 (N_13100,N_12624,N_12191);
or U13101 (N_13101,N_12553,N_12184);
nand U13102 (N_13102,N_12448,N_12289);
nand U13103 (N_13103,N_12203,N_12430);
nor U13104 (N_13104,N_12182,N_12023);
or U13105 (N_13105,N_12235,N_12586);
or U13106 (N_13106,N_12552,N_12299);
and U13107 (N_13107,N_12149,N_12739);
xnor U13108 (N_13108,N_12370,N_12425);
or U13109 (N_13109,N_12162,N_12569);
and U13110 (N_13110,N_12504,N_12186);
xnor U13111 (N_13111,N_12102,N_12143);
nor U13112 (N_13112,N_12720,N_12248);
xnor U13113 (N_13113,N_12717,N_12061);
nor U13114 (N_13114,N_12322,N_12460);
nor U13115 (N_13115,N_12398,N_12531);
and U13116 (N_13116,N_12333,N_12571);
nor U13117 (N_13117,N_12220,N_12528);
nor U13118 (N_13118,N_12103,N_12450);
nor U13119 (N_13119,N_12376,N_12349);
and U13120 (N_13120,N_12321,N_12057);
and U13121 (N_13121,N_12679,N_12622);
xor U13122 (N_13122,N_12080,N_12172);
nor U13123 (N_13123,N_12212,N_12243);
xor U13124 (N_13124,N_12473,N_12083);
or U13125 (N_13125,N_12680,N_12395);
nand U13126 (N_13126,N_12716,N_12291);
or U13127 (N_13127,N_12223,N_12658);
nand U13128 (N_13128,N_12348,N_12608);
or U13129 (N_13129,N_12470,N_12314);
nand U13130 (N_13130,N_12063,N_12257);
or U13131 (N_13131,N_12605,N_12192);
and U13132 (N_13132,N_12316,N_12402);
or U13133 (N_13133,N_12348,N_12178);
xnor U13134 (N_13134,N_12376,N_12719);
or U13135 (N_13135,N_12052,N_12268);
nor U13136 (N_13136,N_12034,N_12214);
or U13137 (N_13137,N_12450,N_12135);
xnor U13138 (N_13138,N_12702,N_12045);
and U13139 (N_13139,N_12169,N_12674);
or U13140 (N_13140,N_12453,N_12209);
or U13141 (N_13141,N_12409,N_12480);
and U13142 (N_13142,N_12369,N_12442);
nand U13143 (N_13143,N_12311,N_12675);
nor U13144 (N_13144,N_12035,N_12401);
xor U13145 (N_13145,N_12284,N_12392);
xnor U13146 (N_13146,N_12499,N_12407);
and U13147 (N_13147,N_12088,N_12598);
xor U13148 (N_13148,N_12181,N_12659);
or U13149 (N_13149,N_12346,N_12227);
and U13150 (N_13150,N_12104,N_12316);
xor U13151 (N_13151,N_12115,N_12376);
nand U13152 (N_13152,N_12320,N_12093);
or U13153 (N_13153,N_12085,N_12361);
nand U13154 (N_13154,N_12336,N_12563);
nand U13155 (N_13155,N_12203,N_12431);
or U13156 (N_13156,N_12241,N_12475);
nand U13157 (N_13157,N_12355,N_12649);
nor U13158 (N_13158,N_12005,N_12305);
xor U13159 (N_13159,N_12556,N_12301);
and U13160 (N_13160,N_12746,N_12481);
xnor U13161 (N_13161,N_12447,N_12159);
or U13162 (N_13162,N_12545,N_12472);
and U13163 (N_13163,N_12310,N_12631);
or U13164 (N_13164,N_12212,N_12013);
xnor U13165 (N_13165,N_12429,N_12410);
and U13166 (N_13166,N_12511,N_12627);
nor U13167 (N_13167,N_12125,N_12590);
or U13168 (N_13168,N_12579,N_12402);
nor U13169 (N_13169,N_12272,N_12584);
or U13170 (N_13170,N_12060,N_12654);
or U13171 (N_13171,N_12484,N_12235);
nand U13172 (N_13172,N_12660,N_12087);
nor U13173 (N_13173,N_12621,N_12341);
xnor U13174 (N_13174,N_12196,N_12258);
and U13175 (N_13175,N_12296,N_12716);
and U13176 (N_13176,N_12129,N_12687);
xnor U13177 (N_13177,N_12088,N_12219);
nand U13178 (N_13178,N_12723,N_12347);
nand U13179 (N_13179,N_12271,N_12745);
nand U13180 (N_13180,N_12061,N_12271);
xor U13181 (N_13181,N_12354,N_12356);
and U13182 (N_13182,N_12625,N_12197);
xor U13183 (N_13183,N_12252,N_12014);
nand U13184 (N_13184,N_12212,N_12347);
or U13185 (N_13185,N_12689,N_12268);
or U13186 (N_13186,N_12209,N_12080);
nor U13187 (N_13187,N_12522,N_12447);
nand U13188 (N_13188,N_12004,N_12215);
and U13189 (N_13189,N_12500,N_12651);
or U13190 (N_13190,N_12491,N_12479);
or U13191 (N_13191,N_12613,N_12033);
xor U13192 (N_13192,N_12642,N_12523);
and U13193 (N_13193,N_12322,N_12666);
nor U13194 (N_13194,N_12205,N_12212);
nand U13195 (N_13195,N_12468,N_12747);
nor U13196 (N_13196,N_12086,N_12534);
and U13197 (N_13197,N_12614,N_12156);
and U13198 (N_13198,N_12016,N_12364);
nor U13199 (N_13199,N_12741,N_12377);
and U13200 (N_13200,N_12083,N_12062);
nor U13201 (N_13201,N_12307,N_12063);
nor U13202 (N_13202,N_12416,N_12715);
nor U13203 (N_13203,N_12342,N_12582);
nand U13204 (N_13204,N_12367,N_12084);
nand U13205 (N_13205,N_12181,N_12141);
or U13206 (N_13206,N_12526,N_12138);
or U13207 (N_13207,N_12735,N_12064);
nor U13208 (N_13208,N_12746,N_12199);
nand U13209 (N_13209,N_12161,N_12348);
xor U13210 (N_13210,N_12326,N_12085);
and U13211 (N_13211,N_12018,N_12116);
xnor U13212 (N_13212,N_12164,N_12708);
nor U13213 (N_13213,N_12178,N_12562);
xor U13214 (N_13214,N_12423,N_12524);
xor U13215 (N_13215,N_12478,N_12041);
xnor U13216 (N_13216,N_12711,N_12440);
or U13217 (N_13217,N_12393,N_12355);
and U13218 (N_13218,N_12648,N_12439);
and U13219 (N_13219,N_12605,N_12004);
nor U13220 (N_13220,N_12241,N_12480);
xnor U13221 (N_13221,N_12576,N_12333);
xor U13222 (N_13222,N_12151,N_12499);
or U13223 (N_13223,N_12472,N_12406);
or U13224 (N_13224,N_12411,N_12079);
nor U13225 (N_13225,N_12393,N_12652);
and U13226 (N_13226,N_12703,N_12063);
or U13227 (N_13227,N_12696,N_12557);
or U13228 (N_13228,N_12627,N_12355);
nor U13229 (N_13229,N_12625,N_12188);
and U13230 (N_13230,N_12175,N_12248);
xnor U13231 (N_13231,N_12317,N_12721);
nand U13232 (N_13232,N_12342,N_12421);
and U13233 (N_13233,N_12548,N_12336);
nand U13234 (N_13234,N_12491,N_12622);
xnor U13235 (N_13235,N_12120,N_12306);
or U13236 (N_13236,N_12494,N_12189);
and U13237 (N_13237,N_12502,N_12217);
nor U13238 (N_13238,N_12674,N_12268);
nand U13239 (N_13239,N_12332,N_12748);
nor U13240 (N_13240,N_12682,N_12733);
nor U13241 (N_13241,N_12209,N_12626);
xor U13242 (N_13242,N_12595,N_12098);
and U13243 (N_13243,N_12422,N_12454);
nand U13244 (N_13244,N_12741,N_12573);
nand U13245 (N_13245,N_12039,N_12501);
and U13246 (N_13246,N_12067,N_12165);
nand U13247 (N_13247,N_12138,N_12428);
xor U13248 (N_13248,N_12219,N_12031);
xor U13249 (N_13249,N_12310,N_12532);
nor U13250 (N_13250,N_12526,N_12028);
nor U13251 (N_13251,N_12009,N_12330);
or U13252 (N_13252,N_12456,N_12557);
nand U13253 (N_13253,N_12363,N_12231);
and U13254 (N_13254,N_12088,N_12639);
or U13255 (N_13255,N_12439,N_12353);
and U13256 (N_13256,N_12188,N_12691);
nor U13257 (N_13257,N_12277,N_12123);
nand U13258 (N_13258,N_12175,N_12680);
nor U13259 (N_13259,N_12027,N_12713);
nor U13260 (N_13260,N_12148,N_12006);
xnor U13261 (N_13261,N_12090,N_12110);
nor U13262 (N_13262,N_12309,N_12650);
and U13263 (N_13263,N_12158,N_12469);
and U13264 (N_13264,N_12058,N_12682);
xnor U13265 (N_13265,N_12176,N_12257);
or U13266 (N_13266,N_12403,N_12419);
or U13267 (N_13267,N_12713,N_12701);
nor U13268 (N_13268,N_12159,N_12606);
nand U13269 (N_13269,N_12130,N_12447);
nand U13270 (N_13270,N_12622,N_12314);
xor U13271 (N_13271,N_12438,N_12056);
or U13272 (N_13272,N_12216,N_12271);
or U13273 (N_13273,N_12228,N_12524);
nand U13274 (N_13274,N_12671,N_12714);
or U13275 (N_13275,N_12619,N_12161);
or U13276 (N_13276,N_12162,N_12699);
nor U13277 (N_13277,N_12529,N_12737);
xor U13278 (N_13278,N_12011,N_12066);
or U13279 (N_13279,N_12657,N_12307);
and U13280 (N_13280,N_12251,N_12672);
xnor U13281 (N_13281,N_12542,N_12172);
nand U13282 (N_13282,N_12183,N_12658);
or U13283 (N_13283,N_12558,N_12740);
and U13284 (N_13284,N_12674,N_12367);
nor U13285 (N_13285,N_12157,N_12596);
xor U13286 (N_13286,N_12179,N_12612);
or U13287 (N_13287,N_12338,N_12053);
and U13288 (N_13288,N_12539,N_12345);
xor U13289 (N_13289,N_12270,N_12596);
xor U13290 (N_13290,N_12599,N_12252);
nand U13291 (N_13291,N_12276,N_12074);
nand U13292 (N_13292,N_12345,N_12428);
or U13293 (N_13293,N_12154,N_12539);
nand U13294 (N_13294,N_12243,N_12223);
and U13295 (N_13295,N_12069,N_12308);
xor U13296 (N_13296,N_12394,N_12090);
nand U13297 (N_13297,N_12509,N_12351);
and U13298 (N_13298,N_12426,N_12462);
xor U13299 (N_13299,N_12517,N_12337);
or U13300 (N_13300,N_12694,N_12591);
or U13301 (N_13301,N_12196,N_12723);
nand U13302 (N_13302,N_12576,N_12658);
xor U13303 (N_13303,N_12083,N_12517);
xor U13304 (N_13304,N_12233,N_12016);
nor U13305 (N_13305,N_12333,N_12037);
nand U13306 (N_13306,N_12568,N_12746);
xnor U13307 (N_13307,N_12074,N_12445);
nand U13308 (N_13308,N_12685,N_12714);
xor U13309 (N_13309,N_12400,N_12025);
xnor U13310 (N_13310,N_12051,N_12510);
xor U13311 (N_13311,N_12251,N_12708);
and U13312 (N_13312,N_12394,N_12592);
and U13313 (N_13313,N_12088,N_12336);
or U13314 (N_13314,N_12628,N_12425);
and U13315 (N_13315,N_12186,N_12346);
or U13316 (N_13316,N_12178,N_12016);
nand U13317 (N_13317,N_12580,N_12069);
or U13318 (N_13318,N_12465,N_12693);
or U13319 (N_13319,N_12195,N_12430);
nand U13320 (N_13320,N_12283,N_12683);
nand U13321 (N_13321,N_12270,N_12257);
and U13322 (N_13322,N_12008,N_12380);
and U13323 (N_13323,N_12073,N_12728);
nand U13324 (N_13324,N_12301,N_12463);
and U13325 (N_13325,N_12335,N_12441);
and U13326 (N_13326,N_12221,N_12148);
nand U13327 (N_13327,N_12524,N_12655);
or U13328 (N_13328,N_12081,N_12445);
or U13329 (N_13329,N_12651,N_12359);
xnor U13330 (N_13330,N_12590,N_12381);
nor U13331 (N_13331,N_12397,N_12143);
nand U13332 (N_13332,N_12491,N_12340);
nor U13333 (N_13333,N_12511,N_12255);
nor U13334 (N_13334,N_12342,N_12558);
and U13335 (N_13335,N_12195,N_12302);
nor U13336 (N_13336,N_12417,N_12635);
xnor U13337 (N_13337,N_12404,N_12344);
or U13338 (N_13338,N_12149,N_12022);
or U13339 (N_13339,N_12446,N_12682);
nand U13340 (N_13340,N_12283,N_12726);
nand U13341 (N_13341,N_12328,N_12700);
nor U13342 (N_13342,N_12187,N_12080);
nand U13343 (N_13343,N_12391,N_12627);
xor U13344 (N_13344,N_12349,N_12022);
nand U13345 (N_13345,N_12376,N_12577);
or U13346 (N_13346,N_12396,N_12163);
nand U13347 (N_13347,N_12122,N_12161);
and U13348 (N_13348,N_12740,N_12242);
nand U13349 (N_13349,N_12709,N_12015);
or U13350 (N_13350,N_12066,N_12509);
nor U13351 (N_13351,N_12652,N_12649);
nor U13352 (N_13352,N_12134,N_12638);
or U13353 (N_13353,N_12279,N_12067);
nor U13354 (N_13354,N_12291,N_12528);
nor U13355 (N_13355,N_12727,N_12244);
and U13356 (N_13356,N_12560,N_12385);
and U13357 (N_13357,N_12289,N_12554);
nand U13358 (N_13358,N_12095,N_12426);
xnor U13359 (N_13359,N_12528,N_12732);
xor U13360 (N_13360,N_12605,N_12387);
or U13361 (N_13361,N_12483,N_12676);
xor U13362 (N_13362,N_12296,N_12147);
nor U13363 (N_13363,N_12617,N_12741);
xnor U13364 (N_13364,N_12246,N_12311);
nand U13365 (N_13365,N_12413,N_12659);
nor U13366 (N_13366,N_12171,N_12121);
nand U13367 (N_13367,N_12349,N_12335);
and U13368 (N_13368,N_12230,N_12484);
nor U13369 (N_13369,N_12231,N_12089);
xor U13370 (N_13370,N_12311,N_12252);
or U13371 (N_13371,N_12016,N_12348);
or U13372 (N_13372,N_12098,N_12597);
or U13373 (N_13373,N_12644,N_12471);
nor U13374 (N_13374,N_12309,N_12655);
xor U13375 (N_13375,N_12649,N_12310);
or U13376 (N_13376,N_12423,N_12425);
nor U13377 (N_13377,N_12090,N_12451);
nand U13378 (N_13378,N_12683,N_12367);
xnor U13379 (N_13379,N_12364,N_12679);
and U13380 (N_13380,N_12224,N_12420);
xor U13381 (N_13381,N_12311,N_12610);
xnor U13382 (N_13382,N_12339,N_12123);
and U13383 (N_13383,N_12546,N_12000);
or U13384 (N_13384,N_12348,N_12106);
nand U13385 (N_13385,N_12446,N_12228);
xnor U13386 (N_13386,N_12229,N_12442);
and U13387 (N_13387,N_12294,N_12424);
and U13388 (N_13388,N_12267,N_12212);
nand U13389 (N_13389,N_12033,N_12403);
nor U13390 (N_13390,N_12698,N_12373);
or U13391 (N_13391,N_12504,N_12628);
and U13392 (N_13392,N_12292,N_12236);
nor U13393 (N_13393,N_12525,N_12744);
and U13394 (N_13394,N_12598,N_12149);
or U13395 (N_13395,N_12229,N_12366);
xor U13396 (N_13396,N_12478,N_12663);
xor U13397 (N_13397,N_12654,N_12634);
xnor U13398 (N_13398,N_12319,N_12426);
nor U13399 (N_13399,N_12588,N_12598);
or U13400 (N_13400,N_12296,N_12176);
xor U13401 (N_13401,N_12041,N_12503);
nand U13402 (N_13402,N_12093,N_12275);
nor U13403 (N_13403,N_12413,N_12669);
nand U13404 (N_13404,N_12552,N_12423);
xnor U13405 (N_13405,N_12657,N_12093);
xnor U13406 (N_13406,N_12064,N_12153);
nor U13407 (N_13407,N_12691,N_12707);
nor U13408 (N_13408,N_12544,N_12657);
or U13409 (N_13409,N_12511,N_12030);
and U13410 (N_13410,N_12738,N_12310);
or U13411 (N_13411,N_12130,N_12363);
and U13412 (N_13412,N_12548,N_12713);
and U13413 (N_13413,N_12327,N_12067);
xor U13414 (N_13414,N_12633,N_12438);
and U13415 (N_13415,N_12581,N_12701);
or U13416 (N_13416,N_12527,N_12605);
xnor U13417 (N_13417,N_12119,N_12508);
or U13418 (N_13418,N_12486,N_12591);
and U13419 (N_13419,N_12355,N_12427);
or U13420 (N_13420,N_12493,N_12485);
or U13421 (N_13421,N_12453,N_12388);
xor U13422 (N_13422,N_12283,N_12252);
or U13423 (N_13423,N_12274,N_12583);
nand U13424 (N_13424,N_12271,N_12251);
nor U13425 (N_13425,N_12517,N_12104);
nor U13426 (N_13426,N_12223,N_12447);
xnor U13427 (N_13427,N_12077,N_12003);
nand U13428 (N_13428,N_12316,N_12208);
or U13429 (N_13429,N_12034,N_12627);
nand U13430 (N_13430,N_12117,N_12749);
nor U13431 (N_13431,N_12522,N_12155);
nor U13432 (N_13432,N_12714,N_12653);
or U13433 (N_13433,N_12106,N_12001);
xnor U13434 (N_13434,N_12110,N_12475);
nor U13435 (N_13435,N_12631,N_12707);
and U13436 (N_13436,N_12643,N_12432);
or U13437 (N_13437,N_12075,N_12703);
or U13438 (N_13438,N_12200,N_12382);
xnor U13439 (N_13439,N_12598,N_12562);
nor U13440 (N_13440,N_12135,N_12591);
or U13441 (N_13441,N_12226,N_12302);
nor U13442 (N_13442,N_12691,N_12138);
and U13443 (N_13443,N_12187,N_12268);
nand U13444 (N_13444,N_12325,N_12730);
nand U13445 (N_13445,N_12642,N_12527);
and U13446 (N_13446,N_12743,N_12089);
nand U13447 (N_13447,N_12046,N_12156);
nand U13448 (N_13448,N_12526,N_12287);
or U13449 (N_13449,N_12193,N_12562);
and U13450 (N_13450,N_12452,N_12671);
and U13451 (N_13451,N_12114,N_12599);
or U13452 (N_13452,N_12717,N_12693);
or U13453 (N_13453,N_12743,N_12233);
nand U13454 (N_13454,N_12543,N_12304);
nand U13455 (N_13455,N_12518,N_12182);
or U13456 (N_13456,N_12175,N_12277);
or U13457 (N_13457,N_12257,N_12064);
nand U13458 (N_13458,N_12589,N_12251);
or U13459 (N_13459,N_12728,N_12662);
or U13460 (N_13460,N_12045,N_12046);
nor U13461 (N_13461,N_12082,N_12482);
and U13462 (N_13462,N_12530,N_12739);
and U13463 (N_13463,N_12715,N_12397);
and U13464 (N_13464,N_12631,N_12207);
nor U13465 (N_13465,N_12009,N_12396);
xor U13466 (N_13466,N_12158,N_12616);
xnor U13467 (N_13467,N_12406,N_12475);
nor U13468 (N_13468,N_12550,N_12593);
nor U13469 (N_13469,N_12268,N_12565);
or U13470 (N_13470,N_12071,N_12681);
xnor U13471 (N_13471,N_12243,N_12319);
or U13472 (N_13472,N_12648,N_12527);
nand U13473 (N_13473,N_12690,N_12743);
xor U13474 (N_13474,N_12054,N_12280);
nand U13475 (N_13475,N_12648,N_12229);
xnor U13476 (N_13476,N_12141,N_12206);
nand U13477 (N_13477,N_12231,N_12364);
nor U13478 (N_13478,N_12587,N_12715);
and U13479 (N_13479,N_12054,N_12019);
xor U13480 (N_13480,N_12045,N_12364);
nand U13481 (N_13481,N_12377,N_12042);
nand U13482 (N_13482,N_12484,N_12172);
or U13483 (N_13483,N_12319,N_12551);
nand U13484 (N_13484,N_12381,N_12205);
or U13485 (N_13485,N_12352,N_12697);
or U13486 (N_13486,N_12548,N_12668);
nor U13487 (N_13487,N_12003,N_12076);
nand U13488 (N_13488,N_12282,N_12612);
or U13489 (N_13489,N_12577,N_12119);
and U13490 (N_13490,N_12413,N_12655);
xor U13491 (N_13491,N_12631,N_12744);
xnor U13492 (N_13492,N_12253,N_12169);
nand U13493 (N_13493,N_12427,N_12088);
or U13494 (N_13494,N_12316,N_12360);
nor U13495 (N_13495,N_12197,N_12343);
nor U13496 (N_13496,N_12742,N_12302);
xor U13497 (N_13497,N_12632,N_12450);
xor U13498 (N_13498,N_12739,N_12681);
nor U13499 (N_13499,N_12685,N_12322);
or U13500 (N_13500,N_13215,N_12830);
xor U13501 (N_13501,N_13091,N_13234);
and U13502 (N_13502,N_13422,N_13315);
xnor U13503 (N_13503,N_13388,N_12809);
xor U13504 (N_13504,N_13105,N_12971);
nand U13505 (N_13505,N_13126,N_13001);
and U13506 (N_13506,N_13272,N_12801);
or U13507 (N_13507,N_13265,N_13482);
xnor U13508 (N_13508,N_13078,N_13411);
and U13509 (N_13509,N_13246,N_13281);
nor U13510 (N_13510,N_13393,N_12914);
nand U13511 (N_13511,N_13174,N_12843);
nor U13512 (N_13512,N_13287,N_13130);
or U13513 (N_13513,N_13071,N_13317);
xnor U13514 (N_13514,N_13445,N_13466);
and U13515 (N_13515,N_13335,N_12845);
nand U13516 (N_13516,N_13183,N_13116);
nor U13517 (N_13517,N_13404,N_12981);
nand U13518 (N_13518,N_12915,N_12821);
or U13519 (N_13519,N_13124,N_13112);
nor U13520 (N_13520,N_12857,N_13024);
xor U13521 (N_13521,N_13353,N_13311);
nor U13522 (N_13522,N_13408,N_12885);
nand U13523 (N_13523,N_13370,N_13048);
nand U13524 (N_13524,N_13182,N_13232);
nand U13525 (N_13525,N_13381,N_13449);
nand U13526 (N_13526,N_13344,N_12965);
and U13527 (N_13527,N_12866,N_12973);
xor U13528 (N_13528,N_13484,N_12775);
nand U13529 (N_13529,N_13131,N_13096);
nor U13530 (N_13530,N_13384,N_13206);
nand U13531 (N_13531,N_13486,N_13268);
and U13532 (N_13532,N_13127,N_13329);
nor U13533 (N_13533,N_12819,N_12774);
or U13534 (N_13534,N_13283,N_13022);
or U13535 (N_13535,N_12756,N_12794);
and U13536 (N_13536,N_13398,N_13495);
or U13537 (N_13537,N_13336,N_12964);
nor U13538 (N_13538,N_13417,N_13029);
or U13539 (N_13539,N_13374,N_13386);
nand U13540 (N_13540,N_12955,N_12936);
or U13541 (N_13541,N_12769,N_13045);
nand U13542 (N_13542,N_13196,N_12968);
xor U13543 (N_13543,N_13397,N_12935);
nand U13544 (N_13544,N_13223,N_13240);
xor U13545 (N_13545,N_12822,N_13144);
nand U13546 (N_13546,N_12842,N_13017);
or U13547 (N_13547,N_12934,N_13054);
nand U13548 (N_13548,N_13178,N_12933);
nand U13549 (N_13549,N_12762,N_12764);
and U13550 (N_13550,N_12940,N_13209);
nor U13551 (N_13551,N_12938,N_13172);
xnor U13552 (N_13552,N_13296,N_13431);
and U13553 (N_13553,N_13103,N_12929);
nor U13554 (N_13554,N_13237,N_12810);
nor U13555 (N_13555,N_13361,N_13138);
xor U13556 (N_13556,N_12758,N_12861);
xnor U13557 (N_13557,N_13396,N_12926);
nor U13558 (N_13558,N_13421,N_13038);
and U13559 (N_13559,N_12972,N_12923);
nor U13560 (N_13560,N_13000,N_12848);
xnor U13561 (N_13561,N_12831,N_12907);
xnor U13562 (N_13562,N_13239,N_13288);
nor U13563 (N_13563,N_12835,N_12948);
or U13564 (N_13564,N_13297,N_13260);
nor U13565 (N_13565,N_13162,N_13390);
and U13566 (N_13566,N_12785,N_13125);
nor U13567 (N_13567,N_13471,N_13301);
nand U13568 (N_13568,N_13492,N_13286);
or U13569 (N_13569,N_13316,N_13064);
xor U13570 (N_13570,N_13053,N_13436);
and U13571 (N_13571,N_13075,N_12913);
nand U13572 (N_13572,N_13101,N_13321);
or U13573 (N_13573,N_13158,N_12751);
and U13574 (N_13574,N_13032,N_12757);
nor U13575 (N_13575,N_13171,N_13472);
nor U13576 (N_13576,N_13226,N_13100);
nand U13577 (N_13577,N_12874,N_13345);
and U13578 (N_13578,N_13199,N_13355);
nor U13579 (N_13579,N_12957,N_12943);
and U13580 (N_13580,N_12966,N_12765);
or U13581 (N_13581,N_13010,N_13469);
or U13582 (N_13582,N_12901,N_13210);
and U13583 (N_13583,N_13496,N_13279);
xor U13584 (N_13584,N_13350,N_12912);
nand U13585 (N_13585,N_13008,N_13155);
and U13586 (N_13586,N_12859,N_13018);
xor U13587 (N_13587,N_12873,N_12868);
xor U13588 (N_13588,N_13136,N_13086);
or U13589 (N_13589,N_13128,N_12827);
nor U13590 (N_13590,N_13446,N_13189);
and U13591 (N_13591,N_13443,N_12939);
nand U13592 (N_13592,N_13147,N_12814);
nand U13593 (N_13593,N_12882,N_12941);
and U13594 (N_13594,N_13019,N_13391);
nand U13595 (N_13595,N_13014,N_12851);
nor U13596 (N_13596,N_12927,N_13269);
nor U13597 (N_13597,N_13457,N_12906);
nor U13598 (N_13598,N_13088,N_13238);
and U13599 (N_13599,N_12790,N_13331);
and U13600 (N_13600,N_13094,N_13490);
and U13601 (N_13601,N_13477,N_13102);
or U13602 (N_13602,N_13049,N_13428);
nand U13603 (N_13603,N_13356,N_13383);
and U13604 (N_13604,N_13399,N_13267);
or U13605 (N_13605,N_13177,N_13221);
nor U13606 (N_13606,N_12904,N_13135);
and U13607 (N_13607,N_12897,N_13072);
and U13608 (N_13608,N_13452,N_12782);
xor U13609 (N_13609,N_12813,N_13407);
nor U13610 (N_13610,N_12766,N_13392);
nor U13611 (N_13611,N_12989,N_13263);
and U13612 (N_13612,N_12777,N_13137);
xor U13613 (N_13613,N_13365,N_12967);
xor U13614 (N_13614,N_13044,N_12750);
nor U13615 (N_13615,N_12911,N_13227);
nor U13616 (N_13616,N_13229,N_13025);
nand U13617 (N_13617,N_13491,N_13465);
nor U13618 (N_13618,N_12807,N_13497);
nor U13619 (N_13619,N_13122,N_12872);
nor U13620 (N_13620,N_13415,N_13203);
nand U13621 (N_13621,N_13430,N_12974);
nand U13622 (N_13622,N_13151,N_13163);
xnor U13623 (N_13623,N_12902,N_13458);
xor U13624 (N_13624,N_13197,N_13222);
or U13625 (N_13625,N_12992,N_13299);
or U13626 (N_13626,N_13358,N_13473);
or U13627 (N_13627,N_12818,N_13323);
and U13628 (N_13628,N_13031,N_13170);
xnor U13629 (N_13629,N_13498,N_12802);
or U13630 (N_13630,N_12773,N_13247);
nor U13631 (N_13631,N_13141,N_13173);
xor U13632 (N_13632,N_12987,N_12894);
nand U13633 (N_13633,N_13184,N_12828);
xor U13634 (N_13634,N_13156,N_13456);
nor U13635 (N_13635,N_12924,N_13195);
nand U13636 (N_13636,N_13461,N_12791);
and U13637 (N_13637,N_12884,N_13132);
nand U13638 (N_13638,N_13190,N_12786);
or U13639 (N_13639,N_13187,N_12772);
xor U13640 (N_13640,N_13035,N_12918);
and U13641 (N_13641,N_13282,N_12792);
or U13642 (N_13642,N_13327,N_13121);
or U13643 (N_13643,N_12886,N_12909);
and U13644 (N_13644,N_13055,N_13328);
and U13645 (N_13645,N_12800,N_13143);
or U13646 (N_13646,N_12853,N_13441);
and U13647 (N_13647,N_13074,N_13146);
and U13648 (N_13648,N_13012,N_12900);
nand U13649 (N_13649,N_13273,N_12789);
nand U13650 (N_13650,N_13319,N_12899);
nor U13651 (N_13651,N_12847,N_13027);
and U13652 (N_13652,N_12783,N_12919);
nand U13653 (N_13653,N_13460,N_12895);
and U13654 (N_13654,N_13409,N_12931);
nand U13655 (N_13655,N_13423,N_13275);
or U13656 (N_13656,N_12759,N_12871);
and U13657 (N_13657,N_13157,N_12763);
xnor U13658 (N_13658,N_13082,N_12865);
nor U13659 (N_13659,N_13050,N_13485);
xor U13660 (N_13660,N_13451,N_13264);
and U13661 (N_13661,N_13167,N_12799);
xor U13662 (N_13662,N_13266,N_13214);
nand U13663 (N_13663,N_13334,N_13410);
nor U13664 (N_13664,N_12905,N_13208);
nand U13665 (N_13665,N_13437,N_12985);
nand U13666 (N_13666,N_13108,N_13230);
nand U13667 (N_13667,N_13258,N_13385);
or U13668 (N_13668,N_12982,N_13198);
xor U13669 (N_13669,N_13016,N_12978);
nor U13670 (N_13670,N_12977,N_13483);
xnor U13671 (N_13671,N_13120,N_13169);
nand U13672 (N_13672,N_13425,N_12846);
and U13673 (N_13673,N_13111,N_13090);
and U13674 (N_13674,N_13148,N_13340);
and U13675 (N_13675,N_13363,N_12999);
nor U13676 (N_13676,N_12979,N_12951);
or U13677 (N_13677,N_12963,N_13481);
or U13678 (N_13678,N_13056,N_13164);
and U13679 (N_13679,N_12770,N_13194);
and U13680 (N_13680,N_12817,N_13207);
xnor U13681 (N_13681,N_13205,N_13073);
or U13682 (N_13682,N_13362,N_13114);
and U13683 (N_13683,N_13305,N_13257);
and U13684 (N_13684,N_12850,N_13252);
or U13685 (N_13685,N_13300,N_12855);
and U13686 (N_13686,N_13290,N_12930);
nand U13687 (N_13687,N_13464,N_13333);
nor U13688 (N_13688,N_12976,N_12984);
xnor U13689 (N_13689,N_12961,N_12944);
or U13690 (N_13690,N_12958,N_13220);
xnor U13691 (N_13691,N_13002,N_13068);
and U13692 (N_13692,N_13318,N_13015);
and U13693 (N_13693,N_13005,N_12754);
and U13694 (N_13694,N_12925,N_13432);
nand U13695 (N_13695,N_13079,N_13285);
xor U13696 (N_13696,N_13134,N_12804);
nor U13697 (N_13697,N_13254,N_13439);
nor U13698 (N_13698,N_13293,N_12761);
nor U13699 (N_13699,N_13342,N_12864);
xor U13700 (N_13700,N_12797,N_13069);
and U13701 (N_13701,N_12863,N_12798);
xor U13702 (N_13702,N_13322,N_12768);
nor U13703 (N_13703,N_13249,N_12760);
and U13704 (N_13704,N_13080,N_12877);
or U13705 (N_13705,N_12771,N_13480);
nor U13706 (N_13706,N_13081,N_13021);
xor U13707 (N_13707,N_13168,N_12780);
and U13708 (N_13708,N_13175,N_12983);
or U13709 (N_13709,N_13089,N_13129);
or U13710 (N_13710,N_13060,N_13034);
nand U13711 (N_13711,N_12858,N_13166);
nand U13712 (N_13712,N_12815,N_12903);
nand U13713 (N_13713,N_12844,N_13104);
and U13714 (N_13714,N_13119,N_12869);
and U13715 (N_13715,N_13487,N_12816);
nor U13716 (N_13716,N_13200,N_13295);
or U13717 (N_13717,N_13244,N_12956);
nor U13718 (N_13718,N_12932,N_13212);
xor U13719 (N_13719,N_13447,N_13113);
or U13720 (N_13720,N_13403,N_13095);
nor U13721 (N_13721,N_13020,N_13133);
xnor U13722 (N_13722,N_13427,N_12753);
and U13723 (N_13723,N_13494,N_12784);
xnor U13724 (N_13724,N_12991,N_13092);
and U13725 (N_13725,N_13354,N_12755);
xor U13726 (N_13726,N_13192,N_13217);
nor U13727 (N_13727,N_12824,N_13476);
or U13728 (N_13728,N_13242,N_13067);
nand U13729 (N_13729,N_13367,N_12937);
xnor U13730 (N_13730,N_12805,N_12996);
nor U13731 (N_13731,N_12995,N_13280);
or U13732 (N_13732,N_12921,N_13314);
and U13733 (N_13733,N_13028,N_12867);
and U13734 (N_13734,N_12825,N_13372);
nor U13735 (N_13735,N_13419,N_12832);
nor U13736 (N_13736,N_13371,N_13085);
nand U13737 (N_13737,N_13413,N_13062);
and U13738 (N_13738,N_12834,N_12849);
xnor U13739 (N_13739,N_13202,N_13026);
xor U13740 (N_13740,N_12969,N_13036);
and U13741 (N_13741,N_13007,N_13400);
xor U13742 (N_13742,N_13270,N_13470);
nor U13743 (N_13743,N_13087,N_12896);
nor U13744 (N_13744,N_13150,N_12793);
xnor U13745 (N_13745,N_13211,N_12854);
xnor U13746 (N_13746,N_13046,N_13377);
xnor U13747 (N_13747,N_13373,N_13149);
xnor U13748 (N_13748,N_13325,N_13330);
or U13749 (N_13749,N_13455,N_13303);
and U13750 (N_13750,N_13023,N_13351);
xnor U13751 (N_13751,N_13180,N_12876);
xnor U13752 (N_13752,N_12988,N_13343);
xor U13753 (N_13753,N_12820,N_13011);
and U13754 (N_13754,N_13219,N_12954);
and U13755 (N_13755,N_12887,N_12891);
and U13756 (N_13756,N_12838,N_12778);
and U13757 (N_13757,N_13145,N_13193);
nor U13758 (N_13758,N_12946,N_13165);
xnor U13759 (N_13759,N_13274,N_13043);
or U13760 (N_13760,N_13488,N_13499);
nor U13761 (N_13761,N_13426,N_12910);
xor U13762 (N_13762,N_13448,N_12898);
xnor U13763 (N_13763,N_12837,N_13294);
nand U13764 (N_13764,N_13152,N_12826);
and U13765 (N_13765,N_13284,N_13115);
nand U13766 (N_13766,N_13106,N_13454);
or U13767 (N_13767,N_12962,N_13123);
and U13768 (N_13768,N_13235,N_12928);
or U13769 (N_13769,N_13204,N_13429);
and U13770 (N_13770,N_13444,N_13277);
xor U13771 (N_13771,N_13218,N_12888);
nor U13772 (N_13772,N_13216,N_12949);
nand U13773 (N_13773,N_13213,N_13379);
and U13774 (N_13774,N_12829,N_13369);
xor U13775 (N_13775,N_13030,N_13324);
nor U13776 (N_13776,N_13360,N_13271);
nor U13777 (N_13777,N_13142,N_12960);
nor U13778 (N_13778,N_13313,N_13406);
or U13779 (N_13779,N_13040,N_13185);
nor U13780 (N_13780,N_12870,N_12908);
nand U13781 (N_13781,N_13364,N_13259);
xor U13782 (N_13782,N_13006,N_13063);
nand U13783 (N_13783,N_13181,N_13424);
nand U13784 (N_13784,N_12840,N_13245);
nand U13785 (N_13785,N_13438,N_13387);
or U13786 (N_13786,N_12920,N_12752);
nand U13787 (N_13787,N_13154,N_13039);
xnor U13788 (N_13788,N_13076,N_13312);
xor U13789 (N_13789,N_12852,N_12875);
nor U13790 (N_13790,N_13179,N_12942);
xor U13791 (N_13791,N_13395,N_13308);
xnor U13792 (N_13792,N_12796,N_13110);
or U13793 (N_13793,N_13394,N_12917);
nor U13794 (N_13794,N_13224,N_13109);
and U13795 (N_13795,N_12880,N_13107);
xor U13796 (N_13796,N_13255,N_13052);
and U13797 (N_13797,N_13401,N_12808);
nand U13798 (N_13798,N_13368,N_12823);
or U13799 (N_13799,N_13070,N_13414);
and U13800 (N_13800,N_12998,N_13186);
nand U13801 (N_13801,N_13346,N_13479);
nor U13802 (N_13802,N_13352,N_12856);
or U13803 (N_13803,N_13066,N_13376);
nor U13804 (N_13804,N_13153,N_13037);
and U13805 (N_13805,N_13118,N_13278);
xor U13806 (N_13806,N_12889,N_13097);
nand U13807 (N_13807,N_13262,N_13047);
xor U13808 (N_13808,N_13468,N_13348);
xor U13809 (N_13809,N_12776,N_12781);
nand U13810 (N_13810,N_13357,N_13004);
nor U13811 (N_13811,N_12881,N_12767);
nor U13812 (N_13812,N_13058,N_13033);
or U13813 (N_13813,N_13292,N_13251);
and U13814 (N_13814,N_12916,N_13420);
xor U13815 (N_13815,N_12980,N_13416);
xnor U13816 (N_13816,N_12860,N_12833);
nor U13817 (N_13817,N_13339,N_13093);
and U13818 (N_13818,N_13326,N_13375);
nand U13819 (N_13819,N_13261,N_12997);
nor U13820 (N_13820,N_13378,N_13276);
and U13821 (N_13821,N_13140,N_13159);
and U13822 (N_13822,N_12879,N_13013);
or U13823 (N_13823,N_12841,N_12788);
and U13824 (N_13824,N_12883,N_12839);
and U13825 (N_13825,N_13440,N_13291);
nor U13826 (N_13826,N_13302,N_13042);
or U13827 (N_13827,N_13338,N_13061);
nor U13828 (N_13828,N_13084,N_12803);
or U13829 (N_13829,N_12953,N_13405);
and U13830 (N_13830,N_12990,N_13057);
nand U13831 (N_13831,N_13304,N_13083);
nor U13832 (N_13832,N_13231,N_13065);
nand U13833 (N_13833,N_13475,N_13160);
nor U13834 (N_13834,N_13478,N_12811);
or U13835 (N_13835,N_12945,N_13117);
nor U13836 (N_13836,N_13453,N_13349);
xor U13837 (N_13837,N_13289,N_13256);
or U13838 (N_13838,N_13382,N_13320);
xnor U13839 (N_13839,N_12959,N_13332);
xnor U13840 (N_13840,N_13248,N_13041);
and U13841 (N_13841,N_13051,N_13139);
xor U13842 (N_13842,N_12806,N_13059);
or U13843 (N_13843,N_13462,N_13307);
or U13844 (N_13844,N_12970,N_12922);
xor U13845 (N_13845,N_13191,N_13493);
and U13846 (N_13846,N_13253,N_13337);
nor U13847 (N_13847,N_13309,N_13298);
and U13848 (N_13848,N_13176,N_12975);
nor U13849 (N_13849,N_12993,N_13380);
nor U13850 (N_13850,N_13236,N_13241);
xnor U13851 (N_13851,N_13161,N_13201);
nor U13852 (N_13852,N_13098,N_13450);
and U13853 (N_13853,N_13435,N_13389);
xnor U13854 (N_13854,N_13233,N_13459);
nand U13855 (N_13855,N_13099,N_12862);
and U13856 (N_13856,N_13228,N_13077);
or U13857 (N_13857,N_13418,N_13366);
xor U13858 (N_13858,N_12812,N_13402);
and U13859 (N_13859,N_12795,N_12878);
nor U13860 (N_13860,N_13442,N_13306);
nand U13861 (N_13861,N_12892,N_12947);
and U13862 (N_13862,N_13467,N_12952);
or U13863 (N_13863,N_13003,N_13250);
and U13864 (N_13864,N_12994,N_13412);
nor U13865 (N_13865,N_12836,N_12950);
nand U13866 (N_13866,N_12986,N_13463);
or U13867 (N_13867,N_13188,N_13347);
or U13868 (N_13868,N_13243,N_13009);
or U13869 (N_13869,N_12787,N_12890);
or U13870 (N_13870,N_12779,N_13310);
or U13871 (N_13871,N_13474,N_13359);
and U13872 (N_13872,N_12893,N_13225);
nand U13873 (N_13873,N_13489,N_13433);
xor U13874 (N_13874,N_13341,N_13434);
xnor U13875 (N_13875,N_13417,N_13297);
or U13876 (N_13876,N_13230,N_12914);
or U13877 (N_13877,N_13112,N_13443);
nor U13878 (N_13878,N_13175,N_13121);
nand U13879 (N_13879,N_13277,N_12761);
or U13880 (N_13880,N_13260,N_12976);
and U13881 (N_13881,N_12797,N_12851);
xor U13882 (N_13882,N_13088,N_13293);
or U13883 (N_13883,N_13461,N_13012);
nor U13884 (N_13884,N_13218,N_13437);
nand U13885 (N_13885,N_13014,N_12857);
xor U13886 (N_13886,N_13393,N_13455);
xnor U13887 (N_13887,N_12966,N_13341);
and U13888 (N_13888,N_12973,N_13480);
nor U13889 (N_13889,N_12922,N_12912);
nor U13890 (N_13890,N_13475,N_13198);
nand U13891 (N_13891,N_12847,N_13366);
xor U13892 (N_13892,N_12927,N_13026);
nor U13893 (N_13893,N_13043,N_12792);
and U13894 (N_13894,N_12806,N_12943);
nand U13895 (N_13895,N_13354,N_13166);
xnor U13896 (N_13896,N_12907,N_12768);
and U13897 (N_13897,N_13465,N_13148);
or U13898 (N_13898,N_13040,N_13427);
nor U13899 (N_13899,N_12773,N_13345);
or U13900 (N_13900,N_13114,N_13299);
nor U13901 (N_13901,N_13189,N_12774);
nand U13902 (N_13902,N_13231,N_13178);
nor U13903 (N_13903,N_13409,N_13203);
or U13904 (N_13904,N_13321,N_12818);
nand U13905 (N_13905,N_13011,N_13329);
and U13906 (N_13906,N_12829,N_13123);
or U13907 (N_13907,N_13423,N_13442);
nand U13908 (N_13908,N_13269,N_13122);
xnor U13909 (N_13909,N_13159,N_13448);
or U13910 (N_13910,N_13410,N_13216);
xor U13911 (N_13911,N_13283,N_12805);
and U13912 (N_13912,N_13170,N_13096);
or U13913 (N_13913,N_13060,N_12779);
nor U13914 (N_13914,N_13068,N_13113);
and U13915 (N_13915,N_13446,N_13237);
or U13916 (N_13916,N_13382,N_13298);
xnor U13917 (N_13917,N_13127,N_13279);
and U13918 (N_13918,N_13396,N_13331);
or U13919 (N_13919,N_13218,N_13446);
nand U13920 (N_13920,N_13104,N_12863);
or U13921 (N_13921,N_13489,N_13366);
xor U13922 (N_13922,N_12775,N_12840);
xnor U13923 (N_13923,N_13027,N_12880);
or U13924 (N_13924,N_13234,N_13228);
and U13925 (N_13925,N_13440,N_13192);
or U13926 (N_13926,N_12974,N_12915);
nand U13927 (N_13927,N_13422,N_13436);
xnor U13928 (N_13928,N_12830,N_13013);
nor U13929 (N_13929,N_12765,N_12755);
xnor U13930 (N_13930,N_13256,N_13170);
nand U13931 (N_13931,N_13460,N_12970);
xnor U13932 (N_13932,N_12780,N_12854);
and U13933 (N_13933,N_13348,N_13128);
nor U13934 (N_13934,N_13399,N_13369);
xnor U13935 (N_13935,N_12983,N_13470);
or U13936 (N_13936,N_13214,N_13199);
nor U13937 (N_13937,N_13242,N_13344);
or U13938 (N_13938,N_13174,N_12840);
nand U13939 (N_13939,N_13404,N_13048);
and U13940 (N_13940,N_12850,N_13352);
nor U13941 (N_13941,N_12781,N_12806);
xnor U13942 (N_13942,N_12856,N_13459);
and U13943 (N_13943,N_13125,N_12780);
nor U13944 (N_13944,N_12813,N_13261);
and U13945 (N_13945,N_12986,N_13253);
xnor U13946 (N_13946,N_13393,N_13360);
and U13947 (N_13947,N_13387,N_12773);
or U13948 (N_13948,N_12813,N_12885);
nand U13949 (N_13949,N_12869,N_13124);
or U13950 (N_13950,N_13072,N_13460);
nor U13951 (N_13951,N_13344,N_13200);
and U13952 (N_13952,N_12837,N_13377);
nand U13953 (N_13953,N_13207,N_12902);
and U13954 (N_13954,N_13092,N_12913);
nand U13955 (N_13955,N_12977,N_13229);
nand U13956 (N_13956,N_13118,N_13090);
or U13957 (N_13957,N_13078,N_13271);
and U13958 (N_13958,N_12926,N_13227);
xor U13959 (N_13959,N_13211,N_12910);
xor U13960 (N_13960,N_12802,N_12893);
or U13961 (N_13961,N_12981,N_12950);
nor U13962 (N_13962,N_12755,N_13288);
xor U13963 (N_13963,N_13377,N_13023);
nor U13964 (N_13964,N_13499,N_12941);
or U13965 (N_13965,N_13320,N_13089);
or U13966 (N_13966,N_13241,N_13060);
nand U13967 (N_13967,N_12995,N_13134);
and U13968 (N_13968,N_13327,N_13220);
or U13969 (N_13969,N_13451,N_12904);
xor U13970 (N_13970,N_13356,N_13281);
nand U13971 (N_13971,N_12998,N_12793);
or U13972 (N_13972,N_13098,N_13483);
or U13973 (N_13973,N_13163,N_13016);
or U13974 (N_13974,N_13391,N_12925);
nand U13975 (N_13975,N_13168,N_12912);
and U13976 (N_13976,N_12937,N_13058);
or U13977 (N_13977,N_12967,N_13061);
and U13978 (N_13978,N_12905,N_13266);
nor U13979 (N_13979,N_12945,N_13101);
nor U13980 (N_13980,N_12759,N_13443);
nand U13981 (N_13981,N_13400,N_13000);
and U13982 (N_13982,N_13058,N_13061);
nor U13983 (N_13983,N_13150,N_13379);
and U13984 (N_13984,N_12981,N_12844);
xnor U13985 (N_13985,N_12947,N_13325);
and U13986 (N_13986,N_13322,N_13302);
or U13987 (N_13987,N_13293,N_12923);
xnor U13988 (N_13988,N_12953,N_13481);
nor U13989 (N_13989,N_12901,N_13251);
nor U13990 (N_13990,N_13070,N_12943);
and U13991 (N_13991,N_12769,N_13233);
nand U13992 (N_13992,N_13024,N_12927);
xnor U13993 (N_13993,N_13345,N_13107);
and U13994 (N_13994,N_13212,N_13236);
and U13995 (N_13995,N_12841,N_13389);
and U13996 (N_13996,N_13497,N_13104);
nand U13997 (N_13997,N_13080,N_13000);
nand U13998 (N_13998,N_12834,N_12940);
and U13999 (N_13999,N_13417,N_13275);
nor U14000 (N_14000,N_13021,N_13206);
xnor U14001 (N_14001,N_13202,N_13187);
nor U14002 (N_14002,N_12787,N_13308);
and U14003 (N_14003,N_13287,N_12900);
or U14004 (N_14004,N_13417,N_12997);
or U14005 (N_14005,N_13052,N_13383);
or U14006 (N_14006,N_13020,N_12848);
or U14007 (N_14007,N_12771,N_12822);
xnor U14008 (N_14008,N_13058,N_13010);
nor U14009 (N_14009,N_13348,N_12880);
nand U14010 (N_14010,N_13163,N_12863);
nand U14011 (N_14011,N_12931,N_12893);
and U14012 (N_14012,N_13253,N_13349);
nor U14013 (N_14013,N_13346,N_13021);
nor U14014 (N_14014,N_13350,N_13311);
nand U14015 (N_14015,N_13367,N_13434);
and U14016 (N_14016,N_13479,N_13445);
or U14017 (N_14017,N_12819,N_13417);
and U14018 (N_14018,N_13475,N_13323);
and U14019 (N_14019,N_13194,N_12900);
or U14020 (N_14020,N_13396,N_13470);
xor U14021 (N_14021,N_13417,N_13289);
or U14022 (N_14022,N_12895,N_13184);
and U14023 (N_14023,N_13193,N_12778);
or U14024 (N_14024,N_12793,N_13123);
or U14025 (N_14025,N_13060,N_13342);
nor U14026 (N_14026,N_13066,N_13308);
or U14027 (N_14027,N_12769,N_12782);
xnor U14028 (N_14028,N_13480,N_12915);
nand U14029 (N_14029,N_13076,N_13188);
and U14030 (N_14030,N_13461,N_12814);
and U14031 (N_14031,N_13303,N_13001);
and U14032 (N_14032,N_12965,N_13052);
nand U14033 (N_14033,N_12981,N_13375);
or U14034 (N_14034,N_13344,N_12839);
nand U14035 (N_14035,N_13346,N_12988);
xor U14036 (N_14036,N_13060,N_13143);
nand U14037 (N_14037,N_13248,N_12939);
nand U14038 (N_14038,N_12774,N_12834);
nor U14039 (N_14039,N_13423,N_13351);
xnor U14040 (N_14040,N_13126,N_13116);
nor U14041 (N_14041,N_13437,N_13085);
nand U14042 (N_14042,N_13199,N_12847);
and U14043 (N_14043,N_12782,N_13323);
xnor U14044 (N_14044,N_12844,N_13145);
nor U14045 (N_14045,N_13396,N_13199);
nand U14046 (N_14046,N_13066,N_13462);
nand U14047 (N_14047,N_12758,N_13388);
nor U14048 (N_14048,N_13181,N_13360);
nand U14049 (N_14049,N_13395,N_13277);
or U14050 (N_14050,N_13426,N_13312);
nand U14051 (N_14051,N_12778,N_13009);
or U14052 (N_14052,N_12835,N_13225);
xor U14053 (N_14053,N_13227,N_12922);
nand U14054 (N_14054,N_13475,N_13453);
xor U14055 (N_14055,N_13207,N_12920);
and U14056 (N_14056,N_12832,N_13198);
and U14057 (N_14057,N_13268,N_13212);
nand U14058 (N_14058,N_13204,N_12920);
nor U14059 (N_14059,N_12929,N_12860);
xnor U14060 (N_14060,N_13461,N_13246);
and U14061 (N_14061,N_12860,N_13315);
or U14062 (N_14062,N_13311,N_13473);
nor U14063 (N_14063,N_12915,N_13196);
nand U14064 (N_14064,N_13171,N_13012);
and U14065 (N_14065,N_13294,N_13256);
nor U14066 (N_14066,N_13005,N_12758);
xor U14067 (N_14067,N_13197,N_13001);
nand U14068 (N_14068,N_13469,N_13499);
or U14069 (N_14069,N_12815,N_12769);
and U14070 (N_14070,N_12754,N_13405);
nor U14071 (N_14071,N_13398,N_12967);
xor U14072 (N_14072,N_13174,N_12899);
nor U14073 (N_14073,N_12937,N_13057);
nor U14074 (N_14074,N_13438,N_13074);
xnor U14075 (N_14075,N_13315,N_12898);
or U14076 (N_14076,N_13018,N_13418);
xor U14077 (N_14077,N_13229,N_13104);
or U14078 (N_14078,N_13234,N_12764);
nor U14079 (N_14079,N_13042,N_12993);
xnor U14080 (N_14080,N_13443,N_13081);
xnor U14081 (N_14081,N_12841,N_13200);
nor U14082 (N_14082,N_13429,N_13478);
xnor U14083 (N_14083,N_13320,N_13240);
xor U14084 (N_14084,N_13194,N_13288);
nand U14085 (N_14085,N_12988,N_13458);
or U14086 (N_14086,N_12821,N_13324);
nor U14087 (N_14087,N_13430,N_13033);
xor U14088 (N_14088,N_12906,N_12910);
or U14089 (N_14089,N_13216,N_13348);
nor U14090 (N_14090,N_13321,N_13018);
xor U14091 (N_14091,N_13234,N_13202);
or U14092 (N_14092,N_13108,N_13245);
nor U14093 (N_14093,N_13308,N_13422);
nor U14094 (N_14094,N_13109,N_13490);
xor U14095 (N_14095,N_12853,N_13148);
or U14096 (N_14096,N_13497,N_13265);
nand U14097 (N_14097,N_13462,N_13487);
nor U14098 (N_14098,N_13245,N_12990);
nand U14099 (N_14099,N_13148,N_12931);
and U14100 (N_14100,N_13434,N_12980);
xnor U14101 (N_14101,N_12840,N_13327);
xor U14102 (N_14102,N_12960,N_12836);
or U14103 (N_14103,N_13435,N_13097);
nor U14104 (N_14104,N_12984,N_12923);
and U14105 (N_14105,N_13423,N_13220);
or U14106 (N_14106,N_12816,N_12760);
or U14107 (N_14107,N_13439,N_12897);
xnor U14108 (N_14108,N_13236,N_13187);
nor U14109 (N_14109,N_12912,N_12802);
nor U14110 (N_14110,N_12882,N_13117);
nor U14111 (N_14111,N_13049,N_13303);
xor U14112 (N_14112,N_13388,N_13298);
xnor U14113 (N_14113,N_12860,N_13285);
nor U14114 (N_14114,N_13189,N_13238);
nor U14115 (N_14115,N_13251,N_13459);
xor U14116 (N_14116,N_13015,N_12903);
or U14117 (N_14117,N_13047,N_12804);
and U14118 (N_14118,N_12888,N_13096);
nor U14119 (N_14119,N_13155,N_12794);
nand U14120 (N_14120,N_12917,N_13284);
or U14121 (N_14121,N_13118,N_13223);
nand U14122 (N_14122,N_13322,N_13190);
nor U14123 (N_14123,N_13049,N_13218);
xor U14124 (N_14124,N_12813,N_12904);
xor U14125 (N_14125,N_13101,N_12798);
and U14126 (N_14126,N_13045,N_13273);
and U14127 (N_14127,N_13409,N_13050);
or U14128 (N_14128,N_13373,N_12853);
xnor U14129 (N_14129,N_13054,N_13091);
xnor U14130 (N_14130,N_13434,N_13497);
nand U14131 (N_14131,N_13025,N_12902);
xor U14132 (N_14132,N_13223,N_13413);
nand U14133 (N_14133,N_12948,N_13066);
xor U14134 (N_14134,N_12793,N_13429);
xor U14135 (N_14135,N_13178,N_13474);
nand U14136 (N_14136,N_13233,N_13044);
xnor U14137 (N_14137,N_13439,N_13045);
nor U14138 (N_14138,N_12912,N_13497);
or U14139 (N_14139,N_13138,N_12928);
nand U14140 (N_14140,N_13069,N_13320);
and U14141 (N_14141,N_12810,N_12894);
or U14142 (N_14142,N_13257,N_12768);
or U14143 (N_14143,N_13329,N_12973);
nand U14144 (N_14144,N_12951,N_13227);
nor U14145 (N_14145,N_13267,N_13150);
xor U14146 (N_14146,N_12868,N_12783);
and U14147 (N_14147,N_12830,N_13409);
nor U14148 (N_14148,N_12950,N_13201);
and U14149 (N_14149,N_12798,N_13056);
nand U14150 (N_14150,N_12809,N_13149);
xnor U14151 (N_14151,N_13087,N_12857);
xnor U14152 (N_14152,N_13138,N_13146);
or U14153 (N_14153,N_13469,N_12923);
nand U14154 (N_14154,N_12976,N_13361);
and U14155 (N_14155,N_12780,N_13204);
nor U14156 (N_14156,N_13138,N_12830);
or U14157 (N_14157,N_13081,N_13156);
nor U14158 (N_14158,N_12999,N_13436);
nor U14159 (N_14159,N_13277,N_13480);
and U14160 (N_14160,N_12915,N_13289);
xor U14161 (N_14161,N_13263,N_12970);
nor U14162 (N_14162,N_13068,N_12767);
xor U14163 (N_14163,N_13175,N_13022);
and U14164 (N_14164,N_13488,N_12938);
and U14165 (N_14165,N_12849,N_12870);
xor U14166 (N_14166,N_13090,N_12770);
nor U14167 (N_14167,N_12835,N_12967);
and U14168 (N_14168,N_12823,N_13310);
and U14169 (N_14169,N_12968,N_12860);
nand U14170 (N_14170,N_12868,N_13233);
nand U14171 (N_14171,N_12846,N_13052);
or U14172 (N_14172,N_13191,N_13164);
nor U14173 (N_14173,N_13147,N_13135);
xor U14174 (N_14174,N_13433,N_12806);
nand U14175 (N_14175,N_12862,N_13360);
xor U14176 (N_14176,N_13487,N_13186);
xor U14177 (N_14177,N_13249,N_13156);
or U14178 (N_14178,N_12795,N_13371);
nand U14179 (N_14179,N_13394,N_13199);
or U14180 (N_14180,N_13111,N_13412);
xnor U14181 (N_14181,N_12837,N_13277);
nor U14182 (N_14182,N_13106,N_12765);
nand U14183 (N_14183,N_12894,N_13457);
nor U14184 (N_14184,N_13000,N_12796);
xor U14185 (N_14185,N_13044,N_12779);
or U14186 (N_14186,N_13161,N_13036);
xor U14187 (N_14187,N_13242,N_13477);
nor U14188 (N_14188,N_13339,N_13075);
and U14189 (N_14189,N_13471,N_13268);
nand U14190 (N_14190,N_13287,N_13292);
nor U14191 (N_14191,N_12908,N_12889);
or U14192 (N_14192,N_12862,N_13045);
nor U14193 (N_14193,N_13118,N_12975);
or U14194 (N_14194,N_13416,N_12858);
xor U14195 (N_14195,N_13452,N_12969);
nand U14196 (N_14196,N_13067,N_13251);
xor U14197 (N_14197,N_13365,N_13288);
nand U14198 (N_14198,N_13405,N_12959);
or U14199 (N_14199,N_13472,N_13183);
or U14200 (N_14200,N_13258,N_12788);
or U14201 (N_14201,N_12762,N_13001);
or U14202 (N_14202,N_13337,N_12790);
and U14203 (N_14203,N_12822,N_13491);
xor U14204 (N_14204,N_12936,N_13176);
nand U14205 (N_14205,N_13166,N_13434);
nand U14206 (N_14206,N_12826,N_13404);
nor U14207 (N_14207,N_12998,N_13043);
nand U14208 (N_14208,N_13194,N_13200);
or U14209 (N_14209,N_12929,N_13416);
nand U14210 (N_14210,N_13293,N_13075);
or U14211 (N_14211,N_13193,N_13180);
or U14212 (N_14212,N_12997,N_13447);
or U14213 (N_14213,N_13123,N_12936);
nor U14214 (N_14214,N_13075,N_13310);
and U14215 (N_14215,N_13145,N_12817);
xnor U14216 (N_14216,N_12888,N_13019);
xor U14217 (N_14217,N_13321,N_13380);
or U14218 (N_14218,N_12836,N_13094);
and U14219 (N_14219,N_12852,N_12938);
nand U14220 (N_14220,N_12845,N_12877);
nand U14221 (N_14221,N_13168,N_13140);
xor U14222 (N_14222,N_12868,N_13272);
nand U14223 (N_14223,N_12924,N_13411);
and U14224 (N_14224,N_13039,N_13067);
and U14225 (N_14225,N_13129,N_13292);
nor U14226 (N_14226,N_12948,N_12804);
or U14227 (N_14227,N_13409,N_12959);
xnor U14228 (N_14228,N_13249,N_13198);
or U14229 (N_14229,N_13335,N_12898);
nand U14230 (N_14230,N_12862,N_13189);
xnor U14231 (N_14231,N_12940,N_13181);
and U14232 (N_14232,N_12980,N_13030);
and U14233 (N_14233,N_13407,N_12954);
or U14234 (N_14234,N_13279,N_13389);
nor U14235 (N_14235,N_13211,N_13360);
nor U14236 (N_14236,N_12905,N_13087);
nand U14237 (N_14237,N_13010,N_12988);
or U14238 (N_14238,N_13135,N_12888);
and U14239 (N_14239,N_12892,N_13260);
nand U14240 (N_14240,N_12947,N_13204);
nor U14241 (N_14241,N_13399,N_13223);
and U14242 (N_14242,N_12902,N_12863);
nand U14243 (N_14243,N_12876,N_13134);
and U14244 (N_14244,N_12789,N_13322);
xor U14245 (N_14245,N_13127,N_13198);
and U14246 (N_14246,N_13347,N_13105);
or U14247 (N_14247,N_13304,N_13156);
nand U14248 (N_14248,N_12822,N_13269);
nor U14249 (N_14249,N_13002,N_12778);
nor U14250 (N_14250,N_13973,N_13505);
or U14251 (N_14251,N_14008,N_13569);
or U14252 (N_14252,N_13638,N_14055);
xor U14253 (N_14253,N_14091,N_13625);
nand U14254 (N_14254,N_13548,N_14038);
or U14255 (N_14255,N_13743,N_14078);
nand U14256 (N_14256,N_13783,N_14037);
nor U14257 (N_14257,N_13864,N_14079);
nand U14258 (N_14258,N_13758,N_13751);
nand U14259 (N_14259,N_13556,N_14180);
nor U14260 (N_14260,N_13666,N_13772);
nand U14261 (N_14261,N_13870,N_13636);
or U14262 (N_14262,N_13926,N_14108);
or U14263 (N_14263,N_14002,N_13782);
nor U14264 (N_14264,N_13920,N_13925);
or U14265 (N_14265,N_13602,N_13650);
nor U14266 (N_14266,N_13992,N_13922);
nor U14267 (N_14267,N_14142,N_13886);
xor U14268 (N_14268,N_13794,N_14094);
nand U14269 (N_14269,N_14068,N_14092);
or U14270 (N_14270,N_14128,N_14131);
or U14271 (N_14271,N_13940,N_14058);
nor U14272 (N_14272,N_13931,N_13934);
and U14273 (N_14273,N_14202,N_13785);
and U14274 (N_14274,N_13739,N_14192);
xor U14275 (N_14275,N_13998,N_14148);
nand U14276 (N_14276,N_13656,N_14171);
nor U14277 (N_14277,N_13781,N_14172);
or U14278 (N_14278,N_13996,N_14122);
nand U14279 (N_14279,N_13628,N_13851);
and U14280 (N_14280,N_14044,N_13849);
nor U14281 (N_14281,N_13584,N_13679);
nand U14282 (N_14282,N_13837,N_13933);
or U14283 (N_14283,N_14035,N_13899);
nand U14284 (N_14284,N_13640,N_13788);
or U14285 (N_14285,N_13552,N_13896);
xnor U14286 (N_14286,N_14211,N_13740);
nand U14287 (N_14287,N_14084,N_13589);
nor U14288 (N_14288,N_13601,N_13507);
or U14289 (N_14289,N_13819,N_13723);
nand U14290 (N_14290,N_13868,N_13972);
xnor U14291 (N_14291,N_13810,N_13800);
or U14292 (N_14292,N_13642,N_14027);
or U14293 (N_14293,N_13906,N_14057);
nor U14294 (N_14294,N_14011,N_13593);
nor U14295 (N_14295,N_14083,N_14232);
nor U14296 (N_14296,N_13790,N_14162);
or U14297 (N_14297,N_13571,N_13750);
nand U14298 (N_14298,N_13921,N_14031);
nand U14299 (N_14299,N_13527,N_14026);
and U14300 (N_14300,N_14135,N_13778);
and U14301 (N_14301,N_13732,N_13809);
or U14302 (N_14302,N_14137,N_13792);
xnor U14303 (N_14303,N_14032,N_13865);
nand U14304 (N_14304,N_14155,N_13560);
or U14305 (N_14305,N_13603,N_14080);
nor U14306 (N_14306,N_13777,N_13923);
nor U14307 (N_14307,N_14163,N_14005);
nand U14308 (N_14308,N_13504,N_13949);
nor U14309 (N_14309,N_13727,N_13699);
or U14310 (N_14310,N_13503,N_13753);
or U14311 (N_14311,N_13850,N_14085);
nor U14312 (N_14312,N_13823,N_13657);
nor U14313 (N_14313,N_13796,N_13890);
nand U14314 (N_14314,N_13918,N_13673);
and U14315 (N_14315,N_13913,N_14081);
xnor U14316 (N_14316,N_14147,N_14129);
nor U14317 (N_14317,N_13565,N_14040);
nand U14318 (N_14318,N_13957,N_13624);
xor U14319 (N_14319,N_14156,N_13787);
nand U14320 (N_14320,N_14048,N_14121);
or U14321 (N_14321,N_14033,N_13547);
or U14322 (N_14322,N_14209,N_13703);
xor U14323 (N_14323,N_13974,N_14064);
and U14324 (N_14324,N_13615,N_13539);
or U14325 (N_14325,N_13822,N_13600);
or U14326 (N_14326,N_13532,N_13844);
nor U14327 (N_14327,N_13861,N_13659);
xor U14328 (N_14328,N_13981,N_14187);
nand U14329 (N_14329,N_14089,N_13932);
nor U14330 (N_14330,N_14186,N_13508);
nand U14331 (N_14331,N_14073,N_13690);
and U14332 (N_14332,N_13830,N_14016);
xor U14333 (N_14333,N_14054,N_13721);
and U14334 (N_14334,N_14175,N_14126);
or U14335 (N_14335,N_14113,N_13522);
nor U14336 (N_14336,N_13775,N_14245);
nor U14337 (N_14337,N_13917,N_13688);
nor U14338 (N_14338,N_13726,N_13509);
xnor U14339 (N_14339,N_13544,N_13856);
and U14340 (N_14340,N_14201,N_13797);
and U14341 (N_14341,N_14169,N_13764);
or U14342 (N_14342,N_13667,N_13660);
or U14343 (N_14343,N_13985,N_14165);
xor U14344 (N_14344,N_13555,N_13528);
and U14345 (N_14345,N_13658,N_13848);
nand U14346 (N_14346,N_13910,N_14190);
and U14347 (N_14347,N_13546,N_14007);
xor U14348 (N_14348,N_14015,N_13828);
xnor U14349 (N_14349,N_14117,N_13859);
nor U14350 (N_14350,N_13754,N_13938);
nand U14351 (N_14351,N_13984,N_13803);
or U14352 (N_14352,N_13802,N_13644);
xnor U14353 (N_14353,N_13761,N_13514);
nor U14354 (N_14354,N_13558,N_13680);
or U14355 (N_14355,N_14109,N_14204);
nor U14356 (N_14356,N_14116,N_13704);
nor U14357 (N_14357,N_14235,N_13986);
and U14358 (N_14358,N_13928,N_13551);
and U14359 (N_14359,N_13676,N_13523);
or U14360 (N_14360,N_13833,N_14191);
and U14361 (N_14361,N_14111,N_14185);
nor U14362 (N_14362,N_13784,N_14206);
and U14363 (N_14363,N_13760,N_13663);
and U14364 (N_14364,N_13637,N_14067);
nor U14365 (N_14365,N_14199,N_14217);
nor U14366 (N_14366,N_14020,N_13767);
nand U14367 (N_14367,N_13643,N_14006);
or U14368 (N_14368,N_13604,N_13633);
nand U14369 (N_14369,N_13613,N_13521);
nor U14370 (N_14370,N_13524,N_13627);
or U14371 (N_14371,N_13831,N_13963);
xnor U14372 (N_14372,N_14249,N_13587);
and U14373 (N_14373,N_13927,N_13813);
or U14374 (N_14374,N_13845,N_13882);
or U14375 (N_14375,N_13606,N_13500);
xor U14376 (N_14376,N_14228,N_13946);
nand U14377 (N_14377,N_14170,N_14150);
nor U14378 (N_14378,N_14241,N_13983);
xnor U14379 (N_14379,N_14203,N_13598);
or U14380 (N_14380,N_13884,N_14237);
or U14381 (N_14381,N_13590,N_13804);
nor U14382 (N_14382,N_14214,N_14159);
or U14383 (N_14383,N_14066,N_13694);
nand U14384 (N_14384,N_13533,N_13881);
nand U14385 (N_14385,N_13857,N_13980);
xor U14386 (N_14386,N_13685,N_13866);
nand U14387 (N_14387,N_13581,N_13592);
nand U14388 (N_14388,N_13780,N_13952);
nor U14389 (N_14389,N_13970,N_14164);
or U14390 (N_14390,N_13623,N_13645);
or U14391 (N_14391,N_14063,N_14166);
xor U14392 (N_14392,N_14174,N_13566);
or U14393 (N_14393,N_13526,N_14098);
xor U14394 (N_14394,N_14173,N_13971);
nor U14395 (N_14395,N_13705,N_13879);
and U14396 (N_14396,N_13510,N_13693);
or U14397 (N_14397,N_13738,N_14042);
nand U14398 (N_14398,N_13907,N_14134);
or U14399 (N_14399,N_13841,N_13537);
nand U14400 (N_14400,N_14012,N_14224);
and U14401 (N_14401,N_13692,N_14047);
nand U14402 (N_14402,N_13817,N_14010);
or U14403 (N_14403,N_13911,N_13735);
or U14404 (N_14404,N_13838,N_14125);
xor U14405 (N_14405,N_14188,N_13502);
nand U14406 (N_14406,N_13737,N_13747);
nand U14407 (N_14407,N_14053,N_13774);
nor U14408 (N_14408,N_14179,N_13540);
nand U14409 (N_14409,N_14160,N_13632);
xor U14410 (N_14410,N_13553,N_13903);
and U14411 (N_14411,N_14141,N_14240);
or U14412 (N_14412,N_13965,N_13814);
nand U14413 (N_14413,N_13531,N_13878);
and U14414 (N_14414,N_13714,N_13852);
nor U14415 (N_14415,N_13889,N_14014);
nor U14416 (N_14416,N_13543,N_13988);
nor U14417 (N_14417,N_13959,N_13815);
xor U14418 (N_14418,N_13924,N_14090);
nor U14419 (N_14419,N_13545,N_13716);
nand U14420 (N_14420,N_14145,N_13939);
nand U14421 (N_14421,N_13710,N_14051);
nand U14422 (N_14422,N_13877,N_13961);
nor U14423 (N_14423,N_13895,N_14039);
or U14424 (N_14424,N_13846,N_13826);
nor U14425 (N_14425,N_14101,N_14074);
and U14426 (N_14426,N_13835,N_14106);
nor U14427 (N_14427,N_14087,N_13630);
nand U14428 (N_14428,N_14236,N_13518);
nand U14429 (N_14429,N_13736,N_14103);
or U14430 (N_14430,N_13978,N_13791);
nor U14431 (N_14431,N_14144,N_13824);
xnor U14432 (N_14432,N_13994,N_14050);
nor U14433 (N_14433,N_14022,N_14231);
and U14434 (N_14434,N_13599,N_14226);
and U14435 (N_14435,N_13652,N_13863);
nor U14436 (N_14436,N_14248,N_13883);
nand U14437 (N_14437,N_13748,N_13893);
nand U14438 (N_14438,N_14157,N_13672);
nor U14439 (N_14439,N_13894,N_14076);
or U14440 (N_14440,N_13585,N_13535);
nand U14441 (N_14441,N_13995,N_13573);
xnor U14442 (N_14442,N_13677,N_14181);
or U14443 (N_14443,N_13745,N_14086);
xor U14444 (N_14444,N_14043,N_13517);
and U14445 (N_14445,N_13648,N_13847);
nand U14446 (N_14446,N_13696,N_13577);
xnor U14447 (N_14447,N_13516,N_13731);
or U14448 (N_14448,N_14239,N_14021);
xnor U14449 (N_14449,N_13608,N_13664);
xor U14450 (N_14450,N_14139,N_14102);
nand U14451 (N_14451,N_14112,N_13975);
xor U14452 (N_14452,N_13687,N_14215);
nor U14453 (N_14453,N_13914,N_13762);
and U14454 (N_14454,N_14029,N_13653);
nand U14455 (N_14455,N_13887,N_13853);
nand U14456 (N_14456,N_14242,N_13897);
or U14457 (N_14457,N_13820,N_13605);
xnor U14458 (N_14458,N_13968,N_13670);
and U14459 (N_14459,N_14189,N_13976);
xnor U14460 (N_14460,N_14210,N_13617);
or U14461 (N_14461,N_14096,N_13987);
xor U14462 (N_14462,N_13832,N_13578);
xor U14463 (N_14463,N_13646,N_14138);
nand U14464 (N_14464,N_14225,N_13712);
or U14465 (N_14465,N_14161,N_13875);
and U14466 (N_14466,N_13549,N_13773);
and U14467 (N_14467,N_13799,N_14220);
or U14468 (N_14468,N_14110,N_14093);
xnor U14469 (N_14469,N_13718,N_14099);
nand U14470 (N_14470,N_13711,N_14072);
or U14471 (N_14471,N_13671,N_13982);
nand U14472 (N_14472,N_13691,N_14182);
or U14473 (N_14473,N_13668,N_13570);
or U14474 (N_14474,N_13834,N_13888);
nand U14475 (N_14475,N_14036,N_13900);
or U14476 (N_14476,N_14213,N_13675);
nor U14477 (N_14477,N_14100,N_13862);
nor U14478 (N_14478,N_13964,N_13786);
xor U14479 (N_14479,N_13873,N_13967);
nand U14480 (N_14480,N_13854,N_13842);
nor U14481 (N_14481,N_14130,N_13811);
and U14482 (N_14482,N_13908,N_13641);
nand U14483 (N_14483,N_14167,N_14077);
nand U14484 (N_14484,N_14219,N_13724);
or U14485 (N_14485,N_13586,N_13542);
xnor U14486 (N_14486,N_13999,N_13947);
nor U14487 (N_14487,N_13611,N_13575);
xor U14488 (N_14488,N_13695,N_13742);
nor U14489 (N_14489,N_13557,N_13867);
or U14490 (N_14490,N_13954,N_13969);
and U14491 (N_14491,N_13622,N_13891);
and U14492 (N_14492,N_14154,N_13770);
nand U14493 (N_14493,N_13639,N_13582);
and U14494 (N_14494,N_13776,N_14003);
and U14495 (N_14495,N_14238,N_13979);
and U14496 (N_14496,N_13808,N_14221);
nand U14497 (N_14497,N_14104,N_13626);
or U14498 (N_14498,N_13956,N_13759);
nand U14499 (N_14499,N_13807,N_13825);
nor U14500 (N_14500,N_13901,N_13752);
or U14501 (N_14501,N_13929,N_13683);
or U14502 (N_14502,N_13567,N_13905);
xnor U14503 (N_14503,N_13525,N_13816);
nand U14504 (N_14504,N_14105,N_14030);
or U14505 (N_14505,N_14009,N_13728);
or U14506 (N_14506,N_13953,N_14024);
nor U14507 (N_14507,N_13620,N_14244);
nor U14508 (N_14508,N_14207,N_13583);
nand U14509 (N_14509,N_13876,N_14124);
nand U14510 (N_14510,N_13915,N_14070);
xnor U14511 (N_14511,N_13840,N_13564);
nand U14512 (N_14512,N_13871,N_14069);
nor U14513 (N_14513,N_14019,N_14034);
nand U14514 (N_14514,N_13669,N_13654);
or U14515 (N_14515,N_13756,N_13950);
nand U14516 (N_14516,N_13719,N_13534);
xor U14517 (N_14517,N_14056,N_13909);
nand U14518 (N_14518,N_14071,N_14059);
xnor U14519 (N_14519,N_13576,N_13839);
and U14520 (N_14520,N_13729,N_13506);
nand U14521 (N_14521,N_13614,N_13530);
nor U14522 (N_14522,N_13741,N_13715);
nor U14523 (N_14523,N_13684,N_13720);
nor U14524 (N_14524,N_14196,N_13789);
and U14525 (N_14525,N_14227,N_13655);
and U14526 (N_14526,N_14229,N_13634);
xor U14527 (N_14527,N_13631,N_13574);
xor U14528 (N_14528,N_13944,N_13513);
nor U14529 (N_14529,N_14133,N_13843);
nor U14530 (N_14530,N_14158,N_13597);
xnor U14531 (N_14531,N_13744,N_14184);
nor U14532 (N_14532,N_13916,N_14143);
or U14533 (N_14533,N_13647,N_13635);
nand U14534 (N_14534,N_13827,N_14178);
xor U14535 (N_14535,N_14004,N_13594);
xnor U14536 (N_14536,N_14119,N_13700);
nand U14537 (N_14537,N_14216,N_13880);
and U14538 (N_14538,N_13769,N_13722);
xnor U14539 (N_14539,N_13689,N_13962);
nor U14540 (N_14540,N_13501,N_14017);
nand U14541 (N_14541,N_14140,N_14061);
and U14542 (N_14542,N_13595,N_13610);
xnor U14543 (N_14543,N_14046,N_14023);
nand U14544 (N_14544,N_13607,N_13919);
xnor U14545 (N_14545,N_13746,N_14049);
or U14546 (N_14546,N_13771,N_13559);
or U14547 (N_14547,N_13580,N_13511);
or U14548 (N_14548,N_13793,N_13733);
xnor U14549 (N_14549,N_13616,N_13755);
nor U14550 (N_14550,N_13730,N_13936);
or U14551 (N_14551,N_14234,N_13795);
nand U14552 (N_14552,N_13538,N_13955);
xor U14553 (N_14553,N_14197,N_14152);
nand U14554 (N_14554,N_13717,N_13713);
nor U14555 (N_14555,N_13621,N_14176);
xnor U14556 (N_14556,N_13554,N_13912);
nor U14557 (N_14557,N_13512,N_13618);
and U14558 (N_14558,N_14120,N_14095);
or U14559 (N_14559,N_13612,N_13763);
or U14560 (N_14560,N_14013,N_13930);
and U14561 (N_14561,N_14243,N_13561);
and U14562 (N_14562,N_14065,N_14075);
nand U14563 (N_14563,N_14149,N_13649);
xnor U14564 (N_14564,N_14233,N_13682);
xnor U14565 (N_14565,N_13536,N_13818);
nor U14566 (N_14566,N_13885,N_14246);
xor U14567 (N_14567,N_13898,N_13609);
nor U14568 (N_14568,N_13662,N_13977);
nand U14569 (N_14569,N_13937,N_14082);
or U14570 (N_14570,N_13706,N_13707);
or U14571 (N_14571,N_14153,N_13997);
nor U14572 (N_14572,N_13945,N_13855);
xnor U14573 (N_14573,N_13562,N_14183);
xnor U14574 (N_14574,N_14045,N_13902);
nand U14575 (N_14575,N_13806,N_13702);
nand U14576 (N_14576,N_14041,N_13686);
xnor U14577 (N_14577,N_14212,N_14107);
nor U14578 (N_14578,N_14200,N_14097);
nor U14579 (N_14579,N_13588,N_14052);
or U14580 (N_14580,N_14198,N_14223);
or U14581 (N_14581,N_13874,N_14193);
and U14582 (N_14582,N_14136,N_13960);
nand U14583 (N_14583,N_13766,N_13768);
and U14584 (N_14584,N_14146,N_13698);
and U14585 (N_14585,N_13579,N_13734);
xnor U14586 (N_14586,N_13519,N_14218);
and U14587 (N_14587,N_14114,N_13674);
or U14588 (N_14588,N_14132,N_13779);
nand U14589 (N_14589,N_14062,N_13941);
nor U14590 (N_14590,N_13801,N_13821);
nor U14591 (N_14591,N_13550,N_13681);
nand U14592 (N_14592,N_14018,N_13951);
and U14593 (N_14593,N_13829,N_14208);
xnor U14594 (N_14594,N_14205,N_13708);
nor U14595 (N_14595,N_13989,N_13591);
or U14596 (N_14596,N_13991,N_13661);
nand U14597 (N_14597,N_13757,N_14088);
nand U14598 (N_14598,N_13869,N_13515);
xor U14599 (N_14599,N_13805,N_13798);
xor U14600 (N_14600,N_13725,N_14194);
xor U14601 (N_14601,N_13765,N_13709);
nor U14602 (N_14602,N_13836,N_13942);
and U14603 (N_14603,N_13563,N_13697);
and U14604 (N_14604,N_13860,N_14001);
or U14605 (N_14605,N_13872,N_13568);
and U14606 (N_14606,N_13958,N_14247);
xnor U14607 (N_14607,N_14025,N_14151);
and U14608 (N_14608,N_13596,N_13904);
xnor U14609 (N_14609,N_13858,N_13572);
nand U14610 (N_14610,N_13943,N_13935);
nand U14611 (N_14611,N_14222,N_14060);
nand U14612 (N_14612,N_13749,N_14195);
xor U14613 (N_14613,N_14118,N_13990);
nor U14614 (N_14614,N_14115,N_13678);
or U14615 (N_14615,N_13651,N_14123);
or U14616 (N_14616,N_13993,N_13520);
and U14617 (N_14617,N_14028,N_13892);
nor U14618 (N_14618,N_14230,N_13665);
and U14619 (N_14619,N_13966,N_14127);
nand U14620 (N_14620,N_13948,N_13529);
or U14621 (N_14621,N_14000,N_13619);
or U14622 (N_14622,N_13812,N_14168);
nand U14623 (N_14623,N_13701,N_13629);
and U14624 (N_14624,N_13541,N_14177);
nand U14625 (N_14625,N_13835,N_14001);
nand U14626 (N_14626,N_14066,N_14207);
and U14627 (N_14627,N_13626,N_13561);
and U14628 (N_14628,N_13604,N_13597);
nand U14629 (N_14629,N_13973,N_14161);
or U14630 (N_14630,N_13727,N_13554);
nor U14631 (N_14631,N_13817,N_13702);
nor U14632 (N_14632,N_13667,N_14208);
or U14633 (N_14633,N_13862,N_13732);
nand U14634 (N_14634,N_13705,N_13785);
or U14635 (N_14635,N_13862,N_13544);
nand U14636 (N_14636,N_13881,N_14109);
nand U14637 (N_14637,N_14169,N_13825);
and U14638 (N_14638,N_13519,N_13973);
or U14639 (N_14639,N_13816,N_13966);
xnor U14640 (N_14640,N_13908,N_14200);
or U14641 (N_14641,N_13903,N_14085);
nand U14642 (N_14642,N_13913,N_13630);
and U14643 (N_14643,N_14125,N_14077);
nor U14644 (N_14644,N_13911,N_14078);
xor U14645 (N_14645,N_13617,N_14168);
and U14646 (N_14646,N_13583,N_13888);
nor U14647 (N_14647,N_13966,N_14092);
nor U14648 (N_14648,N_13990,N_14033);
or U14649 (N_14649,N_14176,N_13875);
nor U14650 (N_14650,N_13640,N_13967);
nand U14651 (N_14651,N_13701,N_13585);
nand U14652 (N_14652,N_14234,N_14097);
and U14653 (N_14653,N_13703,N_13547);
nor U14654 (N_14654,N_13587,N_14093);
nand U14655 (N_14655,N_13754,N_14043);
nand U14656 (N_14656,N_13617,N_13665);
nand U14657 (N_14657,N_13798,N_14209);
or U14658 (N_14658,N_13862,N_14164);
nand U14659 (N_14659,N_13872,N_13690);
or U14660 (N_14660,N_14005,N_14112);
and U14661 (N_14661,N_14067,N_14040);
or U14662 (N_14662,N_13508,N_14201);
and U14663 (N_14663,N_14165,N_13533);
nor U14664 (N_14664,N_13917,N_13995);
and U14665 (N_14665,N_14042,N_13885);
or U14666 (N_14666,N_14074,N_13652);
nand U14667 (N_14667,N_13832,N_14052);
and U14668 (N_14668,N_14016,N_13721);
or U14669 (N_14669,N_13732,N_14033);
nand U14670 (N_14670,N_14100,N_14182);
nand U14671 (N_14671,N_14086,N_13651);
nor U14672 (N_14672,N_13947,N_14232);
nand U14673 (N_14673,N_14132,N_14018);
nor U14674 (N_14674,N_13524,N_13637);
nor U14675 (N_14675,N_14240,N_13964);
nor U14676 (N_14676,N_13812,N_13657);
nand U14677 (N_14677,N_13706,N_13650);
or U14678 (N_14678,N_13655,N_14238);
nand U14679 (N_14679,N_13928,N_13734);
nand U14680 (N_14680,N_14185,N_13543);
xnor U14681 (N_14681,N_14154,N_14189);
nor U14682 (N_14682,N_13965,N_14115);
and U14683 (N_14683,N_14157,N_13886);
or U14684 (N_14684,N_14173,N_13972);
nor U14685 (N_14685,N_13980,N_13839);
xnor U14686 (N_14686,N_14040,N_14037);
and U14687 (N_14687,N_14078,N_13940);
or U14688 (N_14688,N_13776,N_13922);
nor U14689 (N_14689,N_14230,N_13676);
and U14690 (N_14690,N_13907,N_13940);
nor U14691 (N_14691,N_13851,N_14111);
nand U14692 (N_14692,N_13852,N_13848);
xor U14693 (N_14693,N_13774,N_13770);
and U14694 (N_14694,N_14023,N_14066);
xor U14695 (N_14695,N_13893,N_13608);
nand U14696 (N_14696,N_14143,N_14121);
or U14697 (N_14697,N_14173,N_13989);
or U14698 (N_14698,N_13990,N_13596);
nand U14699 (N_14699,N_14198,N_13547);
nor U14700 (N_14700,N_13651,N_13516);
and U14701 (N_14701,N_13653,N_14049);
nor U14702 (N_14702,N_13786,N_13604);
nand U14703 (N_14703,N_14127,N_13531);
xnor U14704 (N_14704,N_13545,N_13877);
xnor U14705 (N_14705,N_14041,N_13924);
or U14706 (N_14706,N_14223,N_14218);
or U14707 (N_14707,N_13641,N_14014);
nor U14708 (N_14708,N_13881,N_13608);
nor U14709 (N_14709,N_14235,N_13635);
xnor U14710 (N_14710,N_14199,N_14082);
xnor U14711 (N_14711,N_13894,N_13982);
and U14712 (N_14712,N_14160,N_13917);
nand U14713 (N_14713,N_13605,N_13771);
xor U14714 (N_14714,N_13623,N_14227);
xor U14715 (N_14715,N_13651,N_13727);
nand U14716 (N_14716,N_13767,N_13929);
or U14717 (N_14717,N_13574,N_13690);
and U14718 (N_14718,N_13648,N_13746);
and U14719 (N_14719,N_13581,N_13672);
xnor U14720 (N_14720,N_13671,N_14136);
and U14721 (N_14721,N_14125,N_13670);
and U14722 (N_14722,N_13817,N_13966);
and U14723 (N_14723,N_14040,N_13619);
nand U14724 (N_14724,N_13518,N_13766);
nor U14725 (N_14725,N_13697,N_14094);
and U14726 (N_14726,N_13825,N_14210);
nor U14727 (N_14727,N_13859,N_14012);
and U14728 (N_14728,N_14171,N_13667);
and U14729 (N_14729,N_13788,N_13668);
nand U14730 (N_14730,N_14211,N_13946);
nor U14731 (N_14731,N_13875,N_13569);
and U14732 (N_14732,N_13833,N_13965);
nor U14733 (N_14733,N_13609,N_14009);
nor U14734 (N_14734,N_14090,N_14248);
nor U14735 (N_14735,N_13985,N_13856);
nor U14736 (N_14736,N_14207,N_14103);
nand U14737 (N_14737,N_13849,N_13816);
nand U14738 (N_14738,N_14009,N_14065);
xor U14739 (N_14739,N_13757,N_14031);
or U14740 (N_14740,N_13854,N_13889);
or U14741 (N_14741,N_13651,N_14163);
and U14742 (N_14742,N_13632,N_13948);
nand U14743 (N_14743,N_14222,N_14035);
or U14744 (N_14744,N_13729,N_14183);
nor U14745 (N_14745,N_14113,N_14013);
and U14746 (N_14746,N_14241,N_13825);
or U14747 (N_14747,N_13872,N_14115);
nand U14748 (N_14748,N_13575,N_13743);
nor U14749 (N_14749,N_13950,N_14182);
nor U14750 (N_14750,N_13789,N_14012);
xnor U14751 (N_14751,N_14060,N_13780);
and U14752 (N_14752,N_13828,N_14190);
or U14753 (N_14753,N_14234,N_13623);
or U14754 (N_14754,N_14183,N_13888);
xor U14755 (N_14755,N_14182,N_14218);
and U14756 (N_14756,N_13855,N_13546);
and U14757 (N_14757,N_13527,N_14244);
nor U14758 (N_14758,N_13535,N_13889);
nor U14759 (N_14759,N_13835,N_13632);
nor U14760 (N_14760,N_13651,N_13515);
and U14761 (N_14761,N_14083,N_14211);
or U14762 (N_14762,N_13820,N_13909);
or U14763 (N_14763,N_14150,N_14198);
nand U14764 (N_14764,N_13953,N_13682);
xor U14765 (N_14765,N_13957,N_13700);
and U14766 (N_14766,N_13616,N_14045);
xor U14767 (N_14767,N_13565,N_13526);
and U14768 (N_14768,N_13754,N_14223);
nand U14769 (N_14769,N_13536,N_14186);
nand U14770 (N_14770,N_13639,N_14142);
and U14771 (N_14771,N_13940,N_13671);
or U14772 (N_14772,N_13990,N_14229);
and U14773 (N_14773,N_14092,N_13550);
nand U14774 (N_14774,N_13660,N_13859);
nand U14775 (N_14775,N_13984,N_13799);
nor U14776 (N_14776,N_14243,N_14087);
xor U14777 (N_14777,N_14184,N_14131);
nor U14778 (N_14778,N_14055,N_14144);
or U14779 (N_14779,N_13881,N_14218);
nand U14780 (N_14780,N_14076,N_13563);
or U14781 (N_14781,N_13734,N_14175);
nand U14782 (N_14782,N_14179,N_14035);
nand U14783 (N_14783,N_14037,N_14076);
xnor U14784 (N_14784,N_13872,N_13821);
nor U14785 (N_14785,N_13860,N_13996);
and U14786 (N_14786,N_13598,N_14174);
nand U14787 (N_14787,N_13809,N_13827);
and U14788 (N_14788,N_14229,N_14137);
or U14789 (N_14789,N_14016,N_14096);
or U14790 (N_14790,N_13514,N_14062);
nor U14791 (N_14791,N_14134,N_14078);
or U14792 (N_14792,N_13940,N_14233);
or U14793 (N_14793,N_13517,N_13791);
and U14794 (N_14794,N_14113,N_13618);
and U14795 (N_14795,N_14140,N_13595);
and U14796 (N_14796,N_14013,N_14210);
nand U14797 (N_14797,N_13515,N_13742);
nand U14798 (N_14798,N_13684,N_14084);
nor U14799 (N_14799,N_13968,N_13839);
and U14800 (N_14800,N_14012,N_14235);
nand U14801 (N_14801,N_13884,N_13761);
or U14802 (N_14802,N_13660,N_13712);
or U14803 (N_14803,N_14019,N_14040);
nand U14804 (N_14804,N_14094,N_14138);
or U14805 (N_14805,N_13661,N_13920);
and U14806 (N_14806,N_13628,N_13753);
xor U14807 (N_14807,N_13640,N_14038);
xnor U14808 (N_14808,N_13820,N_14011);
xnor U14809 (N_14809,N_13862,N_13629);
xnor U14810 (N_14810,N_13546,N_14216);
nand U14811 (N_14811,N_13556,N_14115);
or U14812 (N_14812,N_13525,N_13833);
or U14813 (N_14813,N_13875,N_13836);
and U14814 (N_14814,N_13610,N_14068);
and U14815 (N_14815,N_13696,N_13849);
and U14816 (N_14816,N_13802,N_13882);
xnor U14817 (N_14817,N_13864,N_14119);
and U14818 (N_14818,N_13802,N_13778);
nor U14819 (N_14819,N_13710,N_14050);
nand U14820 (N_14820,N_13571,N_14216);
and U14821 (N_14821,N_14003,N_14222);
xnor U14822 (N_14822,N_13786,N_14098);
xnor U14823 (N_14823,N_14195,N_14072);
nand U14824 (N_14824,N_13628,N_13781);
xor U14825 (N_14825,N_14077,N_13725);
nor U14826 (N_14826,N_14217,N_13706);
nor U14827 (N_14827,N_13942,N_14248);
nand U14828 (N_14828,N_14129,N_13999);
xor U14829 (N_14829,N_13639,N_14195);
nand U14830 (N_14830,N_13796,N_14242);
nor U14831 (N_14831,N_13853,N_14084);
and U14832 (N_14832,N_13951,N_13894);
nand U14833 (N_14833,N_13682,N_13729);
nor U14834 (N_14834,N_14199,N_13757);
and U14835 (N_14835,N_13914,N_14058);
nand U14836 (N_14836,N_14151,N_14037);
nand U14837 (N_14837,N_14002,N_13818);
nand U14838 (N_14838,N_14239,N_13729);
and U14839 (N_14839,N_13776,N_13715);
or U14840 (N_14840,N_13854,N_13527);
xor U14841 (N_14841,N_14009,N_13559);
nand U14842 (N_14842,N_13816,N_13819);
nand U14843 (N_14843,N_13544,N_13627);
or U14844 (N_14844,N_14145,N_13856);
nor U14845 (N_14845,N_13730,N_13569);
or U14846 (N_14846,N_14077,N_13994);
or U14847 (N_14847,N_13689,N_13857);
and U14848 (N_14848,N_13712,N_14183);
nor U14849 (N_14849,N_14204,N_13932);
xor U14850 (N_14850,N_13554,N_13576);
nand U14851 (N_14851,N_13739,N_13780);
xor U14852 (N_14852,N_14148,N_14112);
nor U14853 (N_14853,N_14178,N_13532);
nor U14854 (N_14854,N_13724,N_14227);
and U14855 (N_14855,N_13783,N_14025);
or U14856 (N_14856,N_13533,N_13850);
and U14857 (N_14857,N_13739,N_13851);
xor U14858 (N_14858,N_13894,N_14174);
or U14859 (N_14859,N_13948,N_13868);
xnor U14860 (N_14860,N_13731,N_13761);
nand U14861 (N_14861,N_13508,N_14226);
nand U14862 (N_14862,N_13864,N_14199);
nand U14863 (N_14863,N_13809,N_13585);
xor U14864 (N_14864,N_13717,N_13825);
xnor U14865 (N_14865,N_13708,N_13790);
nor U14866 (N_14866,N_13748,N_14089);
xor U14867 (N_14867,N_13818,N_14092);
or U14868 (N_14868,N_14141,N_13811);
or U14869 (N_14869,N_13970,N_13622);
xor U14870 (N_14870,N_13819,N_13532);
nor U14871 (N_14871,N_13838,N_14149);
and U14872 (N_14872,N_13544,N_13629);
nor U14873 (N_14873,N_14128,N_13882);
xor U14874 (N_14874,N_14234,N_13977);
nor U14875 (N_14875,N_13882,N_13764);
nand U14876 (N_14876,N_13879,N_13809);
nor U14877 (N_14877,N_14178,N_13880);
and U14878 (N_14878,N_14206,N_14091);
xnor U14879 (N_14879,N_13598,N_13664);
nor U14880 (N_14880,N_13655,N_14182);
xnor U14881 (N_14881,N_14078,N_13860);
nor U14882 (N_14882,N_14087,N_13579);
and U14883 (N_14883,N_14131,N_13880);
xnor U14884 (N_14884,N_13893,N_13655);
or U14885 (N_14885,N_14169,N_13783);
xnor U14886 (N_14886,N_14008,N_13857);
nand U14887 (N_14887,N_13764,N_13730);
xor U14888 (N_14888,N_14126,N_14206);
or U14889 (N_14889,N_13791,N_13854);
xnor U14890 (N_14890,N_13909,N_14111);
or U14891 (N_14891,N_14004,N_14093);
xor U14892 (N_14892,N_13525,N_14152);
xor U14893 (N_14893,N_13969,N_13603);
nand U14894 (N_14894,N_13999,N_13655);
nor U14895 (N_14895,N_13598,N_13994);
and U14896 (N_14896,N_14235,N_13676);
nand U14897 (N_14897,N_13955,N_13824);
xor U14898 (N_14898,N_13578,N_14091);
or U14899 (N_14899,N_13760,N_13972);
or U14900 (N_14900,N_13773,N_14153);
xnor U14901 (N_14901,N_13760,N_14188);
and U14902 (N_14902,N_13736,N_14176);
nor U14903 (N_14903,N_13918,N_14178);
xor U14904 (N_14904,N_13810,N_13857);
or U14905 (N_14905,N_14236,N_13711);
or U14906 (N_14906,N_13733,N_13947);
and U14907 (N_14907,N_13682,N_13669);
and U14908 (N_14908,N_14017,N_13507);
or U14909 (N_14909,N_14084,N_13921);
nand U14910 (N_14910,N_13932,N_14102);
xnor U14911 (N_14911,N_13534,N_13985);
nor U14912 (N_14912,N_13645,N_14189);
nor U14913 (N_14913,N_14191,N_14115);
nand U14914 (N_14914,N_13875,N_13898);
and U14915 (N_14915,N_13521,N_13967);
and U14916 (N_14916,N_13747,N_14182);
xor U14917 (N_14917,N_13712,N_14021);
nand U14918 (N_14918,N_13878,N_13965);
nand U14919 (N_14919,N_13693,N_13888);
nand U14920 (N_14920,N_14215,N_14146);
nand U14921 (N_14921,N_13874,N_13970);
and U14922 (N_14922,N_14104,N_14018);
and U14923 (N_14923,N_14013,N_13583);
and U14924 (N_14924,N_13990,N_13722);
nand U14925 (N_14925,N_13792,N_13769);
xnor U14926 (N_14926,N_13579,N_14028);
xor U14927 (N_14927,N_13705,N_13561);
and U14928 (N_14928,N_14237,N_13668);
and U14929 (N_14929,N_13777,N_13598);
xnor U14930 (N_14930,N_13940,N_14113);
and U14931 (N_14931,N_13552,N_13521);
xor U14932 (N_14932,N_13956,N_14158);
and U14933 (N_14933,N_13684,N_14201);
and U14934 (N_14934,N_14222,N_13989);
or U14935 (N_14935,N_13619,N_13740);
nor U14936 (N_14936,N_14193,N_13673);
nand U14937 (N_14937,N_13853,N_13625);
nand U14938 (N_14938,N_13810,N_13828);
nand U14939 (N_14939,N_13514,N_13568);
xor U14940 (N_14940,N_13914,N_13898);
nand U14941 (N_14941,N_13918,N_13601);
nand U14942 (N_14942,N_14244,N_13743);
nand U14943 (N_14943,N_14086,N_13954);
xnor U14944 (N_14944,N_13972,N_14203);
nor U14945 (N_14945,N_13582,N_14072);
nor U14946 (N_14946,N_13850,N_14138);
xor U14947 (N_14947,N_14160,N_14247);
nand U14948 (N_14948,N_14206,N_14089);
or U14949 (N_14949,N_13725,N_13690);
or U14950 (N_14950,N_14141,N_13741);
nor U14951 (N_14951,N_13701,N_14111);
nand U14952 (N_14952,N_14231,N_14128);
nor U14953 (N_14953,N_13639,N_14211);
xor U14954 (N_14954,N_14051,N_14106);
nor U14955 (N_14955,N_14111,N_13597);
or U14956 (N_14956,N_13616,N_14110);
xnor U14957 (N_14957,N_14201,N_13976);
and U14958 (N_14958,N_14180,N_13879);
and U14959 (N_14959,N_13895,N_13507);
nor U14960 (N_14960,N_13509,N_13947);
and U14961 (N_14961,N_14218,N_14007);
nor U14962 (N_14962,N_14021,N_14056);
nor U14963 (N_14963,N_13869,N_14211);
nand U14964 (N_14964,N_13922,N_14214);
nor U14965 (N_14965,N_13682,N_14077);
xor U14966 (N_14966,N_13706,N_13646);
nand U14967 (N_14967,N_13784,N_13686);
nand U14968 (N_14968,N_13978,N_13948);
nor U14969 (N_14969,N_14249,N_13755);
nand U14970 (N_14970,N_14231,N_13629);
nand U14971 (N_14971,N_13974,N_14188);
or U14972 (N_14972,N_13850,N_14003);
and U14973 (N_14973,N_13791,N_13995);
nor U14974 (N_14974,N_13772,N_13981);
or U14975 (N_14975,N_13549,N_14099);
nand U14976 (N_14976,N_13515,N_13600);
nor U14977 (N_14977,N_13603,N_13700);
or U14978 (N_14978,N_14218,N_14185);
nand U14979 (N_14979,N_13511,N_13880);
nor U14980 (N_14980,N_13998,N_13681);
nor U14981 (N_14981,N_13737,N_13509);
xnor U14982 (N_14982,N_13533,N_13895);
xnor U14983 (N_14983,N_13948,N_14020);
or U14984 (N_14984,N_14114,N_14036);
and U14985 (N_14985,N_13753,N_13968);
nand U14986 (N_14986,N_13806,N_13602);
and U14987 (N_14987,N_13890,N_13751);
and U14988 (N_14988,N_14229,N_13724);
nor U14989 (N_14989,N_13783,N_14245);
nand U14990 (N_14990,N_14048,N_14089);
xor U14991 (N_14991,N_13968,N_13653);
nand U14992 (N_14992,N_14007,N_13834);
and U14993 (N_14993,N_14119,N_14226);
xor U14994 (N_14994,N_13753,N_13726);
and U14995 (N_14995,N_14061,N_13922);
nand U14996 (N_14996,N_13577,N_14006);
xor U14997 (N_14997,N_13821,N_13781);
nor U14998 (N_14998,N_13847,N_13774);
xor U14999 (N_14999,N_14202,N_14156);
xnor UO_0 (O_0,N_14543,N_14514);
xor UO_1 (O_1,N_14260,N_14721);
and UO_2 (O_2,N_14571,N_14653);
nand UO_3 (O_3,N_14912,N_14977);
nor UO_4 (O_4,N_14434,N_14658);
and UO_5 (O_5,N_14454,N_14779);
nor UO_6 (O_6,N_14594,N_14686);
or UO_7 (O_7,N_14362,N_14832);
xnor UO_8 (O_8,N_14901,N_14361);
nand UO_9 (O_9,N_14678,N_14944);
or UO_10 (O_10,N_14371,N_14964);
or UO_11 (O_11,N_14682,N_14513);
or UO_12 (O_12,N_14845,N_14254);
and UO_13 (O_13,N_14324,N_14689);
xor UO_14 (O_14,N_14458,N_14975);
nand UO_15 (O_15,N_14479,N_14711);
xor UO_16 (O_16,N_14992,N_14877);
nor UO_17 (O_17,N_14432,N_14282);
nand UO_18 (O_18,N_14546,N_14367);
nor UO_19 (O_19,N_14549,N_14635);
and UO_20 (O_20,N_14690,N_14843);
and UO_21 (O_21,N_14378,N_14696);
and UO_22 (O_22,N_14355,N_14486);
or UO_23 (O_23,N_14259,N_14803);
nand UO_24 (O_24,N_14311,N_14900);
or UO_25 (O_25,N_14467,N_14291);
nor UO_26 (O_26,N_14786,N_14854);
or UO_27 (O_27,N_14494,N_14328);
nor UO_28 (O_28,N_14895,N_14979);
xor UO_29 (O_29,N_14482,N_14499);
nor UO_30 (O_30,N_14988,N_14524);
or UO_31 (O_31,N_14535,N_14436);
or UO_32 (O_32,N_14794,N_14887);
and UO_33 (O_33,N_14585,N_14489);
and UO_34 (O_34,N_14428,N_14683);
nand UO_35 (O_35,N_14953,N_14749);
or UO_36 (O_36,N_14747,N_14639);
nand UO_37 (O_37,N_14927,N_14627);
or UO_38 (O_38,N_14528,N_14560);
or UO_39 (O_39,N_14706,N_14463);
xnor UO_40 (O_40,N_14984,N_14646);
nor UO_41 (O_41,N_14995,N_14965);
or UO_42 (O_42,N_14466,N_14893);
nor UO_43 (O_43,N_14570,N_14347);
or UO_44 (O_44,N_14892,N_14906);
nand UO_45 (O_45,N_14881,N_14600);
xor UO_46 (O_46,N_14304,N_14265);
nor UO_47 (O_47,N_14716,N_14356);
or UO_48 (O_48,N_14337,N_14309);
xnor UO_49 (O_49,N_14816,N_14937);
nand UO_50 (O_50,N_14338,N_14952);
nand UO_51 (O_51,N_14713,N_14631);
nand UO_52 (O_52,N_14939,N_14709);
nand UO_53 (O_53,N_14303,N_14715);
or UO_54 (O_54,N_14766,N_14760);
and UO_55 (O_55,N_14315,N_14781);
or UO_56 (O_56,N_14392,N_14642);
nand UO_57 (O_57,N_14763,N_14358);
or UO_58 (O_58,N_14508,N_14663);
nand UO_59 (O_59,N_14751,N_14902);
nand UO_60 (O_60,N_14401,N_14496);
xor UO_61 (O_61,N_14262,N_14552);
or UO_62 (O_62,N_14411,N_14638);
and UO_63 (O_63,N_14908,N_14534);
or UO_64 (O_64,N_14830,N_14737);
or UO_65 (O_65,N_14274,N_14435);
nand UO_66 (O_66,N_14504,N_14491);
and UO_67 (O_67,N_14280,N_14502);
nand UO_68 (O_68,N_14530,N_14993);
xnor UO_69 (O_69,N_14461,N_14903);
nor UO_70 (O_70,N_14390,N_14550);
or UO_71 (O_71,N_14628,N_14437);
xnor UO_72 (O_72,N_14576,N_14614);
and UO_73 (O_73,N_14449,N_14354);
nand UO_74 (O_74,N_14778,N_14608);
nand UO_75 (O_75,N_14777,N_14569);
nand UO_76 (O_76,N_14308,N_14776);
or UO_77 (O_77,N_14558,N_14899);
nand UO_78 (O_78,N_14724,N_14462);
nand UO_79 (O_79,N_14429,N_14368);
nand UO_80 (O_80,N_14962,N_14349);
or UO_81 (O_81,N_14343,N_14918);
nand UO_82 (O_82,N_14790,N_14798);
nand UO_83 (O_83,N_14404,N_14645);
xor UO_84 (O_84,N_14531,N_14369);
and UO_85 (O_85,N_14523,N_14862);
nand UO_86 (O_86,N_14915,N_14607);
or UO_87 (O_87,N_14399,N_14292);
and UO_88 (O_88,N_14509,N_14443);
nor UO_89 (O_89,N_14850,N_14863);
nor UO_90 (O_90,N_14933,N_14469);
nor UO_91 (O_91,N_14662,N_14701);
or UO_92 (O_92,N_14660,N_14366);
xnor UO_93 (O_93,N_14305,N_14263);
nor UO_94 (O_94,N_14444,N_14698);
nor UO_95 (O_95,N_14795,N_14791);
xor UO_96 (O_96,N_14882,N_14272);
or UO_97 (O_97,N_14568,N_14426);
or UO_98 (O_98,N_14722,N_14782);
xor UO_99 (O_99,N_14768,N_14270);
and UO_100 (O_100,N_14332,N_14708);
xor UO_101 (O_101,N_14799,N_14420);
or UO_102 (O_102,N_14981,N_14670);
xor UO_103 (O_103,N_14400,N_14527);
nand UO_104 (O_104,N_14307,N_14876);
or UO_105 (O_105,N_14754,N_14409);
nor UO_106 (O_106,N_14478,N_14312);
and UO_107 (O_107,N_14599,N_14865);
nand UO_108 (O_108,N_14870,N_14413);
nand UO_109 (O_109,N_14287,N_14624);
or UO_110 (O_110,N_14376,N_14557);
xor UO_111 (O_111,N_14256,N_14334);
nand UO_112 (O_112,N_14565,N_14976);
nand UO_113 (O_113,N_14397,N_14575);
nand UO_114 (O_114,N_14266,N_14316);
nor UO_115 (O_115,N_14446,N_14252);
nand UO_116 (O_116,N_14745,N_14886);
and UO_117 (O_117,N_14298,N_14440);
nor UO_118 (O_118,N_14561,N_14310);
nor UO_119 (O_119,N_14991,N_14926);
xnor UO_120 (O_120,N_14321,N_14767);
nor UO_121 (O_121,N_14871,N_14325);
and UO_122 (O_122,N_14562,N_14520);
nand UO_123 (O_123,N_14615,N_14849);
nor UO_124 (O_124,N_14342,N_14733);
or UO_125 (O_125,N_14694,N_14921);
nor UO_126 (O_126,N_14774,N_14517);
nand UO_127 (O_127,N_14335,N_14880);
nor UO_128 (O_128,N_14403,N_14406);
or UO_129 (O_129,N_14809,N_14554);
nand UO_130 (O_130,N_14590,N_14536);
and UO_131 (O_131,N_14680,N_14636);
or UO_132 (O_132,N_14924,N_14940);
nor UO_133 (O_133,N_14957,N_14885);
nand UO_134 (O_134,N_14839,N_14718);
nor UO_135 (O_135,N_14472,N_14812);
nor UO_136 (O_136,N_14503,N_14556);
and UO_137 (O_137,N_14883,N_14666);
xnor UO_138 (O_138,N_14932,N_14838);
xor UO_139 (O_139,N_14999,N_14699);
xor UO_140 (O_140,N_14969,N_14542);
or UO_141 (O_141,N_14935,N_14842);
xor UO_142 (O_142,N_14405,N_14492);
or UO_143 (O_143,N_14817,N_14414);
nand UO_144 (O_144,N_14518,N_14761);
nor UO_145 (O_145,N_14821,N_14493);
nand UO_146 (O_146,N_14674,N_14521);
nand UO_147 (O_147,N_14593,N_14978);
nor UO_148 (O_148,N_14584,N_14498);
and UO_149 (O_149,N_14424,N_14574);
nor UO_150 (O_150,N_14460,N_14532);
xnor UO_151 (O_151,N_14384,N_14673);
and UO_152 (O_152,N_14294,N_14986);
nand UO_153 (O_153,N_14652,N_14473);
or UO_154 (O_154,N_14529,N_14769);
or UO_155 (O_155,N_14644,N_14859);
and UO_156 (O_156,N_14375,N_14739);
nor UO_157 (O_157,N_14891,N_14329);
and UO_158 (O_158,N_14951,N_14253);
xnor UO_159 (O_159,N_14829,N_14383);
nand UO_160 (O_160,N_14919,N_14973);
nand UO_161 (O_161,N_14731,N_14650);
nor UO_162 (O_162,N_14505,N_14815);
xor UO_163 (O_163,N_14425,N_14630);
xnor UO_164 (O_164,N_14357,N_14626);
and UO_165 (O_165,N_14474,N_14967);
nand UO_166 (O_166,N_14770,N_14544);
xor UO_167 (O_167,N_14833,N_14925);
nor UO_168 (O_168,N_14909,N_14661);
or UO_169 (O_169,N_14704,N_14758);
nor UO_170 (O_170,N_14998,N_14379);
or UO_171 (O_171,N_14856,N_14664);
or UO_172 (O_172,N_14640,N_14730);
and UO_173 (O_173,N_14789,N_14955);
and UO_174 (O_174,N_14396,N_14910);
and UO_175 (O_175,N_14622,N_14364);
and UO_176 (O_176,N_14623,N_14923);
nor UO_177 (O_177,N_14746,N_14330);
nor UO_178 (O_178,N_14668,N_14852);
or UO_179 (O_179,N_14784,N_14495);
or UO_180 (O_180,N_14966,N_14319);
nor UO_181 (O_181,N_14258,N_14267);
xor UO_182 (O_182,N_14756,N_14643);
and UO_183 (O_183,N_14959,N_14277);
nand UO_184 (O_184,N_14372,N_14867);
nor UO_185 (O_185,N_14388,N_14507);
nor UO_186 (O_186,N_14336,N_14344);
xor UO_187 (O_187,N_14665,N_14936);
and UO_188 (O_188,N_14907,N_14641);
nand UO_189 (O_189,N_14846,N_14823);
and UO_190 (O_190,N_14712,N_14942);
and UO_191 (O_191,N_14780,N_14351);
and UO_192 (O_192,N_14452,N_14723);
or UO_193 (O_193,N_14488,N_14945);
nor UO_194 (O_194,N_14551,N_14395);
or UO_195 (O_195,N_14897,N_14922);
and UO_196 (O_196,N_14717,N_14888);
xor UO_197 (O_197,N_14948,N_14787);
nand UO_198 (O_198,N_14439,N_14416);
nand UO_199 (O_199,N_14296,N_14609);
and UO_200 (O_200,N_14281,N_14759);
and UO_201 (O_201,N_14506,N_14847);
nand UO_202 (O_202,N_14598,N_14511);
or UO_203 (O_203,N_14826,N_14719);
nor UO_204 (O_204,N_14648,N_14592);
nor UO_205 (O_205,N_14914,N_14669);
nor UO_206 (O_206,N_14855,N_14676);
and UO_207 (O_207,N_14385,N_14917);
xnor UO_208 (O_208,N_14483,N_14748);
or UO_209 (O_209,N_14697,N_14251);
xnor UO_210 (O_210,N_14456,N_14587);
nand UO_211 (O_211,N_14755,N_14596);
nand UO_212 (O_212,N_14649,N_14582);
and UO_213 (O_213,N_14430,N_14667);
and UO_214 (O_214,N_14726,N_14647);
nand UO_215 (O_215,N_14374,N_14928);
nand UO_216 (O_216,N_14651,N_14920);
xor UO_217 (O_217,N_14286,N_14657);
nor UO_218 (O_218,N_14875,N_14583);
or UO_219 (O_219,N_14470,N_14792);
xnor UO_220 (O_220,N_14797,N_14941);
or UO_221 (O_221,N_14617,N_14677);
nor UO_222 (O_222,N_14806,N_14453);
xnor UO_223 (O_223,N_14382,N_14365);
nand UO_224 (O_224,N_14611,N_14455);
nor UO_225 (O_225,N_14990,N_14700);
xor UO_226 (O_226,N_14771,N_14533);
xnor UO_227 (O_227,N_14872,N_14632);
or UO_228 (O_228,N_14398,N_14864);
and UO_229 (O_229,N_14970,N_14938);
and UO_230 (O_230,N_14442,N_14788);
nor UO_231 (O_231,N_14417,N_14762);
xor UO_232 (O_232,N_14606,N_14386);
nor UO_233 (O_233,N_14659,N_14916);
and UO_234 (O_234,N_14738,N_14515);
xor UO_235 (O_235,N_14595,N_14820);
nand UO_236 (O_236,N_14289,N_14996);
nand UO_237 (O_237,N_14750,N_14773);
xor UO_238 (O_238,N_14714,N_14702);
xnor UO_239 (O_239,N_14960,N_14475);
and UO_240 (O_240,N_14869,N_14500);
and UO_241 (O_241,N_14484,N_14851);
and UO_242 (O_242,N_14612,N_14873);
xnor UO_243 (O_243,N_14800,N_14370);
nand UO_244 (O_244,N_14539,N_14559);
xor UO_245 (O_245,N_14744,N_14448);
nor UO_246 (O_246,N_14301,N_14320);
and UO_247 (O_247,N_14257,N_14471);
nor UO_248 (O_248,N_14477,N_14346);
or UO_249 (O_249,N_14633,N_14273);
nor UO_250 (O_250,N_14250,N_14510);
nand UO_251 (O_251,N_14950,N_14827);
and UO_252 (O_252,N_14637,N_14468);
or UO_253 (O_253,N_14898,N_14465);
or UO_254 (O_254,N_14537,N_14297);
nor UO_255 (O_255,N_14753,N_14949);
and UO_256 (O_256,N_14360,N_14485);
nor UO_257 (O_257,N_14729,N_14866);
and UO_258 (O_258,N_14983,N_14431);
and UO_259 (O_259,N_14904,N_14419);
nor UO_260 (O_260,N_14878,N_14317);
nor UO_261 (O_261,N_14982,N_14389);
nand UO_262 (O_262,N_14591,N_14629);
nor UO_263 (O_263,N_14808,N_14314);
and UO_264 (O_264,N_14688,N_14684);
nor UO_265 (O_265,N_14743,N_14879);
nand UO_266 (O_266,N_14946,N_14796);
or UO_267 (O_267,N_14736,N_14525);
and UO_268 (O_268,N_14693,N_14943);
xnor UO_269 (O_269,N_14802,N_14433);
nor UO_270 (O_270,N_14497,N_14563);
or UO_271 (O_271,N_14377,N_14963);
nand UO_272 (O_272,N_14819,N_14956);
nor UO_273 (O_273,N_14290,N_14302);
and UO_274 (O_274,N_14828,N_14834);
xnor UO_275 (O_275,N_14734,N_14894);
nand UO_276 (O_276,N_14861,N_14288);
xnor UO_277 (O_277,N_14619,N_14387);
nor UO_278 (O_278,N_14540,N_14727);
nand UO_279 (O_279,N_14415,N_14620);
xor UO_280 (O_280,N_14441,N_14974);
nor UO_281 (O_281,N_14997,N_14402);
nand UO_282 (O_282,N_14326,N_14840);
and UO_283 (O_283,N_14732,N_14853);
nand UO_284 (O_284,N_14874,N_14728);
and UO_285 (O_285,N_14793,N_14427);
or UO_286 (O_286,N_14911,N_14654);
and UO_287 (O_287,N_14476,N_14269);
or UO_288 (O_288,N_14451,N_14545);
nand UO_289 (O_289,N_14857,N_14971);
and UO_290 (O_290,N_14352,N_14487);
nand UO_291 (O_291,N_14564,N_14394);
or UO_292 (O_292,N_14618,N_14421);
nor UO_293 (O_293,N_14516,N_14381);
nor UO_294 (O_294,N_14980,N_14621);
and UO_295 (O_295,N_14264,N_14268);
and UO_296 (O_296,N_14602,N_14822);
xnor UO_297 (O_297,N_14541,N_14577);
xor UO_298 (O_298,N_14300,N_14896);
nor UO_299 (O_299,N_14930,N_14831);
nand UO_300 (O_300,N_14438,N_14597);
nand UO_301 (O_301,N_14450,N_14580);
and UO_302 (O_302,N_14691,N_14407);
or UO_303 (O_303,N_14860,N_14858);
nor UO_304 (O_304,N_14445,N_14695);
nor UO_305 (O_305,N_14801,N_14548);
nor UO_306 (O_306,N_14339,N_14934);
nand UO_307 (O_307,N_14757,N_14824);
xnor UO_308 (O_308,N_14848,N_14785);
and UO_309 (O_309,N_14459,N_14687);
or UO_310 (O_310,N_14566,N_14555);
nor UO_311 (O_311,N_14359,N_14567);
nor UO_312 (O_312,N_14447,N_14586);
and UO_313 (O_313,N_14836,N_14783);
and UO_314 (O_314,N_14835,N_14293);
nor UO_315 (O_315,N_14805,N_14295);
nand UO_316 (O_316,N_14710,N_14634);
xnor UO_317 (O_317,N_14481,N_14276);
xor UO_318 (O_318,N_14306,N_14588);
or UO_319 (O_319,N_14380,N_14603);
nor UO_320 (O_320,N_14807,N_14501);
and UO_321 (O_321,N_14720,N_14775);
nand UO_322 (O_322,N_14547,N_14725);
xor UO_323 (O_323,N_14284,N_14604);
nor UO_324 (O_324,N_14283,N_14605);
nand UO_325 (O_325,N_14679,N_14837);
nand UO_326 (O_326,N_14961,N_14348);
and UO_327 (O_327,N_14613,N_14350);
and UO_328 (O_328,N_14279,N_14804);
nor UO_329 (O_329,N_14323,N_14573);
xor UO_330 (O_330,N_14422,N_14844);
or UO_331 (O_331,N_14519,N_14672);
xor UO_332 (O_332,N_14333,N_14740);
nor UO_333 (O_333,N_14811,N_14681);
xnor UO_334 (O_334,N_14929,N_14905);
or UO_335 (O_335,N_14299,N_14341);
xnor UO_336 (O_336,N_14318,N_14322);
xor UO_337 (O_337,N_14589,N_14581);
nand UO_338 (O_338,N_14313,N_14255);
and UO_339 (O_339,N_14764,N_14331);
and UO_340 (O_340,N_14705,N_14363);
nand UO_341 (O_341,N_14825,N_14958);
nor UO_342 (O_342,N_14579,N_14418);
nand UO_343 (O_343,N_14868,N_14671);
nand UO_344 (O_344,N_14741,N_14572);
nor UO_345 (O_345,N_14735,N_14989);
xnor UO_346 (O_346,N_14765,N_14423);
or UO_347 (O_347,N_14814,N_14692);
or UO_348 (O_348,N_14985,N_14954);
or UO_349 (O_349,N_14410,N_14931);
or UO_350 (O_350,N_14675,N_14707);
and UO_351 (O_351,N_14553,N_14841);
xor UO_352 (O_352,N_14373,N_14464);
and UO_353 (O_353,N_14610,N_14703);
and UO_354 (O_354,N_14813,N_14625);
xor UO_355 (O_355,N_14345,N_14616);
xor UO_356 (O_356,N_14994,N_14278);
xor UO_357 (O_357,N_14480,N_14601);
xor UO_358 (O_358,N_14512,N_14947);
nor UO_359 (O_359,N_14810,N_14685);
or UO_360 (O_360,N_14285,N_14890);
nor UO_361 (O_361,N_14393,N_14526);
xnor UO_362 (O_362,N_14968,N_14340);
nand UO_363 (O_363,N_14457,N_14490);
nor UO_364 (O_364,N_14275,N_14889);
or UO_365 (O_365,N_14271,N_14987);
nor UO_366 (O_366,N_14353,N_14538);
nor UO_367 (O_367,N_14522,N_14656);
or UO_368 (O_368,N_14742,N_14391);
or UO_369 (O_369,N_14818,N_14913);
nor UO_370 (O_370,N_14408,N_14655);
nand UO_371 (O_371,N_14578,N_14972);
nor UO_372 (O_372,N_14752,N_14327);
or UO_373 (O_373,N_14412,N_14884);
or UO_374 (O_374,N_14261,N_14772);
or UO_375 (O_375,N_14771,N_14282);
xnor UO_376 (O_376,N_14607,N_14343);
xnor UO_377 (O_377,N_14664,N_14463);
nor UO_378 (O_378,N_14328,N_14587);
nand UO_379 (O_379,N_14351,N_14722);
xnor UO_380 (O_380,N_14566,N_14650);
or UO_381 (O_381,N_14975,N_14459);
nor UO_382 (O_382,N_14885,N_14535);
or UO_383 (O_383,N_14584,N_14908);
xor UO_384 (O_384,N_14918,N_14805);
xnor UO_385 (O_385,N_14338,N_14599);
xor UO_386 (O_386,N_14882,N_14618);
xnor UO_387 (O_387,N_14588,N_14752);
and UO_388 (O_388,N_14913,N_14605);
or UO_389 (O_389,N_14733,N_14596);
nor UO_390 (O_390,N_14939,N_14838);
xnor UO_391 (O_391,N_14840,N_14552);
or UO_392 (O_392,N_14924,N_14633);
xor UO_393 (O_393,N_14951,N_14409);
or UO_394 (O_394,N_14893,N_14694);
and UO_395 (O_395,N_14600,N_14682);
and UO_396 (O_396,N_14961,N_14583);
or UO_397 (O_397,N_14762,N_14648);
and UO_398 (O_398,N_14311,N_14775);
xor UO_399 (O_399,N_14780,N_14515);
nand UO_400 (O_400,N_14273,N_14363);
and UO_401 (O_401,N_14623,N_14678);
nor UO_402 (O_402,N_14936,N_14303);
nand UO_403 (O_403,N_14597,N_14473);
xnor UO_404 (O_404,N_14470,N_14545);
or UO_405 (O_405,N_14729,N_14465);
or UO_406 (O_406,N_14342,N_14397);
nand UO_407 (O_407,N_14291,N_14497);
xor UO_408 (O_408,N_14525,N_14943);
nor UO_409 (O_409,N_14374,N_14568);
or UO_410 (O_410,N_14630,N_14390);
and UO_411 (O_411,N_14413,N_14758);
and UO_412 (O_412,N_14487,N_14357);
or UO_413 (O_413,N_14482,N_14561);
or UO_414 (O_414,N_14389,N_14837);
nor UO_415 (O_415,N_14912,N_14277);
and UO_416 (O_416,N_14304,N_14855);
or UO_417 (O_417,N_14309,N_14679);
nor UO_418 (O_418,N_14977,N_14599);
nor UO_419 (O_419,N_14313,N_14620);
and UO_420 (O_420,N_14534,N_14954);
nand UO_421 (O_421,N_14277,N_14820);
xnor UO_422 (O_422,N_14393,N_14611);
nor UO_423 (O_423,N_14838,N_14541);
nand UO_424 (O_424,N_14795,N_14529);
or UO_425 (O_425,N_14725,N_14644);
and UO_426 (O_426,N_14670,N_14303);
xnor UO_427 (O_427,N_14682,N_14996);
xor UO_428 (O_428,N_14306,N_14548);
nor UO_429 (O_429,N_14333,N_14274);
and UO_430 (O_430,N_14315,N_14601);
xnor UO_431 (O_431,N_14890,N_14898);
or UO_432 (O_432,N_14373,N_14335);
or UO_433 (O_433,N_14502,N_14910);
nor UO_434 (O_434,N_14299,N_14602);
nor UO_435 (O_435,N_14680,N_14446);
nand UO_436 (O_436,N_14413,N_14781);
xor UO_437 (O_437,N_14548,N_14403);
or UO_438 (O_438,N_14872,N_14656);
and UO_439 (O_439,N_14283,N_14874);
xor UO_440 (O_440,N_14744,N_14773);
nand UO_441 (O_441,N_14598,N_14919);
nor UO_442 (O_442,N_14653,N_14735);
xnor UO_443 (O_443,N_14735,N_14611);
nor UO_444 (O_444,N_14426,N_14896);
or UO_445 (O_445,N_14992,N_14261);
nor UO_446 (O_446,N_14343,N_14591);
nand UO_447 (O_447,N_14671,N_14318);
nor UO_448 (O_448,N_14944,N_14725);
and UO_449 (O_449,N_14616,N_14997);
and UO_450 (O_450,N_14841,N_14739);
or UO_451 (O_451,N_14708,N_14432);
or UO_452 (O_452,N_14278,N_14806);
xor UO_453 (O_453,N_14698,N_14669);
nor UO_454 (O_454,N_14804,N_14768);
nor UO_455 (O_455,N_14273,N_14671);
xnor UO_456 (O_456,N_14425,N_14786);
xor UO_457 (O_457,N_14326,N_14504);
xnor UO_458 (O_458,N_14696,N_14310);
nor UO_459 (O_459,N_14288,N_14254);
or UO_460 (O_460,N_14974,N_14692);
and UO_461 (O_461,N_14896,N_14861);
nand UO_462 (O_462,N_14290,N_14372);
nor UO_463 (O_463,N_14337,N_14858);
nand UO_464 (O_464,N_14817,N_14273);
xor UO_465 (O_465,N_14585,N_14898);
nor UO_466 (O_466,N_14715,N_14563);
nand UO_467 (O_467,N_14917,N_14280);
nand UO_468 (O_468,N_14493,N_14794);
and UO_469 (O_469,N_14348,N_14979);
xnor UO_470 (O_470,N_14348,N_14592);
nor UO_471 (O_471,N_14269,N_14661);
xnor UO_472 (O_472,N_14822,N_14717);
or UO_473 (O_473,N_14315,N_14942);
nor UO_474 (O_474,N_14745,N_14473);
or UO_475 (O_475,N_14756,N_14711);
and UO_476 (O_476,N_14445,N_14366);
nand UO_477 (O_477,N_14489,N_14461);
nand UO_478 (O_478,N_14516,N_14527);
and UO_479 (O_479,N_14925,N_14461);
nand UO_480 (O_480,N_14552,N_14461);
nand UO_481 (O_481,N_14977,N_14764);
xnor UO_482 (O_482,N_14834,N_14820);
or UO_483 (O_483,N_14908,N_14404);
and UO_484 (O_484,N_14871,N_14777);
xor UO_485 (O_485,N_14798,N_14878);
nand UO_486 (O_486,N_14542,N_14812);
xnor UO_487 (O_487,N_14697,N_14527);
nand UO_488 (O_488,N_14677,N_14744);
or UO_489 (O_489,N_14634,N_14652);
and UO_490 (O_490,N_14851,N_14505);
nor UO_491 (O_491,N_14513,N_14439);
and UO_492 (O_492,N_14563,N_14607);
xnor UO_493 (O_493,N_14947,N_14993);
or UO_494 (O_494,N_14733,N_14426);
xor UO_495 (O_495,N_14284,N_14711);
or UO_496 (O_496,N_14861,N_14357);
and UO_497 (O_497,N_14797,N_14974);
or UO_498 (O_498,N_14965,N_14691);
or UO_499 (O_499,N_14875,N_14426);
xor UO_500 (O_500,N_14259,N_14451);
nor UO_501 (O_501,N_14783,N_14326);
nor UO_502 (O_502,N_14276,N_14882);
and UO_503 (O_503,N_14296,N_14732);
xnor UO_504 (O_504,N_14992,N_14726);
and UO_505 (O_505,N_14591,N_14564);
and UO_506 (O_506,N_14805,N_14735);
or UO_507 (O_507,N_14496,N_14306);
or UO_508 (O_508,N_14266,N_14350);
or UO_509 (O_509,N_14624,N_14496);
and UO_510 (O_510,N_14401,N_14251);
nand UO_511 (O_511,N_14966,N_14403);
or UO_512 (O_512,N_14530,N_14599);
xnor UO_513 (O_513,N_14407,N_14349);
nand UO_514 (O_514,N_14722,N_14439);
and UO_515 (O_515,N_14640,N_14698);
nor UO_516 (O_516,N_14850,N_14795);
nor UO_517 (O_517,N_14772,N_14380);
xnor UO_518 (O_518,N_14774,N_14612);
xor UO_519 (O_519,N_14410,N_14640);
xnor UO_520 (O_520,N_14899,N_14585);
or UO_521 (O_521,N_14675,N_14597);
nand UO_522 (O_522,N_14848,N_14700);
nand UO_523 (O_523,N_14465,N_14847);
xnor UO_524 (O_524,N_14959,N_14489);
nor UO_525 (O_525,N_14704,N_14639);
nand UO_526 (O_526,N_14808,N_14475);
and UO_527 (O_527,N_14266,N_14803);
nand UO_528 (O_528,N_14939,N_14929);
nor UO_529 (O_529,N_14553,N_14497);
or UO_530 (O_530,N_14861,N_14886);
nand UO_531 (O_531,N_14724,N_14790);
and UO_532 (O_532,N_14916,N_14410);
and UO_533 (O_533,N_14456,N_14887);
xnor UO_534 (O_534,N_14874,N_14931);
and UO_535 (O_535,N_14923,N_14540);
nand UO_536 (O_536,N_14764,N_14941);
or UO_537 (O_537,N_14647,N_14801);
or UO_538 (O_538,N_14808,N_14801);
nand UO_539 (O_539,N_14877,N_14671);
and UO_540 (O_540,N_14989,N_14619);
nor UO_541 (O_541,N_14287,N_14394);
or UO_542 (O_542,N_14808,N_14387);
nand UO_543 (O_543,N_14869,N_14397);
nor UO_544 (O_544,N_14905,N_14330);
and UO_545 (O_545,N_14261,N_14542);
xor UO_546 (O_546,N_14687,N_14255);
and UO_547 (O_547,N_14945,N_14972);
xor UO_548 (O_548,N_14575,N_14861);
and UO_549 (O_549,N_14719,N_14450);
nand UO_550 (O_550,N_14287,N_14653);
and UO_551 (O_551,N_14941,N_14406);
or UO_552 (O_552,N_14465,N_14693);
or UO_553 (O_553,N_14371,N_14587);
xnor UO_554 (O_554,N_14810,N_14901);
nor UO_555 (O_555,N_14772,N_14465);
or UO_556 (O_556,N_14928,N_14620);
xor UO_557 (O_557,N_14687,N_14533);
and UO_558 (O_558,N_14832,N_14763);
nor UO_559 (O_559,N_14256,N_14250);
and UO_560 (O_560,N_14699,N_14867);
xnor UO_561 (O_561,N_14767,N_14897);
or UO_562 (O_562,N_14905,N_14397);
nor UO_563 (O_563,N_14775,N_14729);
or UO_564 (O_564,N_14809,N_14538);
nor UO_565 (O_565,N_14522,N_14809);
and UO_566 (O_566,N_14751,N_14490);
or UO_567 (O_567,N_14711,N_14622);
xor UO_568 (O_568,N_14428,N_14515);
nand UO_569 (O_569,N_14735,N_14498);
or UO_570 (O_570,N_14839,N_14470);
nor UO_571 (O_571,N_14994,N_14644);
nor UO_572 (O_572,N_14509,N_14330);
nor UO_573 (O_573,N_14534,N_14730);
nor UO_574 (O_574,N_14781,N_14617);
nand UO_575 (O_575,N_14675,N_14961);
nand UO_576 (O_576,N_14838,N_14264);
and UO_577 (O_577,N_14731,N_14721);
nand UO_578 (O_578,N_14754,N_14354);
nor UO_579 (O_579,N_14763,N_14379);
nor UO_580 (O_580,N_14260,N_14964);
nand UO_581 (O_581,N_14995,N_14719);
nor UO_582 (O_582,N_14511,N_14668);
and UO_583 (O_583,N_14607,N_14847);
nand UO_584 (O_584,N_14676,N_14627);
xor UO_585 (O_585,N_14938,N_14365);
nor UO_586 (O_586,N_14828,N_14389);
nor UO_587 (O_587,N_14657,N_14857);
nand UO_588 (O_588,N_14383,N_14929);
xnor UO_589 (O_589,N_14364,N_14419);
or UO_590 (O_590,N_14753,N_14342);
nand UO_591 (O_591,N_14605,N_14488);
nor UO_592 (O_592,N_14587,N_14770);
nand UO_593 (O_593,N_14913,N_14986);
and UO_594 (O_594,N_14531,N_14726);
and UO_595 (O_595,N_14852,N_14630);
nand UO_596 (O_596,N_14554,N_14962);
xnor UO_597 (O_597,N_14404,N_14613);
or UO_598 (O_598,N_14697,N_14673);
or UO_599 (O_599,N_14315,N_14608);
nand UO_600 (O_600,N_14772,N_14722);
xor UO_601 (O_601,N_14705,N_14655);
nand UO_602 (O_602,N_14781,N_14508);
and UO_603 (O_603,N_14320,N_14406);
or UO_604 (O_604,N_14583,N_14462);
or UO_605 (O_605,N_14432,N_14636);
nor UO_606 (O_606,N_14951,N_14518);
and UO_607 (O_607,N_14719,N_14449);
and UO_608 (O_608,N_14924,N_14359);
and UO_609 (O_609,N_14802,N_14976);
and UO_610 (O_610,N_14483,N_14304);
nand UO_611 (O_611,N_14838,N_14937);
nor UO_612 (O_612,N_14447,N_14897);
and UO_613 (O_613,N_14876,N_14859);
xnor UO_614 (O_614,N_14581,N_14678);
or UO_615 (O_615,N_14998,N_14814);
or UO_616 (O_616,N_14836,N_14682);
and UO_617 (O_617,N_14855,N_14825);
and UO_618 (O_618,N_14301,N_14787);
nor UO_619 (O_619,N_14251,N_14264);
nand UO_620 (O_620,N_14460,N_14696);
and UO_621 (O_621,N_14593,N_14849);
nand UO_622 (O_622,N_14362,N_14462);
nor UO_623 (O_623,N_14819,N_14984);
or UO_624 (O_624,N_14274,N_14956);
nand UO_625 (O_625,N_14920,N_14370);
nor UO_626 (O_626,N_14363,N_14269);
nand UO_627 (O_627,N_14412,N_14834);
nor UO_628 (O_628,N_14407,N_14709);
xnor UO_629 (O_629,N_14278,N_14955);
xnor UO_630 (O_630,N_14294,N_14735);
and UO_631 (O_631,N_14687,N_14423);
and UO_632 (O_632,N_14352,N_14472);
or UO_633 (O_633,N_14257,N_14616);
or UO_634 (O_634,N_14771,N_14749);
nor UO_635 (O_635,N_14862,N_14555);
and UO_636 (O_636,N_14419,N_14340);
nor UO_637 (O_637,N_14832,N_14830);
nand UO_638 (O_638,N_14320,N_14413);
nand UO_639 (O_639,N_14308,N_14749);
and UO_640 (O_640,N_14632,N_14983);
xnor UO_641 (O_641,N_14730,N_14806);
and UO_642 (O_642,N_14616,N_14642);
nand UO_643 (O_643,N_14626,N_14920);
nor UO_644 (O_644,N_14839,N_14584);
xor UO_645 (O_645,N_14477,N_14876);
or UO_646 (O_646,N_14366,N_14473);
and UO_647 (O_647,N_14348,N_14574);
or UO_648 (O_648,N_14571,N_14747);
nor UO_649 (O_649,N_14357,N_14543);
nor UO_650 (O_650,N_14533,N_14301);
xnor UO_651 (O_651,N_14846,N_14312);
xor UO_652 (O_652,N_14985,N_14573);
nor UO_653 (O_653,N_14892,N_14870);
xor UO_654 (O_654,N_14318,N_14578);
nor UO_655 (O_655,N_14776,N_14252);
and UO_656 (O_656,N_14364,N_14627);
xnor UO_657 (O_657,N_14793,N_14869);
or UO_658 (O_658,N_14538,N_14701);
nor UO_659 (O_659,N_14499,N_14342);
or UO_660 (O_660,N_14310,N_14322);
nand UO_661 (O_661,N_14629,N_14361);
and UO_662 (O_662,N_14958,N_14822);
nor UO_663 (O_663,N_14296,N_14382);
and UO_664 (O_664,N_14965,N_14921);
nor UO_665 (O_665,N_14440,N_14411);
xor UO_666 (O_666,N_14460,N_14392);
nand UO_667 (O_667,N_14977,N_14605);
and UO_668 (O_668,N_14432,N_14544);
xnor UO_669 (O_669,N_14512,N_14951);
nand UO_670 (O_670,N_14538,N_14668);
xnor UO_671 (O_671,N_14697,N_14851);
nor UO_672 (O_672,N_14283,N_14473);
or UO_673 (O_673,N_14991,N_14845);
nand UO_674 (O_674,N_14516,N_14605);
nand UO_675 (O_675,N_14378,N_14807);
or UO_676 (O_676,N_14609,N_14252);
nand UO_677 (O_677,N_14962,N_14886);
or UO_678 (O_678,N_14345,N_14333);
and UO_679 (O_679,N_14255,N_14830);
and UO_680 (O_680,N_14499,N_14604);
nor UO_681 (O_681,N_14559,N_14384);
or UO_682 (O_682,N_14891,N_14383);
nor UO_683 (O_683,N_14518,N_14603);
nor UO_684 (O_684,N_14539,N_14522);
xor UO_685 (O_685,N_14320,N_14297);
or UO_686 (O_686,N_14484,N_14991);
or UO_687 (O_687,N_14837,N_14346);
xnor UO_688 (O_688,N_14809,N_14897);
xor UO_689 (O_689,N_14469,N_14969);
and UO_690 (O_690,N_14745,N_14577);
xor UO_691 (O_691,N_14607,N_14562);
and UO_692 (O_692,N_14404,N_14468);
or UO_693 (O_693,N_14842,N_14464);
nor UO_694 (O_694,N_14586,N_14892);
xnor UO_695 (O_695,N_14699,N_14532);
nor UO_696 (O_696,N_14276,N_14345);
and UO_697 (O_697,N_14583,N_14356);
nand UO_698 (O_698,N_14993,N_14410);
nor UO_699 (O_699,N_14692,N_14825);
and UO_700 (O_700,N_14382,N_14819);
and UO_701 (O_701,N_14972,N_14279);
nor UO_702 (O_702,N_14753,N_14803);
xor UO_703 (O_703,N_14731,N_14669);
or UO_704 (O_704,N_14963,N_14968);
or UO_705 (O_705,N_14268,N_14462);
or UO_706 (O_706,N_14620,N_14828);
and UO_707 (O_707,N_14861,N_14900);
nand UO_708 (O_708,N_14613,N_14846);
xnor UO_709 (O_709,N_14337,N_14853);
or UO_710 (O_710,N_14558,N_14259);
nand UO_711 (O_711,N_14681,N_14471);
nand UO_712 (O_712,N_14910,N_14329);
or UO_713 (O_713,N_14869,N_14944);
xor UO_714 (O_714,N_14825,N_14571);
or UO_715 (O_715,N_14380,N_14575);
xor UO_716 (O_716,N_14792,N_14274);
nor UO_717 (O_717,N_14355,N_14750);
xor UO_718 (O_718,N_14687,N_14765);
nand UO_719 (O_719,N_14387,N_14544);
or UO_720 (O_720,N_14291,N_14603);
nor UO_721 (O_721,N_14337,N_14353);
and UO_722 (O_722,N_14557,N_14672);
xnor UO_723 (O_723,N_14359,N_14840);
or UO_724 (O_724,N_14825,N_14734);
nor UO_725 (O_725,N_14369,N_14952);
nor UO_726 (O_726,N_14376,N_14320);
nand UO_727 (O_727,N_14940,N_14930);
or UO_728 (O_728,N_14531,N_14891);
and UO_729 (O_729,N_14953,N_14519);
nor UO_730 (O_730,N_14743,N_14807);
or UO_731 (O_731,N_14400,N_14958);
nand UO_732 (O_732,N_14882,N_14925);
nand UO_733 (O_733,N_14889,N_14910);
nand UO_734 (O_734,N_14551,N_14366);
nor UO_735 (O_735,N_14357,N_14757);
nand UO_736 (O_736,N_14695,N_14796);
and UO_737 (O_737,N_14710,N_14725);
xnor UO_738 (O_738,N_14771,N_14862);
nand UO_739 (O_739,N_14340,N_14709);
nand UO_740 (O_740,N_14636,N_14670);
or UO_741 (O_741,N_14343,N_14725);
or UO_742 (O_742,N_14956,N_14419);
nand UO_743 (O_743,N_14876,N_14693);
nor UO_744 (O_744,N_14929,N_14841);
or UO_745 (O_745,N_14791,N_14624);
nand UO_746 (O_746,N_14305,N_14990);
xnor UO_747 (O_747,N_14753,N_14390);
nand UO_748 (O_748,N_14534,N_14547);
or UO_749 (O_749,N_14706,N_14924);
and UO_750 (O_750,N_14440,N_14592);
xnor UO_751 (O_751,N_14981,N_14305);
xor UO_752 (O_752,N_14437,N_14410);
and UO_753 (O_753,N_14328,N_14516);
nand UO_754 (O_754,N_14387,N_14899);
or UO_755 (O_755,N_14346,N_14527);
or UO_756 (O_756,N_14889,N_14815);
xor UO_757 (O_757,N_14828,N_14973);
nand UO_758 (O_758,N_14551,N_14593);
nor UO_759 (O_759,N_14563,N_14874);
nor UO_760 (O_760,N_14470,N_14342);
xnor UO_761 (O_761,N_14522,N_14698);
and UO_762 (O_762,N_14590,N_14775);
and UO_763 (O_763,N_14935,N_14892);
nor UO_764 (O_764,N_14777,N_14766);
nor UO_765 (O_765,N_14481,N_14724);
and UO_766 (O_766,N_14860,N_14313);
nor UO_767 (O_767,N_14830,N_14593);
and UO_768 (O_768,N_14801,N_14907);
nand UO_769 (O_769,N_14363,N_14873);
xor UO_770 (O_770,N_14529,N_14584);
nor UO_771 (O_771,N_14735,N_14821);
or UO_772 (O_772,N_14402,N_14264);
or UO_773 (O_773,N_14894,N_14552);
nand UO_774 (O_774,N_14608,N_14914);
nand UO_775 (O_775,N_14730,N_14284);
xnor UO_776 (O_776,N_14436,N_14499);
or UO_777 (O_777,N_14682,N_14790);
or UO_778 (O_778,N_14597,N_14708);
nand UO_779 (O_779,N_14706,N_14775);
nand UO_780 (O_780,N_14731,N_14930);
or UO_781 (O_781,N_14496,N_14331);
nand UO_782 (O_782,N_14472,N_14421);
and UO_783 (O_783,N_14936,N_14446);
nor UO_784 (O_784,N_14706,N_14728);
nor UO_785 (O_785,N_14403,N_14587);
or UO_786 (O_786,N_14280,N_14974);
nand UO_787 (O_787,N_14575,N_14333);
nor UO_788 (O_788,N_14691,N_14280);
nor UO_789 (O_789,N_14362,N_14563);
and UO_790 (O_790,N_14927,N_14672);
nand UO_791 (O_791,N_14526,N_14866);
nor UO_792 (O_792,N_14691,N_14573);
xor UO_793 (O_793,N_14280,N_14706);
or UO_794 (O_794,N_14663,N_14750);
xor UO_795 (O_795,N_14314,N_14844);
nand UO_796 (O_796,N_14338,N_14494);
nand UO_797 (O_797,N_14485,N_14991);
nand UO_798 (O_798,N_14807,N_14791);
nor UO_799 (O_799,N_14460,N_14778);
nand UO_800 (O_800,N_14526,N_14371);
xor UO_801 (O_801,N_14575,N_14902);
and UO_802 (O_802,N_14345,N_14905);
xnor UO_803 (O_803,N_14696,N_14716);
nand UO_804 (O_804,N_14546,N_14532);
nor UO_805 (O_805,N_14360,N_14715);
nand UO_806 (O_806,N_14329,N_14644);
and UO_807 (O_807,N_14383,N_14397);
or UO_808 (O_808,N_14875,N_14517);
xor UO_809 (O_809,N_14393,N_14432);
xnor UO_810 (O_810,N_14613,N_14673);
nor UO_811 (O_811,N_14644,N_14566);
nor UO_812 (O_812,N_14608,N_14296);
or UO_813 (O_813,N_14696,N_14869);
xnor UO_814 (O_814,N_14357,N_14375);
nand UO_815 (O_815,N_14329,N_14404);
nand UO_816 (O_816,N_14278,N_14420);
nand UO_817 (O_817,N_14416,N_14794);
or UO_818 (O_818,N_14259,N_14416);
and UO_819 (O_819,N_14948,N_14319);
nor UO_820 (O_820,N_14484,N_14799);
and UO_821 (O_821,N_14924,N_14414);
and UO_822 (O_822,N_14465,N_14959);
or UO_823 (O_823,N_14952,N_14801);
xnor UO_824 (O_824,N_14528,N_14465);
nand UO_825 (O_825,N_14468,N_14303);
nand UO_826 (O_826,N_14618,N_14685);
xnor UO_827 (O_827,N_14590,N_14790);
and UO_828 (O_828,N_14265,N_14833);
or UO_829 (O_829,N_14947,N_14450);
nand UO_830 (O_830,N_14477,N_14274);
nand UO_831 (O_831,N_14509,N_14976);
nor UO_832 (O_832,N_14550,N_14367);
xor UO_833 (O_833,N_14559,N_14634);
nor UO_834 (O_834,N_14619,N_14474);
nor UO_835 (O_835,N_14981,N_14277);
xor UO_836 (O_836,N_14688,N_14682);
or UO_837 (O_837,N_14284,N_14928);
nor UO_838 (O_838,N_14444,N_14251);
nand UO_839 (O_839,N_14405,N_14655);
nand UO_840 (O_840,N_14869,N_14610);
or UO_841 (O_841,N_14623,N_14738);
or UO_842 (O_842,N_14666,N_14557);
nor UO_843 (O_843,N_14368,N_14518);
and UO_844 (O_844,N_14499,N_14435);
and UO_845 (O_845,N_14649,N_14960);
xor UO_846 (O_846,N_14319,N_14437);
nor UO_847 (O_847,N_14390,N_14750);
xnor UO_848 (O_848,N_14660,N_14362);
xor UO_849 (O_849,N_14918,N_14854);
xor UO_850 (O_850,N_14708,N_14543);
xor UO_851 (O_851,N_14595,N_14846);
xor UO_852 (O_852,N_14790,N_14482);
nor UO_853 (O_853,N_14810,N_14705);
nor UO_854 (O_854,N_14567,N_14846);
and UO_855 (O_855,N_14960,N_14637);
and UO_856 (O_856,N_14899,N_14314);
and UO_857 (O_857,N_14627,N_14256);
or UO_858 (O_858,N_14509,N_14759);
or UO_859 (O_859,N_14494,N_14465);
nor UO_860 (O_860,N_14847,N_14548);
xor UO_861 (O_861,N_14746,N_14825);
nand UO_862 (O_862,N_14690,N_14979);
nor UO_863 (O_863,N_14859,N_14591);
xnor UO_864 (O_864,N_14881,N_14503);
or UO_865 (O_865,N_14450,N_14882);
nand UO_866 (O_866,N_14859,N_14585);
xnor UO_867 (O_867,N_14926,N_14655);
nand UO_868 (O_868,N_14923,N_14777);
or UO_869 (O_869,N_14564,N_14952);
xor UO_870 (O_870,N_14681,N_14884);
or UO_871 (O_871,N_14804,N_14741);
or UO_872 (O_872,N_14444,N_14265);
nand UO_873 (O_873,N_14771,N_14511);
and UO_874 (O_874,N_14865,N_14856);
xor UO_875 (O_875,N_14570,N_14258);
and UO_876 (O_876,N_14341,N_14923);
nand UO_877 (O_877,N_14943,N_14393);
nand UO_878 (O_878,N_14310,N_14727);
or UO_879 (O_879,N_14577,N_14925);
or UO_880 (O_880,N_14928,N_14960);
nand UO_881 (O_881,N_14664,N_14350);
and UO_882 (O_882,N_14522,N_14844);
xnor UO_883 (O_883,N_14649,N_14300);
or UO_884 (O_884,N_14758,N_14841);
nor UO_885 (O_885,N_14353,N_14361);
and UO_886 (O_886,N_14330,N_14987);
and UO_887 (O_887,N_14930,N_14888);
nor UO_888 (O_888,N_14308,N_14700);
xnor UO_889 (O_889,N_14945,N_14799);
and UO_890 (O_890,N_14482,N_14448);
and UO_891 (O_891,N_14401,N_14440);
xor UO_892 (O_892,N_14658,N_14716);
and UO_893 (O_893,N_14489,N_14523);
xnor UO_894 (O_894,N_14452,N_14696);
nand UO_895 (O_895,N_14616,N_14312);
nor UO_896 (O_896,N_14805,N_14957);
nor UO_897 (O_897,N_14615,N_14737);
xor UO_898 (O_898,N_14464,N_14866);
and UO_899 (O_899,N_14978,N_14359);
and UO_900 (O_900,N_14905,N_14608);
nand UO_901 (O_901,N_14486,N_14862);
nor UO_902 (O_902,N_14768,N_14962);
nor UO_903 (O_903,N_14312,N_14567);
or UO_904 (O_904,N_14535,N_14828);
or UO_905 (O_905,N_14388,N_14503);
xor UO_906 (O_906,N_14729,N_14457);
nor UO_907 (O_907,N_14296,N_14357);
and UO_908 (O_908,N_14893,N_14821);
and UO_909 (O_909,N_14713,N_14558);
xor UO_910 (O_910,N_14545,N_14874);
nor UO_911 (O_911,N_14442,N_14700);
nand UO_912 (O_912,N_14399,N_14640);
xor UO_913 (O_913,N_14566,N_14432);
and UO_914 (O_914,N_14437,N_14714);
or UO_915 (O_915,N_14791,N_14627);
nand UO_916 (O_916,N_14281,N_14678);
or UO_917 (O_917,N_14723,N_14518);
and UO_918 (O_918,N_14407,N_14431);
and UO_919 (O_919,N_14323,N_14714);
nor UO_920 (O_920,N_14264,N_14471);
nand UO_921 (O_921,N_14901,N_14697);
nand UO_922 (O_922,N_14335,N_14898);
and UO_923 (O_923,N_14903,N_14939);
nor UO_924 (O_924,N_14505,N_14840);
xor UO_925 (O_925,N_14758,N_14921);
nor UO_926 (O_926,N_14412,N_14288);
xnor UO_927 (O_927,N_14346,N_14791);
nand UO_928 (O_928,N_14917,N_14969);
xnor UO_929 (O_929,N_14932,N_14660);
nand UO_930 (O_930,N_14660,N_14376);
xor UO_931 (O_931,N_14374,N_14415);
xnor UO_932 (O_932,N_14443,N_14740);
xor UO_933 (O_933,N_14554,N_14866);
nand UO_934 (O_934,N_14868,N_14347);
nand UO_935 (O_935,N_14954,N_14467);
nor UO_936 (O_936,N_14708,N_14904);
xor UO_937 (O_937,N_14345,N_14290);
and UO_938 (O_938,N_14752,N_14789);
and UO_939 (O_939,N_14577,N_14250);
nor UO_940 (O_940,N_14592,N_14584);
and UO_941 (O_941,N_14330,N_14941);
xnor UO_942 (O_942,N_14439,N_14980);
xor UO_943 (O_943,N_14919,N_14353);
or UO_944 (O_944,N_14724,N_14456);
nor UO_945 (O_945,N_14889,N_14349);
or UO_946 (O_946,N_14664,N_14970);
xnor UO_947 (O_947,N_14636,N_14714);
nand UO_948 (O_948,N_14708,N_14684);
nand UO_949 (O_949,N_14363,N_14348);
nand UO_950 (O_950,N_14903,N_14516);
and UO_951 (O_951,N_14641,N_14711);
nor UO_952 (O_952,N_14949,N_14264);
nand UO_953 (O_953,N_14339,N_14638);
xor UO_954 (O_954,N_14533,N_14909);
nand UO_955 (O_955,N_14964,N_14746);
nor UO_956 (O_956,N_14870,N_14310);
nor UO_957 (O_957,N_14826,N_14621);
xor UO_958 (O_958,N_14701,N_14469);
and UO_959 (O_959,N_14354,N_14568);
nand UO_960 (O_960,N_14931,N_14644);
xnor UO_961 (O_961,N_14691,N_14576);
nor UO_962 (O_962,N_14406,N_14689);
or UO_963 (O_963,N_14790,N_14349);
or UO_964 (O_964,N_14940,N_14956);
or UO_965 (O_965,N_14608,N_14916);
and UO_966 (O_966,N_14647,N_14351);
nor UO_967 (O_967,N_14296,N_14774);
nand UO_968 (O_968,N_14640,N_14300);
or UO_969 (O_969,N_14979,N_14989);
xor UO_970 (O_970,N_14951,N_14515);
nor UO_971 (O_971,N_14624,N_14979);
or UO_972 (O_972,N_14886,N_14534);
xor UO_973 (O_973,N_14750,N_14308);
nand UO_974 (O_974,N_14523,N_14922);
nand UO_975 (O_975,N_14483,N_14509);
nand UO_976 (O_976,N_14519,N_14499);
nand UO_977 (O_977,N_14659,N_14914);
and UO_978 (O_978,N_14732,N_14852);
nor UO_979 (O_979,N_14908,N_14640);
and UO_980 (O_980,N_14385,N_14802);
nand UO_981 (O_981,N_14863,N_14364);
nand UO_982 (O_982,N_14584,N_14688);
nand UO_983 (O_983,N_14447,N_14873);
or UO_984 (O_984,N_14859,N_14673);
xor UO_985 (O_985,N_14433,N_14403);
and UO_986 (O_986,N_14850,N_14496);
and UO_987 (O_987,N_14745,N_14676);
nor UO_988 (O_988,N_14346,N_14762);
xnor UO_989 (O_989,N_14371,N_14728);
xnor UO_990 (O_990,N_14413,N_14963);
nand UO_991 (O_991,N_14715,N_14543);
and UO_992 (O_992,N_14541,N_14250);
xor UO_993 (O_993,N_14716,N_14887);
or UO_994 (O_994,N_14364,N_14429);
nor UO_995 (O_995,N_14511,N_14314);
and UO_996 (O_996,N_14640,N_14329);
nor UO_997 (O_997,N_14774,N_14520);
nand UO_998 (O_998,N_14398,N_14409);
nand UO_999 (O_999,N_14989,N_14279);
xor UO_1000 (O_1000,N_14618,N_14278);
nand UO_1001 (O_1001,N_14344,N_14740);
nand UO_1002 (O_1002,N_14493,N_14674);
and UO_1003 (O_1003,N_14462,N_14910);
nand UO_1004 (O_1004,N_14804,N_14764);
nand UO_1005 (O_1005,N_14769,N_14962);
and UO_1006 (O_1006,N_14870,N_14336);
nor UO_1007 (O_1007,N_14282,N_14259);
xnor UO_1008 (O_1008,N_14818,N_14348);
nand UO_1009 (O_1009,N_14718,N_14956);
xor UO_1010 (O_1010,N_14370,N_14401);
xor UO_1011 (O_1011,N_14706,N_14739);
or UO_1012 (O_1012,N_14338,N_14791);
and UO_1013 (O_1013,N_14605,N_14403);
xor UO_1014 (O_1014,N_14718,N_14264);
nor UO_1015 (O_1015,N_14566,N_14507);
or UO_1016 (O_1016,N_14963,N_14397);
or UO_1017 (O_1017,N_14879,N_14269);
and UO_1018 (O_1018,N_14415,N_14402);
nor UO_1019 (O_1019,N_14984,N_14356);
nand UO_1020 (O_1020,N_14598,N_14448);
nand UO_1021 (O_1021,N_14957,N_14585);
nand UO_1022 (O_1022,N_14278,N_14472);
nor UO_1023 (O_1023,N_14672,N_14573);
nor UO_1024 (O_1024,N_14875,N_14397);
xnor UO_1025 (O_1025,N_14986,N_14928);
and UO_1026 (O_1026,N_14963,N_14567);
nor UO_1027 (O_1027,N_14933,N_14749);
or UO_1028 (O_1028,N_14289,N_14507);
and UO_1029 (O_1029,N_14589,N_14345);
nand UO_1030 (O_1030,N_14829,N_14909);
nand UO_1031 (O_1031,N_14374,N_14372);
nand UO_1032 (O_1032,N_14791,N_14319);
nor UO_1033 (O_1033,N_14915,N_14618);
or UO_1034 (O_1034,N_14759,N_14960);
nand UO_1035 (O_1035,N_14482,N_14731);
nand UO_1036 (O_1036,N_14625,N_14851);
xor UO_1037 (O_1037,N_14924,N_14363);
xor UO_1038 (O_1038,N_14364,N_14589);
and UO_1039 (O_1039,N_14579,N_14909);
xor UO_1040 (O_1040,N_14740,N_14801);
nor UO_1041 (O_1041,N_14887,N_14654);
and UO_1042 (O_1042,N_14744,N_14447);
xnor UO_1043 (O_1043,N_14795,N_14839);
and UO_1044 (O_1044,N_14509,N_14323);
nor UO_1045 (O_1045,N_14346,N_14906);
xnor UO_1046 (O_1046,N_14616,N_14691);
nand UO_1047 (O_1047,N_14519,N_14689);
or UO_1048 (O_1048,N_14576,N_14584);
or UO_1049 (O_1049,N_14450,N_14886);
xor UO_1050 (O_1050,N_14923,N_14489);
nor UO_1051 (O_1051,N_14893,N_14275);
nand UO_1052 (O_1052,N_14748,N_14798);
or UO_1053 (O_1053,N_14546,N_14535);
or UO_1054 (O_1054,N_14522,N_14424);
nand UO_1055 (O_1055,N_14702,N_14637);
xor UO_1056 (O_1056,N_14307,N_14730);
and UO_1057 (O_1057,N_14690,N_14298);
or UO_1058 (O_1058,N_14991,N_14445);
xor UO_1059 (O_1059,N_14928,N_14775);
or UO_1060 (O_1060,N_14959,N_14809);
and UO_1061 (O_1061,N_14993,N_14784);
or UO_1062 (O_1062,N_14334,N_14916);
or UO_1063 (O_1063,N_14313,N_14833);
nand UO_1064 (O_1064,N_14649,N_14983);
nand UO_1065 (O_1065,N_14380,N_14647);
xnor UO_1066 (O_1066,N_14621,N_14294);
nand UO_1067 (O_1067,N_14698,N_14632);
nand UO_1068 (O_1068,N_14923,N_14691);
or UO_1069 (O_1069,N_14451,N_14873);
and UO_1070 (O_1070,N_14345,N_14736);
nor UO_1071 (O_1071,N_14436,N_14774);
xnor UO_1072 (O_1072,N_14662,N_14832);
xnor UO_1073 (O_1073,N_14626,N_14256);
or UO_1074 (O_1074,N_14691,N_14466);
nand UO_1075 (O_1075,N_14542,N_14476);
and UO_1076 (O_1076,N_14907,N_14716);
nand UO_1077 (O_1077,N_14878,N_14721);
nor UO_1078 (O_1078,N_14475,N_14702);
nand UO_1079 (O_1079,N_14941,N_14961);
nand UO_1080 (O_1080,N_14359,N_14372);
and UO_1081 (O_1081,N_14823,N_14313);
xnor UO_1082 (O_1082,N_14445,N_14685);
nor UO_1083 (O_1083,N_14438,N_14831);
or UO_1084 (O_1084,N_14267,N_14986);
or UO_1085 (O_1085,N_14634,N_14565);
or UO_1086 (O_1086,N_14926,N_14935);
xnor UO_1087 (O_1087,N_14395,N_14829);
and UO_1088 (O_1088,N_14292,N_14780);
xor UO_1089 (O_1089,N_14770,N_14850);
nand UO_1090 (O_1090,N_14708,N_14943);
and UO_1091 (O_1091,N_14305,N_14489);
or UO_1092 (O_1092,N_14771,N_14585);
or UO_1093 (O_1093,N_14900,N_14937);
xnor UO_1094 (O_1094,N_14615,N_14448);
xor UO_1095 (O_1095,N_14313,N_14988);
or UO_1096 (O_1096,N_14300,N_14377);
nand UO_1097 (O_1097,N_14915,N_14334);
and UO_1098 (O_1098,N_14461,N_14366);
and UO_1099 (O_1099,N_14516,N_14488);
nand UO_1100 (O_1100,N_14374,N_14637);
nor UO_1101 (O_1101,N_14913,N_14676);
nor UO_1102 (O_1102,N_14762,N_14362);
or UO_1103 (O_1103,N_14544,N_14996);
nand UO_1104 (O_1104,N_14395,N_14777);
nand UO_1105 (O_1105,N_14524,N_14926);
nand UO_1106 (O_1106,N_14567,N_14655);
xor UO_1107 (O_1107,N_14683,N_14948);
xnor UO_1108 (O_1108,N_14610,N_14794);
or UO_1109 (O_1109,N_14351,N_14774);
and UO_1110 (O_1110,N_14675,N_14339);
nand UO_1111 (O_1111,N_14625,N_14446);
xor UO_1112 (O_1112,N_14251,N_14273);
and UO_1113 (O_1113,N_14958,N_14810);
and UO_1114 (O_1114,N_14637,N_14316);
nor UO_1115 (O_1115,N_14338,N_14414);
nor UO_1116 (O_1116,N_14592,N_14947);
and UO_1117 (O_1117,N_14953,N_14313);
nor UO_1118 (O_1118,N_14427,N_14489);
or UO_1119 (O_1119,N_14359,N_14755);
and UO_1120 (O_1120,N_14997,N_14306);
or UO_1121 (O_1121,N_14666,N_14416);
and UO_1122 (O_1122,N_14497,N_14762);
xor UO_1123 (O_1123,N_14845,N_14407);
or UO_1124 (O_1124,N_14471,N_14437);
nor UO_1125 (O_1125,N_14920,N_14336);
nand UO_1126 (O_1126,N_14587,N_14970);
nor UO_1127 (O_1127,N_14384,N_14751);
or UO_1128 (O_1128,N_14605,N_14941);
and UO_1129 (O_1129,N_14476,N_14486);
xnor UO_1130 (O_1130,N_14604,N_14501);
nand UO_1131 (O_1131,N_14646,N_14588);
nor UO_1132 (O_1132,N_14944,N_14953);
nor UO_1133 (O_1133,N_14315,N_14475);
or UO_1134 (O_1134,N_14993,N_14449);
xor UO_1135 (O_1135,N_14943,N_14346);
or UO_1136 (O_1136,N_14601,N_14856);
nand UO_1137 (O_1137,N_14987,N_14606);
or UO_1138 (O_1138,N_14622,N_14916);
and UO_1139 (O_1139,N_14295,N_14909);
and UO_1140 (O_1140,N_14406,N_14730);
and UO_1141 (O_1141,N_14382,N_14414);
xor UO_1142 (O_1142,N_14616,N_14621);
and UO_1143 (O_1143,N_14979,N_14263);
nor UO_1144 (O_1144,N_14981,N_14752);
xor UO_1145 (O_1145,N_14651,N_14772);
and UO_1146 (O_1146,N_14691,N_14333);
and UO_1147 (O_1147,N_14517,N_14271);
or UO_1148 (O_1148,N_14520,N_14625);
nand UO_1149 (O_1149,N_14934,N_14854);
nor UO_1150 (O_1150,N_14345,N_14539);
and UO_1151 (O_1151,N_14596,N_14917);
and UO_1152 (O_1152,N_14506,N_14451);
and UO_1153 (O_1153,N_14363,N_14854);
xor UO_1154 (O_1154,N_14638,N_14509);
xor UO_1155 (O_1155,N_14924,N_14798);
and UO_1156 (O_1156,N_14774,N_14587);
or UO_1157 (O_1157,N_14509,N_14550);
xor UO_1158 (O_1158,N_14556,N_14791);
nand UO_1159 (O_1159,N_14720,N_14815);
or UO_1160 (O_1160,N_14925,N_14401);
and UO_1161 (O_1161,N_14789,N_14919);
nand UO_1162 (O_1162,N_14273,N_14452);
nor UO_1163 (O_1163,N_14351,N_14630);
nand UO_1164 (O_1164,N_14784,N_14375);
xnor UO_1165 (O_1165,N_14938,N_14649);
and UO_1166 (O_1166,N_14392,N_14940);
nor UO_1167 (O_1167,N_14680,N_14575);
nor UO_1168 (O_1168,N_14429,N_14694);
nand UO_1169 (O_1169,N_14469,N_14276);
nand UO_1170 (O_1170,N_14886,N_14486);
nor UO_1171 (O_1171,N_14964,N_14595);
xor UO_1172 (O_1172,N_14509,N_14400);
and UO_1173 (O_1173,N_14394,N_14811);
nor UO_1174 (O_1174,N_14889,N_14598);
nand UO_1175 (O_1175,N_14815,N_14596);
and UO_1176 (O_1176,N_14307,N_14480);
xnor UO_1177 (O_1177,N_14640,N_14659);
and UO_1178 (O_1178,N_14818,N_14317);
xnor UO_1179 (O_1179,N_14881,N_14410);
nor UO_1180 (O_1180,N_14552,N_14950);
and UO_1181 (O_1181,N_14905,N_14749);
nor UO_1182 (O_1182,N_14342,N_14413);
nand UO_1183 (O_1183,N_14622,N_14952);
xnor UO_1184 (O_1184,N_14581,N_14875);
and UO_1185 (O_1185,N_14973,N_14950);
and UO_1186 (O_1186,N_14820,N_14268);
xnor UO_1187 (O_1187,N_14269,N_14740);
and UO_1188 (O_1188,N_14362,N_14980);
nor UO_1189 (O_1189,N_14750,N_14678);
xor UO_1190 (O_1190,N_14968,N_14300);
and UO_1191 (O_1191,N_14280,N_14461);
or UO_1192 (O_1192,N_14480,N_14267);
or UO_1193 (O_1193,N_14274,N_14960);
nor UO_1194 (O_1194,N_14455,N_14521);
or UO_1195 (O_1195,N_14450,N_14390);
or UO_1196 (O_1196,N_14582,N_14938);
xnor UO_1197 (O_1197,N_14877,N_14635);
and UO_1198 (O_1198,N_14308,N_14622);
nand UO_1199 (O_1199,N_14765,N_14664);
nor UO_1200 (O_1200,N_14486,N_14525);
nand UO_1201 (O_1201,N_14669,N_14465);
and UO_1202 (O_1202,N_14263,N_14705);
or UO_1203 (O_1203,N_14466,N_14990);
or UO_1204 (O_1204,N_14711,N_14950);
nand UO_1205 (O_1205,N_14427,N_14719);
or UO_1206 (O_1206,N_14431,N_14587);
xor UO_1207 (O_1207,N_14525,N_14902);
or UO_1208 (O_1208,N_14917,N_14484);
and UO_1209 (O_1209,N_14567,N_14680);
nand UO_1210 (O_1210,N_14760,N_14558);
and UO_1211 (O_1211,N_14843,N_14764);
and UO_1212 (O_1212,N_14524,N_14393);
nand UO_1213 (O_1213,N_14528,N_14409);
nand UO_1214 (O_1214,N_14314,N_14631);
and UO_1215 (O_1215,N_14513,N_14878);
nor UO_1216 (O_1216,N_14752,N_14486);
nor UO_1217 (O_1217,N_14529,N_14437);
and UO_1218 (O_1218,N_14336,N_14827);
xnor UO_1219 (O_1219,N_14975,N_14704);
nor UO_1220 (O_1220,N_14900,N_14967);
nor UO_1221 (O_1221,N_14273,N_14807);
nor UO_1222 (O_1222,N_14337,N_14454);
or UO_1223 (O_1223,N_14882,N_14270);
nand UO_1224 (O_1224,N_14996,N_14618);
xor UO_1225 (O_1225,N_14914,N_14737);
or UO_1226 (O_1226,N_14849,N_14938);
nand UO_1227 (O_1227,N_14297,N_14252);
nand UO_1228 (O_1228,N_14430,N_14623);
nand UO_1229 (O_1229,N_14678,N_14967);
or UO_1230 (O_1230,N_14550,N_14505);
nand UO_1231 (O_1231,N_14327,N_14943);
xnor UO_1232 (O_1232,N_14761,N_14788);
nand UO_1233 (O_1233,N_14894,N_14256);
nand UO_1234 (O_1234,N_14814,N_14753);
nor UO_1235 (O_1235,N_14556,N_14379);
xnor UO_1236 (O_1236,N_14277,N_14725);
xor UO_1237 (O_1237,N_14939,N_14845);
xor UO_1238 (O_1238,N_14287,N_14830);
nand UO_1239 (O_1239,N_14664,N_14900);
xor UO_1240 (O_1240,N_14870,N_14533);
or UO_1241 (O_1241,N_14636,N_14967);
and UO_1242 (O_1242,N_14792,N_14265);
nand UO_1243 (O_1243,N_14564,N_14865);
or UO_1244 (O_1244,N_14587,N_14594);
nor UO_1245 (O_1245,N_14795,N_14440);
nor UO_1246 (O_1246,N_14588,N_14945);
xnor UO_1247 (O_1247,N_14868,N_14731);
xor UO_1248 (O_1248,N_14308,N_14881);
nor UO_1249 (O_1249,N_14837,N_14895);
nand UO_1250 (O_1250,N_14634,N_14304);
or UO_1251 (O_1251,N_14536,N_14997);
xor UO_1252 (O_1252,N_14274,N_14852);
or UO_1253 (O_1253,N_14592,N_14449);
nor UO_1254 (O_1254,N_14429,N_14433);
nand UO_1255 (O_1255,N_14731,N_14954);
xnor UO_1256 (O_1256,N_14942,N_14908);
nor UO_1257 (O_1257,N_14252,N_14624);
and UO_1258 (O_1258,N_14593,N_14783);
nor UO_1259 (O_1259,N_14867,N_14845);
nor UO_1260 (O_1260,N_14482,N_14768);
and UO_1261 (O_1261,N_14903,N_14712);
xnor UO_1262 (O_1262,N_14257,N_14502);
or UO_1263 (O_1263,N_14251,N_14790);
or UO_1264 (O_1264,N_14633,N_14605);
and UO_1265 (O_1265,N_14278,N_14926);
or UO_1266 (O_1266,N_14717,N_14362);
or UO_1267 (O_1267,N_14682,N_14995);
xnor UO_1268 (O_1268,N_14865,N_14531);
nand UO_1269 (O_1269,N_14716,N_14458);
xnor UO_1270 (O_1270,N_14574,N_14984);
or UO_1271 (O_1271,N_14311,N_14389);
xnor UO_1272 (O_1272,N_14360,N_14365);
or UO_1273 (O_1273,N_14448,N_14901);
or UO_1274 (O_1274,N_14481,N_14934);
or UO_1275 (O_1275,N_14826,N_14625);
and UO_1276 (O_1276,N_14757,N_14335);
nand UO_1277 (O_1277,N_14919,N_14771);
nor UO_1278 (O_1278,N_14631,N_14657);
and UO_1279 (O_1279,N_14512,N_14792);
nor UO_1280 (O_1280,N_14310,N_14700);
and UO_1281 (O_1281,N_14756,N_14456);
nand UO_1282 (O_1282,N_14501,N_14526);
and UO_1283 (O_1283,N_14520,N_14389);
and UO_1284 (O_1284,N_14512,N_14800);
and UO_1285 (O_1285,N_14845,N_14821);
or UO_1286 (O_1286,N_14345,N_14545);
or UO_1287 (O_1287,N_14550,N_14343);
nor UO_1288 (O_1288,N_14619,N_14708);
xnor UO_1289 (O_1289,N_14317,N_14730);
xor UO_1290 (O_1290,N_14424,N_14362);
and UO_1291 (O_1291,N_14897,N_14250);
or UO_1292 (O_1292,N_14498,N_14485);
nand UO_1293 (O_1293,N_14550,N_14314);
or UO_1294 (O_1294,N_14277,N_14416);
xor UO_1295 (O_1295,N_14595,N_14465);
nor UO_1296 (O_1296,N_14316,N_14879);
nor UO_1297 (O_1297,N_14932,N_14717);
and UO_1298 (O_1298,N_14275,N_14593);
nand UO_1299 (O_1299,N_14301,N_14698);
or UO_1300 (O_1300,N_14714,N_14820);
nand UO_1301 (O_1301,N_14632,N_14250);
nand UO_1302 (O_1302,N_14560,N_14343);
and UO_1303 (O_1303,N_14736,N_14529);
nor UO_1304 (O_1304,N_14269,N_14733);
nand UO_1305 (O_1305,N_14525,N_14290);
and UO_1306 (O_1306,N_14691,N_14661);
nand UO_1307 (O_1307,N_14768,N_14845);
nand UO_1308 (O_1308,N_14435,N_14475);
nand UO_1309 (O_1309,N_14349,N_14644);
or UO_1310 (O_1310,N_14383,N_14858);
xor UO_1311 (O_1311,N_14687,N_14382);
nand UO_1312 (O_1312,N_14510,N_14816);
or UO_1313 (O_1313,N_14650,N_14889);
nand UO_1314 (O_1314,N_14666,N_14931);
nor UO_1315 (O_1315,N_14693,N_14867);
and UO_1316 (O_1316,N_14930,N_14960);
nand UO_1317 (O_1317,N_14860,N_14643);
and UO_1318 (O_1318,N_14370,N_14657);
and UO_1319 (O_1319,N_14698,N_14465);
and UO_1320 (O_1320,N_14939,N_14849);
xor UO_1321 (O_1321,N_14772,N_14330);
nand UO_1322 (O_1322,N_14705,N_14524);
or UO_1323 (O_1323,N_14983,N_14630);
or UO_1324 (O_1324,N_14955,N_14292);
nand UO_1325 (O_1325,N_14362,N_14486);
nand UO_1326 (O_1326,N_14581,N_14729);
and UO_1327 (O_1327,N_14302,N_14661);
nand UO_1328 (O_1328,N_14893,N_14939);
nand UO_1329 (O_1329,N_14844,N_14850);
nor UO_1330 (O_1330,N_14607,N_14594);
xnor UO_1331 (O_1331,N_14613,N_14642);
nor UO_1332 (O_1332,N_14881,N_14550);
nand UO_1333 (O_1333,N_14899,N_14778);
nand UO_1334 (O_1334,N_14503,N_14493);
nand UO_1335 (O_1335,N_14795,N_14581);
nand UO_1336 (O_1336,N_14674,N_14555);
xor UO_1337 (O_1337,N_14948,N_14692);
nand UO_1338 (O_1338,N_14848,N_14346);
or UO_1339 (O_1339,N_14353,N_14944);
and UO_1340 (O_1340,N_14518,N_14591);
xor UO_1341 (O_1341,N_14767,N_14343);
nor UO_1342 (O_1342,N_14423,N_14536);
xnor UO_1343 (O_1343,N_14392,N_14799);
or UO_1344 (O_1344,N_14557,N_14795);
or UO_1345 (O_1345,N_14865,N_14286);
or UO_1346 (O_1346,N_14281,N_14541);
nor UO_1347 (O_1347,N_14574,N_14717);
nand UO_1348 (O_1348,N_14687,N_14700);
nand UO_1349 (O_1349,N_14387,N_14791);
and UO_1350 (O_1350,N_14513,N_14802);
or UO_1351 (O_1351,N_14507,N_14705);
and UO_1352 (O_1352,N_14318,N_14688);
nor UO_1353 (O_1353,N_14770,N_14471);
or UO_1354 (O_1354,N_14478,N_14800);
nand UO_1355 (O_1355,N_14855,N_14689);
nand UO_1356 (O_1356,N_14543,N_14525);
or UO_1357 (O_1357,N_14412,N_14610);
and UO_1358 (O_1358,N_14769,N_14541);
nor UO_1359 (O_1359,N_14681,N_14252);
xnor UO_1360 (O_1360,N_14445,N_14460);
nand UO_1361 (O_1361,N_14882,N_14382);
nor UO_1362 (O_1362,N_14437,N_14435);
or UO_1363 (O_1363,N_14416,N_14700);
nor UO_1364 (O_1364,N_14804,N_14655);
and UO_1365 (O_1365,N_14660,N_14593);
xnor UO_1366 (O_1366,N_14972,N_14803);
nor UO_1367 (O_1367,N_14718,N_14372);
xor UO_1368 (O_1368,N_14288,N_14911);
and UO_1369 (O_1369,N_14516,N_14434);
or UO_1370 (O_1370,N_14830,N_14643);
nor UO_1371 (O_1371,N_14535,N_14686);
nor UO_1372 (O_1372,N_14818,N_14862);
and UO_1373 (O_1373,N_14319,N_14392);
and UO_1374 (O_1374,N_14823,N_14606);
or UO_1375 (O_1375,N_14413,N_14816);
or UO_1376 (O_1376,N_14824,N_14386);
and UO_1377 (O_1377,N_14530,N_14652);
nand UO_1378 (O_1378,N_14530,N_14551);
and UO_1379 (O_1379,N_14976,N_14882);
xor UO_1380 (O_1380,N_14387,N_14589);
nand UO_1381 (O_1381,N_14596,N_14701);
nand UO_1382 (O_1382,N_14753,N_14813);
nand UO_1383 (O_1383,N_14424,N_14483);
xor UO_1384 (O_1384,N_14984,N_14832);
or UO_1385 (O_1385,N_14970,N_14315);
or UO_1386 (O_1386,N_14942,N_14672);
xnor UO_1387 (O_1387,N_14408,N_14713);
and UO_1388 (O_1388,N_14972,N_14614);
nand UO_1389 (O_1389,N_14389,N_14729);
nor UO_1390 (O_1390,N_14892,N_14691);
nand UO_1391 (O_1391,N_14835,N_14817);
nor UO_1392 (O_1392,N_14648,N_14514);
or UO_1393 (O_1393,N_14291,N_14932);
and UO_1394 (O_1394,N_14988,N_14526);
and UO_1395 (O_1395,N_14309,N_14705);
nor UO_1396 (O_1396,N_14679,N_14697);
nor UO_1397 (O_1397,N_14556,N_14934);
or UO_1398 (O_1398,N_14286,N_14292);
nor UO_1399 (O_1399,N_14305,N_14879);
nand UO_1400 (O_1400,N_14602,N_14701);
xnor UO_1401 (O_1401,N_14766,N_14681);
or UO_1402 (O_1402,N_14972,N_14454);
nand UO_1403 (O_1403,N_14769,N_14827);
nor UO_1404 (O_1404,N_14500,N_14832);
nand UO_1405 (O_1405,N_14906,N_14928);
nor UO_1406 (O_1406,N_14383,N_14804);
nor UO_1407 (O_1407,N_14258,N_14588);
nor UO_1408 (O_1408,N_14778,N_14672);
and UO_1409 (O_1409,N_14501,N_14483);
xnor UO_1410 (O_1410,N_14398,N_14415);
nor UO_1411 (O_1411,N_14843,N_14576);
or UO_1412 (O_1412,N_14250,N_14743);
nor UO_1413 (O_1413,N_14879,N_14662);
and UO_1414 (O_1414,N_14976,N_14313);
nor UO_1415 (O_1415,N_14621,N_14303);
xnor UO_1416 (O_1416,N_14664,N_14991);
nor UO_1417 (O_1417,N_14987,N_14336);
xnor UO_1418 (O_1418,N_14481,N_14770);
nor UO_1419 (O_1419,N_14459,N_14946);
xnor UO_1420 (O_1420,N_14928,N_14859);
nor UO_1421 (O_1421,N_14682,N_14959);
xnor UO_1422 (O_1422,N_14486,N_14677);
nor UO_1423 (O_1423,N_14259,N_14458);
nor UO_1424 (O_1424,N_14433,N_14798);
nand UO_1425 (O_1425,N_14866,N_14639);
or UO_1426 (O_1426,N_14698,N_14384);
or UO_1427 (O_1427,N_14645,N_14937);
nor UO_1428 (O_1428,N_14452,N_14893);
nor UO_1429 (O_1429,N_14391,N_14291);
xor UO_1430 (O_1430,N_14956,N_14354);
or UO_1431 (O_1431,N_14252,N_14923);
xnor UO_1432 (O_1432,N_14967,N_14584);
nor UO_1433 (O_1433,N_14919,N_14648);
or UO_1434 (O_1434,N_14722,N_14736);
or UO_1435 (O_1435,N_14702,N_14750);
and UO_1436 (O_1436,N_14656,N_14802);
and UO_1437 (O_1437,N_14329,N_14673);
nor UO_1438 (O_1438,N_14765,N_14523);
and UO_1439 (O_1439,N_14835,N_14832);
nand UO_1440 (O_1440,N_14450,N_14904);
or UO_1441 (O_1441,N_14446,N_14971);
xnor UO_1442 (O_1442,N_14496,N_14375);
xnor UO_1443 (O_1443,N_14571,N_14750);
and UO_1444 (O_1444,N_14814,N_14402);
or UO_1445 (O_1445,N_14255,N_14943);
xor UO_1446 (O_1446,N_14277,N_14882);
xnor UO_1447 (O_1447,N_14666,N_14620);
xor UO_1448 (O_1448,N_14420,N_14457);
xor UO_1449 (O_1449,N_14463,N_14704);
and UO_1450 (O_1450,N_14917,N_14792);
xnor UO_1451 (O_1451,N_14354,N_14969);
and UO_1452 (O_1452,N_14973,N_14557);
xnor UO_1453 (O_1453,N_14501,N_14945);
and UO_1454 (O_1454,N_14423,N_14510);
xor UO_1455 (O_1455,N_14594,N_14327);
nor UO_1456 (O_1456,N_14543,N_14323);
and UO_1457 (O_1457,N_14703,N_14604);
nand UO_1458 (O_1458,N_14782,N_14375);
nor UO_1459 (O_1459,N_14337,N_14385);
nor UO_1460 (O_1460,N_14566,N_14712);
nor UO_1461 (O_1461,N_14429,N_14264);
nor UO_1462 (O_1462,N_14778,N_14584);
nor UO_1463 (O_1463,N_14311,N_14404);
nor UO_1464 (O_1464,N_14334,N_14276);
nor UO_1465 (O_1465,N_14498,N_14257);
and UO_1466 (O_1466,N_14882,N_14457);
and UO_1467 (O_1467,N_14434,N_14692);
nand UO_1468 (O_1468,N_14921,N_14485);
xnor UO_1469 (O_1469,N_14515,N_14986);
nand UO_1470 (O_1470,N_14523,N_14422);
nand UO_1471 (O_1471,N_14359,N_14319);
nor UO_1472 (O_1472,N_14375,N_14562);
nor UO_1473 (O_1473,N_14277,N_14313);
xnor UO_1474 (O_1474,N_14771,N_14376);
or UO_1475 (O_1475,N_14753,N_14328);
nand UO_1476 (O_1476,N_14344,N_14737);
xor UO_1477 (O_1477,N_14398,N_14425);
nor UO_1478 (O_1478,N_14637,N_14948);
nand UO_1479 (O_1479,N_14556,N_14983);
or UO_1480 (O_1480,N_14623,N_14778);
nor UO_1481 (O_1481,N_14997,N_14825);
xor UO_1482 (O_1482,N_14382,N_14378);
nand UO_1483 (O_1483,N_14870,N_14858);
nor UO_1484 (O_1484,N_14649,N_14704);
nor UO_1485 (O_1485,N_14531,N_14961);
xor UO_1486 (O_1486,N_14625,N_14608);
nand UO_1487 (O_1487,N_14931,N_14454);
nand UO_1488 (O_1488,N_14474,N_14472);
nor UO_1489 (O_1489,N_14422,N_14647);
xor UO_1490 (O_1490,N_14984,N_14502);
nor UO_1491 (O_1491,N_14341,N_14938);
nor UO_1492 (O_1492,N_14528,N_14535);
nor UO_1493 (O_1493,N_14930,N_14367);
and UO_1494 (O_1494,N_14448,N_14957);
and UO_1495 (O_1495,N_14402,N_14828);
and UO_1496 (O_1496,N_14454,N_14746);
nor UO_1497 (O_1497,N_14271,N_14417);
nand UO_1498 (O_1498,N_14876,N_14811);
or UO_1499 (O_1499,N_14286,N_14411);
nor UO_1500 (O_1500,N_14493,N_14766);
or UO_1501 (O_1501,N_14381,N_14609);
or UO_1502 (O_1502,N_14500,N_14591);
nor UO_1503 (O_1503,N_14324,N_14715);
nor UO_1504 (O_1504,N_14759,N_14641);
xor UO_1505 (O_1505,N_14907,N_14890);
or UO_1506 (O_1506,N_14299,N_14860);
xor UO_1507 (O_1507,N_14496,N_14898);
nor UO_1508 (O_1508,N_14826,N_14597);
nor UO_1509 (O_1509,N_14543,N_14747);
nand UO_1510 (O_1510,N_14614,N_14969);
nand UO_1511 (O_1511,N_14572,N_14609);
xnor UO_1512 (O_1512,N_14621,N_14921);
nor UO_1513 (O_1513,N_14296,N_14355);
nand UO_1514 (O_1514,N_14870,N_14513);
xnor UO_1515 (O_1515,N_14859,N_14490);
or UO_1516 (O_1516,N_14931,N_14959);
xor UO_1517 (O_1517,N_14525,N_14477);
or UO_1518 (O_1518,N_14648,N_14697);
xnor UO_1519 (O_1519,N_14591,N_14606);
and UO_1520 (O_1520,N_14771,N_14548);
xor UO_1521 (O_1521,N_14926,N_14261);
and UO_1522 (O_1522,N_14708,N_14300);
and UO_1523 (O_1523,N_14671,N_14672);
nor UO_1524 (O_1524,N_14271,N_14918);
nand UO_1525 (O_1525,N_14848,N_14402);
nor UO_1526 (O_1526,N_14964,N_14922);
or UO_1527 (O_1527,N_14774,N_14917);
and UO_1528 (O_1528,N_14582,N_14990);
nand UO_1529 (O_1529,N_14724,N_14496);
nor UO_1530 (O_1530,N_14606,N_14686);
xor UO_1531 (O_1531,N_14314,N_14358);
nand UO_1532 (O_1532,N_14788,N_14680);
xor UO_1533 (O_1533,N_14735,N_14872);
and UO_1534 (O_1534,N_14361,N_14728);
nand UO_1535 (O_1535,N_14753,N_14611);
or UO_1536 (O_1536,N_14605,N_14377);
or UO_1537 (O_1537,N_14979,N_14587);
and UO_1538 (O_1538,N_14917,N_14985);
and UO_1539 (O_1539,N_14316,N_14954);
xor UO_1540 (O_1540,N_14259,N_14295);
or UO_1541 (O_1541,N_14405,N_14739);
xor UO_1542 (O_1542,N_14532,N_14667);
nor UO_1543 (O_1543,N_14820,N_14718);
xor UO_1544 (O_1544,N_14664,N_14266);
nand UO_1545 (O_1545,N_14952,N_14868);
xnor UO_1546 (O_1546,N_14550,N_14350);
or UO_1547 (O_1547,N_14892,N_14871);
nand UO_1548 (O_1548,N_14494,N_14545);
and UO_1549 (O_1549,N_14440,N_14859);
nand UO_1550 (O_1550,N_14457,N_14985);
or UO_1551 (O_1551,N_14291,N_14515);
and UO_1552 (O_1552,N_14934,N_14972);
and UO_1553 (O_1553,N_14590,N_14925);
xnor UO_1554 (O_1554,N_14517,N_14747);
nor UO_1555 (O_1555,N_14966,N_14710);
nand UO_1556 (O_1556,N_14600,N_14743);
nor UO_1557 (O_1557,N_14252,N_14653);
nand UO_1558 (O_1558,N_14367,N_14867);
xor UO_1559 (O_1559,N_14329,N_14790);
or UO_1560 (O_1560,N_14406,N_14667);
or UO_1561 (O_1561,N_14573,N_14475);
and UO_1562 (O_1562,N_14441,N_14772);
nor UO_1563 (O_1563,N_14315,N_14933);
nand UO_1564 (O_1564,N_14361,N_14876);
xor UO_1565 (O_1565,N_14770,N_14901);
and UO_1566 (O_1566,N_14374,N_14433);
and UO_1567 (O_1567,N_14821,N_14377);
xor UO_1568 (O_1568,N_14864,N_14467);
xor UO_1569 (O_1569,N_14882,N_14948);
nand UO_1570 (O_1570,N_14751,N_14469);
and UO_1571 (O_1571,N_14445,N_14410);
nor UO_1572 (O_1572,N_14371,N_14441);
or UO_1573 (O_1573,N_14559,N_14968);
or UO_1574 (O_1574,N_14553,N_14289);
and UO_1575 (O_1575,N_14413,N_14402);
or UO_1576 (O_1576,N_14488,N_14639);
or UO_1577 (O_1577,N_14283,N_14448);
and UO_1578 (O_1578,N_14798,N_14318);
nor UO_1579 (O_1579,N_14932,N_14305);
and UO_1580 (O_1580,N_14394,N_14606);
or UO_1581 (O_1581,N_14582,N_14937);
and UO_1582 (O_1582,N_14507,N_14758);
and UO_1583 (O_1583,N_14908,N_14259);
nor UO_1584 (O_1584,N_14523,N_14961);
xnor UO_1585 (O_1585,N_14370,N_14487);
nor UO_1586 (O_1586,N_14839,N_14923);
or UO_1587 (O_1587,N_14839,N_14290);
nand UO_1588 (O_1588,N_14286,N_14521);
xnor UO_1589 (O_1589,N_14769,N_14754);
xor UO_1590 (O_1590,N_14544,N_14318);
nor UO_1591 (O_1591,N_14414,N_14250);
or UO_1592 (O_1592,N_14523,N_14900);
xnor UO_1593 (O_1593,N_14912,N_14493);
nor UO_1594 (O_1594,N_14330,N_14759);
nand UO_1595 (O_1595,N_14306,N_14278);
nor UO_1596 (O_1596,N_14398,N_14355);
nand UO_1597 (O_1597,N_14682,N_14970);
and UO_1598 (O_1598,N_14767,N_14798);
nor UO_1599 (O_1599,N_14326,N_14518);
and UO_1600 (O_1600,N_14934,N_14503);
nand UO_1601 (O_1601,N_14693,N_14636);
or UO_1602 (O_1602,N_14406,N_14685);
nor UO_1603 (O_1603,N_14363,N_14372);
nand UO_1604 (O_1604,N_14658,N_14395);
xor UO_1605 (O_1605,N_14826,N_14734);
or UO_1606 (O_1606,N_14731,N_14436);
and UO_1607 (O_1607,N_14521,N_14485);
and UO_1608 (O_1608,N_14291,N_14695);
nor UO_1609 (O_1609,N_14722,N_14917);
nand UO_1610 (O_1610,N_14937,N_14707);
or UO_1611 (O_1611,N_14974,N_14304);
nand UO_1612 (O_1612,N_14701,N_14746);
or UO_1613 (O_1613,N_14284,N_14304);
or UO_1614 (O_1614,N_14501,N_14458);
nor UO_1615 (O_1615,N_14980,N_14464);
nor UO_1616 (O_1616,N_14951,N_14760);
nor UO_1617 (O_1617,N_14438,N_14643);
nor UO_1618 (O_1618,N_14757,N_14909);
xnor UO_1619 (O_1619,N_14842,N_14461);
and UO_1620 (O_1620,N_14903,N_14587);
nor UO_1621 (O_1621,N_14865,N_14480);
nor UO_1622 (O_1622,N_14317,N_14608);
or UO_1623 (O_1623,N_14592,N_14273);
and UO_1624 (O_1624,N_14342,N_14487);
and UO_1625 (O_1625,N_14349,N_14940);
nand UO_1626 (O_1626,N_14882,N_14991);
xnor UO_1627 (O_1627,N_14285,N_14273);
or UO_1628 (O_1628,N_14871,N_14562);
and UO_1629 (O_1629,N_14695,N_14892);
and UO_1630 (O_1630,N_14491,N_14453);
or UO_1631 (O_1631,N_14260,N_14911);
or UO_1632 (O_1632,N_14681,N_14620);
or UO_1633 (O_1633,N_14817,N_14885);
xnor UO_1634 (O_1634,N_14518,N_14836);
nand UO_1635 (O_1635,N_14256,N_14587);
nand UO_1636 (O_1636,N_14689,N_14282);
nand UO_1637 (O_1637,N_14568,N_14649);
nand UO_1638 (O_1638,N_14341,N_14352);
xnor UO_1639 (O_1639,N_14855,N_14671);
nor UO_1640 (O_1640,N_14926,N_14614);
or UO_1641 (O_1641,N_14569,N_14363);
xor UO_1642 (O_1642,N_14720,N_14816);
nor UO_1643 (O_1643,N_14849,N_14653);
nor UO_1644 (O_1644,N_14870,N_14694);
xnor UO_1645 (O_1645,N_14436,N_14290);
nor UO_1646 (O_1646,N_14361,N_14861);
xor UO_1647 (O_1647,N_14606,N_14278);
or UO_1648 (O_1648,N_14889,N_14636);
nor UO_1649 (O_1649,N_14493,N_14396);
nor UO_1650 (O_1650,N_14919,N_14922);
nand UO_1651 (O_1651,N_14844,N_14594);
and UO_1652 (O_1652,N_14980,N_14653);
nor UO_1653 (O_1653,N_14733,N_14298);
xor UO_1654 (O_1654,N_14283,N_14565);
nand UO_1655 (O_1655,N_14979,N_14795);
nor UO_1656 (O_1656,N_14641,N_14745);
nand UO_1657 (O_1657,N_14705,N_14410);
and UO_1658 (O_1658,N_14478,N_14308);
or UO_1659 (O_1659,N_14769,N_14327);
xnor UO_1660 (O_1660,N_14740,N_14435);
xnor UO_1661 (O_1661,N_14859,N_14781);
or UO_1662 (O_1662,N_14356,N_14731);
xnor UO_1663 (O_1663,N_14380,N_14581);
nand UO_1664 (O_1664,N_14547,N_14326);
xor UO_1665 (O_1665,N_14940,N_14852);
xnor UO_1666 (O_1666,N_14596,N_14397);
or UO_1667 (O_1667,N_14789,N_14324);
nand UO_1668 (O_1668,N_14292,N_14280);
xnor UO_1669 (O_1669,N_14500,N_14272);
xnor UO_1670 (O_1670,N_14952,N_14962);
nor UO_1671 (O_1671,N_14701,N_14613);
nand UO_1672 (O_1672,N_14847,N_14389);
and UO_1673 (O_1673,N_14568,N_14378);
nand UO_1674 (O_1674,N_14925,N_14956);
or UO_1675 (O_1675,N_14656,N_14797);
or UO_1676 (O_1676,N_14375,N_14632);
and UO_1677 (O_1677,N_14624,N_14442);
nor UO_1678 (O_1678,N_14837,N_14364);
nor UO_1679 (O_1679,N_14597,N_14340);
or UO_1680 (O_1680,N_14284,N_14850);
or UO_1681 (O_1681,N_14465,N_14633);
nor UO_1682 (O_1682,N_14687,N_14386);
nor UO_1683 (O_1683,N_14366,N_14817);
nand UO_1684 (O_1684,N_14427,N_14301);
xor UO_1685 (O_1685,N_14895,N_14304);
or UO_1686 (O_1686,N_14475,N_14891);
and UO_1687 (O_1687,N_14995,N_14395);
and UO_1688 (O_1688,N_14683,N_14273);
nand UO_1689 (O_1689,N_14862,N_14298);
nor UO_1690 (O_1690,N_14282,N_14922);
nor UO_1691 (O_1691,N_14553,N_14654);
nor UO_1692 (O_1692,N_14266,N_14709);
nor UO_1693 (O_1693,N_14950,N_14438);
xor UO_1694 (O_1694,N_14420,N_14327);
nor UO_1695 (O_1695,N_14365,N_14549);
or UO_1696 (O_1696,N_14434,N_14584);
or UO_1697 (O_1697,N_14901,N_14915);
xor UO_1698 (O_1698,N_14409,N_14282);
or UO_1699 (O_1699,N_14980,N_14738);
or UO_1700 (O_1700,N_14274,N_14729);
nand UO_1701 (O_1701,N_14798,N_14316);
nor UO_1702 (O_1702,N_14713,N_14387);
nor UO_1703 (O_1703,N_14482,N_14908);
or UO_1704 (O_1704,N_14563,N_14766);
or UO_1705 (O_1705,N_14363,N_14389);
and UO_1706 (O_1706,N_14850,N_14721);
nand UO_1707 (O_1707,N_14310,N_14767);
nor UO_1708 (O_1708,N_14545,N_14832);
nor UO_1709 (O_1709,N_14424,N_14299);
or UO_1710 (O_1710,N_14616,N_14460);
nor UO_1711 (O_1711,N_14619,N_14572);
xnor UO_1712 (O_1712,N_14789,N_14567);
nand UO_1713 (O_1713,N_14862,N_14644);
or UO_1714 (O_1714,N_14753,N_14844);
nand UO_1715 (O_1715,N_14328,N_14557);
or UO_1716 (O_1716,N_14327,N_14287);
xor UO_1717 (O_1717,N_14826,N_14845);
nor UO_1718 (O_1718,N_14514,N_14993);
xor UO_1719 (O_1719,N_14880,N_14446);
xor UO_1720 (O_1720,N_14690,N_14849);
nor UO_1721 (O_1721,N_14808,N_14974);
nor UO_1722 (O_1722,N_14754,N_14687);
nand UO_1723 (O_1723,N_14867,N_14595);
and UO_1724 (O_1724,N_14457,N_14321);
and UO_1725 (O_1725,N_14387,N_14486);
and UO_1726 (O_1726,N_14776,N_14622);
nor UO_1727 (O_1727,N_14913,N_14698);
nand UO_1728 (O_1728,N_14842,N_14823);
nand UO_1729 (O_1729,N_14801,N_14683);
xor UO_1730 (O_1730,N_14913,N_14461);
and UO_1731 (O_1731,N_14438,N_14806);
or UO_1732 (O_1732,N_14889,N_14822);
or UO_1733 (O_1733,N_14809,N_14713);
nor UO_1734 (O_1734,N_14676,N_14431);
nor UO_1735 (O_1735,N_14294,N_14953);
nor UO_1736 (O_1736,N_14610,N_14431);
and UO_1737 (O_1737,N_14653,N_14966);
nand UO_1738 (O_1738,N_14762,N_14602);
or UO_1739 (O_1739,N_14388,N_14937);
nand UO_1740 (O_1740,N_14960,N_14866);
and UO_1741 (O_1741,N_14357,N_14294);
or UO_1742 (O_1742,N_14921,N_14539);
or UO_1743 (O_1743,N_14766,N_14859);
or UO_1744 (O_1744,N_14419,N_14945);
or UO_1745 (O_1745,N_14832,N_14716);
or UO_1746 (O_1746,N_14430,N_14527);
nor UO_1747 (O_1747,N_14466,N_14434);
and UO_1748 (O_1748,N_14285,N_14694);
xor UO_1749 (O_1749,N_14871,N_14658);
or UO_1750 (O_1750,N_14740,N_14391);
nand UO_1751 (O_1751,N_14766,N_14741);
nand UO_1752 (O_1752,N_14255,N_14874);
or UO_1753 (O_1753,N_14670,N_14810);
nor UO_1754 (O_1754,N_14469,N_14860);
xnor UO_1755 (O_1755,N_14757,N_14877);
nand UO_1756 (O_1756,N_14915,N_14632);
xor UO_1757 (O_1757,N_14894,N_14333);
and UO_1758 (O_1758,N_14268,N_14460);
nor UO_1759 (O_1759,N_14626,N_14848);
nor UO_1760 (O_1760,N_14372,N_14387);
nand UO_1761 (O_1761,N_14739,N_14358);
and UO_1762 (O_1762,N_14360,N_14404);
xnor UO_1763 (O_1763,N_14741,N_14532);
nand UO_1764 (O_1764,N_14988,N_14982);
and UO_1765 (O_1765,N_14775,N_14332);
nor UO_1766 (O_1766,N_14768,N_14401);
or UO_1767 (O_1767,N_14398,N_14526);
and UO_1768 (O_1768,N_14450,N_14329);
nor UO_1769 (O_1769,N_14579,N_14942);
and UO_1770 (O_1770,N_14428,N_14975);
nand UO_1771 (O_1771,N_14645,N_14360);
nand UO_1772 (O_1772,N_14817,N_14986);
or UO_1773 (O_1773,N_14982,N_14996);
and UO_1774 (O_1774,N_14634,N_14593);
and UO_1775 (O_1775,N_14653,N_14576);
nand UO_1776 (O_1776,N_14853,N_14362);
or UO_1777 (O_1777,N_14777,N_14639);
xor UO_1778 (O_1778,N_14944,N_14617);
nor UO_1779 (O_1779,N_14684,N_14653);
or UO_1780 (O_1780,N_14772,N_14574);
nand UO_1781 (O_1781,N_14534,N_14680);
xnor UO_1782 (O_1782,N_14671,N_14795);
xnor UO_1783 (O_1783,N_14887,N_14317);
xor UO_1784 (O_1784,N_14383,N_14501);
xor UO_1785 (O_1785,N_14850,N_14761);
nor UO_1786 (O_1786,N_14587,N_14583);
nand UO_1787 (O_1787,N_14710,N_14890);
and UO_1788 (O_1788,N_14599,N_14285);
or UO_1789 (O_1789,N_14533,N_14394);
xor UO_1790 (O_1790,N_14854,N_14956);
nor UO_1791 (O_1791,N_14573,N_14618);
and UO_1792 (O_1792,N_14596,N_14265);
and UO_1793 (O_1793,N_14688,N_14712);
and UO_1794 (O_1794,N_14851,N_14699);
nor UO_1795 (O_1795,N_14306,N_14450);
nand UO_1796 (O_1796,N_14746,N_14772);
nor UO_1797 (O_1797,N_14403,N_14773);
or UO_1798 (O_1798,N_14908,N_14990);
nand UO_1799 (O_1799,N_14902,N_14940);
xnor UO_1800 (O_1800,N_14554,N_14615);
xor UO_1801 (O_1801,N_14697,N_14565);
nor UO_1802 (O_1802,N_14702,N_14616);
or UO_1803 (O_1803,N_14613,N_14409);
and UO_1804 (O_1804,N_14902,N_14272);
and UO_1805 (O_1805,N_14852,N_14856);
nor UO_1806 (O_1806,N_14533,N_14884);
nor UO_1807 (O_1807,N_14540,N_14381);
nor UO_1808 (O_1808,N_14927,N_14609);
nor UO_1809 (O_1809,N_14662,N_14700);
and UO_1810 (O_1810,N_14259,N_14571);
and UO_1811 (O_1811,N_14385,N_14925);
nor UO_1812 (O_1812,N_14579,N_14689);
or UO_1813 (O_1813,N_14975,N_14603);
or UO_1814 (O_1814,N_14879,N_14401);
xnor UO_1815 (O_1815,N_14981,N_14462);
xnor UO_1816 (O_1816,N_14288,N_14656);
and UO_1817 (O_1817,N_14255,N_14785);
nor UO_1818 (O_1818,N_14544,N_14892);
or UO_1819 (O_1819,N_14849,N_14290);
nand UO_1820 (O_1820,N_14304,N_14576);
or UO_1821 (O_1821,N_14439,N_14342);
xnor UO_1822 (O_1822,N_14365,N_14284);
xnor UO_1823 (O_1823,N_14450,N_14563);
and UO_1824 (O_1824,N_14354,N_14517);
nor UO_1825 (O_1825,N_14320,N_14971);
or UO_1826 (O_1826,N_14366,N_14434);
nand UO_1827 (O_1827,N_14566,N_14937);
nor UO_1828 (O_1828,N_14995,N_14773);
nor UO_1829 (O_1829,N_14380,N_14888);
nor UO_1830 (O_1830,N_14273,N_14378);
and UO_1831 (O_1831,N_14842,N_14367);
xnor UO_1832 (O_1832,N_14448,N_14797);
nand UO_1833 (O_1833,N_14657,N_14861);
nand UO_1834 (O_1834,N_14498,N_14800);
and UO_1835 (O_1835,N_14333,N_14436);
nand UO_1836 (O_1836,N_14587,N_14481);
nor UO_1837 (O_1837,N_14805,N_14773);
and UO_1838 (O_1838,N_14381,N_14705);
nand UO_1839 (O_1839,N_14405,N_14627);
or UO_1840 (O_1840,N_14523,N_14440);
nand UO_1841 (O_1841,N_14333,N_14980);
xnor UO_1842 (O_1842,N_14560,N_14896);
nand UO_1843 (O_1843,N_14843,N_14979);
nor UO_1844 (O_1844,N_14396,N_14569);
nand UO_1845 (O_1845,N_14898,N_14696);
nor UO_1846 (O_1846,N_14894,N_14639);
xor UO_1847 (O_1847,N_14700,N_14831);
xnor UO_1848 (O_1848,N_14839,N_14474);
or UO_1849 (O_1849,N_14709,N_14871);
nor UO_1850 (O_1850,N_14654,N_14402);
and UO_1851 (O_1851,N_14573,N_14538);
nand UO_1852 (O_1852,N_14268,N_14747);
and UO_1853 (O_1853,N_14449,N_14754);
nor UO_1854 (O_1854,N_14531,N_14373);
xor UO_1855 (O_1855,N_14671,N_14743);
nand UO_1856 (O_1856,N_14887,N_14925);
xor UO_1857 (O_1857,N_14561,N_14263);
xnor UO_1858 (O_1858,N_14703,N_14699);
or UO_1859 (O_1859,N_14253,N_14506);
and UO_1860 (O_1860,N_14627,N_14703);
nand UO_1861 (O_1861,N_14853,N_14331);
nand UO_1862 (O_1862,N_14747,N_14967);
nor UO_1863 (O_1863,N_14844,N_14762);
nor UO_1864 (O_1864,N_14615,N_14660);
nand UO_1865 (O_1865,N_14668,N_14940);
or UO_1866 (O_1866,N_14869,N_14828);
nor UO_1867 (O_1867,N_14708,N_14409);
or UO_1868 (O_1868,N_14517,N_14535);
nor UO_1869 (O_1869,N_14462,N_14312);
xor UO_1870 (O_1870,N_14925,N_14451);
and UO_1871 (O_1871,N_14616,N_14957);
xor UO_1872 (O_1872,N_14340,N_14994);
nand UO_1873 (O_1873,N_14369,N_14506);
xor UO_1874 (O_1874,N_14569,N_14910);
nor UO_1875 (O_1875,N_14992,N_14620);
xnor UO_1876 (O_1876,N_14771,N_14366);
or UO_1877 (O_1877,N_14841,N_14982);
and UO_1878 (O_1878,N_14351,N_14719);
xor UO_1879 (O_1879,N_14591,N_14270);
nand UO_1880 (O_1880,N_14466,N_14975);
nor UO_1881 (O_1881,N_14390,N_14281);
and UO_1882 (O_1882,N_14763,N_14980);
or UO_1883 (O_1883,N_14799,N_14620);
xnor UO_1884 (O_1884,N_14528,N_14812);
or UO_1885 (O_1885,N_14629,N_14620);
and UO_1886 (O_1886,N_14695,N_14440);
or UO_1887 (O_1887,N_14383,N_14910);
nand UO_1888 (O_1888,N_14461,N_14369);
nand UO_1889 (O_1889,N_14473,N_14292);
or UO_1890 (O_1890,N_14318,N_14454);
or UO_1891 (O_1891,N_14675,N_14290);
nor UO_1892 (O_1892,N_14498,N_14666);
nand UO_1893 (O_1893,N_14787,N_14384);
nand UO_1894 (O_1894,N_14665,N_14909);
nor UO_1895 (O_1895,N_14862,N_14792);
nor UO_1896 (O_1896,N_14385,N_14810);
nor UO_1897 (O_1897,N_14431,N_14863);
xor UO_1898 (O_1898,N_14716,N_14435);
or UO_1899 (O_1899,N_14727,N_14999);
xor UO_1900 (O_1900,N_14629,N_14506);
and UO_1901 (O_1901,N_14993,N_14396);
and UO_1902 (O_1902,N_14808,N_14835);
xnor UO_1903 (O_1903,N_14755,N_14712);
nor UO_1904 (O_1904,N_14462,N_14285);
xor UO_1905 (O_1905,N_14695,N_14612);
or UO_1906 (O_1906,N_14269,N_14505);
and UO_1907 (O_1907,N_14359,N_14795);
xor UO_1908 (O_1908,N_14430,N_14571);
or UO_1909 (O_1909,N_14334,N_14753);
and UO_1910 (O_1910,N_14893,N_14427);
or UO_1911 (O_1911,N_14746,N_14674);
or UO_1912 (O_1912,N_14965,N_14469);
nor UO_1913 (O_1913,N_14854,N_14736);
nand UO_1914 (O_1914,N_14996,N_14647);
nor UO_1915 (O_1915,N_14384,N_14676);
nor UO_1916 (O_1916,N_14501,N_14583);
or UO_1917 (O_1917,N_14851,N_14963);
nor UO_1918 (O_1918,N_14898,N_14982);
nor UO_1919 (O_1919,N_14648,N_14443);
nand UO_1920 (O_1920,N_14258,N_14723);
xnor UO_1921 (O_1921,N_14433,N_14305);
and UO_1922 (O_1922,N_14907,N_14982);
xor UO_1923 (O_1923,N_14340,N_14983);
nor UO_1924 (O_1924,N_14899,N_14990);
and UO_1925 (O_1925,N_14982,N_14262);
nor UO_1926 (O_1926,N_14828,N_14372);
xor UO_1927 (O_1927,N_14475,N_14369);
and UO_1928 (O_1928,N_14341,N_14408);
and UO_1929 (O_1929,N_14972,N_14427);
and UO_1930 (O_1930,N_14567,N_14595);
xnor UO_1931 (O_1931,N_14390,N_14252);
and UO_1932 (O_1932,N_14479,N_14710);
and UO_1933 (O_1933,N_14968,N_14783);
nand UO_1934 (O_1934,N_14927,N_14645);
and UO_1935 (O_1935,N_14414,N_14818);
or UO_1936 (O_1936,N_14883,N_14739);
nor UO_1937 (O_1937,N_14403,N_14485);
nand UO_1938 (O_1938,N_14525,N_14576);
or UO_1939 (O_1939,N_14949,N_14437);
or UO_1940 (O_1940,N_14303,N_14619);
nand UO_1941 (O_1941,N_14483,N_14615);
nor UO_1942 (O_1942,N_14592,N_14850);
nand UO_1943 (O_1943,N_14547,N_14833);
nand UO_1944 (O_1944,N_14339,N_14966);
nand UO_1945 (O_1945,N_14876,N_14854);
nor UO_1946 (O_1946,N_14440,N_14939);
or UO_1947 (O_1947,N_14436,N_14338);
nand UO_1948 (O_1948,N_14893,N_14572);
nand UO_1949 (O_1949,N_14580,N_14351);
xor UO_1950 (O_1950,N_14685,N_14315);
and UO_1951 (O_1951,N_14781,N_14886);
or UO_1952 (O_1952,N_14998,N_14487);
nand UO_1953 (O_1953,N_14912,N_14666);
nor UO_1954 (O_1954,N_14419,N_14428);
or UO_1955 (O_1955,N_14876,N_14567);
or UO_1956 (O_1956,N_14332,N_14834);
or UO_1957 (O_1957,N_14390,N_14658);
or UO_1958 (O_1958,N_14921,N_14653);
and UO_1959 (O_1959,N_14418,N_14265);
nor UO_1960 (O_1960,N_14361,N_14777);
and UO_1961 (O_1961,N_14624,N_14611);
and UO_1962 (O_1962,N_14625,N_14769);
nand UO_1963 (O_1963,N_14327,N_14479);
and UO_1964 (O_1964,N_14746,N_14764);
and UO_1965 (O_1965,N_14982,N_14710);
and UO_1966 (O_1966,N_14279,N_14783);
xnor UO_1967 (O_1967,N_14401,N_14981);
and UO_1968 (O_1968,N_14393,N_14781);
nand UO_1969 (O_1969,N_14540,N_14876);
nand UO_1970 (O_1970,N_14530,N_14564);
or UO_1971 (O_1971,N_14379,N_14489);
xnor UO_1972 (O_1972,N_14753,N_14700);
and UO_1973 (O_1973,N_14921,N_14983);
or UO_1974 (O_1974,N_14732,N_14690);
xor UO_1975 (O_1975,N_14418,N_14415);
nor UO_1976 (O_1976,N_14271,N_14951);
nand UO_1977 (O_1977,N_14831,N_14252);
nand UO_1978 (O_1978,N_14917,N_14754);
nor UO_1979 (O_1979,N_14351,N_14842);
xor UO_1980 (O_1980,N_14361,N_14835);
or UO_1981 (O_1981,N_14612,N_14780);
nand UO_1982 (O_1982,N_14265,N_14483);
nand UO_1983 (O_1983,N_14701,N_14744);
and UO_1984 (O_1984,N_14490,N_14354);
xor UO_1985 (O_1985,N_14932,N_14737);
and UO_1986 (O_1986,N_14843,N_14252);
nand UO_1987 (O_1987,N_14775,N_14921);
xor UO_1988 (O_1988,N_14647,N_14848);
and UO_1989 (O_1989,N_14574,N_14388);
nand UO_1990 (O_1990,N_14853,N_14867);
xor UO_1991 (O_1991,N_14600,N_14390);
nand UO_1992 (O_1992,N_14482,N_14362);
or UO_1993 (O_1993,N_14540,N_14840);
xnor UO_1994 (O_1994,N_14601,N_14314);
or UO_1995 (O_1995,N_14396,N_14977);
nand UO_1996 (O_1996,N_14885,N_14469);
xor UO_1997 (O_1997,N_14842,N_14482);
nand UO_1998 (O_1998,N_14891,N_14262);
and UO_1999 (O_1999,N_14955,N_14775);
endmodule