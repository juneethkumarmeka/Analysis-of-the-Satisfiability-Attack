module basic_1000_10000_1500_4_levels_1xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
or U0 (N_0,In_364,In_844);
and U1 (N_1,In_326,In_622);
and U2 (N_2,In_724,In_866);
and U3 (N_3,In_898,In_182);
and U4 (N_4,In_376,In_715);
and U5 (N_5,In_274,In_15);
or U6 (N_6,In_610,In_913);
and U7 (N_7,In_664,In_946);
nand U8 (N_8,In_737,In_382);
or U9 (N_9,In_648,In_450);
and U10 (N_10,In_720,In_49);
or U11 (N_11,In_84,In_550);
or U12 (N_12,In_782,In_354);
nor U13 (N_13,In_823,In_551);
and U14 (N_14,In_423,In_53);
and U15 (N_15,In_22,In_832);
and U16 (N_16,In_224,In_938);
nand U17 (N_17,In_717,In_620);
or U18 (N_18,In_116,In_411);
and U19 (N_19,In_840,In_583);
or U20 (N_20,In_489,In_691);
nor U21 (N_21,In_799,In_311);
or U22 (N_22,In_833,In_179);
or U23 (N_23,In_345,In_649);
and U24 (N_24,In_632,In_178);
nor U25 (N_25,In_974,In_694);
nand U26 (N_26,In_148,In_5);
nor U27 (N_27,In_779,In_646);
nor U28 (N_28,In_687,In_962);
and U29 (N_29,In_122,In_519);
or U30 (N_30,In_81,In_954);
nand U31 (N_31,In_305,In_18);
nor U32 (N_32,In_984,In_787);
or U33 (N_33,In_983,In_363);
and U34 (N_34,In_212,In_422);
nor U35 (N_35,In_156,In_826);
nor U36 (N_36,In_307,In_706);
nand U37 (N_37,In_856,In_681);
nor U38 (N_38,In_536,In_416);
nand U39 (N_39,In_805,In_410);
nor U40 (N_40,In_758,In_278);
and U41 (N_41,In_668,In_659);
nor U42 (N_42,In_356,In_456);
nor U43 (N_43,In_757,In_524);
and U44 (N_44,In_702,In_930);
and U45 (N_45,In_218,In_552);
nor U46 (N_46,In_786,In_240);
or U47 (N_47,In_636,In_566);
xnor U48 (N_48,In_557,In_697);
or U49 (N_49,In_859,In_986);
and U50 (N_50,In_184,In_812);
nand U51 (N_51,In_993,In_380);
nand U52 (N_52,In_432,In_431);
and U53 (N_53,In_727,In_498);
and U54 (N_54,In_474,In_795);
nand U55 (N_55,In_368,In_868);
nand U56 (N_56,In_997,In_292);
nand U57 (N_57,In_3,In_526);
and U58 (N_58,In_371,In_546);
or U59 (N_59,In_52,In_407);
nor U60 (N_60,In_872,In_186);
nor U61 (N_61,In_471,In_943);
nand U62 (N_62,In_333,In_578);
or U63 (N_63,In_655,In_438);
nand U64 (N_64,In_661,In_304);
nand U65 (N_65,In_281,In_468);
nand U66 (N_66,In_940,In_650);
or U67 (N_67,In_197,In_493);
nor U68 (N_68,In_568,In_637);
nand U69 (N_69,In_521,In_483);
or U70 (N_70,In_205,In_150);
or U71 (N_71,In_486,In_809);
nor U72 (N_72,In_562,In_323);
and U73 (N_73,In_574,In_104);
nor U74 (N_74,In_950,In_109);
or U75 (N_75,In_666,In_751);
nand U76 (N_76,In_452,In_891);
nor U77 (N_77,In_221,In_667);
or U78 (N_78,In_759,In_408);
nand U79 (N_79,In_231,In_630);
nand U80 (N_80,In_417,In_260);
nand U81 (N_81,In_596,In_564);
nor U82 (N_82,In_701,In_634);
or U83 (N_83,In_390,In_282);
nand U84 (N_84,In_245,In_472);
or U85 (N_85,In_905,In_462);
nand U86 (N_86,In_445,In_679);
and U87 (N_87,In_624,In_932);
nor U88 (N_88,In_436,In_537);
and U89 (N_89,In_617,In_527);
and U90 (N_90,In_143,In_230);
nand U91 (N_91,In_480,In_455);
and U92 (N_92,In_154,In_185);
nand U93 (N_93,In_277,In_236);
nor U94 (N_94,In_175,In_645);
and U95 (N_95,In_969,In_688);
nand U96 (N_96,In_439,In_226);
nand U97 (N_97,In_194,In_343);
or U98 (N_98,In_190,In_816);
or U99 (N_99,In_276,In_286);
and U100 (N_100,In_99,In_543);
nand U101 (N_101,In_2,In_61);
nor U102 (N_102,In_640,In_421);
and U103 (N_103,In_373,In_34);
or U104 (N_104,In_324,In_528);
and U105 (N_105,In_766,In_754);
nor U106 (N_106,In_682,In_20);
or U107 (N_107,In_37,In_57);
nor U108 (N_108,In_676,In_894);
nor U109 (N_109,In_935,In_855);
or U110 (N_110,In_394,In_152);
or U111 (N_111,In_616,In_604);
or U112 (N_112,In_302,In_842);
nand U113 (N_113,In_712,In_1);
nor U114 (N_114,In_359,In_794);
nand U115 (N_115,In_476,In_982);
and U116 (N_116,In_163,In_520);
nand U117 (N_117,In_31,In_658);
nand U118 (N_118,In_491,In_405);
and U119 (N_119,In_131,In_987);
and U120 (N_120,In_347,In_931);
or U121 (N_121,In_510,In_698);
and U122 (N_122,In_329,In_248);
or U123 (N_123,In_171,In_815);
and U124 (N_124,In_484,In_871);
nand U125 (N_125,In_770,In_23);
nor U126 (N_126,In_629,In_0);
nand U127 (N_127,In_870,In_889);
and U128 (N_128,In_119,In_523);
and U129 (N_129,In_747,In_796);
and U130 (N_130,In_328,In_80);
nor U131 (N_131,In_27,In_124);
or U132 (N_132,In_399,In_879);
nor U133 (N_133,In_752,In_909);
nand U134 (N_134,In_692,In_587);
nand U135 (N_135,In_780,In_188);
and U136 (N_136,In_541,In_398);
nand U137 (N_137,In_19,In_39);
nand U138 (N_138,In_426,In_440);
or U139 (N_139,In_378,In_482);
or U140 (N_140,In_808,In_584);
or U141 (N_141,In_675,In_334);
nand U142 (N_142,In_25,In_626);
nor U143 (N_143,In_209,In_554);
or U144 (N_144,In_424,In_453);
nor U145 (N_145,In_990,In_743);
nand U146 (N_146,In_252,In_92);
or U147 (N_147,In_975,In_90);
and U148 (N_148,In_967,In_925);
nor U149 (N_149,In_873,In_707);
or U150 (N_150,In_841,In_933);
or U151 (N_151,In_853,In_215);
or U152 (N_152,In_74,In_643);
or U153 (N_153,In_348,In_114);
or U154 (N_154,In_690,In_330);
and U155 (N_155,In_258,In_279);
nand U156 (N_156,In_801,In_362);
or U157 (N_157,In_7,In_538);
and U158 (N_158,In_768,In_798);
and U159 (N_159,In_788,In_415);
or U160 (N_160,In_435,In_242);
nor U161 (N_161,In_511,In_619);
nand U162 (N_162,In_864,In_40);
and U163 (N_163,In_852,In_710);
and U164 (N_164,In_485,In_621);
nor U165 (N_165,In_800,In_953);
and U166 (N_166,In_819,In_729);
nand U167 (N_167,In_265,In_669);
and U168 (N_168,In_944,In_825);
and U169 (N_169,In_641,In_945);
or U170 (N_170,In_180,In_534);
xnor U171 (N_171,In_125,In_571);
or U172 (N_172,In_10,In_822);
or U173 (N_173,In_942,In_294);
or U174 (N_174,In_409,In_761);
nand U175 (N_175,In_771,In_392);
and U176 (N_176,In_911,In_341);
and U177 (N_177,In_48,In_259);
or U178 (N_178,In_60,In_241);
nand U179 (N_179,In_589,In_929);
and U180 (N_180,In_860,In_836);
or U181 (N_181,In_389,In_234);
or U182 (N_182,In_978,In_300);
nand U183 (N_183,In_652,In_593);
nor U184 (N_184,In_777,In_736);
nand U185 (N_185,In_900,In_660);
nand U186 (N_186,In_875,In_906);
nand U187 (N_187,In_530,In_569);
and U188 (N_188,In_420,In_899);
nor U189 (N_189,In_837,In_235);
nand U190 (N_190,In_728,In_463);
xnor U191 (N_191,In_955,In_887);
nor U192 (N_192,In_262,In_169);
and U193 (N_193,In_187,In_916);
or U194 (N_194,In_928,In_360);
nor U195 (N_195,In_673,In_704);
nand U196 (N_196,In_193,In_59);
nand U197 (N_197,In_876,In_293);
and U198 (N_198,In_402,In_817);
nand U199 (N_199,In_988,In_6);
nor U200 (N_200,In_699,In_902);
nor U201 (N_201,In_361,In_981);
and U202 (N_202,In_232,In_159);
and U203 (N_203,In_723,In_778);
or U204 (N_204,In_56,In_772);
nand U205 (N_205,In_83,In_949);
nor U206 (N_206,In_63,In_129);
or U207 (N_207,In_95,In_592);
nor U208 (N_208,In_989,In_760);
nor U209 (N_209,In_920,In_117);
or U210 (N_210,In_722,In_149);
nor U211 (N_211,In_956,In_651);
nor U212 (N_212,In_556,In_830);
nor U213 (N_213,In_708,In_609);
nand U214 (N_214,In_273,In_677);
nand U215 (N_215,In_238,In_448);
nor U216 (N_216,In_884,In_217);
nand U217 (N_217,In_924,In_379);
or U218 (N_218,In_202,In_845);
or U219 (N_219,In_346,In_140);
nor U220 (N_220,In_141,In_525);
and U221 (N_221,In_674,In_544);
nand U222 (N_222,In_665,In_518);
and U223 (N_223,In_883,In_222);
and U224 (N_224,In_45,In_36);
or U225 (N_225,In_607,In_517);
nand U226 (N_226,In_979,In_77);
or U227 (N_227,In_939,In_586);
nand U228 (N_228,In_581,In_384);
nor U229 (N_229,In_266,In_144);
and U230 (N_230,In_357,In_97);
and U231 (N_231,In_671,In_400);
nor U232 (N_232,In_598,In_773);
nor U233 (N_233,In_500,In_613);
nor U234 (N_234,In_765,In_406);
or U235 (N_235,In_921,In_608);
and U236 (N_236,In_730,In_96);
nor U237 (N_237,In_827,In_908);
nand U238 (N_238,In_43,In_66);
nand U239 (N_239,In_216,In_315);
or U240 (N_240,In_804,In_910);
nor U241 (N_241,In_82,In_857);
or U242 (N_242,In_515,In_820);
or U243 (N_243,In_638,In_12);
nor U244 (N_244,In_507,In_907);
nor U245 (N_245,In_385,In_590);
nand U246 (N_246,In_393,In_427);
and U247 (N_247,In_995,In_9);
or U248 (N_248,In_366,In_211);
nor U249 (N_249,In_320,In_28);
nor U250 (N_250,In_433,In_465);
nand U251 (N_251,In_880,In_458);
or U252 (N_252,In_46,In_504);
nor U253 (N_253,In_350,In_107);
nor U254 (N_254,In_247,In_203);
nor U255 (N_255,In_503,In_656);
or U256 (N_256,In_888,In_851);
nand U257 (N_257,In_996,In_775);
nor U258 (N_258,In_631,In_892);
or U259 (N_259,In_767,In_280);
or U260 (N_260,In_404,In_915);
nand U261 (N_261,In_549,In_881);
or U262 (N_262,In_683,In_602);
or U263 (N_263,In_381,In_93);
nor U264 (N_264,In_591,In_901);
and U265 (N_265,In_64,In_336);
or U266 (N_266,In_742,In_897);
nor U267 (N_267,In_719,In_806);
or U268 (N_268,In_460,In_199);
and U269 (N_269,In_110,In_106);
nor U270 (N_270,In_306,In_89);
nor U271 (N_271,In_999,In_615);
nand U272 (N_272,In_600,In_267);
nor U273 (N_273,In_684,In_824);
or U274 (N_274,In_764,In_162);
nor U275 (N_275,In_103,In_250);
nor U276 (N_276,In_792,In_228);
or U277 (N_277,In_223,In_86);
and U278 (N_278,In_29,In_919);
or U279 (N_279,In_867,In_370);
and U280 (N_280,In_173,In_744);
nand U281 (N_281,In_803,In_966);
or U282 (N_282,In_91,In_878);
nand U283 (N_283,In_134,In_755);
or U284 (N_284,In_672,In_700);
or U285 (N_285,In_219,In_58);
nor U286 (N_286,In_992,In_303);
and U287 (N_287,In_575,In_108);
and U288 (N_288,In_735,In_539);
nand U289 (N_289,In_142,In_115);
nor U290 (N_290,In_275,In_255);
nand U291 (N_291,In_101,In_991);
and U292 (N_292,In_998,In_297);
and U293 (N_293,In_290,In_332);
nor U294 (N_294,In_85,In_695);
or U295 (N_295,In_391,In_325);
or U296 (N_296,In_738,In_490);
nand U297 (N_297,In_33,In_831);
or U298 (N_298,In_959,In_44);
and U299 (N_299,In_128,In_963);
or U300 (N_300,In_828,In_951);
or U301 (N_301,In_451,In_196);
nand U302 (N_302,In_685,In_317);
nor U303 (N_303,In_76,In_318);
xor U304 (N_304,In_312,In_877);
nor U305 (N_305,In_781,In_13);
or U306 (N_306,In_567,In_705);
and U307 (N_307,In_477,In_753);
nor U308 (N_308,In_869,In_958);
nor U309 (N_309,In_207,In_288);
or U310 (N_310,In_430,In_8);
nand U311 (N_311,In_383,In_434);
nor U312 (N_312,In_151,In_479);
nor U313 (N_313,In_746,In_352);
nor U314 (N_314,In_941,In_35);
and U315 (N_315,In_721,In_627);
nand U316 (N_316,In_397,In_446);
nand U317 (N_317,In_413,In_818);
or U318 (N_318,In_813,In_338);
nor U319 (N_319,In_88,In_130);
nor U320 (N_320,In_79,In_377);
nor U321 (N_321,In_291,In_54);
nand U322 (N_322,In_139,In_965);
and U323 (N_323,In_917,In_459);
and U324 (N_324,In_32,In_313);
and U325 (N_325,In_111,In_30);
nand U326 (N_326,In_51,In_848);
or U327 (N_327,In_612,In_654);
nor U328 (N_328,In_829,In_309);
or U329 (N_329,In_337,In_740);
nor U330 (N_330,In_895,In_548);
or U331 (N_331,In_4,In_478);
or U332 (N_332,In_138,In_442);
xor U333 (N_333,In_611,In_322);
nand U334 (N_334,In_663,In_834);
nor U335 (N_335,In_153,In_614);
or U336 (N_336,In_69,In_271);
nand U337 (N_337,In_461,In_257);
nand U338 (N_338,In_481,In_789);
nand U339 (N_339,In_172,In_120);
nor U340 (N_340,In_670,In_396);
nand U341 (N_341,In_749,In_146);
nor U342 (N_342,In_268,In_167);
and U343 (N_343,In_263,In_447);
and U344 (N_344,In_387,In_299);
nor U345 (N_345,In_301,In_344);
nor U346 (N_346,In_189,In_662);
and U347 (N_347,In_741,In_952);
and U348 (N_348,In_62,In_308);
and U349 (N_349,In_810,In_201);
or U350 (N_350,In_559,In_145);
and U351 (N_351,In_283,In_846);
and U352 (N_352,In_532,In_168);
and U353 (N_353,In_547,In_386);
nand U354 (N_354,In_985,In_603);
nor U355 (N_355,In_923,In_961);
nand U356 (N_356,In_793,In_594);
or U357 (N_357,In_467,In_914);
and U358 (N_358,In_821,In_797);
nand U359 (N_359,In_229,In_136);
nand U360 (N_360,In_287,In_776);
nor U361 (N_361,In_441,In_748);
nand U362 (N_362,In_769,In_714);
nor U363 (N_363,In_339,In_633);
nor U364 (N_364,In_680,In_335);
nor U365 (N_365,In_936,In_198);
and U366 (N_366,In_284,In_375);
nor U367 (N_367,In_733,In_355);
nand U368 (N_368,In_785,In_165);
and U369 (N_369,In_560,In_783);
or U370 (N_370,In_582,In_542);
or U371 (N_371,In_739,In_960);
or U372 (N_372,In_644,In_105);
nor U373 (N_373,In_157,In_210);
or U374 (N_374,In_395,In_87);
and U375 (N_375,In_270,In_904);
or U376 (N_376,In_55,In_401);
or U377 (N_377,In_573,In_718);
xnor U378 (N_378,In_865,In_327);
nand U379 (N_379,In_170,In_558);
nor U380 (N_380,In_147,In_412);
nor U381 (N_381,In_369,In_516);
nand U382 (N_382,In_725,In_449);
nand U383 (N_383,In_726,In_968);
and U384 (N_384,In_678,In_425);
nand U385 (N_385,In_428,In_206);
nand U386 (N_386,In_686,In_454);
nor U387 (N_387,In_254,In_374);
and U388 (N_388,In_164,In_522);
nand U389 (N_389,In_289,In_264);
nor U390 (N_390,In_545,In_994);
or U391 (N_391,In_903,In_912);
nand U392 (N_392,In_711,In_272);
or U393 (N_393,In_208,In_50);
nor U394 (N_394,In_756,In_811);
nand U395 (N_395,In_488,In_126);
nor U396 (N_396,In_863,In_213);
nor U397 (N_397,In_802,In_296);
nor U398 (N_398,In_38,In_508);
and U399 (N_399,In_937,In_166);
or U400 (N_400,In_763,In_174);
or U401 (N_401,In_750,In_65);
or U402 (N_402,In_703,In_896);
nand U403 (N_403,In_716,In_599);
nand U404 (N_404,In_429,In_495);
and U405 (N_405,In_886,In_403);
or U406 (N_406,In_843,In_319);
nor U407 (N_407,In_595,In_70);
nand U408 (N_408,In_285,In_893);
nand U409 (N_409,In_732,In_580);
and U410 (N_410,In_225,In_100);
nand U411 (N_411,In_367,In_696);
nor U412 (N_412,In_487,In_862);
nand U413 (N_413,In_647,In_689);
nand U414 (N_414,In_890,In_957);
and U415 (N_415,In_635,In_457);
and U416 (N_416,In_256,In_419);
and U417 (N_417,In_657,In_349);
or U418 (N_418,In_734,In_926);
nor U419 (N_419,In_135,In_137);
and U420 (N_420,In_791,In_342);
nand U421 (N_421,In_331,In_239);
or U422 (N_422,In_24,In_466);
nand U423 (N_423,In_494,In_563);
nor U424 (N_424,In_774,In_227);
and U425 (N_425,In_555,In_94);
nand U426 (N_426,In_499,In_623);
nor U427 (N_427,In_358,In_858);
or U428 (N_428,In_964,In_200);
or U429 (N_429,In_314,In_839);
nor U430 (N_430,In_418,In_475);
or U431 (N_431,In_253,In_513);
nor U432 (N_432,In_443,In_132);
nand U433 (N_433,In_73,In_214);
nand U434 (N_434,In_469,In_102);
and U435 (N_435,In_321,In_16);
and U436 (N_436,In_882,In_183);
or U437 (N_437,In_713,In_155);
and U438 (N_438,In_540,In_535);
or U439 (N_439,In_505,In_514);
and U440 (N_440,In_597,In_473);
and U441 (N_441,In_251,In_160);
nand U442 (N_442,In_745,In_161);
and U443 (N_443,In_340,In_181);
nor U444 (N_444,In_11,In_112);
and U445 (N_445,In_195,In_849);
nor U446 (N_446,In_572,In_444);
nor U447 (N_447,In_501,In_237);
nor U448 (N_448,In_204,In_971);
and U449 (N_449,In_977,In_762);
and U450 (N_450,In_533,In_14);
and U451 (N_451,In_17,In_854);
nand U452 (N_452,In_492,In_529);
and U453 (N_453,In_588,In_918);
nor U454 (N_454,In_233,In_192);
and U455 (N_455,In_298,In_470);
nand U456 (N_456,In_497,In_21);
and U457 (N_457,In_606,In_365);
and U458 (N_458,In_191,In_885);
nor U459 (N_459,In_72,In_709);
nand U460 (N_460,In_388,In_220);
nor U461 (N_461,In_577,In_693);
or U462 (N_462,In_553,In_628);
nand U463 (N_463,In_98,In_176);
and U464 (N_464,In_605,In_113);
and U465 (N_465,In_353,In_835);
nor U466 (N_466,In_576,In_78);
nor U467 (N_467,In_243,In_118);
nor U468 (N_468,In_26,In_295);
or U469 (N_469,In_464,In_47);
and U470 (N_470,In_177,In_642);
nand U471 (N_471,In_437,In_506);
nand U472 (N_472,In_639,In_71);
and U473 (N_473,In_316,In_42);
nor U474 (N_474,In_861,In_246);
or U475 (N_475,In_310,In_561);
nand U476 (N_476,In_565,In_133);
nor U477 (N_477,In_947,In_874);
nand U478 (N_478,In_244,In_509);
and U479 (N_479,In_158,In_838);
nand U480 (N_480,In_351,In_625);
nand U481 (N_481,In_414,In_127);
and U482 (N_482,In_123,In_121);
nand U483 (N_483,In_249,In_934);
nor U484 (N_484,In_41,In_653);
or U485 (N_485,In_68,In_922);
and U486 (N_486,In_269,In_790);
nand U487 (N_487,In_512,In_261);
or U488 (N_488,In_372,In_502);
or U489 (N_489,In_847,In_579);
nand U490 (N_490,In_618,In_814);
nor U491 (N_491,In_531,In_927);
nor U492 (N_492,In_585,In_570);
or U493 (N_493,In_948,In_784);
nor U494 (N_494,In_496,In_731);
nor U495 (N_495,In_980,In_976);
xnor U496 (N_496,In_970,In_973);
nand U497 (N_497,In_807,In_75);
and U498 (N_498,In_601,In_67);
nor U499 (N_499,In_850,In_972);
and U500 (N_500,In_5,In_661);
nand U501 (N_501,In_987,In_748);
or U502 (N_502,In_194,In_632);
or U503 (N_503,In_61,In_754);
or U504 (N_504,In_589,In_427);
nor U505 (N_505,In_732,In_507);
and U506 (N_506,In_810,In_270);
and U507 (N_507,In_544,In_371);
and U508 (N_508,In_45,In_385);
or U509 (N_509,In_796,In_195);
nor U510 (N_510,In_845,In_97);
nand U511 (N_511,In_95,In_712);
nor U512 (N_512,In_305,In_642);
nand U513 (N_513,In_649,In_545);
nor U514 (N_514,In_992,In_733);
and U515 (N_515,In_995,In_505);
or U516 (N_516,In_52,In_277);
and U517 (N_517,In_150,In_937);
nand U518 (N_518,In_472,In_285);
nor U519 (N_519,In_948,In_476);
or U520 (N_520,In_580,In_44);
and U521 (N_521,In_404,In_735);
and U522 (N_522,In_178,In_46);
and U523 (N_523,In_313,In_117);
or U524 (N_524,In_519,In_149);
and U525 (N_525,In_43,In_12);
nand U526 (N_526,In_644,In_660);
and U527 (N_527,In_406,In_394);
nor U528 (N_528,In_504,In_839);
or U529 (N_529,In_336,In_253);
and U530 (N_530,In_234,In_690);
xnor U531 (N_531,In_514,In_251);
or U532 (N_532,In_741,In_347);
nand U533 (N_533,In_913,In_164);
nor U534 (N_534,In_446,In_170);
nor U535 (N_535,In_699,In_521);
and U536 (N_536,In_250,In_137);
and U537 (N_537,In_429,In_364);
and U538 (N_538,In_879,In_470);
and U539 (N_539,In_216,In_421);
and U540 (N_540,In_110,In_209);
and U541 (N_541,In_616,In_926);
nand U542 (N_542,In_954,In_460);
nand U543 (N_543,In_636,In_434);
nand U544 (N_544,In_863,In_857);
and U545 (N_545,In_449,In_378);
nand U546 (N_546,In_260,In_518);
and U547 (N_547,In_800,In_119);
xor U548 (N_548,In_51,In_477);
nor U549 (N_549,In_406,In_590);
nor U550 (N_550,In_298,In_815);
and U551 (N_551,In_313,In_165);
and U552 (N_552,In_422,In_867);
or U553 (N_553,In_527,In_802);
nor U554 (N_554,In_231,In_19);
or U555 (N_555,In_640,In_466);
nor U556 (N_556,In_316,In_674);
and U557 (N_557,In_84,In_556);
nand U558 (N_558,In_355,In_462);
or U559 (N_559,In_887,In_655);
nor U560 (N_560,In_644,In_846);
nor U561 (N_561,In_934,In_217);
and U562 (N_562,In_731,In_622);
nand U563 (N_563,In_304,In_314);
or U564 (N_564,In_540,In_135);
or U565 (N_565,In_167,In_329);
or U566 (N_566,In_922,In_375);
nor U567 (N_567,In_749,In_739);
nor U568 (N_568,In_397,In_81);
or U569 (N_569,In_991,In_428);
nor U570 (N_570,In_59,In_353);
xor U571 (N_571,In_137,In_769);
nor U572 (N_572,In_336,In_179);
nand U573 (N_573,In_245,In_225);
nor U574 (N_574,In_661,In_442);
and U575 (N_575,In_857,In_970);
and U576 (N_576,In_534,In_428);
nand U577 (N_577,In_74,In_945);
and U578 (N_578,In_882,In_407);
and U579 (N_579,In_644,In_401);
nand U580 (N_580,In_960,In_625);
nand U581 (N_581,In_429,In_885);
nor U582 (N_582,In_170,In_70);
or U583 (N_583,In_56,In_271);
nand U584 (N_584,In_157,In_84);
nand U585 (N_585,In_533,In_672);
nand U586 (N_586,In_91,In_970);
or U587 (N_587,In_235,In_949);
nand U588 (N_588,In_594,In_230);
nor U589 (N_589,In_611,In_77);
or U590 (N_590,In_86,In_413);
and U591 (N_591,In_878,In_786);
and U592 (N_592,In_361,In_517);
nand U593 (N_593,In_132,In_431);
or U594 (N_594,In_448,In_940);
nand U595 (N_595,In_422,In_555);
and U596 (N_596,In_537,In_434);
and U597 (N_597,In_298,In_278);
or U598 (N_598,In_509,In_471);
nand U599 (N_599,In_430,In_198);
nor U600 (N_600,In_984,In_75);
or U601 (N_601,In_820,In_640);
nor U602 (N_602,In_324,In_614);
or U603 (N_603,In_618,In_232);
or U604 (N_604,In_816,In_457);
and U605 (N_605,In_135,In_565);
nand U606 (N_606,In_313,In_111);
and U607 (N_607,In_571,In_183);
or U608 (N_608,In_600,In_975);
or U609 (N_609,In_967,In_561);
or U610 (N_610,In_864,In_111);
nor U611 (N_611,In_105,In_226);
nand U612 (N_612,In_464,In_232);
or U613 (N_613,In_602,In_700);
nand U614 (N_614,In_935,In_30);
nor U615 (N_615,In_557,In_677);
or U616 (N_616,In_580,In_930);
and U617 (N_617,In_662,In_884);
and U618 (N_618,In_801,In_783);
nor U619 (N_619,In_383,In_905);
nor U620 (N_620,In_190,In_183);
and U621 (N_621,In_516,In_812);
nor U622 (N_622,In_233,In_600);
nand U623 (N_623,In_0,In_56);
nand U624 (N_624,In_544,In_332);
nor U625 (N_625,In_776,In_971);
or U626 (N_626,In_572,In_902);
nand U627 (N_627,In_448,In_648);
nor U628 (N_628,In_639,In_796);
nand U629 (N_629,In_791,In_365);
and U630 (N_630,In_492,In_506);
and U631 (N_631,In_945,In_660);
nand U632 (N_632,In_348,In_154);
nand U633 (N_633,In_830,In_529);
or U634 (N_634,In_438,In_35);
or U635 (N_635,In_643,In_909);
xor U636 (N_636,In_1,In_56);
and U637 (N_637,In_664,In_114);
nand U638 (N_638,In_4,In_492);
nand U639 (N_639,In_345,In_247);
xnor U640 (N_640,In_686,In_791);
or U641 (N_641,In_609,In_491);
nand U642 (N_642,In_871,In_505);
or U643 (N_643,In_578,In_495);
nor U644 (N_644,In_405,In_137);
nor U645 (N_645,In_481,In_439);
nand U646 (N_646,In_313,In_975);
nand U647 (N_647,In_736,In_342);
or U648 (N_648,In_162,In_863);
or U649 (N_649,In_91,In_268);
or U650 (N_650,In_113,In_537);
nand U651 (N_651,In_89,In_773);
nand U652 (N_652,In_41,In_697);
nand U653 (N_653,In_986,In_809);
nor U654 (N_654,In_471,In_44);
or U655 (N_655,In_215,In_198);
nor U656 (N_656,In_137,In_8);
nor U657 (N_657,In_735,In_980);
nand U658 (N_658,In_831,In_656);
nand U659 (N_659,In_215,In_262);
or U660 (N_660,In_375,In_728);
nand U661 (N_661,In_233,In_517);
nor U662 (N_662,In_480,In_266);
nor U663 (N_663,In_709,In_219);
and U664 (N_664,In_147,In_199);
nand U665 (N_665,In_273,In_275);
nor U666 (N_666,In_805,In_251);
nand U667 (N_667,In_783,In_503);
and U668 (N_668,In_574,In_4);
nand U669 (N_669,In_699,In_571);
nor U670 (N_670,In_211,In_87);
or U671 (N_671,In_124,In_230);
or U672 (N_672,In_702,In_167);
nor U673 (N_673,In_626,In_968);
or U674 (N_674,In_364,In_23);
or U675 (N_675,In_746,In_94);
or U676 (N_676,In_447,In_748);
nand U677 (N_677,In_692,In_570);
or U678 (N_678,In_467,In_414);
or U679 (N_679,In_471,In_968);
nor U680 (N_680,In_166,In_973);
nor U681 (N_681,In_241,In_824);
and U682 (N_682,In_584,In_786);
nand U683 (N_683,In_132,In_31);
nor U684 (N_684,In_571,In_408);
nor U685 (N_685,In_342,In_550);
or U686 (N_686,In_318,In_703);
nor U687 (N_687,In_993,In_597);
and U688 (N_688,In_16,In_758);
or U689 (N_689,In_275,In_996);
or U690 (N_690,In_989,In_918);
nand U691 (N_691,In_962,In_942);
or U692 (N_692,In_489,In_84);
nand U693 (N_693,In_349,In_925);
or U694 (N_694,In_211,In_509);
or U695 (N_695,In_727,In_690);
nor U696 (N_696,In_59,In_320);
nor U697 (N_697,In_176,In_328);
and U698 (N_698,In_598,In_116);
or U699 (N_699,In_753,In_166);
nand U700 (N_700,In_206,In_853);
nand U701 (N_701,In_556,In_386);
or U702 (N_702,In_794,In_537);
nor U703 (N_703,In_246,In_734);
and U704 (N_704,In_830,In_558);
or U705 (N_705,In_180,In_679);
or U706 (N_706,In_598,In_204);
or U707 (N_707,In_235,In_2);
or U708 (N_708,In_513,In_844);
nor U709 (N_709,In_55,In_675);
or U710 (N_710,In_207,In_773);
or U711 (N_711,In_177,In_874);
nand U712 (N_712,In_428,In_938);
nor U713 (N_713,In_34,In_156);
nand U714 (N_714,In_331,In_111);
and U715 (N_715,In_16,In_96);
nand U716 (N_716,In_614,In_600);
and U717 (N_717,In_987,In_787);
nor U718 (N_718,In_65,In_180);
nand U719 (N_719,In_269,In_296);
nand U720 (N_720,In_923,In_910);
nand U721 (N_721,In_995,In_713);
nand U722 (N_722,In_639,In_954);
or U723 (N_723,In_140,In_525);
nand U724 (N_724,In_684,In_412);
nand U725 (N_725,In_925,In_172);
or U726 (N_726,In_482,In_798);
and U727 (N_727,In_813,In_710);
or U728 (N_728,In_601,In_53);
and U729 (N_729,In_33,In_887);
nand U730 (N_730,In_581,In_281);
nor U731 (N_731,In_659,In_162);
nor U732 (N_732,In_700,In_746);
and U733 (N_733,In_0,In_224);
nand U734 (N_734,In_911,In_621);
nor U735 (N_735,In_381,In_932);
nor U736 (N_736,In_15,In_813);
or U737 (N_737,In_458,In_246);
nand U738 (N_738,In_921,In_263);
nor U739 (N_739,In_428,In_970);
nand U740 (N_740,In_807,In_162);
nor U741 (N_741,In_39,In_198);
or U742 (N_742,In_578,In_151);
nand U743 (N_743,In_329,In_225);
and U744 (N_744,In_526,In_235);
nor U745 (N_745,In_628,In_720);
or U746 (N_746,In_33,In_885);
nand U747 (N_747,In_505,In_42);
xor U748 (N_748,In_466,In_952);
nand U749 (N_749,In_820,In_551);
nand U750 (N_750,In_508,In_729);
or U751 (N_751,In_85,In_962);
nor U752 (N_752,In_592,In_854);
nand U753 (N_753,In_559,In_898);
nand U754 (N_754,In_772,In_142);
nand U755 (N_755,In_28,In_903);
nand U756 (N_756,In_195,In_529);
nand U757 (N_757,In_403,In_507);
or U758 (N_758,In_619,In_26);
or U759 (N_759,In_627,In_755);
nor U760 (N_760,In_959,In_104);
nand U761 (N_761,In_677,In_684);
nor U762 (N_762,In_816,In_902);
nor U763 (N_763,In_797,In_437);
and U764 (N_764,In_915,In_222);
nor U765 (N_765,In_965,In_499);
nand U766 (N_766,In_90,In_167);
nor U767 (N_767,In_788,In_896);
nand U768 (N_768,In_455,In_719);
nor U769 (N_769,In_166,In_926);
nand U770 (N_770,In_778,In_770);
or U771 (N_771,In_355,In_469);
nor U772 (N_772,In_639,In_15);
and U773 (N_773,In_531,In_273);
and U774 (N_774,In_172,In_439);
nor U775 (N_775,In_721,In_662);
and U776 (N_776,In_890,In_410);
nor U777 (N_777,In_615,In_127);
nand U778 (N_778,In_493,In_771);
nor U779 (N_779,In_950,In_10);
nor U780 (N_780,In_773,In_818);
nor U781 (N_781,In_859,In_409);
xnor U782 (N_782,In_541,In_490);
or U783 (N_783,In_54,In_923);
nand U784 (N_784,In_478,In_874);
nor U785 (N_785,In_310,In_136);
and U786 (N_786,In_335,In_474);
nand U787 (N_787,In_487,In_872);
nand U788 (N_788,In_395,In_10);
nor U789 (N_789,In_279,In_955);
nand U790 (N_790,In_928,In_579);
nor U791 (N_791,In_866,In_689);
and U792 (N_792,In_35,In_746);
nor U793 (N_793,In_470,In_446);
xnor U794 (N_794,In_932,In_808);
nor U795 (N_795,In_872,In_990);
or U796 (N_796,In_683,In_861);
and U797 (N_797,In_386,In_841);
and U798 (N_798,In_259,In_940);
nor U799 (N_799,In_832,In_930);
and U800 (N_800,In_568,In_777);
and U801 (N_801,In_252,In_740);
nand U802 (N_802,In_74,In_279);
nor U803 (N_803,In_813,In_324);
or U804 (N_804,In_141,In_194);
or U805 (N_805,In_196,In_402);
and U806 (N_806,In_377,In_895);
nor U807 (N_807,In_599,In_386);
or U808 (N_808,In_506,In_391);
and U809 (N_809,In_20,In_859);
or U810 (N_810,In_588,In_422);
nor U811 (N_811,In_154,In_51);
and U812 (N_812,In_213,In_535);
nor U813 (N_813,In_748,In_844);
nor U814 (N_814,In_204,In_365);
nor U815 (N_815,In_411,In_51);
nand U816 (N_816,In_178,In_885);
or U817 (N_817,In_877,In_559);
nor U818 (N_818,In_97,In_917);
and U819 (N_819,In_502,In_283);
and U820 (N_820,In_755,In_569);
or U821 (N_821,In_254,In_469);
and U822 (N_822,In_788,In_204);
or U823 (N_823,In_789,In_783);
and U824 (N_824,In_984,In_575);
nor U825 (N_825,In_821,In_449);
or U826 (N_826,In_192,In_433);
or U827 (N_827,In_686,In_250);
or U828 (N_828,In_80,In_899);
or U829 (N_829,In_419,In_682);
and U830 (N_830,In_399,In_248);
nor U831 (N_831,In_708,In_234);
and U832 (N_832,In_618,In_162);
nand U833 (N_833,In_869,In_280);
and U834 (N_834,In_999,In_651);
or U835 (N_835,In_480,In_471);
and U836 (N_836,In_111,In_896);
or U837 (N_837,In_242,In_937);
nand U838 (N_838,In_50,In_844);
and U839 (N_839,In_543,In_669);
nand U840 (N_840,In_740,In_500);
nand U841 (N_841,In_473,In_11);
nand U842 (N_842,In_141,In_839);
xor U843 (N_843,In_326,In_819);
and U844 (N_844,In_701,In_154);
nand U845 (N_845,In_825,In_413);
and U846 (N_846,In_975,In_696);
or U847 (N_847,In_386,In_557);
and U848 (N_848,In_868,In_805);
nand U849 (N_849,In_475,In_235);
nor U850 (N_850,In_899,In_545);
and U851 (N_851,In_347,In_722);
and U852 (N_852,In_370,In_442);
or U853 (N_853,In_144,In_73);
nand U854 (N_854,In_350,In_671);
or U855 (N_855,In_92,In_822);
and U856 (N_856,In_797,In_58);
nor U857 (N_857,In_476,In_608);
nor U858 (N_858,In_109,In_416);
or U859 (N_859,In_335,In_458);
xnor U860 (N_860,In_595,In_452);
nand U861 (N_861,In_451,In_585);
or U862 (N_862,In_773,In_742);
nand U863 (N_863,In_752,In_179);
nor U864 (N_864,In_283,In_914);
or U865 (N_865,In_204,In_250);
nand U866 (N_866,In_169,In_48);
and U867 (N_867,In_268,In_211);
and U868 (N_868,In_685,In_356);
and U869 (N_869,In_410,In_736);
and U870 (N_870,In_336,In_441);
or U871 (N_871,In_411,In_400);
and U872 (N_872,In_93,In_761);
nand U873 (N_873,In_10,In_456);
nor U874 (N_874,In_187,In_802);
or U875 (N_875,In_548,In_659);
or U876 (N_876,In_568,In_590);
and U877 (N_877,In_760,In_826);
and U878 (N_878,In_496,In_774);
nor U879 (N_879,In_589,In_528);
nor U880 (N_880,In_648,In_296);
or U881 (N_881,In_135,In_304);
nand U882 (N_882,In_265,In_545);
or U883 (N_883,In_840,In_94);
nor U884 (N_884,In_358,In_13);
xnor U885 (N_885,In_463,In_864);
nand U886 (N_886,In_503,In_293);
and U887 (N_887,In_403,In_481);
or U888 (N_888,In_359,In_360);
and U889 (N_889,In_124,In_212);
and U890 (N_890,In_989,In_866);
nand U891 (N_891,In_969,In_308);
nor U892 (N_892,In_358,In_58);
and U893 (N_893,In_419,In_468);
and U894 (N_894,In_940,In_559);
nor U895 (N_895,In_997,In_963);
and U896 (N_896,In_67,In_269);
and U897 (N_897,In_567,In_997);
or U898 (N_898,In_522,In_883);
nor U899 (N_899,In_459,In_185);
nor U900 (N_900,In_929,In_866);
and U901 (N_901,In_441,In_655);
or U902 (N_902,In_467,In_979);
and U903 (N_903,In_701,In_849);
nor U904 (N_904,In_744,In_376);
nor U905 (N_905,In_810,In_844);
and U906 (N_906,In_918,In_561);
nand U907 (N_907,In_199,In_382);
and U908 (N_908,In_644,In_456);
or U909 (N_909,In_682,In_189);
or U910 (N_910,In_220,In_569);
nand U911 (N_911,In_283,In_713);
nor U912 (N_912,In_436,In_502);
nand U913 (N_913,In_299,In_480);
and U914 (N_914,In_644,In_541);
and U915 (N_915,In_502,In_653);
nor U916 (N_916,In_797,In_945);
or U917 (N_917,In_580,In_690);
or U918 (N_918,In_760,In_827);
nand U919 (N_919,In_519,In_684);
nand U920 (N_920,In_652,In_335);
nor U921 (N_921,In_922,In_494);
or U922 (N_922,In_258,In_233);
and U923 (N_923,In_746,In_105);
nor U924 (N_924,In_85,In_472);
nor U925 (N_925,In_518,In_95);
nor U926 (N_926,In_931,In_608);
nor U927 (N_927,In_138,In_84);
or U928 (N_928,In_927,In_864);
and U929 (N_929,In_249,In_435);
and U930 (N_930,In_349,In_394);
and U931 (N_931,In_221,In_932);
or U932 (N_932,In_428,In_646);
xnor U933 (N_933,In_36,In_858);
or U934 (N_934,In_803,In_874);
nand U935 (N_935,In_656,In_492);
and U936 (N_936,In_15,In_704);
nand U937 (N_937,In_188,In_311);
or U938 (N_938,In_843,In_175);
nor U939 (N_939,In_360,In_407);
and U940 (N_940,In_565,In_371);
nand U941 (N_941,In_44,In_78);
nand U942 (N_942,In_814,In_437);
or U943 (N_943,In_943,In_322);
and U944 (N_944,In_16,In_119);
or U945 (N_945,In_0,In_327);
nor U946 (N_946,In_364,In_223);
or U947 (N_947,In_111,In_126);
xnor U948 (N_948,In_467,In_524);
nor U949 (N_949,In_112,In_14);
nor U950 (N_950,In_548,In_833);
and U951 (N_951,In_301,In_817);
xnor U952 (N_952,In_818,In_295);
and U953 (N_953,In_838,In_634);
nor U954 (N_954,In_493,In_768);
nand U955 (N_955,In_809,In_44);
nand U956 (N_956,In_360,In_481);
or U957 (N_957,In_644,In_983);
and U958 (N_958,In_173,In_381);
and U959 (N_959,In_727,In_183);
or U960 (N_960,In_283,In_490);
nor U961 (N_961,In_402,In_575);
or U962 (N_962,In_12,In_620);
nand U963 (N_963,In_971,In_602);
and U964 (N_964,In_481,In_28);
nor U965 (N_965,In_815,In_273);
and U966 (N_966,In_836,In_541);
or U967 (N_967,In_67,In_70);
nor U968 (N_968,In_142,In_135);
or U969 (N_969,In_816,In_580);
or U970 (N_970,In_122,In_378);
and U971 (N_971,In_537,In_206);
and U972 (N_972,In_367,In_276);
or U973 (N_973,In_2,In_850);
or U974 (N_974,In_499,In_1);
nor U975 (N_975,In_355,In_544);
or U976 (N_976,In_276,In_464);
xor U977 (N_977,In_281,In_702);
nor U978 (N_978,In_300,In_180);
nor U979 (N_979,In_425,In_46);
nor U980 (N_980,In_169,In_877);
nand U981 (N_981,In_473,In_435);
and U982 (N_982,In_859,In_730);
or U983 (N_983,In_116,In_733);
or U984 (N_984,In_734,In_600);
and U985 (N_985,In_550,In_875);
and U986 (N_986,In_459,In_246);
nor U987 (N_987,In_539,In_556);
nor U988 (N_988,In_0,In_759);
nor U989 (N_989,In_978,In_947);
nand U990 (N_990,In_162,In_534);
nor U991 (N_991,In_373,In_576);
nand U992 (N_992,In_632,In_727);
nor U993 (N_993,In_180,In_115);
nand U994 (N_994,In_654,In_134);
or U995 (N_995,In_471,In_536);
and U996 (N_996,In_229,In_687);
nand U997 (N_997,In_687,In_302);
and U998 (N_998,In_253,In_938);
and U999 (N_999,In_932,In_740);
nor U1000 (N_1000,In_87,In_91);
or U1001 (N_1001,In_42,In_476);
nand U1002 (N_1002,In_91,In_807);
nor U1003 (N_1003,In_504,In_248);
nand U1004 (N_1004,In_196,In_2);
and U1005 (N_1005,In_213,In_567);
and U1006 (N_1006,In_590,In_663);
nor U1007 (N_1007,In_412,In_876);
and U1008 (N_1008,In_395,In_797);
nand U1009 (N_1009,In_902,In_508);
or U1010 (N_1010,In_903,In_599);
nand U1011 (N_1011,In_781,In_648);
or U1012 (N_1012,In_983,In_694);
or U1013 (N_1013,In_848,In_409);
nor U1014 (N_1014,In_938,In_608);
nand U1015 (N_1015,In_982,In_839);
and U1016 (N_1016,In_641,In_401);
nor U1017 (N_1017,In_768,In_390);
nor U1018 (N_1018,In_897,In_994);
nand U1019 (N_1019,In_515,In_189);
and U1020 (N_1020,In_791,In_751);
or U1021 (N_1021,In_971,In_126);
and U1022 (N_1022,In_816,In_712);
or U1023 (N_1023,In_899,In_482);
nand U1024 (N_1024,In_292,In_399);
nor U1025 (N_1025,In_511,In_132);
or U1026 (N_1026,In_705,In_289);
nand U1027 (N_1027,In_189,In_233);
and U1028 (N_1028,In_409,In_361);
or U1029 (N_1029,In_233,In_898);
nand U1030 (N_1030,In_234,In_243);
nor U1031 (N_1031,In_367,In_171);
nor U1032 (N_1032,In_305,In_928);
nor U1033 (N_1033,In_76,In_555);
and U1034 (N_1034,In_92,In_982);
nor U1035 (N_1035,In_201,In_886);
nand U1036 (N_1036,In_377,In_267);
nand U1037 (N_1037,In_320,In_544);
nand U1038 (N_1038,In_317,In_273);
or U1039 (N_1039,In_247,In_33);
and U1040 (N_1040,In_288,In_856);
nand U1041 (N_1041,In_919,In_731);
nand U1042 (N_1042,In_374,In_125);
and U1043 (N_1043,In_433,In_859);
or U1044 (N_1044,In_197,In_896);
nand U1045 (N_1045,In_955,In_642);
nor U1046 (N_1046,In_227,In_915);
and U1047 (N_1047,In_400,In_441);
or U1048 (N_1048,In_199,In_82);
nand U1049 (N_1049,In_80,In_907);
or U1050 (N_1050,In_210,In_220);
or U1051 (N_1051,In_885,In_507);
and U1052 (N_1052,In_230,In_665);
nand U1053 (N_1053,In_809,In_259);
nor U1054 (N_1054,In_940,In_262);
and U1055 (N_1055,In_891,In_999);
nand U1056 (N_1056,In_881,In_363);
or U1057 (N_1057,In_415,In_199);
and U1058 (N_1058,In_163,In_278);
and U1059 (N_1059,In_999,In_5);
nor U1060 (N_1060,In_759,In_405);
nand U1061 (N_1061,In_780,In_499);
nand U1062 (N_1062,In_37,In_983);
nor U1063 (N_1063,In_65,In_970);
or U1064 (N_1064,In_183,In_734);
nor U1065 (N_1065,In_477,In_3);
or U1066 (N_1066,In_886,In_383);
and U1067 (N_1067,In_681,In_393);
or U1068 (N_1068,In_510,In_990);
nor U1069 (N_1069,In_41,In_403);
nor U1070 (N_1070,In_55,In_635);
nand U1071 (N_1071,In_633,In_989);
or U1072 (N_1072,In_710,In_301);
nand U1073 (N_1073,In_473,In_717);
and U1074 (N_1074,In_305,In_933);
and U1075 (N_1075,In_225,In_977);
nor U1076 (N_1076,In_585,In_576);
nand U1077 (N_1077,In_618,In_904);
xnor U1078 (N_1078,In_664,In_30);
or U1079 (N_1079,In_152,In_920);
or U1080 (N_1080,In_686,In_42);
nor U1081 (N_1081,In_593,In_918);
and U1082 (N_1082,In_370,In_884);
nand U1083 (N_1083,In_320,In_619);
nand U1084 (N_1084,In_800,In_754);
or U1085 (N_1085,In_312,In_948);
or U1086 (N_1086,In_878,In_423);
nand U1087 (N_1087,In_372,In_706);
and U1088 (N_1088,In_537,In_358);
nand U1089 (N_1089,In_494,In_400);
or U1090 (N_1090,In_403,In_905);
nand U1091 (N_1091,In_46,In_583);
nor U1092 (N_1092,In_14,In_521);
or U1093 (N_1093,In_166,In_633);
or U1094 (N_1094,In_179,In_921);
nand U1095 (N_1095,In_688,In_483);
nor U1096 (N_1096,In_639,In_806);
and U1097 (N_1097,In_26,In_419);
or U1098 (N_1098,In_374,In_741);
and U1099 (N_1099,In_949,In_428);
nand U1100 (N_1100,In_697,In_546);
or U1101 (N_1101,In_903,In_630);
nor U1102 (N_1102,In_251,In_434);
and U1103 (N_1103,In_623,In_824);
nand U1104 (N_1104,In_248,In_978);
and U1105 (N_1105,In_277,In_481);
and U1106 (N_1106,In_667,In_167);
nand U1107 (N_1107,In_812,In_84);
or U1108 (N_1108,In_473,In_808);
nand U1109 (N_1109,In_810,In_465);
nor U1110 (N_1110,In_270,In_422);
or U1111 (N_1111,In_850,In_738);
nor U1112 (N_1112,In_398,In_860);
nor U1113 (N_1113,In_784,In_329);
and U1114 (N_1114,In_670,In_436);
nand U1115 (N_1115,In_318,In_316);
or U1116 (N_1116,In_774,In_71);
nor U1117 (N_1117,In_361,In_681);
nand U1118 (N_1118,In_928,In_300);
and U1119 (N_1119,In_752,In_766);
nand U1120 (N_1120,In_902,In_909);
nand U1121 (N_1121,In_57,In_990);
nor U1122 (N_1122,In_612,In_249);
and U1123 (N_1123,In_989,In_449);
or U1124 (N_1124,In_88,In_508);
nor U1125 (N_1125,In_672,In_112);
nor U1126 (N_1126,In_781,In_636);
or U1127 (N_1127,In_753,In_68);
nand U1128 (N_1128,In_484,In_672);
and U1129 (N_1129,In_43,In_445);
and U1130 (N_1130,In_96,In_724);
nand U1131 (N_1131,In_988,In_869);
nor U1132 (N_1132,In_906,In_884);
nor U1133 (N_1133,In_806,In_613);
and U1134 (N_1134,In_656,In_197);
and U1135 (N_1135,In_34,In_53);
and U1136 (N_1136,In_25,In_640);
nand U1137 (N_1137,In_22,In_163);
nand U1138 (N_1138,In_206,In_745);
or U1139 (N_1139,In_876,In_620);
or U1140 (N_1140,In_815,In_35);
nand U1141 (N_1141,In_232,In_18);
or U1142 (N_1142,In_648,In_222);
or U1143 (N_1143,In_792,In_441);
and U1144 (N_1144,In_637,In_911);
nand U1145 (N_1145,In_658,In_866);
or U1146 (N_1146,In_835,In_329);
nand U1147 (N_1147,In_811,In_780);
or U1148 (N_1148,In_343,In_362);
nor U1149 (N_1149,In_845,In_738);
nand U1150 (N_1150,In_686,In_5);
nor U1151 (N_1151,In_284,In_817);
or U1152 (N_1152,In_402,In_121);
or U1153 (N_1153,In_199,In_422);
or U1154 (N_1154,In_681,In_869);
or U1155 (N_1155,In_164,In_270);
nand U1156 (N_1156,In_545,In_764);
and U1157 (N_1157,In_705,In_326);
or U1158 (N_1158,In_6,In_104);
or U1159 (N_1159,In_890,In_985);
nand U1160 (N_1160,In_828,In_935);
and U1161 (N_1161,In_35,In_46);
nor U1162 (N_1162,In_879,In_954);
nor U1163 (N_1163,In_929,In_217);
nand U1164 (N_1164,In_284,In_219);
or U1165 (N_1165,In_42,In_589);
or U1166 (N_1166,In_488,In_65);
nand U1167 (N_1167,In_514,In_389);
nand U1168 (N_1168,In_71,In_172);
or U1169 (N_1169,In_878,In_559);
or U1170 (N_1170,In_601,In_763);
or U1171 (N_1171,In_473,In_49);
nand U1172 (N_1172,In_882,In_903);
nor U1173 (N_1173,In_735,In_522);
or U1174 (N_1174,In_862,In_764);
and U1175 (N_1175,In_333,In_33);
nand U1176 (N_1176,In_191,In_329);
nor U1177 (N_1177,In_568,In_332);
nand U1178 (N_1178,In_954,In_477);
nand U1179 (N_1179,In_332,In_540);
nand U1180 (N_1180,In_664,In_766);
and U1181 (N_1181,In_451,In_765);
nor U1182 (N_1182,In_397,In_444);
and U1183 (N_1183,In_662,In_278);
and U1184 (N_1184,In_422,In_966);
or U1185 (N_1185,In_52,In_986);
and U1186 (N_1186,In_315,In_154);
nand U1187 (N_1187,In_604,In_180);
or U1188 (N_1188,In_312,In_249);
nand U1189 (N_1189,In_317,In_415);
nor U1190 (N_1190,In_575,In_969);
nor U1191 (N_1191,In_957,In_279);
or U1192 (N_1192,In_642,In_859);
or U1193 (N_1193,In_868,In_722);
or U1194 (N_1194,In_689,In_914);
and U1195 (N_1195,In_908,In_415);
or U1196 (N_1196,In_674,In_996);
nand U1197 (N_1197,In_834,In_442);
xor U1198 (N_1198,In_940,In_863);
nand U1199 (N_1199,In_372,In_310);
nor U1200 (N_1200,In_149,In_361);
nor U1201 (N_1201,In_615,In_311);
and U1202 (N_1202,In_787,In_208);
or U1203 (N_1203,In_471,In_586);
nand U1204 (N_1204,In_294,In_848);
or U1205 (N_1205,In_276,In_935);
nor U1206 (N_1206,In_466,In_909);
or U1207 (N_1207,In_857,In_589);
and U1208 (N_1208,In_13,In_319);
and U1209 (N_1209,In_656,In_916);
nand U1210 (N_1210,In_624,In_991);
or U1211 (N_1211,In_142,In_332);
nand U1212 (N_1212,In_369,In_268);
and U1213 (N_1213,In_239,In_55);
and U1214 (N_1214,In_193,In_964);
nand U1215 (N_1215,In_458,In_111);
and U1216 (N_1216,In_321,In_86);
or U1217 (N_1217,In_218,In_78);
nand U1218 (N_1218,In_250,In_492);
or U1219 (N_1219,In_294,In_973);
nor U1220 (N_1220,In_287,In_401);
or U1221 (N_1221,In_840,In_101);
or U1222 (N_1222,In_111,In_983);
nor U1223 (N_1223,In_477,In_682);
and U1224 (N_1224,In_668,In_221);
or U1225 (N_1225,In_280,In_27);
nor U1226 (N_1226,In_665,In_714);
and U1227 (N_1227,In_643,In_252);
and U1228 (N_1228,In_257,In_997);
nor U1229 (N_1229,In_777,In_566);
or U1230 (N_1230,In_379,In_314);
nor U1231 (N_1231,In_480,In_461);
or U1232 (N_1232,In_358,In_595);
or U1233 (N_1233,In_196,In_578);
or U1234 (N_1234,In_54,In_378);
and U1235 (N_1235,In_150,In_870);
and U1236 (N_1236,In_51,In_94);
nand U1237 (N_1237,In_137,In_581);
nor U1238 (N_1238,In_475,In_367);
or U1239 (N_1239,In_588,In_178);
and U1240 (N_1240,In_298,In_623);
and U1241 (N_1241,In_235,In_924);
and U1242 (N_1242,In_579,In_919);
and U1243 (N_1243,In_516,In_745);
nor U1244 (N_1244,In_858,In_182);
nor U1245 (N_1245,In_972,In_469);
nand U1246 (N_1246,In_899,In_194);
and U1247 (N_1247,In_265,In_262);
nor U1248 (N_1248,In_550,In_299);
and U1249 (N_1249,In_160,In_854);
nand U1250 (N_1250,In_0,In_185);
and U1251 (N_1251,In_393,In_288);
nand U1252 (N_1252,In_23,In_262);
nor U1253 (N_1253,In_278,In_447);
nor U1254 (N_1254,In_250,In_266);
or U1255 (N_1255,In_694,In_1);
nor U1256 (N_1256,In_829,In_89);
nand U1257 (N_1257,In_449,In_531);
nor U1258 (N_1258,In_48,In_135);
or U1259 (N_1259,In_202,In_54);
nand U1260 (N_1260,In_602,In_519);
or U1261 (N_1261,In_355,In_707);
or U1262 (N_1262,In_173,In_12);
or U1263 (N_1263,In_588,In_536);
nor U1264 (N_1264,In_931,In_828);
nor U1265 (N_1265,In_926,In_119);
or U1266 (N_1266,In_172,In_990);
nand U1267 (N_1267,In_324,In_858);
nand U1268 (N_1268,In_374,In_26);
nand U1269 (N_1269,In_933,In_751);
or U1270 (N_1270,In_115,In_565);
or U1271 (N_1271,In_23,In_777);
nand U1272 (N_1272,In_453,In_409);
or U1273 (N_1273,In_982,In_860);
nand U1274 (N_1274,In_697,In_366);
xnor U1275 (N_1275,In_213,In_693);
and U1276 (N_1276,In_85,In_591);
and U1277 (N_1277,In_445,In_631);
nand U1278 (N_1278,In_142,In_148);
nand U1279 (N_1279,In_282,In_833);
nand U1280 (N_1280,In_33,In_886);
nor U1281 (N_1281,In_33,In_839);
or U1282 (N_1282,In_354,In_538);
nand U1283 (N_1283,In_11,In_216);
and U1284 (N_1284,In_178,In_667);
or U1285 (N_1285,In_989,In_254);
nor U1286 (N_1286,In_689,In_633);
or U1287 (N_1287,In_604,In_98);
nand U1288 (N_1288,In_995,In_411);
or U1289 (N_1289,In_562,In_713);
nor U1290 (N_1290,In_436,In_296);
or U1291 (N_1291,In_744,In_801);
nand U1292 (N_1292,In_951,In_166);
nand U1293 (N_1293,In_756,In_434);
nor U1294 (N_1294,In_481,In_727);
or U1295 (N_1295,In_217,In_287);
and U1296 (N_1296,In_509,In_373);
and U1297 (N_1297,In_945,In_975);
or U1298 (N_1298,In_468,In_188);
or U1299 (N_1299,In_703,In_189);
or U1300 (N_1300,In_200,In_191);
nand U1301 (N_1301,In_293,In_63);
or U1302 (N_1302,In_168,In_9);
and U1303 (N_1303,In_9,In_760);
nand U1304 (N_1304,In_298,In_496);
and U1305 (N_1305,In_835,In_438);
or U1306 (N_1306,In_730,In_114);
or U1307 (N_1307,In_383,In_290);
or U1308 (N_1308,In_720,In_585);
nor U1309 (N_1309,In_692,In_306);
and U1310 (N_1310,In_55,In_874);
nor U1311 (N_1311,In_152,In_314);
nor U1312 (N_1312,In_841,In_413);
nor U1313 (N_1313,In_304,In_779);
or U1314 (N_1314,In_835,In_174);
nand U1315 (N_1315,In_162,In_580);
or U1316 (N_1316,In_935,In_752);
nand U1317 (N_1317,In_473,In_448);
and U1318 (N_1318,In_493,In_40);
nand U1319 (N_1319,In_331,In_81);
or U1320 (N_1320,In_625,In_832);
nor U1321 (N_1321,In_863,In_366);
nand U1322 (N_1322,In_876,In_117);
or U1323 (N_1323,In_247,In_642);
and U1324 (N_1324,In_181,In_830);
nor U1325 (N_1325,In_507,In_212);
or U1326 (N_1326,In_776,In_270);
nor U1327 (N_1327,In_143,In_357);
nor U1328 (N_1328,In_994,In_416);
and U1329 (N_1329,In_140,In_238);
or U1330 (N_1330,In_44,In_664);
or U1331 (N_1331,In_737,In_437);
and U1332 (N_1332,In_12,In_192);
nand U1333 (N_1333,In_547,In_74);
or U1334 (N_1334,In_848,In_618);
nor U1335 (N_1335,In_128,In_957);
nor U1336 (N_1336,In_546,In_75);
and U1337 (N_1337,In_842,In_565);
and U1338 (N_1338,In_391,In_858);
nor U1339 (N_1339,In_8,In_324);
nor U1340 (N_1340,In_818,In_466);
nand U1341 (N_1341,In_588,In_255);
or U1342 (N_1342,In_963,In_877);
nor U1343 (N_1343,In_100,In_845);
nand U1344 (N_1344,In_916,In_300);
or U1345 (N_1345,In_902,In_0);
nor U1346 (N_1346,In_265,In_505);
nand U1347 (N_1347,In_792,In_543);
and U1348 (N_1348,In_845,In_446);
nand U1349 (N_1349,In_266,In_740);
nand U1350 (N_1350,In_464,In_162);
nor U1351 (N_1351,In_401,In_964);
nor U1352 (N_1352,In_212,In_615);
and U1353 (N_1353,In_296,In_92);
nor U1354 (N_1354,In_936,In_859);
and U1355 (N_1355,In_378,In_139);
nor U1356 (N_1356,In_756,In_961);
nor U1357 (N_1357,In_276,In_356);
and U1358 (N_1358,In_376,In_240);
nor U1359 (N_1359,In_818,In_378);
nand U1360 (N_1360,In_24,In_309);
or U1361 (N_1361,In_294,In_161);
and U1362 (N_1362,In_242,In_909);
nand U1363 (N_1363,In_130,In_105);
or U1364 (N_1364,In_543,In_811);
nor U1365 (N_1365,In_812,In_471);
nand U1366 (N_1366,In_106,In_436);
and U1367 (N_1367,In_226,In_48);
and U1368 (N_1368,In_870,In_34);
or U1369 (N_1369,In_513,In_489);
and U1370 (N_1370,In_817,In_848);
and U1371 (N_1371,In_445,In_184);
and U1372 (N_1372,In_952,In_461);
or U1373 (N_1373,In_363,In_908);
and U1374 (N_1374,In_224,In_571);
nand U1375 (N_1375,In_484,In_532);
nand U1376 (N_1376,In_148,In_127);
nor U1377 (N_1377,In_278,In_139);
or U1378 (N_1378,In_509,In_637);
or U1379 (N_1379,In_672,In_396);
nand U1380 (N_1380,In_147,In_59);
xor U1381 (N_1381,In_225,In_389);
nand U1382 (N_1382,In_893,In_729);
or U1383 (N_1383,In_509,In_31);
or U1384 (N_1384,In_611,In_61);
nor U1385 (N_1385,In_644,In_759);
nand U1386 (N_1386,In_718,In_532);
nor U1387 (N_1387,In_535,In_852);
and U1388 (N_1388,In_380,In_368);
nor U1389 (N_1389,In_825,In_954);
or U1390 (N_1390,In_843,In_624);
nor U1391 (N_1391,In_423,In_967);
nand U1392 (N_1392,In_368,In_395);
or U1393 (N_1393,In_310,In_662);
nor U1394 (N_1394,In_321,In_936);
nor U1395 (N_1395,In_448,In_881);
nor U1396 (N_1396,In_970,In_958);
nor U1397 (N_1397,In_787,In_957);
or U1398 (N_1398,In_458,In_830);
or U1399 (N_1399,In_864,In_609);
and U1400 (N_1400,In_81,In_909);
nand U1401 (N_1401,In_868,In_301);
or U1402 (N_1402,In_528,In_836);
or U1403 (N_1403,In_735,In_771);
nor U1404 (N_1404,In_338,In_523);
nor U1405 (N_1405,In_895,In_758);
or U1406 (N_1406,In_937,In_49);
nor U1407 (N_1407,In_535,In_224);
and U1408 (N_1408,In_836,In_745);
nor U1409 (N_1409,In_675,In_810);
nor U1410 (N_1410,In_454,In_100);
and U1411 (N_1411,In_474,In_73);
or U1412 (N_1412,In_271,In_136);
and U1413 (N_1413,In_810,In_240);
nor U1414 (N_1414,In_664,In_502);
nor U1415 (N_1415,In_481,In_637);
nor U1416 (N_1416,In_123,In_189);
or U1417 (N_1417,In_560,In_348);
nand U1418 (N_1418,In_973,In_269);
or U1419 (N_1419,In_425,In_873);
nor U1420 (N_1420,In_66,In_27);
nor U1421 (N_1421,In_235,In_896);
nand U1422 (N_1422,In_953,In_102);
nor U1423 (N_1423,In_531,In_888);
and U1424 (N_1424,In_695,In_535);
and U1425 (N_1425,In_856,In_587);
nand U1426 (N_1426,In_996,In_510);
nor U1427 (N_1427,In_54,In_551);
or U1428 (N_1428,In_736,In_54);
and U1429 (N_1429,In_95,In_257);
nand U1430 (N_1430,In_498,In_468);
or U1431 (N_1431,In_414,In_478);
or U1432 (N_1432,In_670,In_308);
and U1433 (N_1433,In_635,In_927);
or U1434 (N_1434,In_124,In_513);
and U1435 (N_1435,In_689,In_218);
or U1436 (N_1436,In_855,In_325);
and U1437 (N_1437,In_350,In_287);
nand U1438 (N_1438,In_302,In_546);
nand U1439 (N_1439,In_445,In_809);
nand U1440 (N_1440,In_668,In_477);
nand U1441 (N_1441,In_973,In_506);
or U1442 (N_1442,In_210,In_549);
nor U1443 (N_1443,In_901,In_764);
nand U1444 (N_1444,In_815,In_698);
or U1445 (N_1445,In_77,In_691);
nand U1446 (N_1446,In_464,In_312);
nor U1447 (N_1447,In_664,In_900);
or U1448 (N_1448,In_130,In_275);
and U1449 (N_1449,In_217,In_648);
or U1450 (N_1450,In_742,In_652);
and U1451 (N_1451,In_250,In_409);
and U1452 (N_1452,In_788,In_201);
nor U1453 (N_1453,In_157,In_112);
and U1454 (N_1454,In_830,In_204);
nor U1455 (N_1455,In_87,In_272);
and U1456 (N_1456,In_487,In_903);
or U1457 (N_1457,In_558,In_192);
or U1458 (N_1458,In_265,In_510);
and U1459 (N_1459,In_72,In_917);
xor U1460 (N_1460,In_832,In_384);
nand U1461 (N_1461,In_84,In_737);
nor U1462 (N_1462,In_333,In_747);
and U1463 (N_1463,In_269,In_314);
nor U1464 (N_1464,In_944,In_259);
and U1465 (N_1465,In_671,In_53);
and U1466 (N_1466,In_221,In_734);
and U1467 (N_1467,In_64,In_270);
or U1468 (N_1468,In_532,In_264);
nor U1469 (N_1469,In_565,In_287);
and U1470 (N_1470,In_477,In_359);
or U1471 (N_1471,In_939,In_407);
nand U1472 (N_1472,In_41,In_13);
nand U1473 (N_1473,In_539,In_998);
nand U1474 (N_1474,In_93,In_649);
nand U1475 (N_1475,In_454,In_475);
nand U1476 (N_1476,In_212,In_501);
nor U1477 (N_1477,In_128,In_433);
nand U1478 (N_1478,In_161,In_124);
nor U1479 (N_1479,In_576,In_687);
nand U1480 (N_1480,In_535,In_827);
and U1481 (N_1481,In_105,In_377);
nor U1482 (N_1482,In_930,In_762);
nor U1483 (N_1483,In_377,In_885);
nand U1484 (N_1484,In_640,In_200);
and U1485 (N_1485,In_583,In_117);
and U1486 (N_1486,In_530,In_887);
or U1487 (N_1487,In_507,In_667);
nand U1488 (N_1488,In_248,In_929);
and U1489 (N_1489,In_205,In_733);
or U1490 (N_1490,In_305,In_617);
nor U1491 (N_1491,In_830,In_333);
nand U1492 (N_1492,In_925,In_427);
nand U1493 (N_1493,In_783,In_832);
and U1494 (N_1494,In_32,In_13);
nand U1495 (N_1495,In_145,In_181);
or U1496 (N_1496,In_881,In_313);
or U1497 (N_1497,In_471,In_695);
nor U1498 (N_1498,In_18,In_839);
or U1499 (N_1499,In_778,In_987);
nand U1500 (N_1500,In_606,In_762);
nand U1501 (N_1501,In_881,In_582);
or U1502 (N_1502,In_413,In_826);
or U1503 (N_1503,In_28,In_365);
and U1504 (N_1504,In_657,In_694);
or U1505 (N_1505,In_144,In_912);
or U1506 (N_1506,In_180,In_910);
and U1507 (N_1507,In_85,In_407);
nor U1508 (N_1508,In_869,In_338);
or U1509 (N_1509,In_554,In_143);
nand U1510 (N_1510,In_141,In_865);
nand U1511 (N_1511,In_923,In_713);
or U1512 (N_1512,In_115,In_811);
nor U1513 (N_1513,In_509,In_223);
and U1514 (N_1514,In_853,In_27);
or U1515 (N_1515,In_105,In_861);
and U1516 (N_1516,In_43,In_574);
nor U1517 (N_1517,In_832,In_140);
and U1518 (N_1518,In_334,In_214);
and U1519 (N_1519,In_571,In_382);
or U1520 (N_1520,In_268,In_919);
nand U1521 (N_1521,In_263,In_764);
nand U1522 (N_1522,In_947,In_889);
nor U1523 (N_1523,In_267,In_506);
xor U1524 (N_1524,In_215,In_178);
nand U1525 (N_1525,In_904,In_244);
nor U1526 (N_1526,In_334,In_539);
nor U1527 (N_1527,In_556,In_814);
or U1528 (N_1528,In_632,In_866);
and U1529 (N_1529,In_88,In_376);
or U1530 (N_1530,In_716,In_385);
or U1531 (N_1531,In_856,In_764);
and U1532 (N_1532,In_294,In_794);
nand U1533 (N_1533,In_328,In_623);
nand U1534 (N_1534,In_972,In_540);
or U1535 (N_1535,In_970,In_518);
or U1536 (N_1536,In_129,In_81);
nor U1537 (N_1537,In_883,In_126);
nand U1538 (N_1538,In_277,In_584);
and U1539 (N_1539,In_696,In_873);
nand U1540 (N_1540,In_319,In_80);
and U1541 (N_1541,In_604,In_341);
nand U1542 (N_1542,In_637,In_713);
or U1543 (N_1543,In_5,In_831);
nor U1544 (N_1544,In_605,In_755);
and U1545 (N_1545,In_836,In_789);
or U1546 (N_1546,In_924,In_663);
nand U1547 (N_1547,In_799,In_282);
nand U1548 (N_1548,In_807,In_978);
nand U1549 (N_1549,In_552,In_597);
or U1550 (N_1550,In_771,In_569);
or U1551 (N_1551,In_231,In_659);
nand U1552 (N_1552,In_442,In_935);
or U1553 (N_1553,In_32,In_693);
or U1554 (N_1554,In_104,In_92);
nand U1555 (N_1555,In_438,In_517);
or U1556 (N_1556,In_469,In_996);
nand U1557 (N_1557,In_637,In_919);
or U1558 (N_1558,In_630,In_526);
or U1559 (N_1559,In_219,In_697);
or U1560 (N_1560,In_973,In_650);
and U1561 (N_1561,In_718,In_553);
nand U1562 (N_1562,In_296,In_209);
nand U1563 (N_1563,In_489,In_98);
nor U1564 (N_1564,In_753,In_129);
or U1565 (N_1565,In_4,In_10);
and U1566 (N_1566,In_406,In_43);
and U1567 (N_1567,In_846,In_974);
nand U1568 (N_1568,In_179,In_679);
nand U1569 (N_1569,In_60,In_823);
and U1570 (N_1570,In_810,In_288);
nor U1571 (N_1571,In_138,In_59);
nor U1572 (N_1572,In_503,In_274);
or U1573 (N_1573,In_725,In_401);
or U1574 (N_1574,In_825,In_589);
or U1575 (N_1575,In_411,In_26);
and U1576 (N_1576,In_809,In_547);
or U1577 (N_1577,In_667,In_725);
nand U1578 (N_1578,In_737,In_749);
or U1579 (N_1579,In_35,In_244);
nand U1580 (N_1580,In_130,In_734);
and U1581 (N_1581,In_790,In_651);
nor U1582 (N_1582,In_760,In_347);
nor U1583 (N_1583,In_384,In_207);
and U1584 (N_1584,In_120,In_996);
or U1585 (N_1585,In_618,In_725);
nand U1586 (N_1586,In_7,In_574);
or U1587 (N_1587,In_378,In_295);
nand U1588 (N_1588,In_288,In_888);
nand U1589 (N_1589,In_583,In_235);
nor U1590 (N_1590,In_787,In_723);
or U1591 (N_1591,In_929,In_990);
nor U1592 (N_1592,In_628,In_996);
nand U1593 (N_1593,In_94,In_990);
or U1594 (N_1594,In_986,In_70);
and U1595 (N_1595,In_580,In_445);
and U1596 (N_1596,In_694,In_773);
or U1597 (N_1597,In_294,In_137);
nand U1598 (N_1598,In_112,In_20);
nand U1599 (N_1599,In_111,In_409);
nor U1600 (N_1600,In_506,In_583);
nor U1601 (N_1601,In_349,In_289);
or U1602 (N_1602,In_723,In_911);
nor U1603 (N_1603,In_217,In_446);
and U1604 (N_1604,In_870,In_239);
nor U1605 (N_1605,In_950,In_992);
nor U1606 (N_1606,In_940,In_23);
nand U1607 (N_1607,In_353,In_642);
or U1608 (N_1608,In_525,In_701);
and U1609 (N_1609,In_328,In_598);
or U1610 (N_1610,In_222,In_966);
nor U1611 (N_1611,In_943,In_182);
nand U1612 (N_1612,In_858,In_416);
and U1613 (N_1613,In_998,In_339);
nor U1614 (N_1614,In_167,In_484);
or U1615 (N_1615,In_980,In_545);
nor U1616 (N_1616,In_547,In_705);
xnor U1617 (N_1617,In_804,In_273);
nand U1618 (N_1618,In_827,In_543);
nand U1619 (N_1619,In_991,In_92);
or U1620 (N_1620,In_347,In_389);
or U1621 (N_1621,In_501,In_946);
nand U1622 (N_1622,In_657,In_682);
nand U1623 (N_1623,In_127,In_491);
nor U1624 (N_1624,In_559,In_492);
and U1625 (N_1625,In_821,In_322);
nor U1626 (N_1626,In_405,In_860);
nor U1627 (N_1627,In_97,In_783);
and U1628 (N_1628,In_437,In_485);
nand U1629 (N_1629,In_884,In_379);
and U1630 (N_1630,In_478,In_198);
or U1631 (N_1631,In_382,In_670);
nand U1632 (N_1632,In_852,In_111);
or U1633 (N_1633,In_466,In_911);
nor U1634 (N_1634,In_609,In_309);
nor U1635 (N_1635,In_709,In_703);
nor U1636 (N_1636,In_586,In_621);
nand U1637 (N_1637,In_217,In_68);
nand U1638 (N_1638,In_80,In_157);
and U1639 (N_1639,In_309,In_20);
nor U1640 (N_1640,In_777,In_760);
or U1641 (N_1641,In_652,In_462);
or U1642 (N_1642,In_91,In_610);
nor U1643 (N_1643,In_247,In_100);
and U1644 (N_1644,In_341,In_883);
nand U1645 (N_1645,In_893,In_128);
or U1646 (N_1646,In_166,In_505);
nor U1647 (N_1647,In_7,In_34);
nor U1648 (N_1648,In_700,In_302);
nor U1649 (N_1649,In_984,In_159);
or U1650 (N_1650,In_516,In_853);
nor U1651 (N_1651,In_702,In_129);
nand U1652 (N_1652,In_445,In_388);
nor U1653 (N_1653,In_862,In_586);
nor U1654 (N_1654,In_217,In_143);
nand U1655 (N_1655,In_380,In_17);
or U1656 (N_1656,In_11,In_830);
nor U1657 (N_1657,In_834,In_614);
nand U1658 (N_1658,In_166,In_408);
or U1659 (N_1659,In_112,In_121);
or U1660 (N_1660,In_659,In_357);
or U1661 (N_1661,In_835,In_910);
nor U1662 (N_1662,In_96,In_38);
or U1663 (N_1663,In_814,In_60);
nand U1664 (N_1664,In_149,In_457);
nor U1665 (N_1665,In_990,In_236);
and U1666 (N_1666,In_855,In_599);
xnor U1667 (N_1667,In_978,In_959);
and U1668 (N_1668,In_652,In_592);
or U1669 (N_1669,In_796,In_336);
and U1670 (N_1670,In_743,In_133);
nand U1671 (N_1671,In_591,In_343);
or U1672 (N_1672,In_334,In_857);
nand U1673 (N_1673,In_571,In_302);
and U1674 (N_1674,In_694,In_522);
nand U1675 (N_1675,In_639,In_908);
nand U1676 (N_1676,In_805,In_589);
and U1677 (N_1677,In_73,In_98);
or U1678 (N_1678,In_837,In_984);
nand U1679 (N_1679,In_139,In_489);
and U1680 (N_1680,In_88,In_74);
nand U1681 (N_1681,In_241,In_784);
and U1682 (N_1682,In_523,In_752);
or U1683 (N_1683,In_332,In_871);
or U1684 (N_1684,In_965,In_635);
or U1685 (N_1685,In_722,In_950);
and U1686 (N_1686,In_59,In_801);
and U1687 (N_1687,In_633,In_439);
and U1688 (N_1688,In_930,In_701);
nor U1689 (N_1689,In_479,In_298);
or U1690 (N_1690,In_936,In_46);
nor U1691 (N_1691,In_914,In_432);
nor U1692 (N_1692,In_612,In_848);
nand U1693 (N_1693,In_879,In_771);
or U1694 (N_1694,In_267,In_316);
nand U1695 (N_1695,In_741,In_941);
xor U1696 (N_1696,In_114,In_713);
nand U1697 (N_1697,In_0,In_57);
nor U1698 (N_1698,In_949,In_124);
and U1699 (N_1699,In_388,In_131);
and U1700 (N_1700,In_409,In_936);
or U1701 (N_1701,In_663,In_402);
or U1702 (N_1702,In_662,In_251);
and U1703 (N_1703,In_114,In_790);
nand U1704 (N_1704,In_357,In_429);
nor U1705 (N_1705,In_615,In_753);
nor U1706 (N_1706,In_869,In_526);
or U1707 (N_1707,In_989,In_560);
and U1708 (N_1708,In_853,In_400);
or U1709 (N_1709,In_150,In_311);
or U1710 (N_1710,In_660,In_12);
nand U1711 (N_1711,In_290,In_440);
or U1712 (N_1712,In_9,In_824);
or U1713 (N_1713,In_200,In_45);
nor U1714 (N_1714,In_83,In_65);
nand U1715 (N_1715,In_281,In_47);
nand U1716 (N_1716,In_280,In_840);
nor U1717 (N_1717,In_153,In_290);
nor U1718 (N_1718,In_630,In_510);
and U1719 (N_1719,In_843,In_987);
and U1720 (N_1720,In_856,In_230);
nand U1721 (N_1721,In_370,In_408);
nand U1722 (N_1722,In_990,In_643);
and U1723 (N_1723,In_492,In_891);
nand U1724 (N_1724,In_585,In_156);
and U1725 (N_1725,In_211,In_973);
nor U1726 (N_1726,In_676,In_255);
nand U1727 (N_1727,In_629,In_439);
or U1728 (N_1728,In_811,In_303);
and U1729 (N_1729,In_211,In_390);
nand U1730 (N_1730,In_730,In_871);
or U1731 (N_1731,In_95,In_15);
nand U1732 (N_1732,In_36,In_409);
nand U1733 (N_1733,In_27,In_725);
or U1734 (N_1734,In_977,In_133);
nand U1735 (N_1735,In_242,In_762);
nand U1736 (N_1736,In_412,In_249);
nand U1737 (N_1737,In_104,In_763);
and U1738 (N_1738,In_689,In_856);
nor U1739 (N_1739,In_799,In_936);
nand U1740 (N_1740,In_805,In_720);
or U1741 (N_1741,In_911,In_16);
nor U1742 (N_1742,In_147,In_410);
or U1743 (N_1743,In_910,In_532);
nand U1744 (N_1744,In_134,In_59);
nand U1745 (N_1745,In_970,In_683);
and U1746 (N_1746,In_872,In_974);
or U1747 (N_1747,In_798,In_0);
nand U1748 (N_1748,In_109,In_290);
and U1749 (N_1749,In_995,In_790);
nand U1750 (N_1750,In_372,In_475);
or U1751 (N_1751,In_519,In_488);
and U1752 (N_1752,In_480,In_954);
or U1753 (N_1753,In_529,In_86);
nor U1754 (N_1754,In_210,In_906);
nor U1755 (N_1755,In_993,In_553);
nand U1756 (N_1756,In_642,In_848);
nor U1757 (N_1757,In_328,In_34);
nor U1758 (N_1758,In_639,In_623);
nor U1759 (N_1759,In_984,In_835);
and U1760 (N_1760,In_17,In_414);
nor U1761 (N_1761,In_447,In_547);
nand U1762 (N_1762,In_356,In_530);
nor U1763 (N_1763,In_137,In_299);
or U1764 (N_1764,In_383,In_800);
nand U1765 (N_1765,In_57,In_640);
or U1766 (N_1766,In_22,In_484);
and U1767 (N_1767,In_617,In_895);
nand U1768 (N_1768,In_15,In_768);
nor U1769 (N_1769,In_927,In_215);
or U1770 (N_1770,In_811,In_108);
and U1771 (N_1771,In_987,In_193);
nor U1772 (N_1772,In_471,In_494);
nand U1773 (N_1773,In_975,In_107);
nor U1774 (N_1774,In_215,In_477);
nor U1775 (N_1775,In_663,In_601);
or U1776 (N_1776,In_160,In_244);
nor U1777 (N_1777,In_197,In_625);
or U1778 (N_1778,In_18,In_162);
nand U1779 (N_1779,In_2,In_600);
and U1780 (N_1780,In_38,In_937);
nand U1781 (N_1781,In_36,In_690);
and U1782 (N_1782,In_572,In_276);
and U1783 (N_1783,In_615,In_549);
nor U1784 (N_1784,In_408,In_173);
and U1785 (N_1785,In_414,In_901);
nor U1786 (N_1786,In_869,In_729);
nor U1787 (N_1787,In_98,In_263);
or U1788 (N_1788,In_768,In_498);
or U1789 (N_1789,In_16,In_724);
and U1790 (N_1790,In_138,In_105);
nor U1791 (N_1791,In_894,In_572);
or U1792 (N_1792,In_747,In_417);
or U1793 (N_1793,In_686,In_95);
nand U1794 (N_1794,In_340,In_951);
and U1795 (N_1795,In_767,In_45);
nand U1796 (N_1796,In_554,In_684);
or U1797 (N_1797,In_739,In_578);
nand U1798 (N_1798,In_492,In_68);
nor U1799 (N_1799,In_120,In_136);
xnor U1800 (N_1800,In_939,In_319);
nor U1801 (N_1801,In_818,In_122);
and U1802 (N_1802,In_519,In_784);
nor U1803 (N_1803,In_640,In_814);
or U1804 (N_1804,In_495,In_147);
and U1805 (N_1805,In_281,In_549);
and U1806 (N_1806,In_747,In_679);
nand U1807 (N_1807,In_954,In_709);
nor U1808 (N_1808,In_516,In_724);
or U1809 (N_1809,In_304,In_174);
or U1810 (N_1810,In_758,In_327);
and U1811 (N_1811,In_857,In_484);
and U1812 (N_1812,In_751,In_631);
or U1813 (N_1813,In_249,In_665);
nor U1814 (N_1814,In_829,In_493);
nor U1815 (N_1815,In_956,In_77);
nand U1816 (N_1816,In_19,In_403);
and U1817 (N_1817,In_214,In_91);
nor U1818 (N_1818,In_877,In_408);
nand U1819 (N_1819,In_980,In_14);
nand U1820 (N_1820,In_996,In_72);
nor U1821 (N_1821,In_462,In_49);
nor U1822 (N_1822,In_569,In_746);
and U1823 (N_1823,In_889,In_689);
nand U1824 (N_1824,In_735,In_506);
and U1825 (N_1825,In_811,In_185);
or U1826 (N_1826,In_971,In_482);
and U1827 (N_1827,In_170,In_832);
and U1828 (N_1828,In_599,In_33);
and U1829 (N_1829,In_88,In_473);
nand U1830 (N_1830,In_159,In_7);
and U1831 (N_1831,In_993,In_857);
or U1832 (N_1832,In_411,In_167);
nand U1833 (N_1833,In_895,In_476);
nand U1834 (N_1834,In_690,In_96);
or U1835 (N_1835,In_318,In_966);
nor U1836 (N_1836,In_808,In_45);
nand U1837 (N_1837,In_430,In_822);
and U1838 (N_1838,In_637,In_682);
or U1839 (N_1839,In_983,In_112);
and U1840 (N_1840,In_641,In_143);
and U1841 (N_1841,In_383,In_250);
or U1842 (N_1842,In_55,In_154);
nor U1843 (N_1843,In_56,In_650);
and U1844 (N_1844,In_262,In_317);
and U1845 (N_1845,In_831,In_215);
and U1846 (N_1846,In_97,In_791);
and U1847 (N_1847,In_671,In_725);
and U1848 (N_1848,In_976,In_224);
or U1849 (N_1849,In_960,In_39);
and U1850 (N_1850,In_804,In_13);
and U1851 (N_1851,In_672,In_716);
nor U1852 (N_1852,In_880,In_803);
nor U1853 (N_1853,In_945,In_4);
nor U1854 (N_1854,In_577,In_664);
and U1855 (N_1855,In_377,In_346);
xnor U1856 (N_1856,In_75,In_985);
nand U1857 (N_1857,In_124,In_135);
and U1858 (N_1858,In_155,In_983);
nand U1859 (N_1859,In_961,In_281);
and U1860 (N_1860,In_372,In_541);
or U1861 (N_1861,In_86,In_417);
and U1862 (N_1862,In_549,In_292);
nor U1863 (N_1863,In_725,In_952);
nor U1864 (N_1864,In_322,In_636);
nand U1865 (N_1865,In_559,In_944);
nand U1866 (N_1866,In_430,In_990);
nor U1867 (N_1867,In_273,In_748);
or U1868 (N_1868,In_898,In_298);
and U1869 (N_1869,In_409,In_878);
and U1870 (N_1870,In_845,In_75);
nand U1871 (N_1871,In_235,In_627);
or U1872 (N_1872,In_874,In_590);
and U1873 (N_1873,In_400,In_877);
xor U1874 (N_1874,In_15,In_880);
nand U1875 (N_1875,In_946,In_808);
and U1876 (N_1876,In_410,In_986);
and U1877 (N_1877,In_818,In_867);
nand U1878 (N_1878,In_780,In_456);
and U1879 (N_1879,In_309,In_979);
or U1880 (N_1880,In_773,In_969);
or U1881 (N_1881,In_886,In_155);
or U1882 (N_1882,In_515,In_264);
nand U1883 (N_1883,In_645,In_977);
or U1884 (N_1884,In_462,In_713);
nor U1885 (N_1885,In_990,In_598);
or U1886 (N_1886,In_590,In_947);
nand U1887 (N_1887,In_15,In_481);
nand U1888 (N_1888,In_726,In_215);
nor U1889 (N_1889,In_21,In_222);
nand U1890 (N_1890,In_202,In_668);
and U1891 (N_1891,In_730,In_200);
nor U1892 (N_1892,In_624,In_763);
nor U1893 (N_1893,In_75,In_417);
nor U1894 (N_1894,In_965,In_112);
nor U1895 (N_1895,In_982,In_713);
and U1896 (N_1896,In_35,In_855);
nand U1897 (N_1897,In_443,In_902);
and U1898 (N_1898,In_310,In_5);
or U1899 (N_1899,In_143,In_98);
nand U1900 (N_1900,In_770,In_681);
xnor U1901 (N_1901,In_882,In_603);
nor U1902 (N_1902,In_933,In_616);
and U1903 (N_1903,In_179,In_948);
and U1904 (N_1904,In_571,In_324);
nor U1905 (N_1905,In_18,In_524);
nor U1906 (N_1906,In_152,In_823);
and U1907 (N_1907,In_130,In_267);
and U1908 (N_1908,In_269,In_103);
nand U1909 (N_1909,In_373,In_495);
nor U1910 (N_1910,In_537,In_744);
or U1911 (N_1911,In_949,In_886);
or U1912 (N_1912,In_859,In_94);
nand U1913 (N_1913,In_136,In_196);
nor U1914 (N_1914,In_433,In_127);
nand U1915 (N_1915,In_401,In_29);
and U1916 (N_1916,In_335,In_538);
nor U1917 (N_1917,In_51,In_620);
nor U1918 (N_1918,In_576,In_297);
and U1919 (N_1919,In_30,In_406);
or U1920 (N_1920,In_76,In_518);
nor U1921 (N_1921,In_541,In_762);
or U1922 (N_1922,In_822,In_615);
nand U1923 (N_1923,In_171,In_494);
and U1924 (N_1924,In_574,In_445);
and U1925 (N_1925,In_205,In_897);
nand U1926 (N_1926,In_598,In_570);
nor U1927 (N_1927,In_254,In_116);
nor U1928 (N_1928,In_873,In_136);
and U1929 (N_1929,In_335,In_314);
nand U1930 (N_1930,In_401,In_86);
nor U1931 (N_1931,In_886,In_502);
or U1932 (N_1932,In_933,In_354);
or U1933 (N_1933,In_331,In_957);
nand U1934 (N_1934,In_545,In_758);
or U1935 (N_1935,In_215,In_597);
or U1936 (N_1936,In_795,In_876);
nor U1937 (N_1937,In_329,In_269);
nor U1938 (N_1938,In_903,In_985);
nand U1939 (N_1939,In_115,In_204);
or U1940 (N_1940,In_806,In_909);
nand U1941 (N_1941,In_462,In_791);
nand U1942 (N_1942,In_907,In_105);
or U1943 (N_1943,In_282,In_124);
and U1944 (N_1944,In_263,In_636);
or U1945 (N_1945,In_641,In_130);
nor U1946 (N_1946,In_520,In_210);
nor U1947 (N_1947,In_824,In_586);
or U1948 (N_1948,In_573,In_448);
nor U1949 (N_1949,In_913,In_637);
nand U1950 (N_1950,In_417,In_230);
or U1951 (N_1951,In_26,In_262);
nor U1952 (N_1952,In_745,In_932);
nor U1953 (N_1953,In_842,In_44);
and U1954 (N_1954,In_925,In_132);
nand U1955 (N_1955,In_83,In_545);
nand U1956 (N_1956,In_922,In_959);
or U1957 (N_1957,In_340,In_360);
and U1958 (N_1958,In_298,In_122);
and U1959 (N_1959,In_212,In_815);
and U1960 (N_1960,In_802,In_580);
or U1961 (N_1961,In_137,In_502);
and U1962 (N_1962,In_670,In_698);
nand U1963 (N_1963,In_341,In_817);
and U1964 (N_1964,In_111,In_945);
nand U1965 (N_1965,In_570,In_36);
or U1966 (N_1966,In_209,In_233);
and U1967 (N_1967,In_470,In_640);
nand U1968 (N_1968,In_121,In_610);
and U1969 (N_1969,In_851,In_154);
and U1970 (N_1970,In_515,In_32);
nor U1971 (N_1971,In_886,In_92);
nand U1972 (N_1972,In_202,In_361);
and U1973 (N_1973,In_106,In_279);
or U1974 (N_1974,In_690,In_719);
nor U1975 (N_1975,In_979,In_141);
nand U1976 (N_1976,In_436,In_387);
nor U1977 (N_1977,In_229,In_988);
or U1978 (N_1978,In_585,In_177);
or U1979 (N_1979,In_54,In_599);
nand U1980 (N_1980,In_367,In_501);
nor U1981 (N_1981,In_592,In_237);
nand U1982 (N_1982,In_655,In_25);
nand U1983 (N_1983,In_756,In_846);
nor U1984 (N_1984,In_971,In_413);
nor U1985 (N_1985,In_191,In_361);
and U1986 (N_1986,In_561,In_373);
nor U1987 (N_1987,In_664,In_584);
nor U1988 (N_1988,In_476,In_947);
and U1989 (N_1989,In_153,In_527);
or U1990 (N_1990,In_797,In_447);
nand U1991 (N_1991,In_489,In_222);
xor U1992 (N_1992,In_892,In_281);
or U1993 (N_1993,In_739,In_77);
and U1994 (N_1994,In_405,In_301);
nand U1995 (N_1995,In_470,In_664);
and U1996 (N_1996,In_511,In_637);
or U1997 (N_1997,In_379,In_832);
or U1998 (N_1998,In_726,In_498);
nand U1999 (N_1999,In_103,In_549);
nand U2000 (N_2000,In_298,In_577);
and U2001 (N_2001,In_44,In_426);
and U2002 (N_2002,In_759,In_904);
nand U2003 (N_2003,In_340,In_949);
and U2004 (N_2004,In_205,In_759);
nor U2005 (N_2005,In_687,In_718);
nor U2006 (N_2006,In_570,In_125);
nor U2007 (N_2007,In_730,In_731);
or U2008 (N_2008,In_400,In_818);
nand U2009 (N_2009,In_862,In_127);
nor U2010 (N_2010,In_375,In_128);
nand U2011 (N_2011,In_244,In_647);
or U2012 (N_2012,In_610,In_882);
nor U2013 (N_2013,In_285,In_791);
nand U2014 (N_2014,In_974,In_241);
nand U2015 (N_2015,In_101,In_977);
or U2016 (N_2016,In_380,In_149);
or U2017 (N_2017,In_273,In_434);
nand U2018 (N_2018,In_360,In_422);
nand U2019 (N_2019,In_350,In_749);
or U2020 (N_2020,In_930,In_976);
or U2021 (N_2021,In_892,In_8);
nand U2022 (N_2022,In_88,In_736);
or U2023 (N_2023,In_405,In_366);
nor U2024 (N_2024,In_130,In_56);
or U2025 (N_2025,In_516,In_327);
nand U2026 (N_2026,In_825,In_81);
nor U2027 (N_2027,In_314,In_600);
nand U2028 (N_2028,In_573,In_548);
nand U2029 (N_2029,In_404,In_189);
and U2030 (N_2030,In_933,In_893);
or U2031 (N_2031,In_408,In_742);
nor U2032 (N_2032,In_96,In_229);
and U2033 (N_2033,In_94,In_913);
nand U2034 (N_2034,In_441,In_333);
and U2035 (N_2035,In_919,In_323);
nor U2036 (N_2036,In_437,In_592);
nand U2037 (N_2037,In_946,In_254);
or U2038 (N_2038,In_876,In_517);
nand U2039 (N_2039,In_905,In_611);
nand U2040 (N_2040,In_132,In_664);
and U2041 (N_2041,In_490,In_609);
nor U2042 (N_2042,In_613,In_468);
and U2043 (N_2043,In_891,In_341);
nand U2044 (N_2044,In_248,In_252);
and U2045 (N_2045,In_213,In_685);
and U2046 (N_2046,In_31,In_206);
nand U2047 (N_2047,In_318,In_451);
and U2048 (N_2048,In_366,In_610);
nand U2049 (N_2049,In_437,In_210);
nor U2050 (N_2050,In_647,In_527);
nor U2051 (N_2051,In_60,In_232);
or U2052 (N_2052,In_750,In_687);
nor U2053 (N_2053,In_187,In_82);
and U2054 (N_2054,In_37,In_868);
or U2055 (N_2055,In_459,In_245);
xor U2056 (N_2056,In_892,In_54);
nor U2057 (N_2057,In_208,In_980);
nand U2058 (N_2058,In_422,In_516);
and U2059 (N_2059,In_452,In_782);
nand U2060 (N_2060,In_591,In_74);
and U2061 (N_2061,In_631,In_16);
and U2062 (N_2062,In_857,In_193);
or U2063 (N_2063,In_317,In_161);
or U2064 (N_2064,In_176,In_553);
nor U2065 (N_2065,In_19,In_570);
and U2066 (N_2066,In_206,In_276);
nand U2067 (N_2067,In_57,In_649);
and U2068 (N_2068,In_24,In_156);
or U2069 (N_2069,In_817,In_533);
or U2070 (N_2070,In_592,In_8);
or U2071 (N_2071,In_78,In_477);
nand U2072 (N_2072,In_506,In_869);
and U2073 (N_2073,In_281,In_224);
nor U2074 (N_2074,In_170,In_452);
or U2075 (N_2075,In_252,In_854);
and U2076 (N_2076,In_943,In_281);
nand U2077 (N_2077,In_775,In_149);
or U2078 (N_2078,In_667,In_512);
nand U2079 (N_2079,In_644,In_853);
nor U2080 (N_2080,In_751,In_719);
and U2081 (N_2081,In_558,In_190);
and U2082 (N_2082,In_51,In_773);
or U2083 (N_2083,In_940,In_820);
nand U2084 (N_2084,In_934,In_440);
and U2085 (N_2085,In_684,In_440);
and U2086 (N_2086,In_974,In_455);
nand U2087 (N_2087,In_128,In_411);
and U2088 (N_2088,In_199,In_145);
nand U2089 (N_2089,In_187,In_817);
or U2090 (N_2090,In_561,In_678);
or U2091 (N_2091,In_468,In_815);
or U2092 (N_2092,In_815,In_158);
nor U2093 (N_2093,In_506,In_986);
nand U2094 (N_2094,In_909,In_237);
or U2095 (N_2095,In_832,In_472);
nor U2096 (N_2096,In_388,In_812);
and U2097 (N_2097,In_881,In_570);
nand U2098 (N_2098,In_144,In_504);
nor U2099 (N_2099,In_519,In_140);
or U2100 (N_2100,In_220,In_341);
nor U2101 (N_2101,In_227,In_835);
nand U2102 (N_2102,In_10,In_629);
nand U2103 (N_2103,In_297,In_664);
and U2104 (N_2104,In_978,In_856);
nor U2105 (N_2105,In_154,In_604);
nor U2106 (N_2106,In_617,In_182);
nand U2107 (N_2107,In_973,In_571);
nand U2108 (N_2108,In_362,In_436);
nor U2109 (N_2109,In_758,In_250);
and U2110 (N_2110,In_523,In_622);
nand U2111 (N_2111,In_100,In_689);
and U2112 (N_2112,In_74,In_526);
and U2113 (N_2113,In_104,In_252);
nand U2114 (N_2114,In_229,In_772);
or U2115 (N_2115,In_128,In_503);
nor U2116 (N_2116,In_996,In_729);
and U2117 (N_2117,In_439,In_641);
or U2118 (N_2118,In_924,In_165);
or U2119 (N_2119,In_128,In_59);
nand U2120 (N_2120,In_130,In_623);
nor U2121 (N_2121,In_383,In_545);
nand U2122 (N_2122,In_506,In_436);
nor U2123 (N_2123,In_461,In_217);
nand U2124 (N_2124,In_939,In_636);
and U2125 (N_2125,In_724,In_239);
and U2126 (N_2126,In_392,In_536);
nand U2127 (N_2127,In_196,In_291);
or U2128 (N_2128,In_704,In_720);
and U2129 (N_2129,In_39,In_435);
nand U2130 (N_2130,In_787,In_26);
nor U2131 (N_2131,In_632,In_212);
and U2132 (N_2132,In_481,In_748);
nand U2133 (N_2133,In_142,In_363);
and U2134 (N_2134,In_733,In_69);
or U2135 (N_2135,In_149,In_32);
nor U2136 (N_2136,In_327,In_391);
and U2137 (N_2137,In_574,In_64);
nand U2138 (N_2138,In_830,In_441);
or U2139 (N_2139,In_284,In_195);
or U2140 (N_2140,In_502,In_318);
or U2141 (N_2141,In_207,In_166);
or U2142 (N_2142,In_143,In_394);
or U2143 (N_2143,In_725,In_713);
or U2144 (N_2144,In_766,In_129);
or U2145 (N_2145,In_24,In_530);
nor U2146 (N_2146,In_413,In_743);
nand U2147 (N_2147,In_514,In_571);
nor U2148 (N_2148,In_91,In_465);
or U2149 (N_2149,In_642,In_968);
nand U2150 (N_2150,In_645,In_280);
or U2151 (N_2151,In_213,In_646);
or U2152 (N_2152,In_228,In_852);
or U2153 (N_2153,In_383,In_665);
and U2154 (N_2154,In_794,In_971);
nand U2155 (N_2155,In_816,In_85);
nor U2156 (N_2156,In_970,In_231);
or U2157 (N_2157,In_273,In_424);
or U2158 (N_2158,In_184,In_129);
nand U2159 (N_2159,In_503,In_254);
nor U2160 (N_2160,In_470,In_617);
nand U2161 (N_2161,In_64,In_827);
and U2162 (N_2162,In_316,In_692);
nand U2163 (N_2163,In_170,In_384);
nor U2164 (N_2164,In_389,In_62);
nand U2165 (N_2165,In_144,In_790);
nor U2166 (N_2166,In_554,In_740);
and U2167 (N_2167,In_946,In_315);
nand U2168 (N_2168,In_832,In_245);
nor U2169 (N_2169,In_278,In_264);
nand U2170 (N_2170,In_7,In_505);
or U2171 (N_2171,In_601,In_553);
nand U2172 (N_2172,In_759,In_78);
nor U2173 (N_2173,In_269,In_201);
nand U2174 (N_2174,In_447,In_667);
or U2175 (N_2175,In_137,In_212);
nand U2176 (N_2176,In_133,In_289);
and U2177 (N_2177,In_820,In_702);
nor U2178 (N_2178,In_489,In_824);
nor U2179 (N_2179,In_213,In_238);
nand U2180 (N_2180,In_977,In_852);
or U2181 (N_2181,In_499,In_846);
nand U2182 (N_2182,In_855,In_342);
nand U2183 (N_2183,In_419,In_872);
or U2184 (N_2184,In_52,In_157);
nand U2185 (N_2185,In_901,In_937);
nand U2186 (N_2186,In_66,In_391);
nor U2187 (N_2187,In_915,In_927);
or U2188 (N_2188,In_362,In_339);
nor U2189 (N_2189,In_747,In_133);
nor U2190 (N_2190,In_684,In_225);
nor U2191 (N_2191,In_184,In_618);
nor U2192 (N_2192,In_545,In_946);
nor U2193 (N_2193,In_269,In_834);
nand U2194 (N_2194,In_381,In_234);
nand U2195 (N_2195,In_377,In_200);
and U2196 (N_2196,In_485,In_587);
nand U2197 (N_2197,In_228,In_258);
nand U2198 (N_2198,In_877,In_444);
or U2199 (N_2199,In_179,In_197);
nand U2200 (N_2200,In_311,In_483);
nand U2201 (N_2201,In_774,In_220);
and U2202 (N_2202,In_523,In_242);
nand U2203 (N_2203,In_137,In_799);
and U2204 (N_2204,In_599,In_549);
nand U2205 (N_2205,In_303,In_993);
or U2206 (N_2206,In_431,In_420);
nor U2207 (N_2207,In_394,In_604);
and U2208 (N_2208,In_474,In_927);
and U2209 (N_2209,In_771,In_965);
nor U2210 (N_2210,In_36,In_935);
and U2211 (N_2211,In_966,In_932);
and U2212 (N_2212,In_340,In_139);
nor U2213 (N_2213,In_993,In_507);
and U2214 (N_2214,In_628,In_351);
nor U2215 (N_2215,In_59,In_579);
nand U2216 (N_2216,In_634,In_972);
nand U2217 (N_2217,In_617,In_61);
and U2218 (N_2218,In_942,In_512);
nand U2219 (N_2219,In_884,In_339);
and U2220 (N_2220,In_783,In_124);
and U2221 (N_2221,In_664,In_757);
nor U2222 (N_2222,In_910,In_645);
nand U2223 (N_2223,In_927,In_152);
or U2224 (N_2224,In_133,In_890);
nor U2225 (N_2225,In_549,In_457);
or U2226 (N_2226,In_611,In_844);
and U2227 (N_2227,In_270,In_220);
nand U2228 (N_2228,In_804,In_781);
nor U2229 (N_2229,In_470,In_453);
nand U2230 (N_2230,In_670,In_377);
or U2231 (N_2231,In_365,In_465);
nand U2232 (N_2232,In_688,In_565);
and U2233 (N_2233,In_989,In_944);
nand U2234 (N_2234,In_577,In_154);
or U2235 (N_2235,In_277,In_85);
or U2236 (N_2236,In_248,In_957);
nor U2237 (N_2237,In_638,In_604);
and U2238 (N_2238,In_130,In_553);
or U2239 (N_2239,In_990,In_354);
nand U2240 (N_2240,In_940,In_510);
and U2241 (N_2241,In_115,In_554);
nor U2242 (N_2242,In_247,In_852);
or U2243 (N_2243,In_25,In_936);
and U2244 (N_2244,In_650,In_458);
nor U2245 (N_2245,In_908,In_603);
and U2246 (N_2246,In_32,In_205);
or U2247 (N_2247,In_354,In_410);
nor U2248 (N_2248,In_499,In_193);
or U2249 (N_2249,In_604,In_307);
nand U2250 (N_2250,In_125,In_352);
and U2251 (N_2251,In_146,In_436);
nand U2252 (N_2252,In_986,In_662);
and U2253 (N_2253,In_252,In_456);
or U2254 (N_2254,In_343,In_765);
nand U2255 (N_2255,In_628,In_64);
or U2256 (N_2256,In_507,In_404);
and U2257 (N_2257,In_991,In_562);
nand U2258 (N_2258,In_465,In_104);
and U2259 (N_2259,In_831,In_235);
nor U2260 (N_2260,In_118,In_142);
and U2261 (N_2261,In_67,In_734);
and U2262 (N_2262,In_180,In_510);
nor U2263 (N_2263,In_293,In_798);
nor U2264 (N_2264,In_255,In_975);
nor U2265 (N_2265,In_461,In_150);
or U2266 (N_2266,In_723,In_364);
or U2267 (N_2267,In_426,In_785);
or U2268 (N_2268,In_134,In_31);
nand U2269 (N_2269,In_121,In_539);
and U2270 (N_2270,In_190,In_692);
nand U2271 (N_2271,In_281,In_650);
nand U2272 (N_2272,In_859,In_948);
or U2273 (N_2273,In_869,In_627);
and U2274 (N_2274,In_861,In_690);
and U2275 (N_2275,In_141,In_221);
nor U2276 (N_2276,In_923,In_43);
nor U2277 (N_2277,In_911,In_814);
and U2278 (N_2278,In_24,In_916);
or U2279 (N_2279,In_868,In_407);
or U2280 (N_2280,In_719,In_348);
and U2281 (N_2281,In_692,In_449);
or U2282 (N_2282,In_880,In_936);
nor U2283 (N_2283,In_20,In_660);
nand U2284 (N_2284,In_422,In_103);
and U2285 (N_2285,In_860,In_891);
or U2286 (N_2286,In_209,In_593);
nand U2287 (N_2287,In_69,In_118);
or U2288 (N_2288,In_748,In_637);
nand U2289 (N_2289,In_686,In_608);
and U2290 (N_2290,In_951,In_38);
and U2291 (N_2291,In_646,In_264);
or U2292 (N_2292,In_855,In_62);
nand U2293 (N_2293,In_96,In_484);
nand U2294 (N_2294,In_891,In_665);
or U2295 (N_2295,In_131,In_254);
nor U2296 (N_2296,In_600,In_667);
or U2297 (N_2297,In_2,In_907);
nor U2298 (N_2298,In_942,In_751);
or U2299 (N_2299,In_881,In_172);
or U2300 (N_2300,In_457,In_827);
or U2301 (N_2301,In_699,In_109);
and U2302 (N_2302,In_18,In_458);
or U2303 (N_2303,In_226,In_54);
and U2304 (N_2304,In_15,In_436);
nand U2305 (N_2305,In_467,In_585);
nor U2306 (N_2306,In_240,In_189);
nor U2307 (N_2307,In_40,In_166);
xnor U2308 (N_2308,In_285,In_43);
or U2309 (N_2309,In_429,In_655);
and U2310 (N_2310,In_870,In_249);
nor U2311 (N_2311,In_434,In_531);
or U2312 (N_2312,In_60,In_956);
and U2313 (N_2313,In_305,In_681);
or U2314 (N_2314,In_986,In_413);
or U2315 (N_2315,In_281,In_479);
and U2316 (N_2316,In_438,In_75);
nand U2317 (N_2317,In_204,In_448);
or U2318 (N_2318,In_138,In_826);
and U2319 (N_2319,In_825,In_211);
nand U2320 (N_2320,In_101,In_370);
nor U2321 (N_2321,In_860,In_6);
or U2322 (N_2322,In_883,In_420);
and U2323 (N_2323,In_693,In_916);
or U2324 (N_2324,In_14,In_5);
nor U2325 (N_2325,In_407,In_433);
nor U2326 (N_2326,In_813,In_495);
or U2327 (N_2327,In_469,In_773);
nor U2328 (N_2328,In_718,In_343);
or U2329 (N_2329,In_482,In_664);
nor U2330 (N_2330,In_258,In_76);
and U2331 (N_2331,In_446,In_988);
nor U2332 (N_2332,In_370,In_659);
and U2333 (N_2333,In_747,In_583);
nand U2334 (N_2334,In_173,In_790);
or U2335 (N_2335,In_49,In_299);
or U2336 (N_2336,In_341,In_868);
and U2337 (N_2337,In_39,In_963);
xnor U2338 (N_2338,In_746,In_832);
nand U2339 (N_2339,In_568,In_760);
or U2340 (N_2340,In_688,In_370);
and U2341 (N_2341,In_370,In_879);
nand U2342 (N_2342,In_961,In_29);
nor U2343 (N_2343,In_464,In_783);
nor U2344 (N_2344,In_126,In_986);
nor U2345 (N_2345,In_219,In_713);
and U2346 (N_2346,In_968,In_249);
nand U2347 (N_2347,In_290,In_811);
and U2348 (N_2348,In_314,In_728);
nand U2349 (N_2349,In_283,In_155);
nand U2350 (N_2350,In_415,In_778);
and U2351 (N_2351,In_865,In_148);
or U2352 (N_2352,In_281,In_417);
or U2353 (N_2353,In_317,In_285);
or U2354 (N_2354,In_589,In_279);
nand U2355 (N_2355,In_20,In_69);
nor U2356 (N_2356,In_938,In_376);
or U2357 (N_2357,In_804,In_653);
nand U2358 (N_2358,In_971,In_547);
or U2359 (N_2359,In_383,In_319);
or U2360 (N_2360,In_618,In_589);
nor U2361 (N_2361,In_817,In_952);
nand U2362 (N_2362,In_141,In_642);
nand U2363 (N_2363,In_464,In_235);
nor U2364 (N_2364,In_176,In_730);
nand U2365 (N_2365,In_892,In_592);
nand U2366 (N_2366,In_292,In_80);
or U2367 (N_2367,In_789,In_756);
nor U2368 (N_2368,In_90,In_621);
or U2369 (N_2369,In_299,In_411);
or U2370 (N_2370,In_539,In_911);
and U2371 (N_2371,In_77,In_99);
nor U2372 (N_2372,In_556,In_197);
or U2373 (N_2373,In_902,In_174);
nor U2374 (N_2374,In_718,In_661);
or U2375 (N_2375,In_413,In_977);
and U2376 (N_2376,In_195,In_597);
and U2377 (N_2377,In_627,In_749);
and U2378 (N_2378,In_6,In_419);
nand U2379 (N_2379,In_947,In_507);
nor U2380 (N_2380,In_563,In_484);
and U2381 (N_2381,In_596,In_467);
or U2382 (N_2382,In_236,In_879);
nand U2383 (N_2383,In_844,In_711);
nand U2384 (N_2384,In_571,In_428);
nand U2385 (N_2385,In_102,In_722);
and U2386 (N_2386,In_802,In_349);
and U2387 (N_2387,In_947,In_806);
and U2388 (N_2388,In_830,In_635);
or U2389 (N_2389,In_401,In_208);
and U2390 (N_2390,In_563,In_698);
nor U2391 (N_2391,In_830,In_744);
nor U2392 (N_2392,In_981,In_815);
and U2393 (N_2393,In_663,In_640);
nand U2394 (N_2394,In_126,In_580);
and U2395 (N_2395,In_511,In_166);
nand U2396 (N_2396,In_290,In_908);
and U2397 (N_2397,In_273,In_866);
nand U2398 (N_2398,In_511,In_457);
nand U2399 (N_2399,In_243,In_228);
and U2400 (N_2400,In_915,In_515);
or U2401 (N_2401,In_658,In_612);
or U2402 (N_2402,In_492,In_58);
nor U2403 (N_2403,In_528,In_293);
nor U2404 (N_2404,In_175,In_858);
nand U2405 (N_2405,In_576,In_577);
nor U2406 (N_2406,In_336,In_142);
and U2407 (N_2407,In_547,In_900);
nand U2408 (N_2408,In_958,In_803);
nand U2409 (N_2409,In_244,In_884);
nor U2410 (N_2410,In_476,In_258);
nor U2411 (N_2411,In_326,In_972);
nor U2412 (N_2412,In_550,In_885);
nor U2413 (N_2413,In_331,In_329);
or U2414 (N_2414,In_580,In_218);
nand U2415 (N_2415,In_577,In_107);
and U2416 (N_2416,In_606,In_498);
nor U2417 (N_2417,In_971,In_643);
or U2418 (N_2418,In_318,In_243);
or U2419 (N_2419,In_997,In_13);
and U2420 (N_2420,In_801,In_280);
and U2421 (N_2421,In_200,In_108);
nand U2422 (N_2422,In_400,In_981);
nor U2423 (N_2423,In_852,In_498);
nand U2424 (N_2424,In_487,In_431);
and U2425 (N_2425,In_233,In_250);
nand U2426 (N_2426,In_619,In_819);
and U2427 (N_2427,In_535,In_98);
nand U2428 (N_2428,In_45,In_851);
and U2429 (N_2429,In_693,In_634);
and U2430 (N_2430,In_275,In_765);
or U2431 (N_2431,In_847,In_359);
or U2432 (N_2432,In_895,In_292);
nand U2433 (N_2433,In_508,In_51);
or U2434 (N_2434,In_963,In_567);
xnor U2435 (N_2435,In_143,In_206);
xor U2436 (N_2436,In_496,In_271);
nand U2437 (N_2437,In_282,In_322);
nand U2438 (N_2438,In_627,In_575);
nand U2439 (N_2439,In_278,In_619);
nand U2440 (N_2440,In_489,In_845);
nand U2441 (N_2441,In_286,In_786);
or U2442 (N_2442,In_255,In_998);
or U2443 (N_2443,In_366,In_835);
or U2444 (N_2444,In_607,In_997);
and U2445 (N_2445,In_142,In_321);
and U2446 (N_2446,In_318,In_886);
nor U2447 (N_2447,In_216,In_291);
and U2448 (N_2448,In_144,In_64);
nand U2449 (N_2449,In_520,In_122);
nor U2450 (N_2450,In_777,In_918);
and U2451 (N_2451,In_880,In_675);
nand U2452 (N_2452,In_238,In_730);
nand U2453 (N_2453,In_526,In_546);
and U2454 (N_2454,In_792,In_507);
or U2455 (N_2455,In_165,In_573);
nor U2456 (N_2456,In_927,In_908);
nor U2457 (N_2457,In_426,In_562);
nor U2458 (N_2458,In_935,In_886);
or U2459 (N_2459,In_13,In_755);
or U2460 (N_2460,In_129,In_182);
nand U2461 (N_2461,In_887,In_720);
or U2462 (N_2462,In_408,In_448);
or U2463 (N_2463,In_503,In_55);
and U2464 (N_2464,In_213,In_659);
and U2465 (N_2465,In_544,In_252);
nor U2466 (N_2466,In_497,In_923);
or U2467 (N_2467,In_804,In_576);
nor U2468 (N_2468,In_924,In_667);
nor U2469 (N_2469,In_508,In_759);
and U2470 (N_2470,In_159,In_375);
nand U2471 (N_2471,In_426,In_474);
and U2472 (N_2472,In_861,In_435);
nand U2473 (N_2473,In_678,In_819);
and U2474 (N_2474,In_176,In_774);
nand U2475 (N_2475,In_791,In_73);
nand U2476 (N_2476,In_926,In_841);
or U2477 (N_2477,In_908,In_362);
or U2478 (N_2478,In_772,In_919);
and U2479 (N_2479,In_382,In_414);
or U2480 (N_2480,In_778,In_599);
and U2481 (N_2481,In_990,In_244);
or U2482 (N_2482,In_707,In_709);
nand U2483 (N_2483,In_59,In_220);
nor U2484 (N_2484,In_363,In_769);
and U2485 (N_2485,In_88,In_772);
and U2486 (N_2486,In_908,In_355);
xnor U2487 (N_2487,In_876,In_400);
and U2488 (N_2488,In_711,In_57);
and U2489 (N_2489,In_151,In_815);
and U2490 (N_2490,In_645,In_449);
and U2491 (N_2491,In_953,In_774);
or U2492 (N_2492,In_374,In_188);
nand U2493 (N_2493,In_254,In_584);
nor U2494 (N_2494,In_544,In_838);
and U2495 (N_2495,In_936,In_27);
nor U2496 (N_2496,In_316,In_434);
nand U2497 (N_2497,In_118,In_980);
nand U2498 (N_2498,In_383,In_653);
and U2499 (N_2499,In_530,In_280);
or U2500 (N_2500,N_944,N_1310);
and U2501 (N_2501,N_1647,N_502);
and U2502 (N_2502,N_646,N_476);
nand U2503 (N_2503,N_1099,N_1918);
nand U2504 (N_2504,N_1933,N_1235);
and U2505 (N_2505,N_1337,N_1736);
nand U2506 (N_2506,N_2330,N_2213);
nand U2507 (N_2507,N_2272,N_2483);
nand U2508 (N_2508,N_1407,N_1480);
and U2509 (N_2509,N_2306,N_1223);
nand U2510 (N_2510,N_2497,N_330);
or U2511 (N_2511,N_463,N_1590);
or U2512 (N_2512,N_1108,N_131);
or U2513 (N_2513,N_258,N_515);
and U2514 (N_2514,N_1209,N_891);
nand U2515 (N_2515,N_1284,N_1112);
or U2516 (N_2516,N_2311,N_2362);
nand U2517 (N_2517,N_1656,N_2363);
nor U2518 (N_2518,N_1814,N_1988);
nor U2519 (N_2519,N_529,N_2314);
and U2520 (N_2520,N_853,N_435);
or U2521 (N_2521,N_2375,N_2128);
nand U2522 (N_2522,N_1120,N_1174);
nand U2523 (N_2523,N_2287,N_209);
and U2524 (N_2524,N_1558,N_906);
and U2525 (N_2525,N_745,N_554);
or U2526 (N_2526,N_1451,N_2350);
nor U2527 (N_2527,N_1946,N_280);
nand U2528 (N_2528,N_302,N_892);
and U2529 (N_2529,N_1349,N_1793);
nor U2530 (N_2530,N_936,N_367);
or U2531 (N_2531,N_2282,N_14);
nand U2532 (N_2532,N_252,N_1853);
nand U2533 (N_2533,N_2111,N_1963);
nor U2534 (N_2534,N_1043,N_1561);
and U2535 (N_2535,N_2223,N_917);
and U2536 (N_2536,N_1373,N_1138);
or U2537 (N_2537,N_1283,N_378);
nand U2538 (N_2538,N_340,N_632);
or U2539 (N_2539,N_1821,N_911);
nor U2540 (N_2540,N_2388,N_1002);
xnor U2541 (N_2541,N_1828,N_273);
and U2542 (N_2542,N_1471,N_808);
nor U2543 (N_2543,N_1253,N_154);
or U2544 (N_2544,N_2419,N_982);
or U2545 (N_2545,N_348,N_882);
nor U2546 (N_2546,N_1280,N_905);
nor U2547 (N_2547,N_57,N_1484);
nor U2548 (N_2548,N_491,N_2045);
or U2549 (N_2549,N_2087,N_1464);
nand U2550 (N_2550,N_2414,N_2113);
nor U2551 (N_2551,N_2412,N_537);
nor U2552 (N_2552,N_417,N_337);
and U2553 (N_2553,N_2098,N_963);
nand U2554 (N_2554,N_724,N_644);
nor U2555 (N_2555,N_959,N_1585);
nor U2556 (N_2556,N_710,N_188);
nor U2557 (N_2557,N_1629,N_2307);
nand U2558 (N_2558,N_1135,N_2268);
and U2559 (N_2559,N_2329,N_1368);
and U2560 (N_2560,N_1124,N_1431);
nor U2561 (N_2561,N_1939,N_411);
or U2562 (N_2562,N_983,N_2228);
nand U2563 (N_2563,N_689,N_575);
nand U2564 (N_2564,N_1236,N_1808);
nand U2565 (N_2565,N_1667,N_1212);
or U2566 (N_2566,N_1700,N_1718);
and U2567 (N_2567,N_1048,N_2225);
and U2568 (N_2568,N_1723,N_932);
nor U2569 (N_2569,N_1020,N_281);
and U2570 (N_2570,N_1039,N_2477);
and U2571 (N_2571,N_443,N_979);
or U2572 (N_2572,N_2447,N_1579);
or U2573 (N_2573,N_2237,N_1514);
and U2574 (N_2574,N_950,N_759);
nand U2575 (N_2575,N_270,N_940);
and U2576 (N_2576,N_68,N_2031);
nor U2577 (N_2577,N_486,N_1592);
nand U2578 (N_2578,N_1745,N_1444);
nand U2579 (N_2579,N_1887,N_1516);
and U2580 (N_2580,N_2271,N_565);
or U2581 (N_2581,N_1913,N_2364);
nor U2582 (N_2582,N_900,N_432);
or U2583 (N_2583,N_475,N_1547);
or U2584 (N_2584,N_754,N_778);
or U2585 (N_2585,N_2058,N_1684);
or U2586 (N_2586,N_879,N_1565);
and U2587 (N_2587,N_2485,N_1548);
xnor U2588 (N_2588,N_843,N_16);
nand U2589 (N_2589,N_2170,N_1485);
and U2590 (N_2590,N_262,N_223);
or U2591 (N_2591,N_2292,N_2083);
nor U2592 (N_2592,N_2138,N_239);
nor U2593 (N_2593,N_2182,N_1622);
nand U2594 (N_2594,N_1902,N_1080);
nor U2595 (N_2595,N_1178,N_1529);
xor U2596 (N_2596,N_29,N_816);
nor U2597 (N_2597,N_202,N_2298);
nor U2598 (N_2598,N_574,N_288);
and U2599 (N_2599,N_2155,N_1049);
or U2600 (N_2600,N_1783,N_1237);
nor U2601 (N_2601,N_2286,N_647);
nor U2602 (N_2602,N_2246,N_2133);
and U2603 (N_2603,N_1508,N_887);
or U2604 (N_2604,N_2369,N_656);
or U2605 (N_2605,N_1405,N_898);
nor U2606 (N_2606,N_981,N_1299);
nand U2607 (N_2607,N_1470,N_517);
or U2608 (N_2608,N_914,N_1551);
nand U2609 (N_2609,N_572,N_1510);
or U2610 (N_2610,N_445,N_1996);
nand U2611 (N_2611,N_1060,N_2255);
and U2612 (N_2612,N_1006,N_229);
nor U2613 (N_2613,N_2366,N_987);
nor U2614 (N_2614,N_777,N_277);
or U2615 (N_2615,N_1317,N_2227);
nor U2616 (N_2616,N_2251,N_1136);
nand U2617 (N_2617,N_1232,N_649);
nor U2618 (N_2618,N_1104,N_1445);
nor U2619 (N_2619,N_811,N_929);
and U2620 (N_2620,N_1696,N_2168);
nor U2621 (N_2621,N_1570,N_1193);
or U2622 (N_2622,N_79,N_850);
and U2623 (N_2623,N_380,N_1780);
and U2624 (N_2624,N_1642,N_192);
or U2625 (N_2625,N_1705,N_1742);
nand U2626 (N_2626,N_551,N_2498);
nand U2627 (N_2627,N_1482,N_263);
and U2628 (N_2628,N_2342,N_1838);
and U2629 (N_2629,N_1084,N_1989);
nand U2630 (N_2630,N_2095,N_1533);
or U2631 (N_2631,N_2029,N_1532);
xor U2632 (N_2632,N_345,N_1526);
nor U2633 (N_2633,N_1359,N_2124);
and U2634 (N_2634,N_1459,N_1897);
nor U2635 (N_2635,N_1074,N_1129);
nor U2636 (N_2636,N_2266,N_2065);
nor U2637 (N_2637,N_1406,N_47);
nor U2638 (N_2638,N_2037,N_538);
and U2639 (N_2639,N_719,N_1151);
nor U2640 (N_2640,N_919,N_1936);
and U2641 (N_2641,N_424,N_1870);
and U2642 (N_2642,N_1574,N_327);
nand U2643 (N_2643,N_1216,N_878);
and U2644 (N_2644,N_254,N_561);
or U2645 (N_2645,N_21,N_751);
nor U2646 (N_2646,N_827,N_420);
nor U2647 (N_2647,N_2269,N_324);
and U2648 (N_2648,N_138,N_611);
or U2649 (N_2649,N_1382,N_183);
and U2650 (N_2650,N_323,N_98);
and U2651 (N_2651,N_1673,N_2121);
and U2652 (N_2652,N_2338,N_189);
nor U2653 (N_2653,N_592,N_531);
nor U2654 (N_2654,N_2318,N_1586);
and U2655 (N_2655,N_2204,N_361);
or U2656 (N_2656,N_1664,N_809);
and U2657 (N_2657,N_2231,N_795);
nand U2658 (N_2658,N_1844,N_396);
nor U2659 (N_2659,N_266,N_1441);
nor U2660 (N_2660,N_2354,N_2208);
nor U2661 (N_2661,N_1949,N_530);
and U2662 (N_2662,N_688,N_1982);
and U2663 (N_2663,N_899,N_1994);
nand U2664 (N_2664,N_1365,N_1820);
nand U2665 (N_2665,N_1638,N_2226);
or U2666 (N_2666,N_510,N_563);
xnor U2667 (N_2667,N_556,N_526);
nand U2668 (N_2668,N_2179,N_993);
and U2669 (N_2669,N_523,N_1677);
nor U2670 (N_2670,N_506,N_2091);
or U2671 (N_2671,N_1334,N_1383);
and U2672 (N_2672,N_1442,N_1955);
and U2673 (N_2673,N_1619,N_279);
nor U2674 (N_2674,N_1313,N_623);
or U2675 (N_2675,N_2382,N_1720);
nor U2676 (N_2676,N_1220,N_1785);
or U2677 (N_2677,N_86,N_1879);
and U2678 (N_2678,N_1331,N_1651);
or U2679 (N_2679,N_548,N_888);
nor U2680 (N_2680,N_2108,N_824);
and U2681 (N_2681,N_1623,N_326);
nor U2682 (N_2682,N_1266,N_1967);
and U2683 (N_2683,N_19,N_375);
nor U2684 (N_2684,N_1908,N_1273);
or U2685 (N_2685,N_127,N_1324);
or U2686 (N_2686,N_392,N_615);
nand U2687 (N_2687,N_2460,N_1865);
nor U2688 (N_2688,N_1242,N_473);
and U2689 (N_2689,N_37,N_1378);
nor U2690 (N_2690,N_1633,N_1554);
and U2691 (N_2691,N_1875,N_699);
or U2692 (N_2692,N_438,N_143);
nand U2693 (N_2693,N_1974,N_1631);
nor U2694 (N_2694,N_1356,N_139);
nand U2695 (N_2695,N_325,N_2118);
nand U2696 (N_2696,N_2149,N_184);
or U2697 (N_2697,N_663,N_2156);
and U2698 (N_2698,N_756,N_1764);
or U2699 (N_2699,N_1077,N_1542);
or U2700 (N_2700,N_331,N_691);
nand U2701 (N_2701,N_1852,N_1671);
xor U2702 (N_2702,N_175,N_297);
nand U2703 (N_2703,N_1096,N_815);
or U2704 (N_2704,N_2391,N_1265);
and U2705 (N_2705,N_339,N_1797);
and U2706 (N_2706,N_2333,N_1917);
nor U2707 (N_2707,N_1916,N_1371);
nor U2708 (N_2708,N_2064,N_1122);
or U2709 (N_2709,N_2006,N_558);
nand U2710 (N_2710,N_1610,N_149);
and U2711 (N_2711,N_2401,N_1860);
nor U2712 (N_2712,N_2034,N_49);
nand U2713 (N_2713,N_1961,N_1704);
nand U2714 (N_2714,N_772,N_314);
and U2715 (N_2715,N_484,N_187);
nor U2716 (N_2716,N_249,N_1017);
or U2717 (N_2717,N_2267,N_2275);
nand U2718 (N_2718,N_1257,N_419);
or U2719 (N_2719,N_798,N_2043);
and U2720 (N_2720,N_2184,N_1707);
or U2721 (N_2721,N_2476,N_1211);
nor U2722 (N_2722,N_671,N_1630);
and U2723 (N_2723,N_382,N_2377);
nand U2724 (N_2724,N_1244,N_871);
nand U2725 (N_2725,N_1507,N_2056);
nor U2726 (N_2726,N_673,N_557);
nand U2727 (N_2727,N_110,N_1737);
nand U2728 (N_2728,N_1411,N_472);
or U2729 (N_2729,N_594,N_1463);
nor U2730 (N_2730,N_1263,N_2464);
nor U2731 (N_2731,N_1909,N_43);
and U2732 (N_2732,N_122,N_434);
nand U2733 (N_2733,N_525,N_2187);
nand U2734 (N_2734,N_24,N_1825);
nor U2735 (N_2735,N_2063,N_1493);
or U2736 (N_2736,N_2478,N_2299);
nor U2737 (N_2737,N_1256,N_1749);
nand U2738 (N_2738,N_1247,N_1403);
or U2739 (N_2739,N_1952,N_2459);
nor U2740 (N_2740,N_1271,N_825);
nand U2741 (N_2741,N_991,N_1027);
nand U2742 (N_2742,N_1605,N_1474);
nor U2743 (N_2743,N_1338,N_1566);
or U2744 (N_2744,N_1032,N_2067);
nor U2745 (N_2745,N_1289,N_1162);
nor U2746 (N_2746,N_407,N_567);
or U2747 (N_2747,N_1008,N_305);
or U2748 (N_2748,N_489,N_1187);
nor U2749 (N_2749,N_1396,N_1744);
or U2750 (N_2750,N_568,N_1986);
nor U2751 (N_2751,N_95,N_121);
nand U2752 (N_2752,N_1550,N_1709);
nor U2753 (N_2753,N_915,N_1168);
and U2754 (N_2754,N_2172,N_790);
nor U2755 (N_2755,N_528,N_2461);
nand U2756 (N_2756,N_1342,N_294);
and U2757 (N_2757,N_2305,N_2499);
and U2758 (N_2758,N_1130,N_2046);
nor U2759 (N_2759,N_863,N_655);
xnor U2760 (N_2760,N_22,N_2310);
and U2761 (N_2761,N_1859,N_2047);
nand U2762 (N_2762,N_1819,N_1119);
or U2763 (N_2763,N_1221,N_2159);
nand U2764 (N_2764,N_2254,N_383);
and U2765 (N_2765,N_1386,N_2468);
nor U2766 (N_2766,N_1758,N_1056);
nor U2767 (N_2767,N_1454,N_666);
nor U2768 (N_2768,N_821,N_1259);
nand U2769 (N_2769,N_1345,N_2163);
nand U2770 (N_2770,N_1275,N_684);
nor U2771 (N_2771,N_2007,N_1456);
nor U2772 (N_2772,N_350,N_500);
and U2773 (N_2773,N_1302,N_2290);
or U2774 (N_2774,N_69,N_487);
or U2775 (N_2775,N_1213,N_573);
xor U2776 (N_2776,N_217,N_2044);
nand U2777 (N_2777,N_1966,N_1419);
nand U2778 (N_2778,N_2066,N_231);
and U2779 (N_2779,N_1695,N_749);
nand U2780 (N_2780,N_1895,N_2378);
and U2781 (N_2781,N_757,N_1429);
or U2782 (N_2782,N_2090,N_0);
xnor U2783 (N_2783,N_1701,N_837);
nor U2784 (N_2784,N_1766,N_1360);
nand U2785 (N_2785,N_2482,N_1117);
xor U2786 (N_2786,N_1327,N_1457);
or U2787 (N_2787,N_780,N_1890);
nand U2788 (N_2788,N_2001,N_1960);
nand U2789 (N_2789,N_730,N_1079);
nor U2790 (N_2790,N_1069,N_1231);
and U2791 (N_2791,N_1513,N_2114);
nor U2792 (N_2792,N_2315,N_159);
and U2793 (N_2793,N_1922,N_842);
nor U2794 (N_2794,N_2371,N_471);
or U2795 (N_2795,N_2434,N_2014);
nor U2796 (N_2796,N_1931,N_2181);
and U2797 (N_2797,N_1904,N_1925);
and U2798 (N_2798,N_953,N_2220);
nor U2799 (N_2799,N_1277,N_1479);
nor U2800 (N_2800,N_2196,N_61);
nand U2801 (N_2801,N_2348,N_2028);
or U2802 (N_2802,N_1267,N_653);
and U2803 (N_2803,N_627,N_2178);
or U2804 (N_2804,N_716,N_354);
nor U2805 (N_2805,N_1976,N_1401);
or U2806 (N_2806,N_2384,N_507);
or U2807 (N_2807,N_896,N_1617);
nor U2808 (N_2808,N_1580,N_1665);
nor U2809 (N_2809,N_576,N_633);
nand U2810 (N_2810,N_26,N_264);
and U2811 (N_2811,N_614,N_388);
and U2812 (N_2812,N_1173,N_977);
nor U2813 (N_2813,N_2245,N_715);
and U2814 (N_2814,N_1741,N_1735);
nor U2815 (N_2815,N_2444,N_964);
nor U2816 (N_2816,N_315,N_2200);
and U2817 (N_2817,N_2157,N_2092);
or U2818 (N_2818,N_1408,N_1078);
nor U2819 (N_2819,N_714,N_481);
nand U2820 (N_2820,N_233,N_758);
or U2821 (N_2821,N_137,N_1523);
or U2822 (N_2822,N_1274,N_2381);
nand U2823 (N_2823,N_146,N_1927);
or U2824 (N_2824,N_2142,N_775);
nor U2825 (N_2825,N_1544,N_660);
nand U2826 (N_2826,N_2230,N_1815);
nand U2827 (N_2827,N_1702,N_398);
nand U2828 (N_2828,N_1873,N_50);
and U2829 (N_2829,N_616,N_678);
nor U2830 (N_2830,N_2012,N_2295);
nand U2831 (N_2831,N_120,N_1295);
nand U2832 (N_2832,N_519,N_482);
or U2833 (N_2833,N_1082,N_1649);
or U2834 (N_2834,N_1358,N_1447);
nor U2835 (N_2835,N_1298,N_28);
nor U2836 (N_2836,N_74,N_841);
or U2837 (N_2837,N_1553,N_1826);
nand U2838 (N_2838,N_1863,N_358);
nand U2839 (N_2839,N_1330,N_1738);
nor U2840 (N_2840,N_1596,N_694);
or U2841 (N_2841,N_2015,N_789);
nand U2842 (N_2842,N_1545,N_930);
and U2843 (N_2843,N_1321,N_1912);
and U2844 (N_2844,N_776,N_1781);
nor U2845 (N_2845,N_1061,N_2242);
nor U2846 (N_2846,N_2036,N_2259);
nor U2847 (N_2847,N_301,N_1968);
and U2848 (N_2848,N_1070,N_124);
nand U2849 (N_2849,N_1653,N_1498);
and U2850 (N_2850,N_520,N_2248);
nand U2851 (N_2851,N_767,N_640);
and U2852 (N_2852,N_1142,N_590);
nor U2853 (N_2853,N_718,N_2300);
nand U2854 (N_2854,N_588,N_1503);
nand U2855 (N_2855,N_499,N_2235);
xor U2856 (N_2856,N_353,N_2039);
or U2857 (N_2857,N_559,N_620);
or U2858 (N_2858,N_211,N_478);
and U2859 (N_2859,N_2402,N_2211);
or U2860 (N_2860,N_1789,N_13);
or U2861 (N_2861,N_2308,N_117);
or U2862 (N_2862,N_144,N_241);
or U2863 (N_2863,N_1595,N_1455);
or U2864 (N_2864,N_2440,N_1387);
nand U2865 (N_2865,N_2293,N_669);
or U2866 (N_2866,N_785,N_1756);
nor U2867 (N_2867,N_511,N_185);
nand U2868 (N_2868,N_1620,N_30);
or U2869 (N_2869,N_1206,N_1941);
and U2870 (N_2870,N_1800,N_2);
and U2871 (N_2871,N_2408,N_916);
nand U2872 (N_2872,N_1492,N_1995);
nand U2873 (N_2873,N_1971,N_861);
or U2874 (N_2874,N_1903,N_158);
or U2875 (N_2875,N_1593,N_2038);
or U2876 (N_2876,N_1834,N_338);
nand U2877 (N_2877,N_2343,N_849);
nor U2878 (N_2878,N_521,N_1164);
nor U2879 (N_2879,N_1101,N_908);
nor U2880 (N_2880,N_1991,N_2449);
nand U2881 (N_2881,N_1727,N_1448);
and U2882 (N_2882,N_1843,N_114);
nand U2883 (N_2883,N_2262,N_1752);
and U2884 (N_2884,N_2010,N_368);
and U2885 (N_2885,N_1443,N_958);
or U2886 (N_2886,N_729,N_2035);
nand U2887 (N_2887,N_1868,N_1589);
and U2888 (N_2888,N_2099,N_94);
and U2889 (N_2889,N_1639,N_140);
nor U2890 (N_2890,N_2016,N_831);
nor U2891 (N_2891,N_1353,N_1948);
nand U2892 (N_2892,N_1179,N_1849);
nand U2893 (N_2893,N_587,N_935);
or U2894 (N_2894,N_243,N_1978);
nand U2895 (N_2895,N_1940,N_1050);
nand U2896 (N_2896,N_109,N_1753);
and U2897 (N_2897,N_1979,N_840);
nand U2898 (N_2898,N_836,N_852);
nor U2899 (N_2899,N_1509,N_2026);
or U2900 (N_2900,N_226,N_477);
nor U2901 (N_2901,N_1290,N_308);
or U2902 (N_2902,N_1708,N_1817);
and U2903 (N_2903,N_2054,N_1921);
nor U2904 (N_2904,N_2152,N_2337);
xnor U2905 (N_2905,N_2158,N_613);
nor U2906 (N_2906,N_133,N_2078);
or U2907 (N_2907,N_1641,N_583);
nand U2908 (N_2908,N_490,N_2340);
and U2909 (N_2909,N_413,N_404);
or U2910 (N_2910,N_384,N_1427);
nor U2911 (N_2911,N_2024,N_429);
nor U2912 (N_2912,N_1261,N_1021);
or U2913 (N_2913,N_1341,N_251);
nor U2914 (N_2914,N_1739,N_2392);
nor U2915 (N_2915,N_503,N_1367);
nand U2916 (N_2916,N_954,N_1822);
or U2917 (N_2917,N_1538,N_1010);
nor U2918 (N_2918,N_1228,N_1248);
or U2919 (N_2919,N_35,N_479);
nand U2920 (N_2920,N_1915,N_1381);
nor U2921 (N_2921,N_926,N_1306);
and U2922 (N_2922,N_1473,N_459);
nor U2923 (N_2923,N_1732,N_924);
nand U2924 (N_2924,N_1856,N_943);
and U2925 (N_2925,N_1877,N_844);
nor U2926 (N_2926,N_1316,N_2352);
xnor U2927 (N_2927,N_450,N_1567);
and U2928 (N_2928,N_1972,N_1659);
nand U2929 (N_2929,N_1197,N_1461);
xnor U2930 (N_2930,N_1252,N_341);
nand U2931 (N_2931,N_1399,N_2373);
nor U2932 (N_2932,N_464,N_970);
and U2933 (N_2933,N_2471,N_2474);
nand U2934 (N_2934,N_1827,N_2367);
nor U2935 (N_2935,N_379,N_1790);
or U2936 (N_2936,N_2359,N_1878);
or U2937 (N_2937,N_1900,N_1336);
nand U2938 (N_2938,N_2465,N_365);
or U2939 (N_2939,N_1024,N_1158);
and U2940 (N_2940,N_1869,N_2263);
nand U2941 (N_2941,N_976,N_2202);
and U2942 (N_2942,N_1970,N_1160);
nand U2943 (N_2943,N_820,N_71);
nor U2944 (N_2944,N_11,N_769);
and U2945 (N_2945,N_2385,N_2103);
nand U2946 (N_2946,N_2379,N_2195);
and U2947 (N_2947,N_1140,N_135);
nand U2948 (N_2948,N_1133,N_2407);
and U2949 (N_2949,N_1087,N_408);
nand U2950 (N_2950,N_1706,N_693);
nor U2951 (N_2951,N_941,N_1392);
nand U2952 (N_2952,N_171,N_89);
or U2953 (N_2953,N_300,N_2102);
and U2954 (N_2954,N_1249,N_1929);
and U2955 (N_2955,N_664,N_1214);
or U2956 (N_2956,N_97,N_1219);
nor U2957 (N_2957,N_234,N_635);
and U2958 (N_2958,N_46,N_64);
xor U2959 (N_2959,N_1740,N_593);
or U2960 (N_2960,N_247,N_157);
or U2961 (N_2961,N_81,N_578);
and U2962 (N_2962,N_762,N_1395);
nand U2963 (N_2963,N_224,N_359);
and U2964 (N_2964,N_1618,N_322);
nand U2965 (N_2965,N_2361,N_598);
and U2966 (N_2966,N_1511,N_2301);
nor U2967 (N_2967,N_717,N_451);
or U2968 (N_2968,N_2284,N_1530);
nand U2969 (N_2969,N_695,N_1420);
nand U2970 (N_2970,N_1572,N_1291);
and U2971 (N_2971,N_2424,N_961);
nor U2972 (N_2972,N_2072,N_2473);
nand U2973 (N_2973,N_1009,N_1711);
nand U2974 (N_2974,N_999,N_1292);
nor U2975 (N_2975,N_641,N_1985);
or U2976 (N_2976,N_518,N_2140);
nand U2977 (N_2977,N_807,N_1475);
or U2978 (N_2978,N_2396,N_134);
nand U2979 (N_2979,N_2429,N_1217);
nand U2980 (N_2980,N_2096,N_501);
nor U2981 (N_2981,N_989,N_1478);
or U2982 (N_2982,N_1486,N_1015);
and U2983 (N_2983,N_1577,N_1721);
or U2984 (N_2984,N_681,N_208);
and U2985 (N_2985,N_1757,N_1222);
or U2986 (N_2986,N_1801,N_465);
or U2987 (N_2987,N_51,N_351);
and U2988 (N_2988,N_1460,N_768);
nor U2989 (N_2989,N_283,N_2252);
or U2990 (N_2990,N_442,N_33);
xnor U2991 (N_2991,N_53,N_453);
nor U2992 (N_2992,N_357,N_2349);
xnor U2993 (N_2993,N_2319,N_1500);
nor U2994 (N_2994,N_1624,N_744);
nand U2995 (N_2995,N_1597,N_320);
nor U2996 (N_2996,N_921,N_1685);
and U2997 (N_2997,N_458,N_182);
nand U2998 (N_2998,N_8,N_2051);
and U2999 (N_2999,N_1393,N_618);
nand U3000 (N_3000,N_1835,N_1147);
nor U3001 (N_3001,N_1030,N_2475);
and U3002 (N_3002,N_712,N_1855);
nand U3003 (N_3003,N_1811,N_2085);
nand U3004 (N_3004,N_2285,N_2126);
and U3005 (N_3005,N_1172,N_1230);
or U3006 (N_3006,N_237,N_1033);
nand U3007 (N_3007,N_1943,N_103);
or U3008 (N_3008,N_1073,N_723);
nor U3009 (N_3009,N_60,N_2280);
nand U3010 (N_3010,N_260,N_2233);
and U3011 (N_3011,N_130,N_433);
and U3012 (N_3012,N_1866,N_1052);
or U3013 (N_3013,N_1688,N_1525);
and U3014 (N_3014,N_610,N_1805);
nor U3015 (N_3015,N_1458,N_734);
or U3016 (N_3016,N_1376,N_832);
nand U3017 (N_3017,N_2166,N_1575);
and U3018 (N_3018,N_1023,N_148);
and U3019 (N_3019,N_2042,N_771);
and U3020 (N_3020,N_2456,N_441);
or U3021 (N_3021,N_1697,N_48);
xor U3022 (N_3022,N_1759,N_2049);
nand U3023 (N_3023,N_1152,N_910);
nand U3024 (N_3024,N_676,N_1011);
nor U3025 (N_3025,N_1568,N_998);
nand U3026 (N_3026,N_126,N_494);
nor U3027 (N_3027,N_1145,N_1415);
nor U3028 (N_3028,N_731,N_2416);
nor U3029 (N_3029,N_642,N_430);
or U3030 (N_3030,N_2344,N_2372);
and U3031 (N_3031,N_643,N_2404);
nand U3032 (N_3032,N_316,N_55);
and U3033 (N_3033,N_1107,N_282);
or U3034 (N_3034,N_9,N_1307);
nand U3035 (N_3035,N_2450,N_2079);
nand U3036 (N_3036,N_2134,N_697);
nor U3037 (N_3037,N_176,N_2232);
and U3038 (N_3038,N_1932,N_2169);
and U3039 (N_3039,N_569,N_738);
and U3040 (N_3040,N_1086,N_980);
or U3041 (N_3041,N_662,N_1446);
nand U3042 (N_3042,N_1733,N_2281);
nand U3043 (N_3043,N_1830,N_1799);
and U3044 (N_3044,N_612,N_2486);
nor U3045 (N_3045,N_621,N_1874);
and U3046 (N_3046,N_2145,N_77);
and U3047 (N_3047,N_709,N_1973);
or U3048 (N_3048,N_2164,N_1362);
and U3049 (N_3049,N_603,N_740);
or U3050 (N_3050,N_1121,N_1449);
or U3051 (N_3051,N_1300,N_2432);
and U3052 (N_3052,N_819,N_2304);
nand U3053 (N_3053,N_372,N_2057);
and U3054 (N_3054,N_1260,N_2445);
nor U3055 (N_3055,N_2125,N_1784);
nand U3056 (N_3056,N_1689,N_1886);
or U3057 (N_3057,N_1541,N_1176);
nand U3058 (N_3058,N_1926,N_1404);
nand U3059 (N_3059,N_792,N_604);
nor U3060 (N_3060,N_1848,N_2480);
and U3061 (N_3061,N_406,N_2141);
or U3062 (N_3062,N_947,N_1388);
or U3063 (N_3063,N_1934,N_2283);
or U3064 (N_3064,N_457,N_1661);
or U3065 (N_3065,N_1776,N_1036);
or U3066 (N_3066,N_2457,N_1831);
and U3067 (N_3067,N_645,N_205);
and U3068 (N_3068,N_2019,N_1803);
or U3069 (N_3069,N_1177,N_75);
nor U3070 (N_3070,N_1964,N_160);
or U3071 (N_3071,N_774,N_232);
nand U3072 (N_3072,N_100,N_1045);
nor U3073 (N_3073,N_2188,N_978);
nor U3074 (N_3074,N_1004,N_1518);
or U3075 (N_3075,N_363,N_42);
nand U3076 (N_3076,N_1901,N_395);
xor U3077 (N_3077,N_468,N_680);
nand U3078 (N_3078,N_1774,N_2229);
and U3079 (N_3079,N_1847,N_692);
or U3080 (N_3080,N_674,N_2020);
nand U3081 (N_3081,N_1636,N_85);
or U3082 (N_3082,N_736,N_894);
nor U3083 (N_3083,N_1535,N_151);
nand U3084 (N_3084,N_562,N_440);
nand U3085 (N_3085,N_311,N_955);
and U3086 (N_3086,N_230,N_2214);
xnor U3087 (N_3087,N_2219,N_760);
nor U3088 (N_3088,N_2376,N_711);
nor U3089 (N_3089,N_1771,N_1881);
nand U3090 (N_3090,N_1314,N_1604);
xnor U3091 (N_3091,N_1106,N_2277);
and U3092 (N_3092,N_752,N_1258);
nand U3093 (N_3093,N_1889,N_1938);
nor U3094 (N_3094,N_788,N_2455);
or U3095 (N_3095,N_1131,N_342);
or U3096 (N_3096,N_918,N_1218);
and U3097 (N_3097,N_1515,N_737);
nor U3098 (N_3098,N_1188,N_2186);
nand U3099 (N_3099,N_755,N_1522);
and U3100 (N_3100,N_1462,N_1992);
nor U3101 (N_3101,N_1693,N_2481);
or U3102 (N_3102,N_257,N_2139);
nor U3103 (N_3103,N_2041,N_427);
and U3104 (N_3104,N_2100,N_2173);
nand U3105 (N_3105,N_2191,N_2109);
or U3106 (N_3106,N_1416,N_893);
nor U3107 (N_3107,N_1601,N_1680);
nand U3108 (N_3108,N_1180,N_1326);
and U3109 (N_3109,N_2466,N_748);
or U3110 (N_3110,N_626,N_707);
and U3111 (N_3111,N_1722,N_220);
and U3112 (N_3112,N_1846,N_942);
nand U3113 (N_3113,N_560,N_1016);
or U3114 (N_3114,N_512,N_2217);
nor U3115 (N_3115,N_1224,N_1208);
or U3116 (N_3116,N_1001,N_2331);
nor U3117 (N_3117,N_1323,N_966);
nand U3118 (N_3118,N_431,N_397);
nor U3119 (N_3119,N_1748,N_1402);
nand U3120 (N_3120,N_2040,N_1380);
or U3121 (N_3121,N_2296,N_974);
nand U3122 (N_3122,N_497,N_474);
or U3123 (N_3123,N_2291,N_1777);
or U3124 (N_3124,N_3,N_225);
nand U3125 (N_3125,N_992,N_2303);
and U3126 (N_3126,N_2433,N_88);
or U3127 (N_3127,N_2129,N_82);
and U3128 (N_3128,N_1937,N_1872);
nand U3129 (N_3129,N_1433,N_1468);
nor U3130 (N_3130,N_58,N_1864);
or U3131 (N_3131,N_2358,N_1672);
nand U3132 (N_3132,N_829,N_456);
and U3133 (N_3133,N_261,N_1896);
or U3134 (N_3134,N_1318,N_483);
and U3135 (N_3135,N_813,N_199);
nand U3136 (N_3136,N_377,N_1159);
or U3137 (N_3137,N_1254,N_1229);
nor U3138 (N_3138,N_1730,N_248);
and U3139 (N_3139,N_2397,N_245);
or U3140 (N_3140,N_67,N_1987);
and U3141 (N_3141,N_2194,N_1312);
nand U3142 (N_3142,N_2062,N_885);
or U3143 (N_3143,N_389,N_1576);
nand U3144 (N_3144,N_1662,N_1582);
nor U3145 (N_3145,N_1778,N_1578);
and U3146 (N_3146,N_739,N_72);
or U3147 (N_3147,N_1655,N_1348);
or U3148 (N_3148,N_1240,N_1663);
nand U3149 (N_3149,N_786,N_2205);
nand U3150 (N_3150,N_2294,N_1612);
nand U3151 (N_3151,N_968,N_606);
and U3152 (N_3152,N_259,N_371);
nand U3153 (N_3153,N_883,N_32);
nand U3154 (N_3154,N_796,N_54);
and U3155 (N_3155,N_2197,N_2069);
nor U3156 (N_3156,N_884,N_1694);
nand U3157 (N_3157,N_31,N_10);
nor U3158 (N_3158,N_2430,N_2274);
nand U3159 (N_3159,N_838,N_1196);
or U3160 (N_3160,N_1957,N_1779);
or U3161 (N_3161,N_2070,N_508);
nand U3162 (N_3162,N_129,N_939);
and U3163 (N_3163,N_1414,N_638);
nand U3164 (N_3164,N_364,N_1947);
and U3165 (N_3165,N_1022,N_2398);
nand U3166 (N_3166,N_2161,N_2410);
nor U3167 (N_3167,N_833,N_2004);
or U3168 (N_3168,N_101,N_952);
nand U3169 (N_3169,N_1998,N_1374);
and U3170 (N_3170,N_1066,N_125);
nor U3171 (N_3171,N_190,N_65);
nand U3172 (N_3172,N_912,N_1625);
nor U3173 (N_3173,N_1981,N_1198);
or U3174 (N_3174,N_1207,N_96);
or U3175 (N_3175,N_984,N_2399);
or U3176 (N_3176,N_422,N_390);
nand U3177 (N_3177,N_448,N_927);
and U3178 (N_3178,N_988,N_1425);
nor U3179 (N_3179,N_2077,N_1329);
or U3180 (N_3180,N_1763,N_460);
nor U3181 (N_3181,N_1435,N_2446);
or U3182 (N_3182,N_265,N_2346);
nor U3183 (N_3183,N_274,N_2221);
nor U3184 (N_3184,N_99,N_1905);
nand U3185 (N_3185,N_1891,N_1608);
nand U3186 (N_3186,N_228,N_416);
and U3187 (N_3187,N_349,N_1114);
or U3188 (N_3188,N_931,N_2167);
or U3189 (N_3189,N_2258,N_1286);
nand U3190 (N_3190,N_200,N_2151);
and U3191 (N_3191,N_216,N_2413);
nand U3192 (N_3192,N_386,N_1089);
nand U3193 (N_3193,N_2425,N_1282);
nand U3194 (N_3194,N_1363,N_466);
nand U3195 (N_3195,N_1226,N_957);
nor U3196 (N_3196,N_41,N_1432);
nand U3197 (N_3197,N_535,N_179);
or U3198 (N_3198,N_1189,N_1144);
nand U3199 (N_3199,N_91,N_1543);
and U3200 (N_3200,N_2052,N_928);
nor U3201 (N_3201,N_1370,N_1311);
nor U3202 (N_3202,N_447,N_668);
and U3203 (N_3203,N_240,N_1132);
or U3204 (N_3204,N_193,N_1268);
nand U3205 (N_3205,N_112,N_2084);
and U3206 (N_3206,N_1,N_394);
and U3207 (N_3207,N_875,N_1203);
nor U3208 (N_3208,N_2018,N_960);
nand U3209 (N_3209,N_802,N_1339);
nor U3210 (N_3210,N_197,N_2177);
and U3211 (N_3211,N_634,N_1372);
nand U3212 (N_3212,N_761,N_312);
or U3213 (N_3213,N_177,N_2316);
and U3214 (N_3214,N_2198,N_2143);
nor U3215 (N_3215,N_446,N_1666);
nor U3216 (N_3216,N_405,N_2059);
or U3217 (N_3217,N_309,N_972);
or U3218 (N_3218,N_59,N_1417);
and U3219 (N_3219,N_1375,N_1304);
nor U3220 (N_3220,N_2312,N_799);
nor U3221 (N_3221,N_191,N_1424);
nand U3222 (N_3222,N_1717,N_306);
nor U3223 (N_3223,N_1528,N_1481);
nor U3224 (N_3224,N_180,N_461);
or U3225 (N_3225,N_1440,N_2148);
nor U3226 (N_3226,N_945,N_544);
nand U3227 (N_3227,N_1840,N_1186);
and U3228 (N_3228,N_401,N_728);
and U3229 (N_3229,N_1888,N_2288);
nand U3230 (N_3230,N_2276,N_269);
or U3231 (N_3231,N_423,N_412);
and U3232 (N_3232,N_235,N_2247);
and U3233 (N_3233,N_687,N_295);
nor U3234 (N_3234,N_2320,N_1692);
nor U3235 (N_3235,N_2150,N_1762);
and U3236 (N_3236,N_2190,N_690);
xor U3237 (N_3237,N_2009,N_2302);
and U3238 (N_3238,N_470,N_246);
and U3239 (N_3239,N_1190,N_1562);
or U3240 (N_3240,N_1340,N_1149);
nand U3241 (N_3241,N_40,N_2206);
and U3242 (N_3242,N_1942,N_2409);
and U3243 (N_3243,N_132,N_1113);
and U3244 (N_3244,N_1430,N_1269);
nand U3245 (N_3245,N_1687,N_2176);
or U3246 (N_3246,N_168,N_1488);
nand U3247 (N_3247,N_2005,N_344);
nand U3248 (N_3248,N_857,N_1426);
nand U3249 (N_3249,N_1731,N_1679);
xor U3250 (N_3250,N_1495,N_1761);
nor U3251 (N_3251,N_858,N_1320);
or U3252 (N_3252,N_889,N_1650);
nand U3253 (N_3253,N_2406,N_80);
nand U3254 (N_3254,N_1491,N_1239);
or U3255 (N_3255,N_570,N_2132);
nor U3256 (N_3256,N_206,N_2115);
and U3257 (N_3257,N_584,N_600);
nor U3258 (N_3258,N_848,N_381);
or U3259 (N_3259,N_648,N_509);
or U3260 (N_3260,N_1100,N_1109);
or U3261 (N_3261,N_1288,N_128);
nand U3262 (N_3262,N_162,N_1907);
or U3263 (N_3263,N_436,N_2313);
nand U3264 (N_3264,N_155,N_1128);
nor U3265 (N_3265,N_514,N_1308);
and U3266 (N_3266,N_2356,N_2403);
nor U3267 (N_3267,N_93,N_823);
nor U3268 (N_3268,N_1072,N_2193);
nand U3269 (N_3269,N_946,N_343);
nor U3270 (N_3270,N_753,N_1075);
nor U3271 (N_3271,N_1366,N_2309);
nor U3272 (N_3272,N_2105,N_1775);
or U3273 (N_3273,N_1675,N_2355);
or U3274 (N_3274,N_1686,N_174);
or U3275 (N_3275,N_1281,N_2492);
or U3276 (N_3276,N_2345,N_854);
nor U3277 (N_3277,N_1657,N_45);
and U3278 (N_3278,N_352,N_2487);
and U3279 (N_3279,N_696,N_1573);
and U3280 (N_3280,N_659,N_1713);
xnor U3281 (N_3281,N_1914,N_1806);
nor U3282 (N_3282,N_564,N_868);
and U3283 (N_3283,N_683,N_1436);
or U3284 (N_3284,N_161,N_539);
nor U3285 (N_3285,N_1614,N_1270);
nor U3286 (N_3286,N_741,N_2462);
or U3287 (N_3287,N_872,N_1110);
nand U3288 (N_3288,N_369,N_18);
and U3289 (N_3289,N_864,N_1127);
nand U3290 (N_3290,N_2289,N_1726);
and U3291 (N_3291,N_356,N_1081);
or U3292 (N_3292,N_855,N_1531);
or U3293 (N_3293,N_493,N_360);
or U3294 (N_3294,N_846,N_1105);
nand U3295 (N_3295,N_1837,N_421);
nand U3296 (N_3296,N_742,N_1858);
or U3297 (N_3297,N_904,N_1555);
or U3298 (N_3298,N_1769,N_1984);
nand U3299 (N_3299,N_1534,N_1691);
nand U3300 (N_3300,N_1928,N_543);
nand U3301 (N_3301,N_1143,N_402);
and U3302 (N_3302,N_704,N_1598);
and U3303 (N_3303,N_851,N_1357);
and U3304 (N_3304,N_218,N_975);
nor U3305 (N_3305,N_391,N_2008);
nor U3306 (N_3306,N_902,N_1626);
or U3307 (N_3307,N_1071,N_907);
nand U3308 (N_3308,N_1734,N_2467);
nand U3309 (N_3309,N_1681,N_36);
nor U3310 (N_3310,N_585,N_1836);
nor U3311 (N_3311,N_2199,N_1031);
and U3312 (N_3312,N_1450,N_1674);
nor U3313 (N_3313,N_1611,N_1139);
nor U3314 (N_3314,N_1116,N_1502);
and U3315 (N_3315,N_1951,N_1569);
or U3316 (N_3316,N_835,N_39);
nor U3317 (N_3317,N_1898,N_1088);
and U3318 (N_3318,N_2427,N_142);
nand U3319 (N_3319,N_803,N_2463);
nor U3320 (N_3320,N_1581,N_2147);
or U3321 (N_3321,N_867,N_1093);
nand U3322 (N_3322,N_213,N_1871);
and U3323 (N_3323,N_1094,N_1754);
and U3324 (N_3324,N_1710,N_1169);
nand U3325 (N_3325,N_2144,N_1658);
nor U3326 (N_3326,N_886,N_2165);
or U3327 (N_3327,N_682,N_504);
or U3328 (N_3328,N_1791,N_1309);
and U3329 (N_3329,N_2327,N_393);
or U3330 (N_3330,N_781,N_1519);
nand U3331 (N_3331,N_52,N_1018);
nor U3332 (N_3332,N_1044,N_2435);
nor U3333 (N_3333,N_2273,N_2328);
or U3334 (N_3334,N_601,N_2238);
nand U3335 (N_3335,N_1175,N_62);
or U3336 (N_3336,N_675,N_1911);
nor U3337 (N_3337,N_1185,N_1251);
and U3338 (N_3338,N_1210,N_2075);
nand U3339 (N_3339,N_1851,N_107);
nor U3340 (N_3340,N_2278,N_1556);
nor U3341 (N_3341,N_1067,N_366);
nand U3342 (N_3342,N_874,N_1064);
and U3343 (N_3343,N_1098,N_806);
nor U3344 (N_3344,N_527,N_1453);
or U3345 (N_3345,N_496,N_1743);
nand U3346 (N_3346,N_1842,N_577);
and U3347 (N_3347,N_2033,N_1645);
nor U3348 (N_3348,N_1377,N_163);
nand U3349 (N_3349,N_866,N_783);
nand U3350 (N_3350,N_901,N_2137);
and U3351 (N_3351,N_1469,N_136);
nor U3352 (N_3352,N_701,N_2074);
nor U3353 (N_3353,N_1202,N_1483);
nand U3354 (N_3354,N_2479,N_1539);
and U3355 (N_3355,N_310,N_1391);
nor U3356 (N_3356,N_1389,N_292);
and U3357 (N_3357,N_469,N_2394);
nand U3358 (N_3358,N_1810,N_2239);
xnor U3359 (N_3359,N_439,N_1452);
nor U3360 (N_3360,N_1606,N_913);
and U3361 (N_3361,N_549,N_890);
or U3362 (N_3362,N_713,N_1910);
nor U3363 (N_3363,N_333,N_2236);
or U3364 (N_3364,N_1171,N_2260);
and U3365 (N_3365,N_153,N_385);
nor U3366 (N_3366,N_2418,N_194);
nand U3367 (N_3367,N_1920,N_1699);
nor U3368 (N_3368,N_2494,N_2175);
or U3369 (N_3369,N_1950,N_1028);
nor U3370 (N_3370,N_586,N_90);
nand U3371 (N_3371,N_2011,N_286);
and U3372 (N_3372,N_1804,N_1571);
nand U3373 (N_3373,N_1205,N_2073);
nand U3374 (N_3374,N_299,N_722);
nor U3375 (N_3375,N_113,N_1423);
nor U3376 (N_3376,N_1035,N_1170);
xnor U3377 (N_3377,N_631,N_1355);
and U3378 (N_3378,N_1521,N_1584);
nand U3379 (N_3379,N_2326,N_25);
nor U3380 (N_3380,N_1632,N_102);
and U3381 (N_3381,N_2112,N_685);
or U3382 (N_3382,N_658,N_428);
or U3383 (N_3383,N_152,N_1013);
or U3384 (N_3384,N_2089,N_1111);
or U3385 (N_3385,N_2174,N_1634);
or U3386 (N_3386,N_1287,N_2341);
nor U3387 (N_3387,N_547,N_2265);
or U3388 (N_3388,N_1065,N_287);
xor U3389 (N_3389,N_865,N_1476);
nand U3390 (N_3390,N_654,N_2022);
and U3391 (N_3391,N_826,N_1954);
and U3392 (N_3392,N_630,N_1332);
and U3393 (N_3393,N_290,N_66);
and U3394 (N_3394,N_1765,N_12);
nand U3395 (N_3395,N_449,N_373);
nand U3396 (N_3396,N_2347,N_1191);
and U3397 (N_3397,N_1410,N_2076);
nand U3398 (N_3398,N_1690,N_1092);
nand U3399 (N_3399,N_733,N_5);
and U3400 (N_3400,N_705,N_1325);
and U3401 (N_3401,N_845,N_1335);
and U3402 (N_3402,N_1953,N_38);
or U3403 (N_3403,N_859,N_1369);
and U3404 (N_3404,N_732,N_1146);
nand U3405 (N_3405,N_2324,N_236);
nand U3406 (N_3406,N_118,N_2222);
nand U3407 (N_3407,N_2368,N_1520);
or U3408 (N_3408,N_1007,N_2212);
or U3409 (N_3409,N_2421,N_628);
or U3410 (N_3410,N_2122,N_467);
or U3411 (N_3411,N_804,N_948);
nand U3412 (N_3412,N_1893,N_2436);
nand U3413 (N_3413,N_937,N_1643);
nor U3414 (N_3414,N_116,N_743);
or U3415 (N_3415,N_1153,N_178);
nor U3416 (N_3416,N_1194,N_2119);
nor U3417 (N_3417,N_1676,N_765);
and U3418 (N_3418,N_1054,N_1319);
or U3419 (N_3419,N_580,N_2470);
and U3420 (N_3420,N_23,N_1166);
nor U3421 (N_3421,N_2448,N_1428);
and U3422 (N_3422,N_784,N_1880);
nand U3423 (N_3423,N_672,N_702);
nand U3424 (N_3424,N_1635,N_1125);
or U3425 (N_3425,N_1923,N_1344);
and U3426 (N_3426,N_1148,N_2192);
or U3427 (N_3427,N_571,N_141);
nand U3428 (N_3428,N_1293,N_997);
nor U3429 (N_3429,N_255,N_1603);
nor U3430 (N_3430,N_818,N_1014);
or U3431 (N_3431,N_172,N_1421);
nand U3432 (N_3432,N_2423,N_207);
nand U3433 (N_3433,N_2207,N_1379);
nor U3434 (N_3434,N_2351,N_505);
nand U3435 (N_3435,N_203,N_1051);
nor U3436 (N_3436,N_2279,N_1390);
nor U3437 (N_3437,N_1354,N_1123);
or U3438 (N_3438,N_2131,N_860);
nand U3439 (N_3439,N_2032,N_156);
nor U3440 (N_3440,N_1628,N_1246);
or U3441 (N_3441,N_1560,N_1303);
nor U3442 (N_3442,N_455,N_1652);
and U3443 (N_3443,N_169,N_2093);
or U3444 (N_3444,N_595,N_76);
and U3445 (N_3445,N_1241,N_2334);
and U3446 (N_3446,N_1058,N_873);
nand U3447 (N_3447,N_1322,N_801);
nand U3448 (N_3448,N_828,N_1413);
nand U3449 (N_3449,N_534,N_2453);
nor U3450 (N_3450,N_328,N_1591);
and U3451 (N_3451,N_480,N_2234);
nand U3452 (N_3452,N_1466,N_1818);
nand U3453 (N_3453,N_2454,N_2261);
nor U3454 (N_3454,N_108,N_2080);
or U3455 (N_3455,N_735,N_1885);
and U3456 (N_3456,N_1729,N_1057);
or U3457 (N_3457,N_2484,N_869);
nand U3458 (N_3458,N_291,N_542);
nand U3459 (N_3459,N_949,N_533);
nand U3460 (N_3460,N_1802,N_1816);
nor U3461 (N_3461,N_1850,N_1670);
nand U3462 (N_3462,N_746,N_967);
nand U3463 (N_3463,N_1255,N_1422);
nand U3464 (N_3464,N_650,N_1499);
nand U3465 (N_3465,N_210,N_665);
nor U3466 (N_3466,N_1438,N_812);
or U3467 (N_3467,N_271,N_1892);
nor U3468 (N_3468,N_1192,N_933);
and U3469 (N_3469,N_1773,N_1841);
nor U3470 (N_3470,N_1141,N_2420);
and U3471 (N_3471,N_1090,N_2400);
nor U3472 (N_3472,N_111,N_2017);
nor U3473 (N_3473,N_1333,N_410);
or U3474 (N_3474,N_2185,N_238);
nor U3475 (N_3475,N_1068,N_2116);
nor U3476 (N_3476,N_355,N_1439);
nand U3477 (N_3477,N_73,N_2297);
nor U3478 (N_3478,N_2458,N_1627);
and U3479 (N_3479,N_540,N_201);
nor U3480 (N_3480,N_2405,N_293);
nand U3481 (N_3481,N_2431,N_897);
and U3482 (N_3482,N_1724,N_581);
or U3483 (N_3483,N_119,N_2390);
or U3484 (N_3484,N_1894,N_2003);
and U3485 (N_3485,N_965,N_1157);
and U3486 (N_3486,N_2321,N_462);
nand U3487 (N_3487,N_1181,N_1588);
or U3488 (N_3488,N_773,N_994);
nor U3489 (N_3489,N_454,N_1557);
nor U3490 (N_3490,N_834,N_597);
nor U3491 (N_3491,N_1343,N_726);
nand U3492 (N_3492,N_221,N_877);
or U3493 (N_3493,N_2107,N_1496);
nand U3494 (N_3494,N_1549,N_1347);
nand U3495 (N_3495,N_2224,N_727);
or U3496 (N_3496,N_2370,N_1698);
and U3497 (N_3497,N_625,N_1296);
nor U3498 (N_3498,N_370,N_1412);
and U3499 (N_3499,N_2441,N_1297);
and U3500 (N_3500,N_1155,N_605);
and U3501 (N_3501,N_791,N_1115);
or U3502 (N_3502,N_1919,N_1059);
nor U3503 (N_3503,N_1026,N_986);
and U3504 (N_3504,N_2094,N_599);
and U3505 (N_3505,N_2317,N_1583);
or U3506 (N_3506,N_164,N_764);
nand U3507 (N_3507,N_1165,N_2210);
nand U3508 (N_3508,N_1005,N_1600);
nor U3509 (N_3509,N_1062,N_546);
and U3510 (N_3510,N_399,N_387);
nor U3511 (N_3511,N_20,N_1829);
and U3512 (N_3512,N_2130,N_2443);
or U3513 (N_3513,N_1867,N_779);
or U3514 (N_3514,N_962,N_1883);
nor U3515 (N_3515,N_1397,N_1264);
nor U3516 (N_3516,N_1038,N_444);
nor U3517 (N_3517,N_6,N_797);
and U3518 (N_3518,N_214,N_553);
and U3519 (N_3519,N_1409,N_1200);
or U3520 (N_3520,N_1715,N_1227);
nand U3521 (N_3521,N_787,N_170);
or U3522 (N_3522,N_639,N_2120);
or U3523 (N_3523,N_1587,N_1042);
nand U3524 (N_3524,N_2025,N_418);
or U3525 (N_3525,N_215,N_15);
and U3526 (N_3526,N_2323,N_2415);
or U3527 (N_3527,N_698,N_566);
nand U3528 (N_3528,N_2048,N_1714);
nand U3529 (N_3529,N_1315,N_1767);
or U3530 (N_3530,N_782,N_2489);
nor U3531 (N_3531,N_969,N_2339);
and U3532 (N_3532,N_1029,N_922);
or U3533 (N_3533,N_105,N_2030);
or U3534 (N_3534,N_1150,N_2071);
and U3535 (N_3535,N_1095,N_275);
or U3536 (N_3536,N_2438,N_2495);
or U3537 (N_3537,N_2203,N_810);
or U3538 (N_3538,N_212,N_1233);
or U3539 (N_3539,N_250,N_602);
nand U3540 (N_3540,N_1394,N_1184);
nor U3541 (N_3541,N_1276,N_2439);
nand U3542 (N_3542,N_794,N_667);
or U3543 (N_3543,N_1243,N_219);
or U3544 (N_3544,N_2386,N_1037);
and U3545 (N_3545,N_317,N_1305);
or U3546 (N_3546,N_2322,N_485);
nor U3547 (N_3547,N_2123,N_2422);
nand U3548 (N_3548,N_2250,N_876);
nor U3549 (N_3549,N_1854,N_686);
nor U3550 (N_3550,N_706,N_1278);
and U3551 (N_3551,N_1669,N_1944);
or U3552 (N_3552,N_1712,N_1616);
and U3553 (N_3553,N_1882,N_1400);
nor U3554 (N_3554,N_1812,N_1350);
or U3555 (N_3555,N_895,N_2332);
nand U3556 (N_3556,N_1103,N_1126);
and U3557 (N_3557,N_1683,N_725);
and U3558 (N_3558,N_766,N_1824);
or U3559 (N_3559,N_856,N_495);
nor U3560 (N_3560,N_2360,N_44);
or U3561 (N_3561,N_321,N_1225);
nand U3562 (N_3562,N_545,N_2209);
and U3563 (N_3563,N_1167,N_452);
nor U3564 (N_3564,N_304,N_2081);
nor U3565 (N_3565,N_166,N_1238);
nor U3566 (N_3566,N_1489,N_1559);
nand U3567 (N_3567,N_909,N_335);
nor U3568 (N_3568,N_1999,N_923);
nand U3569 (N_3569,N_1536,N_2426);
xnor U3570 (N_3570,N_637,N_296);
nor U3571 (N_3571,N_1563,N_1768);
and U3572 (N_3572,N_2243,N_1613);
nand U3573 (N_3573,N_1646,N_2490);
nand U3574 (N_3574,N_973,N_1465);
and U3575 (N_3575,N_332,N_1301);
nand U3576 (N_3576,N_307,N_1418);
and U3577 (N_3577,N_1876,N_1845);
or U3578 (N_3578,N_2053,N_1472);
nand U3579 (N_3579,N_2437,N_532);
or U3580 (N_3580,N_1751,N_2050);
nor U3581 (N_3581,N_1352,N_376);
and U3582 (N_3582,N_1085,N_1746);
or U3583 (N_3583,N_1000,N_622);
or U3584 (N_3584,N_2153,N_1527);
and U3585 (N_3585,N_2110,N_763);
and U3586 (N_3586,N_996,N_920);
nor U3587 (N_3587,N_839,N_1199);
nand U3588 (N_3588,N_1505,N_1728);
nand U3589 (N_3589,N_541,N_1361);
nor U3590 (N_3590,N_589,N_793);
nor U3591 (N_3591,N_985,N_2216);
nor U3592 (N_3592,N_1621,N_318);
and U3593 (N_3593,N_720,N_204);
and U3594 (N_3594,N_1958,N_552);
nor U3595 (N_3595,N_609,N_2374);
nor U3596 (N_3596,N_1494,N_1602);
and U3597 (N_3597,N_1398,N_123);
nand U3598 (N_3598,N_17,N_145);
nand U3599 (N_3599,N_1437,N_1782);
or U3600 (N_3600,N_1215,N_1137);
or U3601 (N_3601,N_195,N_1935);
or U3602 (N_3602,N_1003,N_1201);
and U3603 (N_3603,N_1385,N_1615);
or U3604 (N_3604,N_426,N_1660);
nand U3605 (N_3605,N_4,N_329);
nor U3606 (N_3606,N_1537,N_2264);
and U3607 (N_3607,N_608,N_1962);
and U3608 (N_3608,N_1993,N_516);
nor U3609 (N_3609,N_1041,N_2162);
nor U3610 (N_3610,N_1977,N_319);
nand U3611 (N_3611,N_1012,N_2428);
nand U3612 (N_3612,N_938,N_253);
or U3613 (N_3613,N_814,N_847);
nand U3614 (N_3614,N_2241,N_1517);
and U3615 (N_3615,N_1809,N_703);
nor U3616 (N_3616,N_1980,N_591);
nand U3617 (N_3617,N_1975,N_1234);
nand U3618 (N_3618,N_2491,N_2452);
or U3619 (N_3619,N_817,N_488);
and U3620 (N_3620,N_2061,N_1434);
nor U3621 (N_3621,N_2395,N_2335);
and U3622 (N_3622,N_2270,N_1351);
nor U3623 (N_3623,N_7,N_721);
nor U3624 (N_3624,N_1899,N_1884);
nand U3625 (N_3625,N_1716,N_1786);
or U3626 (N_3626,N_617,N_1832);
nand U3627 (N_3627,N_1384,N_227);
nand U3628 (N_3628,N_2135,N_1076);
and U3629 (N_3629,N_1546,N_147);
nor U3630 (N_3630,N_652,N_1640);
nor U3631 (N_3631,N_1755,N_242);
and U3632 (N_3632,N_2160,N_2088);
and U3633 (N_3633,N_651,N_1682);
nand U3634 (N_3634,N_1161,N_1564);
nor U3635 (N_3635,N_2357,N_2117);
or U3636 (N_3636,N_925,N_1637);
and U3637 (N_3637,N_1594,N_2218);
nor U3638 (N_3638,N_1861,N_1798);
or U3639 (N_3639,N_1813,N_267);
nand U3640 (N_3640,N_2451,N_1609);
nand U3641 (N_3641,N_1959,N_1156);
and U3642 (N_3642,N_2393,N_1796);
nand U3643 (N_3643,N_1807,N_284);
or U3644 (N_3644,N_524,N_1063);
nor U3645 (N_3645,N_1504,N_115);
or U3646 (N_3646,N_27,N_403);
and U3647 (N_3647,N_2244,N_2106);
or U3648 (N_3648,N_63,N_2013);
nor U3649 (N_3649,N_1055,N_1965);
nand U3650 (N_3650,N_334,N_1477);
or U3651 (N_3651,N_1552,N_186);
xor U3652 (N_3652,N_165,N_1823);
nor U3653 (N_3653,N_2101,N_2365);
or U3654 (N_3654,N_198,N_2097);
nor U3655 (N_3655,N_492,N_2496);
and U3656 (N_3656,N_244,N_2183);
nor U3657 (N_3657,N_2389,N_2180);
or U3658 (N_3658,N_700,N_498);
or U3659 (N_3659,N_629,N_298);
or U3660 (N_3660,N_1501,N_1770);
nand U3661 (N_3661,N_1725,N_550);
nor U3662 (N_3662,N_1346,N_1956);
nor U3663 (N_3663,N_437,N_256);
nand U3664 (N_3664,N_2353,N_167);
or U3665 (N_3665,N_862,N_34);
nor U3666 (N_3666,N_2154,N_951);
nor U3667 (N_3667,N_2127,N_2336);
nand U3668 (N_3668,N_303,N_1034);
nor U3669 (N_3669,N_971,N_83);
and U3670 (N_3670,N_596,N_2021);
nor U3671 (N_3671,N_1857,N_1983);
nand U3672 (N_3672,N_1118,N_1053);
nor U3673 (N_3673,N_150,N_1328);
nor U3674 (N_3674,N_579,N_1182);
and U3675 (N_3675,N_1703,N_1506);
nand U3676 (N_3676,N_2060,N_750);
or U3677 (N_3677,N_2249,N_1930);
nor U3678 (N_3678,N_1990,N_2136);
and U3679 (N_3679,N_1195,N_2493);
nor U3680 (N_3680,N_677,N_285);
and U3681 (N_3681,N_1794,N_1795);
nand U3682 (N_3682,N_880,N_770);
nor U3683 (N_3683,N_1750,N_196);
nand U3684 (N_3684,N_173,N_657);
and U3685 (N_3685,N_1245,N_903);
or U3686 (N_3686,N_1183,N_1648);
or U3687 (N_3687,N_2240,N_2068);
and U3688 (N_3688,N_2000,N_1134);
or U3689 (N_3689,N_289,N_1102);
or U3690 (N_3690,N_1154,N_1747);
nand U3691 (N_3691,N_822,N_870);
or U3692 (N_3692,N_536,N_1862);
nand U3693 (N_3693,N_84,N_747);
nor U3694 (N_3694,N_181,N_313);
nor U3695 (N_3695,N_2189,N_278);
nor U3696 (N_3696,N_661,N_670);
nor U3697 (N_3697,N_934,N_1719);
or U3698 (N_3698,N_800,N_636);
nor U3699 (N_3699,N_1969,N_2171);
or U3700 (N_3700,N_1945,N_1839);
nor U3701 (N_3701,N_2023,N_1788);
or U3702 (N_3702,N_1787,N_276);
or U3703 (N_3703,N_956,N_2215);
or U3704 (N_3704,N_2257,N_1163);
and U3705 (N_3705,N_78,N_2086);
or U3706 (N_3706,N_272,N_1599);
or U3707 (N_3707,N_222,N_2380);
nand U3708 (N_3708,N_1294,N_679);
or U3709 (N_3709,N_1833,N_1760);
and U3710 (N_3710,N_1047,N_1083);
and U3711 (N_3711,N_1490,N_87);
nand U3712 (N_3712,N_1262,N_2411);
and U3713 (N_3713,N_995,N_582);
and U3714 (N_3714,N_400,N_1019);
or U3715 (N_3715,N_414,N_619);
or U3716 (N_3716,N_1097,N_409);
or U3717 (N_3717,N_2256,N_1285);
or U3718 (N_3718,N_106,N_362);
or U3719 (N_3719,N_1772,N_1040);
and U3720 (N_3720,N_805,N_346);
nor U3721 (N_3721,N_425,N_2383);
and U3722 (N_3722,N_1497,N_70);
nor U3723 (N_3723,N_1512,N_2253);
nand U3724 (N_3724,N_555,N_104);
and U3725 (N_3725,N_415,N_522);
nor U3726 (N_3726,N_56,N_2082);
nor U3727 (N_3727,N_624,N_2387);
nor U3728 (N_3728,N_2104,N_830);
nor U3729 (N_3729,N_881,N_1487);
or U3730 (N_3730,N_1091,N_1906);
nand U3731 (N_3731,N_1997,N_1524);
nor U3732 (N_3732,N_336,N_1924);
nand U3733 (N_3733,N_2469,N_92);
and U3734 (N_3734,N_1654,N_2417);
and U3735 (N_3735,N_1025,N_347);
nand U3736 (N_3736,N_2146,N_990);
and U3737 (N_3737,N_1272,N_2472);
and U3738 (N_3738,N_374,N_2488);
xnor U3739 (N_3739,N_268,N_1046);
nand U3740 (N_3740,N_1644,N_2201);
nor U3741 (N_3741,N_2002,N_1204);
nor U3742 (N_3742,N_2055,N_1540);
nand U3743 (N_3743,N_1279,N_1678);
or U3744 (N_3744,N_1250,N_2325);
nand U3745 (N_3745,N_1467,N_513);
or U3746 (N_3746,N_2442,N_607);
nand U3747 (N_3747,N_2027,N_1668);
or U3748 (N_3748,N_1364,N_708);
and U3749 (N_3749,N_1607,N_1792);
nor U3750 (N_3750,N_513,N_736);
and U3751 (N_3751,N_1359,N_1950);
and U3752 (N_3752,N_861,N_1063);
and U3753 (N_3753,N_1386,N_1074);
nor U3754 (N_3754,N_1984,N_2386);
and U3755 (N_3755,N_1545,N_2458);
and U3756 (N_3756,N_390,N_1388);
or U3757 (N_3757,N_229,N_1111);
nor U3758 (N_3758,N_1198,N_1820);
nand U3759 (N_3759,N_109,N_730);
nor U3760 (N_3760,N_1632,N_200);
or U3761 (N_3761,N_1357,N_576);
and U3762 (N_3762,N_362,N_1669);
nor U3763 (N_3763,N_335,N_626);
nor U3764 (N_3764,N_291,N_1360);
or U3765 (N_3765,N_976,N_2346);
or U3766 (N_3766,N_1999,N_1002);
or U3767 (N_3767,N_568,N_1890);
xor U3768 (N_3768,N_183,N_1749);
xnor U3769 (N_3769,N_1707,N_2029);
xor U3770 (N_3770,N_1596,N_331);
or U3771 (N_3771,N_2088,N_191);
nand U3772 (N_3772,N_1615,N_2284);
or U3773 (N_3773,N_1051,N_991);
nand U3774 (N_3774,N_11,N_300);
nor U3775 (N_3775,N_2416,N_1198);
nand U3776 (N_3776,N_1617,N_1409);
nor U3777 (N_3777,N_1246,N_2298);
and U3778 (N_3778,N_2061,N_1887);
or U3779 (N_3779,N_1741,N_1578);
or U3780 (N_3780,N_1209,N_488);
or U3781 (N_3781,N_1598,N_756);
nor U3782 (N_3782,N_131,N_1099);
nand U3783 (N_3783,N_1036,N_2238);
or U3784 (N_3784,N_2434,N_1061);
and U3785 (N_3785,N_1449,N_836);
nand U3786 (N_3786,N_1176,N_1617);
and U3787 (N_3787,N_2213,N_541);
and U3788 (N_3788,N_75,N_715);
and U3789 (N_3789,N_1369,N_212);
nor U3790 (N_3790,N_70,N_889);
nand U3791 (N_3791,N_710,N_265);
nand U3792 (N_3792,N_1848,N_1573);
and U3793 (N_3793,N_1058,N_1253);
and U3794 (N_3794,N_217,N_2355);
nor U3795 (N_3795,N_690,N_2147);
nor U3796 (N_3796,N_1463,N_2090);
nand U3797 (N_3797,N_934,N_2047);
nor U3798 (N_3798,N_308,N_2169);
nor U3799 (N_3799,N_2279,N_283);
nand U3800 (N_3800,N_1387,N_872);
and U3801 (N_3801,N_2299,N_2153);
or U3802 (N_3802,N_1605,N_2123);
nor U3803 (N_3803,N_35,N_605);
nor U3804 (N_3804,N_129,N_2075);
and U3805 (N_3805,N_1460,N_1850);
or U3806 (N_3806,N_1761,N_642);
or U3807 (N_3807,N_2250,N_2103);
and U3808 (N_3808,N_364,N_2092);
nor U3809 (N_3809,N_1106,N_674);
and U3810 (N_3810,N_2204,N_1006);
or U3811 (N_3811,N_1314,N_216);
or U3812 (N_3812,N_1033,N_345);
or U3813 (N_3813,N_892,N_28);
nand U3814 (N_3814,N_877,N_2474);
nor U3815 (N_3815,N_553,N_1277);
or U3816 (N_3816,N_831,N_20);
and U3817 (N_3817,N_2009,N_2303);
or U3818 (N_3818,N_1254,N_2499);
and U3819 (N_3819,N_853,N_935);
nand U3820 (N_3820,N_91,N_1551);
nand U3821 (N_3821,N_271,N_1752);
or U3822 (N_3822,N_723,N_1060);
nand U3823 (N_3823,N_2473,N_2495);
nor U3824 (N_3824,N_1298,N_1947);
or U3825 (N_3825,N_2222,N_1536);
nor U3826 (N_3826,N_463,N_1930);
and U3827 (N_3827,N_595,N_763);
and U3828 (N_3828,N_571,N_2276);
or U3829 (N_3829,N_2298,N_2207);
or U3830 (N_3830,N_306,N_11);
nand U3831 (N_3831,N_1797,N_419);
nor U3832 (N_3832,N_50,N_1412);
nand U3833 (N_3833,N_562,N_806);
nor U3834 (N_3834,N_1285,N_690);
and U3835 (N_3835,N_721,N_719);
or U3836 (N_3836,N_2169,N_16);
nor U3837 (N_3837,N_1492,N_635);
or U3838 (N_3838,N_1762,N_989);
and U3839 (N_3839,N_869,N_1363);
and U3840 (N_3840,N_2434,N_356);
nand U3841 (N_3841,N_1145,N_2042);
or U3842 (N_3842,N_1678,N_1395);
nand U3843 (N_3843,N_1545,N_962);
nand U3844 (N_3844,N_1426,N_2017);
and U3845 (N_3845,N_1577,N_1284);
and U3846 (N_3846,N_718,N_1679);
nand U3847 (N_3847,N_547,N_125);
or U3848 (N_3848,N_522,N_798);
and U3849 (N_3849,N_785,N_1606);
or U3850 (N_3850,N_655,N_1509);
or U3851 (N_3851,N_2408,N_681);
nand U3852 (N_3852,N_2028,N_390);
or U3853 (N_3853,N_2176,N_457);
or U3854 (N_3854,N_2082,N_75);
and U3855 (N_3855,N_403,N_1398);
nor U3856 (N_3856,N_291,N_1829);
or U3857 (N_3857,N_117,N_1880);
and U3858 (N_3858,N_2302,N_399);
and U3859 (N_3859,N_199,N_1631);
and U3860 (N_3860,N_1945,N_140);
nor U3861 (N_3861,N_1273,N_735);
and U3862 (N_3862,N_1049,N_704);
or U3863 (N_3863,N_1473,N_1658);
nor U3864 (N_3864,N_362,N_943);
nor U3865 (N_3865,N_1885,N_416);
nand U3866 (N_3866,N_1486,N_756);
and U3867 (N_3867,N_274,N_1842);
nand U3868 (N_3868,N_1181,N_1524);
or U3869 (N_3869,N_1634,N_2178);
nor U3870 (N_3870,N_1767,N_1881);
or U3871 (N_3871,N_1883,N_1488);
nor U3872 (N_3872,N_1905,N_2485);
nand U3873 (N_3873,N_2448,N_1758);
or U3874 (N_3874,N_1678,N_1550);
nand U3875 (N_3875,N_2433,N_469);
nand U3876 (N_3876,N_362,N_301);
nor U3877 (N_3877,N_538,N_2208);
or U3878 (N_3878,N_1364,N_86);
nor U3879 (N_3879,N_1006,N_1635);
or U3880 (N_3880,N_1590,N_513);
or U3881 (N_3881,N_1096,N_1802);
and U3882 (N_3882,N_2445,N_1615);
nor U3883 (N_3883,N_508,N_1343);
and U3884 (N_3884,N_1021,N_1653);
nor U3885 (N_3885,N_725,N_355);
or U3886 (N_3886,N_2413,N_2060);
or U3887 (N_3887,N_198,N_2124);
nand U3888 (N_3888,N_990,N_2318);
nor U3889 (N_3889,N_965,N_1112);
or U3890 (N_3890,N_1194,N_351);
nand U3891 (N_3891,N_160,N_563);
nor U3892 (N_3892,N_1348,N_1631);
nor U3893 (N_3893,N_1802,N_1903);
nand U3894 (N_3894,N_675,N_37);
or U3895 (N_3895,N_1705,N_1008);
and U3896 (N_3896,N_447,N_753);
and U3897 (N_3897,N_1249,N_794);
and U3898 (N_3898,N_1852,N_2174);
nor U3899 (N_3899,N_109,N_225);
or U3900 (N_3900,N_1793,N_142);
nor U3901 (N_3901,N_928,N_2287);
or U3902 (N_3902,N_983,N_591);
or U3903 (N_3903,N_657,N_698);
nand U3904 (N_3904,N_798,N_2105);
and U3905 (N_3905,N_537,N_448);
nor U3906 (N_3906,N_322,N_2154);
nand U3907 (N_3907,N_71,N_939);
nor U3908 (N_3908,N_694,N_608);
nand U3909 (N_3909,N_208,N_1111);
nand U3910 (N_3910,N_656,N_1751);
and U3911 (N_3911,N_1729,N_1229);
nand U3912 (N_3912,N_1822,N_626);
or U3913 (N_3913,N_1456,N_1993);
nand U3914 (N_3914,N_214,N_903);
nand U3915 (N_3915,N_2445,N_390);
or U3916 (N_3916,N_1814,N_1497);
or U3917 (N_3917,N_868,N_95);
nand U3918 (N_3918,N_1134,N_1398);
nor U3919 (N_3919,N_2170,N_2007);
and U3920 (N_3920,N_1364,N_1297);
nor U3921 (N_3921,N_1613,N_2068);
and U3922 (N_3922,N_818,N_239);
and U3923 (N_3923,N_512,N_584);
nor U3924 (N_3924,N_586,N_112);
nor U3925 (N_3925,N_2122,N_491);
nor U3926 (N_3926,N_604,N_2041);
nor U3927 (N_3927,N_1802,N_2236);
nand U3928 (N_3928,N_1596,N_1217);
and U3929 (N_3929,N_469,N_596);
nand U3930 (N_3930,N_1306,N_2007);
or U3931 (N_3931,N_2276,N_881);
and U3932 (N_3932,N_2220,N_1991);
nand U3933 (N_3933,N_564,N_1044);
nor U3934 (N_3934,N_2417,N_1838);
nor U3935 (N_3935,N_2383,N_300);
nor U3936 (N_3936,N_740,N_273);
nand U3937 (N_3937,N_968,N_1720);
and U3938 (N_3938,N_1049,N_51);
and U3939 (N_3939,N_1892,N_744);
nand U3940 (N_3940,N_27,N_648);
nor U3941 (N_3941,N_856,N_1333);
nor U3942 (N_3942,N_2239,N_1824);
and U3943 (N_3943,N_1591,N_2123);
nand U3944 (N_3944,N_2084,N_39);
or U3945 (N_3945,N_1782,N_142);
and U3946 (N_3946,N_2436,N_1327);
nor U3947 (N_3947,N_1032,N_396);
or U3948 (N_3948,N_882,N_1247);
nand U3949 (N_3949,N_384,N_87);
and U3950 (N_3950,N_2442,N_1812);
nor U3951 (N_3951,N_1664,N_2016);
nand U3952 (N_3952,N_1427,N_1250);
nand U3953 (N_3953,N_2460,N_1465);
nand U3954 (N_3954,N_63,N_338);
nor U3955 (N_3955,N_1919,N_96);
and U3956 (N_3956,N_274,N_517);
nor U3957 (N_3957,N_1993,N_1803);
and U3958 (N_3958,N_2405,N_1475);
or U3959 (N_3959,N_2202,N_2334);
or U3960 (N_3960,N_2460,N_1116);
nor U3961 (N_3961,N_744,N_144);
nand U3962 (N_3962,N_1558,N_428);
or U3963 (N_3963,N_1435,N_2149);
or U3964 (N_3964,N_378,N_1065);
or U3965 (N_3965,N_2051,N_1816);
or U3966 (N_3966,N_609,N_225);
nor U3967 (N_3967,N_1605,N_2288);
xor U3968 (N_3968,N_2009,N_1375);
nor U3969 (N_3969,N_967,N_309);
nand U3970 (N_3970,N_1094,N_2053);
or U3971 (N_3971,N_2475,N_1790);
or U3972 (N_3972,N_510,N_1192);
nor U3973 (N_3973,N_1965,N_136);
or U3974 (N_3974,N_2316,N_2011);
or U3975 (N_3975,N_985,N_269);
and U3976 (N_3976,N_873,N_2070);
nor U3977 (N_3977,N_1189,N_1025);
or U3978 (N_3978,N_577,N_1862);
nor U3979 (N_3979,N_968,N_2021);
nor U3980 (N_3980,N_1261,N_2482);
and U3981 (N_3981,N_179,N_2477);
nand U3982 (N_3982,N_2166,N_1636);
and U3983 (N_3983,N_1484,N_15);
nand U3984 (N_3984,N_567,N_390);
nand U3985 (N_3985,N_2352,N_2336);
nor U3986 (N_3986,N_2170,N_1473);
nor U3987 (N_3987,N_1988,N_369);
nand U3988 (N_3988,N_2022,N_844);
nor U3989 (N_3989,N_2435,N_2091);
and U3990 (N_3990,N_1305,N_325);
and U3991 (N_3991,N_2394,N_1500);
nor U3992 (N_3992,N_372,N_1466);
nand U3993 (N_3993,N_1869,N_71);
nor U3994 (N_3994,N_1393,N_1192);
nor U3995 (N_3995,N_554,N_180);
nand U3996 (N_3996,N_2459,N_174);
nor U3997 (N_3997,N_730,N_1432);
and U3998 (N_3998,N_765,N_2198);
nor U3999 (N_3999,N_2423,N_782);
nor U4000 (N_4000,N_1365,N_2030);
and U4001 (N_4001,N_1275,N_1164);
nor U4002 (N_4002,N_2040,N_2447);
and U4003 (N_4003,N_1226,N_628);
nand U4004 (N_4004,N_1051,N_2486);
or U4005 (N_4005,N_28,N_1438);
or U4006 (N_4006,N_1587,N_779);
nand U4007 (N_4007,N_1021,N_1706);
or U4008 (N_4008,N_1812,N_2434);
and U4009 (N_4009,N_1796,N_1496);
nand U4010 (N_4010,N_418,N_2307);
or U4011 (N_4011,N_382,N_693);
nor U4012 (N_4012,N_2126,N_1553);
nand U4013 (N_4013,N_1095,N_674);
and U4014 (N_4014,N_2087,N_280);
or U4015 (N_4015,N_1601,N_624);
or U4016 (N_4016,N_57,N_288);
or U4017 (N_4017,N_969,N_2073);
nand U4018 (N_4018,N_817,N_992);
and U4019 (N_4019,N_310,N_1484);
and U4020 (N_4020,N_1478,N_1573);
and U4021 (N_4021,N_1509,N_1167);
or U4022 (N_4022,N_2376,N_732);
nor U4023 (N_4023,N_684,N_1918);
nand U4024 (N_4024,N_474,N_1675);
nor U4025 (N_4025,N_1852,N_1419);
nand U4026 (N_4026,N_1969,N_2390);
nor U4027 (N_4027,N_461,N_2459);
nand U4028 (N_4028,N_1528,N_761);
or U4029 (N_4029,N_1644,N_2393);
and U4030 (N_4030,N_2335,N_1260);
nor U4031 (N_4031,N_1237,N_523);
nor U4032 (N_4032,N_1141,N_1435);
and U4033 (N_4033,N_1300,N_1033);
or U4034 (N_4034,N_1229,N_1709);
nor U4035 (N_4035,N_1249,N_982);
nand U4036 (N_4036,N_507,N_115);
nand U4037 (N_4037,N_1867,N_1294);
or U4038 (N_4038,N_2352,N_1043);
or U4039 (N_4039,N_2351,N_1661);
nand U4040 (N_4040,N_261,N_399);
nor U4041 (N_4041,N_1478,N_1880);
nor U4042 (N_4042,N_1249,N_1850);
nand U4043 (N_4043,N_1805,N_169);
and U4044 (N_4044,N_1196,N_354);
or U4045 (N_4045,N_753,N_395);
nor U4046 (N_4046,N_127,N_2463);
or U4047 (N_4047,N_1546,N_1317);
and U4048 (N_4048,N_1831,N_2041);
nor U4049 (N_4049,N_2482,N_1993);
nor U4050 (N_4050,N_1186,N_1756);
or U4051 (N_4051,N_470,N_1029);
nor U4052 (N_4052,N_2269,N_2435);
nand U4053 (N_4053,N_1042,N_2018);
nor U4054 (N_4054,N_1121,N_2107);
and U4055 (N_4055,N_717,N_1865);
or U4056 (N_4056,N_587,N_2273);
and U4057 (N_4057,N_311,N_867);
and U4058 (N_4058,N_1870,N_893);
or U4059 (N_4059,N_101,N_2430);
nand U4060 (N_4060,N_173,N_2011);
and U4061 (N_4061,N_301,N_1631);
and U4062 (N_4062,N_637,N_1713);
and U4063 (N_4063,N_1424,N_993);
nor U4064 (N_4064,N_94,N_1945);
nor U4065 (N_4065,N_132,N_2285);
and U4066 (N_4066,N_1724,N_1338);
or U4067 (N_4067,N_980,N_2470);
nand U4068 (N_4068,N_2065,N_2001);
nor U4069 (N_4069,N_574,N_695);
and U4070 (N_4070,N_2079,N_2375);
nand U4071 (N_4071,N_491,N_1094);
and U4072 (N_4072,N_576,N_613);
nand U4073 (N_4073,N_819,N_736);
nand U4074 (N_4074,N_2086,N_2308);
and U4075 (N_4075,N_760,N_1419);
nand U4076 (N_4076,N_1641,N_952);
and U4077 (N_4077,N_945,N_2408);
and U4078 (N_4078,N_632,N_1999);
nor U4079 (N_4079,N_150,N_2153);
or U4080 (N_4080,N_1431,N_1119);
or U4081 (N_4081,N_924,N_61);
and U4082 (N_4082,N_1771,N_888);
nor U4083 (N_4083,N_2032,N_1315);
nor U4084 (N_4084,N_1030,N_1118);
nand U4085 (N_4085,N_2052,N_466);
nand U4086 (N_4086,N_1531,N_2416);
nor U4087 (N_4087,N_2268,N_39);
nand U4088 (N_4088,N_1721,N_1981);
nand U4089 (N_4089,N_404,N_1684);
and U4090 (N_4090,N_946,N_129);
or U4091 (N_4091,N_1053,N_36);
nand U4092 (N_4092,N_285,N_89);
and U4093 (N_4093,N_1851,N_1732);
or U4094 (N_4094,N_1238,N_1299);
and U4095 (N_4095,N_77,N_185);
nand U4096 (N_4096,N_1170,N_293);
and U4097 (N_4097,N_100,N_2084);
or U4098 (N_4098,N_937,N_163);
and U4099 (N_4099,N_1476,N_2289);
and U4100 (N_4100,N_1001,N_2064);
nor U4101 (N_4101,N_553,N_962);
nand U4102 (N_4102,N_349,N_277);
nor U4103 (N_4103,N_2128,N_727);
or U4104 (N_4104,N_1848,N_765);
or U4105 (N_4105,N_1530,N_1146);
nand U4106 (N_4106,N_380,N_1326);
nor U4107 (N_4107,N_1531,N_70);
or U4108 (N_4108,N_1289,N_2438);
or U4109 (N_4109,N_753,N_556);
or U4110 (N_4110,N_483,N_408);
nor U4111 (N_4111,N_992,N_1399);
nor U4112 (N_4112,N_474,N_1808);
nand U4113 (N_4113,N_726,N_1638);
and U4114 (N_4114,N_1393,N_1218);
and U4115 (N_4115,N_2459,N_1232);
or U4116 (N_4116,N_939,N_1858);
and U4117 (N_4117,N_1009,N_2071);
nor U4118 (N_4118,N_132,N_739);
nor U4119 (N_4119,N_1953,N_293);
nand U4120 (N_4120,N_1088,N_2218);
nor U4121 (N_4121,N_1668,N_1567);
or U4122 (N_4122,N_2153,N_973);
or U4123 (N_4123,N_32,N_2212);
and U4124 (N_4124,N_1652,N_196);
and U4125 (N_4125,N_1440,N_2236);
or U4126 (N_4126,N_2185,N_2346);
nand U4127 (N_4127,N_2258,N_2112);
nor U4128 (N_4128,N_85,N_2430);
nor U4129 (N_4129,N_456,N_2238);
or U4130 (N_4130,N_1598,N_202);
or U4131 (N_4131,N_38,N_821);
and U4132 (N_4132,N_1279,N_1316);
nand U4133 (N_4133,N_1610,N_1344);
and U4134 (N_4134,N_1163,N_1324);
and U4135 (N_4135,N_982,N_329);
or U4136 (N_4136,N_104,N_290);
or U4137 (N_4137,N_1075,N_2024);
and U4138 (N_4138,N_2390,N_771);
xnor U4139 (N_4139,N_1216,N_2157);
and U4140 (N_4140,N_740,N_1441);
or U4141 (N_4141,N_1926,N_804);
nor U4142 (N_4142,N_2428,N_1753);
and U4143 (N_4143,N_317,N_1548);
and U4144 (N_4144,N_35,N_989);
and U4145 (N_4145,N_189,N_412);
nand U4146 (N_4146,N_1991,N_914);
nand U4147 (N_4147,N_1518,N_30);
nor U4148 (N_4148,N_1047,N_1971);
nand U4149 (N_4149,N_2491,N_433);
or U4150 (N_4150,N_1873,N_534);
nand U4151 (N_4151,N_2012,N_1613);
or U4152 (N_4152,N_837,N_2331);
and U4153 (N_4153,N_1726,N_1634);
nor U4154 (N_4154,N_1991,N_2094);
or U4155 (N_4155,N_1,N_152);
xor U4156 (N_4156,N_408,N_1545);
nor U4157 (N_4157,N_2230,N_830);
nor U4158 (N_4158,N_645,N_440);
and U4159 (N_4159,N_582,N_1560);
nor U4160 (N_4160,N_980,N_212);
or U4161 (N_4161,N_2111,N_48);
nor U4162 (N_4162,N_1862,N_80);
and U4163 (N_4163,N_1436,N_2010);
or U4164 (N_4164,N_2055,N_1917);
and U4165 (N_4165,N_1478,N_739);
or U4166 (N_4166,N_1340,N_1488);
and U4167 (N_4167,N_2208,N_649);
and U4168 (N_4168,N_912,N_2081);
nand U4169 (N_4169,N_868,N_2460);
nand U4170 (N_4170,N_1351,N_1048);
nand U4171 (N_4171,N_1805,N_1433);
nor U4172 (N_4172,N_446,N_1078);
or U4173 (N_4173,N_1471,N_594);
nor U4174 (N_4174,N_1842,N_1431);
nand U4175 (N_4175,N_2061,N_2443);
and U4176 (N_4176,N_1637,N_776);
or U4177 (N_4177,N_1384,N_1411);
and U4178 (N_4178,N_153,N_28);
nand U4179 (N_4179,N_1223,N_275);
nand U4180 (N_4180,N_557,N_122);
nor U4181 (N_4181,N_1503,N_2487);
nand U4182 (N_4182,N_2032,N_1685);
nand U4183 (N_4183,N_195,N_618);
or U4184 (N_4184,N_1393,N_2134);
and U4185 (N_4185,N_164,N_1252);
or U4186 (N_4186,N_412,N_75);
and U4187 (N_4187,N_2262,N_1484);
nand U4188 (N_4188,N_2430,N_1449);
or U4189 (N_4189,N_1516,N_326);
nand U4190 (N_4190,N_1381,N_2030);
nor U4191 (N_4191,N_528,N_819);
nor U4192 (N_4192,N_1233,N_1348);
or U4193 (N_4193,N_1731,N_1711);
or U4194 (N_4194,N_1818,N_1442);
and U4195 (N_4195,N_54,N_1460);
or U4196 (N_4196,N_869,N_751);
and U4197 (N_4197,N_2197,N_1832);
or U4198 (N_4198,N_70,N_473);
nand U4199 (N_4199,N_927,N_674);
nor U4200 (N_4200,N_404,N_1781);
and U4201 (N_4201,N_757,N_1599);
nor U4202 (N_4202,N_1487,N_1462);
nand U4203 (N_4203,N_2083,N_958);
nand U4204 (N_4204,N_1934,N_542);
nor U4205 (N_4205,N_1948,N_1151);
nor U4206 (N_4206,N_1072,N_619);
xnor U4207 (N_4207,N_1492,N_1333);
or U4208 (N_4208,N_1473,N_1455);
nor U4209 (N_4209,N_350,N_654);
nand U4210 (N_4210,N_2078,N_761);
nand U4211 (N_4211,N_1545,N_2348);
nand U4212 (N_4212,N_131,N_767);
or U4213 (N_4213,N_2248,N_564);
nor U4214 (N_4214,N_670,N_748);
nand U4215 (N_4215,N_1894,N_2260);
nor U4216 (N_4216,N_2362,N_1183);
nor U4217 (N_4217,N_835,N_1338);
and U4218 (N_4218,N_993,N_1962);
nor U4219 (N_4219,N_762,N_1682);
nor U4220 (N_4220,N_2278,N_1441);
nor U4221 (N_4221,N_1403,N_1330);
nand U4222 (N_4222,N_1994,N_1745);
or U4223 (N_4223,N_1129,N_2416);
or U4224 (N_4224,N_1780,N_875);
and U4225 (N_4225,N_1509,N_226);
or U4226 (N_4226,N_2428,N_136);
nand U4227 (N_4227,N_2201,N_1080);
nor U4228 (N_4228,N_2262,N_1721);
and U4229 (N_4229,N_1207,N_217);
or U4230 (N_4230,N_898,N_975);
and U4231 (N_4231,N_1337,N_2195);
nor U4232 (N_4232,N_1648,N_1496);
nand U4233 (N_4233,N_821,N_731);
or U4234 (N_4234,N_923,N_1659);
xor U4235 (N_4235,N_2346,N_354);
or U4236 (N_4236,N_99,N_1919);
or U4237 (N_4237,N_693,N_903);
and U4238 (N_4238,N_990,N_2472);
and U4239 (N_4239,N_1516,N_2416);
nor U4240 (N_4240,N_696,N_944);
nor U4241 (N_4241,N_995,N_2106);
and U4242 (N_4242,N_577,N_1012);
nand U4243 (N_4243,N_993,N_55);
or U4244 (N_4244,N_640,N_1355);
nand U4245 (N_4245,N_1690,N_1820);
and U4246 (N_4246,N_2276,N_228);
nor U4247 (N_4247,N_2208,N_2118);
nand U4248 (N_4248,N_1889,N_1026);
or U4249 (N_4249,N_478,N_94);
nor U4250 (N_4250,N_93,N_383);
nor U4251 (N_4251,N_1345,N_1341);
nor U4252 (N_4252,N_631,N_889);
or U4253 (N_4253,N_1978,N_194);
or U4254 (N_4254,N_2080,N_1230);
or U4255 (N_4255,N_687,N_97);
nand U4256 (N_4256,N_2438,N_2166);
nand U4257 (N_4257,N_1131,N_638);
nor U4258 (N_4258,N_201,N_1975);
nor U4259 (N_4259,N_359,N_2169);
and U4260 (N_4260,N_510,N_2245);
nand U4261 (N_4261,N_1303,N_2221);
nand U4262 (N_4262,N_2347,N_758);
or U4263 (N_4263,N_960,N_2411);
nor U4264 (N_4264,N_1905,N_1607);
nand U4265 (N_4265,N_1094,N_801);
and U4266 (N_4266,N_161,N_2179);
nor U4267 (N_4267,N_903,N_1665);
and U4268 (N_4268,N_212,N_221);
or U4269 (N_4269,N_989,N_1198);
nand U4270 (N_4270,N_2086,N_731);
nor U4271 (N_4271,N_839,N_1523);
or U4272 (N_4272,N_2309,N_1310);
or U4273 (N_4273,N_2226,N_1840);
or U4274 (N_4274,N_191,N_2012);
nor U4275 (N_4275,N_1843,N_2433);
and U4276 (N_4276,N_2125,N_243);
nor U4277 (N_4277,N_1051,N_421);
or U4278 (N_4278,N_848,N_1229);
nand U4279 (N_4279,N_2206,N_684);
nand U4280 (N_4280,N_2079,N_384);
or U4281 (N_4281,N_273,N_739);
nand U4282 (N_4282,N_408,N_2496);
and U4283 (N_4283,N_144,N_1675);
and U4284 (N_4284,N_393,N_1233);
or U4285 (N_4285,N_1383,N_2064);
and U4286 (N_4286,N_1665,N_1410);
nand U4287 (N_4287,N_2053,N_272);
or U4288 (N_4288,N_252,N_597);
or U4289 (N_4289,N_186,N_2372);
nand U4290 (N_4290,N_1858,N_2067);
or U4291 (N_4291,N_790,N_2469);
nand U4292 (N_4292,N_110,N_1260);
nand U4293 (N_4293,N_2058,N_32);
or U4294 (N_4294,N_2063,N_367);
or U4295 (N_4295,N_2065,N_1462);
nand U4296 (N_4296,N_1285,N_876);
nand U4297 (N_4297,N_1432,N_2295);
and U4298 (N_4298,N_920,N_704);
nand U4299 (N_4299,N_616,N_754);
nand U4300 (N_4300,N_2372,N_1293);
nand U4301 (N_4301,N_1847,N_639);
xnor U4302 (N_4302,N_1117,N_457);
and U4303 (N_4303,N_255,N_2418);
and U4304 (N_4304,N_2367,N_1647);
nand U4305 (N_4305,N_2407,N_502);
nor U4306 (N_4306,N_434,N_2246);
and U4307 (N_4307,N_204,N_2449);
nor U4308 (N_4308,N_1871,N_2245);
nor U4309 (N_4309,N_873,N_2448);
nor U4310 (N_4310,N_1002,N_1743);
nor U4311 (N_4311,N_1760,N_743);
nor U4312 (N_4312,N_1692,N_679);
or U4313 (N_4313,N_1649,N_989);
and U4314 (N_4314,N_2334,N_311);
or U4315 (N_4315,N_2326,N_313);
nor U4316 (N_4316,N_1675,N_826);
nand U4317 (N_4317,N_2184,N_450);
or U4318 (N_4318,N_1452,N_1643);
nand U4319 (N_4319,N_827,N_95);
and U4320 (N_4320,N_256,N_563);
nor U4321 (N_4321,N_979,N_1063);
nor U4322 (N_4322,N_582,N_2235);
nor U4323 (N_4323,N_1996,N_1376);
nor U4324 (N_4324,N_1563,N_944);
nor U4325 (N_4325,N_163,N_159);
nand U4326 (N_4326,N_179,N_425);
and U4327 (N_4327,N_796,N_2101);
nand U4328 (N_4328,N_902,N_559);
or U4329 (N_4329,N_1249,N_1646);
nand U4330 (N_4330,N_992,N_181);
nand U4331 (N_4331,N_2052,N_1849);
or U4332 (N_4332,N_1451,N_2003);
and U4333 (N_4333,N_577,N_2279);
nor U4334 (N_4334,N_689,N_433);
and U4335 (N_4335,N_1875,N_132);
nor U4336 (N_4336,N_2409,N_1729);
nor U4337 (N_4337,N_33,N_1689);
nor U4338 (N_4338,N_1855,N_2390);
nor U4339 (N_4339,N_1626,N_494);
and U4340 (N_4340,N_1975,N_7);
nor U4341 (N_4341,N_1135,N_1021);
nand U4342 (N_4342,N_1830,N_2165);
nand U4343 (N_4343,N_301,N_1644);
and U4344 (N_4344,N_1245,N_2023);
and U4345 (N_4345,N_940,N_1923);
or U4346 (N_4346,N_485,N_2095);
or U4347 (N_4347,N_1744,N_1256);
nor U4348 (N_4348,N_627,N_382);
and U4349 (N_4349,N_2090,N_576);
and U4350 (N_4350,N_503,N_535);
or U4351 (N_4351,N_2321,N_45);
and U4352 (N_4352,N_145,N_35);
nor U4353 (N_4353,N_1386,N_1716);
and U4354 (N_4354,N_1573,N_366);
and U4355 (N_4355,N_182,N_995);
xor U4356 (N_4356,N_381,N_1189);
and U4357 (N_4357,N_2053,N_1604);
or U4358 (N_4358,N_649,N_361);
or U4359 (N_4359,N_1801,N_583);
or U4360 (N_4360,N_1952,N_920);
and U4361 (N_4361,N_1183,N_2234);
or U4362 (N_4362,N_1200,N_632);
or U4363 (N_4363,N_1808,N_1278);
and U4364 (N_4364,N_1879,N_1580);
or U4365 (N_4365,N_1833,N_158);
nand U4366 (N_4366,N_1739,N_2249);
or U4367 (N_4367,N_1620,N_396);
nand U4368 (N_4368,N_162,N_988);
and U4369 (N_4369,N_1043,N_1563);
and U4370 (N_4370,N_1238,N_549);
or U4371 (N_4371,N_798,N_345);
and U4372 (N_4372,N_958,N_1356);
nor U4373 (N_4373,N_1124,N_229);
and U4374 (N_4374,N_1996,N_326);
and U4375 (N_4375,N_67,N_543);
nor U4376 (N_4376,N_972,N_2355);
nand U4377 (N_4377,N_1983,N_709);
nand U4378 (N_4378,N_100,N_3);
nor U4379 (N_4379,N_2172,N_1243);
nand U4380 (N_4380,N_1927,N_33);
nor U4381 (N_4381,N_2020,N_395);
and U4382 (N_4382,N_1546,N_933);
or U4383 (N_4383,N_1466,N_1130);
nand U4384 (N_4384,N_1490,N_1478);
nor U4385 (N_4385,N_1046,N_1433);
nor U4386 (N_4386,N_698,N_1208);
or U4387 (N_4387,N_299,N_2493);
and U4388 (N_4388,N_2318,N_2000);
nor U4389 (N_4389,N_2271,N_229);
nor U4390 (N_4390,N_229,N_77);
and U4391 (N_4391,N_1227,N_1150);
nor U4392 (N_4392,N_1410,N_588);
nand U4393 (N_4393,N_533,N_277);
xnor U4394 (N_4394,N_173,N_18);
or U4395 (N_4395,N_2165,N_1584);
or U4396 (N_4396,N_2151,N_66);
nand U4397 (N_4397,N_656,N_448);
nor U4398 (N_4398,N_2084,N_2174);
or U4399 (N_4399,N_1296,N_373);
or U4400 (N_4400,N_307,N_40);
or U4401 (N_4401,N_1878,N_1912);
nand U4402 (N_4402,N_1235,N_514);
nor U4403 (N_4403,N_777,N_763);
and U4404 (N_4404,N_78,N_432);
nor U4405 (N_4405,N_282,N_60);
xor U4406 (N_4406,N_1033,N_2312);
and U4407 (N_4407,N_1193,N_117);
or U4408 (N_4408,N_109,N_2278);
and U4409 (N_4409,N_946,N_1379);
or U4410 (N_4410,N_915,N_2413);
and U4411 (N_4411,N_1049,N_2252);
nand U4412 (N_4412,N_1425,N_984);
or U4413 (N_4413,N_2286,N_2213);
nand U4414 (N_4414,N_962,N_55);
or U4415 (N_4415,N_600,N_2322);
or U4416 (N_4416,N_5,N_1850);
nand U4417 (N_4417,N_985,N_1940);
nor U4418 (N_4418,N_2474,N_1832);
nor U4419 (N_4419,N_1827,N_888);
nand U4420 (N_4420,N_1033,N_2285);
and U4421 (N_4421,N_1395,N_1292);
nor U4422 (N_4422,N_1182,N_843);
and U4423 (N_4423,N_1357,N_1121);
nor U4424 (N_4424,N_1450,N_960);
nand U4425 (N_4425,N_1606,N_404);
nand U4426 (N_4426,N_1384,N_2245);
nor U4427 (N_4427,N_289,N_1274);
nor U4428 (N_4428,N_2389,N_61);
or U4429 (N_4429,N_541,N_879);
and U4430 (N_4430,N_857,N_1703);
and U4431 (N_4431,N_2129,N_1598);
nand U4432 (N_4432,N_797,N_1554);
or U4433 (N_4433,N_1050,N_1795);
nor U4434 (N_4434,N_1305,N_785);
nand U4435 (N_4435,N_395,N_2482);
nand U4436 (N_4436,N_2210,N_480);
and U4437 (N_4437,N_1194,N_1122);
nand U4438 (N_4438,N_2259,N_886);
nor U4439 (N_4439,N_2420,N_1874);
or U4440 (N_4440,N_2188,N_1481);
nand U4441 (N_4441,N_142,N_1784);
nand U4442 (N_4442,N_1788,N_842);
or U4443 (N_4443,N_533,N_468);
nor U4444 (N_4444,N_1746,N_2357);
and U4445 (N_4445,N_490,N_971);
nand U4446 (N_4446,N_2059,N_145);
nand U4447 (N_4447,N_529,N_249);
and U4448 (N_4448,N_2143,N_1226);
and U4449 (N_4449,N_1507,N_1725);
and U4450 (N_4450,N_981,N_1290);
nand U4451 (N_4451,N_2400,N_317);
nor U4452 (N_4452,N_2238,N_814);
nand U4453 (N_4453,N_1551,N_1576);
or U4454 (N_4454,N_1071,N_257);
and U4455 (N_4455,N_1709,N_1909);
nand U4456 (N_4456,N_173,N_2499);
nor U4457 (N_4457,N_2393,N_877);
nor U4458 (N_4458,N_2487,N_1237);
nand U4459 (N_4459,N_487,N_2467);
nor U4460 (N_4460,N_60,N_1243);
or U4461 (N_4461,N_2414,N_678);
nor U4462 (N_4462,N_37,N_1546);
or U4463 (N_4463,N_1767,N_1775);
nor U4464 (N_4464,N_548,N_149);
nor U4465 (N_4465,N_111,N_1458);
nor U4466 (N_4466,N_1985,N_245);
nor U4467 (N_4467,N_1061,N_2151);
or U4468 (N_4468,N_2359,N_1423);
nand U4469 (N_4469,N_2234,N_88);
and U4470 (N_4470,N_2263,N_1777);
or U4471 (N_4471,N_1380,N_44);
nor U4472 (N_4472,N_2374,N_1100);
or U4473 (N_4473,N_2435,N_102);
nor U4474 (N_4474,N_2261,N_1809);
or U4475 (N_4475,N_1458,N_878);
and U4476 (N_4476,N_224,N_1441);
nor U4477 (N_4477,N_101,N_181);
nand U4478 (N_4478,N_1064,N_1223);
nand U4479 (N_4479,N_728,N_1266);
nor U4480 (N_4480,N_974,N_93);
nand U4481 (N_4481,N_172,N_1775);
or U4482 (N_4482,N_1683,N_818);
or U4483 (N_4483,N_1842,N_1524);
xnor U4484 (N_4484,N_1202,N_690);
and U4485 (N_4485,N_1692,N_1402);
and U4486 (N_4486,N_1074,N_790);
or U4487 (N_4487,N_2114,N_1332);
and U4488 (N_4488,N_1309,N_1866);
nand U4489 (N_4489,N_1622,N_56);
nand U4490 (N_4490,N_73,N_2204);
nand U4491 (N_4491,N_1783,N_1917);
nor U4492 (N_4492,N_2040,N_1508);
or U4493 (N_4493,N_228,N_1038);
nand U4494 (N_4494,N_1026,N_911);
nand U4495 (N_4495,N_1565,N_807);
and U4496 (N_4496,N_856,N_20);
and U4497 (N_4497,N_715,N_2381);
nor U4498 (N_4498,N_1546,N_2246);
and U4499 (N_4499,N_859,N_709);
xnor U4500 (N_4500,N_173,N_258);
nand U4501 (N_4501,N_2044,N_281);
and U4502 (N_4502,N_2186,N_355);
and U4503 (N_4503,N_368,N_1313);
nor U4504 (N_4504,N_1384,N_2092);
nand U4505 (N_4505,N_1111,N_1438);
or U4506 (N_4506,N_1099,N_1162);
or U4507 (N_4507,N_875,N_1403);
and U4508 (N_4508,N_289,N_254);
nor U4509 (N_4509,N_1469,N_1579);
or U4510 (N_4510,N_2010,N_1755);
nand U4511 (N_4511,N_1099,N_1648);
and U4512 (N_4512,N_109,N_158);
or U4513 (N_4513,N_2187,N_942);
nor U4514 (N_4514,N_2337,N_486);
nand U4515 (N_4515,N_649,N_1571);
and U4516 (N_4516,N_1292,N_1279);
nand U4517 (N_4517,N_1588,N_1446);
nand U4518 (N_4518,N_832,N_478);
nand U4519 (N_4519,N_1954,N_931);
or U4520 (N_4520,N_1180,N_211);
or U4521 (N_4521,N_802,N_1908);
nor U4522 (N_4522,N_1761,N_851);
or U4523 (N_4523,N_397,N_1719);
and U4524 (N_4524,N_174,N_2473);
xor U4525 (N_4525,N_1526,N_1024);
nor U4526 (N_4526,N_1675,N_1920);
and U4527 (N_4527,N_2369,N_1083);
and U4528 (N_4528,N_929,N_1870);
nor U4529 (N_4529,N_1191,N_1037);
nand U4530 (N_4530,N_1932,N_2477);
nor U4531 (N_4531,N_1411,N_286);
and U4532 (N_4532,N_1260,N_322);
nand U4533 (N_4533,N_539,N_1001);
nor U4534 (N_4534,N_2223,N_1880);
nor U4535 (N_4535,N_877,N_1583);
nor U4536 (N_4536,N_2232,N_788);
or U4537 (N_4537,N_1726,N_2028);
nor U4538 (N_4538,N_2036,N_446);
nor U4539 (N_4539,N_1926,N_1744);
nor U4540 (N_4540,N_389,N_1558);
or U4541 (N_4541,N_566,N_1255);
nor U4542 (N_4542,N_796,N_1604);
nand U4543 (N_4543,N_1850,N_103);
xnor U4544 (N_4544,N_1674,N_168);
nand U4545 (N_4545,N_1368,N_340);
and U4546 (N_4546,N_886,N_2287);
nor U4547 (N_4547,N_2112,N_189);
nand U4548 (N_4548,N_2075,N_1750);
nor U4549 (N_4549,N_2151,N_1806);
or U4550 (N_4550,N_1017,N_65);
or U4551 (N_4551,N_1100,N_1720);
and U4552 (N_4552,N_981,N_1827);
or U4553 (N_4553,N_1216,N_1964);
xnor U4554 (N_4554,N_1751,N_1522);
or U4555 (N_4555,N_551,N_2101);
nand U4556 (N_4556,N_1882,N_156);
nand U4557 (N_4557,N_947,N_226);
and U4558 (N_4558,N_1172,N_987);
and U4559 (N_4559,N_581,N_1038);
or U4560 (N_4560,N_821,N_1830);
and U4561 (N_4561,N_1897,N_1867);
nand U4562 (N_4562,N_1218,N_1500);
nor U4563 (N_4563,N_190,N_1020);
nand U4564 (N_4564,N_2212,N_990);
and U4565 (N_4565,N_839,N_263);
and U4566 (N_4566,N_1340,N_489);
nor U4567 (N_4567,N_644,N_960);
and U4568 (N_4568,N_1453,N_1682);
nor U4569 (N_4569,N_1271,N_633);
and U4570 (N_4570,N_2391,N_2007);
nor U4571 (N_4571,N_1160,N_2174);
and U4572 (N_4572,N_1030,N_269);
xor U4573 (N_4573,N_1312,N_471);
nand U4574 (N_4574,N_2250,N_668);
nor U4575 (N_4575,N_104,N_40);
nand U4576 (N_4576,N_1510,N_1137);
and U4577 (N_4577,N_157,N_305);
or U4578 (N_4578,N_381,N_423);
nor U4579 (N_4579,N_1894,N_1794);
or U4580 (N_4580,N_375,N_2438);
nand U4581 (N_4581,N_221,N_1016);
nand U4582 (N_4582,N_1820,N_924);
nand U4583 (N_4583,N_1402,N_626);
nor U4584 (N_4584,N_2336,N_1367);
and U4585 (N_4585,N_1716,N_164);
and U4586 (N_4586,N_750,N_1904);
and U4587 (N_4587,N_2033,N_844);
and U4588 (N_4588,N_285,N_1642);
nand U4589 (N_4589,N_275,N_2384);
nand U4590 (N_4590,N_1140,N_681);
or U4591 (N_4591,N_2088,N_263);
and U4592 (N_4592,N_792,N_780);
nand U4593 (N_4593,N_176,N_950);
nand U4594 (N_4594,N_2064,N_1883);
or U4595 (N_4595,N_1412,N_1090);
or U4596 (N_4596,N_2472,N_1140);
nand U4597 (N_4597,N_1160,N_1242);
nor U4598 (N_4598,N_2388,N_1657);
and U4599 (N_4599,N_385,N_176);
and U4600 (N_4600,N_1743,N_2284);
or U4601 (N_4601,N_1112,N_1788);
and U4602 (N_4602,N_1585,N_753);
nor U4603 (N_4603,N_2012,N_911);
and U4604 (N_4604,N_1107,N_2277);
nand U4605 (N_4605,N_711,N_1867);
nand U4606 (N_4606,N_918,N_446);
and U4607 (N_4607,N_2131,N_1144);
or U4608 (N_4608,N_1477,N_1604);
nand U4609 (N_4609,N_2484,N_108);
nor U4610 (N_4610,N_615,N_2400);
or U4611 (N_4611,N_1293,N_2460);
nand U4612 (N_4612,N_2300,N_2283);
nand U4613 (N_4613,N_32,N_852);
nor U4614 (N_4614,N_2146,N_16);
nand U4615 (N_4615,N_2061,N_136);
and U4616 (N_4616,N_852,N_1694);
and U4617 (N_4617,N_770,N_1573);
and U4618 (N_4618,N_164,N_708);
nand U4619 (N_4619,N_80,N_2048);
nor U4620 (N_4620,N_2029,N_1072);
or U4621 (N_4621,N_2337,N_1060);
or U4622 (N_4622,N_275,N_777);
and U4623 (N_4623,N_1518,N_1305);
and U4624 (N_4624,N_2495,N_944);
or U4625 (N_4625,N_1015,N_430);
and U4626 (N_4626,N_1282,N_2061);
and U4627 (N_4627,N_1708,N_1300);
nand U4628 (N_4628,N_212,N_2432);
and U4629 (N_4629,N_1492,N_1052);
or U4630 (N_4630,N_1988,N_497);
nor U4631 (N_4631,N_1447,N_1338);
and U4632 (N_4632,N_1311,N_1872);
and U4633 (N_4633,N_1900,N_1302);
nor U4634 (N_4634,N_419,N_781);
and U4635 (N_4635,N_668,N_2334);
nor U4636 (N_4636,N_741,N_2256);
nand U4637 (N_4637,N_2158,N_976);
or U4638 (N_4638,N_1944,N_177);
nor U4639 (N_4639,N_1524,N_2276);
nand U4640 (N_4640,N_1363,N_959);
and U4641 (N_4641,N_2083,N_1101);
or U4642 (N_4642,N_465,N_1859);
and U4643 (N_4643,N_323,N_2351);
and U4644 (N_4644,N_426,N_2355);
and U4645 (N_4645,N_1420,N_1113);
nor U4646 (N_4646,N_1045,N_2475);
nand U4647 (N_4647,N_2480,N_1269);
nand U4648 (N_4648,N_273,N_817);
nand U4649 (N_4649,N_2052,N_1225);
nor U4650 (N_4650,N_1514,N_288);
xnor U4651 (N_4651,N_1617,N_2493);
or U4652 (N_4652,N_1470,N_897);
nand U4653 (N_4653,N_997,N_2373);
nor U4654 (N_4654,N_93,N_2161);
nor U4655 (N_4655,N_2329,N_1611);
or U4656 (N_4656,N_2453,N_1043);
and U4657 (N_4657,N_1076,N_572);
nand U4658 (N_4658,N_2155,N_2301);
nor U4659 (N_4659,N_829,N_1158);
and U4660 (N_4660,N_1923,N_2412);
nand U4661 (N_4661,N_249,N_1768);
or U4662 (N_4662,N_1080,N_300);
nor U4663 (N_4663,N_1401,N_2008);
or U4664 (N_4664,N_48,N_1971);
or U4665 (N_4665,N_305,N_973);
nand U4666 (N_4666,N_754,N_1587);
nor U4667 (N_4667,N_920,N_627);
and U4668 (N_4668,N_1446,N_915);
or U4669 (N_4669,N_2021,N_1329);
and U4670 (N_4670,N_1296,N_1009);
nand U4671 (N_4671,N_465,N_2381);
nor U4672 (N_4672,N_333,N_786);
nor U4673 (N_4673,N_2299,N_744);
nor U4674 (N_4674,N_1552,N_2037);
nand U4675 (N_4675,N_781,N_13);
or U4676 (N_4676,N_811,N_1353);
and U4677 (N_4677,N_1828,N_2351);
or U4678 (N_4678,N_2048,N_1824);
or U4679 (N_4679,N_2448,N_1663);
nand U4680 (N_4680,N_1373,N_1396);
and U4681 (N_4681,N_2199,N_832);
nor U4682 (N_4682,N_1328,N_57);
nand U4683 (N_4683,N_1423,N_2193);
or U4684 (N_4684,N_0,N_2340);
or U4685 (N_4685,N_1672,N_1740);
nand U4686 (N_4686,N_1860,N_1931);
and U4687 (N_4687,N_982,N_2079);
and U4688 (N_4688,N_1562,N_2469);
nor U4689 (N_4689,N_1713,N_1694);
or U4690 (N_4690,N_929,N_1825);
or U4691 (N_4691,N_79,N_1289);
or U4692 (N_4692,N_694,N_2319);
nand U4693 (N_4693,N_481,N_594);
and U4694 (N_4694,N_181,N_2036);
and U4695 (N_4695,N_1196,N_1191);
and U4696 (N_4696,N_1669,N_1800);
nor U4697 (N_4697,N_1573,N_583);
and U4698 (N_4698,N_990,N_2468);
nand U4699 (N_4699,N_2180,N_1188);
nor U4700 (N_4700,N_2255,N_1694);
and U4701 (N_4701,N_860,N_1953);
nand U4702 (N_4702,N_592,N_551);
nand U4703 (N_4703,N_2172,N_2252);
and U4704 (N_4704,N_1809,N_2335);
nand U4705 (N_4705,N_2034,N_1266);
and U4706 (N_4706,N_2488,N_595);
nor U4707 (N_4707,N_1936,N_1285);
and U4708 (N_4708,N_165,N_898);
nor U4709 (N_4709,N_2256,N_2226);
or U4710 (N_4710,N_2113,N_931);
or U4711 (N_4711,N_760,N_1268);
nor U4712 (N_4712,N_2422,N_2160);
or U4713 (N_4713,N_2192,N_93);
and U4714 (N_4714,N_2404,N_187);
nor U4715 (N_4715,N_1462,N_704);
or U4716 (N_4716,N_1896,N_1255);
and U4717 (N_4717,N_767,N_645);
nor U4718 (N_4718,N_743,N_1668);
nand U4719 (N_4719,N_2113,N_37);
nor U4720 (N_4720,N_1788,N_586);
nand U4721 (N_4721,N_329,N_722);
or U4722 (N_4722,N_2425,N_65);
nand U4723 (N_4723,N_463,N_574);
or U4724 (N_4724,N_2061,N_71);
and U4725 (N_4725,N_2290,N_1506);
nor U4726 (N_4726,N_250,N_128);
and U4727 (N_4727,N_2408,N_592);
or U4728 (N_4728,N_808,N_2150);
or U4729 (N_4729,N_6,N_1819);
and U4730 (N_4730,N_834,N_2091);
and U4731 (N_4731,N_2111,N_563);
and U4732 (N_4732,N_1448,N_440);
or U4733 (N_4733,N_233,N_2122);
nand U4734 (N_4734,N_262,N_2316);
nor U4735 (N_4735,N_2422,N_56);
or U4736 (N_4736,N_14,N_2302);
or U4737 (N_4737,N_1290,N_966);
and U4738 (N_4738,N_1632,N_982);
nor U4739 (N_4739,N_1790,N_787);
and U4740 (N_4740,N_2225,N_2323);
nor U4741 (N_4741,N_431,N_132);
and U4742 (N_4742,N_1294,N_83);
nand U4743 (N_4743,N_2326,N_2126);
or U4744 (N_4744,N_1923,N_1879);
nor U4745 (N_4745,N_1222,N_1503);
nor U4746 (N_4746,N_1591,N_1584);
nand U4747 (N_4747,N_1376,N_1198);
nand U4748 (N_4748,N_381,N_351);
nor U4749 (N_4749,N_2439,N_2124);
or U4750 (N_4750,N_1202,N_949);
nand U4751 (N_4751,N_2171,N_1830);
nor U4752 (N_4752,N_1898,N_1840);
and U4753 (N_4753,N_449,N_319);
and U4754 (N_4754,N_2177,N_1212);
nand U4755 (N_4755,N_585,N_2061);
and U4756 (N_4756,N_1642,N_2444);
and U4757 (N_4757,N_1678,N_2148);
nor U4758 (N_4758,N_139,N_2380);
or U4759 (N_4759,N_1213,N_2210);
nor U4760 (N_4760,N_663,N_202);
or U4761 (N_4761,N_445,N_1799);
nand U4762 (N_4762,N_769,N_2200);
and U4763 (N_4763,N_1745,N_661);
nor U4764 (N_4764,N_278,N_2323);
nor U4765 (N_4765,N_1783,N_757);
nor U4766 (N_4766,N_1805,N_2381);
and U4767 (N_4767,N_501,N_2183);
nor U4768 (N_4768,N_1836,N_2217);
nand U4769 (N_4769,N_2096,N_1626);
nor U4770 (N_4770,N_759,N_244);
nor U4771 (N_4771,N_25,N_1062);
or U4772 (N_4772,N_1997,N_302);
and U4773 (N_4773,N_2100,N_1454);
or U4774 (N_4774,N_1027,N_579);
nand U4775 (N_4775,N_1260,N_2019);
or U4776 (N_4776,N_2170,N_290);
and U4777 (N_4777,N_2360,N_1017);
and U4778 (N_4778,N_1762,N_1298);
and U4779 (N_4779,N_1694,N_1153);
nand U4780 (N_4780,N_356,N_13);
and U4781 (N_4781,N_1151,N_1940);
and U4782 (N_4782,N_2256,N_2480);
and U4783 (N_4783,N_2181,N_1279);
nand U4784 (N_4784,N_2400,N_1549);
nand U4785 (N_4785,N_182,N_1306);
and U4786 (N_4786,N_331,N_2477);
and U4787 (N_4787,N_1682,N_1241);
nor U4788 (N_4788,N_2380,N_906);
nor U4789 (N_4789,N_1390,N_1355);
nor U4790 (N_4790,N_2172,N_1312);
nor U4791 (N_4791,N_1904,N_1786);
nand U4792 (N_4792,N_1724,N_111);
and U4793 (N_4793,N_2365,N_1234);
nand U4794 (N_4794,N_1317,N_438);
or U4795 (N_4795,N_761,N_463);
nor U4796 (N_4796,N_1034,N_2390);
nor U4797 (N_4797,N_2297,N_2304);
nor U4798 (N_4798,N_1407,N_1772);
nand U4799 (N_4799,N_354,N_356);
and U4800 (N_4800,N_320,N_1080);
and U4801 (N_4801,N_2258,N_448);
or U4802 (N_4802,N_31,N_1597);
nor U4803 (N_4803,N_1493,N_1965);
and U4804 (N_4804,N_304,N_1771);
and U4805 (N_4805,N_1455,N_240);
nand U4806 (N_4806,N_843,N_1620);
nor U4807 (N_4807,N_1284,N_2325);
nor U4808 (N_4808,N_1739,N_329);
or U4809 (N_4809,N_238,N_1144);
and U4810 (N_4810,N_207,N_1828);
or U4811 (N_4811,N_2064,N_1675);
and U4812 (N_4812,N_505,N_314);
or U4813 (N_4813,N_514,N_2019);
and U4814 (N_4814,N_308,N_2276);
nand U4815 (N_4815,N_753,N_287);
nand U4816 (N_4816,N_2270,N_1276);
nor U4817 (N_4817,N_868,N_2010);
nand U4818 (N_4818,N_194,N_521);
xor U4819 (N_4819,N_216,N_1583);
nor U4820 (N_4820,N_1499,N_202);
nand U4821 (N_4821,N_400,N_1030);
nor U4822 (N_4822,N_113,N_99);
nor U4823 (N_4823,N_411,N_447);
or U4824 (N_4824,N_989,N_1872);
nor U4825 (N_4825,N_682,N_1840);
nor U4826 (N_4826,N_68,N_2289);
nor U4827 (N_4827,N_1460,N_1194);
nand U4828 (N_4828,N_1651,N_1487);
nand U4829 (N_4829,N_2125,N_78);
nor U4830 (N_4830,N_1837,N_895);
nand U4831 (N_4831,N_2155,N_1819);
and U4832 (N_4832,N_1421,N_197);
and U4833 (N_4833,N_848,N_2264);
or U4834 (N_4834,N_820,N_1769);
nor U4835 (N_4835,N_1093,N_1370);
nor U4836 (N_4836,N_418,N_741);
nor U4837 (N_4837,N_1800,N_431);
and U4838 (N_4838,N_1897,N_693);
nand U4839 (N_4839,N_194,N_774);
and U4840 (N_4840,N_1506,N_2146);
nor U4841 (N_4841,N_99,N_51);
or U4842 (N_4842,N_193,N_1273);
nor U4843 (N_4843,N_290,N_1501);
nand U4844 (N_4844,N_653,N_343);
nand U4845 (N_4845,N_1906,N_1201);
nor U4846 (N_4846,N_2017,N_1643);
or U4847 (N_4847,N_224,N_1042);
and U4848 (N_4848,N_80,N_1022);
nand U4849 (N_4849,N_2222,N_2166);
nand U4850 (N_4850,N_1465,N_10);
nand U4851 (N_4851,N_593,N_522);
or U4852 (N_4852,N_850,N_2082);
and U4853 (N_4853,N_1710,N_724);
and U4854 (N_4854,N_12,N_839);
and U4855 (N_4855,N_1514,N_1305);
or U4856 (N_4856,N_1213,N_839);
nor U4857 (N_4857,N_219,N_1403);
and U4858 (N_4858,N_899,N_1347);
nand U4859 (N_4859,N_1226,N_1458);
or U4860 (N_4860,N_440,N_789);
or U4861 (N_4861,N_1562,N_1178);
or U4862 (N_4862,N_2012,N_1235);
nand U4863 (N_4863,N_2367,N_1228);
and U4864 (N_4864,N_45,N_1253);
and U4865 (N_4865,N_2223,N_15);
and U4866 (N_4866,N_1022,N_1157);
nor U4867 (N_4867,N_2243,N_627);
nor U4868 (N_4868,N_859,N_1418);
nor U4869 (N_4869,N_705,N_460);
nand U4870 (N_4870,N_200,N_2022);
nor U4871 (N_4871,N_791,N_982);
or U4872 (N_4872,N_2196,N_2411);
nand U4873 (N_4873,N_127,N_1566);
or U4874 (N_4874,N_286,N_2347);
and U4875 (N_4875,N_990,N_1628);
nor U4876 (N_4876,N_1000,N_1371);
nand U4877 (N_4877,N_582,N_1252);
or U4878 (N_4878,N_803,N_998);
nand U4879 (N_4879,N_1396,N_119);
nor U4880 (N_4880,N_817,N_1670);
or U4881 (N_4881,N_471,N_2182);
and U4882 (N_4882,N_337,N_308);
or U4883 (N_4883,N_459,N_111);
nor U4884 (N_4884,N_2394,N_599);
or U4885 (N_4885,N_2376,N_677);
nor U4886 (N_4886,N_430,N_524);
nand U4887 (N_4887,N_2469,N_1093);
and U4888 (N_4888,N_8,N_838);
nand U4889 (N_4889,N_1486,N_1272);
and U4890 (N_4890,N_1411,N_1211);
nor U4891 (N_4891,N_2260,N_763);
nor U4892 (N_4892,N_1111,N_1580);
or U4893 (N_4893,N_343,N_2352);
or U4894 (N_4894,N_264,N_241);
nor U4895 (N_4895,N_1838,N_1666);
or U4896 (N_4896,N_1545,N_2257);
and U4897 (N_4897,N_836,N_1736);
nor U4898 (N_4898,N_704,N_564);
and U4899 (N_4899,N_2215,N_203);
xor U4900 (N_4900,N_1524,N_1884);
or U4901 (N_4901,N_225,N_1944);
nor U4902 (N_4902,N_1189,N_1012);
or U4903 (N_4903,N_432,N_1356);
and U4904 (N_4904,N_2419,N_487);
nand U4905 (N_4905,N_1963,N_1421);
and U4906 (N_4906,N_2338,N_707);
or U4907 (N_4907,N_1204,N_1760);
or U4908 (N_4908,N_1874,N_109);
nor U4909 (N_4909,N_1558,N_923);
and U4910 (N_4910,N_1269,N_1970);
nand U4911 (N_4911,N_2411,N_1151);
nor U4912 (N_4912,N_672,N_1527);
or U4913 (N_4913,N_2021,N_2479);
nor U4914 (N_4914,N_2373,N_2023);
nand U4915 (N_4915,N_2261,N_268);
or U4916 (N_4916,N_1161,N_1738);
nand U4917 (N_4917,N_1490,N_601);
and U4918 (N_4918,N_824,N_773);
or U4919 (N_4919,N_2033,N_1962);
nor U4920 (N_4920,N_400,N_1080);
nand U4921 (N_4921,N_2234,N_1715);
or U4922 (N_4922,N_1181,N_222);
nor U4923 (N_4923,N_868,N_395);
or U4924 (N_4924,N_10,N_590);
or U4925 (N_4925,N_772,N_165);
and U4926 (N_4926,N_688,N_425);
and U4927 (N_4927,N_1074,N_2397);
nand U4928 (N_4928,N_1817,N_627);
nand U4929 (N_4929,N_579,N_1869);
or U4930 (N_4930,N_31,N_1616);
or U4931 (N_4931,N_494,N_222);
or U4932 (N_4932,N_1960,N_977);
and U4933 (N_4933,N_289,N_811);
or U4934 (N_4934,N_1684,N_2429);
and U4935 (N_4935,N_1763,N_1439);
nand U4936 (N_4936,N_780,N_1991);
nand U4937 (N_4937,N_302,N_2113);
or U4938 (N_4938,N_1375,N_561);
or U4939 (N_4939,N_362,N_2081);
or U4940 (N_4940,N_2385,N_1707);
or U4941 (N_4941,N_1093,N_2488);
or U4942 (N_4942,N_446,N_380);
nor U4943 (N_4943,N_1180,N_546);
and U4944 (N_4944,N_24,N_2330);
nand U4945 (N_4945,N_1070,N_204);
and U4946 (N_4946,N_610,N_428);
or U4947 (N_4947,N_810,N_1181);
nor U4948 (N_4948,N_2277,N_2320);
nor U4949 (N_4949,N_523,N_265);
and U4950 (N_4950,N_1160,N_509);
nand U4951 (N_4951,N_2062,N_529);
nand U4952 (N_4952,N_483,N_2314);
nand U4953 (N_4953,N_1597,N_2455);
nor U4954 (N_4954,N_1445,N_797);
and U4955 (N_4955,N_1774,N_569);
and U4956 (N_4956,N_1799,N_994);
nand U4957 (N_4957,N_811,N_874);
or U4958 (N_4958,N_747,N_2326);
nand U4959 (N_4959,N_1581,N_686);
nand U4960 (N_4960,N_171,N_1976);
and U4961 (N_4961,N_520,N_654);
or U4962 (N_4962,N_1456,N_181);
and U4963 (N_4963,N_424,N_2390);
nand U4964 (N_4964,N_572,N_1994);
or U4965 (N_4965,N_653,N_1769);
nand U4966 (N_4966,N_2456,N_292);
or U4967 (N_4967,N_1292,N_2195);
nor U4968 (N_4968,N_1513,N_472);
nand U4969 (N_4969,N_725,N_1537);
or U4970 (N_4970,N_1676,N_1981);
and U4971 (N_4971,N_470,N_2449);
nor U4972 (N_4972,N_1473,N_315);
xnor U4973 (N_4973,N_88,N_1616);
or U4974 (N_4974,N_1076,N_467);
and U4975 (N_4975,N_1152,N_582);
and U4976 (N_4976,N_398,N_118);
nor U4977 (N_4977,N_2196,N_2099);
and U4978 (N_4978,N_2389,N_46);
nand U4979 (N_4979,N_1884,N_2072);
or U4980 (N_4980,N_1625,N_164);
and U4981 (N_4981,N_2341,N_962);
nor U4982 (N_4982,N_2272,N_1132);
nor U4983 (N_4983,N_381,N_1447);
nand U4984 (N_4984,N_74,N_1950);
nor U4985 (N_4985,N_1217,N_663);
or U4986 (N_4986,N_605,N_427);
and U4987 (N_4987,N_1485,N_1464);
xor U4988 (N_4988,N_1065,N_1397);
nand U4989 (N_4989,N_1940,N_1254);
nor U4990 (N_4990,N_2272,N_1484);
or U4991 (N_4991,N_1738,N_479);
or U4992 (N_4992,N_2133,N_921);
and U4993 (N_4993,N_494,N_254);
nor U4994 (N_4994,N_302,N_258);
nand U4995 (N_4995,N_1936,N_1572);
or U4996 (N_4996,N_2180,N_1731);
xnor U4997 (N_4997,N_1276,N_935);
nor U4998 (N_4998,N_100,N_2466);
nand U4999 (N_4999,N_1386,N_2367);
and U5000 (N_5000,N_3641,N_4931);
nand U5001 (N_5001,N_3888,N_3497);
nor U5002 (N_5002,N_3133,N_3723);
nand U5003 (N_5003,N_3877,N_4094);
or U5004 (N_5004,N_4993,N_3819);
and U5005 (N_5005,N_4956,N_4191);
nand U5006 (N_5006,N_4824,N_2999);
nand U5007 (N_5007,N_3168,N_2879);
and U5008 (N_5008,N_4489,N_3252);
and U5009 (N_5009,N_2969,N_2997);
nor U5010 (N_5010,N_2900,N_3079);
nor U5011 (N_5011,N_3177,N_2938);
nand U5012 (N_5012,N_4122,N_2635);
and U5013 (N_5013,N_4414,N_4646);
and U5014 (N_5014,N_2606,N_4878);
or U5015 (N_5015,N_4999,N_4220);
and U5016 (N_5016,N_4137,N_4703);
nand U5017 (N_5017,N_4350,N_4452);
and U5018 (N_5018,N_4718,N_4011);
nor U5019 (N_5019,N_3280,N_3323);
or U5020 (N_5020,N_4717,N_4654);
and U5021 (N_5021,N_4057,N_3969);
and U5022 (N_5022,N_2696,N_4208);
nand U5023 (N_5023,N_3044,N_4495);
nor U5024 (N_5024,N_3910,N_2640);
nand U5025 (N_5025,N_3410,N_4987);
nor U5026 (N_5026,N_4830,N_3814);
nand U5027 (N_5027,N_3749,N_3435);
nand U5028 (N_5028,N_3999,N_3930);
or U5029 (N_5029,N_4304,N_3573);
or U5030 (N_5030,N_3450,N_2919);
or U5031 (N_5031,N_2810,N_4986);
and U5032 (N_5032,N_4124,N_3439);
and U5033 (N_5033,N_2745,N_3867);
or U5034 (N_5034,N_4207,N_4473);
nor U5035 (N_5035,N_4801,N_3832);
xor U5036 (N_5036,N_4571,N_3859);
nor U5037 (N_5037,N_4880,N_2828);
xnor U5038 (N_5038,N_3895,N_3717);
and U5039 (N_5039,N_4439,N_2758);
and U5040 (N_5040,N_4021,N_4252);
and U5041 (N_5041,N_4896,N_4580);
or U5042 (N_5042,N_3121,N_4943);
nand U5043 (N_5043,N_2722,N_3100);
or U5044 (N_5044,N_3824,N_4401);
nand U5045 (N_5045,N_2764,N_3889);
nand U5046 (N_5046,N_3583,N_2675);
nand U5047 (N_5047,N_3666,N_4596);
or U5048 (N_5048,N_2930,N_2871);
nor U5049 (N_5049,N_3748,N_3447);
or U5050 (N_5050,N_4831,N_4116);
nand U5051 (N_5051,N_4155,N_4685);
nand U5052 (N_5052,N_2676,N_3791);
or U5053 (N_5053,N_4766,N_3065);
or U5054 (N_5054,N_2870,N_4714);
nor U5055 (N_5055,N_4295,N_4212);
or U5056 (N_5056,N_3746,N_4003);
and U5057 (N_5057,N_3099,N_2680);
nand U5058 (N_5058,N_3524,N_4677);
and U5059 (N_5059,N_3631,N_4935);
and U5060 (N_5060,N_4584,N_4146);
nor U5061 (N_5061,N_3765,N_3549);
or U5062 (N_5062,N_3984,N_2724);
nand U5063 (N_5063,N_4501,N_4805);
and U5064 (N_5064,N_4171,N_4074);
nand U5065 (N_5065,N_4297,N_3325);
or U5066 (N_5066,N_4835,N_3123);
or U5067 (N_5067,N_4623,N_3212);
nor U5068 (N_5068,N_4932,N_4399);
nand U5069 (N_5069,N_3516,N_3001);
nor U5070 (N_5070,N_3764,N_2612);
or U5071 (N_5071,N_4249,N_4921);
nand U5072 (N_5072,N_2562,N_2654);
nand U5073 (N_5073,N_3361,N_3346);
nor U5074 (N_5074,N_2704,N_3394);
and U5075 (N_5075,N_4756,N_4579);
or U5076 (N_5076,N_4325,N_2929);
nand U5077 (N_5077,N_3064,N_3866);
and U5078 (N_5078,N_4451,N_2712);
and U5079 (N_5079,N_4110,N_3973);
nand U5080 (N_5080,N_4474,N_4069);
and U5081 (N_5081,N_3444,N_3313);
and U5082 (N_5082,N_4741,N_3585);
or U5083 (N_5083,N_4416,N_4841);
nand U5084 (N_5084,N_3574,N_4961);
nor U5085 (N_5085,N_4858,N_3070);
and U5086 (N_5086,N_4875,N_3520);
or U5087 (N_5087,N_3779,N_2840);
nand U5088 (N_5088,N_3826,N_4376);
nand U5089 (N_5089,N_4920,N_4668);
or U5090 (N_5090,N_4251,N_4803);
and U5091 (N_5091,N_4839,N_2622);
and U5092 (N_5092,N_4159,N_2743);
nand U5093 (N_5093,N_3965,N_3327);
and U5094 (N_5094,N_4898,N_4335);
and U5095 (N_5095,N_4959,N_2805);
nor U5096 (N_5096,N_2595,N_2974);
nand U5097 (N_5097,N_4713,N_4198);
or U5098 (N_5098,N_4360,N_3699);
or U5099 (N_5099,N_4090,N_2799);
or U5100 (N_5100,N_3363,N_3909);
nor U5101 (N_5101,N_3543,N_3809);
and U5102 (N_5102,N_3425,N_2509);
xor U5103 (N_5103,N_4503,N_4353);
nor U5104 (N_5104,N_3935,N_3982);
nor U5105 (N_5105,N_4022,N_4265);
or U5106 (N_5106,N_2829,N_2859);
or U5107 (N_5107,N_3002,N_4261);
and U5108 (N_5108,N_3802,N_4789);
and U5109 (N_5109,N_4586,N_4050);
and U5110 (N_5110,N_3554,N_3357);
nand U5111 (N_5111,N_2842,N_2520);
or U5112 (N_5112,N_2911,N_2707);
nand U5113 (N_5113,N_2729,N_3382);
and U5114 (N_5114,N_4092,N_3381);
and U5115 (N_5115,N_4924,N_4112);
and U5116 (N_5116,N_4675,N_2699);
nor U5117 (N_5117,N_4427,N_4412);
and U5118 (N_5118,N_2601,N_3372);
or U5119 (N_5119,N_3944,N_3250);
nand U5120 (N_5120,N_4760,N_4462);
and U5121 (N_5121,N_4989,N_4828);
nor U5122 (N_5122,N_3446,N_4711);
nand U5123 (N_5123,N_3249,N_2683);
and U5124 (N_5124,N_4281,N_3436);
or U5125 (N_5125,N_4247,N_4377);
or U5126 (N_5126,N_4380,N_4150);
nand U5127 (N_5127,N_4477,N_3108);
and U5128 (N_5128,N_2695,N_3232);
or U5129 (N_5129,N_3606,N_3753);
nor U5130 (N_5130,N_4197,N_3513);
nand U5131 (N_5131,N_3196,N_3747);
nor U5132 (N_5132,N_4510,N_4779);
nand U5133 (N_5133,N_4179,N_4078);
or U5134 (N_5134,N_4844,N_2822);
or U5135 (N_5135,N_4899,N_2800);
xor U5136 (N_5136,N_3883,N_3928);
nand U5137 (N_5137,N_3651,N_3304);
and U5138 (N_5138,N_4909,N_3676);
nor U5139 (N_5139,N_4188,N_4186);
nand U5140 (N_5140,N_3551,N_2843);
or U5141 (N_5141,N_2978,N_3236);
nand U5142 (N_5142,N_4341,N_3614);
and U5143 (N_5143,N_3616,N_2577);
nand U5144 (N_5144,N_4937,N_2710);
nand U5145 (N_5145,N_2964,N_4973);
or U5146 (N_5146,N_4610,N_4118);
xnor U5147 (N_5147,N_3593,N_2660);
nor U5148 (N_5148,N_3577,N_3563);
and U5149 (N_5149,N_4240,N_2542);
nand U5150 (N_5150,N_4939,N_4772);
or U5151 (N_5151,N_3667,N_3091);
nand U5152 (N_5152,N_2760,N_3953);
or U5153 (N_5153,N_3078,N_3190);
or U5154 (N_5154,N_4838,N_4990);
nor U5155 (N_5155,N_4816,N_3509);
and U5156 (N_5156,N_4859,N_2659);
or U5157 (N_5157,N_2645,N_4199);
nand U5158 (N_5158,N_4933,N_3892);
nand U5159 (N_5159,N_3668,N_3544);
nor U5160 (N_5160,N_3798,N_3061);
nor U5161 (N_5161,N_4854,N_4827);
nor U5162 (N_5162,N_2526,N_4131);
xor U5163 (N_5163,N_4291,N_4100);
nand U5164 (N_5164,N_2567,N_4497);
xor U5165 (N_5165,N_4177,N_3374);
nor U5166 (N_5166,N_4565,N_2573);
nor U5167 (N_5167,N_3929,N_3522);
and U5168 (N_5168,N_2594,N_4324);
nor U5169 (N_5169,N_4244,N_3630);
nand U5170 (N_5170,N_3769,N_2820);
and U5171 (N_5171,N_4869,N_4071);
or U5172 (N_5172,N_3318,N_2797);
nor U5173 (N_5173,N_4782,N_4355);
or U5174 (N_5174,N_4849,N_3501);
nor U5175 (N_5175,N_4085,N_3617);
nor U5176 (N_5176,N_3800,N_4715);
or U5177 (N_5177,N_3299,N_4997);
nor U5178 (N_5178,N_3916,N_3480);
nor U5179 (N_5179,N_2772,N_4306);
or U5180 (N_5180,N_4845,N_4906);
and U5181 (N_5181,N_3947,N_3030);
and U5182 (N_5182,N_4808,N_4576);
nor U5183 (N_5183,N_4905,N_4895);
nand U5184 (N_5184,N_3546,N_4248);
or U5185 (N_5185,N_3339,N_3660);
nor U5186 (N_5186,N_3245,N_3691);
and U5187 (N_5187,N_2623,N_3499);
nand U5188 (N_5188,N_2563,N_3740);
nand U5189 (N_5189,N_3580,N_4445);
nand U5190 (N_5190,N_3156,N_4702);
nor U5191 (N_5191,N_3247,N_2811);
nor U5192 (N_5192,N_2952,N_3828);
or U5193 (N_5193,N_3985,N_4447);
nand U5194 (N_5194,N_3876,N_4228);
nand U5195 (N_5195,N_3907,N_2546);
and U5196 (N_5196,N_3272,N_3251);
or U5197 (N_5197,N_4874,N_4476);
nand U5198 (N_5198,N_2928,N_2987);
nor U5199 (N_5199,N_3602,N_2538);
nor U5200 (N_5200,N_2559,N_3961);
nor U5201 (N_5201,N_4558,N_2806);
or U5202 (N_5202,N_2834,N_4486);
or U5203 (N_5203,N_4384,N_4628);
nand U5204 (N_5204,N_4746,N_4161);
and U5205 (N_5205,N_4561,N_4488);
or U5206 (N_5206,N_4234,N_4075);
and U5207 (N_5207,N_4966,N_3882);
or U5208 (N_5208,N_4542,N_3781);
or U5209 (N_5209,N_2851,N_3636);
nor U5210 (N_5210,N_2715,N_4876);
nor U5211 (N_5211,N_4910,N_4136);
or U5212 (N_5212,N_4152,N_2586);
or U5213 (N_5213,N_3193,N_4867);
and U5214 (N_5214,N_4980,N_3950);
nand U5215 (N_5215,N_3370,N_3209);
and U5216 (N_5216,N_2816,N_3204);
nand U5217 (N_5217,N_4908,N_2548);
or U5218 (N_5218,N_3127,N_2768);
and U5219 (N_5219,N_3017,N_3467);
or U5220 (N_5220,N_4217,N_2697);
or U5221 (N_5221,N_3278,N_4053);
nor U5222 (N_5222,N_4018,N_2592);
nor U5223 (N_5223,N_2847,N_3937);
or U5224 (N_5224,N_4557,N_3797);
nor U5225 (N_5225,N_3763,N_3460);
nor U5226 (N_5226,N_3288,N_4286);
and U5227 (N_5227,N_4115,N_2524);
xnor U5228 (N_5228,N_4870,N_4795);
and U5229 (N_5229,N_2801,N_2527);
and U5230 (N_5230,N_3992,N_2587);
nand U5231 (N_5231,N_2720,N_4688);
or U5232 (N_5232,N_4106,N_3365);
xnor U5233 (N_5233,N_4499,N_3548);
or U5234 (N_5234,N_2866,N_4385);
nand U5235 (N_5235,N_3788,N_3956);
nand U5236 (N_5236,N_4695,N_4241);
nand U5237 (N_5237,N_3322,N_3507);
and U5238 (N_5238,N_4314,N_3377);
or U5239 (N_5239,N_4851,N_4707);
nor U5240 (N_5240,N_2804,N_2609);
nor U5241 (N_5241,N_2510,N_3987);
nand U5242 (N_5242,N_4524,N_4728);
nor U5243 (N_5243,N_3682,N_3508);
nor U5244 (N_5244,N_3649,N_4026);
or U5245 (N_5245,N_2915,N_2709);
and U5246 (N_5246,N_4487,N_3671);
or U5247 (N_5247,N_3561,N_3025);
or U5248 (N_5248,N_3719,N_2888);
nor U5249 (N_5249,N_4305,N_3303);
nor U5250 (N_5250,N_4287,N_4710);
nor U5251 (N_5251,N_3075,N_2717);
and U5252 (N_5252,N_3084,N_4180);
nor U5253 (N_5253,N_2777,N_4783);
and U5254 (N_5254,N_4806,N_4383);
and U5255 (N_5255,N_2955,N_3933);
or U5256 (N_5256,N_3042,N_4464);
nor U5257 (N_5257,N_4166,N_2904);
and U5258 (N_5258,N_4308,N_3292);
nand U5259 (N_5259,N_2590,N_3489);
or U5260 (N_5260,N_4031,N_4968);
nand U5261 (N_5261,N_3459,N_3172);
nor U5262 (N_5262,N_4555,N_4975);
nor U5263 (N_5263,N_2740,N_3035);
and U5264 (N_5264,N_3355,N_3305);
and U5265 (N_5265,N_4818,N_4960);
and U5266 (N_5266,N_4045,N_3423);
or U5267 (N_5267,N_3986,N_4575);
nor U5268 (N_5268,N_4449,N_4523);
and U5269 (N_5269,N_4002,N_2674);
and U5270 (N_5270,N_2534,N_2950);
or U5271 (N_5271,N_3060,N_4914);
nand U5272 (N_5272,N_4658,N_4538);
nand U5273 (N_5273,N_3852,N_3487);
or U5274 (N_5274,N_4769,N_4629);
nor U5275 (N_5275,N_4201,N_3290);
or U5276 (N_5276,N_4420,N_2837);
nand U5277 (N_5277,N_4358,N_4096);
and U5278 (N_5278,N_3286,N_3417);
xor U5279 (N_5279,N_4005,N_3805);
or U5280 (N_5280,N_2815,N_4748);
and U5281 (N_5281,N_4992,N_4700);
nor U5282 (N_5282,N_2626,N_4598);
nand U5283 (N_5283,N_4659,N_4357);
or U5284 (N_5284,N_3197,N_4138);
nand U5285 (N_5285,N_2672,N_3920);
and U5286 (N_5286,N_3003,N_4670);
or U5287 (N_5287,N_3139,N_4024);
nor U5288 (N_5288,N_2727,N_3210);
or U5289 (N_5289,N_4536,N_4940);
or U5290 (N_5290,N_2663,N_4035);
or U5291 (N_5291,N_4267,N_4645);
nor U5292 (N_5292,N_2858,N_3378);
xnor U5293 (N_5293,N_3301,N_3657);
or U5294 (N_5294,N_3687,N_4389);
nor U5295 (N_5295,N_3348,N_2884);
or U5296 (N_5296,N_2536,N_3144);
or U5297 (N_5297,N_4317,N_2632);
nor U5298 (N_5298,N_4437,N_4332);
or U5299 (N_5299,N_4362,N_2909);
nor U5300 (N_5300,N_3309,N_3514);
and U5301 (N_5301,N_4059,N_3437);
nand U5302 (N_5302,N_3547,N_4964);
or U5303 (N_5303,N_3557,N_3398);
or U5304 (N_5304,N_4020,N_4716);
nor U5305 (N_5305,N_4065,N_3505);
or U5306 (N_5306,N_2737,N_3675);
and U5307 (N_5307,N_2962,N_3088);
or U5308 (N_5308,N_4534,N_2949);
and U5309 (N_5309,N_4151,N_3297);
nand U5310 (N_5310,N_4817,N_3506);
or U5311 (N_5311,N_3164,N_4406);
or U5312 (N_5312,N_2782,N_2682);
and U5313 (N_5313,N_4614,N_2725);
or U5314 (N_5314,N_4502,N_4417);
nand U5315 (N_5315,N_4954,N_3594);
and U5316 (N_5316,N_4603,N_4551);
nand U5317 (N_5317,N_4015,N_2633);
or U5318 (N_5318,N_2943,N_4187);
and U5319 (N_5319,N_2893,N_3291);
xnor U5320 (N_5320,N_2570,N_4902);
and U5321 (N_5321,N_3391,N_3692);
nor U5322 (N_5322,N_2852,N_4034);
nand U5323 (N_5323,N_4233,N_2788);
and U5324 (N_5324,N_4919,N_3658);
and U5325 (N_5325,N_3104,N_3120);
nor U5326 (N_5326,N_2784,N_3968);
and U5327 (N_5327,N_3008,N_4855);
and U5328 (N_5328,N_3773,N_4126);
and U5329 (N_5329,N_3142,N_4479);
nor U5330 (N_5330,N_4738,N_4893);
and U5331 (N_5331,N_2838,N_3491);
nor U5332 (N_5332,N_4130,N_4872);
or U5333 (N_5333,N_4843,N_4433);
nor U5334 (N_5334,N_4559,N_3462);
nor U5335 (N_5335,N_2670,N_3218);
nand U5336 (N_5336,N_2880,N_4904);
or U5337 (N_5337,N_3778,N_4776);
and U5338 (N_5338,N_4928,N_4771);
or U5339 (N_5339,N_4732,N_3812);
or U5340 (N_5340,N_4253,N_3205);
and U5341 (N_5341,N_3145,N_4704);
nor U5342 (N_5342,N_2896,N_4435);
nor U5343 (N_5343,N_4913,N_3165);
and U5344 (N_5344,N_4595,N_4095);
and U5345 (N_5345,N_3588,N_3534);
or U5346 (N_5346,N_3858,N_3089);
and U5347 (N_5347,N_4661,N_4923);
nand U5348 (N_5348,N_3068,N_4656);
nand U5349 (N_5349,N_3134,N_4160);
or U5350 (N_5350,N_3693,N_3643);
or U5351 (N_5351,N_4759,N_4349);
nand U5352 (N_5352,N_4519,N_4733);
nor U5353 (N_5353,N_4630,N_2890);
and U5354 (N_5354,N_4381,N_4189);
or U5355 (N_5355,N_3012,N_3380);
nand U5356 (N_5356,N_4513,N_4531);
or U5357 (N_5357,N_3970,N_4864);
nand U5358 (N_5358,N_3344,N_3787);
nand U5359 (N_5359,N_3277,N_4550);
or U5360 (N_5360,N_2667,N_3741);
nor U5361 (N_5361,N_2581,N_2841);
nor U5362 (N_5362,N_3163,N_4901);
and U5363 (N_5363,N_3925,N_3784);
and U5364 (N_5364,N_3045,N_2625);
nand U5365 (N_5365,N_2986,N_3870);
nor U5366 (N_5366,N_4915,N_4810);
and U5367 (N_5367,N_2931,N_4903);
and U5368 (N_5368,N_2600,N_2507);
and U5369 (N_5369,N_2926,N_3449);
nand U5370 (N_5370,N_4345,N_3146);
or U5371 (N_5371,N_2998,N_3285);
nand U5372 (N_5372,N_4846,N_2865);
nor U5373 (N_5373,N_3792,N_3550);
nand U5374 (N_5374,N_2966,N_4283);
nand U5375 (N_5375,N_3751,N_3863);
nand U5376 (N_5376,N_2850,N_3050);
and U5377 (N_5377,N_2604,N_3688);
or U5378 (N_5378,N_4549,N_4509);
nand U5379 (N_5379,N_2647,N_3136);
and U5380 (N_5380,N_2568,N_4952);
and U5381 (N_5381,N_2817,N_4567);
nor U5382 (N_5382,N_2642,N_3011);
or U5383 (N_5383,N_3993,N_4706);
nand U5384 (N_5384,N_4185,N_4403);
nor U5385 (N_5385,N_4260,N_4246);
and U5386 (N_5386,N_3936,N_2982);
xnor U5387 (N_5387,N_3067,N_3623);
and U5388 (N_5388,N_2849,N_4072);
nand U5389 (N_5389,N_3083,N_4883);
and U5390 (N_5390,N_4481,N_4446);
nand U5391 (N_5391,N_3428,N_2924);
or U5392 (N_5392,N_4456,N_4210);
and U5393 (N_5393,N_3371,N_4250);
or U5394 (N_5394,N_3843,N_3541);
nor U5395 (N_5395,N_3161,N_4494);
nor U5396 (N_5396,N_4336,N_4441);
or U5397 (N_5397,N_4418,N_3419);
and U5398 (N_5398,N_2831,N_3319);
nor U5399 (N_5399,N_3845,N_4890);
or U5400 (N_5400,N_3485,N_4434);
nor U5401 (N_5401,N_4684,N_3009);
nor U5402 (N_5402,N_3242,N_4258);
nor U5403 (N_5403,N_2741,N_2878);
nand U5404 (N_5404,N_4483,N_3529);
and U5405 (N_5405,N_3700,N_4237);
or U5406 (N_5406,N_3603,N_4958);
and U5407 (N_5407,N_3744,N_3839);
and U5408 (N_5408,N_4616,N_3235);
and U5409 (N_5409,N_3829,N_4029);
and U5410 (N_5410,N_3048,N_4454);
nor U5411 (N_5411,N_2689,N_4882);
nor U5412 (N_5412,N_2813,N_4653);
nor U5413 (N_5413,N_4626,N_3306);
nand U5414 (N_5414,N_3579,N_3775);
nor U5415 (N_5415,N_4047,N_3424);
nor U5416 (N_5416,N_2554,N_3466);
or U5417 (N_5417,N_4001,N_3810);
and U5418 (N_5418,N_4564,N_3601);
nand U5419 (N_5419,N_3894,N_4916);
nand U5420 (N_5420,N_3659,N_4391);
xor U5421 (N_5421,N_3915,N_4724);
nand U5422 (N_5422,N_2883,N_4066);
or U5423 (N_5423,N_3080,N_4774);
nand U5424 (N_5424,N_3206,N_3654);
nand U5425 (N_5425,N_4832,N_3393);
nor U5426 (N_5426,N_3422,N_4988);
and U5427 (N_5427,N_3931,N_3957);
and U5428 (N_5428,N_4017,N_4930);
or U5429 (N_5429,N_2917,N_3523);
nor U5430 (N_5430,N_3458,N_3640);
and U5431 (N_5431,N_3679,N_4202);
nand U5432 (N_5432,N_4039,N_4415);
nor U5433 (N_5433,N_3217,N_3756);
nor U5434 (N_5434,N_3397,N_2767);
nor U5435 (N_5435,N_4318,N_2996);
or U5436 (N_5436,N_3521,N_3566);
nor U5437 (N_5437,N_2602,N_4691);
or U5438 (N_5438,N_4813,N_3106);
and U5439 (N_5439,N_4148,N_3911);
nand U5440 (N_5440,N_3500,N_3782);
and U5441 (N_5441,N_3502,N_4133);
and U5442 (N_5442,N_3878,N_3663);
and U5443 (N_5443,N_4147,N_3409);
or U5444 (N_5444,N_4641,N_4013);
and U5445 (N_5445,N_3169,N_4238);
nand U5446 (N_5446,N_4804,N_4698);
nor U5447 (N_5447,N_3613,N_4547);
and U5448 (N_5448,N_4461,N_3492);
and U5449 (N_5449,N_4708,N_4327);
nand U5450 (N_5450,N_3567,N_4891);
nor U5451 (N_5451,N_4609,N_3420);
nor U5452 (N_5452,N_4373,N_3312);
or U5453 (N_5453,N_2814,N_4929);
and U5454 (N_5454,N_3538,N_3077);
or U5455 (N_5455,N_2571,N_3542);
nand U5456 (N_5456,N_3022,N_3571);
nand U5457 (N_5457,N_2730,N_2803);
or U5458 (N_5458,N_3401,N_3847);
and U5459 (N_5459,N_4548,N_4101);
and U5460 (N_5460,N_3673,N_4378);
and U5461 (N_5461,N_3618,N_4329);
nand U5462 (N_5462,N_4680,N_3977);
or U5463 (N_5463,N_2525,N_4140);
and U5464 (N_5464,N_2521,N_2518);
or U5465 (N_5465,N_2862,N_4761);
nand U5466 (N_5466,N_4176,N_2948);
and U5467 (N_5467,N_4262,N_3940);
and U5468 (N_5468,N_2603,N_2690);
nor U5469 (N_5469,N_4618,N_3453);
nand U5470 (N_5470,N_3581,N_3978);
nand U5471 (N_5471,N_4064,N_2941);
nand U5472 (N_5472,N_3141,N_3178);
and U5473 (N_5473,N_2531,N_3904);
nand U5474 (N_5474,N_4802,N_3665);
and U5475 (N_5475,N_3803,N_4581);
nand U5476 (N_5476,N_4156,N_2619);
and U5477 (N_5477,N_4173,N_2627);
and U5478 (N_5478,N_4877,N_4834);
nor U5479 (N_5479,N_2759,N_3015);
or U5480 (N_5480,N_3817,N_3490);
and U5481 (N_5481,N_4181,N_4257);
and U5482 (N_5482,N_2711,N_4619);
nor U5483 (N_5483,N_2971,N_4073);
nor U5484 (N_5484,N_4139,N_2618);
nor U5485 (N_5485,N_3572,N_4577);
or U5486 (N_5486,N_4387,N_3421);
nor U5487 (N_5487,N_3816,N_3525);
or U5488 (N_5488,N_4944,N_4742);
nand U5489 (N_5489,N_4585,N_2773);
or U5490 (N_5490,N_4278,N_3708);
or U5491 (N_5491,N_4861,N_4516);
nor U5492 (N_5492,N_4459,N_4276);
and U5493 (N_5493,N_3761,N_4319);
or U5494 (N_5494,N_2989,N_4084);
nand U5495 (N_5495,N_3582,N_3880);
nand U5496 (N_5496,N_4046,N_4563);
and U5497 (N_5497,N_4566,N_2983);
and U5498 (N_5498,N_4282,N_2812);
xnor U5499 (N_5499,N_4442,N_4203);
nand U5500 (N_5500,N_2839,N_3584);
nor U5501 (N_5501,N_4450,N_4272);
nor U5502 (N_5502,N_2646,N_4660);
nand U5503 (N_5503,N_2802,N_4157);
nor U5504 (N_5504,N_3310,N_4044);
and U5505 (N_5505,N_3725,N_2778);
nand U5506 (N_5506,N_2836,N_4361);
nor U5507 (N_5507,N_4570,N_3482);
or U5508 (N_5508,N_4107,N_3590);
or U5509 (N_5509,N_2705,N_2599);
nor U5510 (N_5510,N_3200,N_3884);
nor U5511 (N_5511,N_3256,N_3295);
nand U5512 (N_5512,N_2765,N_2700);
or U5513 (N_5513,N_2844,N_4709);
or U5514 (N_5514,N_4498,N_3294);
nor U5515 (N_5515,N_3387,N_4825);
and U5516 (N_5516,N_2719,N_4763);
nor U5517 (N_5517,N_2968,N_3137);
nor U5518 (N_5518,N_2585,N_3610);
and U5519 (N_5519,N_2713,N_4055);
nand U5520 (N_5520,N_3648,N_2589);
nand U5521 (N_5521,N_4048,N_4104);
and U5522 (N_5522,N_3389,N_2953);
nor U5523 (N_5523,N_3238,N_3345);
nand U5524 (N_5524,N_4730,N_3254);
nor U5525 (N_5525,N_2649,N_4222);
and U5526 (N_5526,N_4162,N_2940);
nor U5527 (N_5527,N_4583,N_3092);
or U5528 (N_5528,N_4167,N_4977);
or U5529 (N_5529,N_4856,N_2565);
nand U5530 (N_5530,N_3634,N_3455);
nand U5531 (N_5531,N_3412,N_3721);
nand U5532 (N_5532,N_4236,N_4799);
nand U5533 (N_5533,N_4099,N_3329);
nand U5534 (N_5534,N_3109,N_4873);
nor U5535 (N_5535,N_2993,N_4322);
nor U5536 (N_5536,N_4945,N_3477);
nand U5537 (N_5537,N_3283,N_4625);
nor U5538 (N_5538,N_3774,N_4164);
nand U5539 (N_5539,N_3066,N_4103);
nand U5540 (N_5540,N_2988,N_2652);
or U5541 (N_5541,N_4971,N_4316);
nor U5542 (N_5542,N_3287,N_3248);
nor U5543 (N_5543,N_4823,N_3979);
or U5544 (N_5544,N_2578,N_3821);
and U5545 (N_5545,N_3441,N_3842);
nand U5546 (N_5546,N_2819,N_2886);
nand U5547 (N_5547,N_4311,N_4109);
or U5548 (N_5548,N_3714,N_3350);
nor U5549 (N_5549,N_4592,N_3358);
nor U5550 (N_5550,N_3997,N_3539);
and U5551 (N_5551,N_3338,N_3352);
and U5552 (N_5552,N_4686,N_3710);
and U5553 (N_5553,N_3359,N_3697);
nand U5554 (N_5554,N_3029,N_4819);
nor U5555 (N_5555,N_3942,N_3101);
nand U5556 (N_5556,N_2770,N_3110);
or U5557 (N_5557,N_4028,N_3072);
or U5558 (N_5558,N_4012,N_3597);
nand U5559 (N_5559,N_4947,N_4996);
and U5560 (N_5560,N_3913,N_4466);
nor U5561 (N_5561,N_2650,N_2543);
nor U5562 (N_5562,N_4200,N_4117);
or U5563 (N_5563,N_4781,N_2925);
and U5564 (N_5564,N_3434,N_3182);
or U5565 (N_5565,N_2617,N_2979);
or U5566 (N_5566,N_3406,N_3735);
nand U5567 (N_5567,N_4484,N_4624);
nor U5568 (N_5568,N_3703,N_3224);
or U5569 (N_5569,N_4229,N_4720);
nand U5570 (N_5570,N_2785,N_3503);
nor U5571 (N_5571,N_3855,N_2681);
and U5572 (N_5572,N_4674,N_3486);
and U5573 (N_5573,N_2532,N_4342);
nand U5574 (N_5574,N_4032,N_4153);
nand U5575 (N_5575,N_2522,N_3515);
nand U5576 (N_5576,N_4347,N_4478);
nand U5577 (N_5577,N_4636,N_3922);
and U5578 (N_5578,N_3368,N_3869);
or U5579 (N_5579,N_3512,N_2608);
nand U5580 (N_5580,N_4469,N_3268);
and U5581 (N_5581,N_4395,N_2756);
or U5582 (N_5582,N_3576,N_3154);
and U5583 (N_5583,N_4729,N_4840);
and U5584 (N_5584,N_3655,N_4797);
and U5585 (N_5585,N_3385,N_3342);
nand U5586 (N_5586,N_3860,N_2854);
nand U5587 (N_5587,N_3062,N_4344);
or U5588 (N_5588,N_2588,N_4313);
nand U5589 (N_5589,N_2977,N_2721);
and U5590 (N_5590,N_3927,N_4633);
or U5591 (N_5591,N_2932,N_4254);
nor U5592 (N_5592,N_3853,N_3632);
or U5593 (N_5593,N_4976,N_4363);
and U5594 (N_5594,N_3715,N_2512);
nand U5595 (N_5595,N_4991,N_2755);
nor U5596 (N_5596,N_3416,N_3426);
nand U5597 (N_5597,N_4950,N_4227);
nor U5598 (N_5598,N_4544,N_3833);
and U5599 (N_5599,N_3240,N_3470);
nand U5600 (N_5600,N_3923,N_2679);
nor U5601 (N_5601,N_2611,N_3518);
or U5602 (N_5602,N_4465,N_4455);
nor U5603 (N_5603,N_4601,N_3672);
nor U5604 (N_5604,N_4209,N_3991);
or U5605 (N_5605,N_4863,N_2872);
and U5606 (N_5606,N_4271,N_4860);
and U5607 (N_5607,N_3071,N_2575);
and U5608 (N_5608,N_4040,N_2726);
nand U5609 (N_5609,N_2651,N_3259);
and U5610 (N_5610,N_3716,N_3914);
nor U5611 (N_5611,N_4632,N_4871);
xnor U5612 (N_5612,N_3625,N_4663);
nor U5613 (N_5613,N_3604,N_3684);
or U5614 (N_5614,N_4673,N_4621);
and U5615 (N_5615,N_4183,N_3258);
nor U5616 (N_5616,N_2656,N_2776);
and U5617 (N_5617,N_2787,N_3478);
and U5618 (N_5618,N_4129,N_4573);
nand U5619 (N_5619,N_3041,N_4836);
and U5620 (N_5620,N_3028,N_3330);
and U5621 (N_5621,N_4517,N_3191);
and U5622 (N_5622,N_2661,N_2639);
or U5623 (N_5623,N_2691,N_3369);
nor U5624 (N_5624,N_4485,N_4400);
or U5625 (N_5625,N_3262,N_4230);
xor U5626 (N_5626,N_4507,N_3140);
or U5627 (N_5627,N_3456,N_3018);
or U5628 (N_5628,N_4879,N_3498);
and U5629 (N_5629,N_3989,N_4552);
nor U5630 (N_5630,N_3027,N_4635);
nand U5631 (N_5631,N_3754,N_2687);
or U5632 (N_5632,N_3900,N_4255);
nand U5633 (N_5633,N_4128,N_2789);
nand U5634 (N_5634,N_3528,N_4374);
or U5635 (N_5635,N_3886,N_3366);
or U5636 (N_5636,N_4290,N_3938);
and U5637 (N_5637,N_4505,N_3463);
nor U5638 (N_5638,N_2994,N_4727);
nor U5639 (N_5639,N_4881,N_4239);
or U5640 (N_5640,N_4942,N_2540);
nand U5641 (N_5641,N_4008,N_4372);
and U5642 (N_5642,N_4812,N_3811);
and U5643 (N_5643,N_3155,N_3995);
nor U5644 (N_5644,N_3021,N_4512);
nor U5645 (N_5645,N_2791,N_4453);
or U5646 (N_5646,N_3750,N_4888);
nand U5647 (N_5647,N_3452,N_3694);
and U5648 (N_5648,N_4590,N_2684);
nand U5649 (N_5649,N_4539,N_4182);
and U5650 (N_5650,N_3527,N_4821);
or U5651 (N_5651,N_4734,N_2808);
or U5652 (N_5652,N_4925,N_2569);
nand U5653 (N_5653,N_3102,N_3559);
or U5654 (N_5654,N_4411,N_3712);
and U5655 (N_5655,N_3536,N_3386);
nand U5656 (N_5656,N_4515,N_3116);
or U5657 (N_5657,N_3234,N_2933);
nor U5658 (N_5658,N_4850,N_4886);
nand U5659 (N_5659,N_4299,N_4206);
and U5660 (N_5660,N_4651,N_3905);
nor U5661 (N_5661,N_2792,N_4574);
and U5662 (N_5662,N_2641,N_3861);
nand U5663 (N_5663,N_4277,N_4528);
and U5664 (N_5664,N_2502,N_4370);
and U5665 (N_5665,N_4736,N_3587);
nor U5666 (N_5666,N_4520,N_4444);
nand U5667 (N_5667,N_4773,N_3768);
or U5668 (N_5668,N_2855,N_2686);
nor U5669 (N_5669,N_2972,N_4682);
nand U5670 (N_5670,N_4853,N_3759);
or U5671 (N_5671,N_3353,N_2832);
or U5672 (N_5672,N_4794,N_3074);
or U5673 (N_5673,N_3646,N_2762);
or U5674 (N_5674,N_3105,N_3239);
or U5675 (N_5675,N_4848,N_3039);
and U5676 (N_5676,N_3388,N_4671);
nor U5677 (N_5677,N_3135,N_4457);
nand U5678 (N_5678,N_2643,N_4936);
and U5679 (N_5679,N_4725,N_4025);
and U5680 (N_5680,N_3427,N_2742);
and U5681 (N_5681,N_2666,N_4052);
nor U5682 (N_5682,N_3052,N_4270);
nand U5683 (N_5683,N_4170,N_4080);
or U5684 (N_5684,N_3608,N_4953);
nor U5685 (N_5685,N_4540,N_2673);
nor U5686 (N_5686,N_3758,N_3082);
or U5687 (N_5687,N_2965,N_3983);
nor U5688 (N_5688,N_4422,N_4303);
nor U5689 (N_5689,N_3595,N_4647);
or U5690 (N_5690,N_3282,N_3117);
nor U5691 (N_5691,N_3570,N_4375);
and U5692 (N_5692,N_3334,N_3152);
and U5693 (N_5693,N_3408,N_4154);
and U5694 (N_5694,N_2942,N_3565);
nand U5695 (N_5695,N_3820,N_3231);
or U5696 (N_5696,N_2769,N_4460);
and U5697 (N_5697,N_3331,N_4897);
and U5698 (N_5698,N_3941,N_4791);
nor U5699 (N_5699,N_3096,N_4889);
nor U5700 (N_5700,N_4884,N_4847);
or U5701 (N_5701,N_2867,N_4144);
or U5702 (N_5702,N_3726,N_3998);
nand U5703 (N_5703,N_3149,N_3849);
nand U5704 (N_5704,N_3734,N_3228);
or U5705 (N_5705,N_3429,N_3376);
nand U5706 (N_5706,N_2937,N_2610);
nand U5707 (N_5707,N_4979,N_3187);
or U5708 (N_5708,N_4852,N_2885);
or U5709 (N_5709,N_3461,N_3639);
and U5710 (N_5710,N_2936,N_4857);
and U5711 (N_5711,N_3879,N_3054);
or U5712 (N_5712,N_3488,N_2500);
nand U5713 (N_5713,N_3107,N_3246);
and U5714 (N_5714,N_2576,N_4405);
or U5715 (N_5715,N_3556,N_2796);
nand U5716 (N_5716,N_3276,N_2749);
nand U5717 (N_5717,N_2550,N_3799);
and U5718 (N_5718,N_2903,N_3519);
or U5719 (N_5719,N_3194,N_3674);
or U5720 (N_5720,N_4696,N_4293);
or U5721 (N_5721,N_4033,N_3864);
or U5722 (N_5722,N_4301,N_3851);
and U5723 (N_5723,N_3037,N_2583);
nand U5724 (N_5724,N_4393,N_4232);
and U5725 (N_5725,N_3848,N_3724);
and U5726 (N_5726,N_2564,N_4600);
nand U5727 (N_5727,N_2959,N_3122);
or U5728 (N_5728,N_3707,N_2856);
nand U5729 (N_5729,N_3830,N_4951);
nor U5730 (N_5730,N_4119,N_4334);
nand U5731 (N_5731,N_3229,N_3990);
and U5732 (N_5732,N_3939,N_3822);
nor U5733 (N_5733,N_2754,N_4587);
nor U5734 (N_5734,N_3119,N_3786);
nor U5735 (N_5735,N_3468,N_4582);
and U5736 (N_5736,N_3945,N_3263);
and U5737 (N_5737,N_4701,N_4086);
or U5738 (N_5738,N_4294,N_3713);
and U5739 (N_5739,N_4588,N_3738);
or U5740 (N_5740,N_3834,N_3016);
or U5741 (N_5741,N_3362,N_4693);
or U5742 (N_5742,N_3085,N_4787);
nand U5743 (N_5743,N_4320,N_3418);
nor U5744 (N_5744,N_4114,N_3340);
or U5745 (N_5745,N_2733,N_2889);
nor U5746 (N_5746,N_3006,N_3215);
nor U5747 (N_5747,N_4125,N_4721);
nor U5748 (N_5748,N_4424,N_3934);
or U5749 (N_5749,N_4767,N_3103);
or U5750 (N_5750,N_3780,N_4744);
or U5751 (N_5751,N_2898,N_2698);
nor U5752 (N_5752,N_4321,N_2818);
nor U5753 (N_5753,N_3948,N_4504);
nand U5754 (N_5754,N_4611,N_3157);
and U5755 (N_5755,N_3611,N_4667);
nand U5756 (N_5756,N_4121,N_3451);
or U5757 (N_5757,N_2596,N_4737);
and U5758 (N_5758,N_3296,N_3411);
nor U5759 (N_5759,N_4527,N_2980);
or U5760 (N_5760,N_4784,N_4428);
and U5761 (N_5761,N_3056,N_3128);
nand U5762 (N_5762,N_3564,N_4762);
and U5763 (N_5763,N_4266,N_2708);
nand U5764 (N_5764,N_4102,N_3532);
nand U5765 (N_5765,N_3924,N_4837);
nand U5766 (N_5766,N_2628,N_4396);
or U5767 (N_5767,N_4016,N_3183);
nand U5768 (N_5768,N_3143,N_3881);
nor U5769 (N_5769,N_2825,N_2976);
nor U5770 (N_5770,N_3599,N_2863);
nor U5771 (N_5771,N_4617,N_3762);
nor U5772 (N_5772,N_3967,N_2739);
nand U5773 (N_5773,N_4007,N_3598);
nand U5774 (N_5774,N_3808,N_2752);
nand U5775 (N_5775,N_4946,N_3202);
or U5776 (N_5776,N_3825,N_2529);
or U5777 (N_5777,N_3827,N_4337);
xor U5778 (N_5778,N_4158,N_2503);
nand U5779 (N_5779,N_3448,N_4274);
nor U5780 (N_5780,N_4205,N_4842);
nand U5781 (N_5781,N_3988,N_4382);
nand U5782 (N_5782,N_3794,N_4612);
and U5783 (N_5783,N_2795,N_3356);
nor U5784 (N_5784,N_3207,N_3328);
and U5785 (N_5785,N_3815,N_2621);
nand U5786 (N_5786,N_3341,N_3772);
or U5787 (N_5787,N_3302,N_4365);
or U5788 (N_5788,N_3150,N_2701);
and U5789 (N_5789,N_2922,N_3266);
and U5790 (N_5790,N_4692,N_3912);
and U5791 (N_5791,N_3629,N_3678);
and U5792 (N_5792,N_4699,N_4726);
nor U5793 (N_5793,N_3901,N_2723);
or U5794 (N_5794,N_3615,N_3545);
nor U5795 (N_5795,N_3495,N_2874);
nor U5796 (N_5796,N_3414,N_3966);
or U5797 (N_5797,N_4687,N_3442);
and U5798 (N_5798,N_2557,N_4087);
or U5799 (N_5799,N_3036,N_2934);
or U5800 (N_5800,N_2973,N_4719);
nor U5801 (N_5801,N_4108,N_4775);
nor U5802 (N_5802,N_4604,N_4785);
nand U5803 (N_5803,N_4004,N_3273);
nand U5804 (N_5804,N_3237,N_4038);
nor U5805 (N_5805,N_3955,N_4640);
and U5806 (N_5806,N_4404,N_4493);
nor U5807 (N_5807,N_4049,N_4900);
nand U5808 (N_5808,N_3689,N_3173);
nor U5809 (N_5809,N_3014,N_3926);
and U5810 (N_5810,N_4471,N_3317);
and U5811 (N_5811,N_4368,N_3138);
nor U5812 (N_5812,N_2957,N_3404);
or U5813 (N_5813,N_3896,N_4068);
nand U5814 (N_5814,N_3586,N_3841);
nand U5815 (N_5815,N_3354,N_4754);
or U5816 (N_5816,N_2916,N_4556);
nand U5817 (N_5817,N_4765,N_3652);
or U5818 (N_5818,N_3776,N_2905);
or U5819 (N_5819,N_2706,N_3094);
and U5820 (N_5820,N_2914,N_4448);
nand U5821 (N_5821,N_3718,N_2860);
or U5822 (N_5822,N_3026,N_4429);
nor U5823 (N_5823,N_2582,N_2636);
nand U5824 (N_5824,N_3494,N_3375);
or U5825 (N_5825,N_3890,N_2620);
nand U5826 (N_5826,N_3701,N_4615);
or U5827 (N_5827,N_3081,N_4364);
or U5828 (N_5828,N_4354,N_4390);
or U5829 (N_5829,N_3223,N_4955);
and U5830 (N_5830,N_2506,N_3257);
or U5831 (N_5831,N_4572,N_2823);
nor U5832 (N_5832,N_4010,N_3186);
or U5833 (N_5833,N_4093,N_2638);
and U5834 (N_5834,N_3131,N_3661);
nand U5835 (N_5835,N_4315,N_3745);
and U5836 (N_5836,N_3269,N_4535);
nor U5837 (N_5837,N_2669,N_4982);
or U5838 (N_5838,N_4338,N_2523);
nor U5839 (N_5839,N_4491,N_3430);
nand U5840 (N_5840,N_3804,N_3115);
or U5841 (N_5841,N_4666,N_3474);
nand U5842 (N_5842,N_3076,N_3343);
nand U5843 (N_5843,N_2881,N_3475);
nand U5844 (N_5844,N_4822,N_4111);
and U5845 (N_5845,N_2945,N_3885);
and U5846 (N_5846,N_2613,N_4907);
nand U5847 (N_5847,N_4545,N_3952);
nor U5848 (N_5848,N_4597,N_3619);
nand U5849 (N_5849,N_4218,N_2703);
or U5850 (N_5850,N_3111,N_4042);
or U5851 (N_5851,N_4149,N_3171);
and U5852 (N_5852,N_2607,N_4712);
or U5853 (N_5853,N_4431,N_3130);
nor U5854 (N_5854,N_2637,N_2809);
or U5855 (N_5855,N_4568,N_4312);
nand U5856 (N_5856,N_4672,N_2946);
and U5857 (N_5857,N_3069,N_3727);
and U5858 (N_5858,N_4269,N_2763);
nor U5859 (N_5859,N_3504,N_3321);
nor U5860 (N_5860,N_3695,N_2954);
or U5861 (N_5861,N_4231,N_4178);
nor U5862 (N_5862,N_2552,N_3255);
nand U5863 (N_5863,N_2793,N_4225);
and U5864 (N_5864,N_4432,N_2566);
and U5865 (N_5865,N_4268,N_3963);
nand U5866 (N_5866,N_3980,N_2960);
nor U5867 (N_5867,N_4408,N_3510);
and U5868 (N_5868,N_4780,N_3949);
and U5869 (N_5869,N_4062,N_4135);
and U5870 (N_5870,N_4941,N_4397);
nand U5871 (N_5871,N_3396,N_4522);
nor U5872 (N_5872,N_2985,N_2653);
or U5873 (N_5873,N_2665,N_4091);
nor U5874 (N_5874,N_4120,N_4560);
or U5875 (N_5875,N_2906,N_3621);
or U5876 (N_5876,N_2751,N_3690);
and U5877 (N_5877,N_4058,N_2584);
nand U5878 (N_5878,N_2882,N_2757);
or U5879 (N_5879,N_3162,N_3176);
nor U5880 (N_5880,N_3698,N_2678);
nand U5881 (N_5881,N_4562,N_3517);
nor U5882 (N_5882,N_4351,N_4132);
and U5883 (N_5883,N_3225,N_4443);
and U5884 (N_5884,N_4285,N_3846);
nor U5885 (N_5885,N_3704,N_4676);
or U5886 (N_5886,N_4974,N_4678);
or U5887 (N_5887,N_2992,N_3650);
nor U5888 (N_5888,N_4690,N_4051);
and U5889 (N_5889,N_2514,N_3818);
nand U5890 (N_5890,N_2901,N_4056);
nand U5891 (N_5891,N_3958,N_4526);
or U5892 (N_5892,N_2894,N_3645);
or U5893 (N_5893,N_4467,N_4463);
nor U5894 (N_5894,N_4665,N_4036);
nor U5895 (N_5895,N_3170,N_2515);
nor U5896 (N_5896,N_3865,N_2738);
nand U5897 (N_5897,N_4829,N_4165);
nand U5898 (N_5898,N_3392,N_3095);
nand U5899 (N_5899,N_4421,N_3951);
and U5900 (N_5900,N_4820,N_4060);
and U5901 (N_5901,N_3783,N_4289);
nor U5902 (N_5902,N_3906,N_3943);
or U5903 (N_5903,N_2827,N_4833);
nand U5904 (N_5904,N_2593,N_4642);
nor U5905 (N_5905,N_3600,N_2513);
nand U5906 (N_5906,N_3669,N_3903);
nor U5907 (N_5907,N_3647,N_4472);
nand U5908 (N_5908,N_3364,N_3605);
nand U5909 (N_5909,N_3271,N_3496);
and U5910 (N_5910,N_2775,N_4885);
or U5911 (N_5911,N_4328,N_3227);
and U5912 (N_5912,N_3540,N_4648);
or U5913 (N_5913,N_4965,N_3457);
nor U5914 (N_5914,N_2519,N_4088);
or U5915 (N_5915,N_4333,N_3919);
and U5916 (N_5916,N_4214,N_3473);
or U5917 (N_5917,N_3644,N_4739);
nor U5918 (N_5918,N_2891,N_3174);
nor U5919 (N_5919,N_3316,N_4371);
nand U5920 (N_5920,N_3899,N_2794);
nor U5921 (N_5921,N_2560,N_3893);
nor U5922 (N_5922,N_2821,N_4346);
and U5923 (N_5923,N_3908,N_3113);
and U5924 (N_5924,N_3129,N_3767);
and U5925 (N_5925,N_3807,N_2897);
or U5926 (N_5926,N_3395,N_4475);
nand U5927 (N_5927,N_4778,N_3592);
nand U5928 (N_5928,N_4492,N_4981);
nand U5929 (N_5929,N_2830,N_3789);
nand U5930 (N_5930,N_4927,N_4809);
nand U5931 (N_5931,N_2746,N_3373);
or U5932 (N_5932,N_3562,N_4777);
nand U5933 (N_5933,N_2826,N_2887);
and U5934 (N_5934,N_3836,N_4348);
nand U5935 (N_5935,N_4938,N_4745);
and U5936 (N_5936,N_4753,N_3049);
or U5937 (N_5937,N_4426,N_2517);
nand U5938 (N_5938,N_3184,N_2630);
xor U5939 (N_5939,N_4511,N_3005);
or U5940 (N_5940,N_3241,N_4413);
and U5941 (N_5941,N_3253,N_3159);
nand U5942 (N_5942,N_3483,N_4957);
or U5943 (N_5943,N_3465,N_4245);
nor U5944 (N_5944,N_2981,N_2631);
nand U5945 (N_5945,N_4352,N_4243);
nor U5946 (N_5946,N_3801,N_2648);
and U5947 (N_5947,N_2664,N_4211);
nor U5948 (N_5948,N_3560,N_4083);
and U5949 (N_5949,N_3153,N_4514);
and U5950 (N_5950,N_2939,N_2657);
or U5951 (N_5951,N_3622,N_3624);
or U5952 (N_5952,N_3315,N_4023);
and U5953 (N_5953,N_2995,N_4063);
and U5954 (N_5954,N_3402,N_4887);
nand U5955 (N_5955,N_3020,N_3856);
nand U5956 (N_5956,N_3445,N_4922);
nor U5957 (N_5957,N_4892,N_4643);
or U5958 (N_5958,N_2580,N_4911);
nor U5959 (N_5959,N_3208,N_3400);
and U5960 (N_5960,N_3055,N_4537);
and U5961 (N_5961,N_3038,N_4868);
nor U5962 (N_5962,N_3664,N_3307);
or U5963 (N_5963,N_2923,N_4054);
nand U5964 (N_5964,N_3031,N_3578);
nor U5965 (N_5965,N_4768,N_4392);
or U5966 (N_5966,N_4367,N_4984);
nand U5967 (N_5967,N_4500,N_4749);
or U5968 (N_5968,N_4482,N_4169);
and U5969 (N_5969,N_2629,N_4263);
and U5970 (N_5970,N_2846,N_2944);
or U5971 (N_5971,N_3383,N_4264);
and U5972 (N_5972,N_3706,N_2558);
nor U5973 (N_5973,N_4506,N_2561);
and U5974 (N_5974,N_2615,N_4340);
and U5975 (N_5975,N_3324,N_4681);
and U5976 (N_5976,N_4425,N_4750);
nor U5977 (N_5977,N_4067,N_3180);
nor U5978 (N_5978,N_4554,N_3233);
and U5979 (N_5979,N_2907,N_2644);
xnor U5980 (N_5980,N_3336,N_4296);
or U5981 (N_5981,N_3959,N_3873);
nor U5982 (N_5982,N_2892,N_3399);
nand U5983 (N_5983,N_4731,N_3267);
or U5984 (N_5984,N_3046,N_4407);
or U5985 (N_5985,N_2501,N_3189);
nor U5986 (N_5986,N_3201,N_3337);
and U5987 (N_5987,N_3837,N_3568);
and U5988 (N_5988,N_4127,N_4076);
nand U5989 (N_5989,N_4219,N_2614);
or U5990 (N_5990,N_2508,N_4541);
nor U5991 (N_5991,N_2783,N_4553);
or U5992 (N_5992,N_2956,N_4983);
nand U5993 (N_5993,N_4969,N_3179);
and U5994 (N_5994,N_4430,N_3033);
nand U5995 (N_5995,N_4097,N_4569);
and U5996 (N_5996,N_3484,N_2539);
nand U5997 (N_5997,N_2591,N_4470);
and U5998 (N_5998,N_3469,N_3535);
nand U5999 (N_5999,N_2798,N_3454);
nand U6000 (N_6000,N_2735,N_2947);
or U6001 (N_6001,N_2970,N_3047);
and U6002 (N_6002,N_4356,N_4223);
nand U6003 (N_6003,N_4593,N_4141);
and U6004 (N_6004,N_4683,N_2790);
nand U6005 (N_6005,N_3000,N_4423);
nand U6006 (N_6006,N_3891,N_3279);
nand U6007 (N_6007,N_4098,N_4866);
nor U6008 (N_6008,N_4934,N_3637);
or U6009 (N_6009,N_3569,N_4142);
nand U6010 (N_6010,N_2597,N_4014);
and U6011 (N_6011,N_2544,N_4388);
nand U6012 (N_6012,N_4259,N_3806);
nor U6013 (N_6013,N_3023,N_4113);
or U6014 (N_6014,N_4235,N_2541);
and U6015 (N_6015,N_3702,N_3898);
and U6016 (N_6016,N_4669,N_2551);
and U6017 (N_6017,N_4722,N_3850);
nand U6018 (N_6018,N_2574,N_4302);
or U6019 (N_6019,N_4546,N_3530);
nor U6020 (N_6020,N_3526,N_4607);
nand U6021 (N_6021,N_3087,N_4798);
nor U6022 (N_6022,N_4190,N_4599);
and U6023 (N_6023,N_2857,N_3032);
or U6024 (N_6024,N_3790,N_3626);
nor U6025 (N_6025,N_4862,N_2702);
or U6026 (N_6026,N_3627,N_4521);
nand U6027 (N_6027,N_3720,N_4027);
and U6028 (N_6028,N_4530,N_3175);
nand U6029 (N_6029,N_3683,N_3760);
and U6030 (N_6030,N_3230,N_4273);
and U6031 (N_6031,N_4508,N_4622);
nand U6032 (N_6032,N_4061,N_3862);
and U6033 (N_6033,N_2750,N_4458);
nand U6034 (N_6034,N_3188,N_3960);
and U6035 (N_6035,N_3320,N_2908);
or U6036 (N_6036,N_3875,N_3932);
xnor U6037 (N_6037,N_4323,N_3981);
and U6038 (N_6038,N_2555,N_3685);
nor U6039 (N_6039,N_3511,N_4735);
nand U6040 (N_6040,N_2598,N_2899);
nor U6041 (N_6041,N_3443,N_2864);
and U6042 (N_6042,N_4770,N_4256);
or U6043 (N_6043,N_3553,N_3838);
nor U6044 (N_6044,N_3243,N_2958);
and U6045 (N_6045,N_3533,N_3620);
nor U6046 (N_6046,N_3220,N_4620);
or U6047 (N_6047,N_3742,N_3946);
nor U6048 (N_6048,N_3493,N_3472);
and U6049 (N_6049,N_3670,N_4359);
nor U6050 (N_6050,N_2835,N_3733);
nor U6051 (N_6051,N_2736,N_2833);
or U6052 (N_6052,N_3918,N_3438);
and U6053 (N_6053,N_2920,N_3531);
and U6054 (N_6054,N_3897,N_4369);
nor U6055 (N_6055,N_2766,N_4755);
nand U6056 (N_6056,N_3058,N_4213);
nor U6057 (N_6057,N_4631,N_2753);
and U6058 (N_6058,N_3098,N_2875);
nor U6059 (N_6059,N_3976,N_3709);
nor U6060 (N_6060,N_2605,N_4608);
nand U6061 (N_6061,N_2616,N_4284);
nand U6062 (N_6062,N_3264,N_4006);
or U6063 (N_6063,N_4292,N_4468);
nand U6064 (N_6064,N_4606,N_3552);
or U6065 (N_6065,N_3195,N_4865);
or U6066 (N_6066,N_3298,N_3766);
and U6067 (N_6067,N_4995,N_4330);
or U6068 (N_6068,N_3185,N_4168);
nor U6069 (N_6069,N_3274,N_2744);
or U6070 (N_6070,N_3040,N_4196);
and U6071 (N_6071,N_2807,N_3696);
and U6072 (N_6072,N_4786,N_4613);
and U6073 (N_6073,N_4650,N_4184);
nand U6074 (N_6074,N_3124,N_2579);
and U6075 (N_6075,N_4963,N_3612);
and U6076 (N_6076,N_3057,N_3390);
nand U6077 (N_6077,N_3823,N_3752);
and U6078 (N_6078,N_3222,N_3596);
nand U6079 (N_6079,N_2918,N_4533);
or U6080 (N_6080,N_2848,N_4331);
or U6081 (N_6081,N_4994,N_3589);
nand U6082 (N_6082,N_4216,N_4814);
or U6083 (N_6083,N_4070,N_2731);
or U6084 (N_6084,N_4917,N_3633);
nand U6085 (N_6085,N_4605,N_3198);
and U6086 (N_6086,N_3415,N_3680);
or U6087 (N_6087,N_3004,N_3203);
nor U6088 (N_6088,N_2984,N_2877);
nor U6089 (N_6089,N_4637,N_3112);
nor U6090 (N_6090,N_2990,N_3705);
or U6091 (N_6091,N_3729,N_3265);
nand U6092 (N_6092,N_2913,N_2537);
nor U6093 (N_6093,N_2692,N_3777);
or U6094 (N_6094,N_3972,N_4275);
or U6095 (N_6095,N_4758,N_3261);
nand U6096 (N_6096,N_3293,N_4019);
nor U6097 (N_6097,N_3656,N_2556);
nand U6098 (N_6098,N_4970,N_2662);
nand U6099 (N_6099,N_4041,N_3974);
nand U6100 (N_6100,N_4030,N_3464);
nor U6101 (N_6101,N_2910,N_4043);
and U6102 (N_6102,N_3755,N_3073);
and U6103 (N_6103,N_4815,N_3440);
and U6104 (N_6104,N_3367,N_3097);
xor U6105 (N_6105,N_4134,N_4743);
and U6106 (N_6106,N_3558,N_3289);
nand U6107 (N_6107,N_3114,N_4790);
or U6108 (N_6108,N_4386,N_2869);
and U6109 (N_6109,N_2786,N_4589);
or U6110 (N_6110,N_4912,N_4288);
nand U6111 (N_6111,N_4998,N_3871);
nor U6112 (N_6112,N_2876,N_3887);
nor U6113 (N_6113,N_4634,N_3093);
nor U6114 (N_6114,N_3730,N_4948);
and U6115 (N_6115,N_2716,N_2634);
and U6116 (N_6116,N_4985,N_4300);
nand U6117 (N_6117,N_3379,N_2747);
nor U6118 (N_6118,N_3432,N_3739);
nand U6119 (N_6119,N_3831,N_2714);
or U6120 (N_6120,N_3854,N_2935);
or U6121 (N_6121,N_3308,N_3125);
and U6122 (N_6122,N_2774,N_4174);
nand U6123 (N_6123,N_4657,N_2951);
nand U6124 (N_6124,N_4082,N_4972);
or U6125 (N_6125,N_4764,N_2845);
nor U6126 (N_6126,N_3662,N_3347);
or U6127 (N_6127,N_4926,N_3244);
nor U6128 (N_6128,N_4105,N_3813);
nand U6129 (N_6129,N_3771,N_3167);
xnor U6130 (N_6130,N_4697,N_3555);
nor U6131 (N_6131,N_3090,N_4221);
or U6132 (N_6132,N_4752,N_2868);
and U6133 (N_6133,N_4529,N_4639);
or U6134 (N_6134,N_2961,N_3628);
and U6135 (N_6135,N_2688,N_3607);
nand U6136 (N_6136,N_3677,N_2967);
nand U6137 (N_6137,N_2771,N_3407);
and U6138 (N_6138,N_2873,N_3019);
nor U6139 (N_6139,N_4751,N_4419);
nor U6140 (N_6140,N_3300,N_2748);
or U6141 (N_6141,N_4279,N_3349);
or U6142 (N_6142,N_4793,N_3059);
nor U6143 (N_6143,N_4402,N_3737);
and U6144 (N_6144,N_3476,N_4811);
and U6145 (N_6145,N_2975,N_4894);
nand U6146 (N_6146,N_4788,N_4543);
nor U6147 (N_6147,N_3635,N_4578);
or U6148 (N_6148,N_2516,N_3537);
nor U6149 (N_6149,N_3736,N_4307);
nor U6150 (N_6150,N_4694,N_3743);
and U6151 (N_6151,N_4343,N_2677);
nand U6152 (N_6152,N_4226,N_3333);
nor U6153 (N_6153,N_4379,N_4644);
nor U6154 (N_6154,N_4757,N_3213);
and U6155 (N_6155,N_2963,N_2853);
nand U6156 (N_6156,N_3181,N_3954);
nor U6157 (N_6157,N_3214,N_4194);
or U6158 (N_6158,N_4490,N_2553);
or U6159 (N_6159,N_4705,N_2504);
and U6160 (N_6160,N_3731,N_2533);
and U6161 (N_6161,N_4655,N_3219);
nor U6162 (N_6162,N_3211,N_3964);
nand U6163 (N_6163,N_4826,N_2779);
nor U6164 (N_6164,N_3975,N_2668);
nand U6165 (N_6165,N_2895,N_2511);
nor U6166 (N_6166,N_3872,N_2728);
nand U6167 (N_6167,N_4591,N_4918);
or U6168 (N_6168,N_4143,N_2824);
or U6169 (N_6169,N_4949,N_3681);
nand U6170 (N_6170,N_4409,N_3043);
nor U6171 (N_6171,N_3844,N_3351);
nor U6172 (N_6172,N_3642,N_3868);
nand U6173 (N_6173,N_3314,N_2718);
nand U6174 (N_6174,N_4195,N_4366);
nand U6175 (N_6175,N_4436,N_3118);
nand U6176 (N_6176,N_3917,N_4962);
or U6177 (N_6177,N_3360,N_4037);
or U6178 (N_6178,N_2921,N_3158);
and U6179 (N_6179,N_3732,N_4310);
and U6180 (N_6180,N_2861,N_4326);
or U6181 (N_6181,N_3199,N_3013);
nor U6182 (N_6182,N_2927,N_3148);
nor U6183 (N_6183,N_3575,N_3126);
or U6184 (N_6184,N_4089,N_4438);
nand U6185 (N_6185,N_3770,N_3840);
nor U6186 (N_6186,N_4480,N_4163);
nor U6187 (N_6187,N_4679,N_3433);
nor U6188 (N_6188,N_3757,N_3332);
and U6189 (N_6189,N_3962,N_3311);
nor U6190 (N_6190,N_3034,N_4077);
nor U6191 (N_6191,N_4740,N_2535);
nor U6192 (N_6192,N_3403,N_3226);
nand U6193 (N_6193,N_2781,N_2734);
and U6194 (N_6194,N_3431,N_3686);
nor U6195 (N_6195,N_4398,N_3221);
nor U6196 (N_6196,N_4747,N_4807);
and U6197 (N_6197,N_3024,N_3481);
nor U6198 (N_6198,N_4172,N_3010);
nor U6199 (N_6199,N_3795,N_3281);
or U6200 (N_6200,N_4192,N_4664);
nor U6201 (N_6201,N_2545,N_3413);
nor U6202 (N_6202,N_4662,N_4638);
and U6203 (N_6203,N_3722,N_4792);
and U6204 (N_6204,N_4594,N_2685);
nor U6205 (N_6205,N_4224,N_3728);
and U6206 (N_6206,N_2780,N_4298);
nor U6207 (N_6207,N_2761,N_3147);
nand U6208 (N_6208,N_3053,N_4978);
nand U6209 (N_6209,N_3160,N_3335);
nor U6210 (N_6210,N_3796,N_3063);
nand U6211 (N_6211,N_3166,N_4518);
nor U6212 (N_6212,N_3479,N_4394);
or U6213 (N_6213,N_3653,N_4204);
or U6214 (N_6214,N_4525,N_3275);
and U6215 (N_6215,N_2912,N_4175);
nor U6216 (N_6216,N_4145,N_2572);
and U6217 (N_6217,N_3151,N_4123);
and U6218 (N_6218,N_3971,N_2732);
and U6219 (N_6219,N_2658,N_2655);
and U6220 (N_6220,N_2547,N_4410);
and U6221 (N_6221,N_3638,N_3857);
nor U6222 (N_6222,N_4723,N_2530);
nor U6223 (N_6223,N_3996,N_3326);
nor U6224 (N_6224,N_4081,N_3591);
nor U6225 (N_6225,N_3192,N_3609);
nor U6226 (N_6226,N_4796,N_4440);
nand U6227 (N_6227,N_4532,N_3711);
or U6228 (N_6228,N_4967,N_4242);
or U6229 (N_6229,N_3994,N_3902);
or U6230 (N_6230,N_3874,N_4496);
or U6231 (N_6231,N_2694,N_4215);
or U6232 (N_6232,N_2902,N_3405);
and U6233 (N_6233,N_4652,N_4309);
nand U6234 (N_6234,N_4079,N_2505);
or U6235 (N_6235,N_4339,N_3785);
or U6236 (N_6236,N_4689,N_3471);
nand U6237 (N_6237,N_4627,N_2549);
nor U6238 (N_6238,N_3270,N_2671);
nor U6239 (N_6239,N_3793,N_3284);
nand U6240 (N_6240,N_4193,N_3132);
and U6241 (N_6241,N_2991,N_3260);
nand U6242 (N_6242,N_2624,N_3216);
or U6243 (N_6243,N_3921,N_3384);
and U6244 (N_6244,N_2528,N_3007);
nand U6245 (N_6245,N_2693,N_4602);
or U6246 (N_6246,N_4649,N_3051);
nor U6247 (N_6247,N_4280,N_4009);
xnor U6248 (N_6248,N_3086,N_4800);
and U6249 (N_6249,N_3835,N_4000);
nand U6250 (N_6250,N_3822,N_3708);
and U6251 (N_6251,N_4165,N_2881);
nor U6252 (N_6252,N_3228,N_4709);
and U6253 (N_6253,N_3470,N_4531);
or U6254 (N_6254,N_4889,N_2835);
and U6255 (N_6255,N_3917,N_3889);
or U6256 (N_6256,N_2857,N_3112);
and U6257 (N_6257,N_3184,N_4966);
and U6258 (N_6258,N_4583,N_3628);
and U6259 (N_6259,N_3588,N_4895);
and U6260 (N_6260,N_3223,N_3554);
or U6261 (N_6261,N_4092,N_4053);
nand U6262 (N_6262,N_2568,N_4321);
nor U6263 (N_6263,N_3507,N_3742);
nor U6264 (N_6264,N_2784,N_2985);
nor U6265 (N_6265,N_3970,N_2698);
or U6266 (N_6266,N_3140,N_4448);
nand U6267 (N_6267,N_2641,N_2954);
nand U6268 (N_6268,N_3625,N_4073);
or U6269 (N_6269,N_2617,N_3889);
and U6270 (N_6270,N_3272,N_2686);
and U6271 (N_6271,N_3769,N_2536);
or U6272 (N_6272,N_4364,N_3238);
nor U6273 (N_6273,N_4519,N_4523);
nand U6274 (N_6274,N_3869,N_4170);
nand U6275 (N_6275,N_3526,N_4084);
and U6276 (N_6276,N_3908,N_4765);
xnor U6277 (N_6277,N_2752,N_3756);
nor U6278 (N_6278,N_3155,N_3099);
or U6279 (N_6279,N_3595,N_2794);
and U6280 (N_6280,N_3906,N_3701);
or U6281 (N_6281,N_4165,N_2939);
nand U6282 (N_6282,N_4664,N_2869);
or U6283 (N_6283,N_2662,N_4299);
nand U6284 (N_6284,N_3425,N_4245);
or U6285 (N_6285,N_3865,N_3076);
or U6286 (N_6286,N_3419,N_3299);
or U6287 (N_6287,N_3313,N_4302);
and U6288 (N_6288,N_3329,N_4344);
or U6289 (N_6289,N_4458,N_3215);
or U6290 (N_6290,N_3853,N_2650);
nand U6291 (N_6291,N_3475,N_3423);
nand U6292 (N_6292,N_3596,N_3738);
nand U6293 (N_6293,N_3129,N_4796);
and U6294 (N_6294,N_4931,N_4897);
and U6295 (N_6295,N_4395,N_3119);
or U6296 (N_6296,N_3039,N_4703);
and U6297 (N_6297,N_3267,N_4456);
nand U6298 (N_6298,N_3590,N_3121);
or U6299 (N_6299,N_2816,N_4475);
nand U6300 (N_6300,N_3601,N_3134);
nor U6301 (N_6301,N_3188,N_3795);
nand U6302 (N_6302,N_3577,N_4938);
nor U6303 (N_6303,N_3082,N_4670);
nor U6304 (N_6304,N_4979,N_4926);
nand U6305 (N_6305,N_3166,N_2885);
nor U6306 (N_6306,N_3764,N_4759);
and U6307 (N_6307,N_3929,N_2924);
or U6308 (N_6308,N_4029,N_4052);
nand U6309 (N_6309,N_3289,N_4054);
nand U6310 (N_6310,N_4963,N_3258);
nand U6311 (N_6311,N_2566,N_3795);
nor U6312 (N_6312,N_4280,N_4252);
and U6313 (N_6313,N_3499,N_3908);
nand U6314 (N_6314,N_3312,N_3136);
nand U6315 (N_6315,N_3208,N_4204);
and U6316 (N_6316,N_4233,N_2921);
or U6317 (N_6317,N_4239,N_4932);
or U6318 (N_6318,N_4567,N_3911);
and U6319 (N_6319,N_4560,N_4330);
nand U6320 (N_6320,N_3947,N_4112);
and U6321 (N_6321,N_4830,N_4228);
or U6322 (N_6322,N_4577,N_4741);
and U6323 (N_6323,N_3628,N_4363);
and U6324 (N_6324,N_2514,N_4404);
nor U6325 (N_6325,N_4076,N_3349);
nand U6326 (N_6326,N_4277,N_3479);
and U6327 (N_6327,N_2544,N_2877);
nand U6328 (N_6328,N_4810,N_2876);
nand U6329 (N_6329,N_3143,N_4330);
nand U6330 (N_6330,N_4683,N_4095);
or U6331 (N_6331,N_3551,N_3717);
nand U6332 (N_6332,N_3838,N_4572);
nor U6333 (N_6333,N_2861,N_3002);
and U6334 (N_6334,N_2900,N_4778);
nor U6335 (N_6335,N_3808,N_3732);
and U6336 (N_6336,N_2666,N_3908);
nor U6337 (N_6337,N_3976,N_4125);
nor U6338 (N_6338,N_3462,N_4619);
nor U6339 (N_6339,N_4567,N_2526);
or U6340 (N_6340,N_3584,N_4262);
nor U6341 (N_6341,N_3001,N_3294);
and U6342 (N_6342,N_2887,N_4779);
nor U6343 (N_6343,N_3974,N_4329);
nor U6344 (N_6344,N_3500,N_2937);
and U6345 (N_6345,N_3734,N_3179);
and U6346 (N_6346,N_4755,N_2800);
and U6347 (N_6347,N_2564,N_3685);
or U6348 (N_6348,N_2539,N_4730);
nor U6349 (N_6349,N_3624,N_3636);
and U6350 (N_6350,N_4292,N_3428);
nand U6351 (N_6351,N_3328,N_4962);
and U6352 (N_6352,N_3861,N_3722);
and U6353 (N_6353,N_3973,N_4047);
and U6354 (N_6354,N_3589,N_4965);
nand U6355 (N_6355,N_3332,N_2792);
nor U6356 (N_6356,N_4330,N_3834);
nor U6357 (N_6357,N_3093,N_4373);
and U6358 (N_6358,N_4257,N_3384);
nor U6359 (N_6359,N_4948,N_2912);
nand U6360 (N_6360,N_2904,N_3862);
and U6361 (N_6361,N_3691,N_4083);
nor U6362 (N_6362,N_4917,N_4799);
or U6363 (N_6363,N_4502,N_3477);
and U6364 (N_6364,N_3812,N_4607);
or U6365 (N_6365,N_4667,N_4029);
nand U6366 (N_6366,N_3319,N_2844);
nand U6367 (N_6367,N_4004,N_3676);
nor U6368 (N_6368,N_4637,N_3705);
or U6369 (N_6369,N_2560,N_3538);
and U6370 (N_6370,N_4439,N_3354);
xor U6371 (N_6371,N_4065,N_4704);
and U6372 (N_6372,N_2650,N_3798);
nor U6373 (N_6373,N_4241,N_3427);
and U6374 (N_6374,N_4860,N_4000);
or U6375 (N_6375,N_2886,N_2973);
or U6376 (N_6376,N_2604,N_4545);
and U6377 (N_6377,N_3779,N_3014);
or U6378 (N_6378,N_3773,N_2701);
and U6379 (N_6379,N_4598,N_2988);
nor U6380 (N_6380,N_3006,N_4681);
and U6381 (N_6381,N_4010,N_3858);
or U6382 (N_6382,N_4595,N_4389);
nor U6383 (N_6383,N_3703,N_4708);
nand U6384 (N_6384,N_3954,N_4031);
or U6385 (N_6385,N_2901,N_3367);
or U6386 (N_6386,N_3178,N_4578);
nor U6387 (N_6387,N_4705,N_4915);
nand U6388 (N_6388,N_2751,N_4734);
and U6389 (N_6389,N_3144,N_4700);
and U6390 (N_6390,N_3339,N_3547);
or U6391 (N_6391,N_2754,N_3165);
or U6392 (N_6392,N_4066,N_4031);
nor U6393 (N_6393,N_3623,N_2889);
nor U6394 (N_6394,N_3450,N_4041);
nand U6395 (N_6395,N_4293,N_4046);
nand U6396 (N_6396,N_2597,N_4517);
or U6397 (N_6397,N_4430,N_4441);
xnor U6398 (N_6398,N_4321,N_3924);
and U6399 (N_6399,N_4752,N_3127);
nand U6400 (N_6400,N_2687,N_3482);
or U6401 (N_6401,N_4799,N_3737);
or U6402 (N_6402,N_2812,N_4206);
and U6403 (N_6403,N_2789,N_3095);
and U6404 (N_6404,N_4000,N_3857);
or U6405 (N_6405,N_3038,N_3206);
nor U6406 (N_6406,N_4556,N_4535);
nand U6407 (N_6407,N_3929,N_3082);
nor U6408 (N_6408,N_4103,N_2816);
or U6409 (N_6409,N_4298,N_3508);
nand U6410 (N_6410,N_4609,N_2714);
nor U6411 (N_6411,N_2812,N_4009);
and U6412 (N_6412,N_4291,N_2939);
nand U6413 (N_6413,N_4104,N_4694);
and U6414 (N_6414,N_2592,N_3094);
nor U6415 (N_6415,N_2583,N_4304);
nor U6416 (N_6416,N_4183,N_3338);
or U6417 (N_6417,N_4409,N_2540);
and U6418 (N_6418,N_3641,N_3744);
nor U6419 (N_6419,N_2662,N_2799);
nor U6420 (N_6420,N_2651,N_4292);
nand U6421 (N_6421,N_2991,N_4712);
nand U6422 (N_6422,N_4532,N_4064);
and U6423 (N_6423,N_4030,N_2920);
nand U6424 (N_6424,N_4322,N_4187);
nor U6425 (N_6425,N_2909,N_3819);
nor U6426 (N_6426,N_2880,N_2529);
nand U6427 (N_6427,N_4361,N_2846);
nand U6428 (N_6428,N_3140,N_3079);
nand U6429 (N_6429,N_3396,N_3111);
nand U6430 (N_6430,N_3608,N_3732);
nor U6431 (N_6431,N_3976,N_3605);
nor U6432 (N_6432,N_4193,N_2641);
and U6433 (N_6433,N_3760,N_3910);
nor U6434 (N_6434,N_4954,N_3923);
and U6435 (N_6435,N_2557,N_4493);
and U6436 (N_6436,N_3976,N_3639);
or U6437 (N_6437,N_4050,N_3337);
nand U6438 (N_6438,N_2503,N_2760);
nor U6439 (N_6439,N_4735,N_3560);
or U6440 (N_6440,N_4183,N_2572);
or U6441 (N_6441,N_3447,N_3380);
nand U6442 (N_6442,N_2908,N_3335);
nor U6443 (N_6443,N_3463,N_4809);
or U6444 (N_6444,N_3328,N_3543);
nor U6445 (N_6445,N_4184,N_3114);
and U6446 (N_6446,N_3916,N_2739);
or U6447 (N_6447,N_3733,N_4696);
nand U6448 (N_6448,N_4780,N_3628);
or U6449 (N_6449,N_3998,N_3245);
nand U6450 (N_6450,N_3411,N_3122);
and U6451 (N_6451,N_3448,N_4721);
nand U6452 (N_6452,N_4387,N_3471);
or U6453 (N_6453,N_2731,N_4663);
nor U6454 (N_6454,N_4507,N_2883);
and U6455 (N_6455,N_4146,N_3458);
or U6456 (N_6456,N_4100,N_3820);
nand U6457 (N_6457,N_2639,N_2771);
nand U6458 (N_6458,N_3560,N_2625);
nand U6459 (N_6459,N_2704,N_4995);
nand U6460 (N_6460,N_3458,N_4310);
or U6461 (N_6461,N_4823,N_3868);
and U6462 (N_6462,N_2855,N_4703);
nand U6463 (N_6463,N_2674,N_4976);
and U6464 (N_6464,N_4519,N_4484);
nand U6465 (N_6465,N_3535,N_2627);
or U6466 (N_6466,N_4050,N_3025);
nand U6467 (N_6467,N_4850,N_3521);
and U6468 (N_6468,N_4787,N_4710);
nor U6469 (N_6469,N_3010,N_4203);
nor U6470 (N_6470,N_3206,N_2563);
and U6471 (N_6471,N_4009,N_2594);
or U6472 (N_6472,N_3482,N_2765);
or U6473 (N_6473,N_2798,N_2508);
or U6474 (N_6474,N_3791,N_3519);
nand U6475 (N_6475,N_4193,N_4124);
or U6476 (N_6476,N_3938,N_4335);
nor U6477 (N_6477,N_3872,N_4956);
and U6478 (N_6478,N_4500,N_4109);
nand U6479 (N_6479,N_2592,N_4658);
or U6480 (N_6480,N_4267,N_3341);
nor U6481 (N_6481,N_2581,N_2817);
and U6482 (N_6482,N_3323,N_4659);
nand U6483 (N_6483,N_3645,N_4584);
and U6484 (N_6484,N_3755,N_3946);
or U6485 (N_6485,N_4730,N_4995);
or U6486 (N_6486,N_4740,N_4508);
nand U6487 (N_6487,N_2797,N_4879);
or U6488 (N_6488,N_2942,N_3231);
and U6489 (N_6489,N_4223,N_2800);
and U6490 (N_6490,N_2666,N_4999);
and U6491 (N_6491,N_4581,N_2653);
and U6492 (N_6492,N_4500,N_4183);
nor U6493 (N_6493,N_4633,N_4918);
nor U6494 (N_6494,N_3144,N_2852);
or U6495 (N_6495,N_4329,N_4628);
nand U6496 (N_6496,N_3428,N_3679);
and U6497 (N_6497,N_4420,N_4341);
nand U6498 (N_6498,N_2592,N_3968);
nor U6499 (N_6499,N_3194,N_3420);
nor U6500 (N_6500,N_2506,N_2826);
nand U6501 (N_6501,N_2593,N_2935);
and U6502 (N_6502,N_3882,N_2533);
nand U6503 (N_6503,N_3818,N_3789);
or U6504 (N_6504,N_4368,N_4614);
and U6505 (N_6505,N_4888,N_4214);
and U6506 (N_6506,N_4385,N_4442);
nor U6507 (N_6507,N_4135,N_4372);
nand U6508 (N_6508,N_4492,N_2732);
and U6509 (N_6509,N_4966,N_3120);
nand U6510 (N_6510,N_3616,N_2971);
nor U6511 (N_6511,N_3897,N_3755);
and U6512 (N_6512,N_3275,N_2622);
nand U6513 (N_6513,N_3784,N_3046);
nand U6514 (N_6514,N_2988,N_4877);
nand U6515 (N_6515,N_3751,N_2745);
nor U6516 (N_6516,N_3576,N_4488);
nand U6517 (N_6517,N_3322,N_4002);
nand U6518 (N_6518,N_2941,N_3125);
or U6519 (N_6519,N_3150,N_3068);
and U6520 (N_6520,N_4960,N_3504);
nand U6521 (N_6521,N_4610,N_4000);
nand U6522 (N_6522,N_4589,N_3313);
nor U6523 (N_6523,N_3831,N_2720);
nor U6524 (N_6524,N_2961,N_4416);
nor U6525 (N_6525,N_4816,N_2906);
and U6526 (N_6526,N_4093,N_4769);
and U6527 (N_6527,N_3514,N_3159);
and U6528 (N_6528,N_3748,N_4008);
or U6529 (N_6529,N_3672,N_3970);
and U6530 (N_6530,N_4394,N_2863);
nor U6531 (N_6531,N_3479,N_3267);
nor U6532 (N_6532,N_4531,N_3498);
or U6533 (N_6533,N_3591,N_3010);
or U6534 (N_6534,N_4897,N_3626);
or U6535 (N_6535,N_2913,N_3060);
or U6536 (N_6536,N_4384,N_2750);
nand U6537 (N_6537,N_2517,N_4411);
nor U6538 (N_6538,N_3696,N_3155);
nand U6539 (N_6539,N_2569,N_4945);
and U6540 (N_6540,N_4825,N_3962);
or U6541 (N_6541,N_4482,N_3043);
or U6542 (N_6542,N_3896,N_4548);
or U6543 (N_6543,N_3820,N_2734);
and U6544 (N_6544,N_3785,N_3624);
and U6545 (N_6545,N_4459,N_4611);
nand U6546 (N_6546,N_3969,N_4810);
or U6547 (N_6547,N_3395,N_3607);
nand U6548 (N_6548,N_3979,N_3165);
and U6549 (N_6549,N_2931,N_3340);
nor U6550 (N_6550,N_3165,N_3331);
and U6551 (N_6551,N_4358,N_3353);
and U6552 (N_6552,N_3743,N_4536);
nor U6553 (N_6553,N_4494,N_3986);
or U6554 (N_6554,N_2503,N_3913);
nor U6555 (N_6555,N_4994,N_4977);
nand U6556 (N_6556,N_3849,N_4791);
nor U6557 (N_6557,N_4655,N_3200);
and U6558 (N_6558,N_2507,N_3294);
and U6559 (N_6559,N_3823,N_3149);
nor U6560 (N_6560,N_3847,N_3851);
and U6561 (N_6561,N_4917,N_3250);
nand U6562 (N_6562,N_4163,N_4872);
or U6563 (N_6563,N_4746,N_3245);
nor U6564 (N_6564,N_3743,N_2695);
nor U6565 (N_6565,N_3446,N_4930);
or U6566 (N_6566,N_3406,N_4271);
nor U6567 (N_6567,N_3723,N_3657);
and U6568 (N_6568,N_3771,N_3839);
and U6569 (N_6569,N_4516,N_2550);
nor U6570 (N_6570,N_4857,N_4304);
and U6571 (N_6571,N_3765,N_3107);
or U6572 (N_6572,N_3628,N_2537);
nor U6573 (N_6573,N_3466,N_2815);
or U6574 (N_6574,N_4494,N_4449);
nor U6575 (N_6575,N_4779,N_4626);
nor U6576 (N_6576,N_3822,N_4948);
or U6577 (N_6577,N_4636,N_4380);
or U6578 (N_6578,N_2530,N_4935);
nor U6579 (N_6579,N_3621,N_3839);
nor U6580 (N_6580,N_4401,N_3260);
nand U6581 (N_6581,N_3149,N_2654);
or U6582 (N_6582,N_3839,N_3241);
and U6583 (N_6583,N_2766,N_3943);
nor U6584 (N_6584,N_3839,N_2781);
or U6585 (N_6585,N_3088,N_2928);
and U6586 (N_6586,N_2751,N_4513);
or U6587 (N_6587,N_3691,N_3181);
nor U6588 (N_6588,N_4996,N_4049);
and U6589 (N_6589,N_2894,N_4241);
nand U6590 (N_6590,N_3762,N_4007);
and U6591 (N_6591,N_3015,N_4584);
or U6592 (N_6592,N_4696,N_2503);
nand U6593 (N_6593,N_3794,N_3438);
and U6594 (N_6594,N_4932,N_3388);
or U6595 (N_6595,N_3467,N_4149);
nor U6596 (N_6596,N_4948,N_4234);
or U6597 (N_6597,N_4981,N_4176);
or U6598 (N_6598,N_2959,N_3637);
nand U6599 (N_6599,N_3684,N_2656);
and U6600 (N_6600,N_4075,N_2926);
nor U6601 (N_6601,N_2698,N_3274);
or U6602 (N_6602,N_4011,N_4423);
nand U6603 (N_6603,N_4508,N_4244);
and U6604 (N_6604,N_3383,N_4636);
nor U6605 (N_6605,N_2893,N_4839);
or U6606 (N_6606,N_3008,N_2677);
xor U6607 (N_6607,N_3774,N_4982);
and U6608 (N_6608,N_3445,N_3118);
and U6609 (N_6609,N_4748,N_4685);
or U6610 (N_6610,N_2984,N_3085);
and U6611 (N_6611,N_4478,N_4486);
nor U6612 (N_6612,N_4900,N_4929);
nor U6613 (N_6613,N_3491,N_2842);
and U6614 (N_6614,N_4136,N_4574);
or U6615 (N_6615,N_3348,N_3818);
nand U6616 (N_6616,N_3596,N_3698);
nand U6617 (N_6617,N_3507,N_4788);
or U6618 (N_6618,N_3774,N_3354);
or U6619 (N_6619,N_4886,N_3783);
or U6620 (N_6620,N_4748,N_4539);
nand U6621 (N_6621,N_4342,N_3786);
or U6622 (N_6622,N_2644,N_3775);
and U6623 (N_6623,N_3648,N_4276);
nor U6624 (N_6624,N_3695,N_3539);
nor U6625 (N_6625,N_3934,N_2529);
or U6626 (N_6626,N_2912,N_3143);
nand U6627 (N_6627,N_3948,N_3188);
or U6628 (N_6628,N_2986,N_2838);
nor U6629 (N_6629,N_3264,N_4955);
or U6630 (N_6630,N_3157,N_4241);
or U6631 (N_6631,N_4623,N_3927);
and U6632 (N_6632,N_4616,N_2586);
nand U6633 (N_6633,N_4958,N_4283);
and U6634 (N_6634,N_2871,N_3794);
nor U6635 (N_6635,N_3177,N_3407);
and U6636 (N_6636,N_4921,N_4815);
xnor U6637 (N_6637,N_3530,N_3787);
or U6638 (N_6638,N_4196,N_3679);
and U6639 (N_6639,N_4032,N_2982);
or U6640 (N_6640,N_3559,N_4369);
or U6641 (N_6641,N_4034,N_3720);
nand U6642 (N_6642,N_4732,N_3409);
xor U6643 (N_6643,N_2819,N_3165);
nand U6644 (N_6644,N_3442,N_3934);
xor U6645 (N_6645,N_4069,N_4021);
or U6646 (N_6646,N_4059,N_2574);
or U6647 (N_6647,N_4396,N_2765);
nor U6648 (N_6648,N_2890,N_3964);
and U6649 (N_6649,N_2720,N_3194);
or U6650 (N_6650,N_3378,N_4432);
and U6651 (N_6651,N_2785,N_4563);
nor U6652 (N_6652,N_4969,N_3469);
nor U6653 (N_6653,N_3176,N_3270);
and U6654 (N_6654,N_4009,N_3868);
nor U6655 (N_6655,N_4718,N_2702);
nor U6656 (N_6656,N_3684,N_2621);
nand U6657 (N_6657,N_3271,N_2906);
nor U6658 (N_6658,N_4990,N_4963);
nand U6659 (N_6659,N_4189,N_3754);
or U6660 (N_6660,N_2541,N_3985);
and U6661 (N_6661,N_3719,N_4327);
and U6662 (N_6662,N_3811,N_4886);
or U6663 (N_6663,N_4415,N_3570);
nor U6664 (N_6664,N_4784,N_3501);
nand U6665 (N_6665,N_3985,N_3041);
nand U6666 (N_6666,N_4511,N_4566);
and U6667 (N_6667,N_3089,N_3984);
or U6668 (N_6668,N_4362,N_3871);
nand U6669 (N_6669,N_3154,N_4497);
nand U6670 (N_6670,N_4826,N_2891);
nand U6671 (N_6671,N_4889,N_3792);
or U6672 (N_6672,N_3165,N_4194);
nand U6673 (N_6673,N_2695,N_4558);
nand U6674 (N_6674,N_3374,N_4071);
or U6675 (N_6675,N_2889,N_2726);
nor U6676 (N_6676,N_4509,N_4268);
and U6677 (N_6677,N_4124,N_4243);
and U6678 (N_6678,N_3515,N_4400);
and U6679 (N_6679,N_4796,N_2509);
nand U6680 (N_6680,N_4597,N_3661);
or U6681 (N_6681,N_3110,N_3252);
or U6682 (N_6682,N_3403,N_2665);
nor U6683 (N_6683,N_4812,N_4234);
nor U6684 (N_6684,N_3530,N_3067);
nand U6685 (N_6685,N_4898,N_2590);
nor U6686 (N_6686,N_2529,N_3553);
nor U6687 (N_6687,N_4813,N_4715);
nand U6688 (N_6688,N_3520,N_2588);
nor U6689 (N_6689,N_4830,N_3592);
nand U6690 (N_6690,N_3970,N_4619);
nand U6691 (N_6691,N_2987,N_2909);
nand U6692 (N_6692,N_2884,N_2736);
and U6693 (N_6693,N_3146,N_3786);
nor U6694 (N_6694,N_3890,N_4580);
and U6695 (N_6695,N_2939,N_3489);
and U6696 (N_6696,N_3160,N_4700);
nand U6697 (N_6697,N_3546,N_4227);
or U6698 (N_6698,N_4258,N_3731);
or U6699 (N_6699,N_3766,N_3399);
and U6700 (N_6700,N_4030,N_2888);
or U6701 (N_6701,N_3353,N_3688);
nor U6702 (N_6702,N_4440,N_2725);
or U6703 (N_6703,N_4244,N_4122);
nand U6704 (N_6704,N_3980,N_3491);
and U6705 (N_6705,N_3844,N_4248);
or U6706 (N_6706,N_2696,N_3184);
nand U6707 (N_6707,N_3809,N_4459);
nand U6708 (N_6708,N_3372,N_4340);
nor U6709 (N_6709,N_3759,N_4074);
and U6710 (N_6710,N_3321,N_2707);
nor U6711 (N_6711,N_3985,N_4216);
nand U6712 (N_6712,N_3892,N_2620);
nor U6713 (N_6713,N_3904,N_4304);
or U6714 (N_6714,N_4175,N_3934);
nand U6715 (N_6715,N_4066,N_4630);
and U6716 (N_6716,N_4929,N_3627);
nor U6717 (N_6717,N_3323,N_3242);
nand U6718 (N_6718,N_3797,N_4015);
nand U6719 (N_6719,N_3776,N_4290);
or U6720 (N_6720,N_2798,N_4261);
nor U6721 (N_6721,N_4078,N_2529);
nor U6722 (N_6722,N_3514,N_4639);
or U6723 (N_6723,N_4042,N_2905);
and U6724 (N_6724,N_4970,N_3458);
nand U6725 (N_6725,N_3030,N_3562);
and U6726 (N_6726,N_4837,N_3166);
nor U6727 (N_6727,N_4427,N_4092);
or U6728 (N_6728,N_4541,N_4457);
nand U6729 (N_6729,N_3913,N_2530);
and U6730 (N_6730,N_3542,N_3278);
nor U6731 (N_6731,N_3465,N_3223);
and U6732 (N_6732,N_2630,N_3169);
nand U6733 (N_6733,N_3445,N_4300);
nand U6734 (N_6734,N_4746,N_2741);
nor U6735 (N_6735,N_3186,N_2883);
nor U6736 (N_6736,N_3486,N_2779);
nor U6737 (N_6737,N_4152,N_2526);
nand U6738 (N_6738,N_4563,N_4455);
nand U6739 (N_6739,N_4939,N_2639);
and U6740 (N_6740,N_3005,N_4419);
nand U6741 (N_6741,N_2847,N_4338);
nand U6742 (N_6742,N_3621,N_3026);
xor U6743 (N_6743,N_4230,N_3501);
and U6744 (N_6744,N_3721,N_2647);
and U6745 (N_6745,N_3416,N_4668);
nand U6746 (N_6746,N_4713,N_3072);
nor U6747 (N_6747,N_2808,N_4344);
and U6748 (N_6748,N_4078,N_2973);
and U6749 (N_6749,N_3365,N_4591);
or U6750 (N_6750,N_3478,N_4049);
nand U6751 (N_6751,N_3514,N_2657);
and U6752 (N_6752,N_4138,N_4946);
or U6753 (N_6753,N_3320,N_2552);
nor U6754 (N_6754,N_3807,N_2661);
and U6755 (N_6755,N_4521,N_4823);
nand U6756 (N_6756,N_4155,N_2543);
nor U6757 (N_6757,N_2857,N_3188);
nor U6758 (N_6758,N_3977,N_2565);
nor U6759 (N_6759,N_3199,N_3169);
nor U6760 (N_6760,N_3866,N_3176);
and U6761 (N_6761,N_3094,N_4465);
and U6762 (N_6762,N_2654,N_3468);
nand U6763 (N_6763,N_3590,N_4632);
nand U6764 (N_6764,N_3348,N_4081);
nand U6765 (N_6765,N_3296,N_2812);
or U6766 (N_6766,N_2712,N_4951);
or U6767 (N_6767,N_4079,N_3841);
or U6768 (N_6768,N_2635,N_4892);
and U6769 (N_6769,N_3178,N_3756);
and U6770 (N_6770,N_3204,N_4156);
nand U6771 (N_6771,N_3802,N_3492);
nor U6772 (N_6772,N_2768,N_4226);
nand U6773 (N_6773,N_4863,N_3003);
nand U6774 (N_6774,N_4528,N_4400);
or U6775 (N_6775,N_2770,N_4548);
nand U6776 (N_6776,N_2597,N_4667);
or U6777 (N_6777,N_4524,N_4700);
nor U6778 (N_6778,N_3188,N_4573);
or U6779 (N_6779,N_3090,N_4267);
or U6780 (N_6780,N_2930,N_3981);
nor U6781 (N_6781,N_4330,N_3496);
or U6782 (N_6782,N_3580,N_2817);
nor U6783 (N_6783,N_2924,N_3941);
nand U6784 (N_6784,N_4940,N_3502);
or U6785 (N_6785,N_2735,N_3984);
nor U6786 (N_6786,N_4206,N_4227);
nor U6787 (N_6787,N_3158,N_3676);
or U6788 (N_6788,N_4101,N_2727);
and U6789 (N_6789,N_2614,N_2793);
or U6790 (N_6790,N_2847,N_3371);
and U6791 (N_6791,N_2578,N_4703);
and U6792 (N_6792,N_4215,N_4602);
or U6793 (N_6793,N_3296,N_3395);
nor U6794 (N_6794,N_4497,N_3854);
nand U6795 (N_6795,N_4157,N_4368);
and U6796 (N_6796,N_4016,N_4175);
nor U6797 (N_6797,N_2726,N_4392);
nor U6798 (N_6798,N_4471,N_4118);
nor U6799 (N_6799,N_2507,N_3688);
nor U6800 (N_6800,N_4404,N_4417);
nor U6801 (N_6801,N_3132,N_3927);
nand U6802 (N_6802,N_3077,N_4945);
nor U6803 (N_6803,N_4621,N_4520);
nor U6804 (N_6804,N_2947,N_3623);
and U6805 (N_6805,N_4232,N_3114);
or U6806 (N_6806,N_3319,N_3939);
and U6807 (N_6807,N_3003,N_3515);
nand U6808 (N_6808,N_2752,N_3784);
nor U6809 (N_6809,N_2849,N_3491);
or U6810 (N_6810,N_4622,N_3070);
or U6811 (N_6811,N_4424,N_3658);
nor U6812 (N_6812,N_3361,N_4410);
nand U6813 (N_6813,N_3130,N_4594);
and U6814 (N_6814,N_4220,N_3388);
nor U6815 (N_6815,N_4054,N_2545);
nor U6816 (N_6816,N_3429,N_4767);
nor U6817 (N_6817,N_4538,N_4424);
nor U6818 (N_6818,N_4079,N_3116);
nor U6819 (N_6819,N_3134,N_4482);
or U6820 (N_6820,N_2650,N_2831);
nand U6821 (N_6821,N_3029,N_3226);
nand U6822 (N_6822,N_4255,N_3926);
or U6823 (N_6823,N_3936,N_4328);
nand U6824 (N_6824,N_3657,N_3540);
nor U6825 (N_6825,N_2574,N_2721);
or U6826 (N_6826,N_3166,N_4272);
and U6827 (N_6827,N_3058,N_3569);
nand U6828 (N_6828,N_3383,N_3096);
nor U6829 (N_6829,N_4064,N_4393);
or U6830 (N_6830,N_4992,N_3380);
and U6831 (N_6831,N_3245,N_3098);
nand U6832 (N_6832,N_2545,N_3985);
nor U6833 (N_6833,N_3850,N_3390);
or U6834 (N_6834,N_3447,N_3102);
or U6835 (N_6835,N_3710,N_3277);
nor U6836 (N_6836,N_4344,N_3750);
and U6837 (N_6837,N_4824,N_3855);
nand U6838 (N_6838,N_3793,N_3307);
or U6839 (N_6839,N_4502,N_3076);
and U6840 (N_6840,N_3895,N_3460);
and U6841 (N_6841,N_4210,N_3851);
nor U6842 (N_6842,N_4384,N_4133);
nor U6843 (N_6843,N_2903,N_2515);
nor U6844 (N_6844,N_2875,N_2867);
and U6845 (N_6845,N_2576,N_2635);
nor U6846 (N_6846,N_2681,N_4377);
nor U6847 (N_6847,N_2509,N_4116);
xor U6848 (N_6848,N_2792,N_3462);
and U6849 (N_6849,N_4350,N_4594);
nand U6850 (N_6850,N_3639,N_4752);
and U6851 (N_6851,N_4360,N_3883);
xnor U6852 (N_6852,N_4358,N_3870);
nor U6853 (N_6853,N_4101,N_2842);
and U6854 (N_6854,N_4111,N_3670);
nor U6855 (N_6855,N_3141,N_3469);
or U6856 (N_6856,N_4037,N_2908);
nand U6857 (N_6857,N_4751,N_4549);
nand U6858 (N_6858,N_2978,N_2882);
nor U6859 (N_6859,N_4196,N_4838);
nor U6860 (N_6860,N_4358,N_2674);
nor U6861 (N_6861,N_2697,N_4174);
and U6862 (N_6862,N_4706,N_4010);
or U6863 (N_6863,N_3093,N_3180);
xnor U6864 (N_6864,N_4478,N_4268);
or U6865 (N_6865,N_2825,N_4357);
nor U6866 (N_6866,N_3104,N_4503);
nand U6867 (N_6867,N_3525,N_2565);
nor U6868 (N_6868,N_3995,N_4712);
and U6869 (N_6869,N_3576,N_2878);
or U6870 (N_6870,N_4180,N_3676);
and U6871 (N_6871,N_2640,N_4536);
nor U6872 (N_6872,N_2638,N_4494);
nand U6873 (N_6873,N_4132,N_2752);
nand U6874 (N_6874,N_3011,N_2870);
nor U6875 (N_6875,N_2913,N_4553);
nand U6876 (N_6876,N_2561,N_4025);
and U6877 (N_6877,N_4608,N_4093);
and U6878 (N_6878,N_2945,N_3647);
and U6879 (N_6879,N_3587,N_2739);
or U6880 (N_6880,N_2718,N_2670);
and U6881 (N_6881,N_3455,N_3864);
and U6882 (N_6882,N_4705,N_4632);
nand U6883 (N_6883,N_4469,N_3821);
and U6884 (N_6884,N_3838,N_4148);
or U6885 (N_6885,N_3894,N_2674);
nor U6886 (N_6886,N_2692,N_4988);
or U6887 (N_6887,N_4676,N_2970);
nor U6888 (N_6888,N_3222,N_4724);
or U6889 (N_6889,N_2723,N_3155);
nor U6890 (N_6890,N_3685,N_4473);
or U6891 (N_6891,N_4075,N_3357);
nand U6892 (N_6892,N_4450,N_2701);
nand U6893 (N_6893,N_2979,N_2952);
nor U6894 (N_6894,N_4230,N_4944);
nor U6895 (N_6895,N_4970,N_2917);
nand U6896 (N_6896,N_3081,N_3900);
nand U6897 (N_6897,N_3854,N_3216);
and U6898 (N_6898,N_3105,N_4504);
or U6899 (N_6899,N_4871,N_2864);
nor U6900 (N_6900,N_4355,N_3511);
or U6901 (N_6901,N_3785,N_4310);
or U6902 (N_6902,N_3404,N_3263);
nor U6903 (N_6903,N_3066,N_2854);
nand U6904 (N_6904,N_2653,N_4450);
nand U6905 (N_6905,N_2869,N_3129);
and U6906 (N_6906,N_3154,N_2955);
nand U6907 (N_6907,N_4286,N_4486);
or U6908 (N_6908,N_3558,N_3839);
nand U6909 (N_6909,N_3528,N_4483);
nor U6910 (N_6910,N_3345,N_3242);
nor U6911 (N_6911,N_2622,N_4597);
and U6912 (N_6912,N_4086,N_4098);
nand U6913 (N_6913,N_4417,N_2615);
nor U6914 (N_6914,N_2592,N_4774);
nand U6915 (N_6915,N_4435,N_3208);
and U6916 (N_6916,N_4052,N_4648);
nand U6917 (N_6917,N_3854,N_4471);
nor U6918 (N_6918,N_2529,N_3113);
nor U6919 (N_6919,N_4708,N_4558);
or U6920 (N_6920,N_4495,N_3452);
and U6921 (N_6921,N_3907,N_3533);
nor U6922 (N_6922,N_4774,N_3090);
and U6923 (N_6923,N_3250,N_2641);
or U6924 (N_6924,N_2989,N_4191);
and U6925 (N_6925,N_3766,N_4788);
nor U6926 (N_6926,N_4943,N_2516);
or U6927 (N_6927,N_3940,N_3781);
nand U6928 (N_6928,N_3607,N_4958);
nor U6929 (N_6929,N_4720,N_4498);
or U6930 (N_6930,N_3814,N_4816);
or U6931 (N_6931,N_4903,N_4211);
and U6932 (N_6932,N_4604,N_2627);
nand U6933 (N_6933,N_3869,N_4203);
and U6934 (N_6934,N_2663,N_3243);
and U6935 (N_6935,N_3452,N_3341);
and U6936 (N_6936,N_4692,N_2520);
or U6937 (N_6937,N_4001,N_4124);
or U6938 (N_6938,N_3771,N_4339);
or U6939 (N_6939,N_2842,N_3879);
or U6940 (N_6940,N_3023,N_4904);
nand U6941 (N_6941,N_4270,N_3315);
nor U6942 (N_6942,N_3588,N_2608);
and U6943 (N_6943,N_4649,N_3732);
nand U6944 (N_6944,N_3344,N_3643);
nor U6945 (N_6945,N_3962,N_2581);
or U6946 (N_6946,N_4782,N_3912);
nor U6947 (N_6947,N_2991,N_3764);
and U6948 (N_6948,N_4737,N_2919);
nor U6949 (N_6949,N_3338,N_2857);
nor U6950 (N_6950,N_3847,N_3729);
nor U6951 (N_6951,N_3120,N_3157);
or U6952 (N_6952,N_4993,N_3379);
and U6953 (N_6953,N_2746,N_2521);
and U6954 (N_6954,N_2555,N_4921);
nor U6955 (N_6955,N_2827,N_3154);
nand U6956 (N_6956,N_3285,N_4519);
nand U6957 (N_6957,N_4583,N_3291);
and U6958 (N_6958,N_3651,N_4928);
and U6959 (N_6959,N_2643,N_3339);
nand U6960 (N_6960,N_2783,N_4101);
nand U6961 (N_6961,N_4326,N_3264);
or U6962 (N_6962,N_2783,N_4804);
nand U6963 (N_6963,N_4631,N_2623);
nor U6964 (N_6964,N_3825,N_4136);
nand U6965 (N_6965,N_4901,N_3883);
and U6966 (N_6966,N_2593,N_4362);
nand U6967 (N_6967,N_4111,N_4785);
nand U6968 (N_6968,N_3483,N_4791);
and U6969 (N_6969,N_3633,N_3535);
or U6970 (N_6970,N_3938,N_3270);
nor U6971 (N_6971,N_3928,N_4567);
nor U6972 (N_6972,N_3336,N_2544);
or U6973 (N_6973,N_2828,N_3114);
nor U6974 (N_6974,N_3006,N_4904);
nor U6975 (N_6975,N_3076,N_2702);
nor U6976 (N_6976,N_4669,N_3943);
or U6977 (N_6977,N_3516,N_3991);
nand U6978 (N_6978,N_3083,N_3662);
or U6979 (N_6979,N_3610,N_3578);
or U6980 (N_6980,N_2781,N_4153);
nand U6981 (N_6981,N_3267,N_3844);
or U6982 (N_6982,N_4190,N_3294);
or U6983 (N_6983,N_3638,N_2681);
or U6984 (N_6984,N_3404,N_3678);
nor U6985 (N_6985,N_3838,N_2857);
nand U6986 (N_6986,N_4238,N_4522);
nand U6987 (N_6987,N_4165,N_4750);
nor U6988 (N_6988,N_2748,N_4251);
or U6989 (N_6989,N_4662,N_3901);
or U6990 (N_6990,N_4771,N_4866);
and U6991 (N_6991,N_2527,N_4047);
or U6992 (N_6992,N_3116,N_3915);
or U6993 (N_6993,N_4092,N_3310);
nor U6994 (N_6994,N_3507,N_3953);
nor U6995 (N_6995,N_4302,N_4665);
and U6996 (N_6996,N_2969,N_4078);
nand U6997 (N_6997,N_4688,N_4491);
nand U6998 (N_6998,N_3528,N_3230);
or U6999 (N_6999,N_2683,N_4627);
and U7000 (N_7000,N_3521,N_4188);
or U7001 (N_7001,N_4863,N_4580);
and U7002 (N_7002,N_3591,N_2742);
nor U7003 (N_7003,N_3521,N_3639);
nor U7004 (N_7004,N_3652,N_3980);
nand U7005 (N_7005,N_4933,N_4222);
or U7006 (N_7006,N_4160,N_2721);
and U7007 (N_7007,N_3402,N_3142);
or U7008 (N_7008,N_3533,N_2739);
or U7009 (N_7009,N_3651,N_3157);
nand U7010 (N_7010,N_2569,N_4285);
or U7011 (N_7011,N_4509,N_2592);
and U7012 (N_7012,N_2734,N_3972);
and U7013 (N_7013,N_2973,N_3054);
or U7014 (N_7014,N_2535,N_3771);
and U7015 (N_7015,N_4459,N_3402);
nand U7016 (N_7016,N_4214,N_4092);
nor U7017 (N_7017,N_4497,N_2743);
nand U7018 (N_7018,N_4246,N_2612);
nor U7019 (N_7019,N_2606,N_2615);
and U7020 (N_7020,N_2699,N_4156);
and U7021 (N_7021,N_3716,N_4769);
xor U7022 (N_7022,N_3608,N_4349);
nand U7023 (N_7023,N_4840,N_4672);
or U7024 (N_7024,N_3484,N_3431);
and U7025 (N_7025,N_3584,N_4312);
nor U7026 (N_7026,N_4710,N_4176);
and U7027 (N_7027,N_3147,N_3825);
nor U7028 (N_7028,N_4283,N_4030);
or U7029 (N_7029,N_4674,N_4367);
nor U7030 (N_7030,N_4656,N_2572);
and U7031 (N_7031,N_3368,N_3628);
or U7032 (N_7032,N_2921,N_3188);
or U7033 (N_7033,N_2626,N_4243);
and U7034 (N_7034,N_3080,N_3532);
nor U7035 (N_7035,N_4457,N_3814);
nand U7036 (N_7036,N_2725,N_4706);
or U7037 (N_7037,N_3809,N_3797);
and U7038 (N_7038,N_3817,N_4805);
nand U7039 (N_7039,N_3173,N_3935);
or U7040 (N_7040,N_3517,N_4531);
nand U7041 (N_7041,N_2547,N_3659);
nand U7042 (N_7042,N_4896,N_4616);
nor U7043 (N_7043,N_3586,N_4126);
and U7044 (N_7044,N_2592,N_2741);
or U7045 (N_7045,N_4138,N_3273);
nand U7046 (N_7046,N_3670,N_3969);
and U7047 (N_7047,N_4002,N_3156);
or U7048 (N_7048,N_2694,N_2912);
nor U7049 (N_7049,N_3797,N_4596);
or U7050 (N_7050,N_4255,N_3614);
nand U7051 (N_7051,N_4009,N_2921);
nand U7052 (N_7052,N_3910,N_4031);
or U7053 (N_7053,N_3562,N_4361);
nand U7054 (N_7054,N_2867,N_2639);
nand U7055 (N_7055,N_3121,N_4449);
and U7056 (N_7056,N_3172,N_3818);
and U7057 (N_7057,N_3035,N_3585);
and U7058 (N_7058,N_3483,N_4563);
or U7059 (N_7059,N_4200,N_4367);
or U7060 (N_7060,N_4196,N_2529);
nand U7061 (N_7061,N_4461,N_2615);
or U7062 (N_7062,N_3737,N_4338);
nand U7063 (N_7063,N_4309,N_4216);
or U7064 (N_7064,N_2812,N_4679);
or U7065 (N_7065,N_4698,N_4722);
and U7066 (N_7066,N_3577,N_2727);
nor U7067 (N_7067,N_4747,N_2552);
nand U7068 (N_7068,N_3242,N_4093);
nor U7069 (N_7069,N_4436,N_4643);
and U7070 (N_7070,N_3483,N_4080);
nor U7071 (N_7071,N_3128,N_4457);
nor U7072 (N_7072,N_2571,N_3646);
or U7073 (N_7073,N_4628,N_3439);
nand U7074 (N_7074,N_4753,N_4009);
and U7075 (N_7075,N_4644,N_4447);
and U7076 (N_7076,N_3657,N_2738);
or U7077 (N_7077,N_2852,N_4619);
or U7078 (N_7078,N_4845,N_2613);
or U7079 (N_7079,N_4472,N_3456);
or U7080 (N_7080,N_3409,N_3649);
nor U7081 (N_7081,N_4385,N_3786);
and U7082 (N_7082,N_3146,N_2664);
and U7083 (N_7083,N_4699,N_4473);
nor U7084 (N_7084,N_3107,N_3611);
nand U7085 (N_7085,N_3363,N_3907);
or U7086 (N_7086,N_4871,N_3444);
xor U7087 (N_7087,N_2690,N_4922);
nor U7088 (N_7088,N_4422,N_4550);
nand U7089 (N_7089,N_4042,N_3444);
nor U7090 (N_7090,N_3948,N_3651);
xor U7091 (N_7091,N_3363,N_4754);
nand U7092 (N_7092,N_4635,N_3293);
or U7093 (N_7093,N_3304,N_4640);
nor U7094 (N_7094,N_2972,N_3729);
and U7095 (N_7095,N_2878,N_4502);
nand U7096 (N_7096,N_4673,N_4745);
or U7097 (N_7097,N_2633,N_4292);
nand U7098 (N_7098,N_3646,N_3578);
nor U7099 (N_7099,N_3065,N_4709);
or U7100 (N_7100,N_3311,N_2917);
nand U7101 (N_7101,N_3394,N_3466);
or U7102 (N_7102,N_3039,N_4281);
nor U7103 (N_7103,N_3381,N_3764);
nor U7104 (N_7104,N_3304,N_4376);
and U7105 (N_7105,N_4307,N_3026);
nand U7106 (N_7106,N_4208,N_3564);
and U7107 (N_7107,N_4054,N_4993);
and U7108 (N_7108,N_3760,N_4581);
or U7109 (N_7109,N_4586,N_3178);
and U7110 (N_7110,N_4169,N_3699);
nor U7111 (N_7111,N_2582,N_3599);
or U7112 (N_7112,N_4736,N_4072);
and U7113 (N_7113,N_3473,N_4234);
nor U7114 (N_7114,N_3923,N_4284);
nand U7115 (N_7115,N_4256,N_2681);
or U7116 (N_7116,N_4876,N_3685);
nand U7117 (N_7117,N_4200,N_4662);
and U7118 (N_7118,N_4193,N_4141);
nor U7119 (N_7119,N_4501,N_4738);
or U7120 (N_7120,N_2699,N_3867);
and U7121 (N_7121,N_2775,N_4587);
and U7122 (N_7122,N_3157,N_3850);
nand U7123 (N_7123,N_4897,N_2578);
nand U7124 (N_7124,N_3802,N_4262);
or U7125 (N_7125,N_2594,N_3883);
nand U7126 (N_7126,N_2565,N_2852);
or U7127 (N_7127,N_2836,N_3119);
nor U7128 (N_7128,N_3874,N_4568);
nand U7129 (N_7129,N_4869,N_3740);
nor U7130 (N_7130,N_2671,N_3394);
nand U7131 (N_7131,N_3395,N_4998);
nand U7132 (N_7132,N_3859,N_4271);
or U7133 (N_7133,N_3670,N_4390);
or U7134 (N_7134,N_2549,N_4365);
nand U7135 (N_7135,N_2816,N_2781);
and U7136 (N_7136,N_3965,N_3953);
nand U7137 (N_7137,N_4206,N_2939);
nor U7138 (N_7138,N_3542,N_2762);
nor U7139 (N_7139,N_3765,N_3563);
nand U7140 (N_7140,N_4713,N_3477);
nand U7141 (N_7141,N_4278,N_3103);
nand U7142 (N_7142,N_2590,N_4573);
and U7143 (N_7143,N_2608,N_4776);
nand U7144 (N_7144,N_4596,N_4162);
nand U7145 (N_7145,N_3382,N_4604);
or U7146 (N_7146,N_2568,N_2732);
nor U7147 (N_7147,N_4141,N_2858);
nor U7148 (N_7148,N_2913,N_3774);
and U7149 (N_7149,N_4898,N_2719);
or U7150 (N_7150,N_3304,N_4853);
nor U7151 (N_7151,N_4963,N_3685);
and U7152 (N_7152,N_4729,N_4546);
and U7153 (N_7153,N_4720,N_2968);
nand U7154 (N_7154,N_4136,N_3141);
or U7155 (N_7155,N_2957,N_4729);
or U7156 (N_7156,N_3716,N_3578);
nor U7157 (N_7157,N_3854,N_2994);
nand U7158 (N_7158,N_3792,N_4075);
nor U7159 (N_7159,N_4106,N_3408);
nor U7160 (N_7160,N_3880,N_4149);
nand U7161 (N_7161,N_4431,N_3035);
or U7162 (N_7162,N_3388,N_4002);
nand U7163 (N_7163,N_3364,N_4265);
nor U7164 (N_7164,N_4467,N_2557);
nand U7165 (N_7165,N_4104,N_4006);
and U7166 (N_7166,N_3701,N_4399);
nand U7167 (N_7167,N_4736,N_4091);
nor U7168 (N_7168,N_4231,N_3453);
or U7169 (N_7169,N_3252,N_4496);
and U7170 (N_7170,N_2749,N_4264);
or U7171 (N_7171,N_4795,N_4289);
and U7172 (N_7172,N_4934,N_4143);
nand U7173 (N_7173,N_2535,N_3615);
and U7174 (N_7174,N_3981,N_4091);
or U7175 (N_7175,N_2659,N_4656);
nor U7176 (N_7176,N_2526,N_3103);
nand U7177 (N_7177,N_2950,N_3755);
nor U7178 (N_7178,N_4016,N_3111);
and U7179 (N_7179,N_3950,N_4563);
and U7180 (N_7180,N_3702,N_4381);
nand U7181 (N_7181,N_4019,N_3601);
or U7182 (N_7182,N_3011,N_3136);
and U7183 (N_7183,N_3650,N_4863);
and U7184 (N_7184,N_3391,N_3207);
nor U7185 (N_7185,N_3956,N_4398);
nand U7186 (N_7186,N_3827,N_4928);
or U7187 (N_7187,N_2943,N_3393);
nand U7188 (N_7188,N_3323,N_2609);
and U7189 (N_7189,N_2781,N_4508);
nand U7190 (N_7190,N_3775,N_4919);
or U7191 (N_7191,N_3010,N_3008);
nand U7192 (N_7192,N_2863,N_3921);
or U7193 (N_7193,N_4962,N_3174);
nor U7194 (N_7194,N_3092,N_4246);
xnor U7195 (N_7195,N_3674,N_4757);
and U7196 (N_7196,N_2934,N_4710);
nor U7197 (N_7197,N_4368,N_4841);
nor U7198 (N_7198,N_4947,N_3490);
or U7199 (N_7199,N_4407,N_4398);
and U7200 (N_7200,N_3326,N_2932);
and U7201 (N_7201,N_4377,N_3059);
nor U7202 (N_7202,N_2721,N_3589);
nand U7203 (N_7203,N_4678,N_2640);
nand U7204 (N_7204,N_3719,N_3169);
nor U7205 (N_7205,N_4870,N_4593);
nand U7206 (N_7206,N_3848,N_4559);
or U7207 (N_7207,N_4252,N_4585);
nand U7208 (N_7208,N_3544,N_4997);
nand U7209 (N_7209,N_3418,N_3261);
nor U7210 (N_7210,N_2710,N_3620);
nand U7211 (N_7211,N_3517,N_4197);
nor U7212 (N_7212,N_2674,N_3890);
nor U7213 (N_7213,N_3928,N_4686);
nand U7214 (N_7214,N_4695,N_4960);
or U7215 (N_7215,N_3564,N_2981);
nor U7216 (N_7216,N_3190,N_3085);
nor U7217 (N_7217,N_4314,N_3854);
nand U7218 (N_7218,N_4774,N_4142);
or U7219 (N_7219,N_4464,N_4941);
nor U7220 (N_7220,N_4744,N_3830);
or U7221 (N_7221,N_3205,N_4890);
nand U7222 (N_7222,N_2819,N_3608);
or U7223 (N_7223,N_2907,N_4208);
and U7224 (N_7224,N_3642,N_4683);
and U7225 (N_7225,N_2637,N_2598);
nor U7226 (N_7226,N_4920,N_3046);
nand U7227 (N_7227,N_3097,N_4437);
and U7228 (N_7228,N_4440,N_4198);
or U7229 (N_7229,N_3895,N_2626);
and U7230 (N_7230,N_3332,N_2510);
and U7231 (N_7231,N_2901,N_4956);
nor U7232 (N_7232,N_3165,N_2905);
and U7233 (N_7233,N_2816,N_3878);
and U7234 (N_7234,N_3288,N_4222);
and U7235 (N_7235,N_4906,N_3153);
nand U7236 (N_7236,N_4051,N_2733);
nor U7237 (N_7237,N_3925,N_3007);
nand U7238 (N_7238,N_2959,N_4925);
and U7239 (N_7239,N_2919,N_4893);
and U7240 (N_7240,N_2951,N_4434);
nand U7241 (N_7241,N_2741,N_4530);
and U7242 (N_7242,N_4050,N_4153);
xor U7243 (N_7243,N_3448,N_3517);
and U7244 (N_7244,N_3658,N_3500);
nor U7245 (N_7245,N_3578,N_4670);
nand U7246 (N_7246,N_4820,N_4196);
nor U7247 (N_7247,N_3424,N_3680);
and U7248 (N_7248,N_4395,N_4418);
and U7249 (N_7249,N_3638,N_3083);
and U7250 (N_7250,N_4754,N_4672);
or U7251 (N_7251,N_4401,N_4887);
nor U7252 (N_7252,N_3321,N_3212);
or U7253 (N_7253,N_3931,N_3654);
nand U7254 (N_7254,N_2596,N_4064);
nand U7255 (N_7255,N_3567,N_4327);
and U7256 (N_7256,N_3293,N_3704);
nor U7257 (N_7257,N_4255,N_3333);
nand U7258 (N_7258,N_4601,N_3586);
nand U7259 (N_7259,N_4214,N_4450);
or U7260 (N_7260,N_2787,N_4382);
or U7261 (N_7261,N_4511,N_2591);
or U7262 (N_7262,N_2600,N_3393);
nor U7263 (N_7263,N_2952,N_3869);
nand U7264 (N_7264,N_2844,N_4025);
or U7265 (N_7265,N_2776,N_3595);
or U7266 (N_7266,N_3965,N_3366);
and U7267 (N_7267,N_4084,N_2750);
or U7268 (N_7268,N_3314,N_4696);
nand U7269 (N_7269,N_4335,N_3303);
nor U7270 (N_7270,N_2891,N_4228);
and U7271 (N_7271,N_3629,N_3975);
and U7272 (N_7272,N_4263,N_3234);
and U7273 (N_7273,N_3717,N_4187);
nor U7274 (N_7274,N_2694,N_4945);
xnor U7275 (N_7275,N_4675,N_4639);
nor U7276 (N_7276,N_4700,N_3395);
and U7277 (N_7277,N_2501,N_3173);
nor U7278 (N_7278,N_3988,N_3539);
nor U7279 (N_7279,N_3744,N_3279);
nor U7280 (N_7280,N_4595,N_3180);
and U7281 (N_7281,N_2886,N_3515);
nand U7282 (N_7282,N_4071,N_4756);
and U7283 (N_7283,N_4535,N_2842);
nor U7284 (N_7284,N_3131,N_3960);
nor U7285 (N_7285,N_4574,N_2847);
nand U7286 (N_7286,N_4025,N_3942);
nor U7287 (N_7287,N_4551,N_4631);
or U7288 (N_7288,N_3332,N_4880);
or U7289 (N_7289,N_2977,N_3817);
and U7290 (N_7290,N_3813,N_4564);
and U7291 (N_7291,N_4251,N_4630);
nor U7292 (N_7292,N_4773,N_2873);
or U7293 (N_7293,N_4466,N_4887);
nor U7294 (N_7294,N_4002,N_4325);
nor U7295 (N_7295,N_3026,N_4428);
nand U7296 (N_7296,N_2604,N_2543);
and U7297 (N_7297,N_4057,N_4497);
and U7298 (N_7298,N_4216,N_3581);
and U7299 (N_7299,N_3750,N_3481);
or U7300 (N_7300,N_4285,N_4722);
or U7301 (N_7301,N_2720,N_3524);
nor U7302 (N_7302,N_3995,N_4820);
and U7303 (N_7303,N_3160,N_3030);
and U7304 (N_7304,N_3548,N_3071);
nand U7305 (N_7305,N_4999,N_4258);
nor U7306 (N_7306,N_3965,N_2787);
and U7307 (N_7307,N_4040,N_3670);
or U7308 (N_7308,N_3220,N_4219);
or U7309 (N_7309,N_4158,N_4292);
and U7310 (N_7310,N_2537,N_3588);
or U7311 (N_7311,N_3017,N_2634);
nor U7312 (N_7312,N_2962,N_4565);
and U7313 (N_7313,N_3655,N_3687);
and U7314 (N_7314,N_3393,N_4819);
or U7315 (N_7315,N_4536,N_3032);
nor U7316 (N_7316,N_4168,N_3729);
and U7317 (N_7317,N_4917,N_2844);
or U7318 (N_7318,N_3318,N_2817);
nor U7319 (N_7319,N_2799,N_4687);
nor U7320 (N_7320,N_4631,N_4172);
nand U7321 (N_7321,N_3442,N_4972);
or U7322 (N_7322,N_3331,N_2669);
nand U7323 (N_7323,N_4352,N_3124);
nor U7324 (N_7324,N_2769,N_3035);
and U7325 (N_7325,N_3602,N_2525);
xor U7326 (N_7326,N_3514,N_4907);
nand U7327 (N_7327,N_2551,N_2545);
or U7328 (N_7328,N_3131,N_3035);
nor U7329 (N_7329,N_2592,N_2615);
or U7330 (N_7330,N_3036,N_3897);
and U7331 (N_7331,N_4599,N_4152);
and U7332 (N_7332,N_3521,N_4974);
nand U7333 (N_7333,N_3652,N_3033);
and U7334 (N_7334,N_4964,N_3348);
or U7335 (N_7335,N_4312,N_3898);
or U7336 (N_7336,N_3536,N_3410);
nand U7337 (N_7337,N_3967,N_3254);
nor U7338 (N_7338,N_3061,N_4188);
nor U7339 (N_7339,N_4045,N_4498);
or U7340 (N_7340,N_4876,N_3786);
nor U7341 (N_7341,N_3489,N_2663);
or U7342 (N_7342,N_3984,N_4035);
or U7343 (N_7343,N_4692,N_4684);
or U7344 (N_7344,N_4497,N_2729);
or U7345 (N_7345,N_3042,N_2994);
nand U7346 (N_7346,N_2684,N_4253);
nand U7347 (N_7347,N_3078,N_2913);
and U7348 (N_7348,N_4630,N_3333);
and U7349 (N_7349,N_4973,N_4191);
or U7350 (N_7350,N_4029,N_2931);
nand U7351 (N_7351,N_3832,N_4166);
nand U7352 (N_7352,N_3173,N_4941);
and U7353 (N_7353,N_3131,N_4024);
nor U7354 (N_7354,N_3151,N_3976);
nand U7355 (N_7355,N_4923,N_4570);
and U7356 (N_7356,N_3092,N_3387);
and U7357 (N_7357,N_3767,N_2884);
nand U7358 (N_7358,N_3106,N_3834);
or U7359 (N_7359,N_3726,N_4809);
or U7360 (N_7360,N_2782,N_4896);
nor U7361 (N_7361,N_2706,N_4198);
or U7362 (N_7362,N_4951,N_2716);
nand U7363 (N_7363,N_4575,N_2550);
or U7364 (N_7364,N_2961,N_3147);
and U7365 (N_7365,N_2767,N_3186);
nor U7366 (N_7366,N_3754,N_4512);
or U7367 (N_7367,N_2629,N_3694);
nor U7368 (N_7368,N_3469,N_4493);
nor U7369 (N_7369,N_3113,N_4922);
nand U7370 (N_7370,N_4970,N_4748);
nand U7371 (N_7371,N_3336,N_2519);
nor U7372 (N_7372,N_3221,N_2932);
nor U7373 (N_7373,N_4167,N_3683);
or U7374 (N_7374,N_3964,N_4765);
and U7375 (N_7375,N_4965,N_4316);
and U7376 (N_7376,N_4089,N_3068);
and U7377 (N_7377,N_4059,N_2807);
or U7378 (N_7378,N_4286,N_2632);
and U7379 (N_7379,N_4189,N_4300);
nand U7380 (N_7380,N_4791,N_4080);
nor U7381 (N_7381,N_4344,N_2556);
and U7382 (N_7382,N_3616,N_2582);
nor U7383 (N_7383,N_4636,N_3485);
nor U7384 (N_7384,N_2561,N_4356);
or U7385 (N_7385,N_3156,N_3135);
or U7386 (N_7386,N_4534,N_4609);
or U7387 (N_7387,N_3971,N_3132);
or U7388 (N_7388,N_3963,N_2973);
and U7389 (N_7389,N_4848,N_4389);
nor U7390 (N_7390,N_3893,N_2590);
nand U7391 (N_7391,N_4659,N_4212);
and U7392 (N_7392,N_2571,N_3093);
nand U7393 (N_7393,N_4518,N_3832);
and U7394 (N_7394,N_4310,N_3464);
and U7395 (N_7395,N_3670,N_4701);
nand U7396 (N_7396,N_3407,N_4826);
nand U7397 (N_7397,N_4271,N_2560);
nand U7398 (N_7398,N_4662,N_4769);
nor U7399 (N_7399,N_2654,N_4716);
nor U7400 (N_7400,N_3055,N_3138);
and U7401 (N_7401,N_2824,N_4262);
nor U7402 (N_7402,N_3123,N_4897);
nand U7403 (N_7403,N_3010,N_3083);
and U7404 (N_7404,N_4253,N_4216);
nor U7405 (N_7405,N_2876,N_2645);
and U7406 (N_7406,N_2961,N_3380);
nand U7407 (N_7407,N_3217,N_4134);
or U7408 (N_7408,N_4363,N_3268);
or U7409 (N_7409,N_3568,N_4618);
and U7410 (N_7410,N_4137,N_4057);
nor U7411 (N_7411,N_4486,N_4258);
and U7412 (N_7412,N_2558,N_4844);
nor U7413 (N_7413,N_3845,N_4833);
nor U7414 (N_7414,N_4692,N_4901);
and U7415 (N_7415,N_3898,N_4611);
and U7416 (N_7416,N_4024,N_3449);
nor U7417 (N_7417,N_2986,N_3001);
nor U7418 (N_7418,N_4791,N_2871);
or U7419 (N_7419,N_3053,N_3510);
and U7420 (N_7420,N_3027,N_2756);
nor U7421 (N_7421,N_4536,N_3197);
nand U7422 (N_7422,N_4634,N_3781);
and U7423 (N_7423,N_4738,N_2933);
nor U7424 (N_7424,N_4136,N_4422);
nor U7425 (N_7425,N_4371,N_3043);
and U7426 (N_7426,N_4994,N_4188);
nand U7427 (N_7427,N_2819,N_3632);
nor U7428 (N_7428,N_3101,N_4664);
nor U7429 (N_7429,N_4754,N_4980);
nor U7430 (N_7430,N_3608,N_2519);
nor U7431 (N_7431,N_3816,N_3726);
nand U7432 (N_7432,N_3828,N_4820);
nor U7433 (N_7433,N_4607,N_2869);
nor U7434 (N_7434,N_3268,N_3948);
and U7435 (N_7435,N_4568,N_3177);
nor U7436 (N_7436,N_2966,N_2747);
and U7437 (N_7437,N_3535,N_3886);
or U7438 (N_7438,N_3569,N_4136);
and U7439 (N_7439,N_3138,N_2824);
nand U7440 (N_7440,N_3981,N_4450);
or U7441 (N_7441,N_3812,N_4309);
or U7442 (N_7442,N_3301,N_4536);
nor U7443 (N_7443,N_3222,N_3719);
or U7444 (N_7444,N_3508,N_2759);
nor U7445 (N_7445,N_3458,N_4670);
and U7446 (N_7446,N_3014,N_4093);
nand U7447 (N_7447,N_4031,N_4931);
nor U7448 (N_7448,N_3520,N_3801);
nor U7449 (N_7449,N_3648,N_4619);
and U7450 (N_7450,N_3145,N_2608);
and U7451 (N_7451,N_2980,N_3852);
nand U7452 (N_7452,N_4756,N_3645);
and U7453 (N_7453,N_3183,N_4415);
nand U7454 (N_7454,N_3580,N_2692);
nand U7455 (N_7455,N_4909,N_4721);
nor U7456 (N_7456,N_3716,N_4793);
and U7457 (N_7457,N_4748,N_2971);
nor U7458 (N_7458,N_2606,N_3234);
nor U7459 (N_7459,N_4928,N_2511);
nand U7460 (N_7460,N_4247,N_4134);
nor U7461 (N_7461,N_3237,N_4095);
nor U7462 (N_7462,N_3816,N_4936);
nor U7463 (N_7463,N_2953,N_2993);
nand U7464 (N_7464,N_3510,N_2854);
or U7465 (N_7465,N_4511,N_3455);
nand U7466 (N_7466,N_2906,N_3152);
nand U7467 (N_7467,N_4802,N_4698);
and U7468 (N_7468,N_3239,N_4872);
and U7469 (N_7469,N_4492,N_2916);
nor U7470 (N_7470,N_3363,N_4661);
and U7471 (N_7471,N_4750,N_4776);
and U7472 (N_7472,N_4943,N_4524);
or U7473 (N_7473,N_3583,N_3398);
and U7474 (N_7474,N_4412,N_4976);
or U7475 (N_7475,N_2586,N_2707);
nor U7476 (N_7476,N_3033,N_4257);
nand U7477 (N_7477,N_4440,N_3884);
nor U7478 (N_7478,N_4039,N_4208);
and U7479 (N_7479,N_4583,N_4079);
and U7480 (N_7480,N_3866,N_3731);
nor U7481 (N_7481,N_4534,N_4568);
nor U7482 (N_7482,N_2875,N_2976);
and U7483 (N_7483,N_4628,N_3182);
nand U7484 (N_7484,N_3595,N_2857);
or U7485 (N_7485,N_4326,N_3633);
or U7486 (N_7486,N_2827,N_4998);
or U7487 (N_7487,N_3439,N_4439);
and U7488 (N_7488,N_4975,N_2511);
and U7489 (N_7489,N_3411,N_2681);
or U7490 (N_7490,N_3698,N_3751);
or U7491 (N_7491,N_3950,N_4976);
or U7492 (N_7492,N_4899,N_4458);
and U7493 (N_7493,N_4996,N_2622);
or U7494 (N_7494,N_3153,N_2864);
and U7495 (N_7495,N_3801,N_3478);
nand U7496 (N_7496,N_4678,N_4264);
or U7497 (N_7497,N_2833,N_4441);
nand U7498 (N_7498,N_3107,N_3961);
nand U7499 (N_7499,N_2579,N_4664);
nor U7500 (N_7500,N_5609,N_6383);
and U7501 (N_7501,N_7234,N_7201);
nor U7502 (N_7502,N_5747,N_7241);
nor U7503 (N_7503,N_5323,N_7403);
and U7504 (N_7504,N_5956,N_6953);
or U7505 (N_7505,N_6710,N_5426);
nor U7506 (N_7506,N_6603,N_5481);
or U7507 (N_7507,N_5041,N_5480);
or U7508 (N_7508,N_6832,N_6633);
and U7509 (N_7509,N_6572,N_6017);
or U7510 (N_7510,N_6778,N_5927);
or U7511 (N_7511,N_7172,N_5406);
nand U7512 (N_7512,N_5219,N_5174);
and U7513 (N_7513,N_7231,N_5212);
or U7514 (N_7514,N_6210,N_7390);
nor U7515 (N_7515,N_6433,N_6137);
and U7516 (N_7516,N_6645,N_7027);
nand U7517 (N_7517,N_7362,N_6942);
and U7518 (N_7518,N_5033,N_6556);
and U7519 (N_7519,N_7113,N_5191);
nor U7520 (N_7520,N_6698,N_5572);
and U7521 (N_7521,N_6764,N_5874);
or U7522 (N_7522,N_7026,N_6273);
and U7523 (N_7523,N_5388,N_7186);
nand U7524 (N_7524,N_5961,N_5692);
nand U7525 (N_7525,N_6179,N_7211);
and U7526 (N_7526,N_5976,N_5830);
or U7527 (N_7527,N_6321,N_6399);
nor U7528 (N_7528,N_6613,N_6684);
nand U7529 (N_7529,N_5706,N_6673);
xnor U7530 (N_7530,N_5040,N_6982);
and U7531 (N_7531,N_6694,N_6824);
and U7532 (N_7532,N_6790,N_6371);
nand U7533 (N_7533,N_5799,N_7347);
nand U7534 (N_7534,N_5889,N_7484);
nor U7535 (N_7535,N_5119,N_7233);
and U7536 (N_7536,N_6238,N_5300);
nor U7537 (N_7537,N_5285,N_6611);
nor U7538 (N_7538,N_5849,N_6742);
nand U7539 (N_7539,N_6812,N_6053);
or U7540 (N_7540,N_5647,N_6249);
nor U7541 (N_7541,N_5812,N_5937);
and U7542 (N_7542,N_5284,N_5657);
nor U7543 (N_7543,N_5535,N_5909);
xor U7544 (N_7544,N_5063,N_6261);
nand U7545 (N_7545,N_5037,N_7358);
and U7546 (N_7546,N_7183,N_7368);
nor U7547 (N_7547,N_5577,N_7245);
and U7548 (N_7548,N_6749,N_7124);
or U7549 (N_7549,N_5146,N_7260);
and U7550 (N_7550,N_6706,N_5842);
or U7551 (N_7551,N_5258,N_5507);
and U7552 (N_7552,N_5316,N_6173);
nand U7553 (N_7553,N_6935,N_5837);
xor U7554 (N_7554,N_6374,N_5147);
nand U7555 (N_7555,N_7248,N_5730);
and U7556 (N_7556,N_7141,N_6796);
or U7557 (N_7557,N_6503,N_5352);
nand U7558 (N_7558,N_6941,N_5006);
nor U7559 (N_7559,N_6366,N_7434);
nand U7560 (N_7560,N_7407,N_6855);
nor U7561 (N_7561,N_6901,N_5638);
or U7562 (N_7562,N_5190,N_5298);
or U7563 (N_7563,N_6203,N_6952);
or U7564 (N_7564,N_7048,N_7262);
nor U7565 (N_7565,N_6422,N_7275);
nand U7566 (N_7566,N_5943,N_7497);
nor U7567 (N_7567,N_6477,N_5169);
nor U7568 (N_7568,N_5014,N_5030);
nand U7569 (N_7569,N_6275,N_7116);
nand U7570 (N_7570,N_6589,N_6816);
nor U7571 (N_7571,N_6489,N_7353);
and U7572 (N_7572,N_5168,N_7273);
or U7573 (N_7573,N_6723,N_5674);
or U7574 (N_7574,N_5189,N_5914);
and U7575 (N_7575,N_6926,N_6154);
nand U7576 (N_7576,N_6637,N_5408);
nor U7577 (N_7577,N_5834,N_6703);
or U7578 (N_7578,N_5630,N_6269);
nor U7579 (N_7579,N_5097,N_5758);
or U7580 (N_7580,N_6232,N_6863);
and U7581 (N_7581,N_5533,N_6482);
and U7582 (N_7582,N_6084,N_5558);
or U7583 (N_7583,N_6991,N_5965);
nor U7584 (N_7584,N_6376,N_5347);
nand U7585 (N_7585,N_6225,N_5788);
nor U7586 (N_7586,N_6534,N_5694);
and U7587 (N_7587,N_7415,N_5962);
nor U7588 (N_7588,N_5115,N_6913);
nand U7589 (N_7589,N_5871,N_6467);
nand U7590 (N_7590,N_6539,N_6256);
nor U7591 (N_7591,N_7418,N_5882);
and U7592 (N_7592,N_6091,N_6971);
nor U7593 (N_7593,N_5492,N_6387);
or U7594 (N_7594,N_7445,N_6357);
nor U7595 (N_7595,N_6214,N_6345);
or U7596 (N_7596,N_7417,N_5083);
or U7597 (N_7597,N_6353,N_6152);
or U7598 (N_7598,N_6653,N_5600);
and U7599 (N_7599,N_7204,N_6454);
nand U7600 (N_7600,N_6903,N_5920);
and U7601 (N_7601,N_7144,N_5958);
nor U7602 (N_7602,N_5755,N_5059);
or U7603 (N_7603,N_5132,N_6831);
nor U7604 (N_7604,N_5238,N_5936);
nand U7605 (N_7605,N_6162,N_6209);
nand U7606 (N_7606,N_7406,N_6530);
and U7607 (N_7607,N_6537,N_5445);
and U7608 (N_7608,N_5699,N_5090);
nor U7609 (N_7609,N_7392,N_6580);
nand U7610 (N_7610,N_7354,N_5534);
and U7611 (N_7611,N_5829,N_5227);
and U7612 (N_7612,N_6986,N_5170);
and U7613 (N_7613,N_6317,N_6533);
nand U7614 (N_7614,N_5813,N_7485);
nand U7615 (N_7615,N_5341,N_5230);
and U7616 (N_7616,N_7261,N_6617);
or U7617 (N_7617,N_6767,N_6818);
nand U7618 (N_7618,N_5269,N_6775);
nor U7619 (N_7619,N_6564,N_6121);
nor U7620 (N_7620,N_5476,N_6429);
or U7621 (N_7621,N_5826,N_7377);
nor U7622 (N_7622,N_7054,N_6751);
or U7623 (N_7623,N_6095,N_6453);
or U7624 (N_7624,N_6964,N_6246);
xor U7625 (N_7625,N_6546,N_6958);
nor U7626 (N_7626,N_7218,N_6829);
and U7627 (N_7627,N_5801,N_7119);
nor U7628 (N_7628,N_6923,N_5360);
nor U7629 (N_7629,N_6891,N_5952);
nand U7630 (N_7630,N_6307,N_6212);
or U7631 (N_7631,N_6948,N_6359);
and U7632 (N_7632,N_5397,N_6583);
or U7633 (N_7633,N_5792,N_6271);
or U7634 (N_7634,N_6610,N_5421);
nand U7635 (N_7635,N_5363,N_5550);
nor U7636 (N_7636,N_6532,N_6318);
or U7637 (N_7637,N_6013,N_5164);
nor U7638 (N_7638,N_6576,N_5683);
nand U7639 (N_7639,N_6126,N_7247);
or U7640 (N_7640,N_6227,N_5396);
nand U7641 (N_7641,N_5586,N_6880);
nor U7642 (N_7642,N_5765,N_7151);
or U7643 (N_7643,N_6919,N_7177);
nand U7644 (N_7644,N_7356,N_7076);
nand U7645 (N_7645,N_5667,N_5422);
nand U7646 (N_7646,N_5085,N_7195);
nand U7647 (N_7647,N_7249,N_6783);
or U7648 (N_7648,N_6067,N_5731);
nand U7649 (N_7649,N_6412,N_5478);
or U7650 (N_7650,N_5263,N_5368);
nand U7651 (N_7651,N_7313,N_5637);
nor U7652 (N_7652,N_5656,N_7022);
nand U7653 (N_7653,N_6635,N_6445);
nor U7654 (N_7654,N_6315,N_7315);
and U7655 (N_7655,N_6608,N_7496);
or U7656 (N_7656,N_5917,N_5622);
or U7657 (N_7657,N_5128,N_7178);
nor U7658 (N_7658,N_6016,N_6255);
nand U7659 (N_7659,N_5262,N_6312);
nor U7660 (N_7660,N_6403,N_5963);
or U7661 (N_7661,N_6064,N_6838);
nand U7662 (N_7662,N_6221,N_6052);
xnor U7663 (N_7663,N_6043,N_7030);
or U7664 (N_7664,N_5562,N_7424);
or U7665 (N_7665,N_7305,N_6878);
nor U7666 (N_7666,N_6171,N_5935);
nand U7667 (N_7667,N_6451,N_5545);
or U7668 (N_7668,N_6093,N_6921);
nor U7669 (N_7669,N_5611,N_5782);
and U7670 (N_7670,N_5948,N_5441);
nor U7671 (N_7671,N_6031,N_5015);
nand U7672 (N_7672,N_5668,N_5252);
nand U7673 (N_7673,N_5618,N_5053);
nand U7674 (N_7674,N_5140,N_6675);
or U7675 (N_7675,N_7345,N_6346);
xnor U7676 (N_7676,N_5530,N_7367);
and U7677 (N_7677,N_6995,N_5631);
nor U7678 (N_7678,N_6023,N_6826);
and U7679 (N_7679,N_6444,N_5867);
or U7680 (N_7680,N_6699,N_7490);
or U7681 (N_7681,N_5444,N_7146);
and U7682 (N_7682,N_5159,N_5746);
nand U7683 (N_7683,N_5399,N_7210);
or U7684 (N_7684,N_6130,N_7499);
nor U7685 (N_7685,N_6365,N_7135);
and U7686 (N_7686,N_6298,N_7012);
nor U7687 (N_7687,N_5760,N_6145);
nor U7688 (N_7688,N_5453,N_6036);
and U7689 (N_7689,N_6224,N_5621);
or U7690 (N_7690,N_6734,N_6394);
nand U7691 (N_7691,N_7366,N_5464);
nand U7692 (N_7692,N_5215,N_7268);
and U7693 (N_7693,N_7306,N_7067);
nor U7694 (N_7694,N_5127,N_6956);
and U7695 (N_7695,N_6614,N_6794);
and U7696 (N_7696,N_7021,N_5903);
nor U7697 (N_7697,N_5019,N_7364);
or U7698 (N_7698,N_6343,N_5954);
nor U7699 (N_7699,N_6989,N_7057);
and U7700 (N_7700,N_6306,N_5922);
or U7701 (N_7701,N_5947,N_7117);
nand U7702 (N_7702,N_6491,N_5243);
and U7703 (N_7703,N_6100,N_6108);
nor U7704 (N_7704,N_5220,N_6175);
or U7705 (N_7705,N_6678,N_5328);
or U7706 (N_7706,N_6417,N_6500);
and U7707 (N_7707,N_6805,N_6178);
nand U7708 (N_7708,N_5780,N_5291);
and U7709 (N_7709,N_6882,N_6239);
nor U7710 (N_7710,N_6372,N_5216);
nor U7711 (N_7711,N_5384,N_5757);
nand U7712 (N_7712,N_5955,N_5725);
nor U7713 (N_7713,N_5723,N_7471);
nand U7714 (N_7714,N_5358,N_7388);
or U7715 (N_7715,N_5701,N_7182);
and U7716 (N_7716,N_5972,N_6801);
and U7717 (N_7717,N_5791,N_5264);
nor U7718 (N_7718,N_7425,N_6927);
nor U7719 (N_7719,N_6643,N_6940);
or U7720 (N_7720,N_7221,N_6630);
nand U7721 (N_7721,N_5563,N_6769);
nand U7722 (N_7722,N_5244,N_6311);
nand U7723 (N_7723,N_6949,N_6076);
and U7724 (N_7724,N_7065,N_5850);
or U7725 (N_7725,N_5382,N_5309);
and U7726 (N_7726,N_6174,N_5373);
and U7727 (N_7727,N_7162,N_7126);
nor U7728 (N_7728,N_6435,N_7108);
nand U7729 (N_7729,N_6048,N_6204);
or U7730 (N_7730,N_7277,N_6468);
nand U7731 (N_7731,N_5715,N_5819);
or U7732 (N_7732,N_5361,N_5815);
nor U7733 (N_7733,N_5769,N_5783);
or U7734 (N_7734,N_7166,N_6811);
nand U7735 (N_7735,N_7045,N_5324);
nand U7736 (N_7736,N_5167,N_5482);
nor U7737 (N_7737,N_6819,N_6757);
and U7738 (N_7738,N_6642,N_7335);
nand U7739 (N_7739,N_7256,N_5392);
and U7740 (N_7740,N_6887,N_5145);
or U7741 (N_7741,N_5932,N_6388);
or U7742 (N_7742,N_7292,N_6127);
nor U7743 (N_7743,N_7395,N_6163);
and U7744 (N_7744,N_5513,N_7034);
and U7745 (N_7745,N_6857,N_5756);
nand U7746 (N_7746,N_6234,N_5455);
nand U7747 (N_7747,N_5185,N_7293);
or U7748 (N_7748,N_6281,N_7495);
nor U7749 (N_7749,N_6763,N_6984);
nor U7750 (N_7750,N_5957,N_5894);
and U7751 (N_7751,N_7372,N_7373);
and U7752 (N_7752,N_7308,N_5696);
or U7753 (N_7753,N_6265,N_5193);
and U7754 (N_7754,N_5865,N_6776);
or U7755 (N_7755,N_6244,N_5036);
nand U7756 (N_7756,N_7160,N_5732);
nand U7757 (N_7757,N_7338,N_6514);
nor U7758 (N_7758,N_6110,N_5854);
or U7759 (N_7759,N_5133,N_5662);
nor U7760 (N_7760,N_6917,N_6449);
or U7761 (N_7761,N_6700,N_6762);
and U7762 (N_7762,N_6338,N_6784);
nand U7763 (N_7763,N_7079,N_6011);
nor U7764 (N_7764,N_7159,N_5497);
or U7765 (N_7765,N_6139,N_5992);
and U7766 (N_7766,N_7174,N_6628);
nor U7767 (N_7767,N_6325,N_5239);
or U7768 (N_7768,N_5259,N_6545);
or U7769 (N_7769,N_7439,N_5110);
and U7770 (N_7770,N_5024,N_6665);
nand U7771 (N_7771,N_6025,N_6791);
and U7772 (N_7772,N_7463,N_6022);
and U7773 (N_7773,N_6492,N_5559);
and U7774 (N_7774,N_6159,N_5817);
nand U7775 (N_7775,N_5364,N_5439);
nor U7776 (N_7776,N_5653,N_6198);
nor U7777 (N_7777,N_7399,N_7036);
xnor U7778 (N_7778,N_7133,N_7384);
nand U7779 (N_7779,N_6360,N_6190);
and U7780 (N_7780,N_5051,N_5606);
and U7781 (N_7781,N_7440,N_6308);
or U7782 (N_7782,N_5357,N_5296);
or U7783 (N_7783,N_5999,N_7237);
or U7784 (N_7784,N_7192,N_5582);
and U7785 (N_7785,N_7123,N_5852);
and U7786 (N_7786,N_5736,N_6124);
and U7787 (N_7787,N_6531,N_5425);
nor U7788 (N_7788,N_7043,N_5861);
nor U7789 (N_7789,N_6578,N_6443);
and U7790 (N_7790,N_5613,N_6994);
and U7791 (N_7791,N_5431,N_7351);
nand U7792 (N_7792,N_7452,N_5248);
or U7793 (N_7793,N_7369,N_5828);
and U7794 (N_7794,N_5002,N_7291);
and U7795 (N_7795,N_6077,N_7120);
nor U7796 (N_7796,N_5569,N_5797);
nand U7797 (N_7797,N_6535,N_5111);
nor U7798 (N_7798,N_5458,N_6418);
and U7799 (N_7799,N_6745,N_6407);
nor U7800 (N_7800,N_7180,N_5411);
or U7801 (N_7801,N_5608,N_5345);
nand U7802 (N_7802,N_6090,N_6020);
nand U7803 (N_7803,N_7431,N_7281);
or U7804 (N_7804,N_7492,N_5934);
or U7805 (N_7805,N_5319,N_7441);
nor U7806 (N_7806,N_5578,N_5054);
or U7807 (N_7807,N_7326,N_5073);
nand U7808 (N_7808,N_6396,N_5317);
xnor U7809 (N_7809,N_6223,N_5071);
and U7810 (N_7810,N_7264,N_6722);
nand U7811 (N_7811,N_6414,N_5135);
nand U7812 (N_7812,N_7299,N_5888);
and U7813 (N_7813,N_5234,N_7413);
or U7814 (N_7814,N_6014,N_5270);
and U7815 (N_7815,N_7469,N_5523);
and U7816 (N_7816,N_7327,N_6266);
nand U7817 (N_7817,N_6992,N_7129);
and U7818 (N_7818,N_7111,N_5099);
nand U7819 (N_7819,N_6285,N_6725);
or U7820 (N_7820,N_5855,N_5104);
nor U7821 (N_7821,N_5078,N_6391);
and U7822 (N_7822,N_7419,N_6447);
or U7823 (N_7823,N_7003,N_6029);
nand U7824 (N_7824,N_5878,N_6632);
nand U7825 (N_7825,N_6355,N_7197);
nor U7826 (N_7826,N_5679,N_5820);
nand U7827 (N_7827,N_7226,N_6129);
nor U7828 (N_7828,N_5579,N_6465);
and U7829 (N_7829,N_5503,N_7489);
nand U7830 (N_7830,N_6334,N_6189);
or U7831 (N_7831,N_6906,N_5225);
nor U7832 (N_7832,N_7296,N_6566);
or U7833 (N_7833,N_5575,N_6715);
or U7834 (N_7834,N_6720,N_5774);
and U7835 (N_7835,N_5824,N_6905);
or U7836 (N_7836,N_7199,N_6263);
nor U7837 (N_7837,N_7018,N_5012);
nor U7838 (N_7838,N_5304,N_5539);
and U7839 (N_7839,N_7069,N_6835);
and U7840 (N_7840,N_7223,N_6044);
and U7841 (N_7841,N_5982,N_7044);
or U7842 (N_7842,N_6647,N_5466);
nand U7843 (N_7843,N_6588,N_5342);
and U7844 (N_7844,N_7483,N_6466);
nand U7845 (N_7845,N_6915,N_6523);
and U7846 (N_7846,N_7041,N_5966);
nand U7847 (N_7847,N_5543,N_5542);
nor U7848 (N_7848,N_5344,N_7193);
or U7849 (N_7849,N_6718,N_7039);
or U7850 (N_7850,N_5351,N_5107);
nor U7851 (N_7851,N_5931,N_6691);
nand U7852 (N_7852,N_6657,N_5869);
and U7853 (N_7853,N_5000,N_5209);
and U7854 (N_7854,N_7167,N_5432);
nand U7855 (N_7855,N_5585,N_6813);
or U7856 (N_7856,N_5899,N_6208);
and U7857 (N_7857,N_5420,N_6547);
nor U7858 (N_7858,N_5506,N_5485);
nand U7859 (N_7859,N_6393,N_6096);
nor U7860 (N_7860,N_7380,N_7114);
nor U7861 (N_7861,N_6881,N_6441);
nor U7862 (N_7862,N_5022,N_5528);
or U7863 (N_7863,N_6030,N_5768);
and U7864 (N_7864,N_6854,N_6335);
nor U7865 (N_7865,N_5138,N_7101);
nand U7866 (N_7866,N_6220,N_5515);
nor U7867 (N_7867,N_6283,N_7215);
or U7868 (N_7868,N_7156,N_6600);
nand U7869 (N_7869,N_5703,N_6770);
nand U7870 (N_7870,N_6962,N_6487);
and U7871 (N_7871,N_6978,N_7360);
xor U7872 (N_7872,N_6302,N_6228);
nand U7873 (N_7873,N_5977,N_5417);
and U7874 (N_7874,N_7206,N_5202);
nor U7875 (N_7875,N_6033,N_5413);
nand U7876 (N_7876,N_7051,N_7448);
or U7877 (N_7877,N_6860,N_7017);
or U7878 (N_7878,N_6106,N_6928);
nor U7879 (N_7879,N_6682,N_7350);
nand U7880 (N_7880,N_7389,N_6512);
or U7881 (N_7881,N_5685,N_6621);
nor U7882 (N_7882,N_5847,N_6649);
nor U7883 (N_7883,N_6596,N_7449);
and U7884 (N_7884,N_7414,N_7361);
nand U7885 (N_7885,N_7333,N_5446);
nand U7886 (N_7886,N_6766,N_5025);
nor U7887 (N_7887,N_5489,N_6158);
nand U7888 (N_7888,N_5483,N_5203);
nand U7889 (N_7889,N_5770,N_5069);
and U7890 (N_7890,N_5772,N_5437);
and U7891 (N_7891,N_6042,N_7427);
or U7892 (N_7892,N_5112,N_5359);
or U7893 (N_7893,N_5374,N_6499);
or U7894 (N_7894,N_5429,N_5367);
and U7895 (N_7895,N_5996,N_6544);
and U7896 (N_7896,N_5863,N_5348);
and U7897 (N_7897,N_6571,N_5557);
nand U7898 (N_7898,N_5192,N_5560);
nor U7899 (N_7899,N_6507,N_7093);
and U7900 (N_7900,N_5139,N_5044);
and U7901 (N_7901,N_6842,N_6303);
or U7902 (N_7902,N_7011,N_5349);
nor U7903 (N_7903,N_5116,N_5880);
or U7904 (N_7904,N_7105,N_6001);
nor U7905 (N_7905,N_5526,N_5405);
nand U7906 (N_7906,N_5516,N_6624);
and U7907 (N_7907,N_5789,N_7229);
nand U7908 (N_7908,N_6666,N_5028);
nor U7909 (N_7909,N_7435,N_5313);
and U7910 (N_7910,N_6756,N_5334);
or U7911 (N_7911,N_6641,N_7236);
and U7912 (N_7912,N_5623,N_5501);
nand U7913 (N_7913,N_5009,N_7410);
and U7914 (N_7914,N_5026,N_6264);
or U7915 (N_7915,N_5096,N_5993);
and U7916 (N_7916,N_6977,N_6932);
and U7917 (N_7917,N_7438,N_6591);
and U7918 (N_7918,N_7409,N_5017);
nand U7919 (N_7919,N_5231,N_5018);
nand U7920 (N_7920,N_5840,N_6494);
xnor U7921 (N_7921,N_7282,N_6340);
and U7922 (N_7922,N_5564,N_5237);
nor U7923 (N_7923,N_6350,N_7283);
or U7924 (N_7924,N_5356,N_5720);
nand U7925 (N_7925,N_6134,N_7266);
and U7926 (N_7926,N_6587,N_6486);
and U7927 (N_7927,N_7478,N_5401);
nor U7928 (N_7928,N_7243,N_5800);
and U7929 (N_7929,N_7019,N_7458);
and U7930 (N_7930,N_6890,N_5551);
or U7931 (N_7931,N_5514,N_5142);
or U7932 (N_7932,N_7295,N_6884);
or U7933 (N_7933,N_5113,N_7175);
nor U7934 (N_7934,N_7009,N_5204);
or U7935 (N_7935,N_5213,N_6205);
and U7936 (N_7936,N_5469,N_7224);
nor U7937 (N_7937,N_5487,N_5643);
and U7938 (N_7938,N_7442,N_7163);
nor U7939 (N_7939,N_5438,N_6735);
or U7940 (N_7940,N_6889,N_6087);
nor U7941 (N_7941,N_5060,N_6605);
and U7942 (N_7942,N_6774,N_6744);
nor U7943 (N_7943,N_6071,N_6851);
and U7944 (N_7944,N_5123,N_5717);
or U7945 (N_7945,N_5652,N_5790);
or U7946 (N_7946,N_6092,N_7063);
and U7947 (N_7947,N_5918,N_6348);
nand U7948 (N_7948,N_5921,N_5404);
and U7949 (N_7949,N_5953,N_5946);
and U7950 (N_7950,N_5214,N_6590);
nor U7951 (N_7951,N_5410,N_7491);
nor U7952 (N_7952,N_5346,N_5177);
nor U7953 (N_7953,N_5959,N_5767);
and U7954 (N_7954,N_7334,N_7055);
nor U7955 (N_7955,N_6434,N_5048);
or U7956 (N_7956,N_5595,N_7397);
nor U7957 (N_7957,N_7066,N_6079);
nand U7958 (N_7958,N_6191,N_6692);
nor U7959 (N_7959,N_7081,N_5058);
or U7960 (N_7960,N_5076,N_6946);
nand U7961 (N_7961,N_7205,N_7278);
or U7962 (N_7962,N_6050,N_5527);
or U7963 (N_7963,N_5089,N_6607);
nand U7964 (N_7964,N_6620,N_7190);
nand U7965 (N_7965,N_6278,N_5763);
and U7966 (N_7966,N_7164,N_5787);
and U7967 (N_7967,N_5891,N_6250);
or U7968 (N_7968,N_6746,N_5495);
nor U7969 (N_7969,N_5010,N_5452);
or U7970 (N_7970,N_5198,N_5141);
nor U7971 (N_7971,N_6823,N_5279);
nor U7972 (N_7972,N_5393,N_5427);
nor U7973 (N_7973,N_6085,N_7060);
nand U7974 (N_7974,N_6408,N_5754);
or U7975 (N_7975,N_6219,N_6475);
or U7976 (N_7976,N_5727,N_7150);
and U7977 (N_7977,N_5713,N_7487);
nor U7978 (N_7978,N_5383,N_5556);
nand U7979 (N_7979,N_5330,N_7212);
or U7980 (N_7980,N_5581,N_5843);
nor U7981 (N_7981,N_5806,N_6019);
nand U7982 (N_7982,N_5504,N_6027);
or U7983 (N_7983,N_7073,N_5565);
and U7984 (N_7984,N_5510,N_5103);
nor U7985 (N_7985,N_5052,N_5978);
or U7986 (N_7986,N_7336,N_5794);
and U7987 (N_7987,N_6845,N_5136);
nor U7988 (N_7988,N_6222,N_6287);
or U7989 (N_7989,N_5289,N_6216);
nor U7990 (N_7990,N_5082,N_7202);
nand U7991 (N_7991,N_6515,N_6146);
nand U7992 (N_7992,N_7421,N_6380);
nand U7993 (N_7993,N_5988,N_6669);
nand U7994 (N_7994,N_5380,N_6332);
or U7995 (N_7995,N_7468,N_7401);
nor U7996 (N_7996,N_7383,N_5066);
or U7997 (N_7997,N_5288,N_7013);
or U7998 (N_7998,N_5120,N_6554);
nand U7999 (N_7999,N_5034,N_6323);
and U8000 (N_8000,N_6858,N_6230);
or U8001 (N_8001,N_6395,N_5302);
and U8002 (N_8002,N_5599,N_5062);
nor U8003 (N_8003,N_7238,N_5315);
nand U8004 (N_8004,N_7128,N_5570);
or U8005 (N_8005,N_5845,N_6284);
nor U8006 (N_8006,N_6663,N_6517);
nor U8007 (N_8007,N_6870,N_5131);
and U8008 (N_8008,N_6289,N_6474);
nand U8009 (N_8009,N_6182,N_7494);
or U8010 (N_8010,N_6728,N_6574);
or U8011 (N_8011,N_7109,N_7284);
nand U8012 (N_8012,N_6985,N_5741);
and U8013 (N_8013,N_6765,N_5661);
nor U8014 (N_8014,N_5877,N_6426);
or U8015 (N_8015,N_6358,N_7118);
nor U8016 (N_8016,N_6555,N_5529);
nand U8017 (N_8017,N_7454,N_6864);
nand U8018 (N_8018,N_7138,N_5496);
nor U8019 (N_8019,N_6593,N_6789);
nor U8020 (N_8020,N_6616,N_6651);
or U8021 (N_8021,N_5463,N_6478);
or U8022 (N_8022,N_7082,N_6413);
and U8023 (N_8023,N_5626,N_6837);
or U8024 (N_8024,N_5998,N_7049);
and U8025 (N_8025,N_7476,N_6912);
nor U8026 (N_8026,N_7290,N_5933);
or U8027 (N_8027,N_5250,N_6111);
and U8028 (N_8028,N_7411,N_5617);
and U8029 (N_8029,N_5841,N_5016);
and U8030 (N_8030,N_6646,N_5566);
nor U8031 (N_8031,N_6595,N_6313);
nor U8032 (N_8032,N_7232,N_6597);
and U8033 (N_8033,N_7404,N_6930);
or U8034 (N_8034,N_6622,N_5636);
or U8035 (N_8035,N_5655,N_6604);
nand U8036 (N_8036,N_6988,N_7267);
nand U8037 (N_8037,N_6821,N_7253);
nor U8038 (N_8038,N_6331,N_5844);
nor U8039 (N_8039,N_5320,N_6015);
nand U8040 (N_8040,N_6918,N_7023);
xnor U8041 (N_8041,N_6501,N_5100);
or U8042 (N_8042,N_5709,N_6141);
or U8043 (N_8043,N_5596,N_6436);
or U8044 (N_8044,N_6834,N_5796);
nand U8045 (N_8045,N_7087,N_7070);
xnor U8046 (N_8046,N_5326,N_6051);
nor U8047 (N_8047,N_7158,N_6636);
or U8048 (N_8048,N_7139,N_5423);
or U8049 (N_8049,N_6367,N_7153);
nand U8050 (N_8050,N_6696,N_6848);
or U8051 (N_8051,N_5748,N_5336);
and U8052 (N_8052,N_5020,N_5218);
or U8053 (N_8053,N_7423,N_5691);
nand U8054 (N_8054,N_5121,N_5378);
nor U8055 (N_8055,N_7272,N_7459);
or U8056 (N_8056,N_6170,N_5277);
or U8057 (N_8057,N_6983,N_6568);
nor U8058 (N_8058,N_5835,N_6828);
and U8059 (N_8059,N_6116,N_6229);
nor U8060 (N_8060,N_6518,N_6114);
and U8061 (N_8061,N_6072,N_6716);
nand U8062 (N_8062,N_5261,N_7325);
nor U8063 (N_8063,N_5211,N_7074);
or U8064 (N_8064,N_5734,N_6800);
and U8065 (N_8065,N_5619,N_5249);
nor U8066 (N_8066,N_6008,N_5182);
nor U8067 (N_8067,N_5587,N_6046);
or U8068 (N_8068,N_5299,N_6965);
and U8069 (N_8069,N_6082,N_6120);
and U8070 (N_8070,N_6438,N_7456);
nor U8071 (N_8071,N_5306,N_5644);
or U8072 (N_8072,N_5648,N_7312);
nor U8073 (N_8073,N_6524,N_6252);
nor U8074 (N_8074,N_6034,N_7317);
nand U8075 (N_8075,N_6902,N_6736);
nand U8076 (N_8076,N_6202,N_7007);
nor U8077 (N_8077,N_6333,N_6615);
and U8078 (N_8078,N_6400,N_6327);
nand U8079 (N_8079,N_5616,N_7077);
nor U8080 (N_8080,N_5005,N_5614);
nand U8081 (N_8081,N_6390,N_7265);
nand U8082 (N_8082,N_5180,N_6183);
or U8083 (N_8083,N_6753,N_5654);
nand U8084 (N_8084,N_6211,N_5640);
nor U8085 (N_8085,N_5130,N_7015);
and U8086 (N_8086,N_6432,N_5229);
nor U8087 (N_8087,N_5050,N_6363);
nand U8088 (N_8088,N_6483,N_5598);
or U8089 (N_8089,N_7447,N_6115);
nor U8090 (N_8090,N_6779,N_6868);
nor U8091 (N_8091,N_6869,N_6458);
or U8092 (N_8092,N_5166,N_6950);
or U8093 (N_8093,N_6101,N_7091);
and U8094 (N_8094,N_6969,N_5549);
or U8095 (N_8095,N_7244,N_7328);
or U8096 (N_8096,N_5908,N_5605);
and U8097 (N_8097,N_5833,N_6683);
or U8098 (N_8098,N_6731,N_7251);
or U8099 (N_8099,N_6577,N_5301);
nor U8100 (N_8100,N_5573,N_7216);
or U8101 (N_8101,N_5707,N_5925);
nor U8102 (N_8102,N_5150,N_5991);
nor U8103 (N_8103,N_6570,N_5199);
and U8104 (N_8104,N_6485,N_7482);
and U8105 (N_8105,N_6504,N_5381);
nor U8106 (N_8106,N_5329,N_6300);
or U8107 (N_8107,N_6098,N_5312);
nor U8108 (N_8108,N_5343,N_6240);
nand U8109 (N_8109,N_5615,N_6733);
or U8110 (N_8110,N_5827,N_5969);
nand U8111 (N_8111,N_6172,N_6398);
nand U8112 (N_8112,N_7155,N_7379);
and U8113 (N_8113,N_7255,N_6527);
nor U8114 (N_8114,N_6908,N_7365);
or U8115 (N_8115,N_6411,N_5532);
or U8116 (N_8116,N_7341,N_7279);
nor U8117 (N_8117,N_5251,N_6370);
and U8118 (N_8118,N_5890,N_6885);
nand U8119 (N_8119,N_6103,N_7280);
nor U8120 (N_8120,N_5292,N_5872);
nand U8121 (N_8121,N_5762,N_6168);
nor U8122 (N_8122,N_6010,N_5162);
and U8123 (N_8123,N_7213,N_6045);
or U8124 (N_8124,N_6195,N_6502);
nor U8125 (N_8125,N_7047,N_6480);
nor U8126 (N_8126,N_6373,N_5117);
or U8127 (N_8127,N_5310,N_7310);
or U8128 (N_8128,N_7214,N_7000);
and U8129 (N_8129,N_6841,N_6909);
and U8130 (N_8130,N_5913,N_5879);
nand U8131 (N_8131,N_6012,N_7330);
nor U8132 (N_8132,N_5857,N_5864);
nor U8133 (N_8133,N_5256,N_5286);
nand U8134 (N_8134,N_6248,N_5101);
nor U8135 (N_8135,N_6118,N_5639);
nor U8136 (N_8136,N_5688,N_7321);
nand U8137 (N_8137,N_7102,N_5807);
or U8138 (N_8138,N_5612,N_6740);
and U8139 (N_8139,N_5490,N_5321);
nand U8140 (N_8140,N_5322,N_7042);
and U8141 (N_8141,N_6618,N_7307);
or U8142 (N_8142,N_6849,N_6213);
nand U8143 (N_8143,N_6799,N_6375);
and U8144 (N_8144,N_5325,N_5148);
or U8145 (N_8145,N_6662,N_5171);
nand U8146 (N_8146,N_5102,N_6296);
and U8147 (N_8147,N_7084,N_5540);
and U8148 (N_8148,N_6939,N_5070);
nor U8149 (N_8149,N_6005,N_7235);
nor U8150 (N_8150,N_5680,N_7004);
and U8151 (N_8151,N_6276,N_6207);
nor U8152 (N_8152,N_6830,N_5942);
nand U8153 (N_8153,N_6493,N_5109);
nand U8154 (N_8154,N_6594,N_5885);
nor U8155 (N_8155,N_6440,N_7161);
or U8156 (N_8156,N_6558,N_5651);
and U8157 (N_8157,N_5949,N_7270);
or U8158 (N_8158,N_6132,N_6112);
nor U8159 (N_8159,N_7443,N_6911);
or U8160 (N_8160,N_5676,N_6685);
or U8161 (N_8161,N_7429,N_6083);
or U8162 (N_8162,N_5369,N_6592);
nand U8163 (N_8163,N_5091,N_5398);
or U8164 (N_8164,N_5311,N_5295);
nor U8165 (N_8165,N_5584,N_7002);
or U8166 (N_8166,N_6707,N_5751);
and U8167 (N_8167,N_5620,N_7112);
or U8168 (N_8168,N_6792,N_7446);
or U8169 (N_8169,N_6461,N_5904);
and U8170 (N_8170,N_5666,N_5678);
nor U8171 (N_8171,N_6538,N_5254);
and U8172 (N_8172,N_7115,N_5475);
and U8173 (N_8173,N_6874,N_5402);
nand U8174 (N_8174,N_6054,N_6852);
or U8175 (N_8175,N_6727,N_7064);
and U8176 (N_8176,N_6959,N_5282);
nor U8177 (N_8177,N_7257,N_5045);
and U8178 (N_8178,N_6184,N_5511);
nor U8179 (N_8179,N_6937,N_5272);
nor U8180 (N_8180,N_5450,N_6135);
nor U8181 (N_8181,N_5047,N_5663);
nor U8182 (N_8182,N_6341,N_6070);
and U8183 (N_8183,N_6575,N_6024);
xor U8184 (N_8184,N_6920,N_6235);
or U8185 (N_8185,N_5087,N_5553);
and U8186 (N_8186,N_5681,N_6658);
or U8187 (N_8187,N_6536,N_5370);
nor U8188 (N_8188,N_5994,N_6385);
nand U8189 (N_8189,N_7457,N_7052);
and U8190 (N_8190,N_5603,N_6187);
nor U8191 (N_8191,N_6409,N_5471);
and U8192 (N_8192,N_5088,N_5985);
nand U8193 (N_8193,N_6297,N_6839);
or U8194 (N_8194,N_6301,N_6859);
nor U8195 (N_8195,N_5951,N_6381);
or U8196 (N_8196,N_5519,N_7035);
nor U8197 (N_8197,N_6640,N_6729);
or U8198 (N_8198,N_5901,N_7349);
nor U8199 (N_8199,N_7184,N_7080);
nand U8200 (N_8200,N_6945,N_5075);
or U8201 (N_8201,N_6427,N_5232);
nor U8202 (N_8202,N_7086,N_6316);
and U8203 (N_8203,N_6802,N_6217);
nor U8204 (N_8204,N_5721,N_6639);
nand U8205 (N_8205,N_6999,N_5906);
and U8206 (N_8206,N_5738,N_6602);
nand U8207 (N_8207,N_5307,N_6542);
or U8208 (N_8208,N_6245,N_7152);
and U8209 (N_8209,N_5479,N_5371);
nor U8210 (N_8210,N_6760,N_6997);
nor U8211 (N_8211,N_5698,N_5448);
nand U8212 (N_8212,N_5517,N_6888);
nand U8213 (N_8213,N_5462,N_6847);
or U8214 (N_8214,N_7393,N_5665);
or U8215 (N_8215,N_5805,N_6452);
and U8216 (N_8216,N_5779,N_7179);
nor U8217 (N_8217,N_6055,N_5353);
nor U8218 (N_8218,N_6149,N_5442);
nor U8219 (N_8219,N_5143,N_5484);
nand U8220 (N_8220,N_5114,N_5297);
and U8221 (N_8221,N_6430,N_5941);
nor U8222 (N_8222,N_6644,N_5576);
or U8223 (N_8223,N_5443,N_5409);
nand U8224 (N_8224,N_5201,N_7194);
nand U8225 (N_8225,N_7263,N_6925);
and U8226 (N_8226,N_5588,N_7165);
and U8227 (N_8227,N_5493,N_6420);
and U8228 (N_8228,N_6748,N_7005);
nand U8229 (N_8229,N_6236,N_7498);
and U8230 (N_8230,N_5851,N_7200);
and U8231 (N_8231,N_7486,N_6460);
nand U8232 (N_8232,N_6257,N_6456);
or U8233 (N_8233,N_6352,N_5915);
nor U8234 (N_8234,N_6362,N_5524);
xor U8235 (N_8235,N_6446,N_7348);
and U8236 (N_8236,N_5094,N_6428);
nand U8237 (N_8237,N_5818,N_6808);
nand U8238 (N_8238,N_5571,N_7096);
xnor U8239 (N_8239,N_6936,N_6755);
nor U8240 (N_8240,N_6660,N_5161);
and U8241 (N_8241,N_6481,N_5278);
nor U8242 (N_8242,N_5305,N_6626);
nor U8243 (N_8243,N_6324,N_5043);
nor U8244 (N_8244,N_7053,N_5038);
or U8245 (N_8245,N_6656,N_6817);
or U8246 (N_8246,N_6865,N_5255);
nand U8247 (N_8247,N_7020,N_6329);
nand U8248 (N_8248,N_6337,N_7294);
nand U8249 (N_8249,N_6462,N_7143);
nor U8250 (N_8250,N_6601,N_6496);
nand U8251 (N_8251,N_5743,N_6843);
and U8252 (N_8252,N_6807,N_5808);
nor U8253 (N_8253,N_5705,N_7339);
and U8254 (N_8254,N_7386,N_7217);
and U8255 (N_8255,N_5752,N_6862);
nand U8256 (N_8256,N_5056,N_6105);
nor U8257 (N_8257,N_5332,N_5428);
nor U8258 (N_8258,N_6177,N_5594);
nor U8259 (N_8259,N_6708,N_7420);
and U8260 (N_8260,N_6719,N_5522);
nand U8261 (N_8261,N_6938,N_6772);
nand U8262 (N_8262,N_5737,N_6850);
nor U8263 (N_8263,N_6369,N_6258);
and U8264 (N_8264,N_6201,N_5803);
nor U8265 (N_8265,N_5391,N_5124);
or U8266 (N_8266,N_7103,N_5804);
and U8267 (N_8267,N_6402,N_5407);
nor U8268 (N_8268,N_7433,N_7432);
nor U8269 (N_8269,N_7426,N_7220);
nand U8270 (N_8270,N_6425,N_5158);
and U8271 (N_8271,N_5035,N_5226);
nand U8272 (N_8272,N_6543,N_6439);
nor U8273 (N_8273,N_5990,N_5008);
or U8274 (N_8274,N_5547,N_6894);
nand U8275 (N_8275,N_6966,N_6876);
or U8276 (N_8276,N_6788,N_5810);
nor U8277 (N_8277,N_5896,N_6199);
nand U8278 (N_8278,N_5293,N_6567);
nor U8279 (N_8279,N_6268,N_5108);
nor U8280 (N_8280,N_7332,N_5887);
and U8281 (N_8281,N_5403,N_5195);
nand U8282 (N_8282,N_6758,N_7181);
nand U8283 (N_8283,N_6039,N_5781);
nor U8284 (N_8284,N_6419,N_6724);
nand U8285 (N_8285,N_6153,N_6705);
nand U8286 (N_8286,N_6164,N_5822);
and U8287 (N_8287,N_5436,N_5669);
nand U8288 (N_8288,N_6416,N_5505);
nand U8289 (N_8289,N_6057,N_7154);
nand U8290 (N_8290,N_5989,N_6021);
nor U8291 (N_8291,N_6294,N_5735);
or U8292 (N_8292,N_6166,N_5197);
nor U8293 (N_8293,N_5635,N_7032);
or U8294 (N_8294,N_5973,N_5811);
and U8295 (N_8295,N_5793,N_5433);
nor U8296 (N_8296,N_6780,N_7173);
and U8297 (N_8297,N_6654,N_7323);
nor U8298 (N_8298,N_5924,N_5155);
nor U8299 (N_8299,N_7240,N_6711);
nand U8300 (N_8300,N_7038,N_5042);
nor U8301 (N_8301,N_5337,N_5950);
nand U8302 (N_8302,N_6389,N_5472);
and U8303 (N_8303,N_6364,N_6061);
and U8304 (N_8304,N_7396,N_7302);
and U8305 (N_8305,N_7416,N_6286);
and U8306 (N_8306,N_6102,N_5394);
nand U8307 (N_8307,N_5494,N_6122);
or U8308 (N_8308,N_7147,N_5686);
or U8309 (N_8309,N_5860,N_6181);
nor U8310 (N_8310,N_5777,N_6063);
nand U8311 (N_8311,N_6078,N_7422);
nor U8312 (N_8312,N_6559,N_7130);
nand U8313 (N_8313,N_6277,N_7408);
and U8314 (N_8314,N_5280,N_6080);
and U8315 (N_8315,N_5412,N_5995);
nand U8316 (N_8316,N_6970,N_6686);
nor U8317 (N_8317,N_7157,N_5816);
nor U8318 (N_8318,N_5625,N_6670);
or U8319 (N_8319,N_6304,N_6954);
nand U8320 (N_8320,N_5930,N_6479);
or U8321 (N_8321,N_7301,N_7359);
xor U8322 (N_8322,N_6827,N_6194);
nor U8323 (N_8323,N_6007,N_6314);
nand U8324 (N_8324,N_6107,N_7046);
nor U8325 (N_8325,N_5137,N_5473);
nor U8326 (N_8326,N_7451,N_7376);
nand U8327 (N_8327,N_5247,N_7300);
nor U8328 (N_8328,N_5695,N_5029);
nand U8329 (N_8329,N_5375,N_5283);
and U8330 (N_8330,N_5149,N_6081);
nor U8331 (N_8331,N_6987,N_5303);
nand U8332 (N_8332,N_6721,N_6584);
or U8333 (N_8333,N_6650,N_5775);
nand U8334 (N_8334,N_6169,N_6963);
or U8335 (N_8335,N_6328,N_5823);
or U8336 (N_8336,N_7191,N_6804);
nor U8337 (N_8337,N_5641,N_6671);
or U8338 (N_8338,N_7187,N_6738);
nand U8339 (N_8339,N_5454,N_6793);
nor U8340 (N_8340,N_7355,N_6437);
nor U8341 (N_8341,N_7461,N_5839);
nor U8342 (N_8342,N_6028,N_5333);
nand U8343 (N_8343,N_6180,N_5499);
nand U8344 (N_8344,N_5773,N_5711);
and U8345 (N_8345,N_6981,N_5294);
nor U8346 (N_8346,N_7134,N_6142);
nand U8347 (N_8347,N_5276,N_5634);
nor U8348 (N_8348,N_6528,N_5821);
nor U8349 (N_8349,N_5983,N_6872);
or U8350 (N_8350,N_7072,N_5061);
nor U8351 (N_8351,N_5945,N_6247);
or U8352 (N_8352,N_6521,N_5486);
nor U8353 (N_8353,N_5592,N_5007);
and U8354 (N_8354,N_6193,N_6856);
nand U8355 (N_8355,N_6659,N_7378);
nand U8356 (N_8356,N_6898,N_5604);
and U8357 (N_8357,N_6704,N_7258);
nand U8358 (N_8358,N_6386,N_6330);
and U8359 (N_8359,N_5555,N_7309);
nor U8360 (N_8360,N_7033,N_7062);
nand U8361 (N_8361,N_7289,N_7346);
nor U8362 (N_8362,N_7208,N_6961);
and U8363 (N_8363,N_5624,N_7297);
nand U8364 (N_8364,N_6464,N_5968);
or U8365 (N_8365,N_5838,N_6410);
nand U8366 (N_8366,N_6104,N_6397);
or U8367 (N_8367,N_6074,N_5400);
or U8368 (N_8368,N_7314,N_5846);
nor U8369 (N_8369,N_7311,N_6717);
nand U8370 (N_8370,N_5236,N_5157);
or U8371 (N_8371,N_5546,N_6516);
nor U8372 (N_8372,N_5628,N_5331);
nor U8373 (N_8373,N_6006,N_6143);
nor U8374 (N_8374,N_5176,N_6871);
nand U8375 (N_8375,N_5567,N_6652);
nand U8376 (N_8376,N_6160,N_7029);
nor U8377 (N_8377,N_5589,N_5905);
or U8378 (N_8378,N_7094,N_6933);
nand U8379 (N_8379,N_5740,N_6648);
nand U8380 (N_8380,N_7085,N_6900);
nor U8381 (N_8381,N_6924,N_7028);
nor U8382 (N_8382,N_5013,N_6914);
or U8383 (N_8383,N_6401,N_5926);
nand U8384 (N_8384,N_5049,N_7196);
nor U8385 (N_8385,N_5677,N_5152);
or U8386 (N_8386,N_7481,N_6833);
and U8387 (N_8387,N_7371,N_5151);
nand U8388 (N_8388,N_5122,N_7071);
nand U8389 (N_8389,N_7246,N_5749);
and U8390 (N_8390,N_7436,N_5753);
and U8391 (N_8391,N_5929,N_6709);
nand U8392 (N_8392,N_7467,N_5911);
nor U8393 (N_8393,N_6929,N_5858);
nor U8394 (N_8394,N_7239,N_7250);
nand U8395 (N_8395,N_5881,N_6009);
and U8396 (N_8396,N_6290,N_6133);
nor U8397 (N_8397,N_5491,N_7242);
or U8398 (N_8398,N_5809,N_7398);
or U8399 (N_8399,N_7455,N_6086);
nand U8400 (N_8400,N_7405,N_5712);
or U8401 (N_8401,N_6732,N_6215);
or U8402 (N_8402,N_5210,N_6553);
and U8403 (N_8403,N_6562,N_6747);
and U8404 (N_8404,N_6907,N_7287);
nand U8405 (N_8405,N_7078,N_7148);
nand U8406 (N_8406,N_6310,N_6844);
or U8407 (N_8407,N_6038,N_7331);
nand U8408 (N_8408,N_6026,N_5776);
nand U8409 (N_8409,N_5178,N_7285);
nand U8410 (N_8410,N_5267,N_6510);
and U8411 (N_8411,N_5986,N_6892);
nand U8412 (N_8412,N_6196,N_6272);
and U8413 (N_8413,N_5689,N_7090);
and U8414 (N_8414,N_6259,N_7168);
and U8415 (N_8415,N_7100,N_5745);
or U8416 (N_8416,N_5645,N_5848);
and U8417 (N_8417,N_7450,N_5474);
nand U8418 (N_8418,N_5488,N_6058);
or U8419 (N_8419,N_5366,N_7352);
and U8420 (N_8420,N_6476,N_6899);
or U8421 (N_8421,N_5451,N_6254);
and U8422 (N_8422,N_5181,N_7188);
nand U8423 (N_8423,N_5928,N_7465);
nor U8424 (N_8424,N_6148,N_5023);
nand U8425 (N_8425,N_5548,N_7428);
or U8426 (N_8426,N_5907,N_6687);
or U8427 (N_8427,N_6282,N_5156);
or U8428 (N_8428,N_6541,N_6161);
and U8429 (N_8429,N_5984,N_7286);
nand U8430 (N_8430,N_5910,N_5221);
nor U8431 (N_8431,N_5095,N_5172);
nand U8432 (N_8432,N_5065,N_5633);
and U8433 (N_8433,N_6979,N_5759);
nand U8434 (N_8434,N_5467,N_5902);
and U8435 (N_8435,N_7370,N_5379);
nor U8436 (N_8436,N_6690,N_7385);
nor U8437 (N_8437,N_7122,N_6934);
or U8438 (N_8438,N_5416,N_7375);
nor U8439 (N_8439,N_6003,N_6505);
nand U8440 (N_8440,N_5081,N_5716);
and U8441 (N_8441,N_6916,N_7132);
or U8442 (N_8442,N_7304,N_5074);
nor U8443 (N_8443,N_6897,N_6125);
or U8444 (N_8444,N_7254,N_7269);
or U8445 (N_8445,N_7444,N_5876);
nand U8446 (N_8446,N_6944,N_7228);
and U8447 (N_8447,N_5602,N_5938);
nor U8448 (N_8448,N_6810,N_5981);
nor U8449 (N_8449,N_6291,N_5866);
nand U8450 (N_8450,N_5960,N_7075);
or U8451 (N_8451,N_5086,N_5160);
nor U8452 (N_8452,N_7106,N_5853);
xor U8453 (N_8453,N_6803,N_5235);
and U8454 (N_8454,N_5536,N_6471);
and U8455 (N_8455,N_5884,N_6218);
or U8456 (N_8456,N_6557,N_7462);
nor U8457 (N_8457,N_6973,N_7121);
and U8458 (N_8458,N_5697,N_6200);
nor U8459 (N_8459,N_5658,N_6138);
or U8460 (N_8460,N_5327,N_5376);
nand U8461 (N_8461,N_5574,N_6032);
or U8462 (N_8462,N_6761,N_5372);
or U8463 (N_8463,N_5129,N_6976);
and U8464 (N_8464,N_6243,N_6548);
nor U8465 (N_8465,N_5233,N_7271);
and U8466 (N_8466,N_7140,N_5456);
and U8467 (N_8467,N_6519,N_7142);
nand U8468 (N_8468,N_6680,N_6797);
nand U8469 (N_8469,N_6785,N_5318);
and U8470 (N_8470,N_7318,N_6404);
and U8471 (N_8471,N_6896,N_5003);
and U8472 (N_8472,N_6097,N_6192);
and U8473 (N_8473,N_6069,N_5271);
nand U8474 (N_8474,N_6156,N_5886);
nand U8475 (N_8475,N_6197,N_6836);
or U8476 (N_8476,N_6910,N_5179);
nand U8477 (N_8477,N_6585,N_6448);
xnor U8478 (N_8478,N_6270,N_5389);
nor U8479 (N_8479,N_5385,N_6569);
nand U8480 (N_8480,N_5314,N_5739);
nand U8481 (N_8481,N_7149,N_5538);
and U8482 (N_8482,N_6463,N_6292);
nand U8483 (N_8483,N_5601,N_6667);
and U8484 (N_8484,N_5627,N_5079);
and U8485 (N_8485,N_5814,N_6701);
nand U8486 (N_8486,N_5093,N_6253);
or U8487 (N_8487,N_5802,N_6943);
or U8488 (N_8488,N_7319,N_5273);
and U8489 (N_8489,N_5714,N_6421);
nor U8490 (N_8490,N_6886,N_6508);
and U8491 (N_8491,N_7329,N_6840);
nor U8492 (N_8492,N_6664,N_6980);
nor U8493 (N_8493,N_5228,N_6472);
nor U8494 (N_8494,N_7008,N_5795);
nor U8495 (N_8495,N_6773,N_7259);
nand U8496 (N_8496,N_6702,N_5987);
nor U8497 (N_8497,N_6579,N_5733);
and U8498 (N_8498,N_6041,N_5154);
and U8499 (N_8499,N_5354,N_5173);
nor U8500 (N_8500,N_6771,N_5365);
and U8501 (N_8501,N_7107,N_6895);
or U8502 (N_8502,N_5568,N_6509);
nand U8503 (N_8503,N_5967,N_6406);
nand U8504 (N_8504,N_5939,N_5971);
nand U8505 (N_8505,N_5039,N_5997);
or U8506 (N_8506,N_6681,N_7363);
or U8507 (N_8507,N_5916,N_6155);
or U8508 (N_8508,N_6431,N_6099);
and U8509 (N_8509,N_6968,N_6377);
or U8510 (N_8510,N_7227,N_6459);
nor U8511 (N_8511,N_7058,N_6782);
and U8512 (N_8512,N_6349,N_7125);
and U8513 (N_8513,N_5447,N_7230);
nor U8514 (N_8514,N_6342,N_6879);
nand U8515 (N_8515,N_5979,N_6674);
or U8516 (N_8516,N_6586,N_6233);
nor U8517 (N_8517,N_5690,N_6450);
nor U8518 (N_8518,N_5241,N_7170);
nand U8519 (N_8519,N_5194,N_5897);
and U8520 (N_8520,N_6877,N_6820);
and U8521 (N_8521,N_5350,N_5032);
nand U8522 (N_8522,N_6560,N_6293);
nor U8523 (N_8523,N_5468,N_5253);
nand U8524 (N_8524,N_7324,N_5208);
nor U8525 (N_8525,N_5335,N_5057);
and U8526 (N_8526,N_6688,N_7357);
nor U8527 (N_8527,N_6623,N_6957);
nand U8528 (N_8528,N_5509,N_5537);
and U8529 (N_8529,N_7037,N_6157);
nand U8530 (N_8530,N_6056,N_5338);
or U8531 (N_8531,N_5722,N_6473);
and U8532 (N_8532,N_7394,N_6378);
or U8533 (N_8533,N_6035,N_6668);
and U8534 (N_8534,N_5508,N_5862);
nor U8535 (N_8535,N_7430,N_7185);
nor U8536 (N_8536,N_5223,N_6299);
nor U8537 (N_8537,N_6131,N_5684);
nor U8538 (N_8538,N_7464,N_7298);
and U8539 (N_8539,N_7316,N_5642);
or U8540 (N_8540,N_6089,N_6288);
or U8541 (N_8541,N_7402,N_5266);
nor U8542 (N_8542,N_5498,N_6960);
or U8543 (N_8543,N_6186,N_5520);
and U8544 (N_8544,N_7099,N_5923);
and U8545 (N_8545,N_7016,N_5590);
and U8546 (N_8546,N_6339,N_7127);
nor U8547 (N_8547,N_6382,N_5593);
and U8548 (N_8548,N_6904,N_5186);
or U8549 (N_8549,N_5418,N_6415);
nand U8550 (N_8550,N_5460,N_6109);
and U8551 (N_8551,N_5021,N_7207);
nand U8552 (N_8552,N_7274,N_7088);
and U8553 (N_8553,N_6809,N_5440);
and U8554 (N_8554,N_6846,N_5525);
and U8555 (N_8555,N_5832,N_5591);
nor U8556 (N_8556,N_5704,N_5873);
nand U8557 (N_8557,N_6442,N_6750);
or U8558 (N_8558,N_5435,N_7474);
or U8559 (N_8559,N_6526,N_5387);
nand U8560 (N_8560,N_5187,N_5084);
nor U8561 (N_8561,N_5672,N_6206);
or U8562 (N_8562,N_6457,N_5597);
or U8563 (N_8563,N_7412,N_5064);
nor U8564 (N_8564,N_6351,N_6470);
and U8565 (N_8565,N_6242,N_6066);
nand U8566 (N_8566,N_5386,N_6754);
or U8567 (N_8567,N_6522,N_5265);
or U8568 (N_8568,N_5118,N_6165);
or U8569 (N_8569,N_5646,N_5892);
and U8570 (N_8570,N_6972,N_7010);
nor U8571 (N_8571,N_5895,N_5274);
and U8572 (N_8572,N_6990,N_5395);
or U8573 (N_8573,N_5554,N_7480);
xnor U8574 (N_8574,N_6000,N_6075);
nand U8575 (N_8575,N_7024,N_7031);
xnor U8576 (N_8576,N_6752,N_5944);
or U8577 (N_8577,N_5257,N_5940);
xnor U8578 (N_8578,N_7061,N_5719);
nor U8579 (N_8579,N_5660,N_6549);
or U8580 (N_8580,N_5682,N_5784);
nor U8581 (N_8581,N_6274,N_5125);
or U8582 (N_8582,N_5355,N_5702);
nand U8583 (N_8583,N_5055,N_5742);
nand U8584 (N_8584,N_5673,N_7387);
nand U8585 (N_8585,N_5290,N_5607);
and U8586 (N_8586,N_7104,N_5027);
nand U8587 (N_8587,N_6693,N_6354);
nor U8588 (N_8588,N_6088,N_7145);
nand U8589 (N_8589,N_5710,N_5900);
or U8590 (N_8590,N_7276,N_6815);
and U8591 (N_8591,N_6759,N_6795);
and U8592 (N_8592,N_6309,N_5377);
xnor U8593 (N_8593,N_7131,N_5975);
nand U8594 (N_8594,N_5541,N_5205);
nand U8595 (N_8595,N_7337,N_6488);
or U8596 (N_8596,N_5728,N_7176);
nand U8597 (N_8597,N_5163,N_5670);
or U8598 (N_8598,N_6525,N_6498);
and U8599 (N_8599,N_7083,N_6128);
or U8600 (N_8600,N_5217,N_6188);
or U8601 (N_8601,N_6825,N_6737);
nor U8602 (N_8602,N_6713,N_5687);
or U8603 (N_8603,N_7340,N_6714);
nand U8604 (N_8604,N_5580,N_7374);
nand U8605 (N_8605,N_5461,N_6511);
and U8606 (N_8606,N_5080,N_7098);
and U8607 (N_8607,N_5552,N_5831);
nor U8608 (N_8608,N_5031,N_7136);
and U8609 (N_8609,N_5465,N_6768);
nand U8610 (N_8610,N_6059,N_5144);
and U8611 (N_8611,N_7222,N_6582);
and U8612 (N_8612,N_6490,N_5726);
nor U8613 (N_8613,N_5106,N_6947);
nor U8614 (N_8614,N_6241,N_5245);
and U8615 (N_8615,N_6002,N_7320);
and U8616 (N_8616,N_6581,N_6049);
nor U8617 (N_8617,N_6806,N_5457);
and U8618 (N_8618,N_6495,N_5544);
nand U8619 (N_8619,N_6787,N_6497);
or U8620 (N_8620,N_6037,N_6743);
nor U8621 (N_8621,N_6741,N_7493);
or U8622 (N_8622,N_6786,N_5134);
or U8623 (N_8623,N_6068,N_6529);
nand U8624 (N_8624,N_6634,N_7025);
and U8625 (N_8625,N_5649,N_6147);
nor U8626 (N_8626,N_6931,N_6320);
nand U8627 (N_8627,N_7203,N_7056);
or U8628 (N_8628,N_6424,N_6672);
xor U8629 (N_8629,N_6777,N_6305);
or U8630 (N_8630,N_5430,N_6619);
or U8631 (N_8631,N_6140,N_5268);
nor U8632 (N_8632,N_6119,N_5004);
and U8633 (N_8633,N_5718,N_5650);
and U8634 (N_8634,N_6712,N_6150);
nand U8635 (N_8635,N_6262,N_6974);
or U8636 (N_8636,N_7466,N_7092);
or U8637 (N_8637,N_6606,N_6922);
or U8638 (N_8638,N_7470,N_5518);
or U8639 (N_8639,N_5362,N_6047);
or U8640 (N_8640,N_6631,N_5708);
or U8641 (N_8641,N_7475,N_6513);
and U8642 (N_8642,N_5856,N_5512);
and U8643 (N_8643,N_5729,N_5200);
nor U8644 (N_8644,N_6996,N_6062);
and U8645 (N_8645,N_6677,N_6520);
or U8646 (N_8646,N_6726,N_5700);
nand U8647 (N_8647,N_6676,N_6469);
or U8648 (N_8648,N_5072,N_5744);
and U8649 (N_8649,N_6998,N_5980);
and U8650 (N_8650,N_7068,N_6280);
nor U8651 (N_8651,N_7110,N_5629);
nand U8652 (N_8652,N_5766,N_6883);
or U8653 (N_8653,N_7479,N_6625);
or U8654 (N_8654,N_6226,N_5153);
nor U8655 (N_8655,N_5502,N_7059);
or U8656 (N_8656,N_6565,N_5242);
nand U8657 (N_8657,N_7097,N_6679);
nor U8658 (N_8658,N_6655,N_5077);
nor U8659 (N_8659,N_6781,N_5470);
nor U8660 (N_8660,N_7169,N_5390);
nor U8661 (N_8661,N_6060,N_6638);
and U8662 (N_8662,N_6167,N_5761);
nor U8663 (N_8663,N_7473,N_6853);
nor U8664 (N_8664,N_5105,N_6540);
or U8665 (N_8665,N_5419,N_5531);
and U8666 (N_8666,N_5126,N_7322);
nor U8667 (N_8667,N_5632,N_6040);
and U8668 (N_8668,N_6004,N_5308);
nand U8669 (N_8669,N_5434,N_6151);
and U8670 (N_8670,N_5224,N_7198);
and U8671 (N_8671,N_5206,N_7381);
nand U8672 (N_8672,N_5883,N_6629);
nand U8673 (N_8673,N_6612,N_5870);
and U8674 (N_8674,N_7095,N_6573);
or U8675 (N_8675,N_5561,N_6561);
or U8676 (N_8676,N_6423,N_5693);
nand U8677 (N_8677,N_6073,N_6866);
nor U8678 (N_8678,N_6951,N_6322);
nor U8679 (N_8679,N_6319,N_5340);
nand U8680 (N_8680,N_6326,N_5011);
nor U8681 (N_8681,N_6361,N_6344);
nand U8682 (N_8682,N_7209,N_7089);
nand U8683 (N_8683,N_6295,N_6867);
nor U8684 (N_8684,N_7219,N_6065);
or U8685 (N_8685,N_6368,N_6018);
or U8686 (N_8686,N_6176,N_5583);
and U8687 (N_8687,N_6609,N_5919);
nand U8688 (N_8688,N_6798,N_6231);
and U8689 (N_8689,N_5898,N_6661);
and U8690 (N_8690,N_5207,N_6379);
nand U8691 (N_8691,N_5786,N_5675);
nand U8692 (N_8692,N_6975,N_6392);
nor U8693 (N_8693,N_5974,N_5970);
nor U8694 (N_8694,N_6955,N_5246);
and U8695 (N_8695,N_6484,N_5724);
nand U8696 (N_8696,N_5415,N_5893);
and U8697 (N_8697,N_5836,N_5868);
and U8698 (N_8698,N_6347,N_7453);
and U8699 (N_8699,N_5240,N_7382);
and U8700 (N_8700,N_6336,N_6185);
nor U8701 (N_8701,N_5196,N_6094);
nor U8702 (N_8702,N_5222,N_6814);
nand U8703 (N_8703,N_5771,N_6861);
and U8704 (N_8704,N_6552,N_7288);
and U8705 (N_8705,N_5281,N_5098);
nor U8706 (N_8706,N_7460,N_5778);
and U8707 (N_8707,N_7001,N_5275);
and U8708 (N_8708,N_7225,N_5610);
or U8709 (N_8709,N_5339,N_6123);
xnor U8710 (N_8710,N_6237,N_7252);
or U8711 (N_8711,N_7391,N_6251);
nand U8712 (N_8712,N_5001,N_6730);
nor U8713 (N_8713,N_5875,N_7014);
or U8714 (N_8714,N_5825,N_5671);
nor U8715 (N_8715,N_5068,N_6993);
and U8716 (N_8716,N_5659,N_7437);
nand U8717 (N_8717,N_6455,N_5859);
and U8718 (N_8718,N_6697,N_6260);
and U8719 (N_8719,N_7189,N_7137);
and U8720 (N_8720,N_7171,N_5521);
or U8721 (N_8721,N_6598,N_5184);
and U8722 (N_8722,N_5912,N_7343);
nor U8723 (N_8723,N_6563,N_7006);
or U8724 (N_8724,N_7400,N_6267);
nor U8725 (N_8725,N_6599,N_6739);
nor U8726 (N_8726,N_5459,N_6356);
nor U8727 (N_8727,N_7488,N_7303);
nand U8728 (N_8728,N_7050,N_6873);
nand U8729 (N_8729,N_7040,N_5424);
nor U8730 (N_8730,N_7477,N_6136);
nand U8731 (N_8731,N_5750,N_6627);
or U8732 (N_8732,N_5785,N_5165);
nor U8733 (N_8733,N_6551,N_5414);
and U8734 (N_8734,N_6893,N_5046);
and U8735 (N_8735,N_6279,N_5664);
and U8736 (N_8736,N_7342,N_5092);
or U8737 (N_8737,N_6405,N_5798);
and U8738 (N_8738,N_5964,N_5764);
nor U8739 (N_8739,N_5260,N_5188);
and U8740 (N_8740,N_6822,N_5175);
nand U8741 (N_8741,N_6875,N_6695);
and U8742 (N_8742,N_5287,N_6113);
and U8743 (N_8743,N_6967,N_6550);
nand U8744 (N_8744,N_6506,N_6144);
and U8745 (N_8745,N_5067,N_5477);
or U8746 (N_8746,N_7472,N_5449);
or U8747 (N_8747,N_6689,N_6117);
nand U8748 (N_8748,N_5183,N_7344);
or U8749 (N_8749,N_5500,N_6384);
and U8750 (N_8750,N_5725,N_7449);
nand U8751 (N_8751,N_5665,N_6264);
nand U8752 (N_8752,N_7492,N_6288);
or U8753 (N_8753,N_5223,N_5913);
nand U8754 (N_8754,N_5847,N_5979);
and U8755 (N_8755,N_7282,N_6671);
and U8756 (N_8756,N_6367,N_7307);
nor U8757 (N_8757,N_5190,N_5756);
or U8758 (N_8758,N_6555,N_7301);
nor U8759 (N_8759,N_6285,N_6566);
nand U8760 (N_8760,N_6640,N_6868);
nor U8761 (N_8761,N_6158,N_5802);
nand U8762 (N_8762,N_6543,N_6150);
nor U8763 (N_8763,N_5990,N_5546);
or U8764 (N_8764,N_5054,N_7192);
nor U8765 (N_8765,N_6650,N_7093);
and U8766 (N_8766,N_7110,N_6758);
and U8767 (N_8767,N_7326,N_5172);
nand U8768 (N_8768,N_5707,N_5173);
nor U8769 (N_8769,N_6869,N_6461);
and U8770 (N_8770,N_6346,N_5675);
and U8771 (N_8771,N_6827,N_7199);
nor U8772 (N_8772,N_6935,N_7307);
nand U8773 (N_8773,N_6149,N_7137);
and U8774 (N_8774,N_7470,N_7184);
nor U8775 (N_8775,N_6416,N_5396);
and U8776 (N_8776,N_5136,N_5583);
nand U8777 (N_8777,N_5193,N_5155);
nor U8778 (N_8778,N_6037,N_6811);
nand U8779 (N_8779,N_6307,N_6952);
and U8780 (N_8780,N_7484,N_7014);
nand U8781 (N_8781,N_5340,N_7382);
or U8782 (N_8782,N_6031,N_6257);
or U8783 (N_8783,N_7295,N_5706);
nor U8784 (N_8784,N_5126,N_6987);
nand U8785 (N_8785,N_6885,N_5008);
nand U8786 (N_8786,N_6353,N_5857);
and U8787 (N_8787,N_5063,N_6487);
nand U8788 (N_8788,N_6115,N_6434);
or U8789 (N_8789,N_7426,N_5346);
and U8790 (N_8790,N_5745,N_6698);
and U8791 (N_8791,N_5759,N_5752);
and U8792 (N_8792,N_6089,N_6394);
and U8793 (N_8793,N_7043,N_7467);
nor U8794 (N_8794,N_6842,N_5226);
and U8795 (N_8795,N_5962,N_5535);
nor U8796 (N_8796,N_6185,N_6985);
nand U8797 (N_8797,N_5197,N_6903);
and U8798 (N_8798,N_5177,N_7272);
or U8799 (N_8799,N_5389,N_6028);
nor U8800 (N_8800,N_7399,N_5746);
nand U8801 (N_8801,N_5527,N_5095);
nor U8802 (N_8802,N_5522,N_6460);
nor U8803 (N_8803,N_6078,N_6235);
and U8804 (N_8804,N_5272,N_6071);
nor U8805 (N_8805,N_6751,N_6393);
or U8806 (N_8806,N_7173,N_7113);
nor U8807 (N_8807,N_6684,N_6416);
nor U8808 (N_8808,N_6595,N_5963);
and U8809 (N_8809,N_6757,N_5650);
nand U8810 (N_8810,N_6615,N_5064);
or U8811 (N_8811,N_5306,N_6662);
and U8812 (N_8812,N_6634,N_6315);
nor U8813 (N_8813,N_6657,N_7432);
nand U8814 (N_8814,N_6564,N_5857);
nor U8815 (N_8815,N_6767,N_5665);
nor U8816 (N_8816,N_7017,N_7094);
nor U8817 (N_8817,N_6547,N_6394);
nand U8818 (N_8818,N_6640,N_6153);
and U8819 (N_8819,N_7417,N_7469);
nand U8820 (N_8820,N_6809,N_7055);
and U8821 (N_8821,N_5234,N_6006);
and U8822 (N_8822,N_7188,N_5444);
nand U8823 (N_8823,N_6378,N_6214);
and U8824 (N_8824,N_5441,N_5449);
or U8825 (N_8825,N_5523,N_5472);
nand U8826 (N_8826,N_5072,N_6446);
and U8827 (N_8827,N_6288,N_5755);
nand U8828 (N_8828,N_5097,N_7195);
nand U8829 (N_8829,N_7160,N_7357);
nand U8830 (N_8830,N_5406,N_6215);
nor U8831 (N_8831,N_5522,N_5857);
nand U8832 (N_8832,N_7294,N_6419);
and U8833 (N_8833,N_6397,N_7250);
nor U8834 (N_8834,N_5600,N_6657);
or U8835 (N_8835,N_5320,N_6461);
nand U8836 (N_8836,N_6877,N_5109);
and U8837 (N_8837,N_6116,N_5869);
and U8838 (N_8838,N_5147,N_6763);
and U8839 (N_8839,N_5265,N_7021);
xnor U8840 (N_8840,N_5227,N_5212);
and U8841 (N_8841,N_5732,N_5356);
nor U8842 (N_8842,N_6119,N_6052);
and U8843 (N_8843,N_7371,N_6827);
nor U8844 (N_8844,N_5239,N_6547);
and U8845 (N_8845,N_5915,N_6863);
and U8846 (N_8846,N_5564,N_6434);
nor U8847 (N_8847,N_5672,N_6838);
and U8848 (N_8848,N_6047,N_5531);
or U8849 (N_8849,N_6229,N_7140);
and U8850 (N_8850,N_6795,N_5211);
and U8851 (N_8851,N_5122,N_6763);
nand U8852 (N_8852,N_7095,N_5933);
and U8853 (N_8853,N_5462,N_6767);
and U8854 (N_8854,N_5234,N_6050);
and U8855 (N_8855,N_5859,N_5954);
nand U8856 (N_8856,N_6122,N_5644);
or U8857 (N_8857,N_6039,N_6206);
or U8858 (N_8858,N_6348,N_5702);
and U8859 (N_8859,N_5505,N_5929);
and U8860 (N_8860,N_6318,N_6884);
or U8861 (N_8861,N_6809,N_6668);
nor U8862 (N_8862,N_7480,N_5787);
and U8863 (N_8863,N_6190,N_6802);
and U8864 (N_8864,N_6110,N_5552);
nor U8865 (N_8865,N_5015,N_6175);
nand U8866 (N_8866,N_7446,N_6898);
and U8867 (N_8867,N_5181,N_5025);
nor U8868 (N_8868,N_6870,N_6719);
or U8869 (N_8869,N_7352,N_6616);
or U8870 (N_8870,N_6337,N_7094);
or U8871 (N_8871,N_6206,N_6950);
nor U8872 (N_8872,N_6875,N_6056);
nand U8873 (N_8873,N_6147,N_5172);
and U8874 (N_8874,N_6379,N_7043);
or U8875 (N_8875,N_6031,N_6627);
nand U8876 (N_8876,N_5194,N_7023);
nand U8877 (N_8877,N_5058,N_6147);
and U8878 (N_8878,N_6336,N_6814);
nor U8879 (N_8879,N_6294,N_6694);
and U8880 (N_8880,N_5822,N_6863);
nand U8881 (N_8881,N_6062,N_5861);
nor U8882 (N_8882,N_7386,N_6629);
or U8883 (N_8883,N_7160,N_6285);
and U8884 (N_8884,N_5195,N_7407);
or U8885 (N_8885,N_6621,N_5288);
nor U8886 (N_8886,N_5141,N_7288);
and U8887 (N_8887,N_6529,N_7199);
nor U8888 (N_8888,N_7079,N_6866);
or U8889 (N_8889,N_5267,N_5927);
and U8890 (N_8890,N_5325,N_6648);
nor U8891 (N_8891,N_5210,N_5116);
or U8892 (N_8892,N_7009,N_6174);
nand U8893 (N_8893,N_5701,N_7041);
nand U8894 (N_8894,N_5928,N_7110);
and U8895 (N_8895,N_5099,N_5537);
or U8896 (N_8896,N_6086,N_7128);
nor U8897 (N_8897,N_6042,N_6912);
nand U8898 (N_8898,N_6145,N_7123);
nor U8899 (N_8899,N_7122,N_5572);
nand U8900 (N_8900,N_7152,N_6752);
or U8901 (N_8901,N_5147,N_6571);
nor U8902 (N_8902,N_7013,N_5183);
nand U8903 (N_8903,N_5159,N_5344);
or U8904 (N_8904,N_5017,N_6449);
nor U8905 (N_8905,N_6256,N_6900);
xnor U8906 (N_8906,N_7449,N_6033);
nand U8907 (N_8907,N_7385,N_6602);
nand U8908 (N_8908,N_7282,N_5910);
nor U8909 (N_8909,N_6479,N_6161);
or U8910 (N_8910,N_6016,N_5029);
or U8911 (N_8911,N_6561,N_6578);
or U8912 (N_8912,N_5046,N_6822);
or U8913 (N_8913,N_6868,N_5697);
and U8914 (N_8914,N_5235,N_6671);
nor U8915 (N_8915,N_5897,N_7474);
nand U8916 (N_8916,N_6185,N_5318);
nand U8917 (N_8917,N_5369,N_5383);
nand U8918 (N_8918,N_7188,N_5434);
and U8919 (N_8919,N_6414,N_6522);
or U8920 (N_8920,N_6733,N_7383);
and U8921 (N_8921,N_5800,N_5139);
and U8922 (N_8922,N_5937,N_7095);
nor U8923 (N_8923,N_6077,N_5841);
or U8924 (N_8924,N_6932,N_6503);
nor U8925 (N_8925,N_7199,N_6304);
nor U8926 (N_8926,N_5115,N_6213);
nand U8927 (N_8927,N_5793,N_6449);
or U8928 (N_8928,N_7493,N_6757);
nor U8929 (N_8929,N_5812,N_5342);
or U8930 (N_8930,N_6692,N_5932);
nor U8931 (N_8931,N_6472,N_5097);
or U8932 (N_8932,N_6049,N_5589);
or U8933 (N_8933,N_7402,N_6573);
and U8934 (N_8934,N_5035,N_6953);
and U8935 (N_8935,N_6272,N_5934);
nand U8936 (N_8936,N_5781,N_6447);
or U8937 (N_8937,N_7365,N_7471);
nor U8938 (N_8938,N_7103,N_5636);
or U8939 (N_8939,N_6777,N_6394);
or U8940 (N_8940,N_5135,N_5959);
and U8941 (N_8941,N_7398,N_7348);
nor U8942 (N_8942,N_7210,N_5908);
and U8943 (N_8943,N_5938,N_7315);
and U8944 (N_8944,N_5704,N_6446);
and U8945 (N_8945,N_6755,N_6836);
and U8946 (N_8946,N_7009,N_5746);
nand U8947 (N_8947,N_6773,N_6032);
nor U8948 (N_8948,N_7380,N_5627);
nand U8949 (N_8949,N_5002,N_6286);
nand U8950 (N_8950,N_5215,N_6995);
or U8951 (N_8951,N_7091,N_5976);
nand U8952 (N_8952,N_6430,N_6426);
nand U8953 (N_8953,N_5372,N_5828);
or U8954 (N_8954,N_6365,N_6637);
nand U8955 (N_8955,N_5543,N_6984);
and U8956 (N_8956,N_6512,N_6783);
or U8957 (N_8957,N_5819,N_7295);
nand U8958 (N_8958,N_5401,N_5208);
and U8959 (N_8959,N_6273,N_7482);
or U8960 (N_8960,N_7089,N_6254);
or U8961 (N_8961,N_6619,N_6426);
and U8962 (N_8962,N_6587,N_6567);
and U8963 (N_8963,N_6719,N_7362);
nor U8964 (N_8964,N_6872,N_5724);
or U8965 (N_8965,N_6758,N_6112);
nor U8966 (N_8966,N_6983,N_5503);
or U8967 (N_8967,N_6505,N_6640);
nand U8968 (N_8968,N_6242,N_6531);
and U8969 (N_8969,N_7388,N_5924);
and U8970 (N_8970,N_5718,N_5954);
nand U8971 (N_8971,N_6520,N_6600);
nor U8972 (N_8972,N_5525,N_5196);
or U8973 (N_8973,N_6884,N_7142);
nor U8974 (N_8974,N_7105,N_6644);
or U8975 (N_8975,N_7117,N_5727);
nand U8976 (N_8976,N_5239,N_5540);
and U8977 (N_8977,N_5494,N_7271);
or U8978 (N_8978,N_6157,N_5779);
nand U8979 (N_8979,N_6913,N_6962);
nor U8980 (N_8980,N_5301,N_5362);
or U8981 (N_8981,N_6049,N_6574);
nor U8982 (N_8982,N_6531,N_7487);
or U8983 (N_8983,N_6141,N_5202);
nor U8984 (N_8984,N_5650,N_6406);
and U8985 (N_8985,N_7055,N_7230);
nand U8986 (N_8986,N_6834,N_7342);
and U8987 (N_8987,N_6254,N_6202);
nand U8988 (N_8988,N_6049,N_5458);
and U8989 (N_8989,N_6890,N_5067);
nor U8990 (N_8990,N_5602,N_6646);
or U8991 (N_8991,N_6320,N_6925);
nand U8992 (N_8992,N_5724,N_5965);
and U8993 (N_8993,N_5360,N_6992);
and U8994 (N_8994,N_5029,N_5244);
nand U8995 (N_8995,N_6711,N_7098);
nor U8996 (N_8996,N_5740,N_6586);
nor U8997 (N_8997,N_7395,N_5693);
nand U8998 (N_8998,N_5250,N_5655);
or U8999 (N_8999,N_7362,N_5335);
or U9000 (N_9000,N_5144,N_7309);
or U9001 (N_9001,N_6082,N_5212);
nand U9002 (N_9002,N_6872,N_7141);
or U9003 (N_9003,N_5150,N_6965);
nor U9004 (N_9004,N_6136,N_6421);
xnor U9005 (N_9005,N_6823,N_5447);
or U9006 (N_9006,N_6916,N_5871);
nor U9007 (N_9007,N_5817,N_5651);
nand U9008 (N_9008,N_5700,N_6767);
nor U9009 (N_9009,N_5361,N_5598);
nor U9010 (N_9010,N_5001,N_6597);
and U9011 (N_9011,N_5435,N_6899);
nand U9012 (N_9012,N_6203,N_6606);
and U9013 (N_9013,N_6390,N_7161);
and U9014 (N_9014,N_5488,N_6610);
nor U9015 (N_9015,N_6026,N_7334);
nor U9016 (N_9016,N_5372,N_6695);
and U9017 (N_9017,N_6517,N_7176);
and U9018 (N_9018,N_6357,N_7177);
nand U9019 (N_9019,N_5426,N_7429);
or U9020 (N_9020,N_6824,N_5619);
nand U9021 (N_9021,N_6472,N_7017);
and U9022 (N_9022,N_5416,N_5176);
nand U9023 (N_9023,N_6365,N_6977);
or U9024 (N_9024,N_6174,N_7482);
or U9025 (N_9025,N_6597,N_5523);
nand U9026 (N_9026,N_5147,N_6807);
or U9027 (N_9027,N_5995,N_7460);
and U9028 (N_9028,N_6813,N_7405);
or U9029 (N_9029,N_6792,N_7027);
or U9030 (N_9030,N_5993,N_7233);
nor U9031 (N_9031,N_5632,N_6039);
nand U9032 (N_9032,N_5222,N_6365);
nor U9033 (N_9033,N_6409,N_5252);
or U9034 (N_9034,N_5194,N_5043);
or U9035 (N_9035,N_6896,N_5150);
and U9036 (N_9036,N_5348,N_7439);
or U9037 (N_9037,N_6356,N_6488);
and U9038 (N_9038,N_6635,N_7140);
or U9039 (N_9039,N_7087,N_5136);
nor U9040 (N_9040,N_5947,N_6862);
or U9041 (N_9041,N_7002,N_7397);
nand U9042 (N_9042,N_7401,N_5501);
nor U9043 (N_9043,N_7288,N_5003);
and U9044 (N_9044,N_6487,N_6271);
and U9045 (N_9045,N_5265,N_6994);
nor U9046 (N_9046,N_6088,N_7456);
and U9047 (N_9047,N_6119,N_6768);
or U9048 (N_9048,N_5310,N_6616);
nor U9049 (N_9049,N_5439,N_7452);
and U9050 (N_9050,N_6616,N_6179);
nand U9051 (N_9051,N_5512,N_5008);
nand U9052 (N_9052,N_7193,N_5612);
and U9053 (N_9053,N_5468,N_5179);
nand U9054 (N_9054,N_6783,N_5932);
nor U9055 (N_9055,N_7075,N_5693);
or U9056 (N_9056,N_5424,N_6664);
and U9057 (N_9057,N_6735,N_5226);
nand U9058 (N_9058,N_6994,N_5984);
nor U9059 (N_9059,N_6891,N_7089);
or U9060 (N_9060,N_5137,N_6682);
nor U9061 (N_9061,N_6494,N_5730);
nor U9062 (N_9062,N_6249,N_6014);
nand U9063 (N_9063,N_6540,N_7331);
nand U9064 (N_9064,N_6995,N_5478);
or U9065 (N_9065,N_6138,N_6572);
nor U9066 (N_9066,N_5463,N_5054);
nand U9067 (N_9067,N_5443,N_6517);
xor U9068 (N_9068,N_6414,N_6176);
or U9069 (N_9069,N_5200,N_5257);
or U9070 (N_9070,N_7128,N_6533);
nor U9071 (N_9071,N_6353,N_6547);
or U9072 (N_9072,N_5879,N_5744);
nor U9073 (N_9073,N_6269,N_6282);
nor U9074 (N_9074,N_7004,N_5940);
nor U9075 (N_9075,N_6263,N_5905);
or U9076 (N_9076,N_6555,N_6744);
or U9077 (N_9077,N_6677,N_6084);
nor U9078 (N_9078,N_5677,N_6735);
nand U9079 (N_9079,N_6202,N_6511);
nand U9080 (N_9080,N_7290,N_7151);
and U9081 (N_9081,N_7023,N_7154);
and U9082 (N_9082,N_6066,N_6605);
nand U9083 (N_9083,N_7222,N_6978);
nor U9084 (N_9084,N_5718,N_5457);
or U9085 (N_9085,N_6619,N_5265);
nand U9086 (N_9086,N_5896,N_6586);
and U9087 (N_9087,N_5071,N_5477);
or U9088 (N_9088,N_7060,N_7217);
nor U9089 (N_9089,N_6066,N_7377);
nand U9090 (N_9090,N_7233,N_7143);
and U9091 (N_9091,N_5853,N_6949);
and U9092 (N_9092,N_6948,N_7317);
nor U9093 (N_9093,N_5923,N_5531);
and U9094 (N_9094,N_5647,N_7114);
nand U9095 (N_9095,N_6824,N_6574);
and U9096 (N_9096,N_6965,N_5503);
and U9097 (N_9097,N_6267,N_6727);
and U9098 (N_9098,N_7352,N_6425);
nor U9099 (N_9099,N_7012,N_5598);
and U9100 (N_9100,N_5614,N_7127);
nor U9101 (N_9101,N_6415,N_5869);
and U9102 (N_9102,N_5726,N_7389);
and U9103 (N_9103,N_7084,N_6628);
or U9104 (N_9104,N_6677,N_5106);
and U9105 (N_9105,N_6261,N_7138);
nor U9106 (N_9106,N_5469,N_6005);
or U9107 (N_9107,N_7253,N_7183);
nor U9108 (N_9108,N_6447,N_6110);
or U9109 (N_9109,N_5546,N_7407);
or U9110 (N_9110,N_7062,N_6616);
and U9111 (N_9111,N_7202,N_6171);
nand U9112 (N_9112,N_7215,N_5850);
nor U9113 (N_9113,N_6886,N_5834);
nand U9114 (N_9114,N_6469,N_5264);
and U9115 (N_9115,N_5221,N_5732);
nor U9116 (N_9116,N_6944,N_6383);
or U9117 (N_9117,N_5770,N_5839);
and U9118 (N_9118,N_5966,N_6401);
nand U9119 (N_9119,N_5084,N_7106);
nor U9120 (N_9120,N_5049,N_5469);
or U9121 (N_9121,N_5984,N_6104);
and U9122 (N_9122,N_5541,N_5045);
nand U9123 (N_9123,N_6900,N_7355);
nor U9124 (N_9124,N_6932,N_7039);
nor U9125 (N_9125,N_6828,N_6305);
or U9126 (N_9126,N_5713,N_5616);
nor U9127 (N_9127,N_7023,N_5553);
xor U9128 (N_9128,N_7431,N_5813);
nor U9129 (N_9129,N_5239,N_7375);
or U9130 (N_9130,N_6865,N_6480);
nor U9131 (N_9131,N_5632,N_5386);
nor U9132 (N_9132,N_5245,N_7448);
and U9133 (N_9133,N_7494,N_5695);
and U9134 (N_9134,N_6529,N_5845);
or U9135 (N_9135,N_5307,N_7469);
nor U9136 (N_9136,N_6293,N_7158);
nand U9137 (N_9137,N_5543,N_7232);
nor U9138 (N_9138,N_6481,N_7114);
or U9139 (N_9139,N_5062,N_6566);
or U9140 (N_9140,N_6305,N_7256);
nand U9141 (N_9141,N_5392,N_6185);
or U9142 (N_9142,N_6645,N_5376);
and U9143 (N_9143,N_7102,N_6282);
xnor U9144 (N_9144,N_5718,N_5541);
nand U9145 (N_9145,N_6608,N_6438);
nor U9146 (N_9146,N_6886,N_6797);
or U9147 (N_9147,N_6259,N_6888);
or U9148 (N_9148,N_6725,N_5361);
nand U9149 (N_9149,N_7074,N_6924);
or U9150 (N_9150,N_5242,N_6926);
or U9151 (N_9151,N_5076,N_6882);
and U9152 (N_9152,N_6595,N_6217);
and U9153 (N_9153,N_5450,N_5797);
or U9154 (N_9154,N_6936,N_5508);
and U9155 (N_9155,N_6457,N_7483);
and U9156 (N_9156,N_5636,N_7287);
nand U9157 (N_9157,N_6112,N_7365);
and U9158 (N_9158,N_6360,N_5707);
or U9159 (N_9159,N_6042,N_6145);
and U9160 (N_9160,N_7484,N_7401);
nor U9161 (N_9161,N_6993,N_5675);
or U9162 (N_9162,N_5105,N_6798);
and U9163 (N_9163,N_5207,N_5906);
nor U9164 (N_9164,N_6405,N_5212);
and U9165 (N_9165,N_6565,N_5213);
or U9166 (N_9166,N_5860,N_5958);
nand U9167 (N_9167,N_5840,N_5395);
or U9168 (N_9168,N_6582,N_6964);
or U9169 (N_9169,N_6744,N_7080);
or U9170 (N_9170,N_6143,N_6827);
and U9171 (N_9171,N_6448,N_5356);
nor U9172 (N_9172,N_5712,N_5221);
nor U9173 (N_9173,N_5353,N_6928);
or U9174 (N_9174,N_7190,N_5122);
and U9175 (N_9175,N_5688,N_7000);
or U9176 (N_9176,N_6035,N_5111);
and U9177 (N_9177,N_5413,N_7226);
and U9178 (N_9178,N_5396,N_5482);
nand U9179 (N_9179,N_6545,N_5307);
nor U9180 (N_9180,N_6292,N_5272);
and U9181 (N_9181,N_5066,N_6115);
and U9182 (N_9182,N_7058,N_7290);
or U9183 (N_9183,N_7163,N_5544);
or U9184 (N_9184,N_7335,N_7378);
nand U9185 (N_9185,N_6524,N_6430);
nand U9186 (N_9186,N_6043,N_5840);
and U9187 (N_9187,N_5801,N_6519);
and U9188 (N_9188,N_6543,N_5736);
nand U9189 (N_9189,N_6693,N_5676);
and U9190 (N_9190,N_6517,N_5373);
nor U9191 (N_9191,N_7131,N_6467);
nand U9192 (N_9192,N_6943,N_7467);
nor U9193 (N_9193,N_6869,N_5878);
nor U9194 (N_9194,N_5951,N_5072);
or U9195 (N_9195,N_6492,N_6579);
nand U9196 (N_9196,N_5267,N_5246);
nor U9197 (N_9197,N_7317,N_6823);
nor U9198 (N_9198,N_5296,N_6572);
nand U9199 (N_9199,N_5424,N_5022);
nor U9200 (N_9200,N_6683,N_5857);
nand U9201 (N_9201,N_5017,N_6319);
nor U9202 (N_9202,N_5373,N_6119);
and U9203 (N_9203,N_5046,N_6674);
nor U9204 (N_9204,N_7400,N_5688);
and U9205 (N_9205,N_7319,N_7017);
and U9206 (N_9206,N_7437,N_6203);
nor U9207 (N_9207,N_7254,N_6881);
or U9208 (N_9208,N_5736,N_6668);
nor U9209 (N_9209,N_7414,N_5552);
nand U9210 (N_9210,N_5760,N_5476);
or U9211 (N_9211,N_7159,N_5161);
nand U9212 (N_9212,N_5679,N_6153);
nor U9213 (N_9213,N_5281,N_5861);
nand U9214 (N_9214,N_6794,N_6704);
or U9215 (N_9215,N_6831,N_6032);
or U9216 (N_9216,N_5306,N_6656);
or U9217 (N_9217,N_6835,N_6679);
and U9218 (N_9218,N_5675,N_5385);
or U9219 (N_9219,N_6374,N_5230);
and U9220 (N_9220,N_6805,N_6349);
or U9221 (N_9221,N_5780,N_6013);
nor U9222 (N_9222,N_7426,N_7337);
or U9223 (N_9223,N_6633,N_5043);
and U9224 (N_9224,N_6733,N_5695);
or U9225 (N_9225,N_5896,N_5711);
nor U9226 (N_9226,N_6274,N_5097);
nand U9227 (N_9227,N_7000,N_5378);
nand U9228 (N_9228,N_6654,N_7455);
nor U9229 (N_9229,N_7276,N_7242);
nor U9230 (N_9230,N_6145,N_6311);
and U9231 (N_9231,N_7103,N_7269);
or U9232 (N_9232,N_6783,N_5107);
xnor U9233 (N_9233,N_6492,N_5689);
and U9234 (N_9234,N_6130,N_6996);
and U9235 (N_9235,N_7102,N_6961);
nor U9236 (N_9236,N_5093,N_7317);
or U9237 (N_9237,N_5887,N_5737);
and U9238 (N_9238,N_6627,N_7351);
and U9239 (N_9239,N_7414,N_6652);
nand U9240 (N_9240,N_6829,N_7138);
and U9241 (N_9241,N_5681,N_7078);
or U9242 (N_9242,N_6122,N_5132);
or U9243 (N_9243,N_5827,N_5983);
nand U9244 (N_9244,N_5017,N_6212);
nand U9245 (N_9245,N_5892,N_5997);
or U9246 (N_9246,N_7407,N_6453);
nor U9247 (N_9247,N_7029,N_6786);
or U9248 (N_9248,N_5821,N_5413);
and U9249 (N_9249,N_6469,N_6163);
nor U9250 (N_9250,N_7476,N_5348);
or U9251 (N_9251,N_6558,N_6437);
nor U9252 (N_9252,N_5297,N_6877);
nor U9253 (N_9253,N_7278,N_6178);
or U9254 (N_9254,N_6509,N_5776);
nand U9255 (N_9255,N_7124,N_6602);
and U9256 (N_9256,N_7397,N_5147);
and U9257 (N_9257,N_5821,N_6221);
and U9258 (N_9258,N_6295,N_5634);
nor U9259 (N_9259,N_6601,N_5084);
nand U9260 (N_9260,N_7031,N_5519);
or U9261 (N_9261,N_5193,N_6687);
or U9262 (N_9262,N_6797,N_7141);
nor U9263 (N_9263,N_6256,N_5537);
nand U9264 (N_9264,N_6901,N_7032);
or U9265 (N_9265,N_7430,N_5746);
or U9266 (N_9266,N_7082,N_5377);
and U9267 (N_9267,N_6495,N_5730);
and U9268 (N_9268,N_5096,N_5328);
and U9269 (N_9269,N_6397,N_6701);
and U9270 (N_9270,N_5557,N_6340);
nor U9271 (N_9271,N_6252,N_5150);
nor U9272 (N_9272,N_5178,N_5555);
and U9273 (N_9273,N_5190,N_7429);
nand U9274 (N_9274,N_7366,N_7084);
or U9275 (N_9275,N_6657,N_6646);
nand U9276 (N_9276,N_6294,N_5478);
nor U9277 (N_9277,N_5000,N_7343);
or U9278 (N_9278,N_6862,N_6494);
nor U9279 (N_9279,N_6432,N_5450);
or U9280 (N_9280,N_6445,N_7214);
nor U9281 (N_9281,N_5914,N_7152);
nand U9282 (N_9282,N_6573,N_5321);
and U9283 (N_9283,N_5724,N_6266);
and U9284 (N_9284,N_6965,N_6667);
or U9285 (N_9285,N_6538,N_5768);
xnor U9286 (N_9286,N_7454,N_6877);
or U9287 (N_9287,N_5645,N_7340);
or U9288 (N_9288,N_6360,N_6176);
and U9289 (N_9289,N_7039,N_7085);
nor U9290 (N_9290,N_6610,N_5963);
nand U9291 (N_9291,N_5468,N_6775);
and U9292 (N_9292,N_6165,N_7401);
and U9293 (N_9293,N_6618,N_7127);
nor U9294 (N_9294,N_6310,N_6993);
nor U9295 (N_9295,N_6972,N_6112);
and U9296 (N_9296,N_5382,N_5279);
and U9297 (N_9297,N_6184,N_6209);
nand U9298 (N_9298,N_5997,N_6499);
xor U9299 (N_9299,N_5079,N_5756);
nand U9300 (N_9300,N_7235,N_6819);
nand U9301 (N_9301,N_6024,N_6399);
nor U9302 (N_9302,N_6770,N_6182);
nand U9303 (N_9303,N_5379,N_6627);
nor U9304 (N_9304,N_6411,N_5620);
nor U9305 (N_9305,N_6057,N_5998);
and U9306 (N_9306,N_6670,N_5610);
or U9307 (N_9307,N_6638,N_5876);
nor U9308 (N_9308,N_5349,N_5300);
nor U9309 (N_9309,N_6174,N_6743);
or U9310 (N_9310,N_6541,N_5238);
nand U9311 (N_9311,N_5248,N_6153);
nor U9312 (N_9312,N_7286,N_6255);
nand U9313 (N_9313,N_6110,N_5067);
nand U9314 (N_9314,N_6252,N_5890);
nor U9315 (N_9315,N_6461,N_7068);
xor U9316 (N_9316,N_5995,N_5970);
or U9317 (N_9317,N_5781,N_6863);
and U9318 (N_9318,N_7310,N_6661);
nor U9319 (N_9319,N_6731,N_6738);
xnor U9320 (N_9320,N_5414,N_5495);
and U9321 (N_9321,N_6822,N_6597);
nand U9322 (N_9322,N_5304,N_6453);
nand U9323 (N_9323,N_5701,N_5951);
nor U9324 (N_9324,N_5364,N_5646);
and U9325 (N_9325,N_6060,N_5673);
nor U9326 (N_9326,N_6132,N_7045);
and U9327 (N_9327,N_7490,N_5508);
or U9328 (N_9328,N_6609,N_7423);
or U9329 (N_9329,N_6362,N_7291);
and U9330 (N_9330,N_6897,N_7409);
and U9331 (N_9331,N_5975,N_5201);
nor U9332 (N_9332,N_6720,N_6088);
and U9333 (N_9333,N_5371,N_5338);
nand U9334 (N_9334,N_5263,N_5506);
or U9335 (N_9335,N_5894,N_5236);
or U9336 (N_9336,N_7142,N_6359);
nand U9337 (N_9337,N_5983,N_6183);
nand U9338 (N_9338,N_6722,N_6070);
and U9339 (N_9339,N_5471,N_6021);
and U9340 (N_9340,N_5267,N_6134);
xnor U9341 (N_9341,N_5621,N_7226);
nand U9342 (N_9342,N_5954,N_5710);
nor U9343 (N_9343,N_6745,N_6785);
nand U9344 (N_9344,N_7164,N_6722);
nor U9345 (N_9345,N_5101,N_5314);
or U9346 (N_9346,N_6037,N_6759);
and U9347 (N_9347,N_5576,N_7423);
or U9348 (N_9348,N_7454,N_5363);
nor U9349 (N_9349,N_5605,N_5731);
nand U9350 (N_9350,N_6451,N_5490);
nand U9351 (N_9351,N_6747,N_5450);
nand U9352 (N_9352,N_5086,N_5623);
and U9353 (N_9353,N_5469,N_7062);
nor U9354 (N_9354,N_7123,N_7486);
nor U9355 (N_9355,N_6941,N_5237);
and U9356 (N_9356,N_6559,N_6365);
and U9357 (N_9357,N_5794,N_6762);
or U9358 (N_9358,N_7013,N_5463);
or U9359 (N_9359,N_6366,N_6041);
nand U9360 (N_9360,N_7142,N_5637);
nand U9361 (N_9361,N_7078,N_6556);
and U9362 (N_9362,N_5272,N_6078);
nor U9363 (N_9363,N_5456,N_5284);
and U9364 (N_9364,N_6111,N_6175);
nor U9365 (N_9365,N_5006,N_6067);
or U9366 (N_9366,N_5645,N_7313);
or U9367 (N_9367,N_5939,N_6918);
or U9368 (N_9368,N_7155,N_5432);
nand U9369 (N_9369,N_5191,N_5097);
nor U9370 (N_9370,N_6489,N_5648);
or U9371 (N_9371,N_6101,N_5346);
nor U9372 (N_9372,N_7037,N_6324);
nor U9373 (N_9373,N_5424,N_6474);
or U9374 (N_9374,N_5271,N_6334);
and U9375 (N_9375,N_6293,N_7238);
nand U9376 (N_9376,N_7454,N_6474);
nor U9377 (N_9377,N_5042,N_7202);
nor U9378 (N_9378,N_5143,N_5641);
and U9379 (N_9379,N_7385,N_6517);
or U9380 (N_9380,N_5452,N_5321);
nand U9381 (N_9381,N_5875,N_7449);
nor U9382 (N_9382,N_6135,N_5297);
and U9383 (N_9383,N_5971,N_5348);
or U9384 (N_9384,N_7024,N_6189);
and U9385 (N_9385,N_6696,N_6447);
or U9386 (N_9386,N_6339,N_6603);
nor U9387 (N_9387,N_5050,N_5510);
nand U9388 (N_9388,N_7013,N_5320);
nor U9389 (N_9389,N_5378,N_6822);
and U9390 (N_9390,N_6365,N_7017);
nand U9391 (N_9391,N_5787,N_5182);
nor U9392 (N_9392,N_7298,N_7209);
and U9393 (N_9393,N_6884,N_5437);
and U9394 (N_9394,N_6358,N_6826);
or U9395 (N_9395,N_7052,N_6772);
or U9396 (N_9396,N_7495,N_6316);
nand U9397 (N_9397,N_5681,N_5045);
nor U9398 (N_9398,N_5043,N_5789);
nor U9399 (N_9399,N_5490,N_5372);
nor U9400 (N_9400,N_6406,N_6988);
and U9401 (N_9401,N_7045,N_7480);
nor U9402 (N_9402,N_6896,N_6061);
nand U9403 (N_9403,N_5298,N_7173);
nand U9404 (N_9404,N_7286,N_5139);
and U9405 (N_9405,N_7459,N_5561);
or U9406 (N_9406,N_5979,N_6841);
xor U9407 (N_9407,N_5374,N_5022);
or U9408 (N_9408,N_6962,N_7405);
nor U9409 (N_9409,N_5844,N_6279);
nand U9410 (N_9410,N_5661,N_7458);
and U9411 (N_9411,N_5748,N_7407);
nand U9412 (N_9412,N_7060,N_6590);
and U9413 (N_9413,N_7227,N_6838);
nand U9414 (N_9414,N_5629,N_7356);
nand U9415 (N_9415,N_5335,N_5330);
and U9416 (N_9416,N_6592,N_6959);
nor U9417 (N_9417,N_5132,N_6922);
and U9418 (N_9418,N_7403,N_7060);
or U9419 (N_9419,N_6835,N_6386);
nor U9420 (N_9420,N_7485,N_5084);
or U9421 (N_9421,N_6835,N_5417);
nor U9422 (N_9422,N_5347,N_6549);
or U9423 (N_9423,N_5885,N_6777);
nand U9424 (N_9424,N_7315,N_5963);
and U9425 (N_9425,N_6448,N_6557);
nand U9426 (N_9426,N_5345,N_6943);
and U9427 (N_9427,N_5430,N_5879);
nand U9428 (N_9428,N_5640,N_5394);
and U9429 (N_9429,N_7142,N_6063);
and U9430 (N_9430,N_6989,N_5580);
and U9431 (N_9431,N_6592,N_5722);
nor U9432 (N_9432,N_6194,N_6168);
and U9433 (N_9433,N_7426,N_5698);
and U9434 (N_9434,N_6859,N_5048);
nand U9435 (N_9435,N_5439,N_5373);
nand U9436 (N_9436,N_7230,N_5115);
nand U9437 (N_9437,N_5263,N_6633);
nand U9438 (N_9438,N_6078,N_6435);
nor U9439 (N_9439,N_5530,N_6585);
nor U9440 (N_9440,N_7121,N_6443);
and U9441 (N_9441,N_5395,N_6803);
nand U9442 (N_9442,N_7113,N_5858);
nor U9443 (N_9443,N_6341,N_6406);
and U9444 (N_9444,N_5029,N_7168);
nor U9445 (N_9445,N_7414,N_5578);
or U9446 (N_9446,N_7337,N_5696);
and U9447 (N_9447,N_6097,N_6821);
nor U9448 (N_9448,N_6082,N_7328);
or U9449 (N_9449,N_5273,N_6281);
and U9450 (N_9450,N_7074,N_6942);
nand U9451 (N_9451,N_7082,N_7475);
or U9452 (N_9452,N_6883,N_5328);
and U9453 (N_9453,N_5662,N_7150);
and U9454 (N_9454,N_6834,N_6630);
and U9455 (N_9455,N_7368,N_5883);
nand U9456 (N_9456,N_5246,N_7269);
or U9457 (N_9457,N_7258,N_7344);
and U9458 (N_9458,N_7411,N_6058);
or U9459 (N_9459,N_7014,N_5347);
nand U9460 (N_9460,N_7313,N_5510);
nor U9461 (N_9461,N_6787,N_5893);
and U9462 (N_9462,N_6859,N_7421);
and U9463 (N_9463,N_5983,N_5720);
nor U9464 (N_9464,N_5883,N_5112);
or U9465 (N_9465,N_6764,N_7395);
nor U9466 (N_9466,N_5371,N_7359);
and U9467 (N_9467,N_5512,N_5506);
nand U9468 (N_9468,N_5826,N_7323);
nand U9469 (N_9469,N_7118,N_6842);
xor U9470 (N_9470,N_6171,N_6347);
and U9471 (N_9471,N_5467,N_5182);
and U9472 (N_9472,N_7245,N_5610);
or U9473 (N_9473,N_5901,N_6431);
and U9474 (N_9474,N_6594,N_6434);
or U9475 (N_9475,N_5924,N_5184);
or U9476 (N_9476,N_5259,N_5042);
and U9477 (N_9477,N_6095,N_6482);
nand U9478 (N_9478,N_6487,N_6702);
or U9479 (N_9479,N_5083,N_5597);
nor U9480 (N_9480,N_6304,N_5442);
and U9481 (N_9481,N_6056,N_5568);
nand U9482 (N_9482,N_7289,N_5974);
and U9483 (N_9483,N_7210,N_6609);
and U9484 (N_9484,N_7027,N_7347);
nand U9485 (N_9485,N_7429,N_6227);
and U9486 (N_9486,N_5419,N_7391);
or U9487 (N_9487,N_6540,N_5236);
nor U9488 (N_9488,N_7186,N_7416);
and U9489 (N_9489,N_6786,N_5865);
or U9490 (N_9490,N_5081,N_5889);
or U9491 (N_9491,N_6036,N_6011);
or U9492 (N_9492,N_5232,N_6790);
nor U9493 (N_9493,N_6407,N_6043);
and U9494 (N_9494,N_6685,N_6498);
or U9495 (N_9495,N_5026,N_5856);
and U9496 (N_9496,N_6686,N_6980);
nor U9497 (N_9497,N_5485,N_6345);
or U9498 (N_9498,N_6165,N_7457);
nor U9499 (N_9499,N_6421,N_5242);
and U9500 (N_9500,N_5405,N_6877);
and U9501 (N_9501,N_5364,N_6642);
or U9502 (N_9502,N_5151,N_5969);
or U9503 (N_9503,N_5213,N_6494);
nand U9504 (N_9504,N_7023,N_6081);
or U9505 (N_9505,N_6479,N_7207);
and U9506 (N_9506,N_5570,N_5929);
and U9507 (N_9507,N_5788,N_6638);
or U9508 (N_9508,N_5941,N_5274);
or U9509 (N_9509,N_6315,N_6390);
nor U9510 (N_9510,N_6193,N_6406);
nor U9511 (N_9511,N_5009,N_6645);
and U9512 (N_9512,N_6191,N_7472);
or U9513 (N_9513,N_6305,N_7146);
and U9514 (N_9514,N_5527,N_6825);
or U9515 (N_9515,N_6931,N_5707);
or U9516 (N_9516,N_5037,N_5102);
nand U9517 (N_9517,N_6060,N_7334);
and U9518 (N_9518,N_5746,N_6047);
or U9519 (N_9519,N_5366,N_5849);
nor U9520 (N_9520,N_5091,N_7474);
or U9521 (N_9521,N_6611,N_5329);
nor U9522 (N_9522,N_5108,N_6428);
or U9523 (N_9523,N_6736,N_5924);
nand U9524 (N_9524,N_7359,N_5529);
nand U9525 (N_9525,N_7137,N_6115);
nor U9526 (N_9526,N_5485,N_5023);
nand U9527 (N_9527,N_5991,N_5661);
and U9528 (N_9528,N_6228,N_7043);
or U9529 (N_9529,N_5533,N_6935);
nor U9530 (N_9530,N_5960,N_5519);
and U9531 (N_9531,N_6813,N_6864);
and U9532 (N_9532,N_7292,N_5334);
nor U9533 (N_9533,N_7235,N_5162);
and U9534 (N_9534,N_7408,N_5610);
nor U9535 (N_9535,N_6972,N_7315);
nand U9536 (N_9536,N_5682,N_7121);
nor U9537 (N_9537,N_6512,N_7147);
and U9538 (N_9538,N_6773,N_6516);
nand U9539 (N_9539,N_5093,N_6603);
or U9540 (N_9540,N_7013,N_5120);
nor U9541 (N_9541,N_5878,N_6577);
and U9542 (N_9542,N_5294,N_6623);
or U9543 (N_9543,N_5905,N_5528);
or U9544 (N_9544,N_6567,N_7021);
nand U9545 (N_9545,N_5558,N_6838);
nor U9546 (N_9546,N_5844,N_7259);
and U9547 (N_9547,N_6140,N_5898);
or U9548 (N_9548,N_6001,N_6164);
nand U9549 (N_9549,N_5282,N_5068);
nand U9550 (N_9550,N_5917,N_6078);
nand U9551 (N_9551,N_6526,N_6506);
nand U9552 (N_9552,N_6937,N_7476);
nand U9553 (N_9553,N_6811,N_5801);
nand U9554 (N_9554,N_5580,N_7326);
nor U9555 (N_9555,N_7448,N_6433);
nor U9556 (N_9556,N_5548,N_7322);
and U9557 (N_9557,N_5859,N_6382);
and U9558 (N_9558,N_5634,N_5944);
and U9559 (N_9559,N_6747,N_6385);
nand U9560 (N_9560,N_6684,N_5188);
nor U9561 (N_9561,N_6006,N_5910);
nor U9562 (N_9562,N_7427,N_6277);
nor U9563 (N_9563,N_5400,N_5497);
or U9564 (N_9564,N_7241,N_5640);
or U9565 (N_9565,N_5255,N_7170);
or U9566 (N_9566,N_5758,N_6702);
nor U9567 (N_9567,N_7104,N_5433);
nor U9568 (N_9568,N_6244,N_5258);
or U9569 (N_9569,N_6407,N_6446);
nand U9570 (N_9570,N_5519,N_6229);
or U9571 (N_9571,N_6789,N_5407);
nand U9572 (N_9572,N_5295,N_6685);
and U9573 (N_9573,N_7456,N_5836);
nand U9574 (N_9574,N_5044,N_7473);
nor U9575 (N_9575,N_5963,N_6802);
and U9576 (N_9576,N_5110,N_6935);
and U9577 (N_9577,N_5368,N_5136);
or U9578 (N_9578,N_5394,N_6507);
and U9579 (N_9579,N_6566,N_7124);
and U9580 (N_9580,N_5308,N_7354);
nor U9581 (N_9581,N_7352,N_5493);
nand U9582 (N_9582,N_6001,N_7143);
nand U9583 (N_9583,N_5852,N_6677);
or U9584 (N_9584,N_6839,N_5294);
and U9585 (N_9585,N_7315,N_6483);
and U9586 (N_9586,N_5877,N_5659);
or U9587 (N_9587,N_5438,N_7480);
nand U9588 (N_9588,N_6079,N_7313);
nor U9589 (N_9589,N_7066,N_5291);
and U9590 (N_9590,N_5043,N_5412);
or U9591 (N_9591,N_5404,N_5887);
nor U9592 (N_9592,N_6880,N_6281);
nand U9593 (N_9593,N_5356,N_7089);
nor U9594 (N_9594,N_6943,N_7255);
and U9595 (N_9595,N_5166,N_7255);
nand U9596 (N_9596,N_6441,N_5949);
and U9597 (N_9597,N_6062,N_7366);
xnor U9598 (N_9598,N_6054,N_6624);
nor U9599 (N_9599,N_6516,N_7494);
and U9600 (N_9600,N_6234,N_7188);
nor U9601 (N_9601,N_5893,N_7258);
or U9602 (N_9602,N_5418,N_6036);
nor U9603 (N_9603,N_6561,N_6843);
or U9604 (N_9604,N_5138,N_5792);
or U9605 (N_9605,N_5211,N_5952);
nand U9606 (N_9606,N_5708,N_7024);
nand U9607 (N_9607,N_6883,N_5431);
nor U9608 (N_9608,N_6587,N_7276);
or U9609 (N_9609,N_5193,N_5683);
or U9610 (N_9610,N_6827,N_7233);
or U9611 (N_9611,N_5088,N_6861);
nand U9612 (N_9612,N_5204,N_6686);
nor U9613 (N_9613,N_5260,N_6568);
nor U9614 (N_9614,N_5318,N_5359);
nand U9615 (N_9615,N_5009,N_6864);
nand U9616 (N_9616,N_5293,N_6859);
nor U9617 (N_9617,N_6471,N_5672);
nand U9618 (N_9618,N_6199,N_6460);
nor U9619 (N_9619,N_6893,N_5859);
nand U9620 (N_9620,N_5506,N_6312);
or U9621 (N_9621,N_6805,N_6827);
nand U9622 (N_9622,N_6860,N_6795);
nand U9623 (N_9623,N_6934,N_6927);
nor U9624 (N_9624,N_6942,N_7090);
and U9625 (N_9625,N_7095,N_6647);
nor U9626 (N_9626,N_5156,N_6308);
nand U9627 (N_9627,N_6174,N_6544);
nor U9628 (N_9628,N_7271,N_6392);
and U9629 (N_9629,N_6841,N_5791);
or U9630 (N_9630,N_5716,N_6451);
and U9631 (N_9631,N_5137,N_5218);
nor U9632 (N_9632,N_5885,N_5276);
and U9633 (N_9633,N_5357,N_6684);
or U9634 (N_9634,N_5340,N_6499);
nor U9635 (N_9635,N_5921,N_6233);
nor U9636 (N_9636,N_6889,N_6944);
nor U9637 (N_9637,N_6837,N_5396);
or U9638 (N_9638,N_6303,N_6656);
and U9639 (N_9639,N_5119,N_5508);
and U9640 (N_9640,N_7096,N_7227);
or U9641 (N_9641,N_6966,N_5102);
or U9642 (N_9642,N_5638,N_5637);
nor U9643 (N_9643,N_5499,N_6902);
nand U9644 (N_9644,N_6655,N_6944);
or U9645 (N_9645,N_7320,N_6640);
nor U9646 (N_9646,N_6474,N_7453);
nand U9647 (N_9647,N_6207,N_5055);
nand U9648 (N_9648,N_7128,N_6634);
nor U9649 (N_9649,N_7383,N_5833);
and U9650 (N_9650,N_5094,N_6589);
and U9651 (N_9651,N_5409,N_7227);
or U9652 (N_9652,N_5193,N_7101);
nand U9653 (N_9653,N_7478,N_5149);
nand U9654 (N_9654,N_7371,N_5435);
and U9655 (N_9655,N_7025,N_5397);
nor U9656 (N_9656,N_6025,N_6028);
or U9657 (N_9657,N_7208,N_6152);
nand U9658 (N_9658,N_6464,N_6401);
and U9659 (N_9659,N_7246,N_5117);
xor U9660 (N_9660,N_6245,N_5196);
or U9661 (N_9661,N_5252,N_5647);
nand U9662 (N_9662,N_6862,N_6068);
nor U9663 (N_9663,N_6031,N_6987);
nor U9664 (N_9664,N_5288,N_6647);
or U9665 (N_9665,N_6991,N_7391);
nand U9666 (N_9666,N_5418,N_6136);
and U9667 (N_9667,N_5452,N_5125);
nand U9668 (N_9668,N_7128,N_6612);
nor U9669 (N_9669,N_5135,N_6861);
nand U9670 (N_9670,N_5559,N_5475);
nor U9671 (N_9671,N_6663,N_5961);
nand U9672 (N_9672,N_5966,N_6785);
nor U9673 (N_9673,N_5555,N_6829);
nand U9674 (N_9674,N_6051,N_6523);
nor U9675 (N_9675,N_5085,N_6026);
and U9676 (N_9676,N_5403,N_6633);
nand U9677 (N_9677,N_5157,N_5421);
or U9678 (N_9678,N_5970,N_6189);
or U9679 (N_9679,N_7105,N_7386);
nand U9680 (N_9680,N_5488,N_5612);
or U9681 (N_9681,N_6156,N_5260);
or U9682 (N_9682,N_5861,N_5946);
and U9683 (N_9683,N_6358,N_5149);
nand U9684 (N_9684,N_7487,N_5686);
and U9685 (N_9685,N_6203,N_5464);
nor U9686 (N_9686,N_7007,N_6226);
nor U9687 (N_9687,N_5688,N_6891);
nor U9688 (N_9688,N_5943,N_5078);
nor U9689 (N_9689,N_6636,N_6995);
nor U9690 (N_9690,N_7151,N_5500);
or U9691 (N_9691,N_5270,N_6342);
nor U9692 (N_9692,N_6613,N_6000);
or U9693 (N_9693,N_6859,N_7253);
and U9694 (N_9694,N_6890,N_6581);
and U9695 (N_9695,N_6974,N_6733);
xnor U9696 (N_9696,N_5830,N_7248);
nor U9697 (N_9697,N_7387,N_6689);
or U9698 (N_9698,N_7179,N_7007);
nand U9699 (N_9699,N_6642,N_5730);
nand U9700 (N_9700,N_5190,N_5132);
nor U9701 (N_9701,N_5717,N_5096);
and U9702 (N_9702,N_5676,N_7307);
nor U9703 (N_9703,N_6245,N_7438);
and U9704 (N_9704,N_7383,N_5460);
or U9705 (N_9705,N_6157,N_6917);
and U9706 (N_9706,N_5733,N_6029);
xor U9707 (N_9707,N_6163,N_5701);
nand U9708 (N_9708,N_6420,N_7132);
and U9709 (N_9709,N_5052,N_5065);
nand U9710 (N_9710,N_5635,N_5420);
nand U9711 (N_9711,N_6344,N_7038);
nand U9712 (N_9712,N_5507,N_6834);
nor U9713 (N_9713,N_6537,N_6693);
nand U9714 (N_9714,N_5932,N_5935);
and U9715 (N_9715,N_5384,N_6880);
or U9716 (N_9716,N_6887,N_5749);
and U9717 (N_9717,N_5272,N_5315);
or U9718 (N_9718,N_6330,N_6304);
nand U9719 (N_9719,N_7148,N_5479);
or U9720 (N_9720,N_5079,N_5903);
nand U9721 (N_9721,N_5835,N_6414);
and U9722 (N_9722,N_5220,N_6485);
nand U9723 (N_9723,N_5145,N_5949);
and U9724 (N_9724,N_5137,N_6087);
and U9725 (N_9725,N_7194,N_5535);
nand U9726 (N_9726,N_7438,N_5011);
and U9727 (N_9727,N_7384,N_5348);
and U9728 (N_9728,N_5869,N_6798);
or U9729 (N_9729,N_6103,N_7369);
or U9730 (N_9730,N_6707,N_6223);
nand U9731 (N_9731,N_5452,N_6726);
or U9732 (N_9732,N_5621,N_7367);
nor U9733 (N_9733,N_6723,N_5707);
and U9734 (N_9734,N_5217,N_5917);
nor U9735 (N_9735,N_6423,N_6922);
nand U9736 (N_9736,N_5003,N_6560);
nor U9737 (N_9737,N_5786,N_7364);
nor U9738 (N_9738,N_5808,N_6642);
or U9739 (N_9739,N_6788,N_6567);
nand U9740 (N_9740,N_5765,N_7385);
and U9741 (N_9741,N_6676,N_6470);
nor U9742 (N_9742,N_6705,N_7269);
and U9743 (N_9743,N_6291,N_7286);
nand U9744 (N_9744,N_6554,N_6652);
or U9745 (N_9745,N_7467,N_6865);
or U9746 (N_9746,N_7231,N_6074);
and U9747 (N_9747,N_5905,N_7305);
nand U9748 (N_9748,N_7329,N_7096);
and U9749 (N_9749,N_6936,N_5549);
and U9750 (N_9750,N_5456,N_5363);
and U9751 (N_9751,N_6747,N_6985);
or U9752 (N_9752,N_6448,N_7431);
nand U9753 (N_9753,N_5636,N_5388);
nand U9754 (N_9754,N_7423,N_5583);
nand U9755 (N_9755,N_5310,N_5813);
or U9756 (N_9756,N_5613,N_5419);
or U9757 (N_9757,N_5770,N_6347);
and U9758 (N_9758,N_5119,N_7381);
nand U9759 (N_9759,N_6990,N_5432);
and U9760 (N_9760,N_5024,N_6272);
nand U9761 (N_9761,N_6323,N_7165);
nor U9762 (N_9762,N_5192,N_6254);
and U9763 (N_9763,N_6397,N_5846);
nand U9764 (N_9764,N_5318,N_6896);
nand U9765 (N_9765,N_6545,N_7287);
and U9766 (N_9766,N_6495,N_5256);
nor U9767 (N_9767,N_5708,N_5563);
or U9768 (N_9768,N_5942,N_5478);
nand U9769 (N_9769,N_5257,N_5588);
or U9770 (N_9770,N_5771,N_5982);
or U9771 (N_9771,N_7252,N_5812);
nand U9772 (N_9772,N_6421,N_5216);
nor U9773 (N_9773,N_5488,N_5556);
or U9774 (N_9774,N_5492,N_6637);
nor U9775 (N_9775,N_5797,N_5275);
and U9776 (N_9776,N_7278,N_5011);
and U9777 (N_9777,N_6861,N_5838);
and U9778 (N_9778,N_5765,N_6709);
or U9779 (N_9779,N_6076,N_7115);
and U9780 (N_9780,N_5294,N_6085);
nand U9781 (N_9781,N_7276,N_7303);
or U9782 (N_9782,N_5360,N_5723);
nand U9783 (N_9783,N_5314,N_7086);
nor U9784 (N_9784,N_6624,N_6108);
or U9785 (N_9785,N_5501,N_6509);
and U9786 (N_9786,N_5982,N_6096);
nand U9787 (N_9787,N_6836,N_6761);
nor U9788 (N_9788,N_7366,N_7153);
nand U9789 (N_9789,N_6202,N_7459);
and U9790 (N_9790,N_5169,N_6338);
nor U9791 (N_9791,N_6919,N_6029);
or U9792 (N_9792,N_5316,N_6681);
nor U9793 (N_9793,N_5937,N_7186);
nor U9794 (N_9794,N_5270,N_7336);
nand U9795 (N_9795,N_6797,N_6981);
and U9796 (N_9796,N_7487,N_7049);
and U9797 (N_9797,N_5543,N_5156);
or U9798 (N_9798,N_6558,N_7202);
or U9799 (N_9799,N_7096,N_6261);
nand U9800 (N_9800,N_5833,N_7019);
nand U9801 (N_9801,N_5786,N_5451);
or U9802 (N_9802,N_6212,N_5772);
nand U9803 (N_9803,N_7290,N_6513);
and U9804 (N_9804,N_5679,N_6622);
nor U9805 (N_9805,N_5415,N_5827);
nand U9806 (N_9806,N_5391,N_5204);
nor U9807 (N_9807,N_6170,N_6068);
nor U9808 (N_9808,N_7483,N_5379);
and U9809 (N_9809,N_7028,N_6470);
and U9810 (N_9810,N_5907,N_6124);
and U9811 (N_9811,N_6893,N_7001);
and U9812 (N_9812,N_6065,N_7495);
nor U9813 (N_9813,N_6549,N_5036);
nand U9814 (N_9814,N_6437,N_6238);
nor U9815 (N_9815,N_6641,N_6416);
nand U9816 (N_9816,N_6013,N_6437);
nand U9817 (N_9817,N_6333,N_5684);
nand U9818 (N_9818,N_5231,N_7480);
nor U9819 (N_9819,N_7287,N_6550);
or U9820 (N_9820,N_6753,N_5432);
nand U9821 (N_9821,N_5651,N_6760);
and U9822 (N_9822,N_6725,N_7413);
nor U9823 (N_9823,N_6937,N_5979);
and U9824 (N_9824,N_6004,N_7420);
nand U9825 (N_9825,N_5209,N_6893);
nor U9826 (N_9826,N_6420,N_7104);
nand U9827 (N_9827,N_5673,N_5913);
and U9828 (N_9828,N_6253,N_6441);
nand U9829 (N_9829,N_5270,N_6205);
nor U9830 (N_9830,N_6731,N_6332);
nand U9831 (N_9831,N_5405,N_5666);
or U9832 (N_9832,N_5334,N_5535);
and U9833 (N_9833,N_7361,N_7464);
nand U9834 (N_9834,N_5973,N_5388);
nand U9835 (N_9835,N_6961,N_6652);
or U9836 (N_9836,N_5634,N_6251);
or U9837 (N_9837,N_5243,N_6588);
or U9838 (N_9838,N_6512,N_6693);
xor U9839 (N_9839,N_5094,N_5195);
nor U9840 (N_9840,N_6604,N_7146);
or U9841 (N_9841,N_5929,N_6633);
nor U9842 (N_9842,N_5275,N_5413);
or U9843 (N_9843,N_6777,N_6549);
nand U9844 (N_9844,N_6807,N_6741);
or U9845 (N_9845,N_5453,N_7056);
and U9846 (N_9846,N_5027,N_5322);
and U9847 (N_9847,N_5637,N_5336);
or U9848 (N_9848,N_5687,N_5369);
nand U9849 (N_9849,N_6723,N_6481);
or U9850 (N_9850,N_6622,N_5920);
or U9851 (N_9851,N_6757,N_6194);
or U9852 (N_9852,N_5414,N_7207);
nand U9853 (N_9853,N_5933,N_5342);
nor U9854 (N_9854,N_5419,N_6987);
and U9855 (N_9855,N_7340,N_7466);
and U9856 (N_9856,N_5075,N_6553);
or U9857 (N_9857,N_7224,N_6888);
nor U9858 (N_9858,N_5128,N_6610);
nor U9859 (N_9859,N_6611,N_5839);
or U9860 (N_9860,N_7394,N_5993);
nand U9861 (N_9861,N_6040,N_7288);
or U9862 (N_9862,N_5477,N_7091);
or U9863 (N_9863,N_6993,N_7050);
or U9864 (N_9864,N_6114,N_6067);
nand U9865 (N_9865,N_5955,N_5848);
and U9866 (N_9866,N_5194,N_7122);
nand U9867 (N_9867,N_6075,N_6900);
nand U9868 (N_9868,N_7148,N_5570);
nor U9869 (N_9869,N_7391,N_5455);
and U9870 (N_9870,N_5460,N_6155);
or U9871 (N_9871,N_5021,N_6486);
nor U9872 (N_9872,N_7159,N_6260);
and U9873 (N_9873,N_5698,N_5237);
nor U9874 (N_9874,N_5329,N_7477);
and U9875 (N_9875,N_6839,N_5169);
or U9876 (N_9876,N_6883,N_7375);
nor U9877 (N_9877,N_5051,N_5346);
or U9878 (N_9878,N_5925,N_5273);
nand U9879 (N_9879,N_6974,N_6207);
nor U9880 (N_9880,N_5111,N_6570);
and U9881 (N_9881,N_5500,N_7295);
nor U9882 (N_9882,N_6514,N_5580);
nand U9883 (N_9883,N_5713,N_5791);
nand U9884 (N_9884,N_7044,N_6265);
and U9885 (N_9885,N_5804,N_6431);
or U9886 (N_9886,N_5663,N_6149);
and U9887 (N_9887,N_6277,N_6587);
and U9888 (N_9888,N_5790,N_6452);
and U9889 (N_9889,N_6632,N_5534);
and U9890 (N_9890,N_6393,N_5754);
and U9891 (N_9891,N_7083,N_7399);
nor U9892 (N_9892,N_5745,N_7360);
nand U9893 (N_9893,N_5774,N_7121);
xnor U9894 (N_9894,N_5177,N_5891);
or U9895 (N_9895,N_5558,N_6938);
or U9896 (N_9896,N_7418,N_6306);
and U9897 (N_9897,N_5980,N_6455);
and U9898 (N_9898,N_5086,N_5763);
nand U9899 (N_9899,N_6743,N_6295);
and U9900 (N_9900,N_5104,N_5008);
nor U9901 (N_9901,N_6817,N_5013);
and U9902 (N_9902,N_6895,N_7352);
nand U9903 (N_9903,N_6514,N_6605);
xnor U9904 (N_9904,N_5315,N_5706);
nor U9905 (N_9905,N_7048,N_6038);
nor U9906 (N_9906,N_7232,N_6238);
nor U9907 (N_9907,N_6174,N_5856);
or U9908 (N_9908,N_6529,N_6610);
nand U9909 (N_9909,N_6108,N_6405);
nor U9910 (N_9910,N_5351,N_6143);
or U9911 (N_9911,N_6488,N_7033);
nand U9912 (N_9912,N_6220,N_5750);
nand U9913 (N_9913,N_5925,N_5732);
and U9914 (N_9914,N_6366,N_6260);
or U9915 (N_9915,N_6802,N_6529);
nand U9916 (N_9916,N_6980,N_5803);
nor U9917 (N_9917,N_5875,N_7352);
or U9918 (N_9918,N_6191,N_5147);
nor U9919 (N_9919,N_6641,N_5312);
nor U9920 (N_9920,N_5139,N_5202);
nand U9921 (N_9921,N_6167,N_6899);
and U9922 (N_9922,N_6322,N_6701);
and U9923 (N_9923,N_5275,N_5740);
and U9924 (N_9924,N_7466,N_6160);
nor U9925 (N_9925,N_5043,N_5330);
and U9926 (N_9926,N_5752,N_5135);
or U9927 (N_9927,N_5300,N_6449);
nand U9928 (N_9928,N_5301,N_6071);
and U9929 (N_9929,N_7432,N_5832);
xnor U9930 (N_9930,N_6336,N_6326);
nand U9931 (N_9931,N_7046,N_6488);
or U9932 (N_9932,N_7015,N_7247);
or U9933 (N_9933,N_6963,N_6437);
or U9934 (N_9934,N_6562,N_6725);
nand U9935 (N_9935,N_5154,N_7408);
nand U9936 (N_9936,N_5941,N_6812);
or U9937 (N_9937,N_6518,N_5928);
nand U9938 (N_9938,N_5513,N_5964);
nand U9939 (N_9939,N_7058,N_5695);
or U9940 (N_9940,N_6511,N_6435);
xnor U9941 (N_9941,N_6199,N_5899);
or U9942 (N_9942,N_5105,N_6388);
and U9943 (N_9943,N_7064,N_5633);
nor U9944 (N_9944,N_5648,N_6189);
nand U9945 (N_9945,N_5617,N_7261);
or U9946 (N_9946,N_5173,N_6932);
and U9947 (N_9947,N_6050,N_6734);
nor U9948 (N_9948,N_5542,N_7466);
nand U9949 (N_9949,N_7307,N_7476);
or U9950 (N_9950,N_5155,N_6169);
or U9951 (N_9951,N_7459,N_6941);
nor U9952 (N_9952,N_6122,N_7388);
nand U9953 (N_9953,N_6346,N_5239);
nor U9954 (N_9954,N_6407,N_5892);
or U9955 (N_9955,N_6393,N_6385);
and U9956 (N_9956,N_5206,N_5090);
nand U9957 (N_9957,N_5847,N_5933);
nor U9958 (N_9958,N_6347,N_6811);
or U9959 (N_9959,N_6989,N_5345);
or U9960 (N_9960,N_7050,N_7387);
nor U9961 (N_9961,N_6464,N_5574);
or U9962 (N_9962,N_6978,N_7085);
nand U9963 (N_9963,N_6885,N_6525);
nor U9964 (N_9964,N_5646,N_5857);
nor U9965 (N_9965,N_7465,N_5580);
or U9966 (N_9966,N_5005,N_5012);
and U9967 (N_9967,N_5716,N_5232);
xor U9968 (N_9968,N_5236,N_6606);
nand U9969 (N_9969,N_5707,N_7317);
nand U9970 (N_9970,N_6806,N_7444);
or U9971 (N_9971,N_5285,N_5394);
nand U9972 (N_9972,N_6933,N_5180);
nor U9973 (N_9973,N_6251,N_6489);
and U9974 (N_9974,N_5738,N_6103);
or U9975 (N_9975,N_7355,N_5688);
and U9976 (N_9976,N_5566,N_7257);
and U9977 (N_9977,N_6201,N_6637);
or U9978 (N_9978,N_6409,N_7274);
nand U9979 (N_9979,N_5140,N_6628);
or U9980 (N_9980,N_5430,N_7307);
xnor U9981 (N_9981,N_5162,N_5659);
nor U9982 (N_9982,N_6141,N_5823);
nor U9983 (N_9983,N_6168,N_5845);
and U9984 (N_9984,N_6774,N_7138);
nand U9985 (N_9985,N_6937,N_5417);
and U9986 (N_9986,N_6258,N_6836);
nor U9987 (N_9987,N_5257,N_6447);
and U9988 (N_9988,N_6946,N_6241);
or U9989 (N_9989,N_5178,N_6383);
and U9990 (N_9990,N_5897,N_5452);
or U9991 (N_9991,N_6659,N_6851);
nand U9992 (N_9992,N_7465,N_7071);
nor U9993 (N_9993,N_6830,N_7209);
and U9994 (N_9994,N_6364,N_6686);
or U9995 (N_9995,N_5356,N_6857);
nand U9996 (N_9996,N_6167,N_5852);
and U9997 (N_9997,N_6032,N_5722);
nand U9998 (N_9998,N_5934,N_5579);
nor U9999 (N_9999,N_5896,N_5104);
and UO_0 (O_0,N_8063,N_7894);
or UO_1 (O_1,N_8065,N_7622);
or UO_2 (O_2,N_8694,N_9818);
nor UO_3 (O_3,N_8992,N_8335);
nand UO_4 (O_4,N_9374,N_9475);
nor UO_5 (O_5,N_7679,N_8200);
or UO_6 (O_6,N_8687,N_9408);
or UO_7 (O_7,N_8744,N_8933);
nor UO_8 (O_8,N_9875,N_9953);
and UO_9 (O_9,N_7658,N_8984);
nand UO_10 (O_10,N_9621,N_9486);
or UO_11 (O_11,N_9306,N_8237);
nor UO_12 (O_12,N_7578,N_9186);
or UO_13 (O_13,N_7627,N_8565);
and UO_14 (O_14,N_8569,N_7870);
nand UO_15 (O_15,N_9791,N_7808);
nand UO_16 (O_16,N_9071,N_8963);
nor UO_17 (O_17,N_9582,N_7783);
nor UO_18 (O_18,N_8322,N_9078);
nor UO_19 (O_19,N_8231,N_9666);
and UO_20 (O_20,N_8124,N_8232);
or UO_21 (O_21,N_8360,N_9052);
or UO_22 (O_22,N_9042,N_7685);
nand UO_23 (O_23,N_8726,N_9131);
nand UO_24 (O_24,N_9377,N_9846);
nor UO_25 (O_25,N_9467,N_8855);
and UO_26 (O_26,N_9149,N_8594);
nor UO_27 (O_27,N_8716,N_8819);
nand UO_28 (O_28,N_8152,N_8284);
or UO_29 (O_29,N_8760,N_7589);
nand UO_30 (O_30,N_9676,N_7601);
or UO_31 (O_31,N_8078,N_7820);
nand UO_32 (O_32,N_9570,N_9119);
nor UO_33 (O_33,N_7941,N_9358);
nor UO_34 (O_34,N_9389,N_7912);
or UO_35 (O_35,N_8737,N_9593);
and UO_36 (O_36,N_8466,N_7514);
or UO_37 (O_37,N_7836,N_7969);
and UO_38 (O_38,N_9060,N_8584);
and UO_39 (O_39,N_8048,N_8325);
nand UO_40 (O_40,N_7799,N_9223);
or UO_41 (O_41,N_9166,N_7961);
nor UO_42 (O_42,N_9103,N_9277);
nand UO_43 (O_43,N_8538,N_9949);
and UO_44 (O_44,N_8923,N_9877);
nor UO_45 (O_45,N_9120,N_7876);
or UO_46 (O_46,N_8457,N_9817);
nor UO_47 (O_47,N_9511,N_9733);
nand UO_48 (O_48,N_9347,N_8695);
and UO_49 (O_49,N_8862,N_9375);
nor UO_50 (O_50,N_9940,N_7992);
nand UO_51 (O_51,N_8488,N_7551);
nor UO_52 (O_52,N_9941,N_8648);
or UO_53 (O_53,N_9616,N_8709);
or UO_54 (O_54,N_9501,N_9221);
nor UO_55 (O_55,N_9516,N_9528);
or UO_56 (O_56,N_9418,N_9252);
nor UO_57 (O_57,N_9228,N_9710);
and UO_58 (O_58,N_9689,N_9019);
nor UO_59 (O_59,N_8261,N_8899);
nor UO_60 (O_60,N_7748,N_9836);
and UO_61 (O_61,N_8921,N_9450);
nand UO_62 (O_62,N_8874,N_8574);
and UO_63 (O_63,N_9635,N_9133);
nor UO_64 (O_64,N_9038,N_8292);
and UO_65 (O_65,N_8494,N_9830);
nor UO_66 (O_66,N_9414,N_9681);
or UO_67 (O_67,N_9719,N_8970);
nor UO_68 (O_68,N_8945,N_7756);
and UO_69 (O_69,N_9466,N_9843);
and UO_70 (O_70,N_9327,N_8712);
nand UO_71 (O_71,N_9139,N_8668);
and UO_72 (O_72,N_8402,N_9683);
or UO_73 (O_73,N_8363,N_9432);
or UO_74 (O_74,N_8293,N_8591);
nor UO_75 (O_75,N_9023,N_9271);
or UO_76 (O_76,N_8980,N_9145);
nor UO_77 (O_77,N_8789,N_8551);
nand UO_78 (O_78,N_7867,N_8122);
nand UO_79 (O_79,N_8143,N_8479);
and UO_80 (O_80,N_8435,N_9615);
or UO_81 (O_81,N_7991,N_9290);
nand UO_82 (O_82,N_8739,N_9455);
nor UO_83 (O_83,N_8442,N_9617);
nand UO_84 (O_84,N_9015,N_9054);
and UO_85 (O_85,N_8334,N_8663);
and UO_86 (O_86,N_9100,N_9239);
and UO_87 (O_87,N_9045,N_9317);
nor UO_88 (O_88,N_9735,N_9481);
or UO_89 (O_89,N_9315,N_8462);
or UO_90 (O_90,N_9938,N_8740);
and UO_91 (O_91,N_7529,N_8405);
and UO_92 (O_92,N_8978,N_8699);
nand UO_93 (O_93,N_8509,N_9955);
and UO_94 (O_94,N_9628,N_8315);
nor UO_95 (O_95,N_7527,N_9208);
and UO_96 (O_96,N_9510,N_7678);
and UO_97 (O_97,N_8491,N_8164);
nor UO_98 (O_98,N_8635,N_9763);
and UO_99 (O_99,N_7895,N_8967);
nand UO_100 (O_100,N_9318,N_7648);
and UO_101 (O_101,N_7614,N_9902);
nor UO_102 (O_102,N_7777,N_9337);
nor UO_103 (O_103,N_8219,N_8428);
nor UO_104 (O_104,N_9709,N_9776);
nand UO_105 (O_105,N_9812,N_8421);
or UO_106 (O_106,N_8367,N_8725);
nand UO_107 (O_107,N_9744,N_8528);
or UO_108 (O_108,N_8066,N_9837);
or UO_109 (O_109,N_9831,N_8746);
nand UO_110 (O_110,N_9329,N_9227);
nor UO_111 (O_111,N_9438,N_8208);
nand UO_112 (O_112,N_8755,N_8041);
xnor UO_113 (O_113,N_7931,N_8424);
and UO_114 (O_114,N_8601,N_9793);
and UO_115 (O_115,N_8481,N_7811);
nor UO_116 (O_116,N_9077,N_9064);
or UO_117 (O_117,N_9099,N_9156);
nor UO_118 (O_118,N_8715,N_7821);
or UO_119 (O_119,N_8936,N_9947);
and UO_120 (O_120,N_9662,N_9323);
nor UO_121 (O_121,N_8043,N_8880);
or UO_122 (O_122,N_9013,N_9185);
and UO_123 (O_123,N_9063,N_9496);
and UO_124 (O_124,N_7520,N_7767);
xnor UO_125 (O_125,N_9310,N_9403);
nand UO_126 (O_126,N_8682,N_8900);
or UO_127 (O_127,N_7906,N_8643);
or UO_128 (O_128,N_8940,N_7759);
xor UO_129 (O_129,N_9820,N_8250);
nand UO_130 (O_130,N_9563,N_9611);
nand UO_131 (O_131,N_9933,N_9762);
nand UO_132 (O_132,N_9379,N_7638);
nand UO_133 (O_133,N_9581,N_9883);
or UO_134 (O_134,N_9730,N_9085);
and UO_135 (O_135,N_7615,N_8196);
nor UO_136 (O_136,N_8621,N_7850);
nor UO_137 (O_137,N_9380,N_9749);
or UO_138 (O_138,N_7889,N_9788);
or UO_139 (O_139,N_9264,N_9650);
or UO_140 (O_140,N_8800,N_8618);
and UO_141 (O_141,N_8177,N_9146);
and UO_142 (O_142,N_9586,N_8109);
or UO_143 (O_143,N_7965,N_7884);
or UO_144 (O_144,N_7878,N_7937);
or UO_145 (O_145,N_8414,N_9716);
or UO_146 (O_146,N_8954,N_7933);
nand UO_147 (O_147,N_8094,N_9661);
nand UO_148 (O_148,N_8696,N_9011);
nand UO_149 (O_149,N_9010,N_9974);
or UO_150 (O_150,N_8438,N_8542);
or UO_151 (O_151,N_8681,N_9360);
nand UO_152 (O_152,N_7893,N_9034);
or UO_153 (O_153,N_7932,N_8549);
and UO_154 (O_154,N_9321,N_8271);
or UO_155 (O_155,N_9936,N_9334);
nor UO_156 (O_156,N_8711,N_7818);
nand UO_157 (O_157,N_9012,N_8127);
nand UO_158 (O_158,N_9811,N_9035);
nor UO_159 (O_159,N_9459,N_7523);
nand UO_160 (O_160,N_8742,N_9538);
nand UO_161 (O_161,N_8516,N_8780);
or UO_162 (O_162,N_8974,N_8863);
and UO_163 (O_163,N_9652,N_8671);
nand UO_164 (O_164,N_8181,N_8782);
and UO_165 (O_165,N_8263,N_7797);
nor UO_166 (O_166,N_8689,N_9690);
and UO_167 (O_167,N_9755,N_9425);
nand UO_168 (O_168,N_8608,N_9111);
nand UO_169 (O_169,N_7812,N_8939);
nor UO_170 (O_170,N_9656,N_7944);
nand UO_171 (O_171,N_8805,N_8583);
nor UO_172 (O_172,N_9249,N_8020);
nor UO_173 (O_173,N_9216,N_9348);
nand UO_174 (O_174,N_7784,N_7707);
nor UO_175 (O_175,N_8257,N_7561);
and UO_176 (O_176,N_8074,N_8265);
and UO_177 (O_177,N_7504,N_8260);
nand UO_178 (O_178,N_7887,N_9961);
nor UO_179 (O_179,N_9922,N_9089);
nor UO_180 (O_180,N_7781,N_9598);
nand UO_181 (O_181,N_8297,N_8145);
nand UO_182 (O_182,N_9928,N_9853);
nor UO_183 (O_183,N_9796,N_9702);
nand UO_184 (O_184,N_8724,N_8114);
nor UO_185 (O_185,N_8501,N_7939);
and UO_186 (O_186,N_8326,N_9125);
and UO_187 (O_187,N_8485,N_8348);
nor UO_188 (O_188,N_9154,N_8330);
nor UO_189 (O_189,N_8318,N_7868);
or UO_190 (O_190,N_9738,N_8075);
or UO_191 (O_191,N_9394,N_8413);
nor UO_192 (O_192,N_9944,N_9578);
nor UO_193 (O_193,N_9000,N_8848);
nand UO_194 (O_194,N_7728,N_8469);
nand UO_195 (O_195,N_8607,N_7628);
or UO_196 (O_196,N_9766,N_8834);
and UO_197 (O_197,N_9498,N_8852);
and UO_198 (O_198,N_8323,N_9020);
and UO_199 (O_199,N_8988,N_7563);
and UO_200 (O_200,N_8387,N_9212);
and UO_201 (O_201,N_9913,N_8173);
and UO_202 (O_202,N_9189,N_9400);
and UO_203 (O_203,N_9905,N_9176);
nor UO_204 (O_204,N_8922,N_9887);
and UO_205 (O_205,N_8233,N_7579);
nor UO_206 (O_206,N_7660,N_7655);
nor UO_207 (O_207,N_8827,N_7830);
and UO_208 (O_208,N_8372,N_9230);
or UO_209 (O_209,N_8407,N_9285);
nor UO_210 (O_210,N_8294,N_8153);
and UO_211 (O_211,N_9959,N_8706);
or UO_212 (O_212,N_9781,N_8768);
or UO_213 (O_213,N_8818,N_8316);
nand UO_214 (O_214,N_9107,N_7843);
or UO_215 (O_215,N_9659,N_8487);
or UO_216 (O_216,N_7949,N_7831);
or UO_217 (O_217,N_8947,N_9967);
and UO_218 (O_218,N_7500,N_7719);
or UO_219 (O_219,N_8203,N_8759);
nand UO_220 (O_220,N_9471,N_9359);
or UO_221 (O_221,N_9059,N_7710);
and UO_222 (O_222,N_8956,N_9428);
nand UO_223 (O_223,N_8125,N_9211);
or UO_224 (O_224,N_8544,N_9219);
or UO_225 (O_225,N_9734,N_8129);
nand UO_226 (O_226,N_9646,N_9838);
or UO_227 (O_227,N_9622,N_9858);
nand UO_228 (O_228,N_7838,N_8167);
nand UO_229 (O_229,N_8082,N_9696);
and UO_230 (O_230,N_8580,N_9047);
nand UO_231 (O_231,N_7715,N_8866);
or UO_232 (O_232,N_9927,N_9200);
or UO_233 (O_233,N_8483,N_7851);
and UO_234 (O_234,N_7700,N_8439);
and UO_235 (O_235,N_7633,N_8459);
xor UO_236 (O_236,N_8680,N_9554);
or UO_237 (O_237,N_8812,N_8207);
and UO_238 (O_238,N_8704,N_8592);
nand UO_239 (O_239,N_8690,N_8398);
and UO_240 (O_240,N_7604,N_7858);
nand UO_241 (O_241,N_9660,N_7559);
and UO_242 (O_242,N_8342,N_9623);
and UO_243 (O_243,N_8385,N_7803);
and UO_244 (O_244,N_9888,N_9536);
nand UO_245 (O_245,N_9725,N_8588);
and UO_246 (O_246,N_8223,N_7856);
nand UO_247 (O_247,N_9302,N_8288);
nor UO_248 (O_248,N_7510,N_7524);
nand UO_249 (O_249,N_8926,N_8225);
nor UO_250 (O_250,N_7751,N_8530);
or UO_251 (O_251,N_9109,N_9405);
nand UO_252 (O_252,N_7652,N_9232);
and UO_253 (O_253,N_7620,N_8037);
and UO_254 (O_254,N_7846,N_8534);
nand UO_255 (O_255,N_9943,N_8981);
and UO_256 (O_256,N_7598,N_8305);
nor UO_257 (O_257,N_9457,N_8380);
nor UO_258 (O_258,N_8304,N_8341);
nor UO_259 (O_259,N_9748,N_8351);
or UO_260 (O_260,N_9409,N_9625);
nor UO_261 (O_261,N_8244,N_8313);
nand UO_262 (O_262,N_9672,N_9585);
and UO_263 (O_263,N_9421,N_9675);
nor UO_264 (O_264,N_7553,N_8099);
nand UO_265 (O_265,N_7888,N_8253);
or UO_266 (O_266,N_7824,N_8498);
and UO_267 (O_267,N_9787,N_9764);
nand UO_268 (O_268,N_9192,N_9021);
or UO_269 (O_269,N_9607,N_9647);
nand UO_270 (O_270,N_7522,N_8475);
nand UO_271 (O_271,N_8888,N_8526);
and UO_272 (O_272,N_9740,N_9053);
nor UO_273 (O_273,N_7706,N_8390);
nand UO_274 (O_274,N_8331,N_9491);
or UO_275 (O_275,N_7535,N_8273);
or UO_276 (O_276,N_8340,N_9859);
or UO_277 (O_277,N_7765,N_8660);
nor UO_278 (O_278,N_9392,N_9483);
nand UO_279 (O_279,N_8279,N_9378);
nand UO_280 (O_280,N_8070,N_7956);
nand UO_281 (O_281,N_7886,N_9182);
nor UO_282 (O_282,N_9284,N_8038);
nand UO_283 (O_283,N_9280,N_7834);
or UO_284 (O_284,N_8091,N_9544);
nand UO_285 (O_285,N_7692,N_9474);
and UO_286 (O_286,N_7792,N_8581);
or UO_287 (O_287,N_7671,N_8280);
nor UO_288 (O_288,N_9116,N_9644);
and UO_289 (O_289,N_9236,N_8803);
and UO_290 (O_290,N_7640,N_9911);
and UO_291 (O_291,N_7902,N_8731);
nand UO_292 (O_292,N_8040,N_9016);
xor UO_293 (O_293,N_9505,N_8238);
nand UO_294 (O_294,N_8134,N_9533);
or UO_295 (O_295,N_7605,N_8717);
and UO_296 (O_296,N_8393,N_9030);
and UO_297 (O_297,N_8461,N_7714);
and UO_298 (O_298,N_8850,N_8150);
xnor UO_299 (O_299,N_8087,N_8242);
or UO_300 (O_300,N_8832,N_9153);
nor UO_301 (O_301,N_7840,N_8444);
or UO_302 (O_302,N_8950,N_7985);
xor UO_303 (O_303,N_9934,N_8067);
nor UO_304 (O_304,N_8171,N_8505);
nor UO_305 (O_305,N_9143,N_7684);
and UO_306 (O_306,N_9760,N_9144);
nor UO_307 (O_307,N_9463,N_8560);
and UO_308 (O_308,N_9614,N_9092);
xnor UO_309 (O_309,N_9084,N_7924);
nor UO_310 (O_310,N_9365,N_8490);
or UO_311 (O_311,N_9398,N_7925);
or UO_312 (O_312,N_8473,N_8061);
nand UO_313 (O_313,N_9209,N_9476);
or UO_314 (O_314,N_7610,N_7546);
nand UO_315 (O_315,N_8376,N_9296);
or UO_316 (O_316,N_9415,N_7790);
nor UO_317 (O_317,N_9461,N_9448);
nor UO_318 (O_318,N_9259,N_8944);
nor UO_319 (O_319,N_8747,N_8112);
nand UO_320 (O_320,N_8670,N_9768);
or UO_321 (O_321,N_7786,N_9436);
or UO_322 (O_322,N_7871,N_9062);
or UO_323 (O_323,N_9799,N_8532);
and UO_324 (O_324,N_9383,N_8873);
or UO_325 (O_325,N_7753,N_8625);
and UO_326 (O_326,N_8707,N_8563);
nor UO_327 (O_327,N_7869,N_8350);
nor UO_328 (O_328,N_9196,N_9835);
xor UO_329 (O_329,N_8861,N_8364);
and UO_330 (O_330,N_7763,N_9619);
and UO_331 (O_331,N_8674,N_9178);
nor UO_332 (O_332,N_9565,N_9344);
and UO_333 (O_333,N_9798,N_8135);
or UO_334 (O_334,N_9736,N_8137);
and UO_335 (O_335,N_8904,N_9231);
nor UO_336 (O_336,N_7711,N_9839);
or UO_337 (O_337,N_9739,N_9433);
nand UO_338 (O_338,N_7810,N_8891);
or UO_339 (O_339,N_9371,N_7505);
nand UO_340 (O_340,N_8176,N_8932);
and UO_341 (O_341,N_8548,N_8266);
or UO_342 (O_342,N_7829,N_7518);
and UO_343 (O_343,N_9468,N_8142);
nor UO_344 (O_344,N_8269,N_9174);
or UO_345 (O_345,N_9564,N_7750);
or UO_346 (O_346,N_8011,N_8056);
and UO_347 (O_347,N_8986,N_9751);
or UO_348 (O_348,N_9566,N_8573);
nand UO_349 (O_349,N_7603,N_8779);
or UO_350 (O_350,N_8029,N_8394);
nor UO_351 (O_351,N_9345,N_7509);
nand UO_352 (O_352,N_8358,N_8039);
or UO_353 (O_353,N_8518,N_9822);
and UO_354 (O_354,N_9643,N_9849);
or UO_355 (O_355,N_8830,N_8352);
nand UO_356 (O_356,N_9477,N_8073);
nand UO_357 (O_357,N_9800,N_9539);
nor UO_358 (O_358,N_8286,N_9807);
and UO_359 (O_359,N_8738,N_8464);
and UO_360 (O_360,N_7915,N_8763);
or UO_361 (O_361,N_9750,N_7882);
and UO_362 (O_362,N_8741,N_8191);
or UO_363 (O_363,N_8282,N_8554);
nor UO_364 (O_364,N_8254,N_7929);
nand UO_365 (O_365,N_9703,N_8034);
or UO_366 (O_366,N_7913,N_7801);
nand UO_367 (O_367,N_7727,N_7754);
nand UO_368 (O_368,N_9233,N_8778);
and UO_369 (O_369,N_9898,N_7585);
or UO_370 (O_370,N_8985,N_7896);
nor UO_371 (O_371,N_8968,N_9523);
nand UO_372 (O_372,N_8001,N_7974);
or UO_373 (O_373,N_8131,N_9097);
nand UO_374 (O_374,N_8605,N_7990);
and UO_375 (O_375,N_9583,N_7789);
or UO_376 (O_376,N_7681,N_8199);
nor UO_377 (O_377,N_9485,N_9832);
nor UO_378 (O_378,N_9269,N_9330);
or UO_379 (O_379,N_7570,N_8033);
nand UO_380 (O_380,N_9235,N_9048);
and UO_381 (O_381,N_9803,N_9439);
and UO_382 (O_382,N_8907,N_8121);
and UO_383 (O_383,N_8453,N_8373);
nor UO_384 (O_384,N_8912,N_8400);
and UO_385 (O_385,N_9074,N_8147);
nor UO_386 (O_386,N_7699,N_9279);
or UO_387 (O_387,N_8628,N_8116);
and UO_388 (O_388,N_7542,N_8432);
and UO_389 (O_389,N_8669,N_8541);
or UO_390 (O_390,N_9805,N_8226);
nand UO_391 (O_391,N_8951,N_7676);
or UO_392 (O_392,N_9075,N_8519);
nand UO_393 (O_393,N_8084,N_8566);
or UO_394 (O_394,N_9923,N_9322);
or UO_395 (O_395,N_7623,N_8013);
or UO_396 (O_396,N_8440,N_8991);
or UO_397 (O_397,N_8126,N_7972);
or UO_398 (O_398,N_8357,N_8813);
and UO_399 (O_399,N_7511,N_8183);
nor UO_400 (O_400,N_8302,N_7764);
nor UO_401 (O_401,N_8536,N_8411);
and UO_402 (O_402,N_9618,N_7650);
nor UO_403 (O_403,N_7634,N_9994);
or UO_404 (O_404,N_7732,N_9281);
and UO_405 (O_405,N_8570,N_9663);
and UO_406 (O_406,N_9188,N_8044);
nor UO_407 (O_407,N_8193,N_9728);
nor UO_408 (O_408,N_8030,N_8616);
and UO_409 (O_409,N_9518,N_9606);
nor UO_410 (O_410,N_8182,N_7586);
and UO_411 (O_411,N_9390,N_9878);
or UO_412 (O_412,N_9568,N_9545);
and UO_413 (O_413,N_9790,N_9134);
nand UO_414 (O_414,N_9896,N_9901);
nand UO_415 (O_415,N_9605,N_8148);
nor UO_416 (O_416,N_9283,N_7668);
nor UO_417 (O_417,N_9863,N_9856);
or UO_418 (O_418,N_7743,N_8369);
nor UO_419 (O_419,N_7530,N_8086);
nand UO_420 (O_420,N_8274,N_7901);
nand UO_421 (O_421,N_9980,N_8977);
nor UO_422 (O_422,N_9458,N_9699);
nand UO_423 (O_423,N_8942,N_9043);
nand UO_424 (O_424,N_7900,N_8027);
nor UO_425 (O_425,N_7861,N_8419);
nand UO_426 (O_426,N_8686,N_8645);
nor UO_427 (O_427,N_9915,N_8692);
nand UO_428 (O_428,N_7568,N_8068);
and UO_429 (O_429,N_8529,N_8816);
and UO_430 (O_430,N_8587,N_9292);
nand UO_431 (O_431,N_8777,N_8615);
nor UO_432 (O_432,N_9478,N_9987);
nand UO_433 (O_433,N_9324,N_9624);
nand UO_434 (O_434,N_9789,N_7675);
and UO_435 (O_435,N_9254,N_8764);
and UO_436 (O_436,N_8258,N_9293);
or UO_437 (O_437,N_8194,N_8093);
or UO_438 (O_438,N_9363,N_9309);
or UO_439 (O_439,N_8051,N_9535);
nand UO_440 (O_440,N_7556,N_7807);
or UO_441 (O_441,N_7921,N_9976);
and UO_442 (O_442,N_9112,N_8654);
nand UO_443 (O_443,N_9253,N_9155);
and UO_444 (O_444,N_7964,N_9350);
nor UO_445 (O_445,N_9008,N_9427);
and UO_446 (O_446,N_8287,N_9833);
or UO_447 (O_447,N_9319,N_8661);
or UO_448 (O_448,N_7892,N_8938);
nor UO_449 (O_449,N_8826,N_8336);
nor UO_450 (O_450,N_8730,N_9198);
and UO_451 (O_451,N_9180,N_8090);
nor UO_452 (O_452,N_8644,N_9199);
or UO_453 (O_453,N_7537,N_7508);
or UO_454 (O_454,N_9096,N_8965);
nor UO_455 (O_455,N_9066,N_7928);
nand UO_456 (O_456,N_8221,N_7963);
nand UO_457 (O_457,N_7664,N_7945);
or UO_458 (O_458,N_8308,N_8512);
or UO_459 (O_459,N_9695,N_7955);
nand UO_460 (O_460,N_7629,N_8290);
nor UO_461 (O_461,N_8455,N_8829);
nor UO_462 (O_462,N_9367,N_9509);
nand UO_463 (O_463,N_7866,N_9720);
or UO_464 (O_464,N_8338,N_8166);
nor UO_465 (O_465,N_9680,N_8750);
nand UO_466 (O_466,N_7547,N_9669);
and UO_467 (O_467,N_8019,N_7890);
nor UO_468 (O_468,N_8211,N_8514);
nor UO_469 (O_469,N_7722,N_9452);
and UO_470 (O_470,N_9993,N_9256);
nor UO_471 (O_471,N_9308,N_8748);
and UO_472 (O_472,N_8130,N_8558);
nand UO_473 (O_473,N_8713,N_7762);
nand UO_474 (O_474,N_8408,N_9816);
nor UO_475 (O_475,N_8396,N_7999);
or UO_476 (O_476,N_8571,N_9828);
or UO_477 (O_477,N_9288,N_8362);
and UO_478 (O_478,N_9207,N_9385);
and UO_479 (O_479,N_8141,N_8477);
and UO_480 (O_480,N_9640,N_9774);
nand UO_481 (O_481,N_8997,N_7857);
nor UO_482 (O_482,N_8049,N_7636);
nor UO_483 (O_483,N_9885,N_7845);
or UO_484 (O_484,N_9912,N_8215);
nor UO_485 (O_485,N_8454,N_8427);
nand UO_486 (O_486,N_9775,N_8655);
and UO_487 (O_487,N_9999,N_9827);
xor UO_488 (O_488,N_7864,N_8468);
nand UO_489 (O_489,N_8420,N_8452);
nor UO_490 (O_490,N_9782,N_8911);
and UO_491 (O_491,N_9704,N_7800);
nand UO_492 (O_492,N_7672,N_8417);
and UO_493 (O_493,N_7959,N_9294);
or UO_494 (O_494,N_7823,N_8597);
and UO_495 (O_495,N_9594,N_9924);
or UO_496 (O_496,N_7981,N_7690);
nor UO_497 (O_497,N_8157,N_8321);
nand UO_498 (O_498,N_9921,N_8783);
nor UO_499 (O_499,N_7539,N_7769);
nor UO_500 (O_500,N_8893,N_9592);
or UO_501 (O_501,N_9470,N_9401);
or UO_502 (O_502,N_7874,N_9102);
nand UO_503 (O_503,N_8267,N_8599);
and UO_504 (O_504,N_7986,N_8472);
nor UO_505 (O_505,N_8179,N_7554);
or UO_506 (O_506,N_8235,N_9270);
nor UO_507 (O_507,N_9201,N_8214);
nand UO_508 (O_508,N_9027,N_8784);
nand UO_509 (O_509,N_8032,N_9537);
and UO_510 (O_510,N_9167,N_9642);
nand UO_511 (O_511,N_7595,N_9958);
or UO_512 (O_512,N_9861,N_8636);
nor UO_513 (O_513,N_8788,N_8898);
and UO_514 (O_514,N_7687,N_8929);
or UO_515 (O_515,N_9808,N_9022);
and UO_516 (O_516,N_9164,N_9806);
nor UO_517 (O_517,N_9229,N_8016);
nor UO_518 (O_518,N_7538,N_9772);
and UO_519 (O_519,N_9173,N_9331);
nor UO_520 (O_520,N_8025,N_7651);
and UO_521 (O_521,N_8720,N_9694);
and UO_522 (O_522,N_8241,N_9834);
or UO_523 (O_523,N_9651,N_8773);
nor UO_524 (O_524,N_8971,N_8679);
nor UO_525 (O_525,N_7766,N_9504);
and UO_526 (O_526,N_7976,N_8328);
or UO_527 (O_527,N_7839,N_8517);
nand UO_528 (O_528,N_8089,N_8224);
or UO_529 (O_529,N_9968,N_8953);
nand UO_530 (O_530,N_7562,N_8678);
or UO_531 (O_531,N_9090,N_8892);
nand UO_532 (O_532,N_9124,N_9426);
or UO_533 (O_533,N_9964,N_8397);
nor UO_534 (O_534,N_8356,N_9101);
or UO_535 (O_535,N_9333,N_9316);
and UO_536 (O_536,N_9892,N_9441);
nand UO_537 (O_537,N_9658,N_8492);
and UO_538 (O_538,N_8955,N_8418);
nand UO_539 (O_539,N_9514,N_9655);
or UO_540 (O_540,N_9397,N_8117);
xor UO_541 (O_541,N_9829,N_8354);
nor UO_542 (O_542,N_8064,N_8353);
or UO_543 (O_543,N_7590,N_9341);
nand UO_544 (O_544,N_7733,N_9711);
or UO_545 (O_545,N_9971,N_9747);
and UO_546 (O_546,N_9984,N_7742);
or UO_547 (O_547,N_9499,N_7593);
and UO_548 (O_548,N_9722,N_8450);
nor UO_549 (O_549,N_9261,N_9900);
nand UO_550 (O_550,N_9464,N_8349);
nor UO_551 (O_551,N_8540,N_8876);
and UO_552 (O_552,N_9036,N_9840);
nand UO_553 (O_553,N_9295,N_7770);
nand UO_554 (O_554,N_7689,N_8482);
nor UO_555 (O_555,N_8794,N_8698);
nor UO_556 (O_556,N_7534,N_9110);
nand UO_557 (O_557,N_8620,N_9982);
nor UO_558 (O_558,N_9416,N_8662);
nor UO_559 (O_559,N_9532,N_7952);
or UO_560 (O_560,N_9244,N_7521);
and UO_561 (O_561,N_9287,N_9274);
nor UO_562 (O_562,N_9141,N_7596);
nor UO_563 (O_563,N_9783,N_8406);
nor UO_564 (O_564,N_8856,N_8787);
nand UO_565 (O_565,N_7677,N_8104);
nand UO_566 (O_566,N_8161,N_7814);
nand UO_567 (O_567,N_9918,N_7573);
nand UO_568 (O_568,N_9298,N_9242);
and UO_569 (O_569,N_7611,N_7680);
and UO_570 (O_570,N_9848,N_9353);
nand UO_571 (O_571,N_9419,N_8486);
and UO_572 (O_572,N_7988,N_8676);
and UO_573 (O_573,N_7854,N_8769);
or UO_574 (O_574,N_9445,N_8295);
nor UO_575 (O_575,N_8825,N_7825);
or UO_576 (O_576,N_8872,N_7572);
or UO_577 (O_577,N_8310,N_9079);
or UO_578 (O_578,N_8600,N_8913);
or UO_579 (O_579,N_9600,N_8256);
and UO_580 (O_580,N_8003,N_7872);
and UO_581 (O_581,N_9714,N_9780);
or UO_582 (O_582,N_8456,N_7798);
or UO_583 (O_583,N_9558,N_7599);
or UO_584 (O_584,N_9108,N_8300);
nand UO_585 (O_585,N_8887,N_8202);
nor UO_586 (O_586,N_9919,N_8626);
nor UO_587 (O_587,N_8236,N_8537);
nor UO_588 (O_588,N_8379,N_7934);
and UO_589 (O_589,N_9263,N_7507);
and UO_590 (O_590,N_9051,N_7855);
and UO_591 (O_591,N_7935,N_9991);
and UO_592 (O_592,N_8885,N_8995);
or UO_593 (O_593,N_8213,N_8586);
nand UO_594 (O_594,N_9275,N_9773);
and UO_595 (O_595,N_8753,N_8010);
nor UO_596 (O_596,N_7755,N_7989);
or UO_597 (O_597,N_9257,N_9524);
nor UO_598 (O_598,N_8579,N_8650);
or UO_599 (O_599,N_8404,N_8053);
and UO_600 (O_600,N_9444,N_9810);
or UO_601 (O_601,N_9983,N_7778);
or UO_602 (O_602,N_7607,N_9429);
nor UO_603 (O_603,N_8503,N_8697);
or UO_604 (O_604,N_8535,N_8701);
or UO_605 (O_605,N_9992,N_8189);
nor UO_606 (O_606,N_8395,N_8602);
and UO_607 (O_607,N_8433,N_8727);
or UO_608 (O_608,N_9930,N_9797);
nor UO_609 (O_609,N_9404,N_9866);
or UO_610 (O_610,N_9137,N_9114);
and UO_611 (O_611,N_9639,N_7583);
and UO_612 (O_612,N_7809,N_8867);
nand UO_613 (O_613,N_8205,N_9721);
xnor UO_614 (O_614,N_9962,N_9098);
or UO_615 (O_615,N_8774,N_7993);
nand UO_616 (O_616,N_8843,N_9884);
nor UO_617 (O_617,N_9815,N_8489);
or UO_618 (O_618,N_8798,N_8632);
and UO_619 (O_619,N_8772,N_8743);
or UO_620 (O_620,N_9894,N_8262);
and UO_621 (O_621,N_7501,N_8658);
nor UO_622 (O_622,N_9028,N_8637);
or UO_623 (O_623,N_8054,N_9777);
or UO_624 (O_624,N_8790,N_8667);
nor UO_625 (O_625,N_8734,N_8903);
and UO_626 (O_626,N_7709,N_8631);
nand UO_627 (O_627,N_9431,N_8268);
nand UO_628 (O_628,N_9396,N_8999);
or UO_629 (O_629,N_9058,N_8799);
nor UO_630 (O_630,N_9248,N_7758);
or UO_631 (O_631,N_9550,N_8555);
or UO_632 (O_632,N_7815,N_9368);
nor UO_633 (O_633,N_9677,N_9931);
and UO_634 (O_634,N_8836,N_9869);
or UO_635 (O_635,N_7922,N_9920);
nand UO_636 (O_636,N_8508,N_8909);
and UO_637 (O_637,N_9771,N_8460);
and UO_638 (O_638,N_8480,N_9472);
nor UO_639 (O_639,N_9487,N_7973);
nor UO_640 (O_640,N_9948,N_9343);
nand UO_641 (O_641,N_9479,N_8144);
nand UO_642 (O_642,N_9700,N_8277);
nand UO_643 (O_643,N_8809,N_7806);
nor UO_644 (O_644,N_8014,N_9332);
nor UO_645 (O_645,N_7844,N_9026);
and UO_646 (O_646,N_9094,N_8841);
and UO_647 (O_647,N_8429,N_9217);
nor UO_648 (O_648,N_7536,N_8659);
nor UO_649 (O_649,N_9105,N_8128);
nand UO_650 (O_650,N_7639,N_9506);
and UO_651 (O_651,N_8627,N_8355);
and UO_652 (O_652,N_7662,N_8785);
nor UO_653 (O_653,N_8722,N_8878);
nor UO_654 (O_654,N_7597,N_9526);
nand UO_655 (O_655,N_9613,N_8415);
or UO_656 (O_656,N_9190,N_7739);
nand UO_657 (O_657,N_9266,N_9399);
and UO_658 (O_658,N_8821,N_8299);
nand UO_659 (O_659,N_8546,N_9304);
and UO_660 (O_660,N_9088,N_9946);
and UO_661 (O_661,N_7950,N_9033);
and UO_662 (O_662,N_8507,N_7517);
nor UO_663 (O_663,N_9040,N_9142);
or UO_664 (O_664,N_8881,N_9183);
or UO_665 (O_665,N_7904,N_8705);
and UO_666 (O_666,N_9165,N_8745);
or UO_667 (O_667,N_9687,N_7665);
nand UO_668 (O_668,N_8639,N_7667);
nor UO_669 (O_669,N_9597,N_8814);
and UO_670 (O_670,N_9851,N_8470);
and UO_671 (O_671,N_8426,N_8613);
and UO_672 (O_672,N_8877,N_9451);
and UO_673 (O_673,N_8212,N_9135);
nor UO_674 (O_674,N_9195,N_8564);
nand UO_675 (O_675,N_8103,N_9130);
or UO_676 (O_676,N_9841,N_9726);
and UO_677 (O_677,N_8500,N_7659);
nand UO_678 (O_678,N_8675,N_9202);
or UO_679 (O_679,N_8666,N_9645);
nor UO_680 (O_680,N_8844,N_7978);
or UO_681 (O_681,N_9073,N_7621);
or UO_682 (O_682,N_9197,N_7567);
nand UO_683 (O_683,N_8108,N_8657);
or UO_684 (O_684,N_7757,N_7788);
nor UO_685 (O_685,N_9328,N_9245);
or UO_686 (O_686,N_9925,N_9630);
or UO_687 (O_687,N_8531,N_8969);
nand UO_688 (O_688,N_8307,N_9589);
or UO_689 (O_689,N_8243,N_9494);
or UO_690 (O_690,N_9002,N_7772);
nand UO_691 (O_691,N_9006,N_9260);
nor UO_692 (O_692,N_8197,N_8311);
nor UO_693 (O_693,N_9599,N_8218);
nand UO_694 (O_694,N_9588,N_8374);
nor UO_695 (O_695,N_7649,N_8045);
nor UO_696 (O_696,N_8239,N_8810);
and UO_697 (O_697,N_8102,N_9147);
or UO_698 (O_698,N_7909,N_8522);
nor UO_699 (O_699,N_7847,N_8998);
and UO_700 (O_700,N_8624,N_9081);
nand UO_701 (O_701,N_8329,N_9080);
nand UO_702 (O_702,N_9286,N_7533);
nor UO_703 (O_703,N_9705,N_8007);
and UO_704 (O_704,N_8240,N_8653);
and UO_705 (O_705,N_9688,N_8860);
and UO_706 (O_706,N_8875,N_9384);
and UO_707 (O_707,N_8806,N_8327);
nor UO_708 (O_708,N_7670,N_8092);
nand UO_709 (O_709,N_7975,N_8762);
nand UO_710 (O_710,N_9276,N_8864);
and UO_711 (O_711,N_8765,N_8736);
nor UO_712 (O_712,N_9157,N_9854);
nor UO_713 (O_713,N_9692,N_7582);
nand UO_714 (O_714,N_9674,N_9864);
or UO_715 (O_715,N_8797,N_9954);
or UO_716 (O_716,N_9671,N_8733);
nand UO_717 (O_717,N_7723,N_9126);
or UO_718 (O_718,N_8412,N_9148);
or UO_719 (O_719,N_9778,N_7606);
or UO_720 (O_720,N_8416,N_8448);
nor UO_721 (O_721,N_8975,N_9272);
or UO_722 (O_722,N_9161,N_7571);
and UO_723 (O_723,N_7673,N_9932);
nor UO_724 (O_724,N_9017,N_7828);
nor UO_725 (O_725,N_7897,N_8050);
or UO_726 (O_726,N_7713,N_8081);
or UO_727 (O_727,N_7575,N_8210);
nand UO_728 (O_728,N_9447,N_9203);
nand UO_729 (O_729,N_7908,N_8732);
nor UO_730 (O_730,N_7644,N_8533);
nor UO_731 (O_731,N_9070,N_9880);
nand UO_732 (O_732,N_9068,N_8609);
or UO_733 (O_733,N_8155,N_7940);
or UO_734 (O_734,N_9779,N_8952);
nand UO_735 (O_735,N_9123,N_7849);
or UO_736 (O_736,N_9372,N_8506);
and UO_737 (O_737,N_8185,N_8008);
or UO_738 (O_738,N_9852,N_8723);
and UO_739 (O_739,N_8664,N_9627);
nand UO_740 (O_740,N_9929,N_8920);
nand UO_741 (O_741,N_8527,N_8343);
nand UO_742 (O_742,N_8031,N_7503);
nand UO_743 (O_743,N_8410,N_7626);
nor UO_744 (O_744,N_7608,N_9179);
and UO_745 (O_745,N_8935,N_9547);
nor UO_746 (O_746,N_8633,N_8757);
nand UO_747 (O_747,N_7780,N_9342);
nor UO_748 (O_748,N_9879,N_8976);
or UO_749 (O_749,N_9957,N_9845);
nor UO_750 (O_750,N_8817,N_8022);
nand UO_751 (O_751,N_9443,N_9795);
or UO_752 (O_752,N_9939,N_8392);
and UO_753 (O_753,N_9193,N_9729);
or UO_754 (O_754,N_8309,N_8917);
or UO_755 (O_755,N_7737,N_9897);
and UO_756 (O_756,N_8002,N_8919);
and UO_757 (O_757,N_7880,N_9802);
nand UO_758 (O_758,N_7749,N_9267);
nand UO_759 (O_759,N_9460,N_9713);
and UO_760 (O_760,N_8296,N_8553);
and UO_761 (O_761,N_8312,N_7995);
nand UO_762 (O_762,N_7705,N_8383);
and UO_763 (O_763,N_9632,N_9065);
nor UO_764 (O_764,N_9278,N_9517);
nor UO_765 (O_765,N_9813,N_7744);
nor UO_766 (O_766,N_9576,N_9819);
or UO_767 (O_767,N_7860,N_9386);
nand UO_768 (O_768,N_9871,N_9548);
or UO_769 (O_769,N_9407,N_7712);
and UO_770 (O_770,N_8495,N_9572);
and UO_771 (O_771,N_7624,N_8577);
nand UO_772 (O_772,N_8857,N_8004);
or UO_773 (O_773,N_8754,N_8198);
nor UO_774 (O_774,N_8523,N_7794);
nor UO_775 (O_775,N_7802,N_8835);
or UO_776 (O_776,N_8937,N_9966);
nand UO_777 (O_777,N_9311,N_8366);
nor UO_778 (O_778,N_8111,N_9886);
nor UO_779 (O_779,N_8647,N_8046);
xor UO_780 (O_780,N_8735,N_8994);
nor UO_781 (O_781,N_9169,N_9500);
or UO_782 (O_782,N_8409,N_7557);
nand UO_783 (O_783,N_9914,N_7837);
and UO_784 (O_784,N_9862,N_8949);
nor UO_785 (O_785,N_9979,N_8915);
nor UO_786 (O_786,N_7580,N_8101);
or UO_787 (O_787,N_9521,N_9525);
or UO_788 (O_788,N_7703,N_8381);
nor UO_789 (O_789,N_8058,N_9488);
or UO_790 (O_790,N_9210,N_8139);
or UO_791 (O_791,N_7776,N_8052);
or UO_792 (O_792,N_8100,N_9654);
or UO_793 (O_793,N_9001,N_8170);
nand UO_794 (O_794,N_9121,N_8567);
nand UO_795 (O_795,N_9893,N_7848);
and UO_796 (O_796,N_8229,N_9743);
nor UO_797 (O_797,N_8281,N_9657);
nand UO_798 (O_798,N_9876,N_9823);
and UO_799 (O_799,N_7666,N_8403);
or UO_800 (O_800,N_7631,N_8786);
and UO_801 (O_801,N_9633,N_8972);
or UO_802 (O_802,N_8222,N_8107);
and UO_803 (O_803,N_7552,N_9435);
and UO_804 (O_804,N_8062,N_9825);
and UO_805 (O_805,N_9357,N_9238);
nand UO_806 (O_806,N_8693,N_8993);
nor UO_807 (O_807,N_8767,N_7835);
nor UO_808 (O_808,N_9691,N_9061);
or UO_809 (O_809,N_9082,N_7804);
nor UO_810 (O_810,N_7745,N_7905);
nand UO_811 (O_811,N_9150,N_7923);
or UO_812 (O_812,N_9527,N_9268);
nand UO_813 (O_813,N_8879,N_7506);
xnor UO_814 (O_814,N_8162,N_7531);
and UO_815 (O_815,N_9804,N_9731);
nor UO_816 (O_816,N_8934,N_9753);
nand UO_817 (O_817,N_9908,N_8234);
nor UO_818 (O_818,N_9243,N_8386);
and UO_819 (O_819,N_9446,N_9981);
or UO_820 (O_820,N_8751,N_8060);
nor UO_821 (O_821,N_7577,N_8391);
or UO_822 (O_822,N_9482,N_7795);
nor UO_823 (O_823,N_7947,N_8612);
and UO_824 (O_824,N_9364,N_7647);
nor UO_825 (O_825,N_9354,N_9678);
nor UO_826 (O_826,N_9072,N_9542);
nor UO_827 (O_827,N_7528,N_8465);
nand UO_828 (O_828,N_8761,N_9320);
and UO_829 (O_829,N_7761,N_8853);
and UO_830 (O_830,N_8979,N_8259);
nor UO_831 (O_831,N_9937,N_9648);
and UO_832 (O_832,N_9250,N_9559);
or UO_833 (O_833,N_9313,N_7632);
xor UO_834 (O_834,N_9106,N_8684);
xor UO_835 (O_835,N_9181,N_8370);
nor UO_836 (O_836,N_7782,N_8160);
or UO_837 (O_837,N_7635,N_8055);
or UO_838 (O_838,N_8346,N_8024);
nor UO_839 (O_839,N_9975,N_8946);
xor UO_840 (O_840,N_8656,N_8285);
nand UO_841 (O_841,N_9140,N_8079);
or UO_842 (O_842,N_9163,N_8948);
and UO_843 (O_843,N_8796,N_9115);
nor UO_844 (O_844,N_8249,N_9665);
nor UO_845 (O_845,N_8962,N_8801);
nor UO_846 (O_846,N_9626,N_8445);
nand UO_847 (O_847,N_9727,N_9503);
nor UO_848 (O_848,N_8672,N_8638);
nand UO_849 (O_849,N_8651,N_9765);
nand UO_850 (O_850,N_9171,N_9136);
nor UO_851 (O_851,N_7979,N_8209);
nand UO_852 (O_852,N_9717,N_7726);
and UO_853 (O_853,N_7694,N_8838);
or UO_854 (O_854,N_9204,N_9234);
nor UO_855 (O_855,N_8823,N_9004);
nor UO_856 (O_856,N_8365,N_8525);
or UO_857 (O_857,N_9706,N_8916);
or UO_858 (O_858,N_8610,N_8561);
nor UO_859 (O_859,N_9502,N_7735);
nor UO_860 (O_860,N_8973,N_8276);
nand UO_861 (O_861,N_9349,N_7695);
and UO_862 (O_862,N_7740,N_9032);
and UO_863 (O_863,N_8437,N_8175);
and UO_864 (O_864,N_8133,N_8009);
or UO_865 (O_865,N_9977,N_9767);
and UO_866 (O_866,N_7686,N_9754);
or UO_867 (O_867,N_8169,N_9963);
and UO_868 (O_868,N_9037,N_9595);
or UO_869 (O_869,N_7891,N_8708);
and UO_870 (O_870,N_8113,N_8186);
nand UO_871 (O_871,N_9590,N_8622);
and UO_872 (O_872,N_8149,N_7865);
nor UO_873 (O_873,N_8015,N_7987);
nor UO_874 (O_874,N_8849,N_8163);
and UO_875 (O_875,N_9041,N_9596);
nand UO_876 (O_876,N_9904,N_9039);
nand UO_877 (O_877,N_9453,N_8228);
nor UO_878 (O_878,N_7502,N_9881);
nor UO_879 (O_879,N_9162,N_7643);
nand UO_880 (O_880,N_9069,N_9220);
nor UO_881 (O_881,N_8339,N_8245);
xor UO_882 (O_882,N_8204,N_8443);
or UO_883 (O_883,N_7591,N_9014);
and UO_884 (O_884,N_9985,N_7584);
nor UO_885 (O_885,N_7613,N_9890);
nor UO_886 (O_886,N_7967,N_9529);
nand UO_887 (O_887,N_7917,N_8384);
nor UO_888 (O_888,N_9462,N_9631);
and UO_889 (O_889,N_9177,N_8703);
nand UO_890 (O_890,N_7752,N_8252);
nand UO_891 (O_891,N_8272,N_9844);
nor UO_892 (O_892,N_9560,N_9745);
or UO_893 (O_893,N_9752,N_8640);
and UO_894 (O_894,N_9067,N_7916);
nor UO_895 (O_895,N_8918,N_7997);
and UO_896 (O_896,N_8598,N_9965);
and UO_897 (O_897,N_7984,N_8539);
nor UO_898 (O_898,N_9870,N_7862);
and UO_899 (O_899,N_8700,N_7953);
and UO_900 (O_900,N_7637,N_8927);
and UO_901 (O_901,N_8021,N_8756);
or UO_902 (O_902,N_8347,N_8822);
or UO_903 (O_903,N_7587,N_9118);
nor UO_904 (O_904,N_9746,N_9373);
nand UO_905 (O_905,N_8520,N_9388);
and UO_906 (O_906,N_8502,N_9297);
or UO_907 (O_907,N_7519,N_7532);
or UO_908 (O_908,N_8382,N_8673);
or UO_909 (O_909,N_8375,N_8989);
and UO_910 (O_910,N_8496,N_7697);
nor UO_911 (O_911,N_8543,N_7957);
nand UO_912 (O_912,N_8154,N_7954);
and UO_913 (O_913,N_7930,N_9603);
or UO_914 (O_914,N_7977,N_9906);
nand UO_915 (O_915,N_9519,N_8172);
nand UO_916 (O_916,N_7787,N_9395);
or UO_917 (O_917,N_9969,N_7525);
nor UO_918 (O_918,N_9707,N_9325);
nand UO_919 (O_919,N_7693,N_8251);
and UO_920 (O_920,N_9552,N_9437);
nand UO_921 (O_921,N_8447,N_7863);
or UO_922 (O_922,N_7817,N_9170);
or UO_923 (O_923,N_8846,N_9387);
or UO_924 (O_924,N_9956,N_7642);
nor UO_925 (O_925,N_7646,N_9995);
and UO_926 (O_926,N_8677,N_8882);
or UO_927 (O_927,N_7970,N_8572);
nor UO_928 (O_928,N_9025,N_9044);
nand UO_929 (O_929,N_9910,N_9515);
nor UO_930 (O_930,N_8896,N_9050);
nand UO_931 (O_931,N_9218,N_9543);
and UO_932 (O_932,N_7741,N_9213);
or UO_933 (O_933,N_8642,N_8925);
and UO_934 (O_934,N_7688,N_9305);
nor UO_935 (O_935,N_8905,N_8959);
and UO_936 (O_936,N_8449,N_9413);
nand UO_937 (O_937,N_7919,N_9935);
or UO_938 (O_938,N_9629,N_9512);
and UO_939 (O_939,N_8590,N_9159);
nand UO_940 (O_940,N_9046,N_9255);
nand UO_941 (O_941,N_9679,N_8702);
or UO_942 (O_942,N_9649,N_9701);
nor UO_943 (O_943,N_9469,N_9758);
and UO_944 (O_944,N_9609,N_8758);
or UO_945 (O_945,N_8776,N_8165);
or UO_946 (O_946,N_7747,N_8623);
or UO_947 (O_947,N_7980,N_8839);
nand UO_948 (O_948,N_9005,N_7819);
nand UO_949 (O_949,N_9338,N_8441);
nand UO_950 (O_950,N_9104,N_8578);
and UO_951 (O_951,N_9346,N_9970);
and UO_952 (O_952,N_7998,N_9215);
nand UO_953 (O_953,N_9352,N_8446);
and UO_954 (O_954,N_9151,N_7826);
and UO_955 (O_955,N_7725,N_8069);
nor UO_956 (O_956,N_9214,N_9653);
and UO_957 (O_957,N_8422,N_9086);
nand UO_958 (O_958,N_9340,N_8156);
or UO_959 (O_959,N_7746,N_9555);
nand UO_960 (O_960,N_7903,N_7565);
nor UO_961 (O_961,N_8201,N_7962);
or UO_962 (O_962,N_9449,N_9095);
nor UO_963 (O_963,N_8721,N_7938);
and UO_964 (O_964,N_9289,N_7718);
and UO_965 (O_965,N_7716,N_7926);
nor UO_966 (O_966,N_7760,N_9821);
and UO_967 (O_967,N_8188,N_9855);
nor UO_968 (O_968,N_9225,N_9222);
or UO_969 (O_969,N_9571,N_9241);
and UO_970 (O_970,N_7555,N_9842);
nor UO_971 (O_971,N_8012,N_8206);
nor UO_972 (O_972,N_8303,N_8691);
nand UO_973 (O_973,N_7996,N_9715);
and UO_974 (O_974,N_8298,N_8080);
and UO_975 (O_975,N_8766,N_9508);
nor UO_976 (O_976,N_9168,N_9770);
xor UO_977 (O_977,N_9434,N_7948);
or UO_978 (O_978,N_7540,N_8106);
or UO_979 (O_979,N_8924,N_8576);
and UO_980 (O_980,N_7720,N_9160);
nand UO_981 (O_981,N_8562,N_8132);
and UO_982 (O_982,N_8585,N_7859);
or UO_983 (O_983,N_9420,N_9546);
nor UO_984 (O_984,N_9366,N_7898);
and UO_985 (O_985,N_9534,N_8718);
or UO_986 (O_986,N_9335,N_9339);
nand UO_987 (O_987,N_9951,N_8178);
or UO_988 (O_988,N_9314,N_8688);
or UO_989 (O_989,N_9391,N_7696);
or UO_990 (O_990,N_8515,N_9003);
and UO_991 (O_991,N_7560,N_8646);
or UO_992 (O_992,N_8781,N_9972);
nand UO_993 (O_993,N_8317,N_8423);
or UO_994 (O_994,N_9336,N_8136);
nand UO_995 (O_995,N_8247,N_8524);
nor UO_996 (O_996,N_8497,N_8504);
nand UO_997 (O_997,N_8547,N_9950);
and UO_998 (O_998,N_8791,N_9637);
nand UO_999 (O_999,N_9299,N_9351);
nor UO_1000 (O_1000,N_8629,N_7771);
nor UO_1001 (O_1001,N_9724,N_7691);
and UO_1002 (O_1002,N_7774,N_9187);
nor UO_1003 (O_1003,N_9917,N_8589);
nor UO_1004 (O_1004,N_8550,N_9698);
nand UO_1005 (O_1005,N_9612,N_9868);
nor UO_1006 (O_1006,N_9742,N_9393);
nand UO_1007 (O_1007,N_9907,N_9769);
nand UO_1008 (O_1008,N_8575,N_9916);
nor UO_1009 (O_1009,N_7663,N_9634);
nor UO_1010 (O_1010,N_9158,N_8871);
and UO_1011 (O_1011,N_8987,N_7612);
nor UO_1012 (O_1012,N_9507,N_8941);
nand UO_1013 (O_1013,N_9786,N_9860);
xor UO_1014 (O_1014,N_9718,N_9608);
and UO_1015 (O_1015,N_8606,N_9117);
nor UO_1016 (O_1016,N_8870,N_8319);
and UO_1017 (O_1017,N_9009,N_7951);
xnor UO_1018 (O_1018,N_7942,N_8255);
or UO_1019 (O_1019,N_9522,N_8088);
and UO_1020 (O_1020,N_7943,N_9480);
nor UO_1021 (O_1021,N_7773,N_8652);
nor UO_1022 (O_1022,N_8603,N_7574);
nor UO_1023 (O_1023,N_7927,N_7910);
nor UO_1024 (O_1024,N_9757,N_8568);
nand UO_1025 (O_1025,N_8095,N_8982);
nand UO_1026 (O_1026,N_9490,N_7657);
nor UO_1027 (O_1027,N_8187,N_9362);
nor UO_1028 (O_1028,N_9574,N_9406);
nand UO_1029 (O_1029,N_8842,N_9091);
and UO_1030 (O_1030,N_8493,N_7946);
and UO_1031 (O_1031,N_9989,N_8184);
xnor UO_1032 (O_1032,N_7630,N_7516);
nand UO_1033 (O_1033,N_9138,N_9152);
and UO_1034 (O_1034,N_9402,N_7564);
nor UO_1035 (O_1035,N_9492,N_9573);
and UO_1036 (O_1036,N_8000,N_8869);
or UO_1037 (O_1037,N_9440,N_9410);
and UO_1038 (O_1038,N_7936,N_9682);
or UO_1039 (O_1039,N_7768,N_8831);
nand UO_1040 (O_1040,N_7619,N_9122);
and UO_1041 (O_1041,N_7645,N_9282);
nand UO_1042 (O_1042,N_9826,N_8168);
and UO_1043 (O_1043,N_7708,N_8815);
nor UO_1044 (O_1044,N_8593,N_8710);
nand UO_1045 (O_1045,N_8807,N_8337);
nand UO_1046 (O_1046,N_8802,N_7731);
nor UO_1047 (O_1047,N_9945,N_7704);
and UO_1048 (O_1048,N_9423,N_8246);
xnor UO_1049 (O_1049,N_8283,N_9454);
nand UO_1050 (O_1050,N_8057,N_8195);
nand UO_1051 (O_1051,N_7833,N_8771);
nor UO_1052 (O_1052,N_9784,N_9610);
nand UO_1053 (O_1053,N_9903,N_9668);
xnor UO_1054 (O_1054,N_7702,N_9356);
nand UO_1055 (O_1055,N_9301,N_8120);
and UO_1056 (O_1056,N_8811,N_9801);
nor UO_1057 (O_1057,N_9899,N_7698);
or UO_1058 (O_1058,N_9240,N_8314);
or UO_1059 (O_1059,N_8604,N_8036);
and UO_1060 (O_1060,N_8115,N_9300);
nand UO_1061 (O_1061,N_7911,N_8930);
or UO_1062 (O_1062,N_7734,N_7617);
nand UO_1063 (O_1063,N_7983,N_8083);
or UO_1064 (O_1064,N_9246,N_7515);
or UO_1065 (O_1065,N_7822,N_8906);
nand UO_1066 (O_1066,N_7785,N_7544);
nor UO_1067 (O_1067,N_8359,N_8476);
nor UO_1068 (O_1068,N_9076,N_8902);
nand UO_1069 (O_1069,N_9670,N_7793);
nand UO_1070 (O_1070,N_7791,N_8344);
nor UO_1071 (O_1071,N_7513,N_7674);
nor UO_1072 (O_1072,N_8552,N_8914);
or UO_1073 (O_1073,N_8096,N_8752);
nand UO_1074 (O_1074,N_8388,N_7616);
nand UO_1075 (O_1075,N_8865,N_9551);
and UO_1076 (O_1076,N_8098,N_8332);
nand UO_1077 (O_1077,N_8521,N_8018);
or UO_1078 (O_1078,N_9891,N_8960);
and UO_1079 (O_1079,N_8775,N_9909);
nand UO_1080 (O_1080,N_7545,N_7592);
nand UO_1081 (O_1081,N_9497,N_8595);
nor UO_1082 (O_1082,N_9620,N_9465);
nand UO_1083 (O_1083,N_8076,N_8828);
and UO_1084 (O_1084,N_7881,N_7594);
nor UO_1085 (O_1085,N_9708,N_9685);
or UO_1086 (O_1086,N_9996,N_7883);
nor UO_1087 (O_1087,N_9326,N_9087);
and UO_1088 (O_1088,N_9531,N_8264);
nand UO_1089 (O_1089,N_8928,N_8957);
or UO_1090 (O_1090,N_9493,N_8028);
or UO_1091 (O_1091,N_7576,N_8248);
and UO_1092 (O_1092,N_8884,N_8105);
nor UO_1093 (O_1093,N_9602,N_7852);
nor UO_1094 (O_1094,N_8619,N_8190);
and UO_1095 (O_1095,N_8306,N_7841);
nor UO_1096 (O_1096,N_7805,N_8614);
and UO_1097 (O_1097,N_9273,N_9684);
and UO_1098 (O_1098,N_7526,N_9132);
or UO_1099 (O_1099,N_9926,N_9175);
and UO_1100 (O_1100,N_7914,N_8159);
or UO_1101 (O_1101,N_8425,N_9604);
nand UO_1102 (O_1102,N_7581,N_8749);
or UO_1103 (O_1103,N_7816,N_7512);
and UO_1104 (O_1104,N_9579,N_8996);
nand UO_1105 (O_1105,N_8484,N_7729);
nand UO_1106 (O_1106,N_8227,N_8545);
nand UO_1107 (O_1107,N_8430,N_9867);
nor UO_1108 (O_1108,N_7796,N_9575);
nor UO_1109 (O_1109,N_8320,N_9998);
or UO_1110 (O_1110,N_7600,N_7550);
and UO_1111 (O_1111,N_7656,N_9553);
or UO_1112 (O_1112,N_8683,N_9247);
nor UO_1113 (O_1113,N_9712,N_8889);
and UO_1114 (O_1114,N_8278,N_7879);
and UO_1115 (O_1115,N_7907,N_7541);
or UO_1116 (O_1116,N_9873,N_9809);
nor UO_1117 (O_1117,N_8361,N_9430);
nand UO_1118 (O_1118,N_9127,N_8026);
and UO_1119 (O_1119,N_8983,N_8858);
or UO_1120 (O_1120,N_8582,N_9986);
nand UO_1121 (O_1121,N_8436,N_7877);
or UO_1122 (O_1122,N_7569,N_8908);
nor UO_1123 (O_1123,N_9442,N_9952);
nor UO_1124 (O_1124,N_7609,N_7885);
and UO_1125 (O_1125,N_8868,N_9549);
or UO_1126 (O_1126,N_7654,N_7827);
nand UO_1127 (O_1127,N_7968,N_9312);
or UO_1128 (O_1128,N_9591,N_8345);
and UO_1129 (O_1129,N_8270,N_9732);
nor UO_1130 (O_1130,N_8630,N_9055);
xnor UO_1131 (O_1131,N_8714,N_9057);
or UO_1132 (O_1132,N_9226,N_7558);
nand UO_1133 (O_1133,N_9584,N_8140);
nor UO_1134 (O_1134,N_9756,N_8275);
nor UO_1135 (O_1135,N_9792,N_7618);
nand UO_1136 (O_1136,N_9412,N_7683);
nor UO_1137 (O_1137,N_9857,N_8931);
or UO_1138 (O_1138,N_9723,N_9664);
or UO_1139 (O_1139,N_9561,N_8085);
or UO_1140 (O_1140,N_8943,N_8006);
nand UO_1141 (O_1141,N_9258,N_9641);
and UO_1142 (O_1142,N_8886,N_9361);
or UO_1143 (O_1143,N_9355,N_9530);
and UO_1144 (O_1144,N_8792,N_9667);
or UO_1145 (O_1145,N_7736,N_7625);
nor UO_1146 (O_1146,N_7994,N_8180);
nor UO_1147 (O_1147,N_8471,N_8301);
and UO_1148 (O_1148,N_7918,N_8793);
nand UO_1149 (O_1149,N_7738,N_7653);
nor UO_1150 (O_1150,N_8119,N_9693);
nand UO_1151 (O_1151,N_8431,N_9381);
or UO_1152 (O_1152,N_7982,N_8118);
and UO_1153 (O_1153,N_8729,N_8072);
and UO_1154 (O_1154,N_9540,N_9113);
or UO_1155 (O_1155,N_9417,N_8077);
or UO_1156 (O_1156,N_9785,N_8217);
nand UO_1157 (O_1157,N_9029,N_9265);
and UO_1158 (O_1158,N_8596,N_9024);
and UO_1159 (O_1159,N_9184,N_8371);
nand UO_1160 (O_1160,N_8399,N_8146);
nor UO_1161 (O_1161,N_9541,N_8649);
nor UO_1162 (O_1162,N_8851,N_7641);
and UO_1163 (O_1163,N_9562,N_9794);
and UO_1164 (O_1164,N_9291,N_8042);
and UO_1165 (O_1165,N_9018,N_7832);
nand UO_1166 (O_1166,N_8833,N_7602);
nor UO_1167 (O_1167,N_9567,N_8897);
nand UO_1168 (O_1168,N_8559,N_8499);
and UO_1169 (O_1169,N_9697,N_8824);
nor UO_1170 (O_1170,N_9580,N_9990);
nor UO_1171 (O_1171,N_9872,N_9456);
nand UO_1172 (O_1172,N_9007,N_8151);
and UO_1173 (O_1173,N_8174,N_8966);
nor UO_1174 (O_1174,N_9850,N_7875);
nand UO_1175 (O_1175,N_8216,N_9814);
nor UO_1176 (O_1176,N_8728,N_7682);
and UO_1177 (O_1177,N_8617,N_8110);
and UO_1178 (O_1178,N_9049,N_9303);
nand UO_1179 (O_1179,N_8071,N_7779);
or UO_1180 (O_1180,N_9224,N_8389);
or UO_1181 (O_1181,N_9262,N_9128);
or UO_1182 (O_1182,N_8513,N_9978);
nor UO_1183 (O_1183,N_7548,N_8719);
nor UO_1184 (O_1184,N_9093,N_8017);
and UO_1185 (O_1185,N_8890,N_8557);
or UO_1186 (O_1186,N_9601,N_8047);
or UO_1187 (O_1187,N_7899,N_9083);
nor UO_1188 (O_1188,N_7701,N_7960);
and UO_1189 (O_1189,N_8123,N_9484);
and UO_1190 (O_1190,N_7842,N_8333);
nand UO_1191 (O_1191,N_9489,N_8192);
and UO_1192 (O_1192,N_9737,N_7566);
or UO_1193 (O_1193,N_9577,N_8859);
or UO_1194 (O_1194,N_8685,N_9942);
nor UO_1195 (O_1195,N_9824,N_7853);
or UO_1196 (O_1196,N_7669,N_8795);
and UO_1197 (O_1197,N_8820,N_9759);
and UO_1198 (O_1198,N_9031,N_8964);
or UO_1199 (O_1199,N_8368,N_9424);
nor UO_1200 (O_1200,N_9638,N_8401);
and UO_1201 (O_1201,N_7920,N_9237);
nand UO_1202 (O_1202,N_9673,N_9370);
nor UO_1203 (O_1203,N_9369,N_8804);
or UO_1204 (O_1204,N_9056,N_8158);
nand UO_1205 (O_1205,N_8289,N_9129);
and UO_1206 (O_1206,N_7543,N_8059);
and UO_1207 (O_1207,N_8035,N_7717);
and UO_1208 (O_1208,N_9556,N_9741);
and UO_1209 (O_1209,N_9686,N_8901);
and UO_1210 (O_1210,N_7721,N_8961);
or UO_1211 (O_1211,N_7588,N_9895);
nand UO_1212 (O_1212,N_9889,N_7724);
nand UO_1213 (O_1213,N_8854,N_8324);
nor UO_1214 (O_1214,N_9495,N_8990);
and UO_1215 (O_1215,N_9997,N_8478);
or UO_1216 (O_1216,N_8840,N_8097);
and UO_1217 (O_1217,N_9636,N_8510);
or UO_1218 (O_1218,N_7549,N_8958);
nand UO_1219 (O_1219,N_9513,N_8894);
nand UO_1220 (O_1220,N_9874,N_8230);
or UO_1221 (O_1221,N_9988,N_9382);
and UO_1222 (O_1222,N_8220,N_9761);
or UO_1223 (O_1223,N_9882,N_8634);
or UO_1224 (O_1224,N_8291,N_8556);
nor UO_1225 (O_1225,N_8467,N_9194);
nand UO_1226 (O_1226,N_7958,N_8474);
nor UO_1227 (O_1227,N_9376,N_8611);
nor UO_1228 (O_1228,N_7730,N_7966);
or UO_1229 (O_1229,N_8138,N_8895);
xor UO_1230 (O_1230,N_9557,N_9587);
or UO_1231 (O_1231,N_8837,N_8378);
and UO_1232 (O_1232,N_8023,N_9422);
nand UO_1233 (O_1233,N_7775,N_9172);
nand UO_1234 (O_1234,N_8463,N_8377);
nor UO_1235 (O_1235,N_9307,N_8883);
and UO_1236 (O_1236,N_9251,N_8845);
or UO_1237 (O_1237,N_8847,N_8511);
or UO_1238 (O_1238,N_9411,N_9973);
and UO_1239 (O_1239,N_9520,N_8451);
nor UO_1240 (O_1240,N_8641,N_8005);
and UO_1241 (O_1241,N_8434,N_7661);
or UO_1242 (O_1242,N_8910,N_7971);
nand UO_1243 (O_1243,N_7813,N_8458);
nor UO_1244 (O_1244,N_9473,N_9206);
or UO_1245 (O_1245,N_9847,N_9960);
or UO_1246 (O_1246,N_9569,N_9865);
nand UO_1247 (O_1247,N_8808,N_7873);
nor UO_1248 (O_1248,N_9205,N_8770);
and UO_1249 (O_1249,N_8665,N_9191);
and UO_1250 (O_1250,N_9877,N_8672);
or UO_1251 (O_1251,N_9915,N_9870);
or UO_1252 (O_1252,N_9440,N_7757);
or UO_1253 (O_1253,N_9643,N_9785);
xnor UO_1254 (O_1254,N_9064,N_7858);
and UO_1255 (O_1255,N_8725,N_9895);
or UO_1256 (O_1256,N_8341,N_9660);
and UO_1257 (O_1257,N_8640,N_8212);
and UO_1258 (O_1258,N_7898,N_7990);
and UO_1259 (O_1259,N_9582,N_9272);
and UO_1260 (O_1260,N_8542,N_8722);
or UO_1261 (O_1261,N_7571,N_8590);
and UO_1262 (O_1262,N_7640,N_7877);
nor UO_1263 (O_1263,N_8700,N_7874);
and UO_1264 (O_1264,N_8370,N_9177);
nand UO_1265 (O_1265,N_8575,N_8001);
or UO_1266 (O_1266,N_7505,N_8438);
nor UO_1267 (O_1267,N_9752,N_8811);
nor UO_1268 (O_1268,N_9576,N_8063);
or UO_1269 (O_1269,N_9591,N_8058);
nand UO_1270 (O_1270,N_9581,N_8196);
or UO_1271 (O_1271,N_7678,N_9035);
nor UO_1272 (O_1272,N_8382,N_8876);
and UO_1273 (O_1273,N_9984,N_9201);
or UO_1274 (O_1274,N_8654,N_9360);
or UO_1275 (O_1275,N_9956,N_7593);
and UO_1276 (O_1276,N_9305,N_8861);
nand UO_1277 (O_1277,N_9402,N_8448);
or UO_1278 (O_1278,N_9702,N_9365);
or UO_1279 (O_1279,N_8303,N_9247);
nand UO_1280 (O_1280,N_7912,N_9019);
nand UO_1281 (O_1281,N_8700,N_9978);
or UO_1282 (O_1282,N_8232,N_7966);
nor UO_1283 (O_1283,N_9432,N_8274);
or UO_1284 (O_1284,N_8548,N_7683);
nor UO_1285 (O_1285,N_9625,N_8826);
nor UO_1286 (O_1286,N_9329,N_7764);
or UO_1287 (O_1287,N_8176,N_9794);
nand UO_1288 (O_1288,N_8466,N_8298);
or UO_1289 (O_1289,N_8122,N_7889);
nand UO_1290 (O_1290,N_8847,N_9419);
and UO_1291 (O_1291,N_7984,N_7658);
and UO_1292 (O_1292,N_8255,N_9957);
and UO_1293 (O_1293,N_9345,N_9634);
nand UO_1294 (O_1294,N_8499,N_8971);
or UO_1295 (O_1295,N_9088,N_8249);
nand UO_1296 (O_1296,N_8299,N_8504);
or UO_1297 (O_1297,N_8865,N_9330);
nand UO_1298 (O_1298,N_9116,N_9213);
or UO_1299 (O_1299,N_8928,N_9889);
nand UO_1300 (O_1300,N_8025,N_9657);
nand UO_1301 (O_1301,N_9503,N_7795);
and UO_1302 (O_1302,N_8727,N_8005);
nand UO_1303 (O_1303,N_9544,N_8995);
and UO_1304 (O_1304,N_8347,N_8299);
and UO_1305 (O_1305,N_8918,N_8520);
and UO_1306 (O_1306,N_7792,N_8962);
or UO_1307 (O_1307,N_9253,N_9077);
nor UO_1308 (O_1308,N_8698,N_7901);
nor UO_1309 (O_1309,N_8924,N_9599);
or UO_1310 (O_1310,N_9903,N_9534);
or UO_1311 (O_1311,N_9139,N_7770);
nor UO_1312 (O_1312,N_7679,N_8921);
nand UO_1313 (O_1313,N_9286,N_9081);
nand UO_1314 (O_1314,N_8293,N_8937);
and UO_1315 (O_1315,N_8519,N_9639);
nor UO_1316 (O_1316,N_9644,N_9189);
and UO_1317 (O_1317,N_9200,N_8971);
nand UO_1318 (O_1318,N_9699,N_7756);
nor UO_1319 (O_1319,N_9209,N_8763);
nor UO_1320 (O_1320,N_9021,N_8598);
nor UO_1321 (O_1321,N_8294,N_8322);
nor UO_1322 (O_1322,N_7579,N_8830);
or UO_1323 (O_1323,N_8881,N_9454);
nor UO_1324 (O_1324,N_8531,N_8639);
and UO_1325 (O_1325,N_9970,N_8899);
or UO_1326 (O_1326,N_8021,N_8097);
nor UO_1327 (O_1327,N_9171,N_8195);
nor UO_1328 (O_1328,N_9109,N_9156);
nand UO_1329 (O_1329,N_8008,N_8670);
nand UO_1330 (O_1330,N_8748,N_9704);
and UO_1331 (O_1331,N_8778,N_8078);
nor UO_1332 (O_1332,N_7955,N_8950);
or UO_1333 (O_1333,N_9181,N_9714);
nor UO_1334 (O_1334,N_9331,N_9884);
and UO_1335 (O_1335,N_9809,N_7920);
or UO_1336 (O_1336,N_9419,N_9753);
and UO_1337 (O_1337,N_7706,N_8412);
and UO_1338 (O_1338,N_8441,N_9087);
and UO_1339 (O_1339,N_9125,N_8275);
nand UO_1340 (O_1340,N_7504,N_9498);
or UO_1341 (O_1341,N_9264,N_9394);
or UO_1342 (O_1342,N_8430,N_8393);
and UO_1343 (O_1343,N_8640,N_7900);
nand UO_1344 (O_1344,N_8645,N_8899);
nor UO_1345 (O_1345,N_9626,N_9349);
or UO_1346 (O_1346,N_7981,N_8656);
or UO_1347 (O_1347,N_8535,N_8823);
nor UO_1348 (O_1348,N_8238,N_8205);
nand UO_1349 (O_1349,N_8781,N_8653);
nor UO_1350 (O_1350,N_8231,N_9320);
nand UO_1351 (O_1351,N_8074,N_8041);
nor UO_1352 (O_1352,N_8050,N_8596);
and UO_1353 (O_1353,N_9262,N_9108);
nor UO_1354 (O_1354,N_9010,N_7749);
nor UO_1355 (O_1355,N_8359,N_8186);
nand UO_1356 (O_1356,N_8870,N_7876);
nand UO_1357 (O_1357,N_9840,N_7707);
and UO_1358 (O_1358,N_7500,N_8103);
and UO_1359 (O_1359,N_8342,N_8472);
nand UO_1360 (O_1360,N_9911,N_7704);
and UO_1361 (O_1361,N_9135,N_8837);
and UO_1362 (O_1362,N_8133,N_7983);
and UO_1363 (O_1363,N_8550,N_9006);
nand UO_1364 (O_1364,N_8275,N_8000);
nor UO_1365 (O_1365,N_8851,N_8775);
and UO_1366 (O_1366,N_8821,N_9452);
and UO_1367 (O_1367,N_7901,N_8184);
and UO_1368 (O_1368,N_8424,N_9600);
nor UO_1369 (O_1369,N_9660,N_7881);
and UO_1370 (O_1370,N_9757,N_8939);
or UO_1371 (O_1371,N_9317,N_7873);
or UO_1372 (O_1372,N_9750,N_8645);
nand UO_1373 (O_1373,N_8763,N_8408);
and UO_1374 (O_1374,N_9627,N_9711);
nand UO_1375 (O_1375,N_8477,N_8104);
nor UO_1376 (O_1376,N_7977,N_7853);
nor UO_1377 (O_1377,N_7519,N_9096);
and UO_1378 (O_1378,N_9217,N_9034);
nor UO_1379 (O_1379,N_9209,N_8471);
nor UO_1380 (O_1380,N_8117,N_8439);
and UO_1381 (O_1381,N_9086,N_8319);
nor UO_1382 (O_1382,N_9063,N_8628);
and UO_1383 (O_1383,N_8365,N_8222);
nand UO_1384 (O_1384,N_8128,N_8607);
nand UO_1385 (O_1385,N_9030,N_9938);
and UO_1386 (O_1386,N_8015,N_9517);
or UO_1387 (O_1387,N_9141,N_7807);
and UO_1388 (O_1388,N_9005,N_8698);
nand UO_1389 (O_1389,N_7733,N_9036);
or UO_1390 (O_1390,N_7810,N_9848);
and UO_1391 (O_1391,N_7545,N_7588);
and UO_1392 (O_1392,N_8979,N_8958);
nor UO_1393 (O_1393,N_8115,N_8791);
and UO_1394 (O_1394,N_9545,N_7554);
and UO_1395 (O_1395,N_8285,N_9278);
nand UO_1396 (O_1396,N_7867,N_8059);
nor UO_1397 (O_1397,N_8686,N_8159);
or UO_1398 (O_1398,N_9798,N_9253);
or UO_1399 (O_1399,N_7764,N_8253);
or UO_1400 (O_1400,N_9309,N_9575);
nand UO_1401 (O_1401,N_9157,N_8238);
and UO_1402 (O_1402,N_9044,N_8626);
or UO_1403 (O_1403,N_9142,N_9765);
or UO_1404 (O_1404,N_8191,N_9489);
nand UO_1405 (O_1405,N_9658,N_7729);
or UO_1406 (O_1406,N_9431,N_9877);
nor UO_1407 (O_1407,N_9644,N_7576);
nand UO_1408 (O_1408,N_8883,N_8019);
and UO_1409 (O_1409,N_8253,N_9483);
nor UO_1410 (O_1410,N_9225,N_8332);
or UO_1411 (O_1411,N_9837,N_7688);
and UO_1412 (O_1412,N_7835,N_8819);
and UO_1413 (O_1413,N_8878,N_8752);
and UO_1414 (O_1414,N_8036,N_7593);
nor UO_1415 (O_1415,N_7985,N_9476);
nor UO_1416 (O_1416,N_9282,N_9689);
nor UO_1417 (O_1417,N_8180,N_9359);
or UO_1418 (O_1418,N_8466,N_8119);
xor UO_1419 (O_1419,N_8772,N_7646);
nand UO_1420 (O_1420,N_8321,N_7541);
and UO_1421 (O_1421,N_7969,N_9486);
or UO_1422 (O_1422,N_8224,N_9006);
or UO_1423 (O_1423,N_8597,N_9300);
nand UO_1424 (O_1424,N_8840,N_9448);
nor UO_1425 (O_1425,N_9424,N_8114);
nand UO_1426 (O_1426,N_9086,N_7840);
or UO_1427 (O_1427,N_9650,N_8916);
or UO_1428 (O_1428,N_8814,N_7776);
nor UO_1429 (O_1429,N_7930,N_7602);
or UO_1430 (O_1430,N_8797,N_9753);
or UO_1431 (O_1431,N_7988,N_8187);
nand UO_1432 (O_1432,N_8171,N_9463);
nand UO_1433 (O_1433,N_8739,N_8559);
and UO_1434 (O_1434,N_8782,N_7857);
or UO_1435 (O_1435,N_9684,N_7741);
and UO_1436 (O_1436,N_8285,N_8524);
or UO_1437 (O_1437,N_7697,N_8801);
nand UO_1438 (O_1438,N_7539,N_8467);
or UO_1439 (O_1439,N_8976,N_7821);
nand UO_1440 (O_1440,N_9214,N_9450);
nand UO_1441 (O_1441,N_9795,N_9486);
or UO_1442 (O_1442,N_9373,N_8361);
or UO_1443 (O_1443,N_9982,N_8694);
or UO_1444 (O_1444,N_7621,N_9806);
and UO_1445 (O_1445,N_8185,N_8336);
and UO_1446 (O_1446,N_9514,N_8670);
nand UO_1447 (O_1447,N_9222,N_9503);
and UO_1448 (O_1448,N_9286,N_7876);
nor UO_1449 (O_1449,N_9708,N_9795);
nand UO_1450 (O_1450,N_8078,N_9138);
nand UO_1451 (O_1451,N_7654,N_7561);
nor UO_1452 (O_1452,N_9767,N_9982);
and UO_1453 (O_1453,N_8513,N_9006);
or UO_1454 (O_1454,N_7978,N_8564);
nand UO_1455 (O_1455,N_9839,N_9111);
nor UO_1456 (O_1456,N_9576,N_8470);
nand UO_1457 (O_1457,N_7782,N_7852);
nand UO_1458 (O_1458,N_9159,N_8656);
nor UO_1459 (O_1459,N_9895,N_9103);
xnor UO_1460 (O_1460,N_7510,N_8639);
or UO_1461 (O_1461,N_9035,N_9803);
and UO_1462 (O_1462,N_7785,N_9074);
nor UO_1463 (O_1463,N_8677,N_8162);
or UO_1464 (O_1464,N_8281,N_7504);
or UO_1465 (O_1465,N_8163,N_9746);
nand UO_1466 (O_1466,N_9620,N_9779);
xor UO_1467 (O_1467,N_8098,N_8695);
or UO_1468 (O_1468,N_9388,N_7573);
nor UO_1469 (O_1469,N_8855,N_9113);
nor UO_1470 (O_1470,N_7669,N_8797);
nor UO_1471 (O_1471,N_9716,N_9491);
nor UO_1472 (O_1472,N_8920,N_8628);
and UO_1473 (O_1473,N_8293,N_9875);
nand UO_1474 (O_1474,N_8717,N_7947);
and UO_1475 (O_1475,N_8324,N_8405);
or UO_1476 (O_1476,N_8801,N_9746);
or UO_1477 (O_1477,N_7629,N_8472);
and UO_1478 (O_1478,N_8715,N_8246);
nor UO_1479 (O_1479,N_8977,N_7989);
xnor UO_1480 (O_1480,N_8390,N_9323);
nand UO_1481 (O_1481,N_9743,N_8194);
nor UO_1482 (O_1482,N_9188,N_9389);
nor UO_1483 (O_1483,N_8703,N_9719);
nor UO_1484 (O_1484,N_9459,N_9542);
and UO_1485 (O_1485,N_7919,N_9861);
or UO_1486 (O_1486,N_8038,N_9547);
and UO_1487 (O_1487,N_8072,N_8922);
or UO_1488 (O_1488,N_9684,N_8375);
and UO_1489 (O_1489,N_9194,N_9846);
nor UO_1490 (O_1490,N_9413,N_9459);
and UO_1491 (O_1491,N_9620,N_9517);
nor UO_1492 (O_1492,N_9034,N_9566);
and UO_1493 (O_1493,N_7648,N_8942);
nand UO_1494 (O_1494,N_8638,N_9358);
or UO_1495 (O_1495,N_8447,N_7943);
and UO_1496 (O_1496,N_8789,N_9807);
nor UO_1497 (O_1497,N_8701,N_9186);
nor UO_1498 (O_1498,N_9806,N_7569);
and UO_1499 (O_1499,N_7907,N_8126);
endmodule