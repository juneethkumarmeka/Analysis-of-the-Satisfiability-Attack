module basic_750_5000_1000_5_levels_1xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
nand U0 (N_0,In_17,In_427);
nand U1 (N_1,In_263,In_456);
and U2 (N_2,In_37,In_526);
or U3 (N_3,In_314,In_642);
nor U4 (N_4,In_599,In_433);
nand U5 (N_5,In_31,In_527);
or U6 (N_6,In_168,In_161);
and U7 (N_7,In_229,In_667);
or U8 (N_8,In_59,In_419);
or U9 (N_9,In_193,In_323);
nand U10 (N_10,In_414,In_256);
nor U11 (N_11,In_26,In_436);
and U12 (N_12,In_151,In_80);
or U13 (N_13,In_465,In_457);
nor U14 (N_14,In_637,In_257);
nand U15 (N_15,In_89,In_500);
or U16 (N_16,In_75,In_696);
nand U17 (N_17,In_681,In_297);
nand U18 (N_18,In_676,In_544);
or U19 (N_19,In_201,In_141);
or U20 (N_20,In_452,In_622);
and U21 (N_21,In_541,In_115);
or U22 (N_22,In_210,In_568);
or U23 (N_23,In_8,In_589);
nand U24 (N_24,In_390,In_357);
and U25 (N_25,In_312,In_84);
and U26 (N_26,In_392,In_209);
nand U27 (N_27,In_643,In_410);
and U28 (N_28,In_25,In_540);
or U29 (N_29,In_422,In_554);
and U30 (N_30,In_721,In_716);
and U31 (N_31,In_566,In_406);
or U32 (N_32,In_601,In_7);
and U33 (N_33,In_579,In_387);
and U34 (N_34,In_735,In_389);
and U35 (N_35,In_81,In_114);
nor U36 (N_36,In_635,In_685);
or U37 (N_37,In_202,In_298);
nor U38 (N_38,In_130,In_92);
nor U39 (N_39,In_638,In_158);
nor U40 (N_40,In_16,In_134);
and U41 (N_41,In_471,In_548);
and U42 (N_42,In_483,In_222);
or U43 (N_43,In_86,In_307);
and U44 (N_44,In_35,In_46);
nand U45 (N_45,In_473,In_309);
nand U46 (N_46,In_9,In_138);
and U47 (N_47,In_77,In_564);
or U48 (N_48,In_632,In_523);
nand U49 (N_49,In_664,In_588);
or U50 (N_50,In_137,In_73);
and U51 (N_51,In_559,In_425);
nand U52 (N_52,In_370,In_475);
or U53 (N_53,In_286,In_394);
or U54 (N_54,In_21,In_22);
nand U55 (N_55,In_591,In_205);
nor U56 (N_56,In_143,In_226);
nand U57 (N_57,In_724,In_520);
or U58 (N_58,In_10,In_654);
and U59 (N_59,In_748,In_482);
or U60 (N_60,In_631,In_79);
xnor U61 (N_61,In_179,In_431);
nand U62 (N_62,In_275,In_194);
nand U63 (N_63,In_491,In_615);
and U64 (N_64,In_479,In_100);
nor U65 (N_65,In_53,In_647);
nor U66 (N_66,In_562,In_693);
nor U67 (N_67,In_238,In_76);
and U68 (N_68,In_156,In_247);
and U69 (N_69,In_274,In_492);
or U70 (N_70,In_393,In_413);
or U71 (N_71,In_509,In_188);
xor U72 (N_72,In_459,In_669);
nand U73 (N_73,In_4,In_60);
and U74 (N_74,In_187,In_411);
or U75 (N_75,In_573,In_352);
or U76 (N_76,In_565,In_214);
nor U77 (N_77,In_489,In_512);
nor U78 (N_78,In_455,In_381);
nor U79 (N_79,In_602,In_233);
and U80 (N_80,In_186,In_169);
nor U81 (N_81,In_407,In_474);
nor U82 (N_82,In_361,In_590);
nor U83 (N_83,In_458,In_490);
or U84 (N_84,In_619,In_386);
or U85 (N_85,In_0,In_269);
or U86 (N_86,In_88,In_362);
nand U87 (N_87,In_120,In_227);
and U88 (N_88,In_358,In_742);
and U89 (N_89,In_196,In_206);
and U90 (N_90,In_747,In_694);
or U91 (N_91,In_118,In_749);
nor U92 (N_92,In_710,In_731);
nand U93 (N_93,In_692,In_396);
nor U94 (N_94,In_466,In_348);
nand U95 (N_95,In_14,In_145);
or U96 (N_96,In_709,In_620);
or U97 (N_97,In_221,In_97);
nand U98 (N_98,In_133,In_20);
nor U99 (N_99,In_658,In_687);
or U100 (N_100,In_231,In_426);
or U101 (N_101,In_714,In_525);
nand U102 (N_102,In_435,In_614);
and U103 (N_103,In_551,In_29);
and U104 (N_104,In_45,In_657);
nand U105 (N_105,In_271,In_488);
and U106 (N_106,In_350,In_572);
nand U107 (N_107,In_325,In_737);
and U108 (N_108,In_424,In_310);
or U109 (N_109,In_360,In_575);
nand U110 (N_110,In_518,In_514);
or U111 (N_111,In_688,In_90);
nor U112 (N_112,In_675,In_237);
nand U113 (N_113,In_660,In_701);
and U114 (N_114,In_713,In_534);
or U115 (N_115,In_241,In_68);
and U116 (N_116,In_404,In_445);
or U117 (N_117,In_101,In_403);
nand U118 (N_118,In_356,In_74);
and U119 (N_119,In_2,In_172);
or U120 (N_120,In_108,In_157);
nor U121 (N_121,In_184,In_159);
and U122 (N_122,In_105,In_618);
nand U123 (N_123,In_400,In_71);
nor U124 (N_124,In_296,In_107);
nor U125 (N_125,In_537,In_715);
or U126 (N_126,In_487,In_434);
nand U127 (N_127,In_417,In_727);
and U128 (N_128,In_596,In_245);
nand U129 (N_129,In_529,In_663);
or U130 (N_130,In_597,In_163);
nor U131 (N_131,In_712,In_177);
or U132 (N_132,In_204,In_498);
and U133 (N_133,In_335,In_379);
nor U134 (N_134,In_524,In_87);
nand U135 (N_135,In_371,In_587);
nor U136 (N_136,In_15,In_480);
or U137 (N_137,In_70,In_305);
nand U138 (N_138,In_251,In_195);
and U139 (N_139,In_98,In_135);
nor U140 (N_140,In_653,In_399);
or U141 (N_141,In_355,In_285);
nand U142 (N_142,In_144,In_418);
nand U143 (N_143,In_125,In_39);
or U144 (N_144,In_671,In_744);
nor U145 (N_145,In_267,In_720);
and U146 (N_146,In_167,In_699);
or U147 (N_147,In_337,In_504);
nand U148 (N_148,In_725,In_136);
nor U149 (N_149,In_13,In_723);
or U150 (N_150,In_333,In_569);
nor U151 (N_151,In_367,In_265);
or U152 (N_152,In_388,In_391);
nand U153 (N_153,In_600,In_303);
nor U154 (N_154,In_516,In_547);
or U155 (N_155,In_545,In_472);
nand U156 (N_156,In_364,In_464);
nand U157 (N_157,In_142,In_260);
and U158 (N_158,In_33,In_690);
nand U159 (N_159,In_299,In_270);
nand U160 (N_160,In_578,In_401);
nor U161 (N_161,In_423,In_734);
and U162 (N_162,In_191,In_543);
or U163 (N_163,In_584,In_372);
or U164 (N_164,In_429,In_652);
and U165 (N_165,In_639,In_273);
nand U166 (N_166,In_28,In_365);
or U167 (N_167,In_738,In_636);
nor U168 (N_168,In_448,In_219);
nor U169 (N_169,In_383,In_533);
and U170 (N_170,In_585,In_746);
nand U171 (N_171,In_557,In_248);
nor U172 (N_172,In_58,In_450);
nand U173 (N_173,In_164,In_683);
nand U174 (N_174,In_449,In_532);
or U175 (N_175,In_155,In_656);
or U176 (N_176,In_609,In_48);
nor U177 (N_177,In_517,In_351);
nand U178 (N_178,In_617,In_535);
or U179 (N_179,In_34,In_294);
and U180 (N_180,In_650,In_625);
or U181 (N_181,In_284,In_166);
and U182 (N_182,In_531,In_339);
and U183 (N_183,In_612,In_123);
nor U184 (N_184,In_463,In_36);
nor U185 (N_185,In_278,In_382);
and U186 (N_186,In_322,In_616);
nand U187 (N_187,In_342,In_662);
or U188 (N_188,In_495,In_152);
nor U189 (N_189,In_373,In_729);
nor U190 (N_190,In_672,In_374);
nor U191 (N_191,In_262,In_363);
nand U192 (N_192,In_192,In_510);
nand U193 (N_193,In_644,In_739);
nor U194 (N_194,In_230,In_319);
nor U195 (N_195,In_728,In_69);
or U196 (N_196,In_508,In_740);
or U197 (N_197,In_344,In_65);
nand U198 (N_198,In_85,In_213);
and U199 (N_199,In_375,In_180);
nor U200 (N_200,In_608,In_212);
and U201 (N_201,In_324,In_522);
and U202 (N_202,In_606,In_234);
nor U203 (N_203,In_235,In_293);
nor U204 (N_204,In_126,In_730);
nor U205 (N_205,In_290,In_592);
or U206 (N_206,In_327,In_397);
and U207 (N_207,In_67,In_261);
or U208 (N_208,In_200,In_6);
nand U209 (N_209,In_674,In_3);
and U210 (N_210,In_502,In_287);
and U211 (N_211,In_160,In_57);
nor U212 (N_212,In_542,In_405);
and U213 (N_213,In_41,In_154);
or U214 (N_214,In_536,In_677);
and U215 (N_215,In_467,In_72);
or U216 (N_216,In_82,In_481);
or U217 (N_217,In_50,In_56);
or U218 (N_218,In_453,In_673);
or U219 (N_219,In_302,In_240);
nor U220 (N_220,In_439,In_150);
nor U221 (N_221,In_678,In_430);
and U222 (N_222,In_232,In_292);
nand U223 (N_223,In_94,In_485);
and U224 (N_224,In_556,In_258);
nor U225 (N_225,In_703,In_96);
or U226 (N_226,In_580,In_477);
nand U227 (N_227,In_165,In_623);
nand U228 (N_228,In_461,In_27);
nor U229 (N_229,In_610,In_613);
nand U230 (N_230,In_661,In_301);
nor U231 (N_231,In_611,In_148);
nor U232 (N_232,In_11,In_468);
and U233 (N_233,In_328,In_507);
nor U234 (N_234,In_268,In_220);
and U235 (N_235,In_546,In_528);
nor U236 (N_236,In_62,In_571);
and U237 (N_237,In_420,In_176);
nor U238 (N_238,In_668,In_207);
nand U239 (N_239,In_377,In_380);
and U240 (N_240,In_32,In_630);
nor U241 (N_241,In_103,In_460);
nand U242 (N_242,In_421,In_651);
or U243 (N_243,In_266,In_259);
nor U244 (N_244,In_501,In_104);
and U245 (N_245,In_570,In_503);
nor U246 (N_246,In_49,In_395);
or U247 (N_247,In_338,In_586);
nor U248 (N_248,In_745,In_462);
and U249 (N_249,In_649,In_93);
nand U250 (N_250,In_311,In_243);
and U251 (N_251,In_254,In_552);
nor U252 (N_252,In_595,In_1);
nand U253 (N_253,In_279,In_320);
nor U254 (N_254,In_282,In_670);
nand U255 (N_255,In_558,In_486);
nand U256 (N_256,In_304,In_128);
or U257 (N_257,In_110,In_249);
and U258 (N_258,In_117,In_624);
and U259 (N_259,In_680,In_646);
or U260 (N_260,In_308,In_366);
nand U261 (N_261,In_55,In_47);
nand U262 (N_262,In_12,In_181);
nor U263 (N_263,In_291,In_695);
nand U264 (N_264,In_122,In_581);
or U265 (N_265,In_216,In_629);
and U266 (N_266,In_689,In_354);
or U267 (N_267,In_655,In_197);
nor U268 (N_268,In_499,In_506);
nor U269 (N_269,In_702,In_444);
or U270 (N_270,In_19,In_341);
nand U271 (N_271,In_470,In_185);
nor U272 (N_272,In_437,In_119);
and U273 (N_273,In_326,In_706);
or U274 (N_274,In_717,In_641);
and U275 (N_275,In_684,In_153);
or U276 (N_276,In_626,In_682);
nor U277 (N_277,In_376,In_255);
nor U278 (N_278,In_183,In_347);
or U279 (N_279,In_561,In_228);
or U280 (N_280,In_147,In_52);
nor U281 (N_281,In_66,In_329);
nor U282 (N_282,In_666,In_321);
and U283 (N_283,In_170,In_345);
or U284 (N_284,In_408,In_44);
nand U285 (N_285,In_440,In_127);
and U286 (N_286,In_574,In_223);
or U287 (N_287,In_99,In_182);
nand U288 (N_288,In_369,In_306);
nor U289 (N_289,In_211,In_61);
and U290 (N_290,In_515,In_604);
nor U291 (N_291,In_733,In_648);
and U292 (N_292,In_332,In_704);
or U293 (N_293,In_679,In_711);
nand U294 (N_294,In_139,In_334);
nand U295 (N_295,In_38,In_553);
and U296 (N_296,In_484,In_109);
and U297 (N_297,In_208,In_594);
and U298 (N_298,In_129,In_598);
or U299 (N_299,In_697,In_83);
nand U300 (N_300,In_313,In_521);
and U301 (N_301,In_628,In_113);
or U302 (N_302,In_719,In_331);
nor U303 (N_303,In_698,In_224);
nand U304 (N_304,In_78,In_640);
or U305 (N_305,In_446,In_63);
or U306 (N_306,In_174,In_132);
nand U307 (N_307,In_634,In_252);
nor U308 (N_308,In_560,In_576);
and U309 (N_309,In_691,In_645);
nand U310 (N_310,In_563,In_218);
or U311 (N_311,In_276,In_494);
or U312 (N_312,In_5,In_368);
nor U313 (N_313,In_316,In_621);
nand U314 (N_314,In_442,In_162);
or U315 (N_315,In_451,In_513);
or U316 (N_316,In_505,In_140);
and U317 (N_317,In_441,In_605);
and U318 (N_318,In_190,In_199);
nand U319 (N_319,In_330,In_443);
nor U320 (N_320,In_732,In_384);
or U321 (N_321,In_705,In_246);
nor U322 (N_322,In_607,In_627);
and U323 (N_323,In_402,In_280);
nor U324 (N_324,In_593,In_359);
nand U325 (N_325,In_64,In_24);
and U326 (N_326,In_454,In_478);
nor U327 (N_327,In_633,In_116);
or U328 (N_328,In_131,In_577);
nand U329 (N_329,In_409,In_198);
nor U330 (N_330,In_283,In_416);
and U331 (N_331,In_530,In_91);
or U332 (N_332,In_18,In_438);
nor U333 (N_333,In_272,In_95);
nand U334 (N_334,In_743,In_686);
nor U335 (N_335,In_295,In_736);
nor U336 (N_336,In_415,In_493);
nor U337 (N_337,In_146,In_555);
nor U338 (N_338,In_121,In_318);
xor U339 (N_339,In_343,In_659);
nand U340 (N_340,In_412,In_708);
nand U341 (N_341,In_242,In_378);
and U342 (N_342,In_349,In_54);
and U343 (N_343,In_432,In_567);
or U344 (N_344,In_289,In_42);
nor U345 (N_345,In_549,In_469);
and U346 (N_346,In_30,In_519);
nand U347 (N_347,In_51,In_281);
nor U348 (N_348,In_511,In_102);
and U349 (N_349,In_497,In_539);
nor U350 (N_350,In_250,In_23);
xor U351 (N_351,In_428,In_665);
and U352 (N_352,In_124,In_244);
nor U353 (N_353,In_496,In_217);
or U354 (N_354,In_277,In_726);
or U355 (N_355,In_353,In_582);
nor U356 (N_356,In_336,In_106);
and U357 (N_357,In_112,In_236);
or U358 (N_358,In_718,In_340);
nor U359 (N_359,In_315,In_40);
or U360 (N_360,In_550,In_189);
nor U361 (N_361,In_225,In_398);
xor U362 (N_362,In_171,In_603);
or U363 (N_363,In_707,In_346);
nand U364 (N_364,In_722,In_215);
nor U365 (N_365,In_700,In_538);
nor U366 (N_366,In_741,In_264);
or U367 (N_367,In_385,In_447);
and U368 (N_368,In_173,In_583);
nor U369 (N_369,In_317,In_175);
nor U370 (N_370,In_239,In_253);
nor U371 (N_371,In_178,In_111);
or U372 (N_372,In_288,In_149);
or U373 (N_373,In_476,In_43);
nand U374 (N_374,In_203,In_300);
nand U375 (N_375,In_368,In_21);
and U376 (N_376,In_494,In_77);
and U377 (N_377,In_119,In_280);
nand U378 (N_378,In_718,In_265);
nand U379 (N_379,In_712,In_57);
nand U380 (N_380,In_696,In_361);
or U381 (N_381,In_430,In_698);
and U382 (N_382,In_215,In_531);
nand U383 (N_383,In_746,In_731);
or U384 (N_384,In_548,In_553);
or U385 (N_385,In_563,In_548);
or U386 (N_386,In_700,In_335);
nand U387 (N_387,In_593,In_297);
nor U388 (N_388,In_251,In_445);
or U389 (N_389,In_14,In_214);
and U390 (N_390,In_481,In_394);
or U391 (N_391,In_622,In_476);
or U392 (N_392,In_360,In_162);
nand U393 (N_393,In_155,In_242);
or U394 (N_394,In_647,In_455);
and U395 (N_395,In_744,In_15);
nand U396 (N_396,In_247,In_71);
or U397 (N_397,In_91,In_316);
nor U398 (N_398,In_685,In_481);
nor U399 (N_399,In_619,In_336);
or U400 (N_400,In_465,In_45);
and U401 (N_401,In_96,In_1);
nand U402 (N_402,In_641,In_83);
nor U403 (N_403,In_378,In_592);
or U404 (N_404,In_163,In_36);
nor U405 (N_405,In_312,In_112);
nand U406 (N_406,In_130,In_598);
nand U407 (N_407,In_749,In_440);
and U408 (N_408,In_137,In_556);
nor U409 (N_409,In_652,In_79);
and U410 (N_410,In_211,In_567);
or U411 (N_411,In_540,In_631);
nor U412 (N_412,In_419,In_123);
nand U413 (N_413,In_363,In_568);
nor U414 (N_414,In_181,In_721);
nand U415 (N_415,In_295,In_407);
nand U416 (N_416,In_436,In_499);
nand U417 (N_417,In_43,In_22);
and U418 (N_418,In_199,In_83);
nand U419 (N_419,In_367,In_488);
or U420 (N_420,In_402,In_723);
nor U421 (N_421,In_40,In_645);
nand U422 (N_422,In_255,In_397);
nand U423 (N_423,In_416,In_475);
nand U424 (N_424,In_257,In_258);
or U425 (N_425,In_235,In_541);
nor U426 (N_426,In_249,In_739);
nand U427 (N_427,In_219,In_156);
or U428 (N_428,In_148,In_476);
or U429 (N_429,In_146,In_480);
and U430 (N_430,In_116,In_75);
nand U431 (N_431,In_267,In_304);
nor U432 (N_432,In_390,In_419);
or U433 (N_433,In_102,In_649);
and U434 (N_434,In_548,In_273);
and U435 (N_435,In_729,In_40);
and U436 (N_436,In_514,In_361);
nand U437 (N_437,In_249,In_63);
nor U438 (N_438,In_163,In_52);
nor U439 (N_439,In_443,In_374);
nand U440 (N_440,In_326,In_554);
nand U441 (N_441,In_744,In_151);
and U442 (N_442,In_377,In_628);
nand U443 (N_443,In_104,In_195);
nand U444 (N_444,In_465,In_588);
and U445 (N_445,In_368,In_9);
or U446 (N_446,In_151,In_568);
and U447 (N_447,In_40,In_507);
and U448 (N_448,In_14,In_77);
nor U449 (N_449,In_334,In_669);
and U450 (N_450,In_99,In_711);
nand U451 (N_451,In_617,In_72);
xnor U452 (N_452,In_410,In_375);
nor U453 (N_453,In_324,In_422);
or U454 (N_454,In_45,In_402);
nand U455 (N_455,In_641,In_499);
nand U456 (N_456,In_220,In_673);
and U457 (N_457,In_669,In_194);
nor U458 (N_458,In_552,In_749);
nand U459 (N_459,In_9,In_142);
or U460 (N_460,In_91,In_635);
nor U461 (N_461,In_489,In_741);
nor U462 (N_462,In_193,In_413);
or U463 (N_463,In_144,In_12);
nor U464 (N_464,In_402,In_485);
nand U465 (N_465,In_376,In_618);
nand U466 (N_466,In_48,In_490);
and U467 (N_467,In_121,In_65);
or U468 (N_468,In_277,In_438);
and U469 (N_469,In_393,In_419);
nor U470 (N_470,In_237,In_264);
nor U471 (N_471,In_8,In_551);
or U472 (N_472,In_644,In_114);
or U473 (N_473,In_33,In_73);
nand U474 (N_474,In_216,In_318);
and U475 (N_475,In_352,In_145);
or U476 (N_476,In_613,In_728);
and U477 (N_477,In_620,In_302);
nand U478 (N_478,In_475,In_71);
or U479 (N_479,In_343,In_167);
nand U480 (N_480,In_453,In_90);
and U481 (N_481,In_205,In_686);
nor U482 (N_482,In_450,In_688);
nand U483 (N_483,In_517,In_344);
and U484 (N_484,In_443,In_457);
nor U485 (N_485,In_109,In_287);
and U486 (N_486,In_56,In_684);
nor U487 (N_487,In_377,In_655);
nor U488 (N_488,In_136,In_294);
nand U489 (N_489,In_56,In_610);
nor U490 (N_490,In_107,In_267);
and U491 (N_491,In_166,In_97);
or U492 (N_492,In_640,In_610);
nor U493 (N_493,In_27,In_175);
or U494 (N_494,In_355,In_146);
and U495 (N_495,In_141,In_549);
nand U496 (N_496,In_324,In_363);
nand U497 (N_497,In_76,In_326);
or U498 (N_498,In_334,In_35);
or U499 (N_499,In_428,In_340);
and U500 (N_500,In_581,In_328);
nor U501 (N_501,In_479,In_334);
and U502 (N_502,In_437,In_152);
nor U503 (N_503,In_482,In_21);
nand U504 (N_504,In_582,In_367);
nand U505 (N_505,In_324,In_610);
or U506 (N_506,In_439,In_310);
nand U507 (N_507,In_36,In_371);
or U508 (N_508,In_38,In_483);
nor U509 (N_509,In_52,In_674);
nand U510 (N_510,In_46,In_277);
nor U511 (N_511,In_685,In_277);
and U512 (N_512,In_612,In_285);
or U513 (N_513,In_278,In_182);
or U514 (N_514,In_78,In_356);
xor U515 (N_515,In_314,In_687);
and U516 (N_516,In_218,In_429);
nor U517 (N_517,In_504,In_165);
or U518 (N_518,In_225,In_343);
and U519 (N_519,In_254,In_616);
nand U520 (N_520,In_524,In_730);
nand U521 (N_521,In_615,In_185);
nor U522 (N_522,In_385,In_428);
and U523 (N_523,In_79,In_430);
nor U524 (N_524,In_14,In_604);
nor U525 (N_525,In_666,In_207);
and U526 (N_526,In_611,In_442);
nand U527 (N_527,In_467,In_458);
and U528 (N_528,In_641,In_438);
nand U529 (N_529,In_175,In_735);
nor U530 (N_530,In_142,In_427);
nand U531 (N_531,In_453,In_677);
nor U532 (N_532,In_630,In_177);
and U533 (N_533,In_277,In_108);
nor U534 (N_534,In_113,In_157);
nand U535 (N_535,In_245,In_463);
or U536 (N_536,In_381,In_742);
or U537 (N_537,In_158,In_284);
nor U538 (N_538,In_287,In_203);
nor U539 (N_539,In_688,In_37);
nand U540 (N_540,In_381,In_94);
xor U541 (N_541,In_342,In_655);
and U542 (N_542,In_425,In_161);
nor U543 (N_543,In_395,In_69);
nand U544 (N_544,In_276,In_638);
and U545 (N_545,In_437,In_608);
and U546 (N_546,In_391,In_549);
nor U547 (N_547,In_108,In_348);
and U548 (N_548,In_211,In_206);
nor U549 (N_549,In_565,In_32);
nand U550 (N_550,In_261,In_175);
or U551 (N_551,In_615,In_664);
or U552 (N_552,In_79,In_76);
nand U553 (N_553,In_370,In_101);
or U554 (N_554,In_624,In_122);
or U555 (N_555,In_627,In_243);
and U556 (N_556,In_476,In_683);
or U557 (N_557,In_624,In_70);
nand U558 (N_558,In_119,In_211);
xor U559 (N_559,In_433,In_267);
nor U560 (N_560,In_160,In_672);
and U561 (N_561,In_57,In_327);
or U562 (N_562,In_163,In_524);
or U563 (N_563,In_240,In_158);
or U564 (N_564,In_16,In_316);
nand U565 (N_565,In_121,In_727);
and U566 (N_566,In_117,In_560);
and U567 (N_567,In_659,In_169);
nor U568 (N_568,In_576,In_325);
and U569 (N_569,In_488,In_647);
nor U570 (N_570,In_740,In_379);
nand U571 (N_571,In_722,In_313);
nor U572 (N_572,In_275,In_334);
and U573 (N_573,In_31,In_406);
and U574 (N_574,In_217,In_328);
nand U575 (N_575,In_568,In_159);
nand U576 (N_576,In_235,In_440);
and U577 (N_577,In_587,In_589);
or U578 (N_578,In_419,In_608);
nor U579 (N_579,In_322,In_381);
or U580 (N_580,In_531,In_245);
or U581 (N_581,In_81,In_123);
or U582 (N_582,In_412,In_125);
nand U583 (N_583,In_687,In_33);
and U584 (N_584,In_88,In_396);
or U585 (N_585,In_477,In_748);
nand U586 (N_586,In_733,In_673);
nor U587 (N_587,In_272,In_35);
nor U588 (N_588,In_544,In_92);
nand U589 (N_589,In_69,In_630);
and U590 (N_590,In_352,In_715);
nand U591 (N_591,In_643,In_508);
nor U592 (N_592,In_126,In_311);
and U593 (N_593,In_228,In_216);
nand U594 (N_594,In_715,In_534);
or U595 (N_595,In_326,In_492);
or U596 (N_596,In_107,In_420);
nor U597 (N_597,In_647,In_295);
or U598 (N_598,In_317,In_567);
nand U599 (N_599,In_379,In_615);
and U600 (N_600,In_562,In_238);
or U601 (N_601,In_728,In_142);
and U602 (N_602,In_368,In_429);
and U603 (N_603,In_82,In_500);
nor U604 (N_604,In_568,In_73);
nand U605 (N_605,In_425,In_89);
nand U606 (N_606,In_208,In_450);
and U607 (N_607,In_258,In_296);
nand U608 (N_608,In_572,In_585);
nand U609 (N_609,In_507,In_593);
nand U610 (N_610,In_106,In_597);
nand U611 (N_611,In_572,In_429);
or U612 (N_612,In_546,In_179);
nor U613 (N_613,In_108,In_48);
nor U614 (N_614,In_168,In_4);
or U615 (N_615,In_430,In_105);
nand U616 (N_616,In_607,In_581);
nand U617 (N_617,In_83,In_426);
or U618 (N_618,In_121,In_555);
nor U619 (N_619,In_701,In_228);
or U620 (N_620,In_546,In_531);
nor U621 (N_621,In_450,In_29);
nor U622 (N_622,In_286,In_115);
nand U623 (N_623,In_381,In_68);
nand U624 (N_624,In_554,In_233);
or U625 (N_625,In_504,In_580);
nor U626 (N_626,In_232,In_580);
or U627 (N_627,In_321,In_137);
nor U628 (N_628,In_745,In_90);
nor U629 (N_629,In_592,In_296);
and U630 (N_630,In_410,In_368);
nand U631 (N_631,In_348,In_2);
and U632 (N_632,In_621,In_114);
and U633 (N_633,In_440,In_745);
or U634 (N_634,In_325,In_504);
nand U635 (N_635,In_238,In_721);
and U636 (N_636,In_45,In_422);
and U637 (N_637,In_450,In_428);
or U638 (N_638,In_0,In_158);
xnor U639 (N_639,In_340,In_329);
nor U640 (N_640,In_169,In_521);
nand U641 (N_641,In_334,In_146);
and U642 (N_642,In_475,In_547);
or U643 (N_643,In_162,In_405);
or U644 (N_644,In_271,In_517);
or U645 (N_645,In_245,In_9);
nor U646 (N_646,In_220,In_477);
and U647 (N_647,In_328,In_228);
nand U648 (N_648,In_629,In_219);
and U649 (N_649,In_707,In_643);
nand U650 (N_650,In_497,In_260);
or U651 (N_651,In_236,In_666);
or U652 (N_652,In_652,In_629);
nand U653 (N_653,In_469,In_653);
nand U654 (N_654,In_705,In_432);
and U655 (N_655,In_491,In_302);
nor U656 (N_656,In_117,In_551);
and U657 (N_657,In_439,In_122);
nor U658 (N_658,In_139,In_191);
and U659 (N_659,In_554,In_136);
and U660 (N_660,In_609,In_679);
nor U661 (N_661,In_524,In_294);
nand U662 (N_662,In_642,In_585);
nand U663 (N_663,In_250,In_110);
nor U664 (N_664,In_145,In_500);
nand U665 (N_665,In_475,In_254);
nand U666 (N_666,In_33,In_301);
or U667 (N_667,In_710,In_71);
nand U668 (N_668,In_330,In_269);
nor U669 (N_669,In_575,In_223);
nor U670 (N_670,In_300,In_322);
and U671 (N_671,In_338,In_306);
nor U672 (N_672,In_117,In_537);
nor U673 (N_673,In_565,In_25);
nor U674 (N_674,In_433,In_437);
nand U675 (N_675,In_697,In_262);
and U676 (N_676,In_136,In_699);
or U677 (N_677,In_98,In_195);
nand U678 (N_678,In_224,In_494);
and U679 (N_679,In_624,In_665);
or U680 (N_680,In_97,In_553);
or U681 (N_681,In_469,In_574);
nor U682 (N_682,In_257,In_691);
and U683 (N_683,In_147,In_577);
nor U684 (N_684,In_219,In_30);
or U685 (N_685,In_249,In_175);
and U686 (N_686,In_309,In_722);
nand U687 (N_687,In_270,In_43);
nor U688 (N_688,In_128,In_463);
and U689 (N_689,In_709,In_655);
nand U690 (N_690,In_327,In_346);
nor U691 (N_691,In_78,In_589);
nand U692 (N_692,In_89,In_460);
and U693 (N_693,In_496,In_232);
nor U694 (N_694,In_566,In_439);
nand U695 (N_695,In_471,In_279);
and U696 (N_696,In_741,In_637);
nor U697 (N_697,In_172,In_514);
or U698 (N_698,In_473,In_99);
nor U699 (N_699,In_332,In_333);
nor U700 (N_700,In_370,In_124);
nand U701 (N_701,In_738,In_243);
and U702 (N_702,In_242,In_708);
and U703 (N_703,In_336,In_198);
and U704 (N_704,In_143,In_139);
or U705 (N_705,In_260,In_636);
nor U706 (N_706,In_728,In_653);
nand U707 (N_707,In_220,In_669);
or U708 (N_708,In_219,In_134);
nand U709 (N_709,In_545,In_368);
nor U710 (N_710,In_27,In_606);
and U711 (N_711,In_731,In_503);
nor U712 (N_712,In_376,In_705);
and U713 (N_713,In_196,In_546);
or U714 (N_714,In_408,In_645);
or U715 (N_715,In_154,In_647);
nor U716 (N_716,In_637,In_152);
nor U717 (N_717,In_131,In_276);
or U718 (N_718,In_420,In_240);
nand U719 (N_719,In_513,In_393);
or U720 (N_720,In_291,In_358);
nor U721 (N_721,In_12,In_471);
and U722 (N_722,In_211,In_130);
nor U723 (N_723,In_18,In_658);
or U724 (N_724,In_131,In_208);
or U725 (N_725,In_688,In_717);
nand U726 (N_726,In_65,In_538);
or U727 (N_727,In_667,In_716);
nand U728 (N_728,In_517,In_127);
nor U729 (N_729,In_395,In_649);
or U730 (N_730,In_337,In_379);
nand U731 (N_731,In_403,In_604);
or U732 (N_732,In_250,In_531);
nor U733 (N_733,In_106,In_406);
nand U734 (N_734,In_370,In_318);
nor U735 (N_735,In_365,In_202);
and U736 (N_736,In_120,In_154);
and U737 (N_737,In_181,In_457);
or U738 (N_738,In_205,In_444);
nor U739 (N_739,In_167,In_68);
nand U740 (N_740,In_460,In_82);
nor U741 (N_741,In_80,In_209);
and U742 (N_742,In_338,In_335);
or U743 (N_743,In_136,In_705);
nor U744 (N_744,In_275,In_85);
nor U745 (N_745,In_694,In_66);
nand U746 (N_746,In_460,In_254);
and U747 (N_747,In_32,In_179);
and U748 (N_748,In_303,In_373);
nor U749 (N_749,In_486,In_580);
nor U750 (N_750,In_286,In_428);
nand U751 (N_751,In_735,In_244);
or U752 (N_752,In_558,In_257);
nor U753 (N_753,In_486,In_121);
nor U754 (N_754,In_83,In_646);
and U755 (N_755,In_133,In_218);
and U756 (N_756,In_267,In_747);
nor U757 (N_757,In_31,In_113);
or U758 (N_758,In_736,In_204);
or U759 (N_759,In_382,In_241);
nand U760 (N_760,In_609,In_373);
nand U761 (N_761,In_733,In_191);
or U762 (N_762,In_319,In_476);
and U763 (N_763,In_350,In_565);
nand U764 (N_764,In_423,In_636);
and U765 (N_765,In_702,In_413);
nor U766 (N_766,In_607,In_519);
nand U767 (N_767,In_737,In_617);
nor U768 (N_768,In_507,In_525);
and U769 (N_769,In_519,In_501);
or U770 (N_770,In_72,In_403);
or U771 (N_771,In_551,In_364);
nand U772 (N_772,In_379,In_511);
and U773 (N_773,In_523,In_238);
nor U774 (N_774,In_146,In_220);
and U775 (N_775,In_362,In_386);
nand U776 (N_776,In_271,In_317);
nor U777 (N_777,In_265,In_100);
and U778 (N_778,In_537,In_365);
or U779 (N_779,In_530,In_640);
nor U780 (N_780,In_708,In_321);
nor U781 (N_781,In_281,In_302);
or U782 (N_782,In_402,In_174);
and U783 (N_783,In_5,In_256);
nor U784 (N_784,In_259,In_65);
nor U785 (N_785,In_211,In_441);
and U786 (N_786,In_643,In_706);
and U787 (N_787,In_565,In_700);
nor U788 (N_788,In_223,In_540);
and U789 (N_789,In_619,In_708);
nor U790 (N_790,In_365,In_564);
or U791 (N_791,In_648,In_148);
nand U792 (N_792,In_312,In_477);
nor U793 (N_793,In_397,In_662);
nand U794 (N_794,In_636,In_476);
or U795 (N_795,In_97,In_691);
xnor U796 (N_796,In_298,In_409);
or U797 (N_797,In_353,In_67);
nor U798 (N_798,In_127,In_360);
or U799 (N_799,In_616,In_455);
or U800 (N_800,In_328,In_494);
and U801 (N_801,In_671,In_246);
nor U802 (N_802,In_695,In_275);
nor U803 (N_803,In_120,In_109);
and U804 (N_804,In_293,In_186);
nor U805 (N_805,In_230,In_713);
nor U806 (N_806,In_738,In_202);
or U807 (N_807,In_679,In_137);
nand U808 (N_808,In_68,In_379);
or U809 (N_809,In_745,In_461);
nor U810 (N_810,In_229,In_588);
and U811 (N_811,In_349,In_571);
nor U812 (N_812,In_661,In_329);
nand U813 (N_813,In_450,In_235);
or U814 (N_814,In_164,In_327);
and U815 (N_815,In_384,In_339);
nand U816 (N_816,In_605,In_266);
or U817 (N_817,In_514,In_4);
or U818 (N_818,In_360,In_482);
nand U819 (N_819,In_405,In_4);
or U820 (N_820,In_387,In_184);
and U821 (N_821,In_438,In_487);
and U822 (N_822,In_267,In_480);
and U823 (N_823,In_704,In_1);
and U824 (N_824,In_558,In_515);
nand U825 (N_825,In_123,In_250);
and U826 (N_826,In_540,In_77);
or U827 (N_827,In_122,In_565);
and U828 (N_828,In_710,In_213);
nand U829 (N_829,In_556,In_282);
nand U830 (N_830,In_86,In_586);
or U831 (N_831,In_402,In_671);
nor U832 (N_832,In_673,In_83);
nor U833 (N_833,In_64,In_262);
and U834 (N_834,In_447,In_648);
or U835 (N_835,In_431,In_559);
or U836 (N_836,In_449,In_465);
or U837 (N_837,In_346,In_680);
nor U838 (N_838,In_115,In_163);
nand U839 (N_839,In_556,In_534);
nor U840 (N_840,In_739,In_654);
nor U841 (N_841,In_178,In_279);
nor U842 (N_842,In_706,In_685);
nor U843 (N_843,In_236,In_517);
nand U844 (N_844,In_109,In_468);
nor U845 (N_845,In_726,In_392);
xnor U846 (N_846,In_114,In_405);
or U847 (N_847,In_453,In_234);
and U848 (N_848,In_148,In_170);
nor U849 (N_849,In_382,In_343);
and U850 (N_850,In_117,In_642);
and U851 (N_851,In_82,In_465);
or U852 (N_852,In_101,In_671);
nor U853 (N_853,In_740,In_283);
nor U854 (N_854,In_119,In_25);
nand U855 (N_855,In_349,In_306);
and U856 (N_856,In_108,In_746);
nand U857 (N_857,In_198,In_730);
nand U858 (N_858,In_92,In_490);
or U859 (N_859,In_42,In_306);
nand U860 (N_860,In_57,In_456);
or U861 (N_861,In_361,In_637);
and U862 (N_862,In_93,In_256);
nor U863 (N_863,In_340,In_43);
and U864 (N_864,In_351,In_202);
and U865 (N_865,In_543,In_295);
or U866 (N_866,In_706,In_92);
nand U867 (N_867,In_510,In_725);
and U868 (N_868,In_682,In_366);
nor U869 (N_869,In_110,In_140);
or U870 (N_870,In_259,In_189);
nor U871 (N_871,In_213,In_596);
or U872 (N_872,In_604,In_312);
or U873 (N_873,In_350,In_684);
nand U874 (N_874,In_622,In_250);
nand U875 (N_875,In_193,In_337);
and U876 (N_876,In_713,In_245);
and U877 (N_877,In_691,In_542);
or U878 (N_878,In_710,In_204);
nor U879 (N_879,In_493,In_462);
and U880 (N_880,In_158,In_281);
nor U881 (N_881,In_158,In_138);
and U882 (N_882,In_529,In_711);
or U883 (N_883,In_130,In_4);
and U884 (N_884,In_77,In_671);
nor U885 (N_885,In_170,In_168);
and U886 (N_886,In_280,In_612);
nand U887 (N_887,In_272,In_317);
nor U888 (N_888,In_607,In_640);
nor U889 (N_889,In_282,In_165);
and U890 (N_890,In_80,In_713);
nand U891 (N_891,In_98,In_106);
and U892 (N_892,In_286,In_259);
or U893 (N_893,In_456,In_726);
nor U894 (N_894,In_473,In_111);
and U895 (N_895,In_144,In_638);
nand U896 (N_896,In_724,In_186);
nand U897 (N_897,In_671,In_112);
nand U898 (N_898,In_662,In_131);
and U899 (N_899,In_439,In_428);
nor U900 (N_900,In_732,In_50);
nand U901 (N_901,In_302,In_7);
nor U902 (N_902,In_520,In_465);
nand U903 (N_903,In_40,In_607);
nand U904 (N_904,In_98,In_228);
nor U905 (N_905,In_109,In_461);
or U906 (N_906,In_494,In_145);
nand U907 (N_907,In_300,In_433);
or U908 (N_908,In_665,In_60);
and U909 (N_909,In_282,In_275);
nand U910 (N_910,In_420,In_648);
nor U911 (N_911,In_329,In_519);
or U912 (N_912,In_0,In_441);
and U913 (N_913,In_235,In_99);
and U914 (N_914,In_666,In_359);
or U915 (N_915,In_73,In_131);
and U916 (N_916,In_688,In_21);
nand U917 (N_917,In_126,In_587);
and U918 (N_918,In_707,In_629);
nand U919 (N_919,In_712,In_107);
nand U920 (N_920,In_499,In_510);
nor U921 (N_921,In_299,In_169);
and U922 (N_922,In_283,In_273);
or U923 (N_923,In_174,In_87);
or U924 (N_924,In_711,In_557);
xnor U925 (N_925,In_553,In_496);
and U926 (N_926,In_138,In_7);
nor U927 (N_927,In_655,In_615);
or U928 (N_928,In_439,In_532);
or U929 (N_929,In_581,In_731);
and U930 (N_930,In_177,In_573);
nor U931 (N_931,In_645,In_51);
xnor U932 (N_932,In_737,In_420);
nor U933 (N_933,In_722,In_97);
nand U934 (N_934,In_229,In_422);
nand U935 (N_935,In_663,In_243);
and U936 (N_936,In_131,In_674);
and U937 (N_937,In_354,In_103);
or U938 (N_938,In_18,In_173);
nand U939 (N_939,In_108,In_375);
or U940 (N_940,In_69,In_137);
nand U941 (N_941,In_719,In_22);
nor U942 (N_942,In_120,In_414);
or U943 (N_943,In_749,In_54);
or U944 (N_944,In_607,In_388);
and U945 (N_945,In_680,In_543);
and U946 (N_946,In_527,In_180);
nor U947 (N_947,In_491,In_123);
nor U948 (N_948,In_654,In_511);
nand U949 (N_949,In_335,In_261);
nor U950 (N_950,In_521,In_103);
nand U951 (N_951,In_363,In_265);
nand U952 (N_952,In_195,In_240);
or U953 (N_953,In_10,In_98);
and U954 (N_954,In_73,In_486);
or U955 (N_955,In_685,In_398);
nor U956 (N_956,In_671,In_296);
and U957 (N_957,In_186,In_17);
nand U958 (N_958,In_184,In_582);
or U959 (N_959,In_565,In_574);
and U960 (N_960,In_619,In_147);
nor U961 (N_961,In_217,In_488);
nor U962 (N_962,In_591,In_117);
nor U963 (N_963,In_456,In_337);
or U964 (N_964,In_461,In_555);
nor U965 (N_965,In_680,In_90);
or U966 (N_966,In_457,In_319);
and U967 (N_967,In_669,In_639);
or U968 (N_968,In_86,In_127);
nor U969 (N_969,In_517,In_294);
xnor U970 (N_970,In_109,In_148);
or U971 (N_971,In_595,In_171);
nor U972 (N_972,In_247,In_468);
nor U973 (N_973,In_229,In_656);
nand U974 (N_974,In_596,In_471);
or U975 (N_975,In_570,In_132);
nor U976 (N_976,In_53,In_477);
or U977 (N_977,In_543,In_132);
or U978 (N_978,In_742,In_62);
nor U979 (N_979,In_206,In_725);
and U980 (N_980,In_472,In_643);
nor U981 (N_981,In_210,In_585);
or U982 (N_982,In_129,In_545);
or U983 (N_983,In_460,In_582);
nand U984 (N_984,In_367,In_354);
and U985 (N_985,In_425,In_743);
and U986 (N_986,In_570,In_49);
nor U987 (N_987,In_676,In_333);
nor U988 (N_988,In_671,In_113);
and U989 (N_989,In_740,In_180);
and U990 (N_990,In_128,In_707);
or U991 (N_991,In_480,In_107);
and U992 (N_992,In_96,In_515);
nor U993 (N_993,In_302,In_293);
nand U994 (N_994,In_206,In_116);
and U995 (N_995,In_136,In_211);
nand U996 (N_996,In_461,In_590);
or U997 (N_997,In_187,In_585);
nor U998 (N_998,In_210,In_492);
or U999 (N_999,In_290,In_599);
or U1000 (N_1000,N_707,N_767);
and U1001 (N_1001,N_241,N_439);
and U1002 (N_1002,N_649,N_729);
nand U1003 (N_1003,N_347,N_365);
or U1004 (N_1004,N_1,N_383);
nor U1005 (N_1005,N_297,N_16);
and U1006 (N_1006,N_318,N_981);
and U1007 (N_1007,N_161,N_534);
or U1008 (N_1008,N_904,N_822);
nor U1009 (N_1009,N_37,N_125);
nand U1010 (N_1010,N_739,N_735);
nand U1011 (N_1011,N_921,N_75);
nand U1012 (N_1012,N_698,N_238);
and U1013 (N_1013,N_793,N_743);
nand U1014 (N_1014,N_758,N_986);
nor U1015 (N_1015,N_127,N_442);
nand U1016 (N_1016,N_109,N_448);
nand U1017 (N_1017,N_403,N_253);
or U1018 (N_1018,N_311,N_36);
nor U1019 (N_1019,N_639,N_540);
nor U1020 (N_1020,N_485,N_126);
nand U1021 (N_1021,N_86,N_688);
nand U1022 (N_1022,N_672,N_531);
nor U1023 (N_1023,N_997,N_953);
or U1024 (N_1024,N_992,N_814);
and U1025 (N_1025,N_665,N_736);
nor U1026 (N_1026,N_434,N_930);
or U1027 (N_1027,N_291,N_595);
nor U1028 (N_1028,N_156,N_709);
nor U1029 (N_1029,N_447,N_101);
and U1030 (N_1030,N_430,N_742);
or U1031 (N_1031,N_611,N_791);
nand U1032 (N_1032,N_298,N_487);
or U1033 (N_1033,N_121,N_287);
or U1034 (N_1034,N_124,N_79);
or U1035 (N_1035,N_932,N_556);
nand U1036 (N_1036,N_280,N_623);
nor U1037 (N_1037,N_535,N_25);
nand U1038 (N_1038,N_105,N_585);
or U1039 (N_1039,N_984,N_372);
and U1040 (N_1040,N_234,N_54);
nor U1041 (N_1041,N_247,N_45);
nor U1042 (N_1042,N_444,N_693);
or U1043 (N_1043,N_482,N_259);
nor U1044 (N_1044,N_393,N_154);
and U1045 (N_1045,N_569,N_972);
nor U1046 (N_1046,N_166,N_660);
and U1047 (N_1047,N_231,N_590);
and U1048 (N_1048,N_870,N_950);
nand U1049 (N_1049,N_301,N_478);
or U1050 (N_1050,N_51,N_788);
nand U1051 (N_1051,N_453,N_613);
nand U1052 (N_1052,N_634,N_469);
or U1053 (N_1053,N_172,N_23);
or U1054 (N_1054,N_865,N_21);
nor U1055 (N_1055,N_420,N_142);
or U1056 (N_1056,N_66,N_371);
or U1057 (N_1057,N_927,N_83);
nor U1058 (N_1058,N_451,N_705);
nor U1059 (N_1059,N_271,N_587);
nand U1060 (N_1060,N_302,N_431);
nand U1061 (N_1061,N_668,N_11);
nor U1062 (N_1062,N_446,N_602);
nand U1063 (N_1063,N_409,N_356);
and U1064 (N_1064,N_770,N_53);
or U1065 (N_1065,N_164,N_237);
or U1066 (N_1066,N_220,N_324);
nor U1067 (N_1067,N_339,N_85);
and U1068 (N_1068,N_648,N_171);
or U1069 (N_1069,N_362,N_454);
nor U1070 (N_1070,N_706,N_143);
and U1071 (N_1071,N_946,N_601);
or U1072 (N_1072,N_240,N_94);
nand U1073 (N_1073,N_527,N_279);
or U1074 (N_1074,N_727,N_398);
or U1075 (N_1075,N_781,N_522);
or U1076 (N_1076,N_110,N_98);
nor U1077 (N_1077,N_797,N_82);
nand U1078 (N_1078,N_348,N_182);
xor U1079 (N_1079,N_394,N_296);
or U1080 (N_1080,N_330,N_22);
nor U1081 (N_1081,N_757,N_428);
or U1082 (N_1082,N_285,N_504);
and U1083 (N_1083,N_103,N_461);
nor U1084 (N_1084,N_881,N_900);
and U1085 (N_1085,N_963,N_913);
nor U1086 (N_1086,N_872,N_708);
or U1087 (N_1087,N_26,N_303);
nor U1088 (N_1088,N_286,N_7);
nand U1089 (N_1089,N_955,N_32);
nor U1090 (N_1090,N_951,N_242);
or U1091 (N_1091,N_979,N_112);
and U1092 (N_1092,N_783,N_333);
nor U1093 (N_1093,N_191,N_670);
and U1094 (N_1094,N_879,N_738);
or U1095 (N_1095,N_939,N_489);
or U1096 (N_1096,N_961,N_857);
nor U1097 (N_1097,N_364,N_580);
or U1098 (N_1098,N_549,N_654);
nor U1099 (N_1099,N_873,N_929);
nor U1100 (N_1100,N_265,N_490);
nand U1101 (N_1101,N_379,N_412);
nand U1102 (N_1102,N_799,N_519);
nand U1103 (N_1103,N_404,N_667);
and U1104 (N_1104,N_185,N_355);
nor U1105 (N_1105,N_871,N_619);
nor U1106 (N_1106,N_565,N_294);
and U1107 (N_1107,N_532,N_254);
nand U1108 (N_1108,N_811,N_851);
and U1109 (N_1109,N_307,N_643);
or U1110 (N_1110,N_530,N_855);
nor U1111 (N_1111,N_924,N_544);
nand U1112 (N_1112,N_69,N_600);
nand U1113 (N_1113,N_861,N_267);
and U1114 (N_1114,N_815,N_392);
nand U1115 (N_1115,N_366,N_903);
nand U1116 (N_1116,N_713,N_244);
nand U1117 (N_1117,N_258,N_422);
or U1118 (N_1118,N_440,N_803);
nor U1119 (N_1119,N_644,N_397);
or U1120 (N_1120,N_503,N_180);
and U1121 (N_1121,N_222,N_141);
nand U1122 (N_1122,N_876,N_9);
and U1123 (N_1123,N_957,N_774);
nor U1124 (N_1124,N_342,N_157);
nand U1125 (N_1125,N_831,N_304);
and U1126 (N_1126,N_889,N_678);
nor U1127 (N_1127,N_306,N_860);
nor U1128 (N_1128,N_849,N_848);
or U1129 (N_1129,N_377,N_862);
nor U1130 (N_1130,N_335,N_223);
nand U1131 (N_1131,N_382,N_612);
nand U1132 (N_1132,N_495,N_173);
nand U1133 (N_1133,N_933,N_64);
and U1134 (N_1134,N_17,N_836);
and U1135 (N_1135,N_571,N_970);
or U1136 (N_1136,N_880,N_31);
or U1137 (N_1137,N_754,N_59);
or U1138 (N_1138,N_943,N_29);
nand U1139 (N_1139,N_91,N_218);
and U1140 (N_1140,N_902,N_61);
nand U1141 (N_1141,N_381,N_895);
nand U1142 (N_1142,N_977,N_15);
and U1143 (N_1143,N_472,N_959);
nand U1144 (N_1144,N_789,N_837);
or U1145 (N_1145,N_133,N_177);
or U1146 (N_1146,N_236,N_329);
nand U1147 (N_1147,N_777,N_87);
and U1148 (N_1148,N_67,N_796);
nor U1149 (N_1149,N_426,N_194);
nand U1150 (N_1150,N_58,N_875);
nor U1151 (N_1151,N_740,N_694);
nor U1152 (N_1152,N_81,N_771);
nor U1153 (N_1153,N_989,N_609);
nor U1154 (N_1154,N_720,N_883);
nand U1155 (N_1155,N_724,N_547);
and U1156 (N_1156,N_856,N_834);
and U1157 (N_1157,N_948,N_456);
nand U1158 (N_1158,N_92,N_846);
nor U1159 (N_1159,N_391,N_923);
or U1160 (N_1160,N_685,N_460);
nor U1161 (N_1161,N_251,N_407);
or U1162 (N_1162,N_671,N_228);
nand U1163 (N_1163,N_471,N_564);
or U1164 (N_1164,N_618,N_443);
nand U1165 (N_1165,N_716,N_317);
or U1166 (N_1166,N_570,N_597);
or U1167 (N_1167,N_212,N_260);
and U1168 (N_1168,N_369,N_589);
nand U1169 (N_1169,N_859,N_802);
nor U1170 (N_1170,N_541,N_683);
nand U1171 (N_1171,N_353,N_293);
and U1172 (N_1172,N_807,N_792);
or U1173 (N_1173,N_195,N_120);
nand U1174 (N_1174,N_512,N_367);
and U1175 (N_1175,N_405,N_40);
or U1176 (N_1176,N_310,N_901);
nand U1177 (N_1177,N_89,N_843);
nor U1178 (N_1178,N_484,N_136);
nand U1179 (N_1179,N_332,N_664);
and U1180 (N_1180,N_388,N_973);
and U1181 (N_1181,N_196,N_213);
nor U1182 (N_1182,N_681,N_906);
nand U1183 (N_1183,N_934,N_731);
nor U1184 (N_1184,N_579,N_548);
nand U1185 (N_1185,N_582,N_290);
and U1186 (N_1186,N_493,N_625);
and U1187 (N_1187,N_780,N_937);
and U1188 (N_1188,N_5,N_123);
nand U1189 (N_1189,N_358,N_4);
nor U1190 (N_1190,N_514,N_555);
or U1191 (N_1191,N_315,N_562);
nor U1192 (N_1192,N_760,N_956);
or U1193 (N_1193,N_275,N_631);
or U1194 (N_1194,N_563,N_877);
xnor U1195 (N_1195,N_737,N_546);
nor U1196 (N_1196,N_113,N_354);
nor U1197 (N_1197,N_827,N_129);
nand U1198 (N_1198,N_536,N_55);
nor U1199 (N_1199,N_622,N_163);
nand U1200 (N_1200,N_425,N_958);
nand U1201 (N_1201,N_656,N_229);
or U1202 (N_1202,N_114,N_516);
and U1203 (N_1203,N_626,N_717);
or U1204 (N_1204,N_429,N_928);
and U1205 (N_1205,N_373,N_918);
or U1206 (N_1206,N_219,N_414);
or U1207 (N_1207,N_752,N_842);
or U1208 (N_1208,N_474,N_349);
nand U1209 (N_1209,N_118,N_363);
and U1210 (N_1210,N_288,N_772);
nor U1211 (N_1211,N_614,N_808);
nand U1212 (N_1212,N_278,N_417);
nor U1213 (N_1213,N_633,N_636);
or U1214 (N_1214,N_581,N_277);
nor U1215 (N_1215,N_104,N_152);
nand U1216 (N_1216,N_554,N_284);
nand U1217 (N_1217,N_497,N_108);
or U1218 (N_1218,N_661,N_838);
or U1219 (N_1219,N_203,N_593);
nor U1220 (N_1220,N_140,N_350);
or U1221 (N_1221,N_520,N_427);
nand U1222 (N_1222,N_413,N_775);
and U1223 (N_1223,N_246,N_73);
nor U1224 (N_1224,N_749,N_224);
or U1225 (N_1225,N_305,N_494);
nor U1226 (N_1226,N_68,N_476);
or U1227 (N_1227,N_227,N_964);
nand U1228 (N_1228,N_620,N_441);
nand U1229 (N_1229,N_756,N_387);
nand U1230 (N_1230,N_262,N_696);
and U1231 (N_1231,N_715,N_276);
and U1232 (N_1232,N_359,N_887);
nand U1233 (N_1233,N_515,N_396);
and U1234 (N_1234,N_337,N_805);
nor U1235 (N_1235,N_35,N_217);
and U1236 (N_1236,N_341,N_647);
nand U1237 (N_1237,N_666,N_886);
nand U1238 (N_1238,N_576,N_817);
or U1239 (N_1239,N_847,N_769);
nor U1240 (N_1240,N_677,N_750);
nand U1241 (N_1241,N_88,N_583);
nor U1242 (N_1242,N_162,N_584);
or U1243 (N_1243,N_763,N_987);
and U1244 (N_1244,N_679,N_949);
or U1245 (N_1245,N_591,N_117);
or U1246 (N_1246,N_281,N_588);
or U1247 (N_1247,N_204,N_50);
nor U1248 (N_1248,N_825,N_607);
nor U1249 (N_1249,N_331,N_719);
or U1250 (N_1250,N_160,N_501);
or U1251 (N_1251,N_675,N_866);
nor U1252 (N_1252,N_410,N_508);
and U1253 (N_1253,N_13,N_197);
and U1254 (N_1254,N_76,N_663);
nand U1255 (N_1255,N_741,N_498);
and U1256 (N_1256,N_914,N_190);
nand U1257 (N_1257,N_971,N_319);
nand U1258 (N_1258,N_380,N_746);
and U1259 (N_1259,N_72,N_833);
or U1260 (N_1260,N_389,N_450);
and U1261 (N_1261,N_878,N_722);
and U1262 (N_1262,N_988,N_435);
nand U1263 (N_1263,N_686,N_189);
nor U1264 (N_1264,N_940,N_481);
nor U1265 (N_1265,N_557,N_506);
nand U1266 (N_1266,N_322,N_139);
nor U1267 (N_1267,N_947,N_261);
and U1268 (N_1268,N_432,N_888);
nor U1269 (N_1269,N_181,N_818);
nor U1270 (N_1270,N_210,N_813);
xor U1271 (N_1271,N_158,N_74);
nor U1272 (N_1272,N_159,N_682);
and U1273 (N_1273,N_151,N_8);
nand U1274 (N_1274,N_526,N_518);
nor U1275 (N_1275,N_840,N_605);
nor U1276 (N_1276,N_399,N_10);
nand U1277 (N_1277,N_952,N_199);
and U1278 (N_1278,N_216,N_457);
or U1279 (N_1279,N_561,N_386);
or U1280 (N_1280,N_823,N_835);
nor U1281 (N_1281,N_0,N_653);
or U1282 (N_1282,N_202,N_437);
nand U1283 (N_1283,N_149,N_603);
and U1284 (N_1284,N_703,N_455);
and U1285 (N_1285,N_909,N_744);
nor U1286 (N_1286,N_673,N_525);
and U1287 (N_1287,N_27,N_18);
nor U1288 (N_1288,N_662,N_300);
nor U1289 (N_1289,N_184,N_931);
nor U1290 (N_1290,N_374,N_965);
nand U1291 (N_1291,N_77,N_991);
nand U1292 (N_1292,N_325,N_637);
nand U1293 (N_1293,N_982,N_336);
or U1294 (N_1294,N_936,N_144);
nor U1295 (N_1295,N_630,N_491);
and U1296 (N_1296,N_542,N_378);
or U1297 (N_1297,N_208,N_274);
nand U1298 (N_1298,N_214,N_560);
nand U1299 (N_1299,N_852,N_776);
or U1300 (N_1300,N_44,N_773);
xnor U1301 (N_1301,N_375,N_523);
or U1302 (N_1302,N_916,N_14);
nor U1303 (N_1303,N_328,N_467);
nand U1304 (N_1304,N_46,N_733);
and U1305 (N_1305,N_463,N_608);
and U1306 (N_1306,N_233,N_211);
nand U1307 (N_1307,N_33,N_985);
nand U1308 (N_1308,N_134,N_48);
nor U1309 (N_1309,N_510,N_850);
and U1310 (N_1310,N_826,N_968);
or U1311 (N_1311,N_480,N_976);
or U1312 (N_1312,N_559,N_445);
nand U1313 (N_1313,N_812,N_568);
nor U1314 (N_1314,N_747,N_941);
nand U1315 (N_1315,N_778,N_995);
nand U1316 (N_1316,N_116,N_295);
nor U1317 (N_1317,N_299,N_500);
nand U1318 (N_1318,N_798,N_408);
or U1319 (N_1319,N_980,N_641);
and U1320 (N_1320,N_243,N_263);
nor U1321 (N_1321,N_321,N_174);
nand U1322 (N_1322,N_470,N_312);
and U1323 (N_1323,N_890,N_192);
nand U1324 (N_1324,N_135,N_674);
or U1325 (N_1325,N_994,N_41);
nand U1326 (N_1326,N_255,N_652);
nand U1327 (N_1327,N_699,N_894);
nor U1328 (N_1328,N_452,N_858);
nand U1329 (N_1329,N_748,N_509);
nor U1330 (N_1330,N_586,N_464);
and U1331 (N_1331,N_96,N_820);
and U1332 (N_1332,N_790,N_640);
or U1333 (N_1333,N_486,N_84);
nor U1334 (N_1334,N_248,N_800);
nor U1335 (N_1335,N_225,N_755);
nand U1336 (N_1336,N_221,N_95);
and U1337 (N_1337,N_567,N_400);
nor U1338 (N_1338,N_621,N_996);
and U1339 (N_1339,N_680,N_70);
or U1340 (N_1340,N_370,N_759);
and U1341 (N_1341,N_701,N_130);
nor U1342 (N_1342,N_944,N_967);
nand U1343 (N_1343,N_465,N_459);
nor U1344 (N_1344,N_659,N_438);
or U1345 (N_1345,N_292,N_642);
or U1346 (N_1346,N_638,N_175);
nand U1347 (N_1347,N_283,N_816);
nand U1348 (N_1348,N_543,N_176);
nor U1349 (N_1349,N_911,N_401);
nor U1350 (N_1350,N_645,N_264);
and U1351 (N_1351,N_726,N_867);
or U1352 (N_1352,N_360,N_115);
and U1353 (N_1353,N_723,N_801);
nor U1354 (N_1354,N_553,N_327);
nand U1355 (N_1355,N_926,N_572);
nor U1356 (N_1356,N_864,N_343);
nor U1357 (N_1357,N_891,N_153);
nor U1358 (N_1358,N_187,N_604);
and U1359 (N_1359,N_962,N_524);
and U1360 (N_1360,N_411,N_492);
nor U1361 (N_1361,N_969,N_80);
nand U1362 (N_1362,N_47,N_28);
nand U1363 (N_1363,N_320,N_999);
or U1364 (N_1364,N_30,N_863);
nor U1365 (N_1365,N_232,N_226);
xor U1366 (N_1366,N_131,N_167);
and U1367 (N_1367,N_517,N_138);
xor U1368 (N_1368,N_155,N_594);
or U1369 (N_1369,N_334,N_821);
nor U1370 (N_1370,N_868,N_71);
nand U1371 (N_1371,N_784,N_687);
nor U1372 (N_1372,N_418,N_178);
and U1373 (N_1373,N_468,N_599);
and U1374 (N_1374,N_819,N_235);
or U1375 (N_1375,N_869,N_462);
nor U1376 (N_1376,N_505,N_270);
nand U1377 (N_1377,N_145,N_632);
nand U1378 (N_1378,N_421,N_122);
nor U1379 (N_1379,N_782,N_201);
nand U1380 (N_1380,N_917,N_628);
nor U1381 (N_1381,N_853,N_545);
or U1382 (N_1382,N_316,N_684);
nand U1383 (N_1383,N_3,N_351);
or U1384 (N_1384,N_575,N_150);
and U1385 (N_1385,N_249,N_690);
nor U1386 (N_1386,N_954,N_97);
nand U1387 (N_1387,N_966,N_577);
nor U1388 (N_1388,N_712,N_179);
or U1389 (N_1389,N_323,N_721);
nor U1390 (N_1390,N_745,N_761);
xor U1391 (N_1391,N_313,N_24);
and U1392 (N_1392,N_925,N_795);
nor U1393 (N_1393,N_436,N_539);
nand U1394 (N_1394,N_475,N_975);
nand U1395 (N_1395,N_344,N_766);
and U1396 (N_1396,N_390,N_193);
and U1397 (N_1397,N_874,N_282);
nand U1398 (N_1398,N_406,N_882);
nor U1399 (N_1399,N_945,N_676);
nand U1400 (N_1400,N_458,N_768);
or U1401 (N_1401,N_49,N_148);
or U1402 (N_1402,N_919,N_692);
and U1403 (N_1403,N_188,N_829);
or U1404 (N_1404,N_206,N_198);
nand U1405 (N_1405,N_424,N_832);
nor U1406 (N_1406,N_93,N_43);
nand U1407 (N_1407,N_751,N_361);
nand U1408 (N_1408,N_786,N_804);
or U1409 (N_1409,N_528,N_938);
nand U1410 (N_1410,N_19,N_466);
nand U1411 (N_1411,N_252,N_896);
nor U1412 (N_1412,N_326,N_186);
and U1413 (N_1413,N_828,N_779);
and U1414 (N_1414,N_376,N_147);
and U1415 (N_1415,N_824,N_764);
or U1416 (N_1416,N_499,N_38);
and U1417 (N_1417,N_57,N_598);
and U1418 (N_1418,N_340,N_230);
or U1419 (N_1419,N_573,N_346);
nor U1420 (N_1420,N_646,N_711);
and U1421 (N_1421,N_689,N_978);
nor U1422 (N_1422,N_107,N_552);
and U1423 (N_1423,N_714,N_200);
nor U1424 (N_1424,N_702,N_566);
nand U1425 (N_1425,N_183,N_841);
nand U1426 (N_1426,N_423,N_592);
and U1427 (N_1427,N_650,N_132);
nand U1428 (N_1428,N_615,N_596);
nand U1429 (N_1429,N_710,N_106);
nand U1430 (N_1430,N_205,N_728);
xor U1431 (N_1431,N_993,N_250);
nand U1432 (N_1432,N_165,N_854);
nor U1433 (N_1433,N_357,N_697);
or U1434 (N_1434,N_990,N_617);
or U1435 (N_1435,N_922,N_257);
and U1436 (N_1436,N_245,N_215);
nand U1437 (N_1437,N_102,N_700);
or U1438 (N_1438,N_695,N_119);
nor U1439 (N_1439,N_496,N_395);
nand U1440 (N_1440,N_2,N_892);
nand U1441 (N_1441,N_60,N_170);
and U1442 (N_1442,N_624,N_998);
and U1443 (N_1443,N_657,N_111);
and U1444 (N_1444,N_146,N_209);
nand U1445 (N_1445,N_907,N_920);
nor U1446 (N_1446,N_785,N_905);
nand U1447 (N_1447,N_345,N_915);
nand U1448 (N_1448,N_90,N_935);
or U1449 (N_1449,N_753,N_551);
or U1450 (N_1450,N_616,N_787);
or U1451 (N_1451,N_488,N_239);
nand U1452 (N_1452,N_558,N_338);
and U1453 (N_1453,N_704,N_884);
nand U1454 (N_1454,N_42,N_734);
nand U1455 (N_1455,N_502,N_266);
nand U1456 (N_1456,N_385,N_610);
or U1457 (N_1457,N_352,N_794);
or U1458 (N_1458,N_899,N_629);
nand U1459 (N_1459,N_537,N_893);
nand U1460 (N_1460,N_691,N_384);
or U1461 (N_1461,N_809,N_730);
nor U1462 (N_1462,N_844,N_273);
xor U1463 (N_1463,N_56,N_433);
nand U1464 (N_1464,N_942,N_269);
nand U1465 (N_1465,N_402,N_62);
or U1466 (N_1466,N_908,N_449);
nor U1467 (N_1467,N_655,N_529);
nor U1468 (N_1468,N_839,N_415);
and U1469 (N_1469,N_479,N_983);
nor U1470 (N_1470,N_898,N_574);
nand U1471 (N_1471,N_272,N_810);
nand U1472 (N_1472,N_416,N_477);
or U1473 (N_1473,N_207,N_765);
nor U1474 (N_1474,N_78,N_606);
or U1475 (N_1475,N_20,N_473);
or U1476 (N_1476,N_6,N_63);
and U1477 (N_1477,N_806,N_39);
nand U1478 (N_1478,N_845,N_513);
nand U1479 (N_1479,N_511,N_635);
and U1480 (N_1480,N_974,N_12);
or U1481 (N_1481,N_578,N_533);
nor U1482 (N_1482,N_169,N_314);
and U1483 (N_1483,N_65,N_137);
nand U1484 (N_1484,N_897,N_669);
or U1485 (N_1485,N_718,N_725);
nor U1486 (N_1486,N_762,N_885);
nand U1487 (N_1487,N_99,N_830);
nor U1488 (N_1488,N_268,N_309);
nand U1489 (N_1489,N_168,N_960);
or U1490 (N_1490,N_289,N_538);
and U1491 (N_1491,N_128,N_483);
or U1492 (N_1492,N_651,N_912);
nor U1493 (N_1493,N_732,N_521);
or U1494 (N_1494,N_419,N_34);
nand U1495 (N_1495,N_368,N_910);
and U1496 (N_1496,N_52,N_256);
nor U1497 (N_1497,N_658,N_627);
nor U1498 (N_1498,N_550,N_100);
or U1499 (N_1499,N_308,N_507);
and U1500 (N_1500,N_565,N_978);
or U1501 (N_1501,N_457,N_616);
xnor U1502 (N_1502,N_374,N_768);
nand U1503 (N_1503,N_260,N_525);
nor U1504 (N_1504,N_32,N_172);
nor U1505 (N_1505,N_118,N_207);
nor U1506 (N_1506,N_786,N_150);
or U1507 (N_1507,N_223,N_143);
nor U1508 (N_1508,N_669,N_787);
or U1509 (N_1509,N_827,N_301);
nand U1510 (N_1510,N_66,N_915);
and U1511 (N_1511,N_323,N_739);
or U1512 (N_1512,N_45,N_28);
and U1513 (N_1513,N_708,N_478);
nand U1514 (N_1514,N_202,N_595);
and U1515 (N_1515,N_505,N_413);
or U1516 (N_1516,N_279,N_840);
nand U1517 (N_1517,N_822,N_350);
nand U1518 (N_1518,N_643,N_876);
nand U1519 (N_1519,N_284,N_736);
nand U1520 (N_1520,N_632,N_38);
nand U1521 (N_1521,N_630,N_485);
and U1522 (N_1522,N_779,N_709);
nor U1523 (N_1523,N_75,N_68);
nor U1524 (N_1524,N_896,N_430);
nand U1525 (N_1525,N_986,N_169);
or U1526 (N_1526,N_833,N_6);
or U1527 (N_1527,N_998,N_436);
or U1528 (N_1528,N_727,N_162);
and U1529 (N_1529,N_47,N_686);
nand U1530 (N_1530,N_111,N_989);
nor U1531 (N_1531,N_460,N_894);
nand U1532 (N_1532,N_385,N_35);
and U1533 (N_1533,N_257,N_284);
and U1534 (N_1534,N_149,N_414);
nand U1535 (N_1535,N_344,N_906);
nand U1536 (N_1536,N_990,N_23);
nand U1537 (N_1537,N_360,N_694);
nand U1538 (N_1538,N_815,N_522);
or U1539 (N_1539,N_114,N_629);
or U1540 (N_1540,N_996,N_498);
nor U1541 (N_1541,N_335,N_402);
nor U1542 (N_1542,N_700,N_524);
nor U1543 (N_1543,N_504,N_365);
or U1544 (N_1544,N_840,N_641);
nand U1545 (N_1545,N_491,N_512);
nand U1546 (N_1546,N_519,N_734);
and U1547 (N_1547,N_849,N_767);
nand U1548 (N_1548,N_511,N_462);
nor U1549 (N_1549,N_32,N_328);
and U1550 (N_1550,N_838,N_377);
or U1551 (N_1551,N_126,N_919);
or U1552 (N_1552,N_582,N_79);
nor U1553 (N_1553,N_31,N_722);
and U1554 (N_1554,N_462,N_89);
and U1555 (N_1555,N_845,N_257);
or U1556 (N_1556,N_137,N_714);
nor U1557 (N_1557,N_45,N_200);
or U1558 (N_1558,N_504,N_216);
xnor U1559 (N_1559,N_639,N_280);
and U1560 (N_1560,N_155,N_471);
nand U1561 (N_1561,N_540,N_28);
or U1562 (N_1562,N_826,N_794);
nand U1563 (N_1563,N_308,N_125);
nor U1564 (N_1564,N_304,N_164);
or U1565 (N_1565,N_554,N_356);
nor U1566 (N_1566,N_913,N_293);
and U1567 (N_1567,N_307,N_238);
or U1568 (N_1568,N_645,N_256);
nand U1569 (N_1569,N_650,N_926);
nor U1570 (N_1570,N_873,N_372);
nand U1571 (N_1571,N_498,N_223);
nor U1572 (N_1572,N_610,N_578);
or U1573 (N_1573,N_135,N_150);
and U1574 (N_1574,N_42,N_724);
or U1575 (N_1575,N_530,N_633);
and U1576 (N_1576,N_196,N_663);
and U1577 (N_1577,N_119,N_158);
and U1578 (N_1578,N_911,N_87);
and U1579 (N_1579,N_890,N_327);
nor U1580 (N_1580,N_84,N_697);
or U1581 (N_1581,N_411,N_285);
nand U1582 (N_1582,N_737,N_407);
nand U1583 (N_1583,N_383,N_958);
and U1584 (N_1584,N_153,N_561);
and U1585 (N_1585,N_974,N_601);
or U1586 (N_1586,N_486,N_311);
nor U1587 (N_1587,N_84,N_786);
or U1588 (N_1588,N_657,N_611);
and U1589 (N_1589,N_339,N_666);
and U1590 (N_1590,N_249,N_129);
nor U1591 (N_1591,N_58,N_291);
nor U1592 (N_1592,N_799,N_316);
nand U1593 (N_1593,N_258,N_830);
and U1594 (N_1594,N_677,N_133);
nor U1595 (N_1595,N_738,N_626);
and U1596 (N_1596,N_797,N_10);
nand U1597 (N_1597,N_965,N_607);
nand U1598 (N_1598,N_959,N_811);
nand U1599 (N_1599,N_859,N_880);
nand U1600 (N_1600,N_116,N_325);
or U1601 (N_1601,N_647,N_467);
or U1602 (N_1602,N_619,N_276);
nor U1603 (N_1603,N_363,N_217);
or U1604 (N_1604,N_242,N_478);
or U1605 (N_1605,N_894,N_131);
and U1606 (N_1606,N_733,N_622);
nor U1607 (N_1607,N_285,N_962);
nand U1608 (N_1608,N_102,N_285);
nor U1609 (N_1609,N_216,N_977);
nor U1610 (N_1610,N_23,N_341);
or U1611 (N_1611,N_175,N_177);
nor U1612 (N_1612,N_440,N_356);
nand U1613 (N_1613,N_782,N_316);
nor U1614 (N_1614,N_941,N_142);
nand U1615 (N_1615,N_513,N_574);
nor U1616 (N_1616,N_489,N_836);
nand U1617 (N_1617,N_3,N_86);
or U1618 (N_1618,N_500,N_292);
and U1619 (N_1619,N_396,N_295);
or U1620 (N_1620,N_969,N_403);
nor U1621 (N_1621,N_120,N_685);
or U1622 (N_1622,N_462,N_442);
nand U1623 (N_1623,N_401,N_773);
or U1624 (N_1624,N_969,N_189);
or U1625 (N_1625,N_801,N_337);
nand U1626 (N_1626,N_199,N_56);
or U1627 (N_1627,N_659,N_100);
nor U1628 (N_1628,N_436,N_616);
or U1629 (N_1629,N_314,N_72);
nand U1630 (N_1630,N_722,N_234);
xor U1631 (N_1631,N_304,N_828);
nand U1632 (N_1632,N_198,N_200);
and U1633 (N_1633,N_467,N_644);
or U1634 (N_1634,N_930,N_110);
and U1635 (N_1635,N_201,N_492);
and U1636 (N_1636,N_180,N_747);
and U1637 (N_1637,N_341,N_829);
nand U1638 (N_1638,N_463,N_73);
or U1639 (N_1639,N_232,N_826);
nor U1640 (N_1640,N_898,N_294);
and U1641 (N_1641,N_943,N_165);
nor U1642 (N_1642,N_814,N_511);
and U1643 (N_1643,N_799,N_541);
and U1644 (N_1644,N_934,N_214);
and U1645 (N_1645,N_686,N_533);
xor U1646 (N_1646,N_775,N_51);
nand U1647 (N_1647,N_980,N_360);
nor U1648 (N_1648,N_397,N_408);
nor U1649 (N_1649,N_854,N_349);
and U1650 (N_1650,N_610,N_954);
nand U1651 (N_1651,N_621,N_298);
nand U1652 (N_1652,N_229,N_727);
nand U1653 (N_1653,N_106,N_540);
nor U1654 (N_1654,N_247,N_15);
nand U1655 (N_1655,N_327,N_22);
or U1656 (N_1656,N_254,N_3);
nor U1657 (N_1657,N_531,N_838);
nor U1658 (N_1658,N_692,N_824);
or U1659 (N_1659,N_101,N_475);
nor U1660 (N_1660,N_343,N_945);
and U1661 (N_1661,N_992,N_223);
and U1662 (N_1662,N_276,N_329);
nor U1663 (N_1663,N_371,N_197);
nor U1664 (N_1664,N_400,N_431);
xor U1665 (N_1665,N_725,N_882);
nand U1666 (N_1666,N_376,N_991);
and U1667 (N_1667,N_997,N_139);
or U1668 (N_1668,N_221,N_958);
nor U1669 (N_1669,N_952,N_898);
nor U1670 (N_1670,N_886,N_888);
nor U1671 (N_1671,N_743,N_543);
or U1672 (N_1672,N_132,N_805);
or U1673 (N_1673,N_953,N_493);
or U1674 (N_1674,N_408,N_709);
or U1675 (N_1675,N_54,N_749);
nand U1676 (N_1676,N_673,N_532);
nor U1677 (N_1677,N_525,N_465);
or U1678 (N_1678,N_949,N_920);
nor U1679 (N_1679,N_348,N_941);
nand U1680 (N_1680,N_833,N_48);
or U1681 (N_1681,N_480,N_173);
nor U1682 (N_1682,N_406,N_211);
nand U1683 (N_1683,N_684,N_958);
nor U1684 (N_1684,N_666,N_707);
nor U1685 (N_1685,N_591,N_822);
nand U1686 (N_1686,N_530,N_78);
nand U1687 (N_1687,N_450,N_37);
or U1688 (N_1688,N_755,N_206);
nand U1689 (N_1689,N_449,N_51);
nor U1690 (N_1690,N_416,N_355);
nor U1691 (N_1691,N_758,N_891);
and U1692 (N_1692,N_303,N_609);
or U1693 (N_1693,N_864,N_773);
or U1694 (N_1694,N_153,N_795);
nor U1695 (N_1695,N_210,N_636);
or U1696 (N_1696,N_433,N_651);
and U1697 (N_1697,N_790,N_653);
or U1698 (N_1698,N_707,N_71);
and U1699 (N_1699,N_143,N_500);
nor U1700 (N_1700,N_625,N_991);
and U1701 (N_1701,N_512,N_456);
and U1702 (N_1702,N_709,N_865);
and U1703 (N_1703,N_80,N_551);
nand U1704 (N_1704,N_945,N_278);
nand U1705 (N_1705,N_858,N_58);
or U1706 (N_1706,N_238,N_781);
or U1707 (N_1707,N_644,N_718);
and U1708 (N_1708,N_976,N_795);
nand U1709 (N_1709,N_72,N_400);
and U1710 (N_1710,N_37,N_744);
nand U1711 (N_1711,N_455,N_789);
xor U1712 (N_1712,N_565,N_192);
or U1713 (N_1713,N_988,N_523);
and U1714 (N_1714,N_666,N_156);
nor U1715 (N_1715,N_202,N_466);
nor U1716 (N_1716,N_864,N_686);
nor U1717 (N_1717,N_28,N_329);
nand U1718 (N_1718,N_240,N_977);
nor U1719 (N_1719,N_418,N_144);
nand U1720 (N_1720,N_318,N_413);
and U1721 (N_1721,N_236,N_234);
nand U1722 (N_1722,N_801,N_351);
nor U1723 (N_1723,N_833,N_845);
nand U1724 (N_1724,N_853,N_286);
nand U1725 (N_1725,N_874,N_983);
nor U1726 (N_1726,N_913,N_555);
or U1727 (N_1727,N_137,N_22);
or U1728 (N_1728,N_865,N_720);
or U1729 (N_1729,N_557,N_641);
or U1730 (N_1730,N_611,N_850);
and U1731 (N_1731,N_403,N_727);
or U1732 (N_1732,N_532,N_456);
nor U1733 (N_1733,N_74,N_277);
and U1734 (N_1734,N_906,N_519);
or U1735 (N_1735,N_413,N_430);
or U1736 (N_1736,N_290,N_610);
or U1737 (N_1737,N_962,N_326);
or U1738 (N_1738,N_328,N_295);
or U1739 (N_1739,N_682,N_687);
xnor U1740 (N_1740,N_454,N_864);
or U1741 (N_1741,N_497,N_104);
nor U1742 (N_1742,N_341,N_527);
or U1743 (N_1743,N_193,N_986);
or U1744 (N_1744,N_363,N_336);
nand U1745 (N_1745,N_901,N_125);
or U1746 (N_1746,N_948,N_789);
nand U1747 (N_1747,N_343,N_73);
xor U1748 (N_1748,N_686,N_829);
and U1749 (N_1749,N_958,N_766);
and U1750 (N_1750,N_301,N_780);
or U1751 (N_1751,N_521,N_937);
nor U1752 (N_1752,N_444,N_666);
nor U1753 (N_1753,N_357,N_191);
and U1754 (N_1754,N_871,N_292);
nor U1755 (N_1755,N_773,N_331);
and U1756 (N_1756,N_570,N_132);
and U1757 (N_1757,N_558,N_269);
nor U1758 (N_1758,N_778,N_83);
and U1759 (N_1759,N_485,N_610);
or U1760 (N_1760,N_781,N_737);
or U1761 (N_1761,N_890,N_755);
nor U1762 (N_1762,N_984,N_163);
nand U1763 (N_1763,N_163,N_951);
nor U1764 (N_1764,N_589,N_615);
xnor U1765 (N_1765,N_920,N_401);
and U1766 (N_1766,N_441,N_796);
and U1767 (N_1767,N_141,N_548);
or U1768 (N_1768,N_125,N_258);
or U1769 (N_1769,N_481,N_649);
and U1770 (N_1770,N_75,N_761);
or U1771 (N_1771,N_334,N_686);
and U1772 (N_1772,N_977,N_6);
or U1773 (N_1773,N_326,N_197);
nand U1774 (N_1774,N_360,N_545);
and U1775 (N_1775,N_709,N_864);
or U1776 (N_1776,N_393,N_181);
and U1777 (N_1777,N_18,N_841);
nand U1778 (N_1778,N_987,N_723);
nor U1779 (N_1779,N_335,N_953);
nand U1780 (N_1780,N_388,N_19);
nor U1781 (N_1781,N_332,N_445);
nand U1782 (N_1782,N_773,N_532);
nor U1783 (N_1783,N_607,N_508);
and U1784 (N_1784,N_432,N_385);
or U1785 (N_1785,N_46,N_706);
nand U1786 (N_1786,N_886,N_200);
and U1787 (N_1787,N_616,N_138);
or U1788 (N_1788,N_464,N_852);
nand U1789 (N_1789,N_799,N_310);
nor U1790 (N_1790,N_442,N_735);
or U1791 (N_1791,N_154,N_266);
nand U1792 (N_1792,N_212,N_711);
nand U1793 (N_1793,N_874,N_128);
nand U1794 (N_1794,N_9,N_197);
and U1795 (N_1795,N_523,N_524);
and U1796 (N_1796,N_879,N_142);
nor U1797 (N_1797,N_171,N_373);
or U1798 (N_1798,N_135,N_884);
nor U1799 (N_1799,N_810,N_648);
and U1800 (N_1800,N_116,N_149);
nand U1801 (N_1801,N_338,N_444);
nand U1802 (N_1802,N_857,N_669);
and U1803 (N_1803,N_791,N_401);
or U1804 (N_1804,N_90,N_554);
nand U1805 (N_1805,N_774,N_813);
nand U1806 (N_1806,N_971,N_74);
nand U1807 (N_1807,N_257,N_156);
or U1808 (N_1808,N_658,N_564);
or U1809 (N_1809,N_733,N_237);
nor U1810 (N_1810,N_644,N_599);
and U1811 (N_1811,N_118,N_569);
nor U1812 (N_1812,N_684,N_242);
or U1813 (N_1813,N_344,N_681);
nor U1814 (N_1814,N_480,N_283);
and U1815 (N_1815,N_330,N_435);
and U1816 (N_1816,N_944,N_453);
and U1817 (N_1817,N_235,N_122);
or U1818 (N_1818,N_690,N_405);
and U1819 (N_1819,N_890,N_594);
nand U1820 (N_1820,N_367,N_913);
nand U1821 (N_1821,N_762,N_62);
nand U1822 (N_1822,N_604,N_132);
and U1823 (N_1823,N_709,N_713);
or U1824 (N_1824,N_895,N_356);
nand U1825 (N_1825,N_172,N_423);
nor U1826 (N_1826,N_636,N_480);
or U1827 (N_1827,N_132,N_876);
nand U1828 (N_1828,N_686,N_446);
nand U1829 (N_1829,N_935,N_579);
nor U1830 (N_1830,N_81,N_836);
nand U1831 (N_1831,N_674,N_33);
and U1832 (N_1832,N_649,N_346);
nand U1833 (N_1833,N_311,N_966);
or U1834 (N_1834,N_994,N_931);
nand U1835 (N_1835,N_2,N_922);
nor U1836 (N_1836,N_710,N_937);
nor U1837 (N_1837,N_604,N_150);
nand U1838 (N_1838,N_486,N_179);
nand U1839 (N_1839,N_460,N_436);
or U1840 (N_1840,N_538,N_668);
and U1841 (N_1841,N_936,N_721);
nor U1842 (N_1842,N_835,N_729);
and U1843 (N_1843,N_464,N_634);
nand U1844 (N_1844,N_984,N_800);
nor U1845 (N_1845,N_214,N_735);
nor U1846 (N_1846,N_112,N_395);
nor U1847 (N_1847,N_40,N_4);
nand U1848 (N_1848,N_113,N_174);
and U1849 (N_1849,N_372,N_35);
and U1850 (N_1850,N_177,N_590);
and U1851 (N_1851,N_458,N_644);
or U1852 (N_1852,N_737,N_617);
or U1853 (N_1853,N_679,N_198);
and U1854 (N_1854,N_889,N_555);
nor U1855 (N_1855,N_569,N_585);
nand U1856 (N_1856,N_55,N_99);
and U1857 (N_1857,N_923,N_109);
nand U1858 (N_1858,N_723,N_667);
or U1859 (N_1859,N_176,N_598);
and U1860 (N_1860,N_94,N_808);
and U1861 (N_1861,N_108,N_78);
nand U1862 (N_1862,N_602,N_285);
nand U1863 (N_1863,N_679,N_637);
nand U1864 (N_1864,N_374,N_644);
or U1865 (N_1865,N_433,N_465);
nor U1866 (N_1866,N_530,N_808);
or U1867 (N_1867,N_717,N_94);
nor U1868 (N_1868,N_637,N_46);
nor U1869 (N_1869,N_690,N_497);
nor U1870 (N_1870,N_453,N_829);
and U1871 (N_1871,N_319,N_817);
and U1872 (N_1872,N_662,N_713);
or U1873 (N_1873,N_104,N_990);
or U1874 (N_1874,N_808,N_874);
and U1875 (N_1875,N_941,N_651);
nor U1876 (N_1876,N_11,N_517);
or U1877 (N_1877,N_521,N_601);
nand U1878 (N_1878,N_402,N_0);
nand U1879 (N_1879,N_916,N_81);
nand U1880 (N_1880,N_948,N_664);
and U1881 (N_1881,N_535,N_600);
or U1882 (N_1882,N_250,N_327);
nand U1883 (N_1883,N_323,N_59);
or U1884 (N_1884,N_249,N_482);
nor U1885 (N_1885,N_439,N_996);
and U1886 (N_1886,N_755,N_20);
or U1887 (N_1887,N_929,N_703);
nand U1888 (N_1888,N_49,N_730);
nand U1889 (N_1889,N_304,N_415);
nor U1890 (N_1890,N_875,N_299);
and U1891 (N_1891,N_240,N_75);
and U1892 (N_1892,N_964,N_29);
nand U1893 (N_1893,N_563,N_791);
nor U1894 (N_1894,N_872,N_346);
or U1895 (N_1895,N_685,N_706);
and U1896 (N_1896,N_312,N_871);
and U1897 (N_1897,N_316,N_168);
and U1898 (N_1898,N_266,N_418);
nor U1899 (N_1899,N_692,N_517);
nor U1900 (N_1900,N_336,N_951);
or U1901 (N_1901,N_702,N_393);
nor U1902 (N_1902,N_725,N_160);
and U1903 (N_1903,N_486,N_771);
nor U1904 (N_1904,N_822,N_951);
and U1905 (N_1905,N_699,N_76);
and U1906 (N_1906,N_98,N_246);
or U1907 (N_1907,N_512,N_742);
and U1908 (N_1908,N_549,N_942);
and U1909 (N_1909,N_691,N_183);
and U1910 (N_1910,N_689,N_486);
and U1911 (N_1911,N_295,N_885);
nor U1912 (N_1912,N_136,N_52);
nand U1913 (N_1913,N_916,N_384);
and U1914 (N_1914,N_902,N_453);
xnor U1915 (N_1915,N_358,N_632);
nand U1916 (N_1916,N_322,N_529);
nor U1917 (N_1917,N_516,N_167);
nand U1918 (N_1918,N_86,N_588);
and U1919 (N_1919,N_121,N_507);
or U1920 (N_1920,N_360,N_713);
nor U1921 (N_1921,N_202,N_482);
nand U1922 (N_1922,N_923,N_679);
nor U1923 (N_1923,N_609,N_122);
nand U1924 (N_1924,N_941,N_880);
nor U1925 (N_1925,N_975,N_280);
and U1926 (N_1926,N_683,N_675);
and U1927 (N_1927,N_941,N_374);
nor U1928 (N_1928,N_449,N_967);
or U1929 (N_1929,N_278,N_309);
or U1930 (N_1930,N_183,N_382);
nor U1931 (N_1931,N_357,N_672);
nor U1932 (N_1932,N_776,N_761);
and U1933 (N_1933,N_480,N_250);
nand U1934 (N_1934,N_557,N_620);
nor U1935 (N_1935,N_947,N_602);
and U1936 (N_1936,N_624,N_422);
or U1937 (N_1937,N_657,N_954);
nor U1938 (N_1938,N_286,N_267);
nor U1939 (N_1939,N_633,N_487);
or U1940 (N_1940,N_149,N_922);
nor U1941 (N_1941,N_881,N_581);
nand U1942 (N_1942,N_456,N_466);
and U1943 (N_1943,N_100,N_731);
and U1944 (N_1944,N_427,N_91);
nor U1945 (N_1945,N_340,N_108);
nor U1946 (N_1946,N_865,N_238);
or U1947 (N_1947,N_348,N_805);
or U1948 (N_1948,N_452,N_655);
and U1949 (N_1949,N_745,N_400);
nor U1950 (N_1950,N_249,N_507);
or U1951 (N_1951,N_2,N_20);
and U1952 (N_1952,N_676,N_380);
or U1953 (N_1953,N_601,N_276);
and U1954 (N_1954,N_172,N_251);
and U1955 (N_1955,N_386,N_820);
and U1956 (N_1956,N_564,N_583);
nor U1957 (N_1957,N_74,N_988);
nor U1958 (N_1958,N_378,N_268);
nor U1959 (N_1959,N_530,N_979);
or U1960 (N_1960,N_883,N_419);
nor U1961 (N_1961,N_208,N_574);
and U1962 (N_1962,N_75,N_19);
nor U1963 (N_1963,N_455,N_600);
nor U1964 (N_1964,N_680,N_168);
or U1965 (N_1965,N_413,N_441);
and U1966 (N_1966,N_763,N_390);
nand U1967 (N_1967,N_198,N_709);
or U1968 (N_1968,N_487,N_613);
and U1969 (N_1969,N_349,N_506);
nand U1970 (N_1970,N_69,N_743);
nor U1971 (N_1971,N_90,N_599);
nand U1972 (N_1972,N_39,N_943);
nor U1973 (N_1973,N_705,N_329);
and U1974 (N_1974,N_73,N_912);
or U1975 (N_1975,N_766,N_0);
and U1976 (N_1976,N_141,N_281);
nand U1977 (N_1977,N_669,N_766);
nor U1978 (N_1978,N_779,N_960);
and U1979 (N_1979,N_833,N_974);
or U1980 (N_1980,N_497,N_565);
nor U1981 (N_1981,N_306,N_583);
and U1982 (N_1982,N_36,N_205);
and U1983 (N_1983,N_887,N_890);
nand U1984 (N_1984,N_238,N_606);
and U1985 (N_1985,N_642,N_550);
nor U1986 (N_1986,N_836,N_980);
and U1987 (N_1987,N_522,N_987);
or U1988 (N_1988,N_495,N_231);
and U1989 (N_1989,N_189,N_154);
and U1990 (N_1990,N_890,N_257);
and U1991 (N_1991,N_515,N_768);
and U1992 (N_1992,N_926,N_978);
or U1993 (N_1993,N_308,N_574);
nor U1994 (N_1994,N_742,N_861);
or U1995 (N_1995,N_578,N_171);
or U1996 (N_1996,N_693,N_145);
nand U1997 (N_1997,N_238,N_354);
nor U1998 (N_1998,N_186,N_901);
nand U1999 (N_1999,N_565,N_510);
or U2000 (N_2000,N_1321,N_1238);
and U2001 (N_2001,N_1060,N_1093);
and U2002 (N_2002,N_1215,N_1863);
or U2003 (N_2003,N_1332,N_1067);
nor U2004 (N_2004,N_1888,N_1902);
nand U2005 (N_2005,N_1778,N_1715);
and U2006 (N_2006,N_1058,N_1887);
nand U2007 (N_2007,N_1520,N_1550);
nand U2008 (N_2008,N_1081,N_1099);
xor U2009 (N_2009,N_1515,N_1757);
and U2010 (N_2010,N_1160,N_1442);
and U2011 (N_2011,N_1454,N_1944);
or U2012 (N_2012,N_1236,N_1175);
nand U2013 (N_2013,N_1849,N_1387);
nand U2014 (N_2014,N_1028,N_1064);
or U2015 (N_2015,N_1304,N_1930);
nor U2016 (N_2016,N_1226,N_1085);
nor U2017 (N_2017,N_1068,N_1114);
and U2018 (N_2018,N_1137,N_1300);
or U2019 (N_2019,N_1980,N_1203);
nor U2020 (N_2020,N_1135,N_1531);
nor U2021 (N_2021,N_1674,N_1499);
nand U2022 (N_2022,N_1760,N_1087);
or U2023 (N_2023,N_1590,N_1517);
nor U2024 (N_2024,N_1919,N_1649);
or U2025 (N_2025,N_1325,N_1637);
nand U2026 (N_2026,N_1726,N_1047);
xnor U2027 (N_2027,N_1889,N_1864);
and U2028 (N_2028,N_1310,N_1982);
and U2029 (N_2029,N_1315,N_1630);
nand U2030 (N_2030,N_1577,N_1861);
or U2031 (N_2031,N_1307,N_1014);
nand U2032 (N_2032,N_1736,N_1992);
nand U2033 (N_2033,N_1822,N_1122);
and U2034 (N_2034,N_1188,N_1783);
nor U2035 (N_2035,N_1032,N_1868);
nand U2036 (N_2036,N_1573,N_1999);
nor U2037 (N_2037,N_1927,N_1460);
and U2038 (N_2038,N_1611,N_1580);
nor U2039 (N_2039,N_1240,N_1554);
nor U2040 (N_2040,N_1616,N_1832);
nor U2041 (N_2041,N_1125,N_1129);
nand U2042 (N_2042,N_1224,N_1324);
or U2043 (N_2043,N_1034,N_1467);
and U2044 (N_2044,N_1192,N_1937);
nor U2045 (N_2045,N_1483,N_1260);
nor U2046 (N_2046,N_1433,N_1190);
nand U2047 (N_2047,N_1294,N_1311);
xor U2048 (N_2048,N_1742,N_1322);
nor U2049 (N_2049,N_1645,N_1801);
nand U2050 (N_2050,N_1660,N_1666);
or U2051 (N_2051,N_1512,N_1052);
nor U2052 (N_2052,N_1024,N_1837);
and U2053 (N_2053,N_1417,N_1705);
or U2054 (N_2054,N_1487,N_1373);
or U2055 (N_2055,N_1116,N_1128);
nor U2056 (N_2056,N_1186,N_1010);
and U2057 (N_2057,N_1316,N_1003);
and U2058 (N_2058,N_1252,N_1039);
nand U2059 (N_2059,N_1143,N_1042);
nand U2060 (N_2060,N_1139,N_1342);
and U2061 (N_2061,N_1273,N_1308);
nand U2062 (N_2062,N_1289,N_1918);
nor U2063 (N_2063,N_1366,N_1117);
nand U2064 (N_2064,N_1400,N_1299);
or U2065 (N_2065,N_1495,N_1473);
and U2066 (N_2066,N_1636,N_1663);
xnor U2067 (N_2067,N_1169,N_1770);
or U2068 (N_2068,N_1870,N_1676);
nand U2069 (N_2069,N_1302,N_1812);
and U2070 (N_2070,N_1256,N_1920);
or U2071 (N_2071,N_1277,N_1865);
or U2072 (N_2072,N_1481,N_1365);
and U2073 (N_2073,N_1205,N_1876);
and U2074 (N_2074,N_1108,N_1838);
nand U2075 (N_2075,N_1072,N_1288);
or U2076 (N_2076,N_1267,N_1173);
nand U2077 (N_2077,N_1560,N_1412);
nand U2078 (N_2078,N_1800,N_1073);
nand U2079 (N_2079,N_1601,N_1303);
or U2080 (N_2080,N_1651,N_1065);
nor U2081 (N_2081,N_1624,N_1947);
nand U2082 (N_2082,N_1654,N_1023);
or U2083 (N_2083,N_1419,N_1562);
nand U2084 (N_2084,N_1568,N_1506);
and U2085 (N_2085,N_1179,N_1095);
or U2086 (N_2086,N_1270,N_1523);
or U2087 (N_2087,N_1713,N_1748);
and U2088 (N_2088,N_1813,N_1350);
nand U2089 (N_2089,N_1048,N_1271);
or U2090 (N_2090,N_1798,N_1153);
nor U2091 (N_2091,N_1700,N_1409);
nand U2092 (N_2092,N_1530,N_1981);
nor U2093 (N_2093,N_1607,N_1677);
and U2094 (N_2094,N_1606,N_1799);
and U2095 (N_2095,N_1111,N_1819);
nand U2096 (N_2096,N_1542,N_1695);
and U2097 (N_2097,N_1437,N_1806);
and U2098 (N_2098,N_1979,N_1132);
and U2099 (N_2099,N_1112,N_1591);
and U2100 (N_2100,N_1599,N_1589);
and U2101 (N_2101,N_1788,N_1848);
nor U2102 (N_2102,N_1885,N_1296);
nor U2103 (N_2103,N_1565,N_1519);
xor U2104 (N_2104,N_1445,N_1418);
and U2105 (N_2105,N_1040,N_1037);
nand U2106 (N_2106,N_1489,N_1723);
nand U2107 (N_2107,N_1490,N_1612);
and U2108 (N_2108,N_1976,N_1811);
or U2109 (N_2109,N_1362,N_1977);
nand U2110 (N_2110,N_1814,N_1435);
nor U2111 (N_2111,N_1463,N_1579);
nor U2112 (N_2112,N_1860,N_1582);
nand U2113 (N_2113,N_1873,N_1856);
nand U2114 (N_2114,N_1521,N_1793);
nor U2115 (N_2115,N_1540,N_1510);
or U2116 (N_2116,N_1056,N_1584);
nor U2117 (N_2117,N_1619,N_1142);
or U2118 (N_2118,N_1284,N_1281);
or U2119 (N_2119,N_1526,N_1767);
and U2120 (N_2120,N_1008,N_1451);
nor U2121 (N_2121,N_1941,N_1692);
nand U2122 (N_2122,N_1576,N_1535);
or U2123 (N_2123,N_1587,N_1368);
or U2124 (N_2124,N_1103,N_1079);
or U2125 (N_2125,N_1201,N_1274);
or U2126 (N_2126,N_1957,N_1853);
nor U2127 (N_2127,N_1675,N_1703);
nor U2128 (N_2128,N_1380,N_1198);
or U2129 (N_2129,N_1269,N_1776);
nand U2130 (N_2130,N_1900,N_1453);
and U2131 (N_2131,N_1007,N_1737);
nor U2132 (N_2132,N_1894,N_1431);
or U2133 (N_2133,N_1381,N_1493);
nor U2134 (N_2134,N_1686,N_1539);
and U2135 (N_2135,N_1295,N_1104);
or U2136 (N_2136,N_1263,N_1759);
and U2137 (N_2137,N_1457,N_1314);
or U2138 (N_2138,N_1815,N_1213);
or U2139 (N_2139,N_1916,N_1563);
or U2140 (N_2140,N_1009,N_1518);
nor U2141 (N_2141,N_1706,N_1633);
and U2142 (N_2142,N_1989,N_1136);
nand U2143 (N_2143,N_1155,N_1420);
nor U2144 (N_2144,N_1988,N_1396);
nor U2145 (N_2145,N_1758,N_1080);
nor U2146 (N_2146,N_1390,N_1209);
or U2147 (N_2147,N_1948,N_1242);
nand U2148 (N_2148,N_1780,N_1398);
or U2149 (N_2149,N_1344,N_1448);
nand U2150 (N_2150,N_1915,N_1212);
and U2151 (N_2151,N_1020,N_1075);
nor U2152 (N_2152,N_1874,N_1120);
or U2153 (N_2153,N_1334,N_1782);
nand U2154 (N_2154,N_1343,N_1702);
nor U2155 (N_2155,N_1346,N_1268);
nor U2156 (N_2156,N_1402,N_1679);
nor U2157 (N_2157,N_1422,N_1652);
nand U2158 (N_2158,N_1728,N_1834);
nor U2159 (N_2159,N_1041,N_1667);
nand U2160 (N_2160,N_1247,N_1393);
and U2161 (N_2161,N_1229,N_1914);
xnor U2162 (N_2162,N_1218,N_1347);
and U2163 (N_2163,N_1817,N_1045);
or U2164 (N_2164,N_1922,N_1985);
nand U2165 (N_2165,N_1846,N_1057);
and U2166 (N_2166,N_1527,N_1119);
nand U2167 (N_2167,N_1880,N_1464);
and U2168 (N_2168,N_1140,N_1642);
nand U2169 (N_2169,N_1000,N_1882);
nand U2170 (N_2170,N_1424,N_1395);
and U2171 (N_2171,N_1839,N_1282);
nand U2172 (N_2172,N_1397,N_1082);
and U2173 (N_2173,N_1069,N_1754);
nand U2174 (N_2174,N_1784,N_1115);
nand U2175 (N_2175,N_1379,N_1671);
and U2176 (N_2176,N_1878,N_1044);
nand U2177 (N_2177,N_1138,N_1995);
nand U2178 (N_2178,N_1908,N_1851);
nand U2179 (N_2179,N_1221,N_1855);
nor U2180 (N_2180,N_1275,N_1070);
or U2181 (N_2181,N_1144,N_1744);
nor U2182 (N_2182,N_1382,N_1475);
or U2183 (N_2183,N_1338,N_1643);
and U2184 (N_2184,N_1570,N_1195);
nor U2185 (N_2185,N_1762,N_1852);
nor U2186 (N_2186,N_1472,N_1792);
and U2187 (N_2187,N_1622,N_1763);
and U2188 (N_2188,N_1408,N_1732);
nor U2189 (N_2189,N_1353,N_1017);
nand U2190 (N_2190,N_1357,N_1216);
nor U2191 (N_2191,N_1638,N_1163);
nand U2192 (N_2192,N_1963,N_1808);
and U2193 (N_2193,N_1731,N_1548);
and U2194 (N_2194,N_1953,N_1339);
and U2195 (N_2195,N_1033,N_1912);
nor U2196 (N_2196,N_1745,N_1162);
nor U2197 (N_2197,N_1993,N_1425);
and U2198 (N_2198,N_1372,N_1447);
and U2199 (N_2199,N_1547,N_1484);
xnor U2200 (N_2200,N_1482,N_1022);
xor U2201 (N_2201,N_1336,N_1287);
or U2202 (N_2202,N_1461,N_1657);
nor U2203 (N_2203,N_1097,N_1553);
nor U2204 (N_2204,N_1413,N_1683);
and U2205 (N_2205,N_1796,N_1025);
and U2206 (N_2206,N_1335,N_1309);
and U2207 (N_2207,N_1363,N_1533);
and U2208 (N_2208,N_1978,N_1086);
nand U2209 (N_2209,N_1313,N_1890);
or U2210 (N_2210,N_1960,N_1439);
nor U2211 (N_2211,N_1791,N_1013);
nand U2212 (N_2212,N_1278,N_1625);
and U2213 (N_2213,N_1525,N_1857);
or U2214 (N_2214,N_1251,N_1771);
nand U2215 (N_2215,N_1248,N_1711);
and U2216 (N_2216,N_1572,N_1183);
or U2217 (N_2217,N_1661,N_1673);
nand U2218 (N_2218,N_1050,N_1756);
nor U2219 (N_2219,N_1426,N_1958);
and U2220 (N_2220,N_1641,N_1089);
nand U2221 (N_2221,N_1168,N_1323);
or U2222 (N_2222,N_1721,N_1502);
nand U2223 (N_2223,N_1741,N_1348);
nand U2224 (N_2224,N_1150,N_1388);
and U2225 (N_2225,N_1234,N_1593);
and U2226 (N_2226,N_1498,N_1018);
nor U2227 (N_2227,N_1789,N_1613);
nand U2228 (N_2228,N_1283,N_1730);
or U2229 (N_2229,N_1773,N_1015);
nand U2230 (N_2230,N_1997,N_1534);
nand U2231 (N_2231,N_1984,N_1991);
nand U2232 (N_2232,N_1739,N_1749);
or U2233 (N_2233,N_1990,N_1961);
and U2234 (N_2234,N_1331,N_1279);
and U2235 (N_2235,N_1765,N_1866);
nand U2236 (N_2236,N_1557,N_1441);
and U2237 (N_2237,N_1559,N_1290);
and U2238 (N_2238,N_1862,N_1006);
nand U2239 (N_2239,N_1516,N_1691);
nor U2240 (N_2240,N_1298,N_1965);
nor U2241 (N_2241,N_1002,N_1507);
nand U2242 (N_2242,N_1858,N_1131);
and U2243 (N_2243,N_1259,N_1219);
and U2244 (N_2244,N_1374,N_1197);
nor U2245 (N_2245,N_1462,N_1962);
and U2246 (N_2246,N_1149,N_1021);
and U2247 (N_2247,N_1297,N_1317);
nand U2248 (N_2248,N_1465,N_1508);
or U2249 (N_2249,N_1176,N_1476);
and U2250 (N_2250,N_1828,N_1090);
and U2251 (N_2251,N_1318,N_1126);
and U2252 (N_2252,N_1719,N_1578);
nand U2253 (N_2253,N_1551,N_1232);
or U2254 (N_2254,N_1102,N_1764);
and U2255 (N_2255,N_1355,N_1621);
or U2256 (N_2256,N_1614,N_1246);
or U2257 (N_2257,N_1967,N_1327);
nor U2258 (N_2258,N_1345,N_1609);
and U2259 (N_2259,N_1514,N_1200);
nand U2260 (N_2260,N_1301,N_1655);
or U2261 (N_2261,N_1955,N_1755);
nor U2262 (N_2262,N_1564,N_1012);
or U2263 (N_2263,N_1685,N_1061);
and U2264 (N_2264,N_1055,N_1471);
nand U2265 (N_2265,N_1959,N_1906);
and U2266 (N_2266,N_1053,N_1043);
and U2267 (N_2267,N_1222,N_1154);
and U2268 (N_2268,N_1171,N_1975);
or U2269 (N_2269,N_1193,N_1810);
nor U2270 (N_2270,N_1807,N_1233);
nand U2271 (N_2271,N_1257,N_1934);
nand U2272 (N_2272,N_1717,N_1123);
nor U2273 (N_2273,N_1932,N_1841);
and U2274 (N_2274,N_1797,N_1653);
xnor U2275 (N_2275,N_1320,N_1477);
nand U2276 (N_2276,N_1921,N_1378);
and U2277 (N_2277,N_1903,N_1091);
or U2278 (N_2278,N_1285,N_1604);
or U2279 (N_2279,N_1011,N_1970);
nor U2280 (N_2280,N_1896,N_1689);
and U2281 (N_2281,N_1805,N_1505);
nor U2282 (N_2282,N_1727,N_1494);
and U2283 (N_2283,N_1610,N_1648);
nand U2284 (N_2284,N_1708,N_1405);
or U2285 (N_2285,N_1913,N_1968);
or U2286 (N_2286,N_1480,N_1943);
and U2287 (N_2287,N_1907,N_1743);
nor U2288 (N_2288,N_1670,N_1062);
and U2289 (N_2289,N_1092,N_1333);
nand U2290 (N_2290,N_1261,N_1561);
and U2291 (N_2291,N_1174,N_1469);
or U2292 (N_2292,N_1650,N_1130);
nor U2293 (N_2293,N_1820,N_1898);
nand U2294 (N_2294,N_1950,N_1360);
xnor U2295 (N_2295,N_1833,N_1938);
nor U2296 (N_2296,N_1740,N_1468);
and U2297 (N_2297,N_1994,N_1133);
nand U2298 (N_2298,N_1196,N_1734);
or U2299 (N_2299,N_1931,N_1904);
or U2300 (N_2300,N_1935,N_1444);
and U2301 (N_2301,N_1694,N_1239);
nor U2302 (N_2302,N_1124,N_1210);
nand U2303 (N_2303,N_1600,N_1850);
nor U2304 (N_2304,N_1394,N_1432);
and U2305 (N_2305,N_1629,N_1871);
or U2306 (N_2306,N_1096,N_1172);
nor U2307 (N_2307,N_1255,N_1241);
nor U2308 (N_2308,N_1597,N_1078);
xor U2309 (N_2309,N_1720,N_1077);
and U2310 (N_2310,N_1501,N_1929);
or U2311 (N_2311,N_1566,N_1249);
or U2312 (N_2312,N_1787,N_1567);
or U2313 (N_2313,N_1485,N_1161);
nand U2314 (N_2314,N_1911,N_1421);
or U2315 (N_2315,N_1724,N_1802);
nand U2316 (N_2316,N_1752,N_1794);
nor U2317 (N_2317,N_1185,N_1735);
and U2318 (N_2318,N_1223,N_1076);
xnor U2319 (N_2319,N_1148,N_1291);
nor U2320 (N_2320,N_1046,N_1329);
or U2321 (N_2321,N_1359,N_1877);
or U2322 (N_2322,N_1410,N_1416);
nor U2323 (N_2323,N_1722,N_1714);
or U2324 (N_2324,N_1423,N_1134);
and U2325 (N_2325,N_1428,N_1971);
nor U2326 (N_2326,N_1987,N_1790);
or U2327 (N_2327,N_1693,N_1404);
xor U2328 (N_2328,N_1180,N_1823);
nand U2329 (N_2329,N_1774,N_1098);
or U2330 (N_2330,N_1225,N_1146);
and U2331 (N_2331,N_1066,N_1664);
nor U2332 (N_2332,N_1588,N_1895);
or U2333 (N_2333,N_1479,N_1503);
or U2334 (N_2334,N_1141,N_1051);
nand U2335 (N_2335,N_1513,N_1628);
and U2336 (N_2336,N_1795,N_1083);
nand U2337 (N_2337,N_1063,N_1030);
and U2338 (N_2338,N_1639,N_1933);
or U2339 (N_2339,N_1228,N_1549);
nor U2340 (N_2340,N_1825,N_1182);
or U2341 (N_2341,N_1556,N_1474);
or U2342 (N_2342,N_1964,N_1826);
nand U2343 (N_2343,N_1881,N_1019);
or U2344 (N_2344,N_1546,N_1293);
nand U2345 (N_2345,N_1376,N_1456);
or U2346 (N_2346,N_1905,N_1986);
nand U2347 (N_2347,N_1843,N_1709);
nor U2348 (N_2348,N_1504,N_1511);
and U2349 (N_2349,N_1227,N_1751);
and U2350 (N_2350,N_1646,N_1678);
nand U2351 (N_2351,N_1998,N_1429);
and U2352 (N_2352,N_1035,N_1330);
nor U2353 (N_2353,N_1319,N_1725);
and U2354 (N_2354,N_1753,N_1384);
and U2355 (N_2355,N_1158,N_1829);
nand U2356 (N_2356,N_1697,N_1258);
nor U2357 (N_2357,N_1237,N_1016);
and U2358 (N_2358,N_1665,N_1552);
and U2359 (N_2359,N_1152,N_1886);
nand U2360 (N_2360,N_1443,N_1687);
and U2361 (N_2361,N_1594,N_1167);
nand U2362 (N_2362,N_1875,N_1436);
nor U2363 (N_2363,N_1371,N_1220);
nor U2364 (N_2364,N_1901,N_1110);
and U2365 (N_2365,N_1956,N_1459);
or U2366 (N_2366,N_1544,N_1264);
and U2367 (N_2367,N_1105,N_1031);
and U2368 (N_2368,N_1383,N_1543);
and U2369 (N_2369,N_1524,N_1411);
nand U2370 (N_2370,N_1470,N_1377);
nand U2371 (N_2371,N_1718,N_1349);
nand U2372 (N_2372,N_1585,N_1969);
nand U2373 (N_2373,N_1541,N_1392);
nor U2374 (N_2374,N_1746,N_1569);
nand U2375 (N_2375,N_1157,N_1214);
nor U2376 (N_2376,N_1004,N_1954);
nand U2377 (N_2377,N_1438,N_1620);
and U2378 (N_2378,N_1681,N_1658);
and U2379 (N_2379,N_1974,N_1088);
nand U2380 (N_2380,N_1684,N_1391);
nand U2381 (N_2381,N_1603,N_1026);
nand U2382 (N_2382,N_1529,N_1450);
nor U2383 (N_2383,N_1364,N_1458);
or U2384 (N_2384,N_1434,N_1272);
nand U2385 (N_2385,N_1945,N_1243);
or U2386 (N_2386,N_1266,N_1352);
nor U2387 (N_2387,N_1199,N_1262);
nor U2388 (N_2388,N_1522,N_1027);
nand U2389 (N_2389,N_1414,N_1265);
or U2390 (N_2390,N_1084,N_1170);
xor U2391 (N_2391,N_1361,N_1254);
or U2392 (N_2392,N_1772,N_1710);
or U2393 (N_2393,N_1698,N_1113);
nor U2394 (N_2394,N_1250,N_1827);
nor U2395 (N_2395,N_1847,N_1761);
nand U2396 (N_2396,N_1049,N_1608);
nand U2397 (N_2397,N_1816,N_1165);
and U2398 (N_2398,N_1403,N_1766);
nor U2399 (N_2399,N_1845,N_1701);
nand U2400 (N_2400,N_1340,N_1151);
or U2401 (N_2401,N_1202,N_1777);
and U2402 (N_2402,N_1804,N_1109);
nand U2403 (N_2403,N_1656,N_1803);
or U2404 (N_2404,N_1926,N_1983);
or U2405 (N_2405,N_1029,N_1189);
nor U2406 (N_2406,N_1939,N_1245);
xnor U2407 (N_2407,N_1370,N_1235);
nor U2408 (N_2408,N_1538,N_1074);
nand U2409 (N_2409,N_1145,N_1107);
and U2410 (N_2410,N_1635,N_1399);
nand U2411 (N_2411,N_1207,N_1127);
nand U2412 (N_2412,N_1617,N_1688);
nor U2413 (N_2413,N_1716,N_1492);
or U2414 (N_2414,N_1821,N_1634);
nor U2415 (N_2415,N_1177,N_1647);
and U2416 (N_2416,N_1389,N_1769);
nand U2417 (N_2417,N_1872,N_1680);
or U2418 (N_2418,N_1292,N_1305);
nor U2419 (N_2419,N_1595,N_1286);
nor U2420 (N_2420,N_1500,N_1244);
nor U2421 (N_2421,N_1786,N_1231);
and U2422 (N_2422,N_1615,N_1312);
nor U2423 (N_2423,N_1101,N_1632);
nor U2424 (N_2424,N_1486,N_1623);
or U2425 (N_2425,N_1738,N_1407);
and U2426 (N_2426,N_1840,N_1528);
nand U2427 (N_2427,N_1672,N_1071);
and U2428 (N_2428,N_1690,N_1859);
nor U2429 (N_2429,N_1893,N_1415);
nor U2430 (N_2430,N_1750,N_1598);
or U2431 (N_2431,N_1488,N_1879);
nand U2432 (N_2432,N_1631,N_1536);
and U2433 (N_2433,N_1586,N_1181);
nand U2434 (N_2434,N_1949,N_1831);
or U2435 (N_2435,N_1712,N_1440);
or U2436 (N_2436,N_1351,N_1747);
or U2437 (N_2437,N_1869,N_1159);
nor U2438 (N_2438,N_1644,N_1166);
nor U2439 (N_2439,N_1618,N_1555);
nor U2440 (N_2440,N_1369,N_1147);
nor U2441 (N_2441,N_1899,N_1054);
and U2442 (N_2442,N_1867,N_1699);
nand U2443 (N_2443,N_1446,N_1537);
or U2444 (N_2444,N_1455,N_1118);
or U2445 (N_2445,N_1669,N_1707);
nand U2446 (N_2446,N_1809,N_1217);
nand U2447 (N_2447,N_1187,N_1972);
and U2448 (N_2448,N_1940,N_1966);
xnor U2449 (N_2449,N_1358,N_1781);
or U2450 (N_2450,N_1936,N_1696);
or U2451 (N_2451,N_1121,N_1592);
or U2452 (N_2452,N_1883,N_1909);
or U2453 (N_2453,N_1532,N_1897);
or U2454 (N_2454,N_1917,N_1306);
nand U2455 (N_2455,N_1640,N_1164);
nand U2456 (N_2456,N_1768,N_1581);
and U2457 (N_2457,N_1626,N_1452);
and U2458 (N_2458,N_1178,N_1005);
or U2459 (N_2459,N_1491,N_1682);
nor U2460 (N_2460,N_1659,N_1923);
nand U2461 (N_2461,N_1824,N_1211);
and U2462 (N_2462,N_1925,N_1558);
or U2463 (N_2463,N_1496,N_1942);
or U2464 (N_2464,N_1466,N_1204);
nor U2465 (N_2465,N_1497,N_1830);
and U2466 (N_2466,N_1337,N_1326);
and U2467 (N_2467,N_1430,N_1779);
nor U2468 (N_2468,N_1662,N_1952);
and U2469 (N_2469,N_1951,N_1844);
or U2470 (N_2470,N_1194,N_1106);
or U2471 (N_2471,N_1574,N_1509);
nor U2472 (N_2472,N_1910,N_1575);
nand U2473 (N_2473,N_1230,N_1094);
nor U2474 (N_2474,N_1733,N_1785);
nor U2475 (N_2475,N_1356,N_1602);
nor U2476 (N_2476,N_1605,N_1924);
or U2477 (N_2477,N_1835,N_1973);
or U2478 (N_2478,N_1818,N_1184);
xnor U2479 (N_2479,N_1253,N_1668);
and U2480 (N_2480,N_1328,N_1100);
and U2481 (N_2481,N_1367,N_1427);
or U2482 (N_2482,N_1996,N_1375);
and U2483 (N_2483,N_1449,N_1156);
and U2484 (N_2484,N_1884,N_1729);
or U2485 (N_2485,N_1627,N_1280);
xnor U2486 (N_2486,N_1036,N_1596);
nor U2487 (N_2487,N_1842,N_1583);
nand U2488 (N_2488,N_1038,N_1775);
or U2489 (N_2489,N_1406,N_1208);
nand U2490 (N_2490,N_1928,N_1341);
nor U2491 (N_2491,N_1892,N_1478);
and U2492 (N_2492,N_1354,N_1059);
nor U2493 (N_2493,N_1891,N_1854);
nor U2494 (N_2494,N_1401,N_1206);
and U2495 (N_2495,N_1836,N_1386);
or U2496 (N_2496,N_1001,N_1545);
or U2497 (N_2497,N_1704,N_1946);
nor U2498 (N_2498,N_1571,N_1191);
or U2499 (N_2499,N_1385,N_1276);
nand U2500 (N_2500,N_1878,N_1885);
or U2501 (N_2501,N_1966,N_1207);
or U2502 (N_2502,N_1081,N_1531);
or U2503 (N_2503,N_1356,N_1244);
nand U2504 (N_2504,N_1901,N_1277);
and U2505 (N_2505,N_1839,N_1235);
nor U2506 (N_2506,N_1335,N_1641);
nor U2507 (N_2507,N_1483,N_1669);
and U2508 (N_2508,N_1261,N_1127);
and U2509 (N_2509,N_1786,N_1176);
or U2510 (N_2510,N_1406,N_1891);
nor U2511 (N_2511,N_1010,N_1307);
or U2512 (N_2512,N_1396,N_1701);
or U2513 (N_2513,N_1868,N_1767);
nor U2514 (N_2514,N_1674,N_1187);
nand U2515 (N_2515,N_1375,N_1353);
nor U2516 (N_2516,N_1100,N_1901);
or U2517 (N_2517,N_1792,N_1571);
and U2518 (N_2518,N_1950,N_1572);
nor U2519 (N_2519,N_1940,N_1583);
or U2520 (N_2520,N_1337,N_1170);
nor U2521 (N_2521,N_1383,N_1717);
nand U2522 (N_2522,N_1701,N_1904);
or U2523 (N_2523,N_1320,N_1506);
and U2524 (N_2524,N_1687,N_1490);
or U2525 (N_2525,N_1617,N_1767);
and U2526 (N_2526,N_1058,N_1190);
nor U2527 (N_2527,N_1835,N_1494);
nor U2528 (N_2528,N_1119,N_1388);
and U2529 (N_2529,N_1267,N_1979);
nand U2530 (N_2530,N_1449,N_1023);
nand U2531 (N_2531,N_1537,N_1015);
or U2532 (N_2532,N_1626,N_1213);
or U2533 (N_2533,N_1369,N_1307);
and U2534 (N_2534,N_1326,N_1739);
and U2535 (N_2535,N_1020,N_1889);
nand U2536 (N_2536,N_1912,N_1734);
or U2537 (N_2537,N_1352,N_1693);
nor U2538 (N_2538,N_1479,N_1238);
nand U2539 (N_2539,N_1706,N_1198);
or U2540 (N_2540,N_1208,N_1575);
and U2541 (N_2541,N_1248,N_1833);
nand U2542 (N_2542,N_1793,N_1517);
nand U2543 (N_2543,N_1427,N_1269);
nand U2544 (N_2544,N_1066,N_1246);
and U2545 (N_2545,N_1625,N_1027);
nand U2546 (N_2546,N_1607,N_1843);
nand U2547 (N_2547,N_1186,N_1916);
and U2548 (N_2548,N_1644,N_1801);
nor U2549 (N_2549,N_1885,N_1943);
or U2550 (N_2550,N_1933,N_1340);
or U2551 (N_2551,N_1670,N_1287);
nand U2552 (N_2552,N_1374,N_1901);
nor U2553 (N_2553,N_1341,N_1815);
xnor U2554 (N_2554,N_1304,N_1574);
nand U2555 (N_2555,N_1651,N_1726);
and U2556 (N_2556,N_1506,N_1153);
nand U2557 (N_2557,N_1411,N_1462);
nor U2558 (N_2558,N_1098,N_1181);
nand U2559 (N_2559,N_1298,N_1245);
nor U2560 (N_2560,N_1415,N_1181);
and U2561 (N_2561,N_1566,N_1956);
or U2562 (N_2562,N_1153,N_1930);
nand U2563 (N_2563,N_1969,N_1532);
or U2564 (N_2564,N_1141,N_1005);
or U2565 (N_2565,N_1613,N_1669);
and U2566 (N_2566,N_1382,N_1198);
nand U2567 (N_2567,N_1902,N_1818);
nor U2568 (N_2568,N_1516,N_1269);
or U2569 (N_2569,N_1178,N_1765);
or U2570 (N_2570,N_1039,N_1404);
nor U2571 (N_2571,N_1985,N_1365);
nor U2572 (N_2572,N_1475,N_1773);
nand U2573 (N_2573,N_1536,N_1761);
nor U2574 (N_2574,N_1551,N_1350);
nand U2575 (N_2575,N_1144,N_1111);
nor U2576 (N_2576,N_1818,N_1448);
and U2577 (N_2577,N_1969,N_1514);
nor U2578 (N_2578,N_1590,N_1533);
nor U2579 (N_2579,N_1977,N_1124);
nand U2580 (N_2580,N_1493,N_1967);
nand U2581 (N_2581,N_1755,N_1514);
or U2582 (N_2582,N_1083,N_1654);
or U2583 (N_2583,N_1084,N_1521);
nand U2584 (N_2584,N_1745,N_1143);
and U2585 (N_2585,N_1093,N_1819);
or U2586 (N_2586,N_1398,N_1544);
nor U2587 (N_2587,N_1295,N_1818);
and U2588 (N_2588,N_1574,N_1906);
and U2589 (N_2589,N_1619,N_1591);
nor U2590 (N_2590,N_1065,N_1339);
and U2591 (N_2591,N_1706,N_1065);
and U2592 (N_2592,N_1499,N_1966);
or U2593 (N_2593,N_1829,N_1376);
and U2594 (N_2594,N_1006,N_1863);
and U2595 (N_2595,N_1247,N_1901);
nand U2596 (N_2596,N_1743,N_1315);
nand U2597 (N_2597,N_1427,N_1701);
nor U2598 (N_2598,N_1003,N_1750);
or U2599 (N_2599,N_1338,N_1767);
and U2600 (N_2600,N_1823,N_1028);
or U2601 (N_2601,N_1058,N_1751);
nand U2602 (N_2602,N_1232,N_1569);
and U2603 (N_2603,N_1583,N_1786);
nand U2604 (N_2604,N_1248,N_1626);
nand U2605 (N_2605,N_1900,N_1538);
and U2606 (N_2606,N_1204,N_1405);
or U2607 (N_2607,N_1522,N_1398);
nand U2608 (N_2608,N_1940,N_1368);
nand U2609 (N_2609,N_1653,N_1832);
xor U2610 (N_2610,N_1843,N_1019);
nand U2611 (N_2611,N_1661,N_1437);
nand U2612 (N_2612,N_1704,N_1796);
nor U2613 (N_2613,N_1118,N_1340);
and U2614 (N_2614,N_1290,N_1574);
and U2615 (N_2615,N_1374,N_1252);
nand U2616 (N_2616,N_1282,N_1602);
nand U2617 (N_2617,N_1808,N_1612);
and U2618 (N_2618,N_1025,N_1844);
or U2619 (N_2619,N_1423,N_1495);
nand U2620 (N_2620,N_1251,N_1855);
or U2621 (N_2621,N_1387,N_1187);
nor U2622 (N_2622,N_1438,N_1944);
and U2623 (N_2623,N_1485,N_1975);
or U2624 (N_2624,N_1231,N_1043);
nand U2625 (N_2625,N_1658,N_1755);
or U2626 (N_2626,N_1578,N_1848);
xnor U2627 (N_2627,N_1491,N_1256);
nor U2628 (N_2628,N_1291,N_1641);
nand U2629 (N_2629,N_1938,N_1158);
nor U2630 (N_2630,N_1026,N_1758);
or U2631 (N_2631,N_1626,N_1950);
nand U2632 (N_2632,N_1712,N_1484);
nor U2633 (N_2633,N_1393,N_1850);
or U2634 (N_2634,N_1408,N_1537);
nand U2635 (N_2635,N_1976,N_1158);
nand U2636 (N_2636,N_1167,N_1473);
and U2637 (N_2637,N_1483,N_1905);
or U2638 (N_2638,N_1176,N_1195);
nand U2639 (N_2639,N_1781,N_1519);
and U2640 (N_2640,N_1747,N_1328);
or U2641 (N_2641,N_1008,N_1554);
nor U2642 (N_2642,N_1878,N_1267);
and U2643 (N_2643,N_1400,N_1481);
nand U2644 (N_2644,N_1080,N_1173);
nor U2645 (N_2645,N_1832,N_1893);
nor U2646 (N_2646,N_1116,N_1243);
nor U2647 (N_2647,N_1667,N_1691);
nand U2648 (N_2648,N_1950,N_1103);
and U2649 (N_2649,N_1547,N_1753);
and U2650 (N_2650,N_1839,N_1769);
nand U2651 (N_2651,N_1236,N_1230);
nand U2652 (N_2652,N_1962,N_1115);
nand U2653 (N_2653,N_1735,N_1240);
or U2654 (N_2654,N_1634,N_1051);
nor U2655 (N_2655,N_1424,N_1695);
and U2656 (N_2656,N_1090,N_1807);
nor U2657 (N_2657,N_1846,N_1563);
or U2658 (N_2658,N_1328,N_1619);
xnor U2659 (N_2659,N_1435,N_1970);
nand U2660 (N_2660,N_1156,N_1992);
or U2661 (N_2661,N_1193,N_1684);
or U2662 (N_2662,N_1667,N_1255);
and U2663 (N_2663,N_1356,N_1897);
and U2664 (N_2664,N_1179,N_1736);
or U2665 (N_2665,N_1264,N_1101);
nor U2666 (N_2666,N_1917,N_1984);
nand U2667 (N_2667,N_1033,N_1168);
or U2668 (N_2668,N_1766,N_1400);
or U2669 (N_2669,N_1437,N_1962);
nand U2670 (N_2670,N_1175,N_1811);
or U2671 (N_2671,N_1767,N_1975);
or U2672 (N_2672,N_1363,N_1737);
and U2673 (N_2673,N_1109,N_1523);
nor U2674 (N_2674,N_1933,N_1501);
or U2675 (N_2675,N_1020,N_1321);
or U2676 (N_2676,N_1996,N_1821);
and U2677 (N_2677,N_1653,N_1563);
and U2678 (N_2678,N_1373,N_1371);
nand U2679 (N_2679,N_1340,N_1961);
and U2680 (N_2680,N_1418,N_1018);
nand U2681 (N_2681,N_1878,N_1167);
or U2682 (N_2682,N_1655,N_1850);
nor U2683 (N_2683,N_1313,N_1943);
or U2684 (N_2684,N_1303,N_1746);
nor U2685 (N_2685,N_1194,N_1879);
and U2686 (N_2686,N_1676,N_1738);
nand U2687 (N_2687,N_1256,N_1735);
nand U2688 (N_2688,N_1356,N_1095);
and U2689 (N_2689,N_1307,N_1709);
nand U2690 (N_2690,N_1750,N_1690);
nand U2691 (N_2691,N_1708,N_1142);
or U2692 (N_2692,N_1623,N_1591);
nor U2693 (N_2693,N_1974,N_1730);
or U2694 (N_2694,N_1263,N_1014);
or U2695 (N_2695,N_1050,N_1945);
or U2696 (N_2696,N_1725,N_1177);
nor U2697 (N_2697,N_1368,N_1435);
nand U2698 (N_2698,N_1077,N_1534);
or U2699 (N_2699,N_1915,N_1730);
nor U2700 (N_2700,N_1616,N_1703);
and U2701 (N_2701,N_1472,N_1755);
nor U2702 (N_2702,N_1897,N_1643);
or U2703 (N_2703,N_1784,N_1155);
nand U2704 (N_2704,N_1950,N_1989);
or U2705 (N_2705,N_1920,N_1269);
and U2706 (N_2706,N_1550,N_1396);
or U2707 (N_2707,N_1314,N_1074);
and U2708 (N_2708,N_1032,N_1362);
nor U2709 (N_2709,N_1949,N_1291);
nand U2710 (N_2710,N_1424,N_1438);
nand U2711 (N_2711,N_1797,N_1337);
or U2712 (N_2712,N_1773,N_1784);
nor U2713 (N_2713,N_1672,N_1524);
and U2714 (N_2714,N_1598,N_1981);
nand U2715 (N_2715,N_1731,N_1071);
and U2716 (N_2716,N_1649,N_1038);
nand U2717 (N_2717,N_1108,N_1876);
or U2718 (N_2718,N_1946,N_1059);
and U2719 (N_2719,N_1947,N_1615);
and U2720 (N_2720,N_1626,N_1418);
nand U2721 (N_2721,N_1176,N_1641);
nor U2722 (N_2722,N_1730,N_1705);
nand U2723 (N_2723,N_1008,N_1686);
or U2724 (N_2724,N_1376,N_1361);
nor U2725 (N_2725,N_1429,N_1800);
and U2726 (N_2726,N_1400,N_1353);
nand U2727 (N_2727,N_1289,N_1038);
nor U2728 (N_2728,N_1551,N_1459);
nor U2729 (N_2729,N_1756,N_1772);
or U2730 (N_2730,N_1812,N_1851);
nand U2731 (N_2731,N_1491,N_1524);
xor U2732 (N_2732,N_1004,N_1963);
nand U2733 (N_2733,N_1977,N_1961);
nand U2734 (N_2734,N_1630,N_1105);
or U2735 (N_2735,N_1074,N_1570);
and U2736 (N_2736,N_1601,N_1127);
nand U2737 (N_2737,N_1808,N_1283);
and U2738 (N_2738,N_1758,N_1042);
nor U2739 (N_2739,N_1248,N_1386);
nand U2740 (N_2740,N_1004,N_1037);
and U2741 (N_2741,N_1205,N_1670);
nor U2742 (N_2742,N_1183,N_1102);
nor U2743 (N_2743,N_1340,N_1788);
nor U2744 (N_2744,N_1557,N_1550);
or U2745 (N_2745,N_1769,N_1170);
or U2746 (N_2746,N_1369,N_1524);
or U2747 (N_2747,N_1328,N_1817);
and U2748 (N_2748,N_1456,N_1977);
nand U2749 (N_2749,N_1401,N_1562);
nand U2750 (N_2750,N_1313,N_1650);
or U2751 (N_2751,N_1804,N_1930);
or U2752 (N_2752,N_1035,N_1637);
nor U2753 (N_2753,N_1247,N_1565);
and U2754 (N_2754,N_1024,N_1003);
and U2755 (N_2755,N_1260,N_1228);
nand U2756 (N_2756,N_1488,N_1640);
nand U2757 (N_2757,N_1761,N_1393);
or U2758 (N_2758,N_1718,N_1358);
or U2759 (N_2759,N_1236,N_1874);
nor U2760 (N_2760,N_1105,N_1076);
or U2761 (N_2761,N_1624,N_1428);
nor U2762 (N_2762,N_1148,N_1667);
nand U2763 (N_2763,N_1078,N_1354);
or U2764 (N_2764,N_1143,N_1609);
or U2765 (N_2765,N_1050,N_1200);
nor U2766 (N_2766,N_1810,N_1666);
or U2767 (N_2767,N_1808,N_1199);
nor U2768 (N_2768,N_1411,N_1221);
or U2769 (N_2769,N_1337,N_1710);
nand U2770 (N_2770,N_1382,N_1754);
and U2771 (N_2771,N_1543,N_1454);
or U2772 (N_2772,N_1689,N_1612);
nor U2773 (N_2773,N_1261,N_1784);
and U2774 (N_2774,N_1209,N_1226);
nand U2775 (N_2775,N_1654,N_1497);
xor U2776 (N_2776,N_1414,N_1793);
nand U2777 (N_2777,N_1209,N_1043);
nor U2778 (N_2778,N_1129,N_1436);
nor U2779 (N_2779,N_1890,N_1045);
nand U2780 (N_2780,N_1348,N_1208);
nor U2781 (N_2781,N_1869,N_1410);
nand U2782 (N_2782,N_1180,N_1557);
nor U2783 (N_2783,N_1595,N_1661);
or U2784 (N_2784,N_1997,N_1363);
nand U2785 (N_2785,N_1270,N_1697);
nand U2786 (N_2786,N_1337,N_1690);
nand U2787 (N_2787,N_1132,N_1225);
nor U2788 (N_2788,N_1107,N_1047);
nor U2789 (N_2789,N_1918,N_1373);
nor U2790 (N_2790,N_1301,N_1294);
or U2791 (N_2791,N_1919,N_1881);
or U2792 (N_2792,N_1353,N_1950);
and U2793 (N_2793,N_1084,N_1189);
or U2794 (N_2794,N_1168,N_1486);
and U2795 (N_2795,N_1871,N_1715);
nor U2796 (N_2796,N_1561,N_1357);
nand U2797 (N_2797,N_1502,N_1770);
nor U2798 (N_2798,N_1613,N_1106);
nor U2799 (N_2799,N_1742,N_1049);
nor U2800 (N_2800,N_1201,N_1185);
nand U2801 (N_2801,N_1120,N_1580);
nand U2802 (N_2802,N_1922,N_1427);
nand U2803 (N_2803,N_1008,N_1155);
nor U2804 (N_2804,N_1190,N_1692);
nor U2805 (N_2805,N_1823,N_1363);
or U2806 (N_2806,N_1214,N_1877);
or U2807 (N_2807,N_1733,N_1619);
or U2808 (N_2808,N_1717,N_1919);
nor U2809 (N_2809,N_1974,N_1995);
and U2810 (N_2810,N_1686,N_1376);
and U2811 (N_2811,N_1650,N_1367);
nor U2812 (N_2812,N_1035,N_1346);
and U2813 (N_2813,N_1332,N_1656);
and U2814 (N_2814,N_1952,N_1027);
and U2815 (N_2815,N_1370,N_1089);
nor U2816 (N_2816,N_1399,N_1996);
and U2817 (N_2817,N_1738,N_1300);
nor U2818 (N_2818,N_1064,N_1519);
nand U2819 (N_2819,N_1500,N_1372);
nor U2820 (N_2820,N_1943,N_1207);
or U2821 (N_2821,N_1478,N_1151);
nand U2822 (N_2822,N_1281,N_1975);
and U2823 (N_2823,N_1228,N_1470);
and U2824 (N_2824,N_1749,N_1853);
or U2825 (N_2825,N_1373,N_1233);
and U2826 (N_2826,N_1035,N_1934);
nor U2827 (N_2827,N_1043,N_1947);
nor U2828 (N_2828,N_1731,N_1130);
nor U2829 (N_2829,N_1393,N_1561);
nor U2830 (N_2830,N_1668,N_1722);
nor U2831 (N_2831,N_1979,N_1644);
or U2832 (N_2832,N_1788,N_1592);
nor U2833 (N_2833,N_1958,N_1414);
or U2834 (N_2834,N_1852,N_1052);
or U2835 (N_2835,N_1906,N_1076);
nor U2836 (N_2836,N_1305,N_1222);
nand U2837 (N_2837,N_1618,N_1380);
or U2838 (N_2838,N_1615,N_1354);
and U2839 (N_2839,N_1192,N_1247);
xnor U2840 (N_2840,N_1925,N_1397);
nand U2841 (N_2841,N_1521,N_1748);
and U2842 (N_2842,N_1087,N_1140);
and U2843 (N_2843,N_1977,N_1610);
nand U2844 (N_2844,N_1575,N_1201);
nand U2845 (N_2845,N_1288,N_1930);
nand U2846 (N_2846,N_1410,N_1669);
or U2847 (N_2847,N_1339,N_1058);
nand U2848 (N_2848,N_1229,N_1950);
and U2849 (N_2849,N_1570,N_1967);
and U2850 (N_2850,N_1131,N_1705);
and U2851 (N_2851,N_1459,N_1838);
or U2852 (N_2852,N_1889,N_1971);
nor U2853 (N_2853,N_1249,N_1466);
nor U2854 (N_2854,N_1498,N_1287);
and U2855 (N_2855,N_1231,N_1447);
or U2856 (N_2856,N_1715,N_1373);
or U2857 (N_2857,N_1441,N_1094);
and U2858 (N_2858,N_1497,N_1317);
or U2859 (N_2859,N_1959,N_1871);
nor U2860 (N_2860,N_1952,N_1442);
or U2861 (N_2861,N_1472,N_1241);
or U2862 (N_2862,N_1894,N_1243);
or U2863 (N_2863,N_1559,N_1205);
and U2864 (N_2864,N_1748,N_1165);
and U2865 (N_2865,N_1181,N_1689);
and U2866 (N_2866,N_1106,N_1758);
and U2867 (N_2867,N_1899,N_1020);
and U2868 (N_2868,N_1508,N_1355);
or U2869 (N_2869,N_1043,N_1201);
nand U2870 (N_2870,N_1886,N_1365);
and U2871 (N_2871,N_1915,N_1430);
and U2872 (N_2872,N_1988,N_1969);
and U2873 (N_2873,N_1996,N_1170);
nor U2874 (N_2874,N_1332,N_1037);
and U2875 (N_2875,N_1889,N_1822);
and U2876 (N_2876,N_1136,N_1564);
nand U2877 (N_2877,N_1150,N_1298);
and U2878 (N_2878,N_1030,N_1032);
or U2879 (N_2879,N_1297,N_1014);
or U2880 (N_2880,N_1774,N_1476);
and U2881 (N_2881,N_1466,N_1782);
or U2882 (N_2882,N_1551,N_1174);
xnor U2883 (N_2883,N_1410,N_1800);
nor U2884 (N_2884,N_1900,N_1029);
or U2885 (N_2885,N_1623,N_1182);
nor U2886 (N_2886,N_1779,N_1965);
and U2887 (N_2887,N_1277,N_1121);
nor U2888 (N_2888,N_1855,N_1319);
nor U2889 (N_2889,N_1823,N_1182);
nor U2890 (N_2890,N_1200,N_1432);
and U2891 (N_2891,N_1374,N_1071);
nand U2892 (N_2892,N_1876,N_1526);
nor U2893 (N_2893,N_1641,N_1162);
nor U2894 (N_2894,N_1760,N_1173);
nor U2895 (N_2895,N_1606,N_1641);
nor U2896 (N_2896,N_1386,N_1157);
and U2897 (N_2897,N_1646,N_1077);
and U2898 (N_2898,N_1742,N_1890);
and U2899 (N_2899,N_1958,N_1041);
and U2900 (N_2900,N_1722,N_1450);
nand U2901 (N_2901,N_1691,N_1525);
nor U2902 (N_2902,N_1151,N_1201);
and U2903 (N_2903,N_1729,N_1986);
nand U2904 (N_2904,N_1262,N_1817);
nand U2905 (N_2905,N_1169,N_1322);
and U2906 (N_2906,N_1741,N_1498);
or U2907 (N_2907,N_1493,N_1531);
nor U2908 (N_2908,N_1747,N_1082);
nor U2909 (N_2909,N_1094,N_1498);
or U2910 (N_2910,N_1609,N_1190);
or U2911 (N_2911,N_1793,N_1825);
nor U2912 (N_2912,N_1090,N_1244);
and U2913 (N_2913,N_1706,N_1346);
or U2914 (N_2914,N_1499,N_1063);
and U2915 (N_2915,N_1258,N_1744);
nand U2916 (N_2916,N_1840,N_1165);
nand U2917 (N_2917,N_1532,N_1306);
nor U2918 (N_2918,N_1900,N_1385);
and U2919 (N_2919,N_1662,N_1705);
or U2920 (N_2920,N_1806,N_1146);
and U2921 (N_2921,N_1274,N_1548);
or U2922 (N_2922,N_1224,N_1561);
and U2923 (N_2923,N_1327,N_1222);
nor U2924 (N_2924,N_1639,N_1494);
nor U2925 (N_2925,N_1412,N_1133);
xnor U2926 (N_2926,N_1981,N_1883);
nand U2927 (N_2927,N_1052,N_1580);
nor U2928 (N_2928,N_1679,N_1200);
nand U2929 (N_2929,N_1127,N_1768);
nand U2930 (N_2930,N_1607,N_1771);
nand U2931 (N_2931,N_1473,N_1870);
and U2932 (N_2932,N_1918,N_1048);
nand U2933 (N_2933,N_1284,N_1464);
or U2934 (N_2934,N_1631,N_1630);
xnor U2935 (N_2935,N_1379,N_1779);
nor U2936 (N_2936,N_1689,N_1338);
nand U2937 (N_2937,N_1414,N_1734);
nor U2938 (N_2938,N_1022,N_1883);
nor U2939 (N_2939,N_1829,N_1226);
and U2940 (N_2940,N_1947,N_1579);
or U2941 (N_2941,N_1203,N_1190);
or U2942 (N_2942,N_1957,N_1500);
nand U2943 (N_2943,N_1355,N_1291);
and U2944 (N_2944,N_1345,N_1865);
and U2945 (N_2945,N_1401,N_1972);
or U2946 (N_2946,N_1052,N_1073);
or U2947 (N_2947,N_1997,N_1158);
nand U2948 (N_2948,N_1385,N_1272);
and U2949 (N_2949,N_1351,N_1051);
and U2950 (N_2950,N_1072,N_1661);
and U2951 (N_2951,N_1990,N_1095);
nand U2952 (N_2952,N_1678,N_1902);
nor U2953 (N_2953,N_1783,N_1735);
and U2954 (N_2954,N_1368,N_1055);
nand U2955 (N_2955,N_1093,N_1529);
nand U2956 (N_2956,N_1225,N_1474);
and U2957 (N_2957,N_1415,N_1025);
nand U2958 (N_2958,N_1820,N_1388);
and U2959 (N_2959,N_1614,N_1178);
nand U2960 (N_2960,N_1466,N_1606);
nor U2961 (N_2961,N_1604,N_1806);
nand U2962 (N_2962,N_1989,N_1110);
nor U2963 (N_2963,N_1721,N_1386);
nor U2964 (N_2964,N_1222,N_1799);
and U2965 (N_2965,N_1793,N_1480);
and U2966 (N_2966,N_1767,N_1780);
nand U2967 (N_2967,N_1410,N_1321);
or U2968 (N_2968,N_1868,N_1161);
or U2969 (N_2969,N_1613,N_1378);
and U2970 (N_2970,N_1141,N_1636);
nand U2971 (N_2971,N_1541,N_1815);
nand U2972 (N_2972,N_1431,N_1993);
nor U2973 (N_2973,N_1285,N_1353);
and U2974 (N_2974,N_1769,N_1066);
or U2975 (N_2975,N_1413,N_1223);
nand U2976 (N_2976,N_1784,N_1292);
nor U2977 (N_2977,N_1027,N_1526);
nand U2978 (N_2978,N_1577,N_1839);
and U2979 (N_2979,N_1301,N_1026);
and U2980 (N_2980,N_1460,N_1889);
and U2981 (N_2981,N_1847,N_1957);
nor U2982 (N_2982,N_1560,N_1780);
or U2983 (N_2983,N_1451,N_1025);
nand U2984 (N_2984,N_1103,N_1412);
nand U2985 (N_2985,N_1327,N_1690);
nand U2986 (N_2986,N_1523,N_1976);
and U2987 (N_2987,N_1138,N_1816);
or U2988 (N_2988,N_1500,N_1574);
or U2989 (N_2989,N_1054,N_1298);
or U2990 (N_2990,N_1270,N_1559);
and U2991 (N_2991,N_1416,N_1354);
and U2992 (N_2992,N_1917,N_1563);
nand U2993 (N_2993,N_1043,N_1926);
and U2994 (N_2994,N_1523,N_1376);
or U2995 (N_2995,N_1204,N_1238);
or U2996 (N_2996,N_1197,N_1288);
and U2997 (N_2997,N_1087,N_1223);
and U2998 (N_2998,N_1679,N_1124);
or U2999 (N_2999,N_1174,N_1418);
nand U3000 (N_3000,N_2752,N_2334);
nor U3001 (N_3001,N_2384,N_2834);
and U3002 (N_3002,N_2741,N_2558);
or U3003 (N_3003,N_2579,N_2943);
nor U3004 (N_3004,N_2540,N_2407);
or U3005 (N_3005,N_2264,N_2439);
nor U3006 (N_3006,N_2648,N_2401);
or U3007 (N_3007,N_2268,N_2779);
nand U3008 (N_3008,N_2363,N_2232);
nor U3009 (N_3009,N_2772,N_2761);
nor U3010 (N_3010,N_2388,N_2866);
or U3011 (N_3011,N_2470,N_2117);
or U3012 (N_3012,N_2021,N_2510);
or U3013 (N_3013,N_2272,N_2915);
nand U3014 (N_3014,N_2602,N_2437);
nor U3015 (N_3015,N_2152,N_2405);
and U3016 (N_3016,N_2408,N_2968);
and U3017 (N_3017,N_2603,N_2592);
or U3018 (N_3018,N_2684,N_2469);
nor U3019 (N_3019,N_2835,N_2840);
or U3020 (N_3020,N_2795,N_2420);
and U3021 (N_3021,N_2061,N_2243);
nor U3022 (N_3022,N_2577,N_2262);
or U3023 (N_3023,N_2294,N_2621);
nand U3024 (N_3024,N_2079,N_2986);
and U3025 (N_3025,N_2385,N_2862);
nor U3026 (N_3026,N_2998,N_2837);
and U3027 (N_3027,N_2547,N_2685);
nand U3028 (N_3028,N_2398,N_2534);
and U3029 (N_3029,N_2906,N_2351);
nand U3030 (N_3030,N_2654,N_2151);
and U3031 (N_3031,N_2967,N_2652);
nand U3032 (N_3032,N_2074,N_2567);
nand U3033 (N_3033,N_2644,N_2389);
or U3034 (N_3034,N_2184,N_2280);
and U3035 (N_3035,N_2699,N_2759);
and U3036 (N_3036,N_2970,N_2670);
and U3037 (N_3037,N_2748,N_2872);
and U3038 (N_3038,N_2609,N_2478);
or U3039 (N_3039,N_2108,N_2030);
or U3040 (N_3040,N_2919,N_2853);
nor U3041 (N_3041,N_2423,N_2500);
nor U3042 (N_3042,N_2690,N_2817);
nor U3043 (N_3043,N_2126,N_2382);
or U3044 (N_3044,N_2963,N_2371);
nor U3045 (N_3045,N_2991,N_2627);
nand U3046 (N_3046,N_2634,N_2890);
and U3047 (N_3047,N_2367,N_2839);
nand U3048 (N_3048,N_2629,N_2873);
and U3049 (N_3049,N_2448,N_2164);
nor U3050 (N_3050,N_2016,N_2357);
nand U3051 (N_3051,N_2181,N_2324);
and U3052 (N_3052,N_2196,N_2551);
and U3053 (N_3053,N_2910,N_2810);
and U3054 (N_3054,N_2929,N_2374);
or U3055 (N_3055,N_2664,N_2391);
nor U3056 (N_3056,N_2908,N_2696);
or U3057 (N_3057,N_2564,N_2452);
nor U3058 (N_3058,N_2335,N_2987);
nor U3059 (N_3059,N_2446,N_2559);
or U3060 (N_3060,N_2372,N_2697);
nand U3061 (N_3061,N_2803,N_2005);
and U3062 (N_3062,N_2179,N_2733);
nand U3063 (N_3063,N_2430,N_2312);
and U3064 (N_3064,N_2956,N_2059);
and U3065 (N_3065,N_2740,N_2786);
nor U3066 (N_3066,N_2975,N_2868);
xnor U3067 (N_3067,N_2698,N_2843);
nand U3068 (N_3068,N_2680,N_2502);
or U3069 (N_3069,N_2332,N_2516);
and U3070 (N_3070,N_2345,N_2091);
or U3071 (N_3071,N_2322,N_2583);
xor U3072 (N_3072,N_2090,N_2932);
and U3073 (N_3073,N_2897,N_2617);
nor U3074 (N_3074,N_2316,N_2895);
xnor U3075 (N_3075,N_2594,N_2934);
nor U3076 (N_3076,N_2051,N_2971);
nand U3077 (N_3077,N_2749,N_2404);
nor U3078 (N_3078,N_2637,N_2154);
nand U3079 (N_3079,N_2505,N_2015);
nor U3080 (N_3080,N_2158,N_2467);
nor U3081 (N_3081,N_2459,N_2283);
nor U3082 (N_3082,N_2033,N_2160);
or U3083 (N_3083,N_2801,N_2736);
or U3084 (N_3084,N_2330,N_2891);
nor U3085 (N_3085,N_2624,N_2918);
or U3086 (N_3086,N_2520,N_2366);
nor U3087 (N_3087,N_2096,N_2974);
or U3088 (N_3088,N_2847,N_2568);
nor U3089 (N_3089,N_2443,N_2493);
nand U3090 (N_3090,N_2732,N_2017);
nor U3091 (N_3091,N_2599,N_2124);
nand U3092 (N_3092,N_2498,N_2923);
nand U3093 (N_3093,N_2327,N_2978);
nor U3094 (N_3094,N_2197,N_2219);
and U3095 (N_3095,N_2421,N_2047);
nand U3096 (N_3096,N_2576,N_2192);
nand U3097 (N_3097,N_2212,N_2658);
nor U3098 (N_3098,N_2622,N_2605);
xnor U3099 (N_3099,N_2585,N_2319);
and U3100 (N_3100,N_2566,N_2859);
nand U3101 (N_3101,N_2722,N_2643);
nor U3102 (N_3102,N_2589,N_2782);
nand U3103 (N_3103,N_2341,N_2720);
and U3104 (N_3104,N_2905,N_2705);
nand U3105 (N_3105,N_2311,N_2836);
or U3106 (N_3106,N_2453,N_2745);
nor U3107 (N_3107,N_2318,N_2953);
or U3108 (N_3108,N_2216,N_2930);
and U3109 (N_3109,N_2365,N_2601);
and U3110 (N_3110,N_2813,N_2024);
nor U3111 (N_3111,N_2776,N_2396);
or U3112 (N_3112,N_2375,N_2727);
or U3113 (N_3113,N_2076,N_2921);
nor U3114 (N_3114,N_2048,N_2191);
or U3115 (N_3115,N_2689,N_2506);
or U3116 (N_3116,N_2440,N_2981);
nand U3117 (N_3117,N_2220,N_2710);
nor U3118 (N_3118,N_2307,N_2753);
or U3119 (N_3119,N_2422,N_2744);
nand U3120 (N_3120,N_2792,N_2802);
or U3121 (N_3121,N_2807,N_2392);
or U3122 (N_3122,N_2266,N_2008);
and U3123 (N_3123,N_2263,N_2018);
or U3124 (N_3124,N_2153,N_2823);
nor U3125 (N_3125,N_2468,N_2914);
or U3126 (N_3126,N_2509,N_2434);
nand U3127 (N_3127,N_2298,N_2961);
nor U3128 (N_3128,N_2785,N_2623);
and U3129 (N_3129,N_2309,N_2042);
nand U3130 (N_3130,N_2373,N_2193);
nand U3131 (N_3131,N_2412,N_2189);
or U3132 (N_3132,N_2185,N_2530);
nand U3133 (N_3133,N_2994,N_2147);
and U3134 (N_3134,N_2766,N_2588);
nand U3135 (N_3135,N_2271,N_2166);
nor U3136 (N_3136,N_2286,N_2116);
nand U3137 (N_3137,N_2217,N_2764);
and U3138 (N_3138,N_2234,N_2701);
nand U3139 (N_3139,N_2569,N_2023);
and U3140 (N_3140,N_2708,N_2763);
nor U3141 (N_3141,N_2672,N_2436);
nor U3142 (N_3142,N_2820,N_2040);
nor U3143 (N_3143,N_2927,N_2134);
nor U3144 (N_3144,N_2833,N_2240);
or U3145 (N_3145,N_2521,N_2931);
nand U3146 (N_3146,N_2874,N_2797);
nand U3147 (N_3147,N_2094,N_2209);
and U3148 (N_3148,N_2425,N_2593);
nand U3149 (N_3149,N_2328,N_2228);
nand U3150 (N_3150,N_2128,N_2711);
and U3151 (N_3151,N_2080,N_2635);
or U3152 (N_3152,N_2514,N_2747);
nor U3153 (N_3153,N_2288,N_2660);
and U3154 (N_3154,N_2380,N_2246);
nor U3155 (N_3155,N_2778,N_2253);
nor U3156 (N_3156,N_2653,N_2402);
nand U3157 (N_3157,N_2242,N_2084);
nand U3158 (N_3158,N_2053,N_2554);
nor U3159 (N_3159,N_2983,N_2118);
or U3160 (N_3160,N_2360,N_2565);
nand U3161 (N_3161,N_2111,N_2317);
nand U3162 (N_3162,N_2162,N_2461);
and U3163 (N_3163,N_2177,N_2175);
or U3164 (N_3164,N_2916,N_2642);
and U3165 (N_3165,N_2533,N_2171);
nand U3166 (N_3166,N_2636,N_2002);
nand U3167 (N_3167,N_2362,N_2662);
or U3168 (N_3168,N_2085,N_2581);
and U3169 (N_3169,N_2526,N_2876);
or U3170 (N_3170,N_2631,N_2945);
and U3171 (N_3171,N_2950,N_2052);
or U3172 (N_3172,N_2225,N_2344);
nand U3173 (N_3173,N_2898,N_2867);
and U3174 (N_3174,N_2768,N_2145);
or U3175 (N_3175,N_2007,N_2615);
xor U3176 (N_3176,N_2349,N_2414);
nor U3177 (N_3177,N_2523,N_2980);
nand U3178 (N_3178,N_2203,N_2716);
nor U3179 (N_3179,N_2438,N_2825);
and U3180 (N_3180,N_2009,N_2003);
nor U3181 (N_3181,N_2669,N_2731);
or U3182 (N_3182,N_2495,N_2512);
nand U3183 (N_3183,N_2917,N_2432);
nand U3184 (N_3184,N_2251,N_2904);
and U3185 (N_3185,N_2427,N_2992);
xor U3186 (N_3186,N_2046,N_2058);
and U3187 (N_3187,N_2681,N_2686);
xnor U3188 (N_3188,N_2954,N_2400);
and U3189 (N_3189,N_2186,N_2248);
and U3190 (N_3190,N_2651,N_2337);
or U3191 (N_3191,N_2471,N_2014);
xnor U3192 (N_3192,N_2688,N_2088);
nor U3193 (N_3193,N_2838,N_2522);
and U3194 (N_3194,N_2537,N_2034);
and U3195 (N_3195,N_2123,N_2714);
or U3196 (N_3196,N_2993,N_2394);
nand U3197 (N_3197,N_2227,N_2715);
or U3198 (N_3198,N_2896,N_2972);
and U3199 (N_3199,N_2352,N_2205);
or U3200 (N_3200,N_2036,N_2235);
or U3201 (N_3201,N_2739,N_2083);
or U3202 (N_3202,N_2561,N_2417);
and U3203 (N_3203,N_2730,N_2667);
nand U3204 (N_3204,N_2517,N_2806);
nor U3205 (N_3205,N_2831,N_2233);
or U3206 (N_3206,N_2463,N_2295);
nand U3207 (N_3207,N_2210,N_2411);
or U3208 (N_3208,N_2814,N_2762);
nor U3209 (N_3209,N_2290,N_2525);
nor U3210 (N_3210,N_2570,N_2297);
and U3211 (N_3211,N_2960,N_2458);
or U3212 (N_3212,N_2155,N_2499);
or U3213 (N_3213,N_2329,N_2137);
nor U3214 (N_3214,N_2850,N_2195);
nand U3215 (N_3215,N_2805,N_2238);
nand U3216 (N_3216,N_2004,N_2142);
nor U3217 (N_3217,N_2611,N_2383);
or U3218 (N_3218,N_2812,N_2072);
nor U3219 (N_3219,N_2449,N_2479);
or U3220 (N_3220,N_2139,N_2369);
and U3221 (N_3221,N_2695,N_2466);
and U3222 (N_3222,N_2557,N_2031);
or U3223 (N_3223,N_2755,N_2082);
and U3224 (N_3224,N_2893,N_2877);
nor U3225 (N_3225,N_2097,N_2223);
nor U3226 (N_3226,N_2856,N_2911);
and U3227 (N_3227,N_2338,N_2800);
nand U3228 (N_3228,N_2997,N_2996);
or U3229 (N_3229,N_2650,N_2846);
and U3230 (N_3230,N_2426,N_2144);
or U3231 (N_3231,N_2169,N_2190);
or U3232 (N_3232,N_2325,N_2633);
nand U3233 (N_3233,N_2789,N_2952);
nor U3234 (N_3234,N_2958,N_2719);
nand U3235 (N_3235,N_2482,N_2880);
nand U3236 (N_3236,N_2870,N_2492);
or U3237 (N_3237,N_2553,N_2531);
and U3238 (N_3238,N_2069,N_2536);
or U3239 (N_3239,N_2901,N_2683);
nand U3240 (N_3240,N_2279,N_2455);
and U3241 (N_3241,N_2161,N_2773);
nor U3242 (N_3242,N_2851,N_2550);
nor U3243 (N_3243,N_2377,N_2150);
nand U3244 (N_3244,N_2092,N_2995);
nand U3245 (N_3245,N_2584,N_2457);
nor U3246 (N_3246,N_2703,N_2379);
nand U3247 (N_3247,N_2855,N_2343);
and U3248 (N_3248,N_2590,N_2026);
nor U3249 (N_3249,N_2140,N_2114);
nor U3250 (N_3250,N_2415,N_2940);
nand U3251 (N_3251,N_2176,N_2157);
nor U3252 (N_3252,N_2045,N_2725);
or U3253 (N_3253,N_2019,N_2068);
or U3254 (N_3254,N_2255,N_2798);
and U3255 (N_3255,N_2949,N_2545);
and U3256 (N_3256,N_2666,N_2700);
nand U3257 (N_3257,N_2723,N_2707);
nand U3258 (N_3258,N_2572,N_2323);
nor U3259 (N_3259,N_2965,N_2256);
or U3260 (N_3260,N_2291,N_2252);
or U3261 (N_3261,N_2555,N_2065);
and U3262 (N_3262,N_2926,N_2767);
and U3263 (N_3263,N_2340,N_2848);
or U3264 (N_3264,N_2032,N_2883);
and U3265 (N_3265,N_2244,N_2784);
and U3266 (N_3266,N_2765,N_2081);
nor U3267 (N_3267,N_2267,N_2884);
nand U3268 (N_3268,N_2429,N_2717);
nand U3269 (N_3269,N_2416,N_2845);
nand U3270 (N_3270,N_2827,N_2156);
nand U3271 (N_3271,N_2909,N_2665);
nand U3272 (N_3272,N_2793,N_2000);
nand U3273 (N_3273,N_2390,N_2273);
and U3274 (N_3274,N_2882,N_2413);
nor U3275 (N_3275,N_2087,N_2277);
nor U3276 (N_3276,N_2507,N_2063);
nor U3277 (N_3277,N_2738,N_2957);
or U3278 (N_3278,N_2503,N_2649);
nor U3279 (N_3279,N_2481,N_2539);
nor U3280 (N_3280,N_2130,N_2326);
and U3281 (N_3281,N_2973,N_2287);
nand U3282 (N_3282,N_2102,N_2442);
or U3283 (N_3283,N_2889,N_2066);
or U3284 (N_3284,N_2726,N_2535);
nor U3285 (N_3285,N_2808,N_2788);
nor U3286 (N_3286,N_2308,N_2497);
and U3287 (N_3287,N_2001,N_2936);
and U3288 (N_3288,N_2702,N_2491);
nor U3289 (N_3289,N_2067,N_2475);
nor U3290 (N_3290,N_2485,N_2606);
and U3291 (N_3291,N_2979,N_2368);
nand U3292 (N_3292,N_2346,N_2777);
nor U3293 (N_3293,N_2488,N_2706);
and U3294 (N_3294,N_2025,N_2818);
or U3295 (N_3295,N_2760,N_2620);
nor U3296 (N_3296,N_2815,N_2071);
and U3297 (N_3297,N_2933,N_2358);
nand U3298 (N_3298,N_2946,N_2822);
nand U3299 (N_3299,N_2541,N_2924);
or U3300 (N_3300,N_2598,N_2410);
or U3301 (N_3301,N_2182,N_2419);
or U3302 (N_3302,N_2292,N_2278);
or U3303 (N_3303,N_2679,N_2245);
or U3304 (N_3304,N_2206,N_2180);
nand U3305 (N_3305,N_2928,N_2202);
nand U3306 (N_3306,N_2902,N_2573);
nand U3307 (N_3307,N_2194,N_2050);
nand U3308 (N_3308,N_2103,N_2799);
or U3309 (N_3309,N_2456,N_2676);
or U3310 (N_3310,N_2613,N_2241);
nand U3311 (N_3311,N_2628,N_2112);
or U3312 (N_3312,N_2821,N_2878);
and U3313 (N_3313,N_2213,N_2393);
nand U3314 (N_3314,N_2054,N_2148);
nor U3315 (N_3315,N_2941,N_2062);
nor U3316 (N_3316,N_2757,N_2043);
and U3317 (N_3317,N_2673,N_2113);
or U3318 (N_3318,N_2020,N_2885);
or U3319 (N_3319,N_2355,N_2208);
nor U3320 (N_3320,N_2424,N_2804);
or U3321 (N_3321,N_2824,N_2064);
nand U3322 (N_3322,N_2729,N_2661);
and U3323 (N_3323,N_2655,N_2480);
nand U3324 (N_3324,N_2378,N_2899);
or U3325 (N_3325,N_2811,N_2037);
and U3326 (N_3326,N_2574,N_2938);
nand U3327 (N_3327,N_2663,N_2659);
and U3328 (N_3328,N_2881,N_2274);
and U3329 (N_3329,N_2472,N_2886);
and U3330 (N_3330,N_2832,N_2314);
nor U3331 (N_3331,N_2445,N_2988);
nor U3332 (N_3332,N_2022,N_2301);
or U3333 (N_3333,N_2751,N_2675);
and U3334 (N_3334,N_2582,N_2006);
nor U3335 (N_3335,N_2168,N_2029);
or U3336 (N_3336,N_2863,N_2447);
nand U3337 (N_3337,N_2462,N_2041);
nand U3338 (N_3338,N_2104,N_2571);
and U3339 (N_3339,N_2922,N_2289);
and U3340 (N_3340,N_2913,N_2406);
or U3341 (N_3341,N_2721,N_2348);
and U3342 (N_3342,N_2907,N_2619);
nand U3343 (N_3343,N_2183,N_2854);
nand U3344 (N_3344,N_2562,N_2826);
nor U3345 (N_3345,N_2494,N_2787);
nor U3346 (N_3346,N_2524,N_2556);
nor U3347 (N_3347,N_2451,N_2258);
and U3348 (N_3348,N_2159,N_2333);
and U3349 (N_3349,N_2955,N_2671);
or U3350 (N_3350,N_2486,N_2830);
nand U3351 (N_3351,N_2433,N_2364);
nand U3352 (N_3352,N_2310,N_2563);
or U3353 (N_3353,N_2109,N_2450);
or U3354 (N_3354,N_2270,N_2129);
or U3355 (N_3355,N_2200,N_2039);
nor U3356 (N_3356,N_2120,N_2011);
nor U3357 (N_3357,N_2548,N_2070);
nor U3358 (N_3358,N_2305,N_2474);
or U3359 (N_3359,N_2496,N_2115);
nor U3360 (N_3360,N_2709,N_2887);
and U3361 (N_3361,N_2875,N_2399);
and U3362 (N_3362,N_2418,N_2100);
or U3363 (N_3363,N_2852,N_2912);
and U3364 (N_3364,N_2674,N_2790);
and U3365 (N_3365,N_2300,N_2131);
and U3366 (N_3366,N_2597,N_2187);
nor U3367 (N_3367,N_2057,N_2049);
nor U3368 (N_3368,N_2086,N_2580);
or U3369 (N_3369,N_2269,N_2939);
or U3370 (N_3370,N_2894,N_2527);
nor U3371 (N_3371,N_2038,N_2315);
and U3372 (N_3372,N_2101,N_2409);
nor U3373 (N_3373,N_2473,N_2694);
nor U3374 (N_3374,N_2078,N_2865);
nor U3375 (N_3375,N_2110,N_2724);
nand U3376 (N_3376,N_2376,N_2604);
nor U3377 (N_3377,N_2483,N_2060);
xor U3378 (N_3378,N_2098,N_2511);
nor U3379 (N_3379,N_2610,N_2712);
and U3380 (N_3380,N_2920,N_2682);
or U3381 (N_3381,N_2221,N_2302);
nor U3382 (N_3382,N_2395,N_2387);
nor U3383 (N_3383,N_2677,N_2095);
or U3384 (N_3384,N_2645,N_2758);
nor U3385 (N_3385,N_2935,N_2199);
or U3386 (N_3386,N_2073,N_2331);
or U3387 (N_3387,N_2359,N_2796);
nor U3388 (N_3388,N_2892,N_2861);
nor U3389 (N_3389,N_2578,N_2614);
or U3390 (N_3390,N_2947,N_2127);
nor U3391 (N_3391,N_2099,N_2948);
and U3392 (N_3392,N_2035,N_2214);
nand U3393 (N_3393,N_2816,N_2428);
nand U3394 (N_3394,N_2704,N_2728);
or U3395 (N_3395,N_2713,N_2828);
or U3396 (N_3396,N_2299,N_2632);
nand U3397 (N_3397,N_2769,N_2218);
nand U3398 (N_3398,N_2237,N_2444);
nand U3399 (N_3399,N_2303,N_2869);
or U3400 (N_3400,N_2211,N_2260);
nor U3401 (N_3401,N_2841,N_2771);
and U3402 (N_3402,N_2249,N_2276);
and U3403 (N_3403,N_2075,N_2575);
nand U3404 (N_3404,N_2012,N_2141);
or U3405 (N_3405,N_2844,N_2172);
and U3406 (N_3406,N_2028,N_2959);
nand U3407 (N_3407,N_2107,N_2135);
or U3408 (N_3408,N_2487,N_2925);
nor U3409 (N_3409,N_2431,N_2513);
or U3410 (N_3410,N_2657,N_2229);
or U3411 (N_3411,N_2361,N_2639);
and U3412 (N_3412,N_2693,N_2595);
and U3413 (N_3413,N_2586,N_2044);
nor U3414 (N_3414,N_2122,N_2989);
and U3415 (N_3415,N_2587,N_2275);
or U3416 (N_3416,N_2386,N_2608);
nand U3417 (N_3417,N_2809,N_2010);
and U3418 (N_3418,N_2860,N_2515);
or U3419 (N_3419,N_2600,N_2903);
and U3420 (N_3420,N_2842,N_2656);
or U3421 (N_3421,N_2165,N_2982);
nor U3422 (N_3422,N_2465,N_2607);
and U3423 (N_3423,N_2774,N_2692);
nor U3424 (N_3424,N_2770,N_2077);
and U3425 (N_3425,N_2976,N_2207);
and U3426 (N_3426,N_2125,N_2239);
and U3427 (N_3427,N_2163,N_2638);
or U3428 (N_3428,N_2261,N_2143);
and U3429 (N_3429,N_2178,N_2735);
nand U3430 (N_3430,N_2504,N_2625);
nand U3431 (N_3431,N_2791,N_2977);
nand U3432 (N_3432,N_2687,N_2612);
and U3433 (N_3433,N_2691,N_2170);
nor U3434 (N_3434,N_2321,N_2259);
or U3435 (N_3435,N_2236,N_2538);
nor U3436 (N_3436,N_2013,N_2951);
xor U3437 (N_3437,N_2354,N_2678);
nor U3438 (N_3438,N_2201,N_2089);
and U3439 (N_3439,N_2105,N_2544);
or U3440 (N_3440,N_2149,N_2350);
nor U3441 (N_3441,N_2641,N_2056);
or U3442 (N_3442,N_2306,N_2490);
and U3443 (N_3443,N_2027,N_2093);
and U3444 (N_3444,N_2508,N_2136);
or U3445 (N_3445,N_2226,N_2794);
and U3446 (N_3446,N_2281,N_2756);
nor U3447 (N_3447,N_2858,N_2985);
or U3448 (N_3448,N_2167,N_2626);
nand U3449 (N_3449,N_2138,N_2146);
nor U3450 (N_3450,N_2339,N_2984);
nand U3451 (N_3451,N_2055,N_2630);
nand U3452 (N_3452,N_2743,N_2937);
and U3453 (N_3453,N_2403,N_2640);
xnor U3454 (N_3454,N_2231,N_2737);
and U3455 (N_3455,N_2477,N_2964);
nor U3456 (N_3456,N_2254,N_2460);
and U3457 (N_3457,N_2247,N_2174);
and U3458 (N_3458,N_2618,N_2519);
and U3459 (N_3459,N_2222,N_2173);
nand U3460 (N_3460,N_2829,N_2293);
and U3461 (N_3461,N_2549,N_2888);
and U3462 (N_3462,N_2336,N_2864);
and U3463 (N_3463,N_2501,N_2198);
or U3464 (N_3464,N_2999,N_2518);
nand U3465 (N_3465,N_2119,N_2879);
nand U3466 (N_3466,N_2265,N_2990);
nand U3467 (N_3467,N_2370,N_2204);
and U3468 (N_3468,N_2282,N_2250);
nand U3469 (N_3469,N_2647,N_2132);
and U3470 (N_3470,N_2754,N_2529);
or U3471 (N_3471,N_2476,N_2532);
nor U3472 (N_3472,N_2121,N_2347);
nand U3473 (N_3473,N_2106,N_2969);
nand U3474 (N_3474,N_2435,N_2489);
nand U3475 (N_3475,N_2284,N_2304);
nor U3476 (N_3476,N_2783,N_2342);
nand U3477 (N_3477,N_2718,N_2746);
or U3478 (N_3478,N_2781,N_2775);
or U3479 (N_3479,N_2454,N_2871);
nor U3480 (N_3480,N_2962,N_2397);
nand U3481 (N_3481,N_2542,N_2484);
and U3482 (N_3482,N_2296,N_2552);
nand U3483 (N_3483,N_2734,N_2857);
nand U3484 (N_3484,N_2285,N_2849);
or U3485 (N_3485,N_2543,N_2616);
and U3486 (N_3486,N_2596,N_2819);
or U3487 (N_3487,N_2224,N_2900);
or U3488 (N_3488,N_2742,N_2966);
nor U3489 (N_3489,N_2546,N_2320);
nor U3490 (N_3490,N_2560,N_2528);
nand U3491 (N_3491,N_2591,N_2441);
nand U3492 (N_3492,N_2944,N_2313);
nor U3493 (N_3493,N_2464,N_2780);
nor U3494 (N_3494,N_2750,N_2133);
nand U3495 (N_3495,N_2257,N_2356);
or U3496 (N_3496,N_2942,N_2353);
nor U3497 (N_3497,N_2215,N_2188);
nor U3498 (N_3498,N_2646,N_2230);
nand U3499 (N_3499,N_2668,N_2381);
nand U3500 (N_3500,N_2094,N_2009);
or U3501 (N_3501,N_2469,N_2493);
and U3502 (N_3502,N_2562,N_2819);
and U3503 (N_3503,N_2298,N_2829);
or U3504 (N_3504,N_2160,N_2475);
and U3505 (N_3505,N_2098,N_2170);
nor U3506 (N_3506,N_2055,N_2348);
nand U3507 (N_3507,N_2293,N_2088);
nor U3508 (N_3508,N_2594,N_2229);
nor U3509 (N_3509,N_2816,N_2992);
nand U3510 (N_3510,N_2057,N_2941);
and U3511 (N_3511,N_2904,N_2053);
nor U3512 (N_3512,N_2504,N_2942);
or U3513 (N_3513,N_2092,N_2112);
and U3514 (N_3514,N_2343,N_2798);
or U3515 (N_3515,N_2431,N_2691);
nand U3516 (N_3516,N_2605,N_2959);
nor U3517 (N_3517,N_2242,N_2730);
nor U3518 (N_3518,N_2728,N_2769);
or U3519 (N_3519,N_2185,N_2885);
nand U3520 (N_3520,N_2081,N_2249);
and U3521 (N_3521,N_2903,N_2061);
nand U3522 (N_3522,N_2202,N_2609);
and U3523 (N_3523,N_2457,N_2997);
nor U3524 (N_3524,N_2973,N_2250);
and U3525 (N_3525,N_2831,N_2680);
nor U3526 (N_3526,N_2294,N_2747);
or U3527 (N_3527,N_2680,N_2736);
nand U3528 (N_3528,N_2785,N_2174);
and U3529 (N_3529,N_2176,N_2111);
or U3530 (N_3530,N_2375,N_2288);
nor U3531 (N_3531,N_2286,N_2250);
or U3532 (N_3532,N_2675,N_2154);
nand U3533 (N_3533,N_2360,N_2474);
and U3534 (N_3534,N_2954,N_2591);
and U3535 (N_3535,N_2423,N_2390);
nor U3536 (N_3536,N_2832,N_2345);
or U3537 (N_3537,N_2318,N_2264);
or U3538 (N_3538,N_2146,N_2166);
and U3539 (N_3539,N_2712,N_2458);
nor U3540 (N_3540,N_2537,N_2585);
and U3541 (N_3541,N_2962,N_2885);
nor U3542 (N_3542,N_2281,N_2381);
or U3543 (N_3543,N_2902,N_2596);
nor U3544 (N_3544,N_2659,N_2759);
nor U3545 (N_3545,N_2173,N_2158);
nand U3546 (N_3546,N_2529,N_2368);
or U3547 (N_3547,N_2191,N_2170);
nor U3548 (N_3548,N_2330,N_2055);
or U3549 (N_3549,N_2491,N_2900);
nor U3550 (N_3550,N_2851,N_2699);
nor U3551 (N_3551,N_2877,N_2517);
nand U3552 (N_3552,N_2309,N_2590);
or U3553 (N_3553,N_2579,N_2181);
nor U3554 (N_3554,N_2451,N_2618);
nor U3555 (N_3555,N_2365,N_2761);
nand U3556 (N_3556,N_2969,N_2198);
and U3557 (N_3557,N_2500,N_2492);
nor U3558 (N_3558,N_2068,N_2909);
and U3559 (N_3559,N_2582,N_2208);
or U3560 (N_3560,N_2425,N_2963);
nor U3561 (N_3561,N_2769,N_2829);
or U3562 (N_3562,N_2027,N_2573);
and U3563 (N_3563,N_2559,N_2963);
nand U3564 (N_3564,N_2699,N_2714);
nor U3565 (N_3565,N_2133,N_2499);
and U3566 (N_3566,N_2936,N_2792);
nand U3567 (N_3567,N_2672,N_2664);
and U3568 (N_3568,N_2340,N_2713);
or U3569 (N_3569,N_2749,N_2804);
or U3570 (N_3570,N_2992,N_2982);
nor U3571 (N_3571,N_2593,N_2323);
or U3572 (N_3572,N_2300,N_2788);
nor U3573 (N_3573,N_2160,N_2777);
and U3574 (N_3574,N_2199,N_2167);
or U3575 (N_3575,N_2017,N_2679);
and U3576 (N_3576,N_2960,N_2538);
and U3577 (N_3577,N_2372,N_2404);
nor U3578 (N_3578,N_2246,N_2360);
and U3579 (N_3579,N_2950,N_2217);
or U3580 (N_3580,N_2468,N_2353);
and U3581 (N_3581,N_2512,N_2255);
and U3582 (N_3582,N_2138,N_2745);
and U3583 (N_3583,N_2867,N_2128);
nor U3584 (N_3584,N_2984,N_2133);
nand U3585 (N_3585,N_2204,N_2899);
nor U3586 (N_3586,N_2422,N_2643);
or U3587 (N_3587,N_2117,N_2745);
nand U3588 (N_3588,N_2755,N_2257);
or U3589 (N_3589,N_2851,N_2522);
nand U3590 (N_3590,N_2895,N_2112);
or U3591 (N_3591,N_2210,N_2865);
nand U3592 (N_3592,N_2991,N_2604);
and U3593 (N_3593,N_2478,N_2751);
nor U3594 (N_3594,N_2694,N_2326);
and U3595 (N_3595,N_2832,N_2784);
and U3596 (N_3596,N_2019,N_2219);
nand U3597 (N_3597,N_2059,N_2150);
nor U3598 (N_3598,N_2398,N_2937);
nor U3599 (N_3599,N_2818,N_2241);
nor U3600 (N_3600,N_2382,N_2654);
nand U3601 (N_3601,N_2325,N_2409);
nor U3602 (N_3602,N_2425,N_2759);
nand U3603 (N_3603,N_2083,N_2716);
or U3604 (N_3604,N_2023,N_2196);
or U3605 (N_3605,N_2735,N_2240);
nor U3606 (N_3606,N_2777,N_2337);
nand U3607 (N_3607,N_2975,N_2745);
nor U3608 (N_3608,N_2864,N_2018);
or U3609 (N_3609,N_2275,N_2517);
nor U3610 (N_3610,N_2457,N_2213);
and U3611 (N_3611,N_2384,N_2652);
or U3612 (N_3612,N_2835,N_2551);
nand U3613 (N_3613,N_2211,N_2811);
and U3614 (N_3614,N_2161,N_2048);
nand U3615 (N_3615,N_2531,N_2626);
or U3616 (N_3616,N_2846,N_2698);
nor U3617 (N_3617,N_2501,N_2041);
nand U3618 (N_3618,N_2058,N_2070);
and U3619 (N_3619,N_2368,N_2019);
nand U3620 (N_3620,N_2624,N_2264);
nor U3621 (N_3621,N_2579,N_2268);
nor U3622 (N_3622,N_2542,N_2099);
nor U3623 (N_3623,N_2094,N_2853);
and U3624 (N_3624,N_2598,N_2379);
and U3625 (N_3625,N_2093,N_2576);
nor U3626 (N_3626,N_2364,N_2321);
nor U3627 (N_3627,N_2562,N_2322);
and U3628 (N_3628,N_2210,N_2584);
nand U3629 (N_3629,N_2436,N_2250);
and U3630 (N_3630,N_2762,N_2234);
nor U3631 (N_3631,N_2161,N_2836);
nor U3632 (N_3632,N_2805,N_2061);
and U3633 (N_3633,N_2621,N_2325);
or U3634 (N_3634,N_2144,N_2181);
nand U3635 (N_3635,N_2397,N_2944);
or U3636 (N_3636,N_2343,N_2683);
and U3637 (N_3637,N_2349,N_2710);
and U3638 (N_3638,N_2907,N_2797);
nor U3639 (N_3639,N_2043,N_2023);
nand U3640 (N_3640,N_2330,N_2231);
or U3641 (N_3641,N_2974,N_2875);
nor U3642 (N_3642,N_2468,N_2645);
nand U3643 (N_3643,N_2282,N_2556);
and U3644 (N_3644,N_2096,N_2783);
nor U3645 (N_3645,N_2027,N_2262);
or U3646 (N_3646,N_2580,N_2076);
or U3647 (N_3647,N_2433,N_2622);
nand U3648 (N_3648,N_2840,N_2151);
and U3649 (N_3649,N_2363,N_2066);
and U3650 (N_3650,N_2884,N_2867);
and U3651 (N_3651,N_2102,N_2023);
or U3652 (N_3652,N_2174,N_2739);
nor U3653 (N_3653,N_2972,N_2916);
nor U3654 (N_3654,N_2168,N_2960);
and U3655 (N_3655,N_2912,N_2307);
nor U3656 (N_3656,N_2256,N_2279);
or U3657 (N_3657,N_2173,N_2424);
nand U3658 (N_3658,N_2084,N_2143);
or U3659 (N_3659,N_2800,N_2429);
and U3660 (N_3660,N_2590,N_2839);
and U3661 (N_3661,N_2370,N_2782);
and U3662 (N_3662,N_2631,N_2661);
nand U3663 (N_3663,N_2632,N_2598);
nor U3664 (N_3664,N_2045,N_2861);
and U3665 (N_3665,N_2971,N_2889);
or U3666 (N_3666,N_2942,N_2546);
nand U3667 (N_3667,N_2810,N_2199);
nand U3668 (N_3668,N_2827,N_2008);
and U3669 (N_3669,N_2749,N_2447);
and U3670 (N_3670,N_2706,N_2285);
or U3671 (N_3671,N_2210,N_2406);
nand U3672 (N_3672,N_2830,N_2721);
and U3673 (N_3673,N_2593,N_2377);
nor U3674 (N_3674,N_2785,N_2101);
or U3675 (N_3675,N_2330,N_2999);
nand U3676 (N_3676,N_2757,N_2418);
or U3677 (N_3677,N_2643,N_2364);
and U3678 (N_3678,N_2189,N_2075);
nor U3679 (N_3679,N_2835,N_2942);
or U3680 (N_3680,N_2030,N_2541);
or U3681 (N_3681,N_2152,N_2628);
or U3682 (N_3682,N_2963,N_2521);
nor U3683 (N_3683,N_2818,N_2184);
and U3684 (N_3684,N_2549,N_2594);
and U3685 (N_3685,N_2458,N_2793);
or U3686 (N_3686,N_2347,N_2592);
or U3687 (N_3687,N_2918,N_2238);
nand U3688 (N_3688,N_2486,N_2230);
nor U3689 (N_3689,N_2464,N_2420);
nand U3690 (N_3690,N_2217,N_2040);
and U3691 (N_3691,N_2482,N_2199);
and U3692 (N_3692,N_2724,N_2587);
nand U3693 (N_3693,N_2804,N_2656);
or U3694 (N_3694,N_2073,N_2321);
nor U3695 (N_3695,N_2998,N_2589);
nand U3696 (N_3696,N_2161,N_2426);
or U3697 (N_3697,N_2874,N_2457);
and U3698 (N_3698,N_2189,N_2582);
or U3699 (N_3699,N_2608,N_2946);
and U3700 (N_3700,N_2084,N_2442);
and U3701 (N_3701,N_2141,N_2726);
and U3702 (N_3702,N_2288,N_2158);
and U3703 (N_3703,N_2129,N_2333);
nor U3704 (N_3704,N_2880,N_2942);
or U3705 (N_3705,N_2316,N_2750);
or U3706 (N_3706,N_2047,N_2764);
nand U3707 (N_3707,N_2685,N_2106);
and U3708 (N_3708,N_2742,N_2525);
nor U3709 (N_3709,N_2048,N_2501);
and U3710 (N_3710,N_2499,N_2767);
xor U3711 (N_3711,N_2194,N_2507);
and U3712 (N_3712,N_2176,N_2977);
and U3713 (N_3713,N_2420,N_2186);
or U3714 (N_3714,N_2018,N_2375);
or U3715 (N_3715,N_2225,N_2244);
or U3716 (N_3716,N_2327,N_2191);
or U3717 (N_3717,N_2471,N_2344);
or U3718 (N_3718,N_2825,N_2321);
and U3719 (N_3719,N_2839,N_2656);
or U3720 (N_3720,N_2242,N_2231);
or U3721 (N_3721,N_2963,N_2226);
nand U3722 (N_3722,N_2865,N_2478);
and U3723 (N_3723,N_2815,N_2571);
or U3724 (N_3724,N_2200,N_2137);
nand U3725 (N_3725,N_2054,N_2168);
or U3726 (N_3726,N_2085,N_2102);
and U3727 (N_3727,N_2159,N_2241);
or U3728 (N_3728,N_2350,N_2472);
and U3729 (N_3729,N_2218,N_2061);
and U3730 (N_3730,N_2828,N_2945);
nand U3731 (N_3731,N_2705,N_2113);
nor U3732 (N_3732,N_2368,N_2787);
or U3733 (N_3733,N_2339,N_2296);
nand U3734 (N_3734,N_2688,N_2013);
nor U3735 (N_3735,N_2537,N_2555);
and U3736 (N_3736,N_2914,N_2091);
or U3737 (N_3737,N_2937,N_2465);
or U3738 (N_3738,N_2981,N_2045);
nand U3739 (N_3739,N_2104,N_2226);
nand U3740 (N_3740,N_2156,N_2281);
and U3741 (N_3741,N_2779,N_2381);
nor U3742 (N_3742,N_2385,N_2306);
and U3743 (N_3743,N_2400,N_2699);
xnor U3744 (N_3744,N_2161,N_2019);
nor U3745 (N_3745,N_2600,N_2729);
nor U3746 (N_3746,N_2723,N_2256);
nor U3747 (N_3747,N_2126,N_2702);
and U3748 (N_3748,N_2025,N_2634);
or U3749 (N_3749,N_2079,N_2813);
or U3750 (N_3750,N_2632,N_2677);
or U3751 (N_3751,N_2602,N_2109);
and U3752 (N_3752,N_2067,N_2217);
nand U3753 (N_3753,N_2975,N_2479);
nand U3754 (N_3754,N_2933,N_2031);
nor U3755 (N_3755,N_2591,N_2484);
and U3756 (N_3756,N_2208,N_2173);
and U3757 (N_3757,N_2157,N_2910);
nand U3758 (N_3758,N_2391,N_2198);
and U3759 (N_3759,N_2031,N_2431);
nor U3760 (N_3760,N_2101,N_2918);
nand U3761 (N_3761,N_2220,N_2013);
nand U3762 (N_3762,N_2444,N_2228);
or U3763 (N_3763,N_2483,N_2785);
and U3764 (N_3764,N_2078,N_2142);
and U3765 (N_3765,N_2964,N_2880);
nor U3766 (N_3766,N_2159,N_2553);
or U3767 (N_3767,N_2167,N_2624);
nor U3768 (N_3768,N_2257,N_2293);
or U3769 (N_3769,N_2471,N_2040);
or U3770 (N_3770,N_2949,N_2716);
or U3771 (N_3771,N_2141,N_2885);
nand U3772 (N_3772,N_2043,N_2646);
nand U3773 (N_3773,N_2304,N_2336);
nor U3774 (N_3774,N_2495,N_2207);
or U3775 (N_3775,N_2147,N_2454);
nand U3776 (N_3776,N_2390,N_2582);
or U3777 (N_3777,N_2045,N_2559);
and U3778 (N_3778,N_2225,N_2295);
nand U3779 (N_3779,N_2750,N_2042);
or U3780 (N_3780,N_2538,N_2758);
nor U3781 (N_3781,N_2330,N_2211);
or U3782 (N_3782,N_2339,N_2276);
or U3783 (N_3783,N_2084,N_2113);
and U3784 (N_3784,N_2784,N_2515);
nand U3785 (N_3785,N_2184,N_2445);
nor U3786 (N_3786,N_2886,N_2712);
xor U3787 (N_3787,N_2438,N_2921);
and U3788 (N_3788,N_2810,N_2267);
nand U3789 (N_3789,N_2611,N_2421);
or U3790 (N_3790,N_2294,N_2708);
nor U3791 (N_3791,N_2220,N_2193);
nand U3792 (N_3792,N_2622,N_2930);
and U3793 (N_3793,N_2969,N_2092);
and U3794 (N_3794,N_2904,N_2278);
and U3795 (N_3795,N_2583,N_2622);
or U3796 (N_3796,N_2693,N_2532);
nor U3797 (N_3797,N_2431,N_2832);
or U3798 (N_3798,N_2499,N_2462);
and U3799 (N_3799,N_2696,N_2370);
nand U3800 (N_3800,N_2876,N_2540);
xor U3801 (N_3801,N_2086,N_2044);
or U3802 (N_3802,N_2245,N_2364);
nor U3803 (N_3803,N_2810,N_2077);
or U3804 (N_3804,N_2579,N_2792);
or U3805 (N_3805,N_2123,N_2996);
xor U3806 (N_3806,N_2322,N_2579);
nand U3807 (N_3807,N_2573,N_2112);
and U3808 (N_3808,N_2947,N_2271);
and U3809 (N_3809,N_2709,N_2559);
and U3810 (N_3810,N_2027,N_2656);
and U3811 (N_3811,N_2437,N_2783);
or U3812 (N_3812,N_2933,N_2870);
nand U3813 (N_3813,N_2983,N_2975);
nor U3814 (N_3814,N_2194,N_2211);
and U3815 (N_3815,N_2892,N_2129);
nand U3816 (N_3816,N_2562,N_2075);
nand U3817 (N_3817,N_2000,N_2269);
nand U3818 (N_3818,N_2991,N_2448);
nor U3819 (N_3819,N_2185,N_2845);
nand U3820 (N_3820,N_2787,N_2774);
and U3821 (N_3821,N_2576,N_2632);
nor U3822 (N_3822,N_2524,N_2967);
nor U3823 (N_3823,N_2494,N_2918);
or U3824 (N_3824,N_2535,N_2843);
xnor U3825 (N_3825,N_2294,N_2373);
nand U3826 (N_3826,N_2731,N_2396);
or U3827 (N_3827,N_2346,N_2117);
nor U3828 (N_3828,N_2914,N_2752);
and U3829 (N_3829,N_2198,N_2442);
nand U3830 (N_3830,N_2658,N_2508);
nor U3831 (N_3831,N_2948,N_2334);
or U3832 (N_3832,N_2647,N_2967);
nor U3833 (N_3833,N_2996,N_2565);
or U3834 (N_3834,N_2796,N_2391);
nand U3835 (N_3835,N_2278,N_2566);
and U3836 (N_3836,N_2183,N_2343);
nand U3837 (N_3837,N_2705,N_2749);
or U3838 (N_3838,N_2154,N_2615);
nor U3839 (N_3839,N_2445,N_2021);
or U3840 (N_3840,N_2341,N_2528);
nand U3841 (N_3841,N_2056,N_2321);
or U3842 (N_3842,N_2957,N_2884);
or U3843 (N_3843,N_2950,N_2371);
or U3844 (N_3844,N_2412,N_2449);
nand U3845 (N_3845,N_2326,N_2749);
and U3846 (N_3846,N_2751,N_2465);
nand U3847 (N_3847,N_2604,N_2066);
nand U3848 (N_3848,N_2268,N_2256);
nand U3849 (N_3849,N_2630,N_2411);
nand U3850 (N_3850,N_2585,N_2083);
nand U3851 (N_3851,N_2521,N_2275);
or U3852 (N_3852,N_2757,N_2357);
nor U3853 (N_3853,N_2352,N_2592);
nor U3854 (N_3854,N_2344,N_2764);
nor U3855 (N_3855,N_2492,N_2407);
nand U3856 (N_3856,N_2239,N_2713);
nor U3857 (N_3857,N_2638,N_2355);
or U3858 (N_3858,N_2935,N_2631);
and U3859 (N_3859,N_2829,N_2937);
nor U3860 (N_3860,N_2060,N_2907);
nor U3861 (N_3861,N_2601,N_2568);
xnor U3862 (N_3862,N_2848,N_2888);
nor U3863 (N_3863,N_2970,N_2141);
nor U3864 (N_3864,N_2869,N_2865);
and U3865 (N_3865,N_2792,N_2532);
and U3866 (N_3866,N_2423,N_2744);
and U3867 (N_3867,N_2443,N_2143);
and U3868 (N_3868,N_2086,N_2067);
nand U3869 (N_3869,N_2936,N_2970);
or U3870 (N_3870,N_2239,N_2992);
xnor U3871 (N_3871,N_2832,N_2400);
nand U3872 (N_3872,N_2645,N_2143);
nor U3873 (N_3873,N_2846,N_2527);
or U3874 (N_3874,N_2044,N_2632);
nor U3875 (N_3875,N_2081,N_2910);
and U3876 (N_3876,N_2330,N_2997);
nand U3877 (N_3877,N_2336,N_2168);
nor U3878 (N_3878,N_2612,N_2261);
nor U3879 (N_3879,N_2695,N_2665);
or U3880 (N_3880,N_2057,N_2532);
nor U3881 (N_3881,N_2770,N_2944);
and U3882 (N_3882,N_2777,N_2411);
or U3883 (N_3883,N_2564,N_2148);
and U3884 (N_3884,N_2346,N_2560);
or U3885 (N_3885,N_2464,N_2121);
and U3886 (N_3886,N_2296,N_2438);
or U3887 (N_3887,N_2828,N_2595);
nor U3888 (N_3888,N_2574,N_2329);
or U3889 (N_3889,N_2999,N_2782);
and U3890 (N_3890,N_2407,N_2841);
nand U3891 (N_3891,N_2694,N_2018);
nor U3892 (N_3892,N_2567,N_2725);
nand U3893 (N_3893,N_2107,N_2567);
and U3894 (N_3894,N_2647,N_2871);
nor U3895 (N_3895,N_2816,N_2353);
nor U3896 (N_3896,N_2395,N_2425);
nand U3897 (N_3897,N_2826,N_2330);
nor U3898 (N_3898,N_2947,N_2641);
or U3899 (N_3899,N_2843,N_2858);
nand U3900 (N_3900,N_2759,N_2078);
nand U3901 (N_3901,N_2853,N_2149);
and U3902 (N_3902,N_2828,N_2056);
nor U3903 (N_3903,N_2239,N_2838);
nand U3904 (N_3904,N_2004,N_2928);
or U3905 (N_3905,N_2311,N_2820);
nand U3906 (N_3906,N_2594,N_2255);
and U3907 (N_3907,N_2900,N_2677);
nand U3908 (N_3908,N_2111,N_2164);
and U3909 (N_3909,N_2439,N_2618);
nand U3910 (N_3910,N_2059,N_2585);
or U3911 (N_3911,N_2851,N_2768);
and U3912 (N_3912,N_2676,N_2205);
and U3913 (N_3913,N_2249,N_2336);
and U3914 (N_3914,N_2581,N_2128);
or U3915 (N_3915,N_2849,N_2127);
and U3916 (N_3916,N_2538,N_2325);
nand U3917 (N_3917,N_2219,N_2308);
and U3918 (N_3918,N_2762,N_2060);
or U3919 (N_3919,N_2176,N_2044);
nor U3920 (N_3920,N_2950,N_2808);
nand U3921 (N_3921,N_2126,N_2794);
and U3922 (N_3922,N_2025,N_2898);
or U3923 (N_3923,N_2430,N_2574);
xor U3924 (N_3924,N_2635,N_2296);
nand U3925 (N_3925,N_2413,N_2075);
nand U3926 (N_3926,N_2281,N_2172);
and U3927 (N_3927,N_2580,N_2798);
and U3928 (N_3928,N_2165,N_2971);
nor U3929 (N_3929,N_2687,N_2213);
or U3930 (N_3930,N_2526,N_2613);
or U3931 (N_3931,N_2836,N_2193);
nor U3932 (N_3932,N_2101,N_2710);
or U3933 (N_3933,N_2336,N_2586);
or U3934 (N_3934,N_2302,N_2030);
and U3935 (N_3935,N_2108,N_2513);
nor U3936 (N_3936,N_2220,N_2991);
nand U3937 (N_3937,N_2641,N_2608);
or U3938 (N_3938,N_2668,N_2693);
nor U3939 (N_3939,N_2718,N_2204);
or U3940 (N_3940,N_2389,N_2326);
nand U3941 (N_3941,N_2285,N_2618);
or U3942 (N_3942,N_2896,N_2981);
or U3943 (N_3943,N_2779,N_2066);
nand U3944 (N_3944,N_2080,N_2430);
nor U3945 (N_3945,N_2480,N_2291);
nor U3946 (N_3946,N_2390,N_2106);
and U3947 (N_3947,N_2978,N_2124);
nand U3948 (N_3948,N_2150,N_2275);
nor U3949 (N_3949,N_2817,N_2645);
nand U3950 (N_3950,N_2266,N_2733);
or U3951 (N_3951,N_2732,N_2259);
and U3952 (N_3952,N_2763,N_2862);
or U3953 (N_3953,N_2609,N_2796);
nand U3954 (N_3954,N_2149,N_2197);
or U3955 (N_3955,N_2763,N_2247);
or U3956 (N_3956,N_2183,N_2990);
nor U3957 (N_3957,N_2558,N_2953);
or U3958 (N_3958,N_2834,N_2358);
or U3959 (N_3959,N_2777,N_2723);
nor U3960 (N_3960,N_2423,N_2447);
and U3961 (N_3961,N_2660,N_2907);
or U3962 (N_3962,N_2035,N_2716);
nand U3963 (N_3963,N_2339,N_2329);
nor U3964 (N_3964,N_2134,N_2656);
nand U3965 (N_3965,N_2231,N_2895);
or U3966 (N_3966,N_2655,N_2001);
and U3967 (N_3967,N_2356,N_2669);
nand U3968 (N_3968,N_2610,N_2411);
nor U3969 (N_3969,N_2030,N_2143);
nor U3970 (N_3970,N_2187,N_2118);
nand U3971 (N_3971,N_2590,N_2919);
nand U3972 (N_3972,N_2271,N_2416);
or U3973 (N_3973,N_2048,N_2816);
and U3974 (N_3974,N_2760,N_2646);
nand U3975 (N_3975,N_2865,N_2265);
nand U3976 (N_3976,N_2399,N_2781);
nand U3977 (N_3977,N_2699,N_2457);
and U3978 (N_3978,N_2758,N_2431);
nor U3979 (N_3979,N_2731,N_2698);
nor U3980 (N_3980,N_2841,N_2761);
and U3981 (N_3981,N_2292,N_2960);
nor U3982 (N_3982,N_2217,N_2720);
or U3983 (N_3983,N_2354,N_2697);
nor U3984 (N_3984,N_2529,N_2876);
nor U3985 (N_3985,N_2421,N_2928);
and U3986 (N_3986,N_2933,N_2694);
or U3987 (N_3987,N_2347,N_2021);
nor U3988 (N_3988,N_2231,N_2521);
nand U3989 (N_3989,N_2949,N_2989);
or U3990 (N_3990,N_2529,N_2891);
or U3991 (N_3991,N_2537,N_2172);
nor U3992 (N_3992,N_2074,N_2017);
or U3993 (N_3993,N_2388,N_2899);
or U3994 (N_3994,N_2770,N_2570);
nor U3995 (N_3995,N_2797,N_2004);
and U3996 (N_3996,N_2902,N_2140);
or U3997 (N_3997,N_2926,N_2540);
or U3998 (N_3998,N_2354,N_2525);
nand U3999 (N_3999,N_2612,N_2918);
or U4000 (N_4000,N_3407,N_3146);
nor U4001 (N_4001,N_3937,N_3985);
and U4002 (N_4002,N_3173,N_3723);
nand U4003 (N_4003,N_3817,N_3300);
nor U4004 (N_4004,N_3968,N_3672);
nor U4005 (N_4005,N_3707,N_3896);
nand U4006 (N_4006,N_3581,N_3919);
nor U4007 (N_4007,N_3386,N_3075);
nor U4008 (N_4008,N_3463,N_3219);
and U4009 (N_4009,N_3340,N_3806);
nand U4010 (N_4010,N_3390,N_3466);
or U4011 (N_4011,N_3876,N_3766);
nand U4012 (N_4012,N_3415,N_3002);
nor U4013 (N_4013,N_3825,N_3811);
or U4014 (N_4014,N_3755,N_3349);
and U4015 (N_4015,N_3622,N_3813);
nand U4016 (N_4016,N_3409,N_3064);
nor U4017 (N_4017,N_3408,N_3007);
nor U4018 (N_4018,N_3229,N_3322);
or U4019 (N_4019,N_3240,N_3363);
or U4020 (N_4020,N_3104,N_3788);
nand U4021 (N_4021,N_3258,N_3579);
nand U4022 (N_4022,N_3112,N_3997);
nor U4023 (N_4023,N_3973,N_3103);
and U4024 (N_4024,N_3865,N_3017);
nand U4025 (N_4025,N_3126,N_3656);
nor U4026 (N_4026,N_3781,N_3278);
nand U4027 (N_4027,N_3892,N_3936);
nand U4028 (N_4028,N_3701,N_3617);
or U4029 (N_4029,N_3334,N_3124);
xor U4030 (N_4030,N_3204,N_3249);
nor U4031 (N_4031,N_3547,N_3418);
nand U4032 (N_4032,N_3900,N_3506);
nor U4033 (N_4033,N_3612,N_3795);
nand U4034 (N_4034,N_3444,N_3142);
nor U4035 (N_4035,N_3328,N_3930);
or U4036 (N_4036,N_3089,N_3712);
or U4037 (N_4037,N_3306,N_3776);
nand U4038 (N_4038,N_3875,N_3551);
nor U4039 (N_4039,N_3646,N_3824);
nor U4040 (N_4040,N_3207,N_3090);
and U4041 (N_4041,N_3108,N_3560);
or U4042 (N_4042,N_3220,N_3375);
or U4043 (N_4043,N_3161,N_3574);
nor U4044 (N_4044,N_3593,N_3880);
nand U4045 (N_4045,N_3762,N_3016);
nor U4046 (N_4046,N_3800,N_3809);
nand U4047 (N_4047,N_3969,N_3518);
nand U4048 (N_4048,N_3623,N_3804);
nor U4049 (N_4049,N_3264,N_3354);
nand U4050 (N_4050,N_3828,N_3699);
and U4051 (N_4051,N_3736,N_3850);
or U4052 (N_4052,N_3199,N_3535);
nand U4053 (N_4053,N_3761,N_3129);
nand U4054 (N_4054,N_3687,N_3834);
nor U4055 (N_4055,N_3096,N_3905);
nand U4056 (N_4056,N_3397,N_3269);
or U4057 (N_4057,N_3820,N_3056);
and U4058 (N_4058,N_3946,N_3150);
and U4059 (N_4059,N_3521,N_3226);
nor U4060 (N_4060,N_3185,N_3356);
nor U4061 (N_4061,N_3830,N_3838);
and U4062 (N_4062,N_3121,N_3291);
nand U4063 (N_4063,N_3345,N_3095);
and U4064 (N_4064,N_3538,N_3401);
or U4065 (N_4065,N_3643,N_3495);
or U4066 (N_4066,N_3792,N_3323);
nand U4067 (N_4067,N_3829,N_3594);
or U4068 (N_4068,N_3853,N_3637);
or U4069 (N_4069,N_3517,N_3505);
or U4070 (N_4070,N_3391,N_3476);
nand U4071 (N_4071,N_3599,N_3998);
and U4072 (N_4072,N_3042,N_3948);
nor U4073 (N_4073,N_3995,N_3198);
and U4074 (N_4074,N_3533,N_3667);
or U4075 (N_4075,N_3182,N_3071);
and U4076 (N_4076,N_3559,N_3057);
and U4077 (N_4077,N_3421,N_3496);
or U4078 (N_4078,N_3326,N_3670);
or U4079 (N_4079,N_3065,N_3282);
and U4080 (N_4080,N_3172,N_3020);
and U4081 (N_4081,N_3629,N_3888);
nand U4082 (N_4082,N_3293,N_3426);
and U4083 (N_4083,N_3636,N_3965);
and U4084 (N_4084,N_3436,N_3718);
and U4085 (N_4085,N_3531,N_3890);
nor U4086 (N_4086,N_3159,N_3926);
nand U4087 (N_4087,N_3835,N_3131);
and U4088 (N_4088,N_3215,N_3524);
or U4089 (N_4089,N_3493,N_3190);
or U4090 (N_4090,N_3125,N_3152);
nor U4091 (N_4091,N_3414,N_3992);
nand U4092 (N_4092,N_3254,N_3674);
nor U4093 (N_4093,N_3200,N_3743);
nand U4094 (N_4094,N_3605,N_3251);
nand U4095 (N_4095,N_3324,N_3958);
and U4096 (N_4096,N_3649,N_3727);
or U4097 (N_4097,N_3522,N_3194);
nor U4098 (N_4098,N_3230,N_3309);
or U4099 (N_4099,N_3592,N_3255);
or U4100 (N_4100,N_3253,N_3641);
nand U4101 (N_4101,N_3999,N_3782);
and U4102 (N_4102,N_3840,N_3621);
and U4103 (N_4103,N_3877,N_3740);
nand U4104 (N_4104,N_3256,N_3777);
or U4105 (N_4105,N_3549,N_3921);
or U4106 (N_4106,N_3779,N_3537);
xor U4107 (N_4107,N_3044,N_3805);
nor U4108 (N_4108,N_3856,N_3686);
nand U4109 (N_4109,N_3205,N_3529);
or U4110 (N_4110,N_3899,N_3303);
and U4111 (N_4111,N_3675,N_3050);
and U4112 (N_4112,N_3376,N_3515);
nand U4113 (N_4113,N_3177,N_3758);
nor U4114 (N_4114,N_3232,N_3962);
nor U4115 (N_4115,N_3127,N_3508);
and U4116 (N_4116,N_3210,N_3261);
and U4117 (N_4117,N_3315,N_3677);
nand U4118 (N_4118,N_3960,N_3000);
nor U4119 (N_4119,N_3704,N_3783);
and U4120 (N_4120,N_3941,N_3548);
nor U4121 (N_4121,N_3787,N_3541);
nor U4122 (N_4122,N_3473,N_3650);
or U4123 (N_4123,N_3332,N_3380);
nand U4124 (N_4124,N_3149,N_3713);
or U4125 (N_4125,N_3456,N_3437);
nor U4126 (N_4126,N_3932,N_3903);
nor U4127 (N_4127,N_3005,N_3336);
nand U4128 (N_4128,N_3063,N_3308);
nor U4129 (N_4129,N_3383,N_3494);
and U4130 (N_4130,N_3355,N_3491);
nor U4131 (N_4131,N_3534,N_3582);
nor U4132 (N_4132,N_3250,N_3163);
and U4133 (N_4133,N_3079,N_3981);
and U4134 (N_4134,N_3708,N_3441);
or U4135 (N_4135,N_3902,N_3123);
nand U4136 (N_4136,N_3242,N_3399);
or U4137 (N_4137,N_3682,N_3994);
or U4138 (N_4138,N_3180,N_3618);
nand U4139 (N_4139,N_3338,N_3731);
nor U4140 (N_4140,N_3717,N_3480);
or U4141 (N_4141,N_3514,N_3839);
nor U4142 (N_4142,N_3128,N_3223);
and U4143 (N_4143,N_3798,N_3891);
xnor U4144 (N_4144,N_3351,N_3595);
nand U4145 (N_4145,N_3344,N_3848);
nor U4146 (N_4146,N_3162,N_3633);
nand U4147 (N_4147,N_3187,N_3241);
nand U4148 (N_4148,N_3353,N_3728);
or U4149 (N_4149,N_3741,N_3272);
nor U4150 (N_4150,N_3849,N_3091);
and U4151 (N_4151,N_3923,N_3909);
nor U4152 (N_4152,N_3852,N_3043);
nand U4153 (N_4153,N_3745,N_3742);
xor U4154 (N_4154,N_3014,N_3673);
nand U4155 (N_4155,N_3765,N_3558);
and U4156 (N_4156,N_3305,N_3319);
nor U4157 (N_4157,N_3572,N_3959);
nand U4158 (N_4158,N_3233,N_3512);
nor U4159 (N_4159,N_3317,N_3274);
nor U4160 (N_4160,N_3485,N_3081);
nand U4161 (N_4161,N_3341,N_3078);
xor U4162 (N_4162,N_3647,N_3614);
nand U4163 (N_4163,N_3598,N_3964);
nor U4164 (N_4164,N_3296,N_3939);
nand U4165 (N_4165,N_3520,N_3024);
nor U4166 (N_4166,N_3843,N_3752);
and U4167 (N_4167,N_3097,N_3329);
and U4168 (N_4168,N_3694,N_3860);
and U4169 (N_4169,N_3294,N_3312);
nand U4170 (N_4170,N_3733,N_3734);
nand U4171 (N_4171,N_3299,N_3597);
nand U4172 (N_4172,N_3883,N_3420);
nor U4173 (N_4173,N_3797,N_3577);
nand U4174 (N_4174,N_3974,N_3009);
or U4175 (N_4175,N_3822,N_3952);
and U4176 (N_4176,N_3991,N_3271);
nor U4177 (N_4177,N_3661,N_3279);
and U4178 (N_4178,N_3318,N_3311);
nor U4179 (N_4179,N_3055,N_3034);
and U4180 (N_4180,N_3568,N_3789);
and U4181 (N_4181,N_3449,N_3113);
nor U4182 (N_4182,N_3403,N_3133);
or U4183 (N_4183,N_3450,N_3513);
nand U4184 (N_4184,N_3640,N_3543);
nor U4185 (N_4185,N_3720,N_3243);
or U4186 (N_4186,N_3735,N_3083);
nor U4187 (N_4187,N_3553,N_3845);
and U4188 (N_4188,N_3955,N_3949);
and U4189 (N_4189,N_3008,N_3033);
and U4190 (N_4190,N_3257,N_3151);
and U4191 (N_4191,N_3897,N_3417);
nor U4192 (N_4192,N_3693,N_3924);
nor U4193 (N_4193,N_3362,N_3881);
nor U4194 (N_4194,N_3051,N_3756);
nor U4195 (N_4195,N_3760,N_3287);
nor U4196 (N_4196,N_3611,N_3490);
and U4197 (N_4197,N_3389,N_3392);
or U4198 (N_4198,N_3655,N_3346);
nor U4199 (N_4199,N_3327,N_3596);
or U4200 (N_4200,N_3459,N_3382);
nand U4201 (N_4201,N_3228,N_3801);
nor U4202 (N_4202,N_3950,N_3681);
nand U4203 (N_4203,N_3747,N_3422);
nand U4204 (N_4204,N_3715,N_3953);
and U4205 (N_4205,N_3556,N_3912);
nor U4206 (N_4206,N_3966,N_3486);
nor U4207 (N_4207,N_3904,N_3343);
nand U4208 (N_4208,N_3405,N_3685);
and U4209 (N_4209,N_3542,N_3583);
or U4210 (N_4210,N_3385,N_3202);
nand U4211 (N_4211,N_3726,N_3652);
nor U4212 (N_4212,N_3604,N_3144);
xnor U4213 (N_4213,N_3893,N_3359);
nor U4214 (N_4214,N_3206,N_3624);
or U4215 (N_4215,N_3259,N_3642);
nand U4216 (N_4216,N_3276,N_3455);
and U4217 (N_4217,N_3679,N_3431);
and U4218 (N_4218,N_3908,N_3290);
nand U4219 (N_4219,N_3245,N_3213);
and U4220 (N_4220,N_3406,N_3680);
or U4221 (N_4221,N_3361,N_3504);
nand U4222 (N_4222,N_3688,N_3561);
and U4223 (N_4223,N_3136,N_3193);
and U4224 (N_4224,N_3895,N_3234);
nand U4225 (N_4225,N_3634,N_3333);
and U4226 (N_4226,N_3662,N_3286);
nand U4227 (N_4227,N_3010,N_3140);
or U4228 (N_4228,N_3979,N_3778);
or U4229 (N_4229,N_3393,N_3868);
and U4230 (N_4230,N_3698,N_3690);
nand U4231 (N_4231,N_3130,N_3748);
nor U4232 (N_4232,N_3217,N_3192);
or U4233 (N_4233,N_3993,N_3818);
nand U4234 (N_4234,N_3411,N_3982);
and U4235 (N_4235,N_3608,N_3247);
nand U4236 (N_4236,N_3567,N_3196);
or U4237 (N_4237,N_3216,N_3874);
nand U4238 (N_4238,N_3587,N_3030);
nor U4239 (N_4239,N_3181,N_3358);
or U4240 (N_4240,N_3158,N_3188);
nand U4241 (N_4241,N_3739,N_3153);
nand U4242 (N_4242,N_3102,N_3208);
nand U4243 (N_4243,N_3658,N_3238);
and U4244 (N_4244,N_3350,N_3252);
nand U4245 (N_4245,N_3387,N_3475);
nor U4246 (N_4246,N_3714,N_3638);
nor U4247 (N_4247,N_3951,N_3934);
or U4248 (N_4248,N_3148,N_3211);
nor U4249 (N_4249,N_3544,N_3184);
and U4250 (N_4250,N_3432,N_3100);
and U4251 (N_4251,N_3085,N_3447);
nor U4252 (N_4252,N_3773,N_3659);
and U4253 (N_4253,N_3786,N_3471);
and U4254 (N_4254,N_3774,N_3566);
or U4255 (N_4255,N_3157,N_3092);
nor U4256 (N_4256,N_3764,N_3225);
nand U4257 (N_4257,N_3283,N_3369);
or U4258 (N_4258,N_3268,N_3942);
and U4259 (N_4259,N_3983,N_3218);
nand U4260 (N_4260,N_3027,N_3052);
nor U4261 (N_4261,N_3702,N_3001);
nor U4262 (N_4262,N_3678,N_3469);
or U4263 (N_4263,N_3844,N_3878);
nand U4264 (N_4264,N_3691,N_3070);
xnor U4265 (N_4265,N_3719,N_3928);
or U4266 (N_4266,N_3546,N_3540);
or U4267 (N_4267,N_3458,N_3668);
nor U4268 (N_4268,N_3137,N_3562);
nor U4269 (N_4269,N_3307,N_3370);
nor U4270 (N_4270,N_3442,N_3313);
and U4271 (N_4271,N_3922,N_3780);
nand U4272 (N_4272,N_3488,N_3262);
or U4273 (N_4273,N_3413,N_3607);
nor U4274 (N_4274,N_3115,N_3901);
nor U4275 (N_4275,N_3267,N_3224);
nor U4276 (N_4276,N_3302,N_3298);
and U4277 (N_4277,N_3933,N_3569);
and U4278 (N_4278,N_3189,N_3074);
and U4279 (N_4279,N_3671,N_3796);
and U4280 (N_4280,N_3601,N_3976);
nor U4281 (N_4281,N_3894,N_3703);
nor U4282 (N_4282,N_3613,N_3626);
nor U4283 (N_4283,N_3222,N_3402);
nor U4284 (N_4284,N_3335,N_3147);
nor U4285 (N_4285,N_3037,N_3816);
and U4286 (N_4286,N_3470,N_3235);
and U4287 (N_4287,N_3460,N_3859);
xnor U4288 (N_4288,N_3168,N_3648);
and U4289 (N_4289,N_3114,N_3700);
or U4290 (N_4290,N_3156,N_3676);
and U4291 (N_4291,N_3132,N_3653);
or U4292 (N_4292,N_3011,N_3482);
and U4293 (N_4293,N_3221,N_3812);
nor U4294 (N_4294,N_3663,N_3575);
or U4295 (N_4295,N_3590,N_3101);
nor U4296 (N_4296,N_3454,N_3012);
nor U4297 (N_4297,N_3526,N_3589);
or U4298 (N_4298,N_3031,N_3209);
nand U4299 (N_4299,N_3093,N_3425);
nand U4300 (N_4300,N_3077,N_3275);
nor U4301 (N_4301,N_3368,N_3725);
and U4302 (N_4302,N_3372,N_3836);
nand U4303 (N_4303,N_3578,N_3944);
or U4304 (N_4304,N_3635,N_3381);
or U4305 (N_4305,N_3863,N_3873);
or U4306 (N_4306,N_3987,N_3183);
nand U4307 (N_4307,N_3082,N_3374);
and U4308 (N_4308,N_3195,N_3918);
and U4309 (N_4309,N_3956,N_3775);
or U4310 (N_4310,N_3054,N_3957);
nand U4311 (N_4311,N_3419,N_3111);
nor U4312 (N_4312,N_3706,N_3310);
nand U4313 (N_4313,N_3348,N_3019);
and U4314 (N_4314,N_3331,N_3400);
nand U4315 (N_4315,N_3632,N_3477);
nor U4316 (N_4316,N_3472,N_3439);
nor U4317 (N_4317,N_3889,N_3174);
or U4318 (N_4318,N_3378,N_3554);
nand U4319 (N_4319,N_3099,N_3525);
or U4320 (N_4320,N_3297,N_3815);
nor U4321 (N_4321,N_3076,N_3106);
nand U4322 (N_4322,N_3823,N_3519);
nand U4323 (N_4323,N_3316,N_3068);
and U4324 (N_4324,N_3060,N_3277);
nor U4325 (N_4325,N_3032,N_3048);
nor U4326 (N_4326,N_3847,N_3248);
or U4327 (N_4327,N_3730,N_3620);
or U4328 (N_4328,N_3175,N_3664);
and U4329 (N_4329,N_3457,N_3138);
nand U4330 (N_4330,N_3872,N_3869);
nand U4331 (N_4331,N_3013,N_3810);
and U4332 (N_4332,N_3603,N_3487);
nand U4333 (N_4333,N_3141,N_3084);
nor U4334 (N_4334,N_3281,N_3026);
nor U4335 (N_4335,N_3588,N_3885);
nor U4336 (N_4336,N_3186,N_3263);
or U4337 (N_4337,N_3862,N_3201);
nand U4338 (N_4338,N_3479,N_3120);
and U4339 (N_4339,N_3073,N_3749);
nand U4340 (N_4340,N_3285,N_3062);
nand U4341 (N_4341,N_3631,N_3669);
and U4342 (N_4342,N_3584,N_3814);
or U4343 (N_4343,N_3036,N_3967);
nand U4344 (N_4344,N_3139,N_3645);
or U4345 (N_4345,N_3492,N_3040);
nand U4346 (N_4346,N_3970,N_3750);
nor U4347 (N_4347,N_3438,N_3284);
nor U4348 (N_4348,N_3006,N_3925);
nor U4349 (N_4349,N_3705,N_3366);
or U4350 (N_4350,N_3906,N_3627);
nor U4351 (N_4351,N_3695,N_3122);
or U4352 (N_4352,N_3791,N_3398);
nand U4353 (N_4353,N_3940,N_3088);
or U4354 (N_4354,N_3882,N_3029);
or U4355 (N_4355,N_3511,N_3164);
nand U4356 (N_4356,N_3325,N_3550);
nand U4357 (N_4357,N_3018,N_3746);
or U4358 (N_4358,N_3377,N_3565);
or U4359 (N_4359,N_3364,N_3167);
and U4360 (N_4360,N_3692,N_3320);
nor U4361 (N_4361,N_3683,N_3769);
nor U4362 (N_4362,N_3911,N_3292);
and U4363 (N_4363,N_3654,N_3119);
and U4364 (N_4364,N_3722,N_3059);
or U4365 (N_4365,N_3500,N_3360);
nand U4366 (N_4366,N_3929,N_3996);
or U4367 (N_4367,N_3003,N_3841);
nand U4368 (N_4368,N_3481,N_3468);
and U4369 (N_4369,N_3857,N_3799);
and U4370 (N_4370,N_3528,N_3886);
nor U4371 (N_4371,N_3023,N_3977);
and U4372 (N_4372,N_3552,N_3523);
nor U4373 (N_4373,N_3423,N_3047);
nor U4374 (N_4374,N_3467,N_3980);
nor U4375 (N_4375,N_3434,N_3866);
and U4376 (N_4376,N_3465,N_3270);
nor U4377 (N_4377,N_3831,N_3166);
or U4378 (N_4378,N_3709,N_3619);
nand U4379 (N_4379,N_3931,N_3972);
nand U4380 (N_4380,N_3767,N_3118);
or U4381 (N_4381,N_3913,N_3807);
and U4382 (N_4382,N_3260,N_3171);
nor U4383 (N_4383,N_3445,N_3753);
nand U4384 (N_4384,N_3867,N_3563);
or U4385 (N_4385,N_3819,N_3330);
nor U4386 (N_4386,N_3833,N_3802);
nand U4387 (N_4387,N_3046,N_3484);
and U4388 (N_4388,N_3105,N_3038);
and U4389 (N_4389,N_3295,N_3134);
nand U4390 (N_4390,N_3145,N_3094);
nand U4391 (N_4391,N_3989,N_3160);
nand U4392 (N_4392,N_3304,N_3975);
nor U4393 (N_4393,N_3532,N_3770);
nor U4394 (N_4394,N_3069,N_3696);
nor U4395 (N_4395,N_3015,N_3665);
or U4396 (N_4396,N_3751,N_3724);
or U4397 (N_4397,N_3342,N_3729);
nor U4398 (N_4398,N_3971,N_3864);
and U4399 (N_4399,N_3154,N_3887);
or U4400 (N_4400,N_3428,N_3367);
or U4401 (N_4401,N_3625,N_3738);
nand U4402 (N_4402,N_3388,N_3314);
and U4403 (N_4403,N_3280,N_3808);
nor U4404 (N_4404,N_3214,N_3914);
and U4405 (N_4405,N_3396,N_3961);
or U4406 (N_4406,N_3510,N_3516);
nor U4407 (N_4407,N_3938,N_3754);
or U4408 (N_4408,N_3539,N_3412);
or U4409 (N_4409,N_3203,N_3087);
nand U4410 (N_4410,N_3462,N_3630);
nand U4411 (N_4411,N_3854,N_3498);
and U4412 (N_4412,N_3502,N_3446);
nand U4413 (N_4413,N_3440,N_3404);
and U4414 (N_4414,N_3337,N_3651);
nor U4415 (N_4415,N_3710,N_3107);
nand U4416 (N_4416,N_3321,N_3945);
nor U4417 (N_4417,N_3288,N_3947);
or U4418 (N_4418,N_3116,N_3497);
or U4419 (N_4419,N_3430,N_3022);
or U4420 (N_4420,N_3616,N_3759);
or U4421 (N_4421,N_3155,N_3035);
or U4422 (N_4422,N_3803,N_3237);
nand U4423 (N_4423,N_3489,N_3602);
nor U4424 (N_4424,N_3564,N_3433);
nand U4425 (N_4425,N_3744,N_3339);
or U4426 (N_4426,N_3884,N_3660);
nor U4427 (N_4427,N_3273,N_3898);
nand U4428 (N_4428,N_3684,N_3570);
xor U4429 (N_4429,N_3110,N_3143);
and U4430 (N_4430,N_3394,N_3178);
and U4431 (N_4431,N_3794,N_3169);
or U4432 (N_4432,N_3067,N_3785);
or U4433 (N_4433,N_3371,N_3827);
nand U4434 (N_4434,N_3666,N_3086);
nand U4435 (N_4435,N_3191,N_3910);
and U4436 (N_4436,N_3545,N_3427);
and U4437 (N_4437,N_3080,N_3429);
nor U4438 (N_4438,N_3793,N_3301);
or U4439 (N_4439,N_3609,N_3265);
or U4440 (N_4440,N_3176,N_3557);
or U4441 (N_4441,N_3049,N_3855);
or U4442 (N_4442,N_3451,N_3870);
nand U4443 (N_4443,N_3984,N_3117);
or U4444 (N_4444,N_3165,N_3935);
nand U4445 (N_4445,N_3580,N_3507);
and U4446 (N_4446,N_3058,N_3025);
nor U4447 (N_4447,N_3066,N_3053);
nand U4448 (N_4448,N_3555,N_3461);
or U4449 (N_4449,N_3072,N_3536);
nor U4450 (N_4450,N_3790,N_3721);
nand U4451 (N_4451,N_3435,N_3763);
nand U4452 (N_4452,N_3907,N_3347);
xor U4453 (N_4453,N_3639,N_3716);
nand U4454 (N_4454,N_3109,N_3606);
nand U4455 (N_4455,N_3576,N_3448);
and U4456 (N_4456,N_3920,N_3135);
or U4457 (N_4457,N_3990,N_3615);
and U4458 (N_4458,N_3917,N_3499);
nand U4459 (N_4459,N_3657,N_3357);
nand U4460 (N_4460,N_3028,N_3530);
or U4461 (N_4461,N_3197,N_3021);
nand U4462 (N_4462,N_3689,N_3861);
and U4463 (N_4463,N_3464,N_3978);
nand U4464 (N_4464,N_3098,N_3170);
nor U4465 (N_4465,N_3986,N_3289);
nor U4466 (N_4466,N_3503,N_3943);
or U4467 (N_4467,N_3711,N_3352);
nor U4468 (N_4468,N_3610,N_3478);
or U4469 (N_4469,N_3585,N_3227);
nor U4470 (N_4470,N_3879,N_3179);
nor U4471 (N_4471,N_3244,N_3365);
or U4472 (N_4472,N_3821,N_3266);
nand U4473 (N_4473,N_3384,N_3916);
nand U4474 (N_4474,N_3246,N_3483);
nand U4475 (N_4475,N_3474,N_3039);
nor U4476 (N_4476,N_3963,N_3732);
and U4477 (N_4477,N_3527,N_3954);
nand U4478 (N_4478,N_3600,N_3239);
nand U4479 (N_4479,N_3988,N_3644);
nor U4480 (N_4480,N_3915,N_3737);
or U4481 (N_4481,N_3768,N_3443);
and U4482 (N_4482,N_3846,N_3373);
nand U4483 (N_4483,N_3772,N_3452);
nand U4484 (N_4484,N_3591,N_3571);
or U4485 (N_4485,N_3041,N_3231);
or U4486 (N_4486,N_3379,N_3927);
nand U4487 (N_4487,N_3424,N_3832);
nand U4488 (N_4488,N_3453,N_3395);
and U4489 (N_4489,N_3236,N_3771);
nand U4490 (N_4490,N_3509,N_3871);
nor U4491 (N_4491,N_3501,N_3586);
nor U4492 (N_4492,N_3628,N_3858);
nand U4493 (N_4493,N_3837,N_3842);
or U4494 (N_4494,N_3410,N_3757);
and U4495 (N_4495,N_3061,N_3045);
nor U4496 (N_4496,N_3416,N_3784);
and U4497 (N_4497,N_3697,N_3851);
nor U4498 (N_4498,N_3573,N_3212);
nand U4499 (N_4499,N_3004,N_3826);
and U4500 (N_4500,N_3432,N_3101);
or U4501 (N_4501,N_3826,N_3179);
and U4502 (N_4502,N_3127,N_3437);
or U4503 (N_4503,N_3499,N_3444);
nand U4504 (N_4504,N_3475,N_3247);
and U4505 (N_4505,N_3232,N_3173);
and U4506 (N_4506,N_3095,N_3335);
and U4507 (N_4507,N_3422,N_3139);
or U4508 (N_4508,N_3955,N_3605);
or U4509 (N_4509,N_3980,N_3893);
and U4510 (N_4510,N_3731,N_3780);
nor U4511 (N_4511,N_3281,N_3506);
nor U4512 (N_4512,N_3588,N_3308);
and U4513 (N_4513,N_3906,N_3269);
nand U4514 (N_4514,N_3587,N_3144);
or U4515 (N_4515,N_3442,N_3696);
nor U4516 (N_4516,N_3323,N_3845);
or U4517 (N_4517,N_3201,N_3633);
nor U4518 (N_4518,N_3289,N_3422);
nand U4519 (N_4519,N_3638,N_3892);
nor U4520 (N_4520,N_3164,N_3589);
nand U4521 (N_4521,N_3209,N_3935);
xor U4522 (N_4522,N_3715,N_3199);
or U4523 (N_4523,N_3784,N_3950);
or U4524 (N_4524,N_3496,N_3327);
or U4525 (N_4525,N_3816,N_3629);
or U4526 (N_4526,N_3146,N_3928);
nor U4527 (N_4527,N_3764,N_3624);
nand U4528 (N_4528,N_3475,N_3168);
and U4529 (N_4529,N_3111,N_3921);
nand U4530 (N_4530,N_3769,N_3090);
nor U4531 (N_4531,N_3585,N_3347);
nand U4532 (N_4532,N_3224,N_3014);
nand U4533 (N_4533,N_3860,N_3195);
nand U4534 (N_4534,N_3472,N_3172);
nor U4535 (N_4535,N_3093,N_3810);
nand U4536 (N_4536,N_3998,N_3333);
nor U4537 (N_4537,N_3127,N_3214);
nor U4538 (N_4538,N_3749,N_3554);
nor U4539 (N_4539,N_3272,N_3665);
or U4540 (N_4540,N_3632,N_3753);
nor U4541 (N_4541,N_3721,N_3676);
nand U4542 (N_4542,N_3570,N_3897);
nor U4543 (N_4543,N_3365,N_3254);
nand U4544 (N_4544,N_3332,N_3089);
and U4545 (N_4545,N_3831,N_3872);
or U4546 (N_4546,N_3580,N_3357);
nor U4547 (N_4547,N_3462,N_3081);
or U4548 (N_4548,N_3244,N_3339);
nor U4549 (N_4549,N_3527,N_3516);
nor U4550 (N_4550,N_3967,N_3802);
or U4551 (N_4551,N_3384,N_3180);
or U4552 (N_4552,N_3552,N_3916);
nand U4553 (N_4553,N_3149,N_3857);
nor U4554 (N_4554,N_3939,N_3617);
nand U4555 (N_4555,N_3591,N_3503);
or U4556 (N_4556,N_3663,N_3578);
nand U4557 (N_4557,N_3610,N_3681);
and U4558 (N_4558,N_3442,N_3227);
or U4559 (N_4559,N_3932,N_3331);
nor U4560 (N_4560,N_3331,N_3489);
nor U4561 (N_4561,N_3979,N_3585);
or U4562 (N_4562,N_3588,N_3909);
nand U4563 (N_4563,N_3330,N_3629);
or U4564 (N_4564,N_3230,N_3773);
and U4565 (N_4565,N_3724,N_3513);
nor U4566 (N_4566,N_3641,N_3955);
and U4567 (N_4567,N_3185,N_3121);
and U4568 (N_4568,N_3370,N_3715);
nand U4569 (N_4569,N_3967,N_3267);
and U4570 (N_4570,N_3912,N_3213);
or U4571 (N_4571,N_3016,N_3157);
nand U4572 (N_4572,N_3351,N_3196);
nand U4573 (N_4573,N_3782,N_3686);
or U4574 (N_4574,N_3189,N_3290);
nand U4575 (N_4575,N_3331,N_3497);
or U4576 (N_4576,N_3006,N_3225);
and U4577 (N_4577,N_3275,N_3676);
nand U4578 (N_4578,N_3584,N_3508);
nand U4579 (N_4579,N_3727,N_3746);
nor U4580 (N_4580,N_3942,N_3726);
or U4581 (N_4581,N_3102,N_3944);
nand U4582 (N_4582,N_3272,N_3189);
nor U4583 (N_4583,N_3319,N_3318);
and U4584 (N_4584,N_3716,N_3880);
nand U4585 (N_4585,N_3899,N_3956);
or U4586 (N_4586,N_3707,N_3668);
nor U4587 (N_4587,N_3006,N_3252);
nand U4588 (N_4588,N_3292,N_3964);
or U4589 (N_4589,N_3603,N_3797);
or U4590 (N_4590,N_3876,N_3648);
xnor U4591 (N_4591,N_3350,N_3775);
and U4592 (N_4592,N_3272,N_3086);
or U4593 (N_4593,N_3286,N_3627);
nor U4594 (N_4594,N_3635,N_3425);
nand U4595 (N_4595,N_3303,N_3456);
and U4596 (N_4596,N_3193,N_3705);
and U4597 (N_4597,N_3171,N_3462);
and U4598 (N_4598,N_3090,N_3180);
nor U4599 (N_4599,N_3400,N_3872);
or U4600 (N_4600,N_3090,N_3071);
nand U4601 (N_4601,N_3666,N_3507);
and U4602 (N_4602,N_3605,N_3384);
nor U4603 (N_4603,N_3627,N_3899);
and U4604 (N_4604,N_3848,N_3392);
nor U4605 (N_4605,N_3689,N_3743);
nor U4606 (N_4606,N_3504,N_3730);
nor U4607 (N_4607,N_3727,N_3788);
or U4608 (N_4608,N_3818,N_3824);
or U4609 (N_4609,N_3045,N_3995);
nor U4610 (N_4610,N_3899,N_3905);
nand U4611 (N_4611,N_3006,N_3996);
nand U4612 (N_4612,N_3115,N_3644);
nand U4613 (N_4613,N_3838,N_3199);
nand U4614 (N_4614,N_3301,N_3970);
nand U4615 (N_4615,N_3817,N_3981);
nor U4616 (N_4616,N_3291,N_3118);
or U4617 (N_4617,N_3382,N_3134);
xnor U4618 (N_4618,N_3505,N_3824);
nand U4619 (N_4619,N_3737,N_3849);
and U4620 (N_4620,N_3747,N_3723);
nor U4621 (N_4621,N_3961,N_3841);
nor U4622 (N_4622,N_3242,N_3472);
nor U4623 (N_4623,N_3368,N_3762);
nor U4624 (N_4624,N_3700,N_3453);
and U4625 (N_4625,N_3683,N_3544);
nor U4626 (N_4626,N_3981,N_3532);
nor U4627 (N_4627,N_3151,N_3790);
or U4628 (N_4628,N_3238,N_3841);
and U4629 (N_4629,N_3700,N_3083);
nand U4630 (N_4630,N_3179,N_3761);
and U4631 (N_4631,N_3759,N_3586);
nand U4632 (N_4632,N_3104,N_3077);
nor U4633 (N_4633,N_3505,N_3362);
nor U4634 (N_4634,N_3340,N_3195);
nor U4635 (N_4635,N_3065,N_3207);
nand U4636 (N_4636,N_3933,N_3367);
nor U4637 (N_4637,N_3395,N_3809);
nand U4638 (N_4638,N_3934,N_3900);
or U4639 (N_4639,N_3165,N_3114);
or U4640 (N_4640,N_3358,N_3497);
or U4641 (N_4641,N_3623,N_3889);
and U4642 (N_4642,N_3916,N_3046);
nor U4643 (N_4643,N_3812,N_3948);
nor U4644 (N_4644,N_3530,N_3954);
or U4645 (N_4645,N_3377,N_3234);
and U4646 (N_4646,N_3024,N_3806);
nor U4647 (N_4647,N_3337,N_3017);
or U4648 (N_4648,N_3814,N_3989);
nand U4649 (N_4649,N_3689,N_3585);
nand U4650 (N_4650,N_3539,N_3929);
or U4651 (N_4651,N_3977,N_3400);
and U4652 (N_4652,N_3371,N_3569);
nor U4653 (N_4653,N_3837,N_3434);
and U4654 (N_4654,N_3472,N_3245);
xnor U4655 (N_4655,N_3833,N_3770);
nor U4656 (N_4656,N_3313,N_3779);
and U4657 (N_4657,N_3110,N_3330);
or U4658 (N_4658,N_3266,N_3964);
nor U4659 (N_4659,N_3257,N_3255);
or U4660 (N_4660,N_3702,N_3309);
or U4661 (N_4661,N_3656,N_3279);
or U4662 (N_4662,N_3615,N_3131);
nor U4663 (N_4663,N_3803,N_3187);
or U4664 (N_4664,N_3662,N_3912);
or U4665 (N_4665,N_3343,N_3071);
and U4666 (N_4666,N_3237,N_3566);
or U4667 (N_4667,N_3963,N_3195);
and U4668 (N_4668,N_3000,N_3371);
and U4669 (N_4669,N_3050,N_3960);
nor U4670 (N_4670,N_3771,N_3020);
nand U4671 (N_4671,N_3131,N_3535);
or U4672 (N_4672,N_3652,N_3159);
nor U4673 (N_4673,N_3886,N_3650);
or U4674 (N_4674,N_3643,N_3821);
or U4675 (N_4675,N_3579,N_3268);
and U4676 (N_4676,N_3793,N_3411);
and U4677 (N_4677,N_3063,N_3053);
nor U4678 (N_4678,N_3870,N_3179);
nor U4679 (N_4679,N_3093,N_3802);
or U4680 (N_4680,N_3140,N_3914);
or U4681 (N_4681,N_3627,N_3299);
or U4682 (N_4682,N_3891,N_3464);
and U4683 (N_4683,N_3906,N_3166);
and U4684 (N_4684,N_3742,N_3835);
nor U4685 (N_4685,N_3596,N_3138);
or U4686 (N_4686,N_3185,N_3312);
nor U4687 (N_4687,N_3185,N_3985);
nand U4688 (N_4688,N_3094,N_3609);
and U4689 (N_4689,N_3265,N_3197);
nand U4690 (N_4690,N_3952,N_3602);
nor U4691 (N_4691,N_3540,N_3846);
nor U4692 (N_4692,N_3964,N_3902);
or U4693 (N_4693,N_3570,N_3058);
nand U4694 (N_4694,N_3107,N_3086);
nor U4695 (N_4695,N_3961,N_3430);
nor U4696 (N_4696,N_3497,N_3837);
and U4697 (N_4697,N_3398,N_3980);
and U4698 (N_4698,N_3482,N_3789);
nand U4699 (N_4699,N_3497,N_3574);
nand U4700 (N_4700,N_3822,N_3108);
nor U4701 (N_4701,N_3876,N_3395);
and U4702 (N_4702,N_3860,N_3390);
and U4703 (N_4703,N_3127,N_3315);
nor U4704 (N_4704,N_3927,N_3690);
and U4705 (N_4705,N_3647,N_3030);
or U4706 (N_4706,N_3335,N_3100);
nor U4707 (N_4707,N_3334,N_3653);
or U4708 (N_4708,N_3412,N_3830);
and U4709 (N_4709,N_3341,N_3257);
nand U4710 (N_4710,N_3639,N_3948);
nor U4711 (N_4711,N_3429,N_3484);
and U4712 (N_4712,N_3767,N_3348);
xor U4713 (N_4713,N_3946,N_3424);
and U4714 (N_4714,N_3120,N_3142);
nor U4715 (N_4715,N_3275,N_3829);
and U4716 (N_4716,N_3165,N_3733);
nand U4717 (N_4717,N_3535,N_3990);
or U4718 (N_4718,N_3900,N_3420);
or U4719 (N_4719,N_3200,N_3907);
and U4720 (N_4720,N_3440,N_3826);
or U4721 (N_4721,N_3491,N_3166);
or U4722 (N_4722,N_3087,N_3374);
or U4723 (N_4723,N_3134,N_3072);
nand U4724 (N_4724,N_3156,N_3720);
or U4725 (N_4725,N_3085,N_3520);
nand U4726 (N_4726,N_3234,N_3793);
and U4727 (N_4727,N_3766,N_3277);
xnor U4728 (N_4728,N_3095,N_3349);
or U4729 (N_4729,N_3927,N_3953);
or U4730 (N_4730,N_3572,N_3138);
nor U4731 (N_4731,N_3570,N_3918);
or U4732 (N_4732,N_3788,N_3889);
and U4733 (N_4733,N_3416,N_3816);
and U4734 (N_4734,N_3165,N_3765);
and U4735 (N_4735,N_3677,N_3234);
nor U4736 (N_4736,N_3325,N_3832);
xor U4737 (N_4737,N_3481,N_3860);
and U4738 (N_4738,N_3929,N_3779);
nand U4739 (N_4739,N_3185,N_3524);
or U4740 (N_4740,N_3215,N_3638);
or U4741 (N_4741,N_3891,N_3662);
and U4742 (N_4742,N_3967,N_3258);
xnor U4743 (N_4743,N_3682,N_3987);
nor U4744 (N_4744,N_3094,N_3007);
nor U4745 (N_4745,N_3657,N_3514);
or U4746 (N_4746,N_3389,N_3051);
and U4747 (N_4747,N_3715,N_3623);
nor U4748 (N_4748,N_3431,N_3573);
and U4749 (N_4749,N_3740,N_3110);
and U4750 (N_4750,N_3292,N_3971);
nor U4751 (N_4751,N_3614,N_3281);
nor U4752 (N_4752,N_3467,N_3701);
and U4753 (N_4753,N_3814,N_3827);
nand U4754 (N_4754,N_3996,N_3762);
nand U4755 (N_4755,N_3949,N_3748);
and U4756 (N_4756,N_3917,N_3491);
and U4757 (N_4757,N_3969,N_3260);
or U4758 (N_4758,N_3542,N_3545);
or U4759 (N_4759,N_3738,N_3641);
or U4760 (N_4760,N_3538,N_3739);
nor U4761 (N_4761,N_3901,N_3540);
nor U4762 (N_4762,N_3374,N_3568);
xnor U4763 (N_4763,N_3885,N_3339);
nor U4764 (N_4764,N_3672,N_3311);
and U4765 (N_4765,N_3567,N_3395);
and U4766 (N_4766,N_3896,N_3956);
or U4767 (N_4767,N_3817,N_3722);
nor U4768 (N_4768,N_3228,N_3009);
nor U4769 (N_4769,N_3766,N_3719);
or U4770 (N_4770,N_3274,N_3239);
or U4771 (N_4771,N_3549,N_3920);
or U4772 (N_4772,N_3780,N_3298);
nor U4773 (N_4773,N_3746,N_3034);
nor U4774 (N_4774,N_3321,N_3015);
and U4775 (N_4775,N_3184,N_3100);
nand U4776 (N_4776,N_3023,N_3109);
and U4777 (N_4777,N_3920,N_3269);
or U4778 (N_4778,N_3876,N_3472);
and U4779 (N_4779,N_3912,N_3283);
and U4780 (N_4780,N_3290,N_3887);
xnor U4781 (N_4781,N_3915,N_3443);
and U4782 (N_4782,N_3523,N_3568);
and U4783 (N_4783,N_3199,N_3423);
nor U4784 (N_4784,N_3622,N_3243);
or U4785 (N_4785,N_3077,N_3134);
nand U4786 (N_4786,N_3817,N_3172);
or U4787 (N_4787,N_3761,N_3571);
or U4788 (N_4788,N_3819,N_3728);
or U4789 (N_4789,N_3076,N_3289);
and U4790 (N_4790,N_3191,N_3613);
nand U4791 (N_4791,N_3431,N_3642);
nor U4792 (N_4792,N_3304,N_3171);
xnor U4793 (N_4793,N_3996,N_3999);
nor U4794 (N_4794,N_3450,N_3278);
or U4795 (N_4795,N_3490,N_3958);
nand U4796 (N_4796,N_3432,N_3776);
nor U4797 (N_4797,N_3186,N_3379);
nand U4798 (N_4798,N_3872,N_3623);
nand U4799 (N_4799,N_3191,N_3882);
and U4800 (N_4800,N_3880,N_3672);
nand U4801 (N_4801,N_3867,N_3333);
and U4802 (N_4802,N_3108,N_3460);
xnor U4803 (N_4803,N_3108,N_3791);
nand U4804 (N_4804,N_3849,N_3431);
and U4805 (N_4805,N_3389,N_3432);
or U4806 (N_4806,N_3793,N_3609);
nand U4807 (N_4807,N_3525,N_3084);
and U4808 (N_4808,N_3665,N_3107);
or U4809 (N_4809,N_3061,N_3190);
or U4810 (N_4810,N_3313,N_3154);
and U4811 (N_4811,N_3976,N_3684);
nor U4812 (N_4812,N_3130,N_3937);
or U4813 (N_4813,N_3539,N_3548);
nor U4814 (N_4814,N_3989,N_3231);
nand U4815 (N_4815,N_3046,N_3724);
nand U4816 (N_4816,N_3311,N_3113);
nand U4817 (N_4817,N_3381,N_3602);
and U4818 (N_4818,N_3214,N_3078);
or U4819 (N_4819,N_3954,N_3821);
nand U4820 (N_4820,N_3993,N_3529);
nor U4821 (N_4821,N_3648,N_3959);
nand U4822 (N_4822,N_3770,N_3869);
nor U4823 (N_4823,N_3184,N_3504);
nor U4824 (N_4824,N_3145,N_3483);
or U4825 (N_4825,N_3192,N_3644);
and U4826 (N_4826,N_3494,N_3367);
and U4827 (N_4827,N_3361,N_3797);
nor U4828 (N_4828,N_3945,N_3546);
and U4829 (N_4829,N_3681,N_3877);
and U4830 (N_4830,N_3607,N_3934);
and U4831 (N_4831,N_3457,N_3182);
or U4832 (N_4832,N_3430,N_3482);
nand U4833 (N_4833,N_3923,N_3938);
and U4834 (N_4834,N_3923,N_3215);
or U4835 (N_4835,N_3936,N_3501);
or U4836 (N_4836,N_3446,N_3073);
or U4837 (N_4837,N_3811,N_3594);
nor U4838 (N_4838,N_3465,N_3724);
nor U4839 (N_4839,N_3728,N_3317);
nor U4840 (N_4840,N_3382,N_3483);
nand U4841 (N_4841,N_3230,N_3980);
and U4842 (N_4842,N_3337,N_3589);
nor U4843 (N_4843,N_3545,N_3134);
nor U4844 (N_4844,N_3328,N_3493);
nand U4845 (N_4845,N_3988,N_3795);
nor U4846 (N_4846,N_3226,N_3085);
nor U4847 (N_4847,N_3233,N_3862);
nand U4848 (N_4848,N_3122,N_3222);
nand U4849 (N_4849,N_3717,N_3971);
or U4850 (N_4850,N_3735,N_3257);
and U4851 (N_4851,N_3460,N_3962);
or U4852 (N_4852,N_3109,N_3272);
nand U4853 (N_4853,N_3475,N_3346);
nand U4854 (N_4854,N_3321,N_3372);
nor U4855 (N_4855,N_3327,N_3853);
or U4856 (N_4856,N_3504,N_3832);
nor U4857 (N_4857,N_3213,N_3312);
or U4858 (N_4858,N_3384,N_3443);
and U4859 (N_4859,N_3259,N_3878);
or U4860 (N_4860,N_3639,N_3453);
nor U4861 (N_4861,N_3774,N_3097);
or U4862 (N_4862,N_3402,N_3462);
and U4863 (N_4863,N_3828,N_3792);
nand U4864 (N_4864,N_3571,N_3528);
nor U4865 (N_4865,N_3280,N_3054);
nor U4866 (N_4866,N_3973,N_3781);
or U4867 (N_4867,N_3418,N_3916);
nand U4868 (N_4868,N_3536,N_3403);
or U4869 (N_4869,N_3495,N_3233);
nand U4870 (N_4870,N_3235,N_3244);
nand U4871 (N_4871,N_3948,N_3127);
nand U4872 (N_4872,N_3772,N_3844);
and U4873 (N_4873,N_3526,N_3576);
or U4874 (N_4874,N_3589,N_3043);
nand U4875 (N_4875,N_3744,N_3808);
and U4876 (N_4876,N_3202,N_3063);
nand U4877 (N_4877,N_3008,N_3591);
or U4878 (N_4878,N_3096,N_3033);
and U4879 (N_4879,N_3124,N_3836);
or U4880 (N_4880,N_3393,N_3789);
and U4881 (N_4881,N_3023,N_3597);
and U4882 (N_4882,N_3434,N_3336);
or U4883 (N_4883,N_3690,N_3351);
or U4884 (N_4884,N_3932,N_3547);
or U4885 (N_4885,N_3334,N_3406);
and U4886 (N_4886,N_3028,N_3892);
nor U4887 (N_4887,N_3482,N_3592);
or U4888 (N_4888,N_3265,N_3263);
nand U4889 (N_4889,N_3514,N_3993);
nand U4890 (N_4890,N_3014,N_3594);
or U4891 (N_4891,N_3713,N_3891);
and U4892 (N_4892,N_3297,N_3779);
or U4893 (N_4893,N_3582,N_3093);
nand U4894 (N_4894,N_3960,N_3292);
or U4895 (N_4895,N_3725,N_3261);
and U4896 (N_4896,N_3172,N_3088);
nand U4897 (N_4897,N_3765,N_3627);
and U4898 (N_4898,N_3024,N_3359);
nand U4899 (N_4899,N_3108,N_3429);
and U4900 (N_4900,N_3734,N_3615);
or U4901 (N_4901,N_3686,N_3962);
nand U4902 (N_4902,N_3400,N_3556);
nand U4903 (N_4903,N_3323,N_3933);
and U4904 (N_4904,N_3712,N_3221);
nand U4905 (N_4905,N_3853,N_3229);
nor U4906 (N_4906,N_3053,N_3980);
or U4907 (N_4907,N_3461,N_3651);
or U4908 (N_4908,N_3346,N_3702);
and U4909 (N_4909,N_3396,N_3757);
or U4910 (N_4910,N_3006,N_3756);
nand U4911 (N_4911,N_3528,N_3568);
nand U4912 (N_4912,N_3674,N_3695);
nand U4913 (N_4913,N_3592,N_3823);
nand U4914 (N_4914,N_3191,N_3654);
nand U4915 (N_4915,N_3527,N_3555);
nor U4916 (N_4916,N_3061,N_3140);
or U4917 (N_4917,N_3392,N_3263);
and U4918 (N_4918,N_3236,N_3743);
or U4919 (N_4919,N_3462,N_3827);
and U4920 (N_4920,N_3419,N_3566);
nor U4921 (N_4921,N_3319,N_3279);
and U4922 (N_4922,N_3096,N_3679);
nand U4923 (N_4923,N_3135,N_3683);
or U4924 (N_4924,N_3243,N_3123);
and U4925 (N_4925,N_3431,N_3181);
nor U4926 (N_4926,N_3876,N_3128);
and U4927 (N_4927,N_3882,N_3198);
and U4928 (N_4928,N_3426,N_3583);
nor U4929 (N_4929,N_3979,N_3864);
or U4930 (N_4930,N_3972,N_3438);
nor U4931 (N_4931,N_3789,N_3139);
nand U4932 (N_4932,N_3825,N_3531);
nand U4933 (N_4933,N_3920,N_3899);
nor U4934 (N_4934,N_3279,N_3858);
and U4935 (N_4935,N_3069,N_3356);
nor U4936 (N_4936,N_3922,N_3865);
nand U4937 (N_4937,N_3680,N_3962);
nand U4938 (N_4938,N_3997,N_3790);
and U4939 (N_4939,N_3967,N_3301);
nand U4940 (N_4940,N_3207,N_3210);
nor U4941 (N_4941,N_3940,N_3205);
nor U4942 (N_4942,N_3276,N_3694);
and U4943 (N_4943,N_3215,N_3889);
nor U4944 (N_4944,N_3615,N_3287);
and U4945 (N_4945,N_3888,N_3765);
or U4946 (N_4946,N_3451,N_3999);
nand U4947 (N_4947,N_3589,N_3995);
nand U4948 (N_4948,N_3514,N_3711);
and U4949 (N_4949,N_3855,N_3823);
nor U4950 (N_4950,N_3435,N_3994);
and U4951 (N_4951,N_3777,N_3525);
nor U4952 (N_4952,N_3311,N_3310);
nand U4953 (N_4953,N_3898,N_3129);
and U4954 (N_4954,N_3291,N_3887);
nor U4955 (N_4955,N_3223,N_3243);
nor U4956 (N_4956,N_3302,N_3841);
nor U4957 (N_4957,N_3499,N_3580);
and U4958 (N_4958,N_3002,N_3269);
nor U4959 (N_4959,N_3177,N_3915);
or U4960 (N_4960,N_3661,N_3028);
nor U4961 (N_4961,N_3040,N_3353);
nand U4962 (N_4962,N_3266,N_3519);
nor U4963 (N_4963,N_3865,N_3076);
and U4964 (N_4964,N_3927,N_3420);
nand U4965 (N_4965,N_3036,N_3064);
and U4966 (N_4966,N_3038,N_3194);
nor U4967 (N_4967,N_3393,N_3804);
xor U4968 (N_4968,N_3047,N_3210);
nand U4969 (N_4969,N_3636,N_3114);
nor U4970 (N_4970,N_3812,N_3497);
and U4971 (N_4971,N_3049,N_3708);
or U4972 (N_4972,N_3350,N_3103);
nand U4973 (N_4973,N_3276,N_3545);
and U4974 (N_4974,N_3532,N_3133);
nor U4975 (N_4975,N_3722,N_3457);
nand U4976 (N_4976,N_3561,N_3455);
nor U4977 (N_4977,N_3797,N_3431);
or U4978 (N_4978,N_3619,N_3366);
nor U4979 (N_4979,N_3092,N_3875);
and U4980 (N_4980,N_3998,N_3765);
nand U4981 (N_4981,N_3655,N_3148);
nor U4982 (N_4982,N_3521,N_3202);
nor U4983 (N_4983,N_3486,N_3340);
nand U4984 (N_4984,N_3192,N_3797);
nor U4985 (N_4985,N_3060,N_3120);
nor U4986 (N_4986,N_3559,N_3781);
or U4987 (N_4987,N_3787,N_3633);
nor U4988 (N_4988,N_3877,N_3204);
and U4989 (N_4989,N_3405,N_3476);
nand U4990 (N_4990,N_3153,N_3593);
or U4991 (N_4991,N_3215,N_3532);
nor U4992 (N_4992,N_3037,N_3440);
and U4993 (N_4993,N_3903,N_3589);
nor U4994 (N_4994,N_3407,N_3331);
or U4995 (N_4995,N_3685,N_3441);
nor U4996 (N_4996,N_3184,N_3625);
or U4997 (N_4997,N_3408,N_3706);
nand U4998 (N_4998,N_3341,N_3804);
or U4999 (N_4999,N_3648,N_3301);
or UO_0 (O_0,N_4446,N_4621);
nor UO_1 (O_1,N_4116,N_4338);
nor UO_2 (O_2,N_4540,N_4155);
nand UO_3 (O_3,N_4662,N_4686);
nand UO_4 (O_4,N_4997,N_4164);
and UO_5 (O_5,N_4249,N_4421);
and UO_6 (O_6,N_4439,N_4141);
or UO_7 (O_7,N_4576,N_4587);
or UO_8 (O_8,N_4330,N_4352);
or UO_9 (O_9,N_4056,N_4749);
nand UO_10 (O_10,N_4893,N_4429);
and UO_11 (O_11,N_4567,N_4925);
nor UO_12 (O_12,N_4591,N_4565);
or UO_13 (O_13,N_4039,N_4530);
nand UO_14 (O_14,N_4709,N_4379);
or UO_15 (O_15,N_4940,N_4644);
and UO_16 (O_16,N_4852,N_4057);
or UO_17 (O_17,N_4428,N_4127);
nand UO_18 (O_18,N_4906,N_4669);
or UO_19 (O_19,N_4776,N_4802);
or UO_20 (O_20,N_4745,N_4696);
nand UO_21 (O_21,N_4605,N_4501);
and UO_22 (O_22,N_4457,N_4792);
nor UO_23 (O_23,N_4831,N_4939);
nor UO_24 (O_24,N_4528,N_4158);
nand UO_25 (O_25,N_4729,N_4445);
nor UO_26 (O_26,N_4606,N_4740);
nand UO_27 (O_27,N_4685,N_4920);
or UO_28 (O_28,N_4645,N_4904);
nand UO_29 (O_29,N_4130,N_4609);
nand UO_30 (O_30,N_4803,N_4364);
and UO_31 (O_31,N_4118,N_4044);
and UO_32 (O_32,N_4007,N_4458);
nor UO_33 (O_33,N_4666,N_4817);
and UO_34 (O_34,N_4835,N_4734);
and UO_35 (O_35,N_4225,N_4550);
nand UO_36 (O_36,N_4449,N_4974);
nand UO_37 (O_37,N_4062,N_4703);
or UO_38 (O_38,N_4423,N_4728);
and UO_39 (O_39,N_4046,N_4913);
and UO_40 (O_40,N_4403,N_4089);
nand UO_41 (O_41,N_4038,N_4579);
and UO_42 (O_42,N_4244,N_4406);
or UO_43 (O_43,N_4190,N_4950);
or UO_44 (O_44,N_4508,N_4498);
nand UO_45 (O_45,N_4689,N_4743);
nor UO_46 (O_46,N_4842,N_4131);
or UO_47 (O_47,N_4861,N_4582);
and UO_48 (O_48,N_4369,N_4034);
nand UO_49 (O_49,N_4425,N_4959);
nor UO_50 (O_50,N_4409,N_4443);
nor UO_51 (O_51,N_4794,N_4286);
nor UO_52 (O_52,N_4004,N_4500);
nand UO_53 (O_53,N_4397,N_4161);
nor UO_54 (O_54,N_4739,N_4642);
or UO_55 (O_55,N_4777,N_4005);
and UO_56 (O_56,N_4494,N_4477);
nor UO_57 (O_57,N_4836,N_4226);
nor UO_58 (O_58,N_4882,N_4807);
and UO_59 (O_59,N_4150,N_4117);
nor UO_60 (O_60,N_4614,N_4144);
and UO_61 (O_61,N_4979,N_4393);
and UO_62 (O_62,N_4073,N_4931);
and UO_63 (O_63,N_4377,N_4595);
nor UO_64 (O_64,N_4557,N_4600);
or UO_65 (O_65,N_4754,N_4868);
nand UO_66 (O_66,N_4020,N_4140);
nand UO_67 (O_67,N_4715,N_4091);
nor UO_68 (O_68,N_4598,N_4748);
or UO_69 (O_69,N_4726,N_4744);
or UO_70 (O_70,N_4334,N_4783);
nand UO_71 (O_71,N_4195,N_4465);
and UO_72 (O_72,N_4980,N_4548);
and UO_73 (O_73,N_4264,N_4752);
or UO_74 (O_74,N_4160,N_4615);
and UO_75 (O_75,N_4751,N_4525);
and UO_76 (O_76,N_4450,N_4771);
nand UO_77 (O_77,N_4681,N_4536);
and UO_78 (O_78,N_4658,N_4217);
and UO_79 (O_79,N_4901,N_4510);
and UO_80 (O_80,N_4516,N_4961);
and UO_81 (O_81,N_4848,N_4215);
or UO_82 (O_82,N_4832,N_4098);
nor UO_83 (O_83,N_4176,N_4378);
nand UO_84 (O_84,N_4203,N_4755);
and UO_85 (O_85,N_4736,N_4635);
and UO_86 (O_86,N_4052,N_4341);
nor UO_87 (O_87,N_4630,N_4623);
and UO_88 (O_88,N_4616,N_4361);
nand UO_89 (O_89,N_4907,N_4679);
nand UO_90 (O_90,N_4461,N_4927);
nand UO_91 (O_91,N_4275,N_4420);
or UO_92 (O_92,N_4829,N_4012);
nor UO_93 (O_93,N_4732,N_4181);
nor UO_94 (O_94,N_4174,N_4143);
nor UO_95 (O_95,N_4408,N_4710);
xor UO_96 (O_96,N_4018,N_4188);
or UO_97 (O_97,N_4357,N_4462);
nand UO_98 (O_98,N_4655,N_4256);
nor UO_99 (O_99,N_4723,N_4555);
or UO_100 (O_100,N_4311,N_4358);
and UO_101 (O_101,N_4231,N_4796);
nand UO_102 (O_102,N_4934,N_4197);
nor UO_103 (O_103,N_4660,N_4454);
nor UO_104 (O_104,N_4452,N_4339);
or UO_105 (O_105,N_4066,N_4845);
nand UO_106 (O_106,N_4324,N_4208);
and UO_107 (O_107,N_4284,N_4086);
nand UO_108 (O_108,N_4879,N_4192);
nand UO_109 (O_109,N_4973,N_4093);
or UO_110 (O_110,N_4948,N_4105);
nor UO_111 (O_111,N_4871,N_4430);
and UO_112 (O_112,N_4031,N_4546);
and UO_113 (O_113,N_4781,N_4575);
and UO_114 (O_114,N_4810,N_4825);
or UO_115 (O_115,N_4714,N_4663);
or UO_116 (O_116,N_4884,N_4800);
and UO_117 (O_117,N_4684,N_4075);
nor UO_118 (O_118,N_4992,N_4081);
nor UO_119 (O_119,N_4488,N_4382);
nor UO_120 (O_120,N_4148,N_4756);
or UO_121 (O_121,N_4386,N_4270);
nor UO_122 (O_122,N_4125,N_4727);
and UO_123 (O_123,N_4482,N_4337);
nand UO_124 (O_124,N_4100,N_4307);
nand UO_125 (O_125,N_4444,N_4077);
or UO_126 (O_126,N_4724,N_4889);
and UO_127 (O_127,N_4479,N_4050);
or UO_128 (O_128,N_4849,N_4881);
nand UO_129 (O_129,N_4115,N_4157);
or UO_130 (O_130,N_4599,N_4122);
nor UO_131 (O_131,N_4613,N_4064);
nand UO_132 (O_132,N_4700,N_4344);
or UO_133 (O_133,N_4798,N_4787);
and UO_134 (O_134,N_4985,N_4129);
nor UO_135 (O_135,N_4702,N_4293);
or UO_136 (O_136,N_4704,N_4819);
and UO_137 (O_137,N_4198,N_4111);
or UO_138 (O_138,N_4618,N_4890);
and UO_139 (O_139,N_4410,N_4022);
and UO_140 (O_140,N_4041,N_4232);
or UO_141 (O_141,N_4123,N_4059);
and UO_142 (O_142,N_4413,N_4417);
nand UO_143 (O_143,N_4559,N_4163);
or UO_144 (O_144,N_4806,N_4513);
and UO_145 (O_145,N_4366,N_4023);
nand UO_146 (O_146,N_4469,N_4265);
and UO_147 (O_147,N_4492,N_4603);
nor UO_148 (O_148,N_4253,N_4763);
and UO_149 (O_149,N_4389,N_4201);
and UO_150 (O_150,N_4731,N_4717);
nand UO_151 (O_151,N_4705,N_4333);
and UO_152 (O_152,N_4189,N_4987);
and UO_153 (O_153,N_4813,N_4643);
and UO_154 (O_154,N_4107,N_4965);
or UO_155 (O_155,N_4321,N_4119);
and UO_156 (O_156,N_4486,N_4251);
and UO_157 (O_157,N_4580,N_4675);
nor UO_158 (O_158,N_4894,N_4986);
nor UO_159 (O_159,N_4902,N_4432);
or UO_160 (O_160,N_4024,N_4531);
nand UO_161 (O_161,N_4308,N_4033);
and UO_162 (O_162,N_4362,N_4011);
nor UO_163 (O_163,N_4495,N_4407);
nand UO_164 (O_164,N_4697,N_4526);
nor UO_165 (O_165,N_4360,N_4995);
or UO_166 (O_166,N_4693,N_4607);
or UO_167 (O_167,N_4891,N_4095);
and UO_168 (O_168,N_4147,N_4078);
and UO_169 (O_169,N_4677,N_4317);
or UO_170 (O_170,N_4213,N_4636);
nor UO_171 (O_171,N_4481,N_4910);
and UO_172 (O_172,N_4416,N_4601);
nor UO_173 (O_173,N_4941,N_4560);
or UO_174 (O_174,N_4242,N_4657);
nor UO_175 (O_175,N_4937,N_4730);
nand UO_176 (O_176,N_4678,N_4053);
nand UO_177 (O_177,N_4017,N_4110);
and UO_178 (O_178,N_4822,N_4072);
nand UO_179 (O_179,N_4517,N_4000);
nand UO_180 (O_180,N_4099,N_4993);
and UO_181 (O_181,N_4653,N_4047);
xor UO_182 (O_182,N_4563,N_4532);
and UO_183 (O_183,N_4071,N_4074);
nand UO_184 (O_184,N_4302,N_4343);
nand UO_185 (O_185,N_4399,N_4065);
nor UO_186 (O_186,N_4674,N_4272);
and UO_187 (O_187,N_4826,N_4789);
nand UO_188 (O_188,N_4040,N_4594);
xor UO_189 (O_189,N_4422,N_4448);
and UO_190 (O_190,N_4772,N_4656);
or UO_191 (O_191,N_4058,N_4999);
or UO_192 (O_192,N_4647,N_4261);
nand UO_193 (O_193,N_4692,N_4294);
or UO_194 (O_194,N_4552,N_4042);
nand UO_195 (O_195,N_4566,N_4619);
nor UO_196 (O_196,N_4841,N_4298);
or UO_197 (O_197,N_4903,N_4460);
or UO_198 (O_198,N_4808,N_4875);
or UO_199 (O_199,N_4196,N_4026);
nor UO_200 (O_200,N_4759,N_4648);
nor UO_201 (O_201,N_4924,N_4476);
and UO_202 (O_202,N_4069,N_4778);
nand UO_203 (O_203,N_4610,N_4112);
and UO_204 (O_204,N_4350,N_4390);
and UO_205 (O_205,N_4035,N_4870);
nor UO_206 (O_206,N_4394,N_4912);
nand UO_207 (O_207,N_4336,N_4021);
and UO_208 (O_208,N_4082,N_4706);
nand UO_209 (O_209,N_4451,N_4793);
nand UO_210 (O_210,N_4142,N_4843);
or UO_211 (O_211,N_4132,N_4243);
or UO_212 (O_212,N_4942,N_4279);
nand UO_213 (O_213,N_4049,N_4167);
nand UO_214 (O_214,N_4897,N_4782);
nand UO_215 (O_215,N_4888,N_4541);
or UO_216 (O_216,N_4914,N_4694);
or UO_217 (O_217,N_4542,N_4585);
and UO_218 (O_218,N_4911,N_4551);
and UO_219 (O_219,N_4101,N_4162);
nand UO_220 (O_220,N_4984,N_4856);
and UO_221 (O_221,N_4471,N_4316);
nand UO_222 (O_222,N_4654,N_4951);
or UO_223 (O_223,N_4774,N_4166);
and UO_224 (O_224,N_4179,N_4983);
or UO_225 (O_225,N_4175,N_4876);
nand UO_226 (O_226,N_4263,N_4757);
or UO_227 (O_227,N_4722,N_4593);
or UO_228 (O_228,N_4988,N_4060);
and UO_229 (O_229,N_4627,N_4529);
and UO_230 (O_230,N_4949,N_4400);
or UO_231 (O_231,N_4079,N_4652);
or UO_232 (O_232,N_4972,N_4106);
and UO_233 (O_233,N_4741,N_4797);
and UO_234 (O_234,N_4153,N_4313);
nand UO_235 (O_235,N_4823,N_4083);
nand UO_236 (O_236,N_4886,N_4260);
nand UO_237 (O_237,N_4246,N_4649);
or UO_238 (O_238,N_4391,N_4345);
and UO_239 (O_239,N_4571,N_4045);
or UO_240 (O_240,N_4833,N_4535);
or UO_241 (O_241,N_4365,N_4511);
nor UO_242 (O_242,N_4312,N_4145);
or UO_243 (O_243,N_4447,N_4222);
nand UO_244 (O_244,N_4464,N_4638);
nand UO_245 (O_245,N_4964,N_4561);
nand UO_246 (O_246,N_4229,N_4837);
nor UO_247 (O_247,N_4608,N_4314);
nor UO_248 (O_248,N_4114,N_4712);
nand UO_249 (O_249,N_4699,N_4947);
nor UO_250 (O_250,N_4154,N_4281);
nand UO_251 (O_251,N_4151,N_4385);
and UO_252 (O_252,N_4507,N_4388);
nor UO_253 (O_253,N_4853,N_4664);
nor UO_254 (O_254,N_4297,N_4804);
xor UO_255 (O_255,N_4258,N_4758);
nor UO_256 (O_256,N_4880,N_4342);
and UO_257 (O_257,N_4520,N_4885);
or UO_258 (O_258,N_4493,N_4269);
nand UO_259 (O_259,N_4067,N_4381);
and UO_260 (O_260,N_4646,N_4172);
and UO_261 (O_261,N_4440,N_4780);
or UO_262 (O_262,N_4918,N_4183);
or UO_263 (O_263,N_4892,N_4866);
nor UO_264 (O_264,N_4376,N_4383);
or UO_265 (O_265,N_4718,N_4919);
and UO_266 (O_266,N_4199,N_4568);
or UO_267 (O_267,N_4641,N_4087);
or UO_268 (O_268,N_4746,N_4356);
and UO_269 (O_269,N_4205,N_4267);
and UO_270 (O_270,N_4953,N_4522);
nor UO_271 (O_271,N_4467,N_4969);
and UO_272 (O_272,N_4773,N_4682);
nand UO_273 (O_273,N_4504,N_4725);
nor UO_274 (O_274,N_4887,N_4765);
xnor UO_275 (O_275,N_4926,N_4801);
or UO_276 (O_276,N_4135,N_4489);
nand UO_277 (O_277,N_4236,N_4665);
nand UO_278 (O_278,N_4917,N_4288);
nor UO_279 (O_279,N_4475,N_4761);
nand UO_280 (O_280,N_4255,N_4588);
nand UO_281 (O_281,N_4013,N_4335);
or UO_282 (O_282,N_4878,N_4304);
or UO_283 (O_283,N_4431,N_4946);
nand UO_284 (O_284,N_4436,N_4938);
and UO_285 (O_285,N_4325,N_4977);
nor UO_286 (O_286,N_4786,N_4570);
nand UO_287 (O_287,N_4036,N_4496);
or UO_288 (O_288,N_4137,N_4412);
nand UO_289 (O_289,N_4204,N_4340);
or UO_290 (O_290,N_4503,N_4327);
or UO_291 (O_291,N_4349,N_4967);
and UO_292 (O_292,N_4289,N_4028);
and UO_293 (O_293,N_4241,N_4633);
and UO_294 (O_294,N_4016,N_4572);
nor UO_295 (O_295,N_4943,N_4387);
and UO_296 (O_296,N_4224,N_4667);
nand UO_297 (O_297,N_4770,N_4695);
nor UO_298 (O_298,N_4126,N_4976);
and UO_299 (O_299,N_4207,N_4309);
and UO_300 (O_300,N_4867,N_4380);
or UO_301 (O_301,N_4586,N_4480);
and UO_302 (O_302,N_4830,N_4003);
and UO_303 (O_303,N_4634,N_4472);
nor UO_304 (O_304,N_4068,N_4219);
nand UO_305 (O_305,N_4355,N_4367);
nand UO_306 (O_306,N_4612,N_4900);
xor UO_307 (O_307,N_4030,N_4169);
or UO_308 (O_308,N_4002,N_4405);
and UO_309 (O_309,N_4374,N_4538);
nor UO_310 (O_310,N_4485,N_4945);
nor UO_311 (O_311,N_4076,N_4001);
and UO_312 (O_312,N_4146,N_4805);
or UO_313 (O_313,N_4839,N_4063);
nor UO_314 (O_314,N_4814,N_4159);
nor UO_315 (O_315,N_4418,N_4274);
nor UO_316 (O_316,N_4930,N_4860);
nor UO_317 (O_317,N_4533,N_4171);
nand UO_318 (O_318,N_4438,N_4015);
nand UO_319 (O_319,N_4055,N_4096);
or UO_320 (O_320,N_4982,N_4518);
or UO_321 (O_321,N_4968,N_4899);
nor UO_322 (O_322,N_4173,N_4483);
nor UO_323 (O_323,N_4519,N_4212);
nand UO_324 (O_324,N_4515,N_4434);
nand UO_325 (O_325,N_4426,N_4323);
or UO_326 (O_326,N_4922,N_4872);
nand UO_327 (O_327,N_4760,N_4221);
or UO_328 (O_328,N_4459,N_4617);
nand UO_329 (O_329,N_4564,N_4254);
nand UO_330 (O_330,N_4611,N_4240);
and UO_331 (O_331,N_4456,N_4916);
and UO_332 (O_332,N_4818,N_4955);
xor UO_333 (O_333,N_4602,N_4553);
nand UO_334 (O_334,N_4296,N_4354);
and UO_335 (O_335,N_4401,N_4248);
nor UO_336 (O_336,N_4547,N_4283);
nand UO_337 (O_337,N_4840,N_4441);
nor UO_338 (O_338,N_4750,N_4628);
nand UO_339 (O_339,N_4855,N_4989);
nor UO_340 (O_340,N_4534,N_4120);
nor UO_341 (O_341,N_4487,N_4103);
nand UO_342 (O_342,N_4252,N_4184);
nor UO_343 (O_343,N_4250,N_4008);
or UO_344 (O_344,N_4187,N_4775);
nand UO_345 (O_345,N_4211,N_4978);
nand UO_346 (O_346,N_4562,N_4716);
nand UO_347 (O_347,N_4210,N_4202);
or UO_348 (O_348,N_4554,N_4168);
nor UO_349 (O_349,N_4929,N_4549);
nand UO_350 (O_350,N_4411,N_4747);
and UO_351 (O_351,N_4398,N_4811);
or UO_352 (O_352,N_4453,N_4276);
and UO_353 (O_353,N_4220,N_4956);
nand UO_354 (O_354,N_4239,N_4990);
or UO_355 (O_355,N_4303,N_4733);
or UO_356 (O_356,N_4414,N_4719);
and UO_357 (O_357,N_4372,N_4766);
nor UO_358 (O_358,N_4185,N_4680);
and UO_359 (O_359,N_4996,N_4315);
nor UO_360 (O_360,N_4514,N_4795);
and UO_361 (O_361,N_4944,N_4788);
nand UO_362 (O_362,N_4051,N_4102);
and UO_363 (O_363,N_4720,N_4402);
or UO_364 (O_364,N_4847,N_4424);
nand UO_365 (O_365,N_4006,N_4597);
and UO_366 (O_366,N_4824,N_4178);
nor UO_367 (O_367,N_4857,N_4259);
nand UO_368 (O_368,N_4673,N_4152);
xnor UO_369 (O_369,N_4933,N_4359);
nor UO_370 (O_370,N_4524,N_4713);
and UO_371 (O_371,N_4701,N_4027);
and UO_372 (O_372,N_4604,N_4156);
and UO_373 (O_373,N_4351,N_4404);
or UO_374 (O_374,N_4865,N_4668);
and UO_375 (O_375,N_4962,N_4468);
and UO_376 (O_376,N_4375,N_4133);
or UO_377 (O_377,N_4874,N_4898);
nand UO_378 (O_378,N_4622,N_4182);
or UO_379 (O_379,N_4257,N_4273);
and UO_380 (O_380,N_4139,N_4373);
nor UO_381 (O_381,N_4767,N_4009);
nand UO_382 (O_382,N_4478,N_4828);
and UO_383 (O_383,N_4671,N_4558);
nor UO_384 (O_384,N_4932,N_4280);
or UO_385 (O_385,N_4991,N_4512);
or UO_386 (O_386,N_4584,N_4543);
nor UO_387 (O_387,N_4165,N_4909);
and UO_388 (O_388,N_4735,N_4966);
nand UO_389 (O_389,N_4683,N_4295);
nand UO_390 (O_390,N_4556,N_4523);
or UO_391 (O_391,N_4869,N_4592);
or UO_392 (O_392,N_4278,N_4659);
nand UO_393 (O_393,N_4676,N_4640);
or UO_394 (O_394,N_4484,N_4812);
nand UO_395 (O_395,N_4180,N_4491);
nor UO_396 (O_396,N_4862,N_4437);
nand UO_397 (O_397,N_4905,N_4569);
and UO_398 (O_398,N_4539,N_4816);
or UO_399 (O_399,N_4191,N_4502);
nor UO_400 (O_400,N_4858,N_4200);
and UO_401 (O_401,N_4277,N_4234);
or UO_402 (O_402,N_4300,N_4670);
and UO_403 (O_403,N_4799,N_4509);
nand UO_404 (O_404,N_4707,N_4291);
nor UO_405 (O_405,N_4844,N_4209);
and UO_406 (O_406,N_4639,N_4194);
nand UO_407 (O_407,N_4753,N_4820);
and UO_408 (O_408,N_4328,N_4473);
or UO_409 (O_409,N_4084,N_4353);
or UO_410 (O_410,N_4080,N_4688);
xnor UO_411 (O_411,N_4923,N_4791);
nand UO_412 (O_412,N_4010,N_4994);
and UO_413 (O_413,N_4223,N_4505);
nor UO_414 (O_414,N_4287,N_4237);
and UO_415 (O_415,N_4415,N_4632);
and UO_416 (O_416,N_4238,N_4227);
nor UO_417 (O_417,N_4474,N_4092);
nand UO_418 (O_418,N_4850,N_4690);
nand UO_419 (O_419,N_4691,N_4113);
nor UO_420 (O_420,N_4768,N_4625);
nand UO_421 (O_421,N_4497,N_4319);
and UO_422 (O_422,N_4711,N_4433);
nor UO_423 (O_423,N_4214,N_4245);
nand UO_424 (O_424,N_4136,N_4935);
or UO_425 (O_425,N_4014,N_4032);
nand UO_426 (O_426,N_4463,N_4370);
or UO_427 (O_427,N_4998,N_4466);
xor UO_428 (O_428,N_4624,N_4698);
or UO_429 (O_429,N_4435,N_4419);
and UO_430 (O_430,N_4838,N_4672);
nand UO_431 (O_431,N_4455,N_4331);
or UO_432 (O_432,N_4233,N_4368);
and UO_433 (O_433,N_4170,N_4544);
nor UO_434 (O_434,N_4128,N_4427);
nand UO_435 (O_435,N_4521,N_4651);
nor UO_436 (O_436,N_4915,N_4310);
and UO_437 (O_437,N_4661,N_4506);
nor UO_438 (O_438,N_4851,N_4025);
nand UO_439 (O_439,N_4769,N_4442);
or UO_440 (O_440,N_4596,N_4545);
and UO_441 (O_441,N_4527,N_4177);
and UO_442 (O_442,N_4883,N_4193);
or UO_443 (O_443,N_4864,N_4785);
or UO_444 (O_444,N_4371,N_4859);
nor UO_445 (O_445,N_4762,N_4346);
or UO_446 (O_446,N_4846,N_4908);
nand UO_447 (O_447,N_4764,N_4981);
and UO_448 (O_448,N_4301,N_4957);
and UO_449 (O_449,N_4285,N_4332);
nor UO_450 (O_450,N_4054,N_4088);
nor UO_451 (O_451,N_4206,N_4737);
nand UO_452 (O_452,N_4895,N_4395);
and UO_453 (O_453,N_4305,N_4186);
and UO_454 (O_454,N_4363,N_4896);
nand UO_455 (O_455,N_4104,N_4952);
or UO_456 (O_456,N_4809,N_4230);
nor UO_457 (O_457,N_4970,N_4048);
nor UO_458 (O_458,N_4134,N_4928);
nand UO_459 (O_459,N_4626,N_4218);
and UO_460 (O_460,N_4590,N_4090);
nor UO_461 (O_461,N_4499,N_4790);
nor UO_462 (O_462,N_4124,N_4348);
nor UO_463 (O_463,N_4687,N_4268);
or UO_464 (O_464,N_4854,N_4779);
or UO_465 (O_465,N_4149,N_4347);
nor UO_466 (O_466,N_4960,N_4708);
or UO_467 (O_467,N_4070,N_4085);
and UO_468 (O_468,N_4108,N_4742);
nor UO_469 (O_469,N_4537,N_4581);
and UO_470 (O_470,N_4589,N_4320);
nand UO_471 (O_471,N_4299,N_4019);
or UO_472 (O_472,N_4721,N_4877);
and UO_473 (O_473,N_4228,N_4247);
or UO_474 (O_474,N_4963,N_4827);
nand UO_475 (O_475,N_4784,N_4834);
nand UO_476 (O_476,N_4873,N_4631);
nor UO_477 (O_477,N_4863,N_4216);
or UO_478 (O_478,N_4282,N_4384);
nor UO_479 (O_479,N_4292,N_4094);
nor UO_480 (O_480,N_4573,N_4971);
or UO_481 (O_481,N_4577,N_4821);
nand UO_482 (O_482,N_4306,N_4235);
nand UO_483 (O_483,N_4470,N_4574);
and UO_484 (O_484,N_4392,N_4138);
and UO_485 (O_485,N_4266,N_4650);
or UO_486 (O_486,N_4322,N_4975);
nand UO_487 (O_487,N_4109,N_4936);
and UO_488 (O_488,N_4578,N_4954);
and UO_489 (O_489,N_4262,N_4583);
nand UO_490 (O_490,N_4815,N_4329);
and UO_491 (O_491,N_4029,N_4061);
nor UO_492 (O_492,N_4121,N_4490);
or UO_493 (O_493,N_4620,N_4043);
and UO_494 (O_494,N_4738,N_4396);
nand UO_495 (O_495,N_4271,N_4318);
or UO_496 (O_496,N_4037,N_4326);
and UO_497 (O_497,N_4097,N_4290);
nor UO_498 (O_498,N_4921,N_4637);
nand UO_499 (O_499,N_4958,N_4629);
or UO_500 (O_500,N_4712,N_4321);
or UO_501 (O_501,N_4415,N_4590);
nor UO_502 (O_502,N_4312,N_4028);
nor UO_503 (O_503,N_4799,N_4925);
and UO_504 (O_504,N_4676,N_4042);
and UO_505 (O_505,N_4194,N_4924);
nand UO_506 (O_506,N_4696,N_4760);
nor UO_507 (O_507,N_4554,N_4049);
and UO_508 (O_508,N_4720,N_4055);
and UO_509 (O_509,N_4994,N_4922);
nand UO_510 (O_510,N_4366,N_4969);
or UO_511 (O_511,N_4322,N_4226);
and UO_512 (O_512,N_4064,N_4151);
or UO_513 (O_513,N_4483,N_4777);
nand UO_514 (O_514,N_4029,N_4948);
and UO_515 (O_515,N_4470,N_4589);
or UO_516 (O_516,N_4046,N_4997);
or UO_517 (O_517,N_4039,N_4155);
and UO_518 (O_518,N_4016,N_4291);
nor UO_519 (O_519,N_4706,N_4694);
nor UO_520 (O_520,N_4652,N_4889);
nor UO_521 (O_521,N_4496,N_4890);
or UO_522 (O_522,N_4506,N_4789);
nand UO_523 (O_523,N_4149,N_4391);
and UO_524 (O_524,N_4423,N_4575);
nor UO_525 (O_525,N_4128,N_4926);
nor UO_526 (O_526,N_4390,N_4292);
or UO_527 (O_527,N_4071,N_4377);
nor UO_528 (O_528,N_4074,N_4066);
nor UO_529 (O_529,N_4496,N_4313);
nand UO_530 (O_530,N_4535,N_4372);
and UO_531 (O_531,N_4267,N_4186);
or UO_532 (O_532,N_4164,N_4994);
nand UO_533 (O_533,N_4654,N_4596);
nand UO_534 (O_534,N_4458,N_4702);
or UO_535 (O_535,N_4673,N_4515);
nor UO_536 (O_536,N_4752,N_4859);
nand UO_537 (O_537,N_4000,N_4499);
nand UO_538 (O_538,N_4127,N_4910);
nand UO_539 (O_539,N_4098,N_4163);
nor UO_540 (O_540,N_4821,N_4724);
nor UO_541 (O_541,N_4644,N_4882);
and UO_542 (O_542,N_4712,N_4053);
nand UO_543 (O_543,N_4905,N_4782);
or UO_544 (O_544,N_4877,N_4648);
nand UO_545 (O_545,N_4447,N_4085);
and UO_546 (O_546,N_4157,N_4355);
nand UO_547 (O_547,N_4542,N_4765);
nand UO_548 (O_548,N_4837,N_4513);
nand UO_549 (O_549,N_4113,N_4792);
nor UO_550 (O_550,N_4189,N_4624);
nand UO_551 (O_551,N_4091,N_4830);
and UO_552 (O_552,N_4641,N_4873);
nand UO_553 (O_553,N_4349,N_4573);
nor UO_554 (O_554,N_4191,N_4372);
nor UO_555 (O_555,N_4547,N_4994);
nor UO_556 (O_556,N_4950,N_4422);
nor UO_557 (O_557,N_4238,N_4184);
nor UO_558 (O_558,N_4871,N_4149);
nor UO_559 (O_559,N_4233,N_4681);
or UO_560 (O_560,N_4630,N_4773);
and UO_561 (O_561,N_4471,N_4032);
nor UO_562 (O_562,N_4811,N_4458);
nand UO_563 (O_563,N_4452,N_4347);
or UO_564 (O_564,N_4288,N_4625);
and UO_565 (O_565,N_4613,N_4023);
and UO_566 (O_566,N_4636,N_4571);
nor UO_567 (O_567,N_4015,N_4566);
or UO_568 (O_568,N_4369,N_4679);
nand UO_569 (O_569,N_4813,N_4561);
nor UO_570 (O_570,N_4410,N_4834);
and UO_571 (O_571,N_4017,N_4829);
nand UO_572 (O_572,N_4679,N_4900);
or UO_573 (O_573,N_4673,N_4173);
nand UO_574 (O_574,N_4878,N_4835);
or UO_575 (O_575,N_4354,N_4833);
or UO_576 (O_576,N_4003,N_4929);
nand UO_577 (O_577,N_4606,N_4381);
or UO_578 (O_578,N_4427,N_4945);
or UO_579 (O_579,N_4469,N_4895);
nand UO_580 (O_580,N_4069,N_4426);
nand UO_581 (O_581,N_4643,N_4569);
nand UO_582 (O_582,N_4043,N_4965);
nor UO_583 (O_583,N_4094,N_4203);
and UO_584 (O_584,N_4290,N_4576);
nor UO_585 (O_585,N_4140,N_4438);
or UO_586 (O_586,N_4381,N_4546);
and UO_587 (O_587,N_4727,N_4011);
and UO_588 (O_588,N_4183,N_4025);
and UO_589 (O_589,N_4861,N_4933);
nand UO_590 (O_590,N_4960,N_4489);
nand UO_591 (O_591,N_4710,N_4159);
nand UO_592 (O_592,N_4429,N_4089);
or UO_593 (O_593,N_4699,N_4207);
nand UO_594 (O_594,N_4484,N_4669);
and UO_595 (O_595,N_4518,N_4885);
nor UO_596 (O_596,N_4664,N_4151);
or UO_597 (O_597,N_4075,N_4808);
nand UO_598 (O_598,N_4177,N_4005);
nand UO_599 (O_599,N_4362,N_4391);
xor UO_600 (O_600,N_4153,N_4595);
and UO_601 (O_601,N_4140,N_4754);
or UO_602 (O_602,N_4718,N_4486);
nand UO_603 (O_603,N_4293,N_4610);
or UO_604 (O_604,N_4675,N_4707);
nor UO_605 (O_605,N_4294,N_4151);
and UO_606 (O_606,N_4091,N_4408);
nor UO_607 (O_607,N_4296,N_4272);
nor UO_608 (O_608,N_4516,N_4160);
or UO_609 (O_609,N_4987,N_4497);
and UO_610 (O_610,N_4638,N_4773);
nand UO_611 (O_611,N_4734,N_4883);
nor UO_612 (O_612,N_4975,N_4239);
nand UO_613 (O_613,N_4177,N_4047);
nor UO_614 (O_614,N_4002,N_4224);
nor UO_615 (O_615,N_4816,N_4634);
and UO_616 (O_616,N_4155,N_4243);
nor UO_617 (O_617,N_4436,N_4935);
nand UO_618 (O_618,N_4205,N_4574);
nand UO_619 (O_619,N_4524,N_4971);
nand UO_620 (O_620,N_4075,N_4235);
nand UO_621 (O_621,N_4727,N_4295);
and UO_622 (O_622,N_4491,N_4319);
or UO_623 (O_623,N_4488,N_4598);
nand UO_624 (O_624,N_4756,N_4005);
or UO_625 (O_625,N_4634,N_4680);
or UO_626 (O_626,N_4680,N_4545);
nand UO_627 (O_627,N_4776,N_4970);
or UO_628 (O_628,N_4826,N_4852);
and UO_629 (O_629,N_4207,N_4687);
and UO_630 (O_630,N_4700,N_4234);
or UO_631 (O_631,N_4969,N_4927);
or UO_632 (O_632,N_4006,N_4026);
and UO_633 (O_633,N_4479,N_4828);
and UO_634 (O_634,N_4189,N_4522);
and UO_635 (O_635,N_4247,N_4311);
or UO_636 (O_636,N_4796,N_4228);
and UO_637 (O_637,N_4574,N_4461);
xor UO_638 (O_638,N_4527,N_4418);
and UO_639 (O_639,N_4119,N_4104);
nor UO_640 (O_640,N_4598,N_4092);
xnor UO_641 (O_641,N_4646,N_4085);
or UO_642 (O_642,N_4623,N_4879);
nor UO_643 (O_643,N_4481,N_4032);
and UO_644 (O_644,N_4598,N_4571);
or UO_645 (O_645,N_4552,N_4351);
nand UO_646 (O_646,N_4680,N_4757);
or UO_647 (O_647,N_4456,N_4323);
nor UO_648 (O_648,N_4579,N_4496);
or UO_649 (O_649,N_4655,N_4398);
or UO_650 (O_650,N_4490,N_4540);
nand UO_651 (O_651,N_4065,N_4446);
nor UO_652 (O_652,N_4074,N_4936);
nand UO_653 (O_653,N_4611,N_4566);
nand UO_654 (O_654,N_4443,N_4810);
and UO_655 (O_655,N_4406,N_4277);
or UO_656 (O_656,N_4688,N_4010);
nor UO_657 (O_657,N_4553,N_4150);
nor UO_658 (O_658,N_4482,N_4819);
and UO_659 (O_659,N_4023,N_4655);
nor UO_660 (O_660,N_4148,N_4423);
or UO_661 (O_661,N_4549,N_4642);
and UO_662 (O_662,N_4492,N_4240);
nand UO_663 (O_663,N_4984,N_4174);
nand UO_664 (O_664,N_4003,N_4110);
and UO_665 (O_665,N_4530,N_4085);
nor UO_666 (O_666,N_4419,N_4121);
and UO_667 (O_667,N_4495,N_4749);
nor UO_668 (O_668,N_4663,N_4841);
nand UO_669 (O_669,N_4457,N_4423);
and UO_670 (O_670,N_4895,N_4099);
nand UO_671 (O_671,N_4705,N_4307);
nor UO_672 (O_672,N_4523,N_4932);
and UO_673 (O_673,N_4569,N_4965);
and UO_674 (O_674,N_4356,N_4568);
nor UO_675 (O_675,N_4412,N_4500);
or UO_676 (O_676,N_4201,N_4732);
nor UO_677 (O_677,N_4953,N_4749);
nor UO_678 (O_678,N_4647,N_4868);
or UO_679 (O_679,N_4056,N_4184);
or UO_680 (O_680,N_4521,N_4692);
nand UO_681 (O_681,N_4538,N_4610);
and UO_682 (O_682,N_4351,N_4027);
and UO_683 (O_683,N_4114,N_4038);
and UO_684 (O_684,N_4760,N_4905);
and UO_685 (O_685,N_4180,N_4370);
and UO_686 (O_686,N_4278,N_4804);
and UO_687 (O_687,N_4890,N_4125);
or UO_688 (O_688,N_4292,N_4895);
nor UO_689 (O_689,N_4629,N_4853);
and UO_690 (O_690,N_4028,N_4987);
nor UO_691 (O_691,N_4239,N_4424);
and UO_692 (O_692,N_4696,N_4084);
and UO_693 (O_693,N_4711,N_4756);
or UO_694 (O_694,N_4464,N_4087);
and UO_695 (O_695,N_4536,N_4492);
and UO_696 (O_696,N_4577,N_4197);
or UO_697 (O_697,N_4074,N_4807);
or UO_698 (O_698,N_4117,N_4109);
nor UO_699 (O_699,N_4365,N_4123);
nor UO_700 (O_700,N_4228,N_4807);
or UO_701 (O_701,N_4822,N_4807);
or UO_702 (O_702,N_4199,N_4554);
nor UO_703 (O_703,N_4768,N_4281);
nor UO_704 (O_704,N_4981,N_4855);
and UO_705 (O_705,N_4310,N_4912);
nor UO_706 (O_706,N_4329,N_4612);
nand UO_707 (O_707,N_4539,N_4004);
or UO_708 (O_708,N_4923,N_4115);
and UO_709 (O_709,N_4030,N_4900);
or UO_710 (O_710,N_4960,N_4748);
and UO_711 (O_711,N_4124,N_4864);
and UO_712 (O_712,N_4677,N_4340);
nor UO_713 (O_713,N_4532,N_4916);
nand UO_714 (O_714,N_4017,N_4096);
nor UO_715 (O_715,N_4000,N_4068);
or UO_716 (O_716,N_4842,N_4746);
or UO_717 (O_717,N_4526,N_4178);
nand UO_718 (O_718,N_4585,N_4257);
and UO_719 (O_719,N_4618,N_4908);
nor UO_720 (O_720,N_4094,N_4338);
and UO_721 (O_721,N_4969,N_4210);
and UO_722 (O_722,N_4245,N_4539);
or UO_723 (O_723,N_4775,N_4644);
and UO_724 (O_724,N_4235,N_4946);
nor UO_725 (O_725,N_4661,N_4525);
and UO_726 (O_726,N_4571,N_4435);
nor UO_727 (O_727,N_4437,N_4050);
nor UO_728 (O_728,N_4587,N_4169);
nor UO_729 (O_729,N_4597,N_4058);
nor UO_730 (O_730,N_4981,N_4324);
nand UO_731 (O_731,N_4156,N_4891);
and UO_732 (O_732,N_4607,N_4065);
and UO_733 (O_733,N_4649,N_4089);
or UO_734 (O_734,N_4263,N_4406);
nor UO_735 (O_735,N_4553,N_4960);
and UO_736 (O_736,N_4994,N_4863);
nor UO_737 (O_737,N_4012,N_4133);
or UO_738 (O_738,N_4996,N_4257);
nand UO_739 (O_739,N_4102,N_4530);
or UO_740 (O_740,N_4284,N_4596);
or UO_741 (O_741,N_4836,N_4531);
or UO_742 (O_742,N_4245,N_4104);
or UO_743 (O_743,N_4787,N_4709);
nor UO_744 (O_744,N_4535,N_4119);
or UO_745 (O_745,N_4090,N_4171);
nor UO_746 (O_746,N_4671,N_4316);
nor UO_747 (O_747,N_4873,N_4524);
and UO_748 (O_748,N_4159,N_4023);
or UO_749 (O_749,N_4656,N_4588);
or UO_750 (O_750,N_4854,N_4157);
or UO_751 (O_751,N_4302,N_4713);
and UO_752 (O_752,N_4797,N_4285);
and UO_753 (O_753,N_4095,N_4443);
nand UO_754 (O_754,N_4485,N_4895);
and UO_755 (O_755,N_4823,N_4792);
and UO_756 (O_756,N_4432,N_4494);
nor UO_757 (O_757,N_4588,N_4745);
and UO_758 (O_758,N_4877,N_4660);
nor UO_759 (O_759,N_4043,N_4142);
nor UO_760 (O_760,N_4263,N_4044);
nor UO_761 (O_761,N_4833,N_4832);
nor UO_762 (O_762,N_4710,N_4838);
or UO_763 (O_763,N_4341,N_4464);
and UO_764 (O_764,N_4419,N_4219);
nand UO_765 (O_765,N_4357,N_4823);
nand UO_766 (O_766,N_4503,N_4827);
or UO_767 (O_767,N_4447,N_4937);
or UO_768 (O_768,N_4563,N_4775);
nand UO_769 (O_769,N_4931,N_4157);
nand UO_770 (O_770,N_4586,N_4706);
or UO_771 (O_771,N_4847,N_4197);
and UO_772 (O_772,N_4553,N_4747);
nand UO_773 (O_773,N_4629,N_4991);
nor UO_774 (O_774,N_4109,N_4523);
nor UO_775 (O_775,N_4493,N_4434);
nand UO_776 (O_776,N_4091,N_4201);
nand UO_777 (O_777,N_4276,N_4109);
or UO_778 (O_778,N_4303,N_4115);
or UO_779 (O_779,N_4059,N_4330);
or UO_780 (O_780,N_4753,N_4869);
and UO_781 (O_781,N_4259,N_4300);
nand UO_782 (O_782,N_4365,N_4921);
or UO_783 (O_783,N_4534,N_4725);
and UO_784 (O_784,N_4209,N_4141);
nand UO_785 (O_785,N_4711,N_4088);
nor UO_786 (O_786,N_4754,N_4311);
or UO_787 (O_787,N_4898,N_4347);
or UO_788 (O_788,N_4206,N_4456);
and UO_789 (O_789,N_4398,N_4934);
or UO_790 (O_790,N_4437,N_4799);
or UO_791 (O_791,N_4112,N_4449);
nor UO_792 (O_792,N_4413,N_4948);
nor UO_793 (O_793,N_4738,N_4070);
and UO_794 (O_794,N_4886,N_4584);
and UO_795 (O_795,N_4814,N_4013);
nand UO_796 (O_796,N_4282,N_4169);
xnor UO_797 (O_797,N_4256,N_4843);
and UO_798 (O_798,N_4278,N_4415);
and UO_799 (O_799,N_4976,N_4206);
and UO_800 (O_800,N_4453,N_4590);
or UO_801 (O_801,N_4538,N_4256);
nor UO_802 (O_802,N_4196,N_4114);
and UO_803 (O_803,N_4154,N_4935);
nand UO_804 (O_804,N_4318,N_4067);
or UO_805 (O_805,N_4952,N_4334);
and UO_806 (O_806,N_4049,N_4251);
nor UO_807 (O_807,N_4610,N_4866);
and UO_808 (O_808,N_4597,N_4135);
or UO_809 (O_809,N_4345,N_4355);
nor UO_810 (O_810,N_4574,N_4328);
and UO_811 (O_811,N_4313,N_4651);
and UO_812 (O_812,N_4091,N_4387);
nand UO_813 (O_813,N_4412,N_4326);
or UO_814 (O_814,N_4615,N_4458);
nor UO_815 (O_815,N_4631,N_4100);
and UO_816 (O_816,N_4361,N_4445);
nand UO_817 (O_817,N_4403,N_4704);
nor UO_818 (O_818,N_4142,N_4002);
and UO_819 (O_819,N_4588,N_4551);
nor UO_820 (O_820,N_4430,N_4226);
nor UO_821 (O_821,N_4342,N_4677);
and UO_822 (O_822,N_4261,N_4065);
nand UO_823 (O_823,N_4713,N_4179);
nor UO_824 (O_824,N_4253,N_4110);
nor UO_825 (O_825,N_4028,N_4936);
nand UO_826 (O_826,N_4014,N_4145);
or UO_827 (O_827,N_4199,N_4642);
nand UO_828 (O_828,N_4276,N_4760);
nand UO_829 (O_829,N_4682,N_4438);
and UO_830 (O_830,N_4770,N_4390);
and UO_831 (O_831,N_4797,N_4614);
nand UO_832 (O_832,N_4836,N_4891);
or UO_833 (O_833,N_4126,N_4423);
nand UO_834 (O_834,N_4032,N_4075);
or UO_835 (O_835,N_4516,N_4523);
or UO_836 (O_836,N_4283,N_4961);
and UO_837 (O_837,N_4136,N_4392);
and UO_838 (O_838,N_4866,N_4678);
nand UO_839 (O_839,N_4183,N_4244);
and UO_840 (O_840,N_4078,N_4903);
nand UO_841 (O_841,N_4168,N_4652);
and UO_842 (O_842,N_4409,N_4254);
or UO_843 (O_843,N_4101,N_4650);
and UO_844 (O_844,N_4727,N_4761);
and UO_845 (O_845,N_4499,N_4793);
xor UO_846 (O_846,N_4279,N_4774);
nor UO_847 (O_847,N_4711,N_4011);
and UO_848 (O_848,N_4207,N_4887);
nor UO_849 (O_849,N_4027,N_4083);
nand UO_850 (O_850,N_4561,N_4521);
and UO_851 (O_851,N_4316,N_4928);
nand UO_852 (O_852,N_4507,N_4161);
nor UO_853 (O_853,N_4788,N_4025);
nand UO_854 (O_854,N_4274,N_4048);
nand UO_855 (O_855,N_4058,N_4047);
or UO_856 (O_856,N_4217,N_4525);
nor UO_857 (O_857,N_4530,N_4880);
or UO_858 (O_858,N_4716,N_4566);
or UO_859 (O_859,N_4891,N_4909);
and UO_860 (O_860,N_4499,N_4700);
nor UO_861 (O_861,N_4189,N_4947);
nand UO_862 (O_862,N_4036,N_4646);
or UO_863 (O_863,N_4727,N_4452);
and UO_864 (O_864,N_4344,N_4993);
nor UO_865 (O_865,N_4090,N_4118);
nand UO_866 (O_866,N_4202,N_4937);
nor UO_867 (O_867,N_4074,N_4049);
or UO_868 (O_868,N_4095,N_4981);
and UO_869 (O_869,N_4397,N_4745);
nand UO_870 (O_870,N_4145,N_4112);
nand UO_871 (O_871,N_4902,N_4773);
nor UO_872 (O_872,N_4957,N_4124);
nor UO_873 (O_873,N_4694,N_4593);
xnor UO_874 (O_874,N_4107,N_4859);
or UO_875 (O_875,N_4048,N_4334);
nor UO_876 (O_876,N_4885,N_4829);
or UO_877 (O_877,N_4816,N_4348);
nand UO_878 (O_878,N_4428,N_4634);
nor UO_879 (O_879,N_4923,N_4038);
nand UO_880 (O_880,N_4889,N_4609);
or UO_881 (O_881,N_4994,N_4025);
and UO_882 (O_882,N_4466,N_4086);
or UO_883 (O_883,N_4528,N_4055);
nand UO_884 (O_884,N_4996,N_4849);
nand UO_885 (O_885,N_4564,N_4092);
or UO_886 (O_886,N_4174,N_4959);
and UO_887 (O_887,N_4479,N_4812);
nand UO_888 (O_888,N_4119,N_4339);
and UO_889 (O_889,N_4689,N_4957);
nor UO_890 (O_890,N_4626,N_4185);
and UO_891 (O_891,N_4585,N_4984);
nand UO_892 (O_892,N_4440,N_4249);
and UO_893 (O_893,N_4988,N_4546);
and UO_894 (O_894,N_4436,N_4526);
nor UO_895 (O_895,N_4419,N_4964);
nor UO_896 (O_896,N_4934,N_4222);
nor UO_897 (O_897,N_4157,N_4908);
nand UO_898 (O_898,N_4806,N_4521);
nor UO_899 (O_899,N_4567,N_4049);
nor UO_900 (O_900,N_4139,N_4573);
nand UO_901 (O_901,N_4352,N_4581);
and UO_902 (O_902,N_4175,N_4430);
nor UO_903 (O_903,N_4327,N_4676);
nor UO_904 (O_904,N_4311,N_4159);
nor UO_905 (O_905,N_4367,N_4433);
or UO_906 (O_906,N_4865,N_4193);
xnor UO_907 (O_907,N_4482,N_4634);
or UO_908 (O_908,N_4022,N_4259);
or UO_909 (O_909,N_4231,N_4015);
and UO_910 (O_910,N_4468,N_4357);
and UO_911 (O_911,N_4725,N_4256);
nand UO_912 (O_912,N_4402,N_4319);
or UO_913 (O_913,N_4503,N_4493);
nor UO_914 (O_914,N_4801,N_4459);
nand UO_915 (O_915,N_4405,N_4062);
and UO_916 (O_916,N_4770,N_4319);
and UO_917 (O_917,N_4821,N_4953);
and UO_918 (O_918,N_4784,N_4467);
nand UO_919 (O_919,N_4773,N_4169);
nand UO_920 (O_920,N_4636,N_4154);
or UO_921 (O_921,N_4547,N_4020);
and UO_922 (O_922,N_4031,N_4685);
nor UO_923 (O_923,N_4841,N_4876);
and UO_924 (O_924,N_4629,N_4278);
nor UO_925 (O_925,N_4967,N_4880);
or UO_926 (O_926,N_4552,N_4095);
and UO_927 (O_927,N_4987,N_4083);
nor UO_928 (O_928,N_4342,N_4068);
nor UO_929 (O_929,N_4291,N_4855);
nor UO_930 (O_930,N_4959,N_4515);
or UO_931 (O_931,N_4428,N_4377);
nand UO_932 (O_932,N_4714,N_4552);
nand UO_933 (O_933,N_4232,N_4824);
nand UO_934 (O_934,N_4381,N_4648);
and UO_935 (O_935,N_4965,N_4600);
and UO_936 (O_936,N_4301,N_4519);
and UO_937 (O_937,N_4223,N_4150);
or UO_938 (O_938,N_4840,N_4072);
nor UO_939 (O_939,N_4564,N_4928);
and UO_940 (O_940,N_4175,N_4080);
nand UO_941 (O_941,N_4968,N_4550);
or UO_942 (O_942,N_4080,N_4253);
nand UO_943 (O_943,N_4996,N_4294);
nor UO_944 (O_944,N_4508,N_4931);
or UO_945 (O_945,N_4454,N_4947);
and UO_946 (O_946,N_4295,N_4953);
nor UO_947 (O_947,N_4187,N_4870);
nand UO_948 (O_948,N_4352,N_4656);
nor UO_949 (O_949,N_4441,N_4686);
and UO_950 (O_950,N_4970,N_4123);
and UO_951 (O_951,N_4934,N_4141);
nor UO_952 (O_952,N_4971,N_4892);
or UO_953 (O_953,N_4063,N_4529);
nor UO_954 (O_954,N_4994,N_4717);
and UO_955 (O_955,N_4685,N_4563);
or UO_956 (O_956,N_4860,N_4054);
and UO_957 (O_957,N_4123,N_4105);
nor UO_958 (O_958,N_4325,N_4573);
and UO_959 (O_959,N_4202,N_4300);
nand UO_960 (O_960,N_4995,N_4465);
nor UO_961 (O_961,N_4437,N_4342);
and UO_962 (O_962,N_4958,N_4214);
nor UO_963 (O_963,N_4106,N_4555);
and UO_964 (O_964,N_4328,N_4350);
nand UO_965 (O_965,N_4991,N_4392);
nor UO_966 (O_966,N_4365,N_4496);
nand UO_967 (O_967,N_4403,N_4578);
nor UO_968 (O_968,N_4194,N_4396);
or UO_969 (O_969,N_4321,N_4943);
nor UO_970 (O_970,N_4970,N_4688);
or UO_971 (O_971,N_4522,N_4541);
xor UO_972 (O_972,N_4370,N_4545);
or UO_973 (O_973,N_4656,N_4329);
nand UO_974 (O_974,N_4113,N_4482);
or UO_975 (O_975,N_4146,N_4504);
and UO_976 (O_976,N_4273,N_4972);
or UO_977 (O_977,N_4924,N_4022);
and UO_978 (O_978,N_4185,N_4216);
nor UO_979 (O_979,N_4154,N_4006);
nor UO_980 (O_980,N_4818,N_4492);
and UO_981 (O_981,N_4474,N_4248);
or UO_982 (O_982,N_4726,N_4761);
and UO_983 (O_983,N_4889,N_4776);
nand UO_984 (O_984,N_4673,N_4885);
xnor UO_985 (O_985,N_4220,N_4710);
nor UO_986 (O_986,N_4420,N_4800);
nor UO_987 (O_987,N_4659,N_4611);
nor UO_988 (O_988,N_4301,N_4130);
nand UO_989 (O_989,N_4250,N_4372);
or UO_990 (O_990,N_4745,N_4008);
nand UO_991 (O_991,N_4145,N_4030);
nand UO_992 (O_992,N_4042,N_4860);
nor UO_993 (O_993,N_4728,N_4541);
and UO_994 (O_994,N_4501,N_4059);
nor UO_995 (O_995,N_4984,N_4751);
and UO_996 (O_996,N_4914,N_4490);
nand UO_997 (O_997,N_4791,N_4985);
nand UO_998 (O_998,N_4755,N_4072);
nand UO_999 (O_999,N_4412,N_4985);
endmodule